// Benchmark "top" written by ABC on Fri Jun 21 17:49:24 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n141_, new_new_n142_, new_new_n143_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1033_, new_new_n1034_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  OR4        g0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g0067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  NO2        g0068(.A(new_new_n89_), .B(new_new_n90_), .Y(new_new_n91_));
  OAI210     g0069(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n91_), .Y(new_new_n92_));
  NAi21      g0070(.An(i_6_), .B(i_10_), .Y(new_new_n93_));
  NA2        g0071(.A(i_6_), .B(i_9_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n93_), .B0(new_new_n64_), .Y(new_new_n95_));
  NA2        g0073(.A(i_2_), .B(i_6_), .Y(new_new_n96_));
  INV        g0074(.A(new_new_n95_), .Y(new_new_n97_));
  AOI210     g0075(.A0(new_new_n97_), .A1(new_new_n92_), .B0(new_new_n81_), .Y(new_new_n98_));
  AN3        g0076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n99_));
  NAi21      g0077(.An(i_6_), .B(i_11_), .Y(new_new_n100_));
  NO2        g0078(.A(i_5_), .B(i_8_), .Y(new_new_n101_));
  NOi21      g0079(.An(new_new_n101_), .B(new_new_n100_), .Y(new_new_n102_));
  AOI220     g0080(.A0(new_new_n102_), .A1(new_new_n63_), .B0(new_new_n99_), .B1(new_new_n32_), .Y(new_new_n103_));
  INV        g0081(.A(i_7_), .Y(new_new_n104_));
  NA2        g0082(.A(new_new_n47_), .B(new_new_n104_), .Y(new_new_n105_));
  NO2        g0083(.A(i_0_), .B(i_5_), .Y(new_new_n106_));
  NO2        g0084(.A(new_new_n106_), .B(new_new_n87_), .Y(new_new_n107_));
  NA2        g0085(.A(i_12_), .B(i_3_), .Y(new_new_n108_));
  INV        g0086(.A(new_new_n108_), .Y(new_new_n109_));
  NA3        g0087(.A(new_new_n109_), .B(new_new_n107_), .C(new_new_n105_), .Y(new_new_n110_));
  NAi21      g0088(.An(i_7_), .B(i_11_), .Y(new_new_n111_));
  NO3        g0089(.A(new_new_n111_), .B(new_new_n93_), .C(new_new_n54_), .Y(new_new_n112_));
  AN2        g0090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g0091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g0092(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n115_));
  NO2        g0093(.A(i_8_), .B(new_new_n104_), .Y(new_new_n116_));
  NO3        g0094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g0095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g0097(.A(i_11_), .B(i_12_), .Y(new_new_n120_));
  INV        g0098(.A(new_new_n120_), .Y(new_new_n121_));
  NO2        g0099(.A(new_new_n121_), .B(new_new_n117_), .Y(new_new_n122_));
  NAi41      g0100(.An(new_new_n112_), .B(new_new_n122_), .C(new_new_n110_), .D(new_new_n103_), .Y(new_new_n123_));
  NOi21      g0101(.An(i_1_), .B(i_5_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(i_11_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n126_));
  NA2        g0104(.A(i_7_), .B(new_new_n25_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n127_), .B(new_new_n126_), .Y(new_new_n128_));
  NO2        g0106(.A(new_new_n128_), .B(new_new_n47_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n94_), .B(new_new_n93_), .Y(new_new_n130_));
  NAi21      g0108(.An(i_3_), .B(i_8_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n131_), .B(new_new_n63_), .Y(new_new_n132_));
  NOi31      g0110(.An(new_new_n132_), .B(new_new_n130_), .C(new_new_n129_), .Y(new_new_n133_));
  NO2        g0111(.A(i_1_), .B(new_new_n87_), .Y(new_new_n134_));
  NO2        g0112(.A(i_6_), .B(i_5_), .Y(new_new_n135_));
  NA2        g0113(.A(new_new_n135_), .B(i_3_), .Y(new_new_n136_));
  AO210      g0114(.A0(new_new_n136_), .A1(new_new_n48_), .B0(new_new_n134_), .Y(new_new_n137_));
  OAI220     g0115(.A0(new_new_n137_), .A1(new_new_n111_), .B0(new_new_n133_), .B1(new_new_n125_), .Y(new_new_n138_));
  NO3        g0116(.A(new_new_n138_), .B(new_new_n123_), .C(new_new_n98_), .Y(new_new_n139_));
  NA3        g0117(.A(new_new_n139_), .B(new_new_n80_), .C(new_new_n57_), .Y(mai2));
  NO2        g0118(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n141_));
  NA2        g0119(.A(i_6_), .B(new_new_n25_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(new_new_n141_), .Y(new_new_n143_));
  NA4        g0121(.A(new_new_n143_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(mai0));
  AN2        g0122(.A(i_8_), .B(i_7_), .Y(new_new_n145_));
  NA2        g0123(.A(new_new_n145_), .B(i_6_), .Y(new_new_n146_));
  NO2        g0124(.A(i_12_), .B(i_13_), .Y(new_new_n147_));
  NAi21      g0125(.An(i_5_), .B(i_11_), .Y(new_new_n148_));
  NOi21      g0126(.An(new_new_n147_), .B(new_new_n148_), .Y(new_new_n149_));
  NO2        g0127(.A(i_0_), .B(i_1_), .Y(new_new_n150_));
  NA2        g0128(.A(i_2_), .B(i_3_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(i_4_), .Y(new_new_n152_));
  NA3        g0130(.A(new_new_n152_), .B(new_new_n150_), .C(new_new_n149_), .Y(new_new_n153_));
  AN2        g0131(.A(new_new_n147_), .B(new_new_n84_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n154_), .B(new_new_n27_), .Y(new_new_n155_));
  NA2        g0133(.A(i_1_), .B(i_5_), .Y(new_new_n156_));
  NO2        g0134(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n157_));
  NA2        g0135(.A(new_new_n157_), .B(new_new_n36_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n156_), .C(new_new_n155_), .Y(new_new_n159_));
  OR2        g0137(.A(i_0_), .B(i_1_), .Y(new_new_n160_));
  NO3        g0138(.A(new_new_n160_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n161_));
  NAi32      g0139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n162_));
  NAi21      g0140(.An(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  NOi21      g0141(.An(i_4_), .B(i_10_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n40_), .Y(new_new_n165_));
  NO2        g0143(.A(i_3_), .B(i_5_), .Y(new_new_n166_));
  NO3        g0144(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n167_));
  NA2        g0145(.A(new_new_n167_), .B(new_new_n166_), .Y(new_new_n168_));
  OAI210     g0146(.A0(new_new_n168_), .A1(new_new_n165_), .B0(new_new_n163_), .Y(new_new_n169_));
  NO2        g0147(.A(new_new_n169_), .B(new_new_n159_), .Y(new_new_n170_));
  AOI210     g0148(.A0(new_new_n170_), .A1(new_new_n153_), .B0(new_new_n146_), .Y(new_new_n171_));
  NA3        g0149(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n172_));
  NA2        g0150(.A(i_3_), .B(new_new_n49_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_4_), .B(i_9_), .Y(new_new_n174_));
  NOi21      g0152(.An(i_11_), .B(i_13_), .Y(new_new_n175_));
  NA2        g0153(.A(new_new_n175_), .B(new_new_n174_), .Y(new_new_n176_));
  OR2        g0154(.A(new_new_n176_), .B(new_new_n173_), .Y(new_new_n177_));
  NO2        g0155(.A(i_4_), .B(i_5_), .Y(new_new_n178_));
  NAi21      g0156(.An(i_12_), .B(i_11_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n179_), .B(i_13_), .Y(new_new_n180_));
  NA3        g0158(.A(new_new_n180_), .B(new_new_n178_), .C(new_new_n84_), .Y(new_new_n181_));
  AOI210     g0159(.A0(new_new_n181_), .A1(new_new_n177_), .B0(new_new_n172_), .Y(new_new_n182_));
  NO2        g0160(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n183_));
  INV        g0161(.A(new_new_n183_), .Y(new_new_n184_));
  NA2        g0162(.A(new_new_n36_), .B(i_5_), .Y(new_new_n185_));
  NAi31      g0163(.An(new_new_n185_), .B(new_new_n154_), .C(i_11_), .Y(new_new_n186_));
  NA2        g0164(.A(i_3_), .B(i_5_), .Y(new_new_n187_));
  OR2        g0165(.A(new_new_n187_), .B(new_new_n176_), .Y(new_new_n188_));
  AOI210     g0166(.A0(new_new_n188_), .A1(new_new_n186_), .B0(new_new_n184_), .Y(new_new_n189_));
  NO2        g0167(.A(new_new_n74_), .B(i_5_), .Y(new_new_n190_));
  NO2        g0168(.A(i_13_), .B(i_10_), .Y(new_new_n191_));
  NA3        g0169(.A(new_new_n191_), .B(new_new_n190_), .C(new_new_n45_), .Y(new_new_n192_));
  NO2        g0170(.A(i_2_), .B(i_1_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_3_), .Y(new_new_n194_));
  NAi21      g0172(.An(i_4_), .B(i_12_), .Y(new_new_n195_));
  NO3        g0173(.A(new_new_n194_), .B(new_new_n192_), .C(new_new_n25_), .Y(new_new_n196_));
  NO3        g0174(.A(new_new_n196_), .B(new_new_n189_), .C(new_new_n182_), .Y(new_new_n197_));
  INV        g0175(.A(i_8_), .Y(new_new_n198_));
  NO2        g0176(.A(new_new_n198_), .B(i_7_), .Y(new_new_n199_));
  NA2        g0177(.A(new_new_n199_), .B(i_6_), .Y(new_new_n200_));
  NO3        g0178(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n201_));
  NA2        g0179(.A(new_new_n201_), .B(new_new_n116_), .Y(new_new_n202_));
  NO3        g0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n203_));
  NA3        g0181(.A(new_new_n203_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n204_));
  NO3        g0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n205_));
  OAI210     g0183(.A0(new_new_n99_), .A1(i_12_), .B0(new_new_n205_), .Y(new_new_n206_));
  AOI210     g0184(.A0(new_new_n206_), .A1(new_new_n204_), .B0(new_new_n202_), .Y(new_new_n207_));
  NO2        g0185(.A(i_3_), .B(i_8_), .Y(new_new_n208_));
  NO3        g0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n209_));
  NO2        g0187(.A(new_new_n106_), .B(new_new_n59_), .Y(new_new_n210_));
  NO2        g0188(.A(i_13_), .B(i_9_), .Y(new_new_n211_));
  NA3        g0189(.A(new_new_n211_), .B(i_6_), .C(new_new_n198_), .Y(new_new_n212_));
  NAi21      g0190(.An(i_12_), .B(i_3_), .Y(new_new_n213_));
  OR2        g0191(.A(new_new_n213_), .B(new_new_n212_), .Y(new_new_n214_));
  NO2        g0192(.A(new_new_n45_), .B(i_5_), .Y(new_new_n215_));
  NO3        g0193(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n216_));
  NA2        g0194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n217_), .B(new_new_n214_), .Y(new_new_n218_));
  NO2        g0196(.A(new_new_n218_), .B(new_new_n207_), .Y(new_new_n219_));
  OAI220     g0197(.A0(new_new_n219_), .A1(i_4_), .B0(new_new_n200_), .B1(new_new_n197_), .Y(new_new_n220_));
  NAi21      g0198(.An(i_12_), .B(i_7_), .Y(new_new_n221_));
  NA3        g0199(.A(i_13_), .B(new_new_n198_), .C(i_10_), .Y(new_new_n222_));
  NA2        g0200(.A(i_0_), .B(i_5_), .Y(new_new_n223_));
  NAi31      g0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n225_));
  INV        g0203(.A(i_13_), .Y(new_new_n226_));
  NO2        g0204(.A(i_12_), .B(new_new_n226_), .Y(new_new_n227_));
  NO2        g0205(.A(i_12_), .B(new_new_n37_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n187_), .B(i_4_), .Y(new_new_n229_));
  NA2        g0207(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n230_));
  OR2        g0208(.A(i_8_), .B(i_7_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n231_), .B(new_new_n87_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n54_), .B(i_1_), .Y(new_new_n233_));
  NA2        g0211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  INV        g0212(.A(i_12_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n45_), .B(new_new_n235_), .Y(new_new_n236_));
  NO3        g0214(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n237_));
  NA2        g0215(.A(i_2_), .B(i_1_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n234_), .B(new_new_n230_), .Y(new_new_n239_));
  NO3        g0217(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n240_));
  NAi21      g0218(.An(i_4_), .B(i_3_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n241_), .B(new_new_n76_), .Y(new_new_n242_));
  NO2        g0220(.A(i_0_), .B(i_6_), .Y(new_new_n243_));
  NOi41      g0221(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n244_));
  NA2        g0222(.A(new_new_n244_), .B(new_new_n243_), .Y(new_new_n245_));
  NO2        g0223(.A(new_new_n238_), .B(new_new_n187_), .Y(new_new_n246_));
  NAi21      g0224(.An(new_new_n245_), .B(new_new_n246_), .Y(new_new_n247_));
  INV        g0225(.A(new_new_n247_), .Y(new_new_n248_));
  AOI210     g0226(.A0(new_new_n248_), .A1(new_new_n40_), .B0(new_new_n239_), .Y(new_new_n249_));
  NO2        g0227(.A(i_11_), .B(new_new_n226_), .Y(new_new_n250_));
  NOi21      g0228(.An(i_1_), .B(i_6_), .Y(new_new_n251_));
  NAi21      g0229(.An(i_3_), .B(i_7_), .Y(new_new_n252_));
  NA2        g0230(.A(new_new_n235_), .B(i_9_), .Y(new_new_n253_));
  OR4        g0231(.A(new_new_n253_), .B(new_new_n252_), .C(new_new_n251_), .D(new_new_n190_), .Y(new_new_n254_));
  NO2        g0232(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n255_));
  NO2        g0233(.A(i_12_), .B(i_3_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n74_), .B(i_5_), .Y(new_new_n257_));
  NA2        g0235(.A(i_3_), .B(i_9_), .Y(new_new_n258_));
  NAi21      g0236(.An(i_7_), .B(i_10_), .Y(new_new_n259_));
  NO2        g0237(.A(new_new_n259_), .B(new_new_n258_), .Y(new_new_n260_));
  NA3        g0238(.A(new_new_n260_), .B(new_new_n257_), .C(new_new_n65_), .Y(new_new_n261_));
  NA2        g0239(.A(new_new_n261_), .B(new_new_n254_), .Y(new_new_n262_));
  NA3        g0240(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n263_));
  INV        g0241(.A(new_new_n146_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n235_), .B(i_13_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n76_), .Y(new_new_n266_));
  AOI220     g0244(.A0(new_new_n266_), .A1(new_new_n264_), .B0(new_new_n262_), .B1(new_new_n250_), .Y(new_new_n267_));
  NO2        g0245(.A(new_new_n231_), .B(new_new_n37_), .Y(new_new_n268_));
  NA2        g0246(.A(i_12_), .B(i_6_), .Y(new_new_n269_));
  OR2        g0247(.A(i_13_), .B(i_9_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n241_), .B(i_2_), .Y(new_new_n271_));
  NA2        g0249(.A(new_new_n250_), .B(i_9_), .Y(new_new_n272_));
  NA2        g0250(.A(new_new_n157_), .B(new_new_n64_), .Y(new_new_n273_));
  NO3        g0251(.A(i_11_), .B(new_new_n226_), .C(new_new_n25_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n252_), .B(i_8_), .Y(new_new_n275_));
  NO2        g0253(.A(i_6_), .B(new_new_n49_), .Y(new_new_n276_));
  NA3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n274_), .Y(new_new_n277_));
  NO3        g0255(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n278_));
  NA3        g0256(.A(new_new_n278_), .B(new_new_n268_), .C(new_new_n227_), .Y(new_new_n279_));
  AOI210     g0257(.A0(new_new_n279_), .A1(new_new_n277_), .B0(new_new_n273_), .Y(new_new_n280_));
  INV        g0258(.A(new_new_n280_), .Y(new_new_n281_));
  NA3        g0259(.A(new_new_n281_), .B(new_new_n267_), .C(new_new_n249_), .Y(new_new_n282_));
  NO3        g0260(.A(i_12_), .B(new_new_n226_), .C(new_new_n37_), .Y(new_new_n283_));
  INV        g0261(.A(new_new_n283_), .Y(new_new_n284_));
  NA2        g0262(.A(i_8_), .B(new_new_n104_), .Y(new_new_n285_));
  NOi21      g0263(.An(new_new_n166_), .B(new_new_n87_), .Y(new_new_n286_));
  NO3        g0264(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n287_));
  AOI220     g0265(.A0(new_new_n287_), .A1(new_new_n201_), .B0(new_new_n286_), .B1(new_new_n233_), .Y(new_new_n288_));
  NO2        g0266(.A(new_new_n288_), .B(new_new_n285_), .Y(new_new_n289_));
  NO2        g0267(.A(new_new_n238_), .B(i_0_), .Y(new_new_n290_));
  NA2        g0268(.A(i_0_), .B(i_1_), .Y(new_new_n291_));
  NO2        g0269(.A(new_new_n291_), .B(i_2_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n60_), .B(i_6_), .Y(new_new_n293_));
  NA3        g0271(.A(new_new_n293_), .B(new_new_n292_), .C(new_new_n166_), .Y(new_new_n294_));
  OAI210     g0272(.A0(new_new_n168_), .A1(new_new_n146_), .B0(new_new_n294_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n295_), .B(new_new_n289_), .Y(new_new_n296_));
  NO2        g0274(.A(i_3_), .B(i_10_), .Y(new_new_n297_));
  NA3        g0275(.A(new_new_n297_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n298_));
  NO2        g0276(.A(i_2_), .B(new_new_n104_), .Y(new_new_n299_));
  NA2        g0277(.A(i_1_), .B(new_new_n36_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n300_), .B(i_8_), .Y(new_new_n301_));
  NOi21      g0279(.An(new_new_n223_), .B(new_new_n106_), .Y(new_new_n302_));
  NA3        g0280(.A(new_new_n302_), .B(new_new_n301_), .C(new_new_n299_), .Y(new_new_n303_));
  AN2        g0281(.A(i_3_), .B(i_10_), .Y(new_new_n304_));
  NA4        g0282(.A(new_new_n304_), .B(new_new_n203_), .C(new_new_n180_), .D(new_new_n178_), .Y(new_new_n305_));
  NO2        g0283(.A(i_5_), .B(new_new_n37_), .Y(new_new_n306_));
  NO2        g0284(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n307_));
  OR2        g0285(.A(new_new_n303_), .B(new_new_n298_), .Y(new_new_n308_));
  OAI220     g0286(.A0(new_new_n308_), .A1(i_6_), .B0(new_new_n296_), .B1(new_new_n284_), .Y(new_new_n309_));
  NO4        g0287(.A(new_new_n309_), .B(new_new_n282_), .C(new_new_n220_), .D(new_new_n171_), .Y(new_new_n310_));
  NO3        g0288(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n311_));
  NO2        g0289(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n312_));
  NA2        g0290(.A(new_new_n290_), .B(new_new_n312_), .Y(new_new_n313_));
  NO3        g0291(.A(i_6_), .B(new_new_n198_), .C(i_7_), .Y(new_new_n314_));
  NA2        g0292(.A(new_new_n314_), .B(new_new_n203_), .Y(new_new_n315_));
  AOI210     g0293(.A0(new_new_n315_), .A1(new_new_n313_), .B0(new_new_n173_), .Y(new_new_n316_));
  NO2        g0294(.A(i_2_), .B(i_3_), .Y(new_new_n317_));
  OR2        g0295(.A(i_0_), .B(i_5_), .Y(new_new_n318_));
  NA2        g0296(.A(new_new_n223_), .B(new_new_n318_), .Y(new_new_n319_));
  NA4        g0297(.A(new_new_n319_), .B(new_new_n232_), .C(new_new_n317_), .D(i_1_), .Y(new_new_n320_));
  NA3        g0298(.A(new_new_n290_), .B(new_new_n286_), .C(new_new_n116_), .Y(new_new_n321_));
  NAi21      g0299(.An(i_8_), .B(i_7_), .Y(new_new_n322_));
  NO2        g0300(.A(new_new_n322_), .B(i_6_), .Y(new_new_n323_));
  NO2        g0301(.A(new_new_n160_), .B(new_new_n47_), .Y(new_new_n324_));
  NA3        g0302(.A(new_new_n324_), .B(new_new_n323_), .C(new_new_n166_), .Y(new_new_n325_));
  NA3        g0303(.A(new_new_n325_), .B(new_new_n321_), .C(new_new_n320_), .Y(new_new_n326_));
  OAI210     g0304(.A0(new_new_n326_), .A1(new_new_n316_), .B0(i_4_), .Y(new_new_n327_));
  NO2        g0305(.A(i_12_), .B(i_10_), .Y(new_new_n328_));
  NOi21      g0306(.An(i_5_), .B(i_0_), .Y(new_new_n329_));
  NA4        g0307(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n330_));
  NO2        g0308(.A(i_6_), .B(i_8_), .Y(new_new_n331_));
  NOi21      g0309(.An(i_0_), .B(i_2_), .Y(new_new_n332_));
  AN2        g0310(.A(new_new_n332_), .B(new_new_n331_), .Y(new_new_n333_));
  NO2        g0311(.A(i_1_), .B(i_7_), .Y(new_new_n334_));
  AO220      g0312(.A0(new_new_n334_), .A1(new_new_n333_), .B0(new_new_n323_), .B1(new_new_n233_), .Y(new_new_n335_));
  NA2        g0313(.A(new_new_n335_), .B(new_new_n42_), .Y(new_new_n336_));
  NA2        g0314(.A(new_new_n336_), .B(new_new_n327_), .Y(new_new_n337_));
  NO3        g0315(.A(new_new_n231_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n338_));
  NO3        g0316(.A(new_new_n322_), .B(i_2_), .C(i_1_), .Y(new_new_n339_));
  OAI210     g0317(.A0(new_new_n339_), .A1(new_new_n338_), .B0(i_6_), .Y(new_new_n340_));
  NO2        g0318(.A(new_new_n340_), .B(new_new_n319_), .Y(new_new_n341_));
  NOi21      g0319(.An(new_new_n156_), .B(new_new_n107_), .Y(new_new_n342_));
  NO2        g0320(.A(new_new_n342_), .B(new_new_n127_), .Y(new_new_n343_));
  OAI210     g0321(.A0(new_new_n343_), .A1(new_new_n341_), .B0(i_3_), .Y(new_new_n344_));
  INV        g0322(.A(new_new_n85_), .Y(new_new_n345_));
  NO2        g0323(.A(new_new_n291_), .B(new_new_n82_), .Y(new_new_n346_));
  NA2        g0324(.A(new_new_n346_), .B(new_new_n135_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n96_), .B(new_new_n198_), .Y(new_new_n348_));
  NA3        g0326(.A(new_new_n302_), .B(new_new_n348_), .C(new_new_n64_), .Y(new_new_n349_));
  AOI210     g0327(.A0(new_new_n349_), .A1(new_new_n347_), .B0(new_new_n345_), .Y(new_new_n350_));
  NO2        g0328(.A(new_new_n198_), .B(i_9_), .Y(new_new_n351_));
  NA2        g0329(.A(new_new_n351_), .B(new_new_n210_), .Y(new_new_n352_));
  NO2        g0330(.A(new_new_n352_), .B(new_new_n47_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n353_), .B(new_new_n350_), .Y(new_new_n354_));
  AOI210     g0332(.A0(new_new_n354_), .A1(new_new_n344_), .B0(new_new_n165_), .Y(new_new_n355_));
  AOI210     g0333(.A0(new_new_n337_), .A1(new_new_n311_), .B0(new_new_n355_), .Y(new_new_n356_));
  NOi32      g0334(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n357_));
  INV        g0335(.A(new_new_n357_), .Y(new_new_n358_));
  NAi21      g0336(.An(i_0_), .B(i_6_), .Y(new_new_n359_));
  NAi21      g0337(.An(i_1_), .B(i_5_), .Y(new_new_n360_));
  NA2        g0338(.A(new_new_n360_), .B(new_new_n359_), .Y(new_new_n361_));
  NA2        g0339(.A(new_new_n361_), .B(new_new_n25_), .Y(new_new_n362_));
  OAI210     g0340(.A0(new_new_n362_), .A1(new_new_n162_), .B0(new_new_n245_), .Y(new_new_n363_));
  NAi41      g0341(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n364_));
  OAI220     g0342(.A0(new_new_n364_), .A1(new_new_n360_), .B0(new_new_n224_), .B1(new_new_n162_), .Y(new_new_n365_));
  NO2        g0343(.A(new_new_n162_), .B(new_new_n160_), .Y(new_new_n366_));
  NOi32      g0344(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n367_));
  NAi21      g0345(.An(i_6_), .B(i_1_), .Y(new_new_n368_));
  NA3        g0346(.A(new_new_n368_), .B(new_new_n367_), .C(new_new_n47_), .Y(new_new_n369_));
  NO2        g0347(.A(new_new_n369_), .B(i_0_), .Y(new_new_n370_));
  OR3        g0348(.A(new_new_n370_), .B(new_new_n366_), .C(new_new_n365_), .Y(new_new_n371_));
  NO2        g0349(.A(i_1_), .B(new_new_n104_), .Y(new_new_n372_));
  NAi21      g0350(.An(i_3_), .B(i_4_), .Y(new_new_n373_));
  NO2        g0351(.A(new_new_n373_), .B(i_9_), .Y(new_new_n374_));
  AN2        g0352(.A(i_6_), .B(i_7_), .Y(new_new_n375_));
  OAI210     g0353(.A0(new_new_n375_), .A1(new_new_n372_), .B0(new_new_n374_), .Y(new_new_n376_));
  NA2        g0354(.A(i_2_), .B(i_7_), .Y(new_new_n377_));
  NO2        g0355(.A(new_new_n373_), .B(i_10_), .Y(new_new_n378_));
  NO2        g0356(.A(new_new_n376_), .B(new_new_n190_), .Y(new_new_n379_));
  AOI210     g0357(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n380_));
  OAI210     g0358(.A0(new_new_n380_), .A1(new_new_n193_), .B0(new_new_n378_), .Y(new_new_n381_));
  AOI220     g0359(.A0(new_new_n378_), .A1(new_new_n334_), .B0(new_new_n237_), .B1(new_new_n193_), .Y(new_new_n382_));
  AOI210     g0360(.A0(new_new_n382_), .A1(new_new_n381_), .B0(i_5_), .Y(new_new_n383_));
  NO4        g0361(.A(new_new_n383_), .B(new_new_n379_), .C(new_new_n371_), .D(new_new_n363_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n384_), .B(new_new_n358_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n386_));
  AN2        g0364(.A(i_12_), .B(i_5_), .Y(new_new_n387_));
  NO2        g0365(.A(i_4_), .B(new_new_n26_), .Y(new_new_n388_));
  INV        g0366(.A(new_new_n387_), .Y(new_new_n389_));
  NO2        g0367(.A(i_11_), .B(i_6_), .Y(new_new_n390_));
  NO2        g0368(.A(new_new_n241_), .B(i_5_), .Y(new_new_n391_));
  NO2        g0369(.A(i_5_), .B(i_10_), .Y(new_new_n392_));
  AOI220     g0370(.A0(new_new_n392_), .A1(new_new_n271_), .B0(new_new_n391_), .B1(new_new_n203_), .Y(new_new_n393_));
  NA2        g0371(.A(new_new_n147_), .B(new_new_n46_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n394_), .B(new_new_n393_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n395_), .B(new_new_n386_), .Y(new_new_n396_));
  NO2        g0374(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n397_));
  NO3        g0375(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n398_));
  NO2        g0376(.A(i_11_), .B(i_12_), .Y(new_new_n399_));
  NA3        g0377(.A(new_new_n116_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n400_), .B(new_new_n224_), .Y(new_new_n401_));
  NAi21      g0379(.An(i_13_), .B(i_0_), .Y(new_new_n402_));
  NO2        g0380(.A(new_new_n402_), .B(new_new_n238_), .Y(new_new_n403_));
  NA2        g0381(.A(new_new_n401_), .B(new_new_n403_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n404_), .B(new_new_n396_), .Y(new_new_n405_));
  NO2        g0383(.A(i_0_), .B(i_11_), .Y(new_new_n406_));
  INV        g0384(.A(i_5_), .Y(new_new_n407_));
  AN2        g0385(.A(i_1_), .B(i_6_), .Y(new_new_n408_));
  NOi21      g0386(.An(i_2_), .B(i_12_), .Y(new_new_n409_));
  NA2        g0387(.A(new_new_n409_), .B(new_new_n408_), .Y(new_new_n410_));
  NO2        g0388(.A(new_new_n410_), .B(new_new_n407_), .Y(new_new_n411_));
  NA2        g0389(.A(new_new_n145_), .B(i_9_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n412_), .B(i_4_), .Y(new_new_n413_));
  NA2        g0391(.A(new_new_n411_), .B(new_new_n413_), .Y(new_new_n414_));
  NAi21      g0392(.An(i_9_), .B(i_4_), .Y(new_new_n415_));
  OR2        g0393(.A(i_13_), .B(i_10_), .Y(new_new_n416_));
  NO3        g0394(.A(new_new_n416_), .B(new_new_n120_), .C(new_new_n415_), .Y(new_new_n417_));
  OR2        g0395(.A(new_new_n222_), .B(new_new_n221_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n104_), .B(new_new_n25_), .Y(new_new_n419_));
  NA2        g0397(.A(new_new_n283_), .B(new_new_n419_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n276_), .B(new_new_n216_), .Y(new_new_n421_));
  OAI220     g0399(.A0(new_new_n421_), .A1(new_new_n418_), .B0(new_new_n420_), .B1(new_new_n342_), .Y(new_new_n422_));
  INV        g0400(.A(new_new_n422_), .Y(new_new_n423_));
  AOI210     g0401(.A0(new_new_n423_), .A1(new_new_n414_), .B0(new_new_n26_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n321_), .B(new_new_n320_), .Y(new_new_n425_));
  AOI220     g0403(.A0(new_new_n293_), .A1(new_new_n287_), .B0(new_new_n290_), .B1(new_new_n312_), .Y(new_new_n426_));
  NO2        g0404(.A(new_new_n426_), .B(new_new_n173_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n187_), .B(new_new_n87_), .Y(new_new_n428_));
  AOI220     g0406(.A0(new_new_n428_), .A1(new_new_n292_), .B0(new_new_n278_), .B1(new_new_n216_), .Y(new_new_n429_));
  NO2        g0407(.A(new_new_n429_), .B(new_new_n285_), .Y(new_new_n430_));
  NO3        g0408(.A(new_new_n430_), .B(new_new_n427_), .C(new_new_n425_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n201_), .B(new_new_n99_), .Y(new_new_n432_));
  NA3        g0410(.A(new_new_n324_), .B(new_new_n166_), .C(new_new_n87_), .Y(new_new_n433_));
  AOI210     g0411(.A0(new_new_n433_), .A1(new_new_n432_), .B0(new_new_n322_), .Y(new_new_n434_));
  NA2        g0412(.A(new_new_n198_), .B(i_10_), .Y(new_new_n435_));
  NA3        g0413(.A(new_new_n257_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n436_));
  NA2        g0414(.A(new_new_n293_), .B(new_new_n233_), .Y(new_new_n437_));
  OAI220     g0415(.A0(new_new_n437_), .A1(new_new_n187_), .B0(new_new_n436_), .B1(new_new_n435_), .Y(new_new_n438_));
  NO2        g0416(.A(i_3_), .B(new_new_n49_), .Y(new_new_n439_));
  NA3        g0417(.A(new_new_n334_), .B(new_new_n333_), .C(new_new_n439_), .Y(new_new_n440_));
  NA2        g0418(.A(new_new_n314_), .B(new_new_n319_), .Y(new_new_n441_));
  OAI210     g0419(.A0(new_new_n441_), .A1(new_new_n194_), .B0(new_new_n440_), .Y(new_new_n442_));
  NO3        g0420(.A(new_new_n442_), .B(new_new_n438_), .C(new_new_n434_), .Y(new_new_n443_));
  AOI210     g0421(.A0(new_new_n443_), .A1(new_new_n431_), .B0(new_new_n272_), .Y(new_new_n444_));
  NO4        g0422(.A(new_new_n444_), .B(new_new_n424_), .C(new_new_n405_), .D(new_new_n385_), .Y(new_new_n445_));
  NO2        g0423(.A(new_new_n64_), .B(i_4_), .Y(new_new_n446_));
  NO2        g0424(.A(new_new_n74_), .B(i_13_), .Y(new_new_n447_));
  NA3        g0425(.A(new_new_n447_), .B(new_new_n446_), .C(i_2_), .Y(new_new_n448_));
  NO2        g0426(.A(i_10_), .B(i_9_), .Y(new_new_n449_));
  NAi21      g0427(.An(i_12_), .B(i_8_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n450_), .B(i_3_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n451_), .B(new_new_n449_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n47_), .B(i_4_), .Y(new_new_n453_));
  NO2        g0431(.A(new_new_n452_), .B(new_new_n448_), .Y(new_new_n454_));
  NA2        g0432(.A(new_new_n307_), .B(i_0_), .Y(new_new_n455_));
  NO3        g0433(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n456_));
  NA2        g0434(.A(new_new_n269_), .B(new_new_n100_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n457_), .B(new_new_n456_), .Y(new_new_n458_));
  NA2        g0436(.A(i_8_), .B(i_9_), .Y(new_new_n459_));
  NO2        g0437(.A(new_new_n458_), .B(new_new_n455_), .Y(new_new_n460_));
  NA2        g0438(.A(new_new_n250_), .B(new_new_n306_), .Y(new_new_n461_));
  NO3        g0439(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n462_));
  INV        g0440(.A(new_new_n462_), .Y(new_new_n463_));
  NA3        g0441(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n464_));
  NA4        g0442(.A(new_new_n148_), .B(new_new_n119_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n465_));
  OAI220     g0443(.A0(new_new_n465_), .A1(new_new_n464_), .B0(new_new_n463_), .B1(new_new_n461_), .Y(new_new_n466_));
  NO3        g0444(.A(new_new_n466_), .B(new_new_n460_), .C(new_new_n454_), .Y(new_new_n467_));
  NA2        g0445(.A(new_new_n292_), .B(new_new_n111_), .Y(new_new_n468_));
  OR2        g0446(.A(new_new_n468_), .B(new_new_n212_), .Y(new_new_n469_));
  OA210      g0447(.A0(new_new_n352_), .A1(new_new_n104_), .B0(new_new_n294_), .Y(new_new_n470_));
  OA220      g0448(.A0(new_new_n470_), .A1(new_new_n165_), .B0(new_new_n469_), .B1(new_new_n230_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n99_), .B(i_13_), .Y(new_new_n472_));
  NO2        g0450(.A(i_2_), .B(i_13_), .Y(new_new_n473_));
  NO3        g0451(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n474_));
  NO2        g0452(.A(i_6_), .B(i_7_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n475_), .B(new_new_n474_), .Y(new_new_n476_));
  NO2        g0454(.A(i_11_), .B(i_1_), .Y(new_new_n477_));
  NO2        g0455(.A(new_new_n74_), .B(i_3_), .Y(new_new_n478_));
  OR2        g0456(.A(i_11_), .B(i_8_), .Y(new_new_n479_));
  NOi21      g0457(.An(i_2_), .B(i_7_), .Y(new_new_n480_));
  NAi31      g0458(.An(new_new_n479_), .B(new_new_n480_), .C(new_new_n478_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n416_), .B(i_6_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n482_), .B(new_new_n446_), .Y(new_new_n483_));
  NO2        g0461(.A(new_new_n483_), .B(new_new_n481_), .Y(new_new_n484_));
  NO2        g0462(.A(i_3_), .B(new_new_n198_), .Y(new_new_n485_));
  NO2        g0463(.A(i_6_), .B(i_10_), .Y(new_new_n486_));
  NA4        g0464(.A(new_new_n486_), .B(new_new_n311_), .C(new_new_n485_), .D(new_new_n235_), .Y(new_new_n487_));
  NO2        g0465(.A(new_new_n487_), .B(new_new_n158_), .Y(new_new_n488_));
  NA3        g0466(.A(new_new_n244_), .B(new_new_n175_), .C(new_new_n135_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n490_));
  NO2        g0468(.A(new_new_n160_), .B(i_3_), .Y(new_new_n491_));
  NAi31      g0469(.An(new_new_n490_), .B(new_new_n491_), .C(new_new_n227_), .Y(new_new_n492_));
  NA3        g0470(.A(new_new_n397_), .B(new_new_n183_), .C(new_new_n152_), .Y(new_new_n493_));
  NA3        g0471(.A(new_new_n493_), .B(new_new_n492_), .C(new_new_n489_), .Y(new_new_n494_));
  NO3        g0472(.A(new_new_n494_), .B(new_new_n488_), .C(new_new_n484_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n456_), .B(new_new_n387_), .Y(new_new_n496_));
  NAi21      g0474(.An(new_new_n222_), .B(new_new_n399_), .Y(new_new_n497_));
  NO2        g0475(.A(new_new_n26_), .B(i_5_), .Y(new_new_n498_));
  NO2        g0476(.A(i_0_), .B(new_new_n87_), .Y(new_new_n499_));
  NA3        g0477(.A(new_new_n499_), .B(new_new_n498_), .C(new_new_n145_), .Y(new_new_n500_));
  OR3        g0478(.A(new_new_n300_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n501_));
  NO2        g0479(.A(new_new_n501_), .B(new_new_n500_), .Y(new_new_n502_));
  NA2        g0480(.A(new_new_n27_), .B(i_10_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n311_), .B(new_new_n237_), .Y(new_new_n504_));
  OAI220     g0482(.A0(new_new_n504_), .A1(new_new_n436_), .B0(new_new_n503_), .B1(new_new_n472_), .Y(new_new_n505_));
  NA4        g0483(.A(new_new_n304_), .B(new_new_n225_), .C(new_new_n74_), .D(new_new_n235_), .Y(new_new_n506_));
  NO2        g0484(.A(new_new_n506_), .B(new_new_n476_), .Y(new_new_n507_));
  NO3        g0485(.A(new_new_n507_), .B(new_new_n505_), .C(new_new_n502_), .Y(new_new_n508_));
  NA4        g0486(.A(new_new_n508_), .B(new_new_n495_), .C(new_new_n471_), .D(new_new_n467_), .Y(new_new_n509_));
  NA3        g0487(.A(new_new_n304_), .B(new_new_n180_), .C(new_new_n178_), .Y(new_new_n510_));
  OAI210     g0488(.A0(new_new_n298_), .A1(new_new_n185_), .B0(new_new_n510_), .Y(new_new_n511_));
  AN2        g0489(.A(new_new_n287_), .B(new_new_n232_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n512_), .B(new_new_n511_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n311_), .B(new_new_n167_), .Y(new_new_n514_));
  OAI210     g0492(.A0(new_new_n514_), .A1(new_new_n230_), .B0(new_new_n305_), .Y(new_new_n515_));
  NA2        g0493(.A(new_new_n515_), .B(new_new_n323_), .Y(new_new_n516_));
  NA4        g0494(.A(new_new_n447_), .B(new_new_n446_), .C(new_new_n208_), .D(i_2_), .Y(new_new_n517_));
  INV        g0495(.A(new_new_n517_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n387_), .B(new_new_n226_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n357_), .B(new_new_n74_), .Y(new_new_n520_));
  NA2        g0498(.A(new_new_n375_), .B(new_new_n367_), .Y(new_new_n521_));
  OR2        g0499(.A(new_new_n519_), .B(new_new_n521_), .Y(new_new_n522_));
  NO2        g0500(.A(new_new_n36_), .B(i_8_), .Y(new_new_n523_));
  NAi41      g0501(.An(new_new_n520_), .B(new_new_n486_), .C(new_new_n523_), .D(new_new_n47_), .Y(new_new_n524_));
  AOI210     g0502(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n417_), .Y(new_new_n525_));
  NA3        g0503(.A(new_new_n525_), .B(new_new_n524_), .C(new_new_n522_), .Y(new_new_n526_));
  AOI210     g0504(.A0(new_new_n518_), .A1(new_new_n209_), .B0(new_new_n526_), .Y(new_new_n527_));
  AOI210     g0505(.A0(new_new_n199_), .A1(i_9_), .B0(new_new_n268_), .Y(new_new_n528_));
  NO2        g0506(.A(new_new_n528_), .B(new_new_n204_), .Y(new_new_n529_));
  NO2        g0507(.A(new_new_n187_), .B(new_new_n87_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n530_), .B(new_new_n529_), .Y(new_new_n531_));
  NA4        g0509(.A(new_new_n531_), .B(new_new_n527_), .C(new_new_n516_), .D(new_new_n513_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n391_), .B(new_new_n292_), .Y(new_new_n533_));
  OAI210     g0511(.A0(new_new_n389_), .A1(new_new_n172_), .B0(new_new_n533_), .Y(new_new_n534_));
  NO2        g0512(.A(i_12_), .B(new_new_n198_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n535_), .B(new_new_n226_), .Y(new_new_n536_));
  NO3        g0514(.A(new_new_n1033_), .B(new_new_n536_), .C(new_new_n468_), .Y(new_new_n537_));
  NOi31      g0515(.An(new_new_n314_), .B(new_new_n416_), .C(new_new_n38_), .Y(new_new_n538_));
  OAI210     g0516(.A0(new_new_n538_), .A1(new_new_n537_), .B0(new_new_n534_), .Y(new_new_n539_));
  NO2        g0517(.A(i_8_), .B(i_7_), .Y(new_new_n540_));
  OAI210     g0518(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n541_));
  NA2        g0519(.A(new_new_n541_), .B(new_new_n225_), .Y(new_new_n542_));
  AOI220     g0520(.A0(new_new_n324_), .A1(new_new_n40_), .B0(new_new_n233_), .B1(new_new_n211_), .Y(new_new_n543_));
  OAI220     g0521(.A0(new_new_n543_), .A1(new_new_n187_), .B0(new_new_n542_), .B1(new_new_n241_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n45_), .B(i_10_), .Y(new_new_n545_));
  NO2        g0523(.A(new_new_n545_), .B(i_6_), .Y(new_new_n546_));
  NA3        g0524(.A(new_new_n546_), .B(new_new_n544_), .C(new_new_n540_), .Y(new_new_n547_));
  NO2        g0525(.A(new_new_n472_), .B(new_new_n136_), .Y(new_new_n548_));
  NA2        g0526(.A(new_new_n548_), .B(new_new_n268_), .Y(new_new_n549_));
  NOi31      g0527(.An(new_new_n290_), .B(new_new_n298_), .C(new_new_n185_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n550_), .B(new_new_n462_), .Y(new_new_n551_));
  NA4        g0529(.A(new_new_n551_), .B(new_new_n549_), .C(new_new_n547_), .D(new_new_n539_), .Y(new_new_n552_));
  NA3        g0530(.A(new_new_n223_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n283_), .B(new_new_n85_), .Y(new_new_n554_));
  AOI210     g0532(.A0(new_new_n553_), .A1(new_new_n347_), .B0(new_new_n554_), .Y(new_new_n555_));
  NA2        g0533(.A(new_new_n293_), .B(new_new_n287_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n556_), .B(new_new_n177_), .Y(new_new_n557_));
  AOI210     g0535(.A0(new_new_n368_), .A1(new_new_n47_), .B0(new_new_n372_), .Y(new_new_n558_));
  NA2        g0536(.A(i_0_), .B(new_new_n49_), .Y(new_new_n559_));
  NA3        g0537(.A(new_new_n535_), .B(new_new_n274_), .C(new_new_n559_), .Y(new_new_n560_));
  NO2        g0538(.A(new_new_n558_), .B(new_new_n560_), .Y(new_new_n561_));
  NO3        g0539(.A(new_new_n561_), .B(new_new_n557_), .C(new_new_n555_), .Y(new_new_n562_));
  NO4        g0540(.A(new_new_n251_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n563_));
  NO3        g0541(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n564_));
  NO2        g0542(.A(new_new_n231_), .B(new_new_n36_), .Y(new_new_n565_));
  AN2        g0543(.A(new_new_n565_), .B(new_new_n564_), .Y(new_new_n566_));
  OA210      g0544(.A0(new_new_n566_), .A1(new_new_n563_), .B0(new_new_n357_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n416_), .B(i_1_), .Y(new_new_n568_));
  NOi31      g0546(.An(new_new_n568_), .B(new_new_n457_), .C(new_new_n74_), .Y(new_new_n569_));
  AN4        g0547(.A(new_new_n569_), .B(new_new_n413_), .C(new_new_n498_), .D(i_2_), .Y(new_new_n570_));
  NO2        g0548(.A(new_new_n426_), .B(new_new_n181_), .Y(new_new_n571_));
  NO3        g0549(.A(new_new_n571_), .B(new_new_n570_), .C(new_new_n567_), .Y(new_new_n572_));
  NOi21      g0550(.An(i_10_), .B(i_6_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n575_));
  NA2        g0553(.A(new_new_n314_), .B(new_new_n167_), .Y(new_new_n576_));
  AOI220     g0554(.A0(new_new_n576_), .A1(new_new_n437_), .B0(new_new_n188_), .B1(new_new_n186_), .Y(new_new_n577_));
  NO2        g0555(.A(new_new_n203_), .B(new_new_n37_), .Y(new_new_n578_));
  NOi31      g0556(.An(new_new_n149_), .B(new_new_n578_), .C(new_new_n330_), .Y(new_new_n579_));
  NO2        g0557(.A(new_new_n579_), .B(new_new_n577_), .Y(new_new_n580_));
  INV        g0558(.A(new_new_n317_), .Y(new_new_n581_));
  NO2        g0559(.A(i_12_), .B(new_new_n87_), .Y(new_new_n582_));
  NA2        g0560(.A(new_new_n178_), .B(i_0_), .Y(new_new_n583_));
  NO3        g0561(.A(new_new_n583_), .B(new_new_n340_), .C(new_new_n298_), .Y(new_new_n584_));
  OR2        g0562(.A(i_2_), .B(i_5_), .Y(new_new_n585_));
  OR2        g0563(.A(new_new_n585_), .B(new_new_n408_), .Y(new_new_n586_));
  AOI210     g0564(.A0(new_new_n377_), .A1(new_new_n243_), .B0(new_new_n203_), .Y(new_new_n587_));
  AOI210     g0565(.A0(new_new_n587_), .A1(new_new_n586_), .B0(new_new_n497_), .Y(new_new_n588_));
  NO2        g0566(.A(new_new_n588_), .B(new_new_n584_), .Y(new_new_n589_));
  NA4        g0567(.A(new_new_n589_), .B(new_new_n580_), .C(new_new_n572_), .D(new_new_n562_), .Y(new_new_n590_));
  NO4        g0568(.A(new_new_n590_), .B(new_new_n552_), .C(new_new_n532_), .D(new_new_n509_), .Y(new_new_n591_));
  NA4        g0569(.A(new_new_n591_), .B(new_new_n445_), .C(new_new_n356_), .D(new_new_n310_), .Y(mai7));
  NO2        g0570(.A(new_new_n96_), .B(new_new_n55_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n111_), .B(new_new_n93_), .Y(new_new_n594_));
  NA2        g0572(.A(new_new_n388_), .B(new_new_n594_), .Y(new_new_n595_));
  NA2        g0573(.A(new_new_n486_), .B(new_new_n85_), .Y(new_new_n596_));
  NA2        g0574(.A(i_11_), .B(new_new_n198_), .Y(new_new_n597_));
  NA2        g0575(.A(new_new_n147_), .B(new_new_n597_), .Y(new_new_n598_));
  OAI210     g0576(.A0(new_new_n598_), .A1(new_new_n596_), .B0(new_new_n595_), .Y(new_new_n599_));
  NA3        g0577(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n600_));
  NO2        g0578(.A(new_new_n235_), .B(i_4_), .Y(new_new_n601_));
  NA2        g0579(.A(new_new_n601_), .B(i_8_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n108_), .B(new_new_n600_), .Y(new_new_n603_));
  NA2        g0581(.A(i_2_), .B(new_new_n87_), .Y(new_new_n604_));
  OAI210     g0582(.A0(new_new_n90_), .A1(new_new_n208_), .B0(new_new_n209_), .Y(new_new_n605_));
  NO2        g0583(.A(i_7_), .B(new_new_n37_), .Y(new_new_n606_));
  NA2        g0584(.A(i_4_), .B(i_8_), .Y(new_new_n607_));
  AOI210     g0585(.A0(new_new_n607_), .A1(new_new_n304_), .B0(new_new_n606_), .Y(new_new_n608_));
  OAI220     g0586(.A0(new_new_n608_), .A1(new_new_n604_), .B0(new_new_n605_), .B1(i_13_), .Y(new_new_n609_));
  NO4        g0587(.A(new_new_n609_), .B(new_new_n603_), .C(new_new_n599_), .D(new_new_n593_), .Y(new_new_n610_));
  AOI210     g0588(.A0(new_new_n131_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n611_));
  AOI210     g0589(.A0(new_new_n611_), .A1(new_new_n235_), .B0(new_new_n164_), .Y(new_new_n612_));
  OR2        g0590(.A(i_6_), .B(i_10_), .Y(new_new_n613_));
  NO2        g0591(.A(new_new_n613_), .B(new_new_n23_), .Y(new_new_n614_));
  OR3        g0592(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n615_));
  NO3        g0593(.A(new_new_n615_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n616_));
  INV        g0594(.A(new_new_n205_), .Y(new_new_n617_));
  NO2        g0595(.A(new_new_n616_), .B(new_new_n614_), .Y(new_new_n618_));
  OA220      g0596(.A0(new_new_n618_), .A1(new_new_n581_), .B0(new_new_n612_), .B1(new_new_n270_), .Y(new_new_n619_));
  AOI210     g0597(.A0(new_new_n619_), .A1(new_new_n610_), .B0(new_new_n64_), .Y(new_new_n620_));
  NOi21      g0598(.An(i_11_), .B(i_7_), .Y(new_new_n621_));
  AO210      g0599(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n622_));
  NO2        g0600(.A(new_new_n622_), .B(new_new_n621_), .Y(new_new_n623_));
  NA2        g0601(.A(new_new_n623_), .B(new_new_n211_), .Y(new_new_n624_));
  NA3        g0602(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n625_));
  NO2        g0603(.A(new_new_n624_), .B(new_new_n64_), .Y(new_new_n626_));
  NA2        g0604(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n627_));
  AO210      g0605(.A0(new_new_n627_), .A1(new_new_n382_), .B0(new_new_n41_), .Y(new_new_n628_));
  NA2        g0606(.A(new_new_n227_), .B(new_new_n64_), .Y(new_new_n629_));
  NO2        g0607(.A(new_new_n64_), .B(i_9_), .Y(new_new_n630_));
  NO2        g0608(.A(i_1_), .B(i_12_), .Y(new_new_n631_));
  NA3        g0609(.A(new_new_n631_), .B(new_new_n113_), .C(new_new_n24_), .Y(new_new_n632_));
  BUFFER     g0610(.A(new_new_n632_), .Y(new_new_n633_));
  NA3        g0611(.A(new_new_n633_), .B(new_new_n629_), .C(new_new_n628_), .Y(new_new_n634_));
  OAI210     g0612(.A0(new_new_n634_), .A1(new_new_n626_), .B0(i_6_), .Y(new_new_n635_));
  NO2        g0613(.A(new_new_n625_), .B(new_new_n111_), .Y(new_new_n636_));
  NA2        g0614(.A(new_new_n636_), .B(new_new_n582_), .Y(new_new_n637_));
  NO2        g0615(.A(i_6_), .B(i_11_), .Y(new_new_n638_));
  NA2        g0616(.A(new_new_n637_), .B(new_new_n458_), .Y(new_new_n639_));
  NO4        g0617(.A(new_new_n221_), .B(new_new_n131_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n640_));
  NA2        g0618(.A(new_new_n640_), .B(new_new_n630_), .Y(new_new_n641_));
  NA2        g0619(.A(new_new_n235_), .B(i_6_), .Y(new_new_n642_));
  NA2        g0620(.A(i_1_), .B(new_new_n260_), .Y(new_new_n643_));
  OAI210     g0621(.A0(new_new_n643_), .A1(new_new_n45_), .B0(new_new_n641_), .Y(new_new_n644_));
  INV        g0622(.A(i_2_), .Y(new_new_n645_));
  NA2        g0623(.A(new_new_n141_), .B(i_9_), .Y(new_new_n646_));
  NA3        g0624(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n47_), .B(i_1_), .Y(new_new_n648_));
  NA3        g0626(.A(new_new_n648_), .B(new_new_n269_), .C(new_new_n45_), .Y(new_new_n649_));
  OAI220     g0627(.A0(new_new_n649_), .A1(new_new_n647_), .B0(new_new_n646_), .B1(new_new_n645_), .Y(new_new_n650_));
  NA3        g0628(.A(new_new_n630_), .B(new_new_n317_), .C(i_6_), .Y(new_new_n651_));
  NO2        g0629(.A(new_new_n651_), .B(new_new_n23_), .Y(new_new_n652_));
  AOI210     g0630(.A0(new_new_n477_), .A1(new_new_n419_), .B0(new_new_n240_), .Y(new_new_n653_));
  NO2        g0631(.A(new_new_n653_), .B(new_new_n604_), .Y(new_new_n654_));
  NO2        g0632(.A(i_11_), .B(new_new_n37_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n655_), .B(new_new_n24_), .Y(new_new_n656_));
  OR3        g0634(.A(new_new_n654_), .B(new_new_n652_), .C(new_new_n650_), .Y(new_new_n657_));
  NO3        g0635(.A(new_new_n657_), .B(new_new_n644_), .C(new_new_n639_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n235_), .B(new_new_n104_), .Y(new_new_n659_));
  NO2        g0637(.A(new_new_n659_), .B(new_new_n621_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n660_), .B(i_1_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n661_), .B(new_new_n615_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n415_), .B(new_new_n87_), .Y(new_new_n663_));
  NA2        g0641(.A(new_new_n662_), .B(new_new_n47_), .Y(new_new_n664_));
  NA2        g0642(.A(i_3_), .B(new_new_n198_), .Y(new_new_n665_));
  NO2        g0643(.A(new_new_n665_), .B(new_new_n118_), .Y(new_new_n666_));
  AN2        g0644(.A(new_new_n666_), .B(new_new_n546_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n231_), .B(new_new_n45_), .Y(new_new_n668_));
  NO3        g0646(.A(new_new_n668_), .B(new_new_n307_), .C(new_new_n236_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n120_), .B(new_new_n37_), .Y(new_new_n670_));
  NO2        g0648(.A(new_new_n670_), .B(i_6_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n87_), .B(i_9_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n672_), .B(new_new_n64_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n673_), .B(new_new_n631_), .Y(new_new_n674_));
  NO4        g0652(.A(new_new_n674_), .B(new_new_n671_), .C(new_new_n669_), .D(i_4_), .Y(new_new_n675_));
  NA2        g0653(.A(i_1_), .B(i_3_), .Y(new_new_n676_));
  NO2        g0654(.A(new_new_n459_), .B(new_new_n96_), .Y(new_new_n677_));
  AOI210     g0655(.A0(new_new_n668_), .A1(new_new_n573_), .B0(new_new_n677_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n678_), .B(new_new_n676_), .Y(new_new_n679_));
  NO3        g0657(.A(new_new_n679_), .B(new_new_n675_), .C(new_new_n667_), .Y(new_new_n680_));
  NA4        g0658(.A(new_new_n680_), .B(new_new_n664_), .C(new_new_n658_), .D(new_new_n635_), .Y(new_new_n681_));
  AN2        g0659(.A(new_new_n244_), .B(new_new_n87_), .Y(new_new_n682_));
  NA2        g0660(.A(new_new_n375_), .B(new_new_n374_), .Y(new_new_n683_));
  INV        g0661(.A(new_new_n683_), .Y(new_new_n684_));
  OAI210     g0662(.A0(new_new_n684_), .A1(new_new_n682_), .B0(i_1_), .Y(new_new_n685_));
  AOI210     g0663(.A0(new_new_n269_), .A1(new_new_n100_), .B0(i_1_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n373_), .B(i_2_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n687_), .B(new_new_n686_), .Y(new_new_n688_));
  OAI210     g0666(.A0(new_new_n651_), .A1(new_new_n450_), .B0(new_new_n688_), .Y(new_new_n689_));
  INV        g0667(.A(new_new_n689_), .Y(new_new_n690_));
  AOI210     g0668(.A0(new_new_n690_), .A1(new_new_n685_), .B0(i_13_), .Y(new_new_n691_));
  OR2        g0669(.A(i_11_), .B(i_7_), .Y(new_new_n692_));
  NA3        g0670(.A(new_new_n692_), .B(new_new_n109_), .C(new_new_n141_), .Y(new_new_n693_));
  AOI220     g0671(.A0(new_new_n473_), .A1(new_new_n164_), .B0(new_new_n453_), .B1(new_new_n141_), .Y(new_new_n694_));
  OAI210     g0672(.A0(new_new_n694_), .A1(new_new_n45_), .B0(new_new_n693_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n55_), .B(i_12_), .Y(new_new_n696_));
  INV        g0674(.A(new_new_n696_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n480_), .B(new_new_n24_), .Y(new_new_n698_));
  AOI220     g0676(.A0(new_new_n698_), .A1(new_new_n663_), .B0(new_new_n244_), .B1(new_new_n134_), .Y(new_new_n699_));
  OAI220     g0677(.A0(new_new_n699_), .A1(new_new_n41_), .B0(new_new_n697_), .B1(new_new_n96_), .Y(new_new_n700_));
  AOI210     g0678(.A0(new_new_n695_), .A1(new_new_n331_), .B0(new_new_n700_), .Y(new_new_n701_));
  INV        g0679(.A(new_new_n118_), .Y(new_new_n702_));
  AOI220     g0680(.A0(new_new_n702_), .A1(new_new_n73_), .B0(new_new_n390_), .B1(new_new_n648_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n703_), .B(new_new_n241_), .Y(new_new_n704_));
  AOI210     g0682(.A0(new_new_n450_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n705_));
  NOi31      g0683(.An(new_new_n705_), .B(new_new_n596_), .C(new_new_n45_), .Y(new_new_n706_));
  NA2        g0684(.A(new_new_n130_), .B(i_13_), .Y(new_new_n707_));
  NO2        g0685(.A(new_new_n647_), .B(new_new_n118_), .Y(new_new_n708_));
  INV        g0686(.A(new_new_n708_), .Y(new_new_n709_));
  OAI220     g0687(.A0(new_new_n709_), .A1(new_new_n72_), .B0(new_new_n707_), .B1(new_new_n686_), .Y(new_new_n710_));
  NO3        g0688(.A(new_new_n72_), .B(new_new_n32_), .C(new_new_n104_), .Y(new_new_n711_));
  NA2        g0689(.A(new_new_n26_), .B(new_new_n198_), .Y(new_new_n712_));
  NA2        g0690(.A(new_new_n712_), .B(i_7_), .Y(new_new_n713_));
  NO3        g0691(.A(new_new_n480_), .B(new_new_n235_), .C(new_new_n87_), .Y(new_new_n714_));
  AOI210     g0692(.A0(new_new_n714_), .A1(new_new_n713_), .B0(new_new_n711_), .Y(new_new_n715_));
  AOI220     g0693(.A0(new_new_n390_), .A1(new_new_n648_), .B0(new_new_n95_), .B1(new_new_n105_), .Y(new_new_n716_));
  OAI220     g0694(.A0(new_new_n716_), .A1(new_new_n602_), .B0(new_new_n715_), .B1(new_new_n617_), .Y(new_new_n717_));
  NO4        g0695(.A(new_new_n717_), .B(new_new_n710_), .C(new_new_n706_), .D(new_new_n704_), .Y(new_new_n718_));
  OR2        g0696(.A(i_11_), .B(i_6_), .Y(new_new_n719_));
  NA3        g0697(.A(new_new_n601_), .B(new_new_n712_), .C(i_7_), .Y(new_new_n720_));
  AOI210     g0698(.A0(new_new_n720_), .A1(new_new_n709_), .B0(new_new_n719_), .Y(new_new_n721_));
  NA3        g0699(.A(new_new_n409_), .B(new_new_n606_), .C(new_new_n100_), .Y(new_new_n722_));
  NA2        g0700(.A(new_new_n638_), .B(i_13_), .Y(new_new_n723_));
  NAi21      g0701(.An(i_11_), .B(i_12_), .Y(new_new_n724_));
  NOi41      g0702(.An(new_new_n114_), .B(new_new_n724_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n725_));
  NO3        g0703(.A(new_new_n480_), .B(new_new_n582_), .C(new_new_n607_), .Y(new_new_n726_));
  AOI220     g0704(.A0(new_new_n726_), .A1(new_new_n311_), .B0(new_new_n725_), .B1(new_new_n47_), .Y(new_new_n727_));
  NA3        g0705(.A(new_new_n727_), .B(new_new_n723_), .C(new_new_n722_), .Y(new_new_n728_));
  OAI210     g0706(.A0(new_new_n728_), .A1(new_new_n721_), .B0(new_new_n64_), .Y(new_new_n729_));
  NO2        g0707(.A(i_2_), .B(i_12_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n372_), .B(new_new_n730_), .Y(new_new_n731_));
  NA2        g0709(.A(i_8_), .B(new_new_n25_), .Y(new_new_n732_));
  NO3        g0710(.A(new_new_n732_), .B(new_new_n388_), .C(new_new_n601_), .Y(new_new_n733_));
  OAI210     g0711(.A0(new_new_n733_), .A1(new_new_n374_), .B0(new_new_n372_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n131_), .B(i_2_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n735_), .B(new_new_n631_), .Y(new_new_n736_));
  NA3        g0714(.A(new_new_n736_), .B(new_new_n734_), .C(new_new_n731_), .Y(new_new_n737_));
  NA3        g0715(.A(new_new_n737_), .B(new_new_n46_), .C(new_new_n226_), .Y(new_new_n738_));
  NA4        g0716(.A(new_new_n738_), .B(new_new_n729_), .C(new_new_n718_), .D(new_new_n701_), .Y(new_new_n739_));
  OR4        g0717(.A(new_new_n739_), .B(new_new_n691_), .C(new_new_n681_), .D(new_new_n620_), .Y(mai5));
  NA2        g0718(.A(new_new_n660_), .B(new_new_n271_), .Y(new_new_n741_));
  AN2        g0719(.A(new_new_n24_), .B(i_10_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n742_), .B(new_new_n730_), .C(new_new_n111_), .Y(new_new_n743_));
  NO2        g0721(.A(new_new_n602_), .B(i_11_), .Y(new_new_n744_));
  NA2        g0722(.A(new_new_n90_), .B(new_new_n744_), .Y(new_new_n745_));
  NA3        g0723(.A(new_new_n745_), .B(new_new_n743_), .C(new_new_n741_), .Y(new_new_n746_));
  NO3        g0724(.A(i_11_), .B(new_new_n235_), .C(i_13_), .Y(new_new_n747_));
  NO2        g0725(.A(new_new_n127_), .B(new_new_n23_), .Y(new_new_n748_));
  NA2        g0726(.A(i_12_), .B(i_8_), .Y(new_new_n749_));
  OAI210     g0727(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n749_), .Y(new_new_n750_));
  INV        g0728(.A(new_new_n449_), .Y(new_new_n751_));
  AOI220     g0729(.A0(new_new_n317_), .A1(new_new_n575_), .B0(new_new_n750_), .B1(new_new_n748_), .Y(new_new_n752_));
  INV        g0730(.A(new_new_n752_), .Y(new_new_n753_));
  NO2        g0731(.A(new_new_n753_), .B(new_new_n746_), .Y(new_new_n754_));
  INV        g0732(.A(new_new_n175_), .Y(new_new_n755_));
  INV        g0733(.A(new_new_n244_), .Y(new_new_n756_));
  OAI210     g0734(.A0(new_new_n687_), .A1(new_new_n451_), .B0(new_new_n114_), .Y(new_new_n757_));
  AOI210     g0735(.A0(new_new_n757_), .A1(new_new_n756_), .B0(new_new_n755_), .Y(new_new_n758_));
  NO2        g0736(.A(new_new_n459_), .B(new_new_n26_), .Y(new_new_n759_));
  NO2        g0737(.A(new_new_n759_), .B(new_new_n419_), .Y(new_new_n760_));
  NA2        g0738(.A(new_new_n760_), .B(i_2_), .Y(new_new_n761_));
  INV        g0739(.A(new_new_n761_), .Y(new_new_n762_));
  AOI210     g0740(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n416_), .Y(new_new_n763_));
  AOI210     g0741(.A0(new_new_n763_), .A1(new_new_n762_), .B0(new_new_n758_), .Y(new_new_n764_));
  NO2        g0742(.A(new_new_n195_), .B(new_new_n128_), .Y(new_new_n765_));
  OAI210     g0743(.A0(new_new_n765_), .A1(new_new_n748_), .B0(i_2_), .Y(new_new_n766_));
  INV        g0744(.A(new_new_n176_), .Y(new_new_n767_));
  NO3        g0745(.A(new_new_n622_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n768_));
  AOI210     g0746(.A0(new_new_n767_), .A1(new_new_n90_), .B0(new_new_n768_), .Y(new_new_n769_));
  AOI210     g0747(.A0(new_new_n769_), .A1(new_new_n766_), .B0(new_new_n198_), .Y(new_new_n770_));
  OA210      g0748(.A0(new_new_n623_), .A1(new_new_n129_), .B0(i_13_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n205_), .B(new_new_n208_), .Y(new_new_n772_));
  NA2        g0750(.A(new_new_n154_), .B(new_new_n597_), .Y(new_new_n773_));
  AOI210     g0751(.A0(new_new_n773_), .A1(new_new_n772_), .B0(new_new_n377_), .Y(new_new_n774_));
  AOI210     g0752(.A0(new_new_n213_), .A1(new_new_n151_), .B0(new_new_n523_), .Y(new_new_n775_));
  NA2        g0753(.A(new_new_n775_), .B(new_new_n419_), .Y(new_new_n776_));
  NO2        g0754(.A(new_new_n105_), .B(new_new_n45_), .Y(new_new_n777_));
  INV        g0755(.A(new_new_n299_), .Y(new_new_n778_));
  NA4        g0756(.A(new_new_n778_), .B(new_new_n304_), .C(new_new_n127_), .D(new_new_n43_), .Y(new_new_n779_));
  OAI210     g0757(.A0(new_new_n779_), .A1(new_new_n777_), .B0(new_new_n776_), .Y(new_new_n780_));
  NO4        g0758(.A(new_new_n780_), .B(new_new_n774_), .C(new_new_n771_), .D(new_new_n770_), .Y(new_new_n781_));
  NA2        g0759(.A(new_new_n575_), .B(new_new_n28_), .Y(new_new_n782_));
  NA2        g0760(.A(new_new_n747_), .B(new_new_n275_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(new_new_n782_), .Y(new_new_n784_));
  NO2        g0762(.A(new_new_n63_), .B(i_12_), .Y(new_new_n785_));
  NO2        g0763(.A(new_new_n785_), .B(new_new_n129_), .Y(new_new_n786_));
  NO2        g0764(.A(new_new_n786_), .B(new_new_n597_), .Y(new_new_n787_));
  AOI220     g0765(.A0(new_new_n787_), .A1(new_new_n36_), .B0(new_new_n784_), .B1(new_new_n47_), .Y(new_new_n788_));
  NA4        g0766(.A(new_new_n788_), .B(new_new_n781_), .C(new_new_n764_), .D(new_new_n754_), .Y(mai6));
  NO3        g0767(.A(new_new_n255_), .B(new_new_n306_), .C(i_1_), .Y(new_new_n790_));
  NO2        g0768(.A(new_new_n190_), .B(new_new_n142_), .Y(new_new_n791_));
  OAI210     g0769(.A0(new_new_n791_), .A1(new_new_n790_), .B0(new_new_n735_), .Y(new_new_n792_));
  NA4        g0770(.A(new_new_n392_), .B(new_new_n485_), .C(new_new_n72_), .D(new_new_n104_), .Y(new_new_n793_));
  INV        g0771(.A(new_new_n793_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n224_), .B(new_new_n490_), .Y(new_new_n795_));
  NO2        g0773(.A(i_11_), .B(i_9_), .Y(new_new_n796_));
  NO2        g0774(.A(new_new_n794_), .B(new_new_n329_), .Y(new_new_n797_));
  AO210      g0775(.A0(new_new_n797_), .A1(new_new_n792_), .B0(i_12_), .Y(new_new_n798_));
  NA2        g0776(.A(new_new_n378_), .B(new_new_n334_), .Y(new_new_n799_));
  NA2        g0777(.A(new_new_n582_), .B(new_new_n64_), .Y(new_new_n800_));
  BUFFER     g0778(.A(new_new_n627_), .Y(new_new_n801_));
  NA3        g0779(.A(new_new_n801_), .B(new_new_n800_), .C(new_new_n799_), .Y(new_new_n802_));
  INV        g0780(.A(new_new_n202_), .Y(new_new_n803_));
  AOI220     g0781(.A0(new_new_n803_), .A1(new_new_n796_), .B0(new_new_n802_), .B1(new_new_n74_), .Y(new_new_n804_));
  INV        g0782(.A(new_new_n328_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n76_), .B(new_new_n134_), .Y(new_new_n806_));
  INV        g0784(.A(new_new_n127_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n807_), .B(new_new_n47_), .Y(new_new_n808_));
  AOI210     g0786(.A0(new_new_n808_), .A1(new_new_n806_), .B0(new_new_n805_), .Y(new_new_n809_));
  NO2        g0787(.A(new_new_n251_), .B(i_9_), .Y(new_new_n810_));
  NA2        g0788(.A(new_new_n810_), .B(new_new_n785_), .Y(new_new_n811_));
  AOI210     g0789(.A0(new_new_n811_), .A1(new_new_n521_), .B0(new_new_n190_), .Y(new_new_n812_));
  NO2        g0790(.A(new_new_n32_), .B(i_11_), .Y(new_new_n813_));
  NAi32      g0791(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n814_));
  NO2        g0792(.A(new_new_n719_), .B(new_new_n814_), .Y(new_new_n815_));
  OR3        g0793(.A(new_new_n815_), .B(new_new_n812_), .C(new_new_n809_), .Y(new_new_n816_));
  NO2        g0794(.A(new_new_n692_), .B(i_2_), .Y(new_new_n817_));
  NA2        g0795(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n818_));
  NO2        g0796(.A(new_new_n818_), .B(new_new_n408_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n819_), .B(new_new_n817_), .Y(new_new_n820_));
  AO220      g0798(.A0(new_new_n361_), .A1(new_new_n351_), .B0(new_new_n398_), .B1(new_new_n597_), .Y(new_new_n821_));
  NA3        g0799(.A(new_new_n821_), .B(new_new_n256_), .C(i_7_), .Y(new_new_n822_));
  OR2        g0800(.A(new_new_n623_), .B(new_new_n451_), .Y(new_new_n823_));
  NA3        g0801(.A(new_new_n823_), .B(new_new_n150_), .C(new_new_n70_), .Y(new_new_n824_));
  OR2        g0802(.A(new_new_n751_), .B(new_new_n36_), .Y(new_new_n825_));
  NA4        g0803(.A(new_new_n825_), .B(new_new_n824_), .C(new_new_n822_), .D(new_new_n820_), .Y(new_new_n826_));
  OAI210     g0804(.A0(i_6_), .A1(i_11_), .B0(new_new_n88_), .Y(new_new_n827_));
  AOI220     g0805(.A0(new_new_n827_), .A1(new_new_n564_), .B0(new_new_n795_), .B1(new_new_n713_), .Y(new_new_n828_));
  NA2        g0806(.A(new_new_n398_), .B(new_new_n71_), .Y(new_new_n829_));
  NA3        g0807(.A(new_new_n829_), .B(new_new_n828_), .C(new_new_n605_), .Y(new_new_n830_));
  AO210      g0808(.A0(new_new_n523_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n831_));
  NA3        g0809(.A(new_new_n831_), .B(new_new_n486_), .C(new_new_n223_), .Y(new_new_n832_));
  AOI210     g0810(.A0(new_new_n451_), .A1(new_new_n449_), .B0(new_new_n563_), .Y(new_new_n833_));
  NO2        g0811(.A(new_new_n613_), .B(new_new_n105_), .Y(new_new_n834_));
  OAI210     g0812(.A0(new_new_n834_), .A1(new_new_n115_), .B0(new_new_n406_), .Y(new_new_n835_));
  INV        g0813(.A(new_new_n586_), .Y(new_new_n836_));
  NA3        g0814(.A(new_new_n836_), .B(new_new_n328_), .C(i_7_), .Y(new_new_n837_));
  NA4        g0815(.A(new_new_n837_), .B(new_new_n835_), .C(new_new_n833_), .D(new_new_n832_), .Y(new_new_n838_));
  NO4        g0816(.A(new_new_n838_), .B(new_new_n830_), .C(new_new_n826_), .D(new_new_n816_), .Y(new_new_n839_));
  NA4        g0817(.A(new_new_n839_), .B(new_new_n804_), .C(new_new_n798_), .D(new_new_n384_), .Y(mai3));
  NA2        g0818(.A(i_6_), .B(i_7_), .Y(new_new_n841_));
  NO2        g0819(.A(new_new_n841_), .B(i_0_), .Y(new_new_n842_));
  NO2        g0820(.A(i_11_), .B(new_new_n235_), .Y(new_new_n843_));
  OAI210     g0821(.A0(new_new_n842_), .A1(new_new_n290_), .B0(new_new_n843_), .Y(new_new_n844_));
  NO2        g0822(.A(new_new_n844_), .B(new_new_n198_), .Y(new_new_n845_));
  NO3        g0823(.A(new_new_n455_), .B(new_new_n93_), .C(new_new_n45_), .Y(new_new_n846_));
  OA210      g0824(.A0(new_new_n846_), .A1(new_new_n845_), .B0(new_new_n178_), .Y(new_new_n847_));
  NOi21      g0825(.An(new_new_n99_), .B(new_new_n760_), .Y(new_new_n848_));
  NA2        g0826(.A(new_new_n409_), .B(new_new_n46_), .Y(new_new_n849_));
  AN2        g0827(.A(new_new_n457_), .B(new_new_n56_), .Y(new_new_n850_));
  NO2        g0828(.A(new_new_n850_), .B(new_new_n848_), .Y(new_new_n851_));
  NO2        g0829(.A(new_new_n851_), .B(new_new_n49_), .Y(new_new_n852_));
  NO4        g0830(.A(new_new_n380_), .B(new_new_n387_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n190_), .B(new_new_n573_), .Y(new_new_n854_));
  NOi21      g0832(.An(new_new_n854_), .B(new_new_n853_), .Y(new_new_n855_));
  NA2        g0833(.A(new_new_n705_), .B(new_new_n672_), .Y(new_new_n856_));
  NA2        g0834(.A(new_new_n332_), .B(new_new_n439_), .Y(new_new_n857_));
  OAI220     g0835(.A0(new_new_n857_), .A1(new_new_n856_), .B0(new_new_n855_), .B1(new_new_n64_), .Y(new_new_n858_));
  NOi21      g0836(.An(i_5_), .B(i_9_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n859_), .B(new_new_n447_), .Y(new_new_n860_));
  BUFFER     g0838(.A(new_new_n269_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n861_), .B(new_new_n477_), .Y(new_new_n862_));
  NO3        g0840(.A(new_new_n412_), .B(new_new_n269_), .C(new_new_n74_), .Y(new_new_n863_));
  NO2        g0841(.A(new_new_n179_), .B(new_new_n151_), .Y(new_new_n864_));
  AOI210     g0842(.A0(new_new_n864_), .A1(new_new_n243_), .B0(new_new_n863_), .Y(new_new_n865_));
  OAI220     g0843(.A0(new_new_n865_), .A1(new_new_n185_), .B0(new_new_n862_), .B1(new_new_n860_), .Y(new_new_n866_));
  NO4        g0844(.A(new_new_n866_), .B(new_new_n858_), .C(new_new_n852_), .D(new_new_n847_), .Y(new_new_n867_));
  NA2        g0845(.A(new_new_n190_), .B(new_new_n24_), .Y(new_new_n868_));
  NO2        g0846(.A(new_new_n670_), .B(new_new_n594_), .Y(new_new_n869_));
  NO2        g0847(.A(new_new_n869_), .B(new_new_n868_), .Y(new_new_n870_));
  INV        g0848(.A(new_new_n870_), .Y(new_new_n871_));
  NO2        g0849(.A(new_new_n392_), .B(new_new_n291_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n872_), .B(new_new_n708_), .Y(new_new_n873_));
  NA2        g0851(.A(new_new_n574_), .B(i_0_), .Y(new_new_n874_));
  NO4        g0852(.A(new_new_n585_), .B(new_new_n221_), .C(new_new_n416_), .D(new_new_n408_), .Y(new_new_n875_));
  NA2        g0853(.A(new_new_n875_), .B(i_11_), .Y(new_new_n876_));
  AN2        g0854(.A(new_new_n99_), .B(new_new_n242_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n747_), .B(new_new_n329_), .Y(new_new_n878_));
  AOI210     g0856(.A0(new_new_n486_), .A1(new_new_n90_), .B0(new_new_n59_), .Y(new_new_n879_));
  OAI220     g0857(.A0(new_new_n879_), .A1(new_new_n878_), .B0(new_new_n656_), .B1(new_new_n542_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n253_), .B(new_new_n156_), .Y(new_new_n881_));
  NA2        g0859(.A(i_0_), .B(i_10_), .Y(new_new_n882_));
  INV        g0860(.A(new_new_n545_), .Y(new_new_n883_));
  NO4        g0861(.A(new_new_n118_), .B(new_new_n59_), .C(new_new_n665_), .D(i_5_), .Y(new_new_n884_));
  AO220      g0862(.A0(new_new_n884_), .A1(new_new_n883_), .B0(new_new_n881_), .B1(i_6_), .Y(new_new_n885_));
  AOI220     g0863(.A0(new_new_n332_), .A1(new_new_n101_), .B0(new_new_n190_), .B1(new_new_n85_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n568_), .B(i_4_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n193_), .B(new_new_n208_), .Y(new_new_n888_));
  OAI220     g0866(.A0(new_new_n888_), .A1(new_new_n878_), .B0(new_new_n887_), .B1(new_new_n886_), .Y(new_new_n889_));
  NO4        g0867(.A(new_new_n889_), .B(new_new_n885_), .C(new_new_n880_), .D(new_new_n877_), .Y(new_new_n890_));
  NA4        g0868(.A(new_new_n890_), .B(new_new_n876_), .C(new_new_n873_), .D(new_new_n871_), .Y(new_new_n891_));
  NA2        g0869(.A(i_11_), .B(i_9_), .Y(new_new_n892_));
  NO2        g0870(.A(new_new_n49_), .B(i_7_), .Y(new_new_n893_));
  NA2        g0871(.A(new_new_n397_), .B(new_new_n183_), .Y(new_new_n894_));
  NA2        g0872(.A(new_new_n894_), .B(new_new_n163_), .Y(new_new_n895_));
  NO2        g0873(.A(new_new_n892_), .B(new_new_n74_), .Y(new_new_n896_));
  NO2        g0874(.A(new_new_n179_), .B(i_0_), .Y(new_new_n897_));
  INV        g0875(.A(new_new_n897_), .Y(new_new_n898_));
  NA2        g0876(.A(new_new_n475_), .B(new_new_n229_), .Y(new_new_n899_));
  NA2        g0877(.A(new_new_n375_), .B(new_new_n42_), .Y(new_new_n900_));
  OAI220     g0878(.A0(new_new_n900_), .A1(new_new_n860_), .B0(new_new_n899_), .B1(new_new_n898_), .Y(new_new_n901_));
  NO2        g0879(.A(new_new_n901_), .B(new_new_n895_), .Y(new_new_n902_));
  NA2        g0880(.A(new_new_n655_), .B(new_new_n124_), .Y(new_new_n903_));
  NO2        g0881(.A(i_6_), .B(new_new_n903_), .Y(new_new_n904_));
  AOI210     g0882(.A0(new_new_n450_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n175_), .B(new_new_n106_), .Y(new_new_n906_));
  NOi32      g0884(.An(new_new_n905_), .Bn(new_new_n193_), .C(new_new_n906_), .Y(new_new_n907_));
  NA2        g0885(.A(new_new_n606_), .B(new_new_n329_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n908_), .B(new_new_n849_), .Y(new_new_n909_));
  NO3        g0887(.A(new_new_n909_), .B(new_new_n907_), .C(new_new_n904_), .Y(new_new_n910_));
  NOi21      g0888(.An(i_7_), .B(i_5_), .Y(new_new_n911_));
  OR2        g0889(.A(new_new_n906_), .B(new_new_n521_), .Y(new_new_n912_));
  NO3        g0890(.A(new_new_n402_), .B(new_new_n364_), .C(new_new_n360_), .Y(new_new_n913_));
  NO2        g0891(.A(new_new_n263_), .B(new_new_n318_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n724_), .B(new_new_n258_), .Y(new_new_n915_));
  AOI210     g0893(.A0(new_new_n915_), .A1(new_new_n914_), .B0(new_new_n913_), .Y(new_new_n916_));
  NA4        g0894(.A(new_new_n916_), .B(new_new_n912_), .C(new_new_n910_), .D(new_new_n902_), .Y(new_new_n917_));
  NO2        g0895(.A(new_new_n868_), .B(new_new_n238_), .Y(new_new_n918_));
  AN2        g0896(.A(new_new_n331_), .B(new_new_n329_), .Y(new_new_n919_));
  AN2        g0897(.A(new_new_n919_), .B(new_new_n864_), .Y(new_new_n920_));
  OAI210     g0898(.A0(new_new_n920_), .A1(new_new_n918_), .B0(i_10_), .Y(new_new_n921_));
  OA210      g0899(.A0(new_new_n475_), .A1(new_new_n225_), .B0(new_new_n474_), .Y(new_new_n922_));
  NA2        g0900(.A(new_new_n896_), .B(new_new_n304_), .Y(new_new_n923_));
  OAI210     g0901(.A0(i_2_), .A1(new_new_n192_), .B0(new_new_n923_), .Y(new_new_n924_));
  NA2        g0902(.A(new_new_n924_), .B(new_new_n475_), .Y(new_new_n925_));
  NO3        g0903(.A(new_new_n585_), .B(new_new_n359_), .C(new_new_n24_), .Y(new_new_n926_));
  INV        g0904(.A(new_new_n926_), .Y(new_new_n927_));
  NAi21      g0905(.An(i_9_), .B(i_5_), .Y(new_new_n928_));
  NO2        g0906(.A(new_new_n928_), .B(new_new_n402_), .Y(new_new_n929_));
  NO2        g0907(.A(new_new_n600_), .B(new_new_n108_), .Y(new_new_n930_));
  AOI220     g0908(.A0(new_new_n930_), .A1(i_0_), .B0(new_new_n929_), .B1(new_new_n623_), .Y(new_new_n931_));
  OAI220     g0909(.A0(new_new_n931_), .A1(new_new_n87_), .B0(new_new_n927_), .B1(new_new_n176_), .Y(new_new_n932_));
  NO2        g0910(.A(new_new_n932_), .B(new_new_n526_), .Y(new_new_n933_));
  NA3        g0911(.A(new_new_n933_), .B(new_new_n925_), .C(new_new_n921_), .Y(new_new_n934_));
  NO3        g0912(.A(new_new_n934_), .B(new_new_n917_), .C(new_new_n891_), .Y(new_new_n935_));
  NO2        g0913(.A(i_0_), .B(new_new_n724_), .Y(new_new_n936_));
  NA2        g0914(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n937_));
  INV        g0915(.A(new_new_n937_), .Y(new_new_n938_));
  NO3        g0916(.A(new_new_n108_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n939_));
  AO220      g0917(.A0(new_new_n939_), .A1(new_new_n938_), .B0(new_new_n936_), .B1(new_new_n178_), .Y(new_new_n940_));
  AOI210     g0918(.A0(new_new_n800_), .A1(new_new_n683_), .B0(new_new_n906_), .Y(new_new_n941_));
  AOI210     g0919(.A0(new_new_n940_), .A1(new_new_n348_), .B0(new_new_n941_), .Y(new_new_n942_));
  NA2        g0920(.A(new_new_n735_), .B(new_new_n149_), .Y(new_new_n943_));
  INV        g0921(.A(new_new_n943_), .Y(new_new_n944_));
  NA3        g0922(.A(new_new_n944_), .B(new_new_n672_), .C(new_new_n74_), .Y(new_new_n945_));
  NA3        g0923(.A(new_new_n842_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n946_));
  NA2        g0924(.A(new_new_n843_), .B(i_9_), .Y(new_new_n947_));
  AOI210     g0925(.A0(new_new_n946_), .A1(new_new_n500_), .B0(new_new_n947_), .Y(new_new_n948_));
  OAI210     g0926(.A0(new_new_n243_), .A1(i_9_), .B0(new_new_n228_), .Y(new_new_n949_));
  AOI210     g0927(.A0(new_new_n949_), .A1(new_new_n874_), .B0(new_new_n156_), .Y(new_new_n950_));
  NO2        g0928(.A(new_new_n950_), .B(new_new_n948_), .Y(new_new_n951_));
  NA3        g0929(.A(new_new_n951_), .B(new_new_n945_), .C(new_new_n942_), .Y(new_new_n952_));
  NA2        g0930(.A(new_new_n919_), .B(new_new_n377_), .Y(new_new_n953_));
  AOI210     g0931(.A0(new_new_n298_), .A1(new_new_n165_), .B0(new_new_n953_), .Y(new_new_n954_));
  NA3        g0932(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n955_));
  NA2        g0933(.A(new_new_n893_), .B(new_new_n491_), .Y(new_new_n956_));
  AOI210     g0934(.A0(new_new_n955_), .A1(new_new_n165_), .B0(new_new_n956_), .Y(new_new_n957_));
  NO2        g0935(.A(new_new_n957_), .B(new_new_n954_), .Y(new_new_n958_));
  NO3        g0936(.A(new_new_n882_), .B(new_new_n859_), .C(new_new_n195_), .Y(new_new_n959_));
  AOI220     g0937(.A0(new_new_n959_), .A1(i_11_), .B0(new_new_n569_), .B1(new_new_n76_), .Y(new_new_n960_));
  NO3        g0938(.A(new_new_n215_), .B(new_new_n387_), .C(i_0_), .Y(new_new_n961_));
  OAI210     g0939(.A0(new_new_n961_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n962_));
  INV        g0940(.A(new_new_n223_), .Y(new_new_n963_));
  OAI220     g0941(.A0(new_new_n536_), .A1(new_new_n142_), .B0(new_new_n642_), .B1(new_new_n617_), .Y(new_new_n964_));
  NA3        g0942(.A(new_new_n964_), .B(new_new_n1034_), .C(new_new_n963_), .Y(new_new_n965_));
  NA4        g0943(.A(new_new_n965_), .B(new_new_n962_), .C(new_new_n960_), .D(new_new_n958_), .Y(new_new_n966_));
  INV        g0944(.A(new_new_n112_), .Y(new_new_n967_));
  AOI220     g0945(.A0(new_new_n911_), .A1(new_new_n491_), .B0(new_new_n842_), .B1(new_new_n166_), .Y(new_new_n968_));
  NA2        g0946(.A(new_new_n351_), .B(new_new_n180_), .Y(new_new_n969_));
  OA220      g0947(.A0(new_new_n969_), .A1(new_new_n968_), .B0(new_new_n967_), .B1(i_5_), .Y(new_new_n970_));
  AOI210     g0948(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n179_), .Y(new_new_n971_));
  NA2        g0949(.A(new_new_n971_), .B(new_new_n922_), .Y(new_new_n972_));
  NA3        g0950(.A(new_new_n614_), .B(new_new_n190_), .C(new_new_n85_), .Y(new_new_n973_));
  INV        g0951(.A(new_new_n973_), .Y(new_new_n974_));
  NO3        g0952(.A(new_new_n849_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n975_));
  NA2        g0953(.A(new_new_n496_), .B(new_new_n489_), .Y(new_new_n976_));
  NO3        g0954(.A(new_new_n976_), .B(new_new_n975_), .C(new_new_n974_), .Y(new_new_n977_));
  NA3        g0955(.A(new_new_n893_), .B(new_new_n290_), .C(new_new_n228_), .Y(new_new_n978_));
  INV        g0956(.A(new_new_n978_), .Y(new_new_n979_));
  NOi31      g0957(.An(new_new_n391_), .B(new_new_n937_), .C(new_new_n238_), .Y(new_new_n980_));
  NO3        g0958(.A(new_new_n892_), .B(new_new_n223_), .C(new_new_n195_), .Y(new_new_n981_));
  NO3        g0959(.A(new_new_n981_), .B(new_new_n980_), .C(new_new_n979_), .Y(new_new_n982_));
  NA4        g0960(.A(new_new_n982_), .B(new_new_n977_), .C(new_new_n972_), .D(new_new_n970_), .Y(new_new_n983_));
  INV        g0961(.A(new_new_n616_), .Y(new_new_n984_));
  NO3        g0962(.A(new_new_n984_), .B(new_new_n559_), .C(new_new_n345_), .Y(new_new_n985_));
  INV        g0963(.A(new_new_n985_), .Y(new_new_n986_));
  NA2        g0964(.A(new_new_n794_), .B(new_new_n180_), .Y(new_new_n987_));
  NA3        g0965(.A(new_new_n101_), .B(new_new_n573_), .C(i_11_), .Y(new_new_n988_));
  NO2        g0966(.A(new_new_n988_), .B(new_new_n158_), .Y(new_new_n989_));
  INV        g0967(.A(new_new_n989_), .Y(new_new_n990_));
  NA3        g0968(.A(new_new_n990_), .B(new_new_n987_), .C(new_new_n986_), .Y(new_new_n991_));
  NO4        g0969(.A(new_new_n991_), .B(new_new_n983_), .C(new_new_n966_), .D(new_new_n952_), .Y(new_new_n992_));
  OAI210     g0970(.A0(new_new_n817_), .A1(new_new_n813_), .B0(new_new_n37_), .Y(new_new_n993_));
  NA3        g0971(.A(new_new_n905_), .B(new_new_n372_), .C(i_5_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n994_), .B(new_new_n993_), .C(new_new_n612_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n995_), .B(new_new_n211_), .Y(new_new_n996_));
  AN2        g0974(.A(new_new_n692_), .B(new_new_n373_), .Y(new_new_n997_));
  NA2        g0975(.A(new_new_n191_), .B(new_new_n193_), .Y(new_new_n998_));
  AO210      g0976(.A0(new_new_n997_), .A1(new_new_n33_), .B0(new_new_n998_), .Y(new_new_n999_));
  OAI210     g0977(.A0(new_new_n616_), .A1(new_new_n614_), .B0(new_new_n317_), .Y(new_new_n1000_));
  NAi31      g0978(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1001_));
  NO2        g0979(.A(new_new_n71_), .B(new_new_n1001_), .Y(new_new_n1002_));
  INV        g0980(.A(new_new_n1002_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n1003_), .B(new_new_n1000_), .C(new_new_n999_), .Y(new_new_n1004_));
  NO2        g0982(.A(new_new_n464_), .B(new_new_n269_), .Y(new_new_n1005_));
  NO4        g0983(.A(new_new_n231_), .B(new_new_n148_), .C(new_new_n676_), .D(new_new_n37_), .Y(new_new_n1006_));
  NO3        g0984(.A(new_new_n1006_), .B(new_new_n1005_), .C(new_new_n875_), .Y(new_new_n1007_));
  OAI210     g0985(.A0(new_new_n988_), .A1(new_new_n151_), .B0(new_new_n1007_), .Y(new_new_n1008_));
  AOI210     g0986(.A0(new_new_n1004_), .A1(new_new_n49_), .B0(new_new_n1008_), .Y(new_new_n1009_));
  AOI210     g0987(.A0(new_new_n1009_), .A1(new_new_n996_), .B0(new_new_n74_), .Y(new_new_n1010_));
  NO2        g0988(.A(new_new_n566_), .B(new_new_n383_), .Y(new_new_n1011_));
  NO2        g0989(.A(new_new_n1011_), .B(new_new_n755_), .Y(new_new_n1012_));
  NA2        g0990(.A(new_new_n263_), .B(new_new_n58_), .Y(new_new_n1013_));
  AOI220     g0991(.A0(new_new_n1013_), .A1(new_new_n77_), .B0(new_new_n346_), .B1(new_new_n255_), .Y(new_new_n1014_));
  NO2        g0992(.A(new_new_n1014_), .B(new_new_n235_), .Y(new_new_n1015_));
  NA3        g0993(.A(new_new_n99_), .B(new_new_n306_), .C(new_new_n31_), .Y(new_new_n1016_));
  INV        g0994(.A(new_new_n1016_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n1017_), .B(new_new_n1015_), .Y(new_new_n1018_));
  NA2        g0996(.A(new_new_n607_), .B(new_new_n221_), .Y(new_new_n1019_));
  OAI210     g0997(.A0(new_new_n1019_), .A1(new_new_n905_), .B0(new_new_n211_), .Y(new_new_n1020_));
  NA2        g0998(.A(new_new_n167_), .B(i_5_), .Y(new_new_n1021_));
  NO2        g0999(.A(new_new_n1020_), .B(new_new_n1021_), .Y(new_new_n1022_));
  NO4        g1000(.A(new_new_n928_), .B(new_new_n479_), .C(new_new_n252_), .D(new_new_n251_), .Y(new_new_n1023_));
  NO2        g1001(.A(new_new_n1023_), .B(new_new_n563_), .Y(new_new_n1024_));
  INV        g1002(.A(new_new_n365_), .Y(new_new_n1025_));
  AOI210     g1003(.A0(new_new_n1025_), .A1(new_new_n1024_), .B0(new_new_n41_), .Y(new_new_n1026_));
  NO2        g1004(.A(new_new_n1026_), .B(new_new_n1022_), .Y(new_new_n1027_));
  OAI210     g1005(.A0(new_new_n1018_), .A1(i_4_), .B0(new_new_n1027_), .Y(new_new_n1028_));
  NO3        g1006(.A(new_new_n1028_), .B(new_new_n1012_), .C(new_new_n1010_), .Y(new_new_n1029_));
  NA4        g1007(.A(new_new_n1029_), .B(new_new_n992_), .C(new_new_n935_), .D(new_new_n867_), .Y(mai4));
  INV        g1008(.A(new_new_n486_), .Y(new_new_n1033_));
  INV        g1009(.A(i_3_), .Y(new_new_n1034_));
endmodule


