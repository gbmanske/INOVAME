library verilog;
use verilog.vl_types.all;
entity tb_mac is
end tb_mac;
