//Benchmark atmr_9sym_175_0.0313

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n172_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  NA2        o002(.A(i_4_), .B(ori_ori_n12_), .Y(ori_ori_n13_));
  INV        o003(.A(i_5_), .Y(ori_ori_n14_));
  NOi21      o004(.An(i_3_), .B(i_7_), .Y(ori_ori_n15_));
  NA3        o005(.A(ori_ori_n15_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n16_));
  INV        o006(.A(i_0_), .Y(ori_ori_n17_));
  NOi21      o007(.An(i_1_), .B(i_3_), .Y(ori_ori_n18_));
  NO2        o008(.A(ori_ori_n16_), .B(ori_ori_n13_), .Y(ori_ori_n19_));
  INV        o009(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o010(.A(i_0_), .B(ori_ori_n20_), .Y(ori_ori_n21_));
  INV        o011(.A(i_7_), .Y(ori_ori_n22_));
  NA3        o012(.A(i_6_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n23_));
  NOi21      o013(.An(i_8_), .B(i_6_), .Y(ori_ori_n24_));
  NOi21      o014(.An(i_1_), .B(i_8_), .Y(ori_ori_n25_));
  AOI220     o015(.A0(ori_ori_n25_), .A1(i_2_), .B0(ori_ori_n24_), .B1(i_5_), .Y(ori_ori_n26_));
  AOI210     o016(.A0(ori_ori_n26_), .A1(ori_ori_n23_), .B0(ori_ori_n21_), .Y(ori_ori_n27_));
  AOI210     o017(.A0(ori_ori_n27_), .A1(ori_ori_n11_), .B0(ori_ori_n19_), .Y(ori_ori_n28_));
  NA2        o018(.A(i_0_), .B(ori_ori_n14_), .Y(ori_ori_n29_));
  NA2        o019(.A(ori_ori_n17_), .B(i_5_), .Y(ori_ori_n30_));
  NO2        o020(.A(i_2_), .B(i_4_), .Y(ori_ori_n31_));
  NA3        o021(.A(ori_ori_n31_), .B(i_6_), .C(i_8_), .Y(ori_ori_n32_));
  AOI210     o022(.A0(ori_ori_n30_), .A1(ori_ori_n29_), .B0(ori_ori_n32_), .Y(ori_ori_n33_));
  INV        o023(.A(i_2_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_5_), .B(i_0_), .Y(ori_ori_n35_));
  NOi21      o025(.An(i_6_), .B(i_8_), .Y(ori_ori_n36_));
  NOi21      o026(.An(i_7_), .B(i_1_), .Y(ori_ori_n37_));
  NOi21      o027(.An(i_5_), .B(i_6_), .Y(ori_ori_n38_));
  AOI220     o028(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n36_), .B1(ori_ori_n35_), .Y(ori_ori_n39_));
  NO3        o029(.A(ori_ori_n39_), .B(ori_ori_n34_), .C(i_4_), .Y(ori_ori_n40_));
  NOi21      o030(.An(i_0_), .B(i_4_), .Y(ori_ori_n41_));
  XO2        o031(.A(i_1_), .B(i_3_), .Y(ori_ori_n42_));
  NOi21      o032(.An(i_7_), .B(i_5_), .Y(ori_ori_n43_));
  AN3        o033(.A(ori_ori_n43_), .B(ori_ori_n42_), .C(ori_ori_n41_), .Y(ori_ori_n44_));
  INV        o034(.A(i_1_), .Y(ori_ori_n45_));
  NOi21      o035(.An(i_3_), .B(i_0_), .Y(ori_ori_n46_));
  NA2        o036(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o037(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n48_));
  NO4        o038(.A(ori_ori_n48_), .B(ori_ori_n44_), .C(ori_ori_n40_), .D(ori_ori_n33_), .Y(ori_ori_n49_));
  NOi21      o039(.An(i_4_), .B(i_0_), .Y(ori_ori_n50_));
  NO2        o040(.A(ori_ori_n24_), .B(ori_ori_n15_), .Y(ori_ori_n51_));
  NA2        o041(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n52_));
  NOi21      o042(.An(i_2_), .B(i_8_), .Y(ori_ori_n53_));
  NO2        o043(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n54_));
  NO3        o044(.A(ori_ori_n54_), .B(ori_ori_n52_), .C(ori_ori_n51_), .Y(ori_ori_n55_));
  INV        o045(.A(ori_ori_n55_), .Y(ori_ori_n56_));
  NOi31      o046(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n57_));
  NA2        o047(.A(ori_ori_n57_), .B(i_0_), .Y(ori_ori_n58_));
  NOi21      o048(.An(i_4_), .B(i_3_), .Y(ori_ori_n59_));
  NOi21      o049(.An(i_1_), .B(i_4_), .Y(ori_ori_n60_));
  OAI210     o050(.A0(ori_ori_n60_), .A1(ori_ori_n59_), .B0(ori_ori_n53_), .Y(ori_ori_n61_));
  NA2        o051(.A(ori_ori_n61_), .B(ori_ori_n58_), .Y(ori_ori_n62_));
  AN2        o052(.A(i_8_), .B(i_7_), .Y(ori_ori_n63_));
  INV        o053(.A(ori_ori_n63_), .Y(ori_ori_n64_));
  NOi21      o054(.An(i_8_), .B(i_7_), .Y(ori_ori_n65_));
  NA3        o055(.A(ori_ori_n65_), .B(ori_ori_n59_), .C(i_6_), .Y(ori_ori_n66_));
  OAI210     o056(.A0(ori_ori_n64_), .A1(ori_ori_n52_), .B0(ori_ori_n66_), .Y(ori_ori_n67_));
  AOI220     o057(.A0(ori_ori_n67_), .A1(ori_ori_n34_), .B0(ori_ori_n62_), .B1(ori_ori_n38_), .Y(ori_ori_n68_));
  NA4        o058(.A(ori_ori_n68_), .B(ori_ori_n56_), .C(ori_ori_n49_), .D(ori_ori_n28_), .Y(ori_ori_n69_));
  NA2        o059(.A(i_8_), .B(i_7_), .Y(ori_ori_n70_));
  NO2        o060(.A(ori_ori_n70_), .B(i_1_), .Y(ori_ori_n71_));
  NA2        o061(.A(i_8_), .B(ori_ori_n22_), .Y(ori_ori_n72_));
  AOI220     o062(.A0(ori_ori_n46_), .A1(i_1_), .B0(ori_ori_n42_), .B1(i_2_), .Y(ori_ori_n73_));
  NOi21      o063(.An(i_1_), .B(i_2_), .Y(ori_ori_n74_));
  NO2        o064(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n75_));
  OAI210     o065(.A0(ori_ori_n75_), .A1(ori_ori_n71_), .B0(ori_ori_n14_), .Y(ori_ori_n76_));
  NA3        o066(.A(ori_ori_n65_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n77_));
  NA2        o067(.A(ori_ori_n25_), .B(ori_ori_n14_), .Y(ori_ori_n78_));
  NA2        o068(.A(ori_ori_n78_), .B(ori_ori_n77_), .Y(ori_ori_n79_));
  NA2        o069(.A(ori_ori_n18_), .B(i_6_), .Y(ori_ori_n80_));
  INV        o070(.A(ori_ori_n80_), .Y(ori_ori_n81_));
  INV        o071(.A(i_0_), .Y(ori_ori_n82_));
  AOI220     o072(.A0(ori_ori_n82_), .A1(ori_ori_n81_), .B0(ori_ori_n79_), .B1(ori_ori_n59_), .Y(ori_ori_n83_));
  NA2        o073(.A(ori_ori_n83_), .B(ori_ori_n76_), .Y(ori_ori_n84_));
  NA2        o074(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n85_));
  NOi21      o075(.An(i_7_), .B(i_8_), .Y(ori_ori_n86_));
  NOi21      o076(.An(i_6_), .B(i_5_), .Y(ori_ori_n87_));
  AOI210     o077(.A0(ori_ori_n86_), .A1(ori_ori_n12_), .B0(ori_ori_n87_), .Y(ori_ori_n88_));
  OAI210     o078(.A0(ori_ori_n88_), .A1(ori_ori_n11_), .B0(ori_ori_n85_), .Y(ori_ori_n89_));
  NA2        o079(.A(ori_ori_n89_), .B(ori_ori_n74_), .Y(ori_ori_n90_));
  AOI220     o080(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n18_), .B1(ori_ori_n34_), .Y(ori_ori_n91_));
  NA3        o081(.A(ori_ori_n20_), .B(i_5_), .C(i_7_), .Y(ori_ori_n92_));
  NO2        o082(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  INV        o083(.A(ori_ori_n93_), .Y(ori_ori_n94_));
  NA3        o084(.A(ori_ori_n65_), .B(ori_ori_n34_), .C(i_3_), .Y(ori_ori_n95_));
  NA2        o085(.A(ori_ori_n45_), .B(i_6_), .Y(ori_ori_n96_));
  AOI210     o086(.A0(ori_ori_n96_), .A1(ori_ori_n21_), .B0(ori_ori_n95_), .Y(ori_ori_n97_));
  NOi21      o087(.An(i_2_), .B(i_1_), .Y(ori_ori_n98_));
  AN3        o088(.A(ori_ori_n86_), .B(ori_ori_n98_), .C(ori_ori_n50_), .Y(ori_ori_n99_));
  NAi21      o089(.An(i_6_), .B(i_0_), .Y(ori_ori_n100_));
  NA3        o090(.A(ori_ori_n60_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n101_));
  NOi21      o091(.An(i_4_), .B(i_6_), .Y(ori_ori_n102_));
  NOi21      o092(.An(i_5_), .B(i_3_), .Y(ori_ori_n103_));
  NA3        o093(.A(ori_ori_n103_), .B(ori_ori_n74_), .C(ori_ori_n102_), .Y(ori_ori_n104_));
  OAI210     o094(.A0(ori_ori_n101_), .A1(ori_ori_n100_), .B0(ori_ori_n104_), .Y(ori_ori_n105_));
  NA2        o095(.A(ori_ori_n74_), .B(ori_ori_n36_), .Y(ori_ori_n106_));
  NO3        o096(.A(ori_ori_n105_), .B(ori_ori_n99_), .C(ori_ori_n97_), .Y(ori_ori_n107_));
  NOi21      o097(.An(i_6_), .B(i_1_), .Y(ori_ori_n108_));
  AOI220     o098(.A0(ori_ori_n108_), .A1(i_7_), .B0(ori_ori_n24_), .B1(i_5_), .Y(ori_ori_n109_));
  NOi31      o099(.An(ori_ori_n50_), .B(ori_ori_n109_), .C(i_2_), .Y(ori_ori_n110_));
  NA2        o100(.A(ori_ori_n65_), .B(ori_ori_n12_), .Y(ori_ori_n111_));
  NA2        o101(.A(ori_ori_n36_), .B(ori_ori_n14_), .Y(ori_ori_n112_));
  NOi21      o102(.An(i_3_), .B(i_1_), .Y(ori_ori_n113_));
  NA2        o103(.A(ori_ori_n113_), .B(i_4_), .Y(ori_ori_n114_));
  AOI210     o104(.A0(ori_ori_n112_), .A1(ori_ori_n111_), .B0(ori_ori_n114_), .Y(ori_ori_n115_));
  NOi31      o105(.An(ori_ori_n46_), .B(i_5_), .C(ori_ori_n34_), .Y(ori_ori_n116_));
  NO3        o106(.A(ori_ori_n116_), .B(ori_ori_n115_), .C(ori_ori_n110_), .Y(ori_ori_n117_));
  NA4        o107(.A(ori_ori_n117_), .B(ori_ori_n107_), .C(ori_ori_n94_), .D(ori_ori_n90_), .Y(ori_ori_n118_));
  NOi31      o108(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n119_));
  NOi31      o109(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n120_));
  OAI210     o110(.A0(ori_ori_n120_), .A1(ori_ori_n119_), .B0(i_7_), .Y(ori_ori_n121_));
  NA2        o111(.A(ori_ori_n36_), .B(ori_ori_n14_), .Y(ori_ori_n122_));
  NA3        o112(.A(ori_ori_n122_), .B(ori_ori_n121_), .C(ori_ori_n106_), .Y(ori_ori_n123_));
  NA2        o113(.A(ori_ori_n123_), .B(ori_ori_n41_), .Y(ori_ori_n124_));
  NA2        o114(.A(ori_ori_n59_), .B(ori_ori_n37_), .Y(ori_ori_n125_));
  AOI210     o115(.A0(ori_ori_n125_), .A1(ori_ori_n77_), .B0(ori_ori_n30_), .Y(ori_ori_n126_));
  NA3        o116(.A(ori_ori_n63_), .B(ori_ori_n17_), .C(ori_ori_n12_), .Y(ori_ori_n127_));
  NAi31      o117(.An(ori_ori_n100_), .B(ori_ori_n86_), .C(ori_ori_n98_), .Y(ori_ori_n128_));
  NA3        o118(.A(ori_ori_n65_), .B(ori_ori_n57_), .C(i_6_), .Y(ori_ori_n129_));
  NA3        o119(.A(ori_ori_n129_), .B(ori_ori_n128_), .C(ori_ori_n127_), .Y(ori_ori_n130_));
  NOi21      o120(.An(i_0_), .B(i_2_), .Y(ori_ori_n131_));
  NA3        o121(.A(ori_ori_n131_), .B(ori_ori_n37_), .C(ori_ori_n102_), .Y(ori_ori_n132_));
  NOi32      o122(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n133_));
  NA2        o123(.A(ori_ori_n133_), .B(ori_ori_n119_), .Y(ori_ori_n134_));
  NA3        o124(.A(ori_ori_n131_), .B(ori_ori_n59_), .C(ori_ori_n36_), .Y(ori_ori_n135_));
  NA3        o125(.A(ori_ori_n135_), .B(ori_ori_n134_), .C(ori_ori_n132_), .Y(ori_ori_n136_));
  NA4        o126(.A(ori_ori_n57_), .B(i_6_), .C(ori_ori_n14_), .D(i_7_), .Y(ori_ori_n137_));
  NA4        o127(.A(ori_ori_n60_), .B(ori_ori_n46_), .C(i_5_), .D(ori_ori_n22_), .Y(ori_ori_n138_));
  NA2        o128(.A(ori_ori_n138_), .B(ori_ori_n137_), .Y(ori_ori_n139_));
  NO4        o129(.A(ori_ori_n139_), .B(ori_ori_n136_), .C(ori_ori_n130_), .D(ori_ori_n126_), .Y(ori_ori_n140_));
  NOi21      o130(.An(i_5_), .B(i_2_), .Y(ori_ori_n141_));
  AOI220     o131(.A0(ori_ori_n141_), .A1(ori_ori_n86_), .B0(ori_ori_n63_), .B1(ori_ori_n31_), .Y(ori_ori_n142_));
  NO2        o132(.A(ori_ori_n142_), .B(ori_ori_n96_), .Y(ori_ori_n143_));
  NO4        o133(.A(i_2_), .B(ori_ori_n20_), .C(ori_ori_n11_), .D(ori_ori_n14_), .Y(ori_ori_n144_));
  NA2        o134(.A(i_2_), .B(i_4_), .Y(ori_ori_n145_));
  INV        o135(.A(ori_ori_n145_), .Y(ori_ori_n146_));
  NO2        o136(.A(i_8_), .B(i_7_), .Y(ori_ori_n147_));
  OA210      o137(.A0(ori_ori_n146_), .A1(ori_ori_n144_), .B0(ori_ori_n147_), .Y(ori_ori_n148_));
  NA4        o138(.A(ori_ori_n113_), .B(i_0_), .C(i_5_), .D(ori_ori_n22_), .Y(ori_ori_n149_));
  NO2        o139(.A(ori_ori_n149_), .B(i_4_), .Y(ori_ori_n150_));
  NO3        o140(.A(ori_ori_n150_), .B(ori_ori_n148_), .C(ori_ori_n143_), .Y(ori_ori_n151_));
  NA2        o141(.A(ori_ori_n86_), .B(ori_ori_n12_), .Y(ori_ori_n152_));
  NA3        o142(.A(i_2_), .B(i_1_), .C(ori_ori_n14_), .Y(ori_ori_n153_));
  NA2        o143(.A(ori_ori_n50_), .B(i_3_), .Y(ori_ori_n154_));
  AOI210     o144(.A0(ori_ori_n154_), .A1(ori_ori_n153_), .B0(ori_ori_n152_), .Y(ori_ori_n155_));
  NA3        o145(.A(ori_ori_n131_), .B(ori_ori_n65_), .C(ori_ori_n102_), .Y(ori_ori_n156_));
  OAI210     o146(.A0(ori_ori_n95_), .A1(ori_ori_n30_), .B0(ori_ori_n156_), .Y(ori_ori_n157_));
  NA4        o147(.A(ori_ori_n103_), .B(ori_ori_n63_), .C(ori_ori_n45_), .D(ori_ori_n20_), .Y(ori_ori_n158_));
  NA2        o148(.A(ori_ori_n53_), .B(ori_ori_n15_), .Y(ori_ori_n159_));
  NOi31      o149(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n160_));
  NA2        o150(.A(ori_ori_n133_), .B(ori_ori_n160_), .Y(ori_ori_n161_));
  NA3        o151(.A(ori_ori_n161_), .B(ori_ori_n159_), .C(ori_ori_n158_), .Y(ori_ori_n162_));
  NO3        o152(.A(ori_ori_n162_), .B(ori_ori_n157_), .C(ori_ori_n155_), .Y(ori_ori_n163_));
  NA4        o153(.A(ori_ori_n163_), .B(ori_ori_n151_), .C(ori_ori_n140_), .D(ori_ori_n124_), .Y(ori_ori_n164_));
  OR4        o154(.A(ori_ori_n164_), .B(ori_ori_n118_), .C(ori_ori_n84_), .D(ori_ori_n69_), .Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  INV        m005(.A(i_0_), .Y(mai_mai_n16_));
  NOi21      m006(.An(i_1_), .B(i_3_), .Y(mai_mai_n17_));
  NA3        m007(.A(mai_mai_n17_), .B(mai_mai_n16_), .C(i_2_), .Y(mai_mai_n18_));
  NO2        m008(.A(mai_mai_n18_), .B(mai_mai_n13_), .Y(mai_mai_n19_));
  INV        m009(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m010(.A(i_0_), .B(mai_mai_n20_), .Y(mai_mai_n21_));
  INV        m011(.A(i_7_), .Y(mai_mai_n22_));
  NA3        m012(.A(i_6_), .B(i_5_), .C(mai_mai_n22_), .Y(mai_mai_n23_));
  NOi21      m013(.An(i_8_), .B(i_6_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_1_), .B(i_8_), .Y(mai_mai_n25_));
  AOI220     m015(.A0(mai_mai_n25_), .A1(i_2_), .B0(mai_mai_n24_), .B1(i_5_), .Y(mai_mai_n26_));
  AOI210     m016(.A0(mai_mai_n26_), .A1(mai_mai_n23_), .B0(mai_mai_n21_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n27_), .A1(mai_mai_n11_), .B0(mai_mai_n19_), .Y(mai_mai_n28_));
  NA2        m018(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n29_));
  NA2        m019(.A(mai_mai_n16_), .B(i_5_), .Y(mai_mai_n30_));
  NO2        m020(.A(i_2_), .B(i_4_), .Y(mai_mai_n31_));
  NA3        m021(.A(mai_mai_n31_), .B(i_6_), .C(i_8_), .Y(mai_mai_n32_));
  AOI210     m022(.A0(mai_mai_n30_), .A1(mai_mai_n29_), .B0(mai_mai_n32_), .Y(mai_mai_n33_));
  INV        m023(.A(i_2_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_5_), .B(i_0_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_6_), .B(i_8_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_7_), .B(i_1_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_5_), .B(i_6_), .Y(mai_mai_n38_));
  AOI220     m028(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n36_), .B1(mai_mai_n35_), .Y(mai_mai_n39_));
  NO3        m029(.A(mai_mai_n39_), .B(mai_mai_n34_), .C(i_4_), .Y(mai_mai_n40_));
  NOi21      m030(.An(i_0_), .B(i_4_), .Y(mai_mai_n41_));
  XO2        m031(.A(i_1_), .B(i_3_), .Y(mai_mai_n42_));
  NOi21      m032(.An(i_7_), .B(i_5_), .Y(mai_mai_n43_));
  AN3        m033(.A(mai_mai_n43_), .B(mai_mai_n42_), .C(mai_mai_n41_), .Y(mai_mai_n44_));
  INV        m034(.A(i_1_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_3_), .B(i_0_), .Y(mai_mai_n46_));
  NO3        m036(.A(mai_mai_n44_), .B(mai_mai_n40_), .C(mai_mai_n33_), .Y(mai_mai_n47_));
  INV        m037(.A(i_8_), .Y(mai_mai_n48_));
  NA2        m038(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n49_));
  NO4        m039(.A(mai_mai_n49_), .B(mai_mai_n29_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n50_));
  NOi21      m040(.An(i_4_), .B(i_0_), .Y(mai_mai_n51_));
  AOI210     m041(.A0(mai_mai_n51_), .A1(mai_mai_n24_), .B0(mai_mai_n15_), .Y(mai_mai_n52_));
  NA2        m042(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n53_));
  NOi21      m043(.An(i_2_), .B(i_8_), .Y(mai_mai_n54_));
  NO3        m044(.A(mai_mai_n54_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai_mai_n55_));
  NO3        m045(.A(mai_mai_n55_), .B(mai_mai_n53_), .C(mai_mai_n52_), .Y(mai_mai_n56_));
  NO2        m046(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n57_));
  NOi31      m047(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n58_));
  NA2        m048(.A(mai_mai_n58_), .B(i_0_), .Y(mai_mai_n59_));
  NOi21      m049(.An(i_4_), .B(i_3_), .Y(mai_mai_n60_));
  NOi21      m050(.An(i_1_), .B(i_4_), .Y(mai_mai_n61_));
  OAI210     m051(.A0(mai_mai_n61_), .A1(mai_mai_n60_), .B0(mai_mai_n54_), .Y(mai_mai_n62_));
  NA2        m052(.A(mai_mai_n62_), .B(mai_mai_n59_), .Y(mai_mai_n63_));
  AN2        m053(.A(i_8_), .B(i_7_), .Y(mai_mai_n64_));
  NA2        m054(.A(mai_mai_n64_), .B(mai_mai_n12_), .Y(mai_mai_n65_));
  NOi21      m055(.An(i_8_), .B(i_7_), .Y(mai_mai_n66_));
  NA3        m056(.A(mai_mai_n66_), .B(mai_mai_n60_), .C(i_6_), .Y(mai_mai_n67_));
  OAI210     m057(.A0(mai_mai_n65_), .A1(mai_mai_n53_), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m058(.A0(mai_mai_n68_), .A1(mai_mai_n34_), .B0(mai_mai_n63_), .B1(mai_mai_n38_), .Y(mai_mai_n69_));
  NA4        m059(.A(mai_mai_n69_), .B(mai_mai_n57_), .C(mai_mai_n47_), .D(mai_mai_n28_), .Y(mai_mai_n70_));
  NA2        m060(.A(i_8_), .B(mai_mai_n22_), .Y(mai_mai_n71_));
  AOI220     m061(.A0(mai_mai_n46_), .A1(i_1_), .B0(mai_mai_n42_), .B1(i_2_), .Y(mai_mai_n72_));
  NOi21      m062(.An(i_1_), .B(i_2_), .Y(mai_mai_n73_));
  NO2        m063(.A(mai_mai_n72_), .B(mai_mai_n71_), .Y(mai_mai_n74_));
  NA2        m064(.A(mai_mai_n74_), .B(mai_mai_n14_), .Y(mai_mai_n75_));
  NA2        m065(.A(mai_mai_n66_), .B(i_2_), .Y(mai_mai_n76_));
  NA3        m066(.A(mai_mai_n25_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n77_));
  INV        m067(.A(mai_mai_n77_), .Y(mai_mai_n78_));
  NOi32      m068(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n79_));
  NA2        m069(.A(mai_mai_n79_), .B(i_3_), .Y(mai_mai_n80_));
  NA3        m070(.A(mai_mai_n17_), .B(i_2_), .C(i_6_), .Y(mai_mai_n81_));
  NA2        m071(.A(mai_mai_n81_), .B(mai_mai_n80_), .Y(mai_mai_n82_));
  NO2        m072(.A(i_0_), .B(i_4_), .Y(mai_mai_n83_));
  AOI220     m073(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n78_), .B1(mai_mai_n60_), .Y(mai_mai_n84_));
  NA2        m074(.A(mai_mai_n84_), .B(mai_mai_n75_), .Y(mai_mai_n85_));
  NAi21      m075(.An(i_3_), .B(i_6_), .Y(mai_mai_n86_));
  NO3        m076(.A(mai_mai_n86_), .B(i_0_), .C(mai_mai_n48_), .Y(mai_mai_n87_));
  NA2        m077(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n88_));
  NOi21      m078(.An(i_7_), .B(i_8_), .Y(mai_mai_n89_));
  NOi31      m079(.An(i_6_), .B(i_5_), .C(i_7_), .Y(mai_mai_n90_));
  AOI210     m080(.A0(mai_mai_n89_), .A1(mai_mai_n12_), .B0(mai_mai_n90_), .Y(mai_mai_n91_));
  OAI210     m081(.A0(mai_mai_n91_), .A1(mai_mai_n11_), .B0(mai_mai_n88_), .Y(mai_mai_n92_));
  OAI210     m082(.A0(mai_mai_n92_), .A1(mai_mai_n87_), .B0(mai_mai_n73_), .Y(mai_mai_n93_));
  NA3        m083(.A(mai_mai_n24_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n94_));
  AOI210     m084(.A0(mai_mai_n21_), .A1(mai_mai_n49_), .B0(mai_mai_n94_), .Y(mai_mai_n95_));
  AOI220     m085(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n17_), .B1(mai_mai_n34_), .Y(mai_mai_n96_));
  NA3        m086(.A(mai_mai_n20_), .B(i_5_), .C(i_7_), .Y(mai_mai_n97_));
  NO2        m087(.A(mai_mai_n97_), .B(mai_mai_n96_), .Y(mai_mai_n98_));
  NO2        m088(.A(mai_mai_n98_), .B(mai_mai_n95_), .Y(mai_mai_n99_));
  NA3        m089(.A(mai_mai_n66_), .B(mai_mai_n34_), .C(i_3_), .Y(mai_mai_n100_));
  NA2        m090(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n101_));
  AOI210     m091(.A0(mai_mai_n101_), .A1(mai_mai_n21_), .B0(mai_mai_n100_), .Y(mai_mai_n102_));
  NAi21      m092(.An(i_6_), .B(i_0_), .Y(mai_mai_n103_));
  NA3        m093(.A(mai_mai_n61_), .B(i_5_), .C(mai_mai_n22_), .Y(mai_mai_n104_));
  NOi21      m094(.An(i_4_), .B(i_6_), .Y(mai_mai_n105_));
  NOi21      m095(.An(i_5_), .B(i_3_), .Y(mai_mai_n106_));
  NA3        m096(.A(mai_mai_n106_), .B(mai_mai_n73_), .C(mai_mai_n105_), .Y(mai_mai_n107_));
  OAI210     m097(.A0(mai_mai_n104_), .A1(mai_mai_n103_), .B0(mai_mai_n107_), .Y(mai_mai_n108_));
  NA2        m098(.A(mai_mai_n73_), .B(mai_mai_n36_), .Y(mai_mai_n109_));
  NOi21      m099(.An(mai_mai_n43_), .B(mai_mai_n109_), .Y(mai_mai_n110_));
  NO3        m100(.A(mai_mai_n110_), .B(mai_mai_n108_), .C(mai_mai_n102_), .Y(mai_mai_n111_));
  NOi21      m101(.An(i_6_), .B(i_1_), .Y(mai_mai_n112_));
  AOI210     m102(.A0(mai_mai_n112_), .A1(i_7_), .B0(mai_mai_n24_), .Y(mai_mai_n113_));
  NOi31      m103(.An(mai_mai_n51_), .B(mai_mai_n113_), .C(i_2_), .Y(mai_mai_n114_));
  NOi21      m104(.An(i_3_), .B(i_1_), .Y(mai_mai_n115_));
  NA2        m105(.A(mai_mai_n115_), .B(i_4_), .Y(mai_mai_n116_));
  NO2        m106(.A(i_6_), .B(mai_mai_n116_), .Y(mai_mai_n117_));
  NA2        m107(.A(mai_mai_n89_), .B(mai_mai_n14_), .Y(mai_mai_n118_));
  NOi31      m108(.An(mai_mai_n46_), .B(mai_mai_n118_), .C(mai_mai_n34_), .Y(mai_mai_n119_));
  NO3        m109(.A(mai_mai_n119_), .B(mai_mai_n117_), .C(mai_mai_n114_), .Y(mai_mai_n120_));
  NA4        m110(.A(mai_mai_n120_), .B(mai_mai_n111_), .C(mai_mai_n99_), .D(mai_mai_n93_), .Y(mai_mai_n121_));
  NA2        m111(.A(mai_mai_n54_), .B(mai_mai_n15_), .Y(mai_mai_n122_));
  NOi31      m112(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n123_));
  NA2        m113(.A(mai_mai_n123_), .B(i_7_), .Y(mai_mai_n124_));
  NA3        m114(.A(mai_mai_n36_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n125_));
  NA4        m115(.A(mai_mai_n125_), .B(mai_mai_n124_), .C(mai_mai_n122_), .D(mai_mai_n109_), .Y(mai_mai_n126_));
  NA2        m116(.A(mai_mai_n126_), .B(mai_mai_n41_), .Y(mai_mai_n127_));
  NA2        m117(.A(mai_mai_n60_), .B(mai_mai_n37_), .Y(mai_mai_n128_));
  AOI210     m118(.A0(mai_mai_n128_), .A1(mai_mai_n76_), .B0(mai_mai_n30_), .Y(mai_mai_n129_));
  NA3        m119(.A(mai_mai_n66_), .B(mai_mai_n58_), .C(i_6_), .Y(mai_mai_n130_));
  INV        m120(.A(mai_mai_n130_), .Y(mai_mai_n131_));
  NA3        m121(.A(mai_mai_n51_), .B(mai_mai_n43_), .C(mai_mai_n17_), .Y(mai_mai_n132_));
  NA2        m122(.A(mai_mai_n60_), .B(mai_mai_n36_), .Y(mai_mai_n133_));
  NA2        m123(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n134_));
  NA3        m124(.A(mai_mai_n58_), .B(mai_mai_n14_), .C(i_7_), .Y(mai_mai_n135_));
  NA4        m125(.A(mai_mai_n61_), .B(mai_mai_n38_), .C(mai_mai_n16_), .D(i_8_), .Y(mai_mai_n136_));
  NA2        m126(.A(mai_mai_n136_), .B(mai_mai_n135_), .Y(mai_mai_n137_));
  NO4        m127(.A(mai_mai_n137_), .B(mai_mai_n134_), .C(mai_mai_n131_), .D(mai_mai_n129_), .Y(mai_mai_n138_));
  AOI210     m128(.A0(mai_mai_n64_), .A1(mai_mai_n31_), .B0(mai_mai_n89_), .Y(mai_mai_n139_));
  AOI210     m129(.A0(mai_mai_n139_), .A1(mai_mai_n122_), .B0(mai_mai_n101_), .Y(mai_mai_n140_));
  NO3        m130(.A(i_2_), .B(mai_mai_n20_), .C(mai_mai_n11_), .Y(mai_mai_n141_));
  NA2        m131(.A(i_2_), .B(i_4_), .Y(mai_mai_n142_));
  NO2        m132(.A(mai_mai_n103_), .B(mai_mai_n142_), .Y(mai_mai_n143_));
  NO2        m133(.A(i_8_), .B(i_7_), .Y(mai_mai_n144_));
  OA210      m134(.A0(mai_mai_n143_), .A1(mai_mai_n141_), .B0(mai_mai_n144_), .Y(mai_mai_n145_));
  NA3        m135(.A(mai_mai_n115_), .B(i_0_), .C(mai_mai_n22_), .Y(mai_mai_n146_));
  NO2        m136(.A(mai_mai_n146_), .B(i_4_), .Y(mai_mai_n147_));
  NO3        m137(.A(mai_mai_n147_), .B(mai_mai_n145_), .C(mai_mai_n140_), .Y(mai_mai_n148_));
  NA2        m138(.A(mai_mai_n89_), .B(mai_mai_n12_), .Y(mai_mai_n149_));
  NA2        m139(.A(i_2_), .B(mai_mai_n14_), .Y(mai_mai_n150_));
  NA2        m140(.A(mai_mai_n51_), .B(i_3_), .Y(mai_mai_n151_));
  AOI210     m141(.A0(mai_mai_n151_), .A1(mai_mai_n150_), .B0(mai_mai_n149_), .Y(mai_mai_n152_));
  NA2        m142(.A(mai_mai_n66_), .B(mai_mai_n105_), .Y(mai_mai_n153_));
  INV        m143(.A(mai_mai_n153_), .Y(mai_mai_n154_));
  NA4        m144(.A(mai_mai_n106_), .B(mai_mai_n64_), .C(mai_mai_n45_), .D(mai_mai_n20_), .Y(mai_mai_n155_));
  NA2        m145(.A(mai_mai_n35_), .B(mai_mai_n15_), .Y(mai_mai_n156_));
  NOi31      m146(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n157_));
  OAI210     m147(.A0(i_4_), .A1(mai_mai_n79_), .B0(mai_mai_n157_), .Y(mai_mai_n158_));
  NA3        m148(.A(mai_mai_n158_), .B(mai_mai_n156_), .C(mai_mai_n155_), .Y(mai_mai_n159_));
  NO3        m149(.A(mai_mai_n159_), .B(mai_mai_n154_), .C(mai_mai_n152_), .Y(mai_mai_n160_));
  NA4        m150(.A(mai_mai_n160_), .B(mai_mai_n148_), .C(mai_mai_n138_), .D(mai_mai_n127_), .Y(mai_mai_n161_));
  OR4        m151(.A(mai_mai_n161_), .B(mai_mai_n121_), .C(mai_mai_n85_), .D(mai_mai_n70_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NA3        u013(.A(i_6_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n24_));
  NOi21      u014(.An(i_8_), .B(i_6_), .Y(men_men_n25_));
  AOI210     u015(.A0(men_men_n172_), .A1(men_men_n24_), .B0(men_men_n22_), .Y(men_men_n26_));
  AOI210     u016(.A0(men_men_n26_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n27_));
  NA2        u017(.A(men_men_n17_), .B(i_5_), .Y(men_men_n28_));
  NO2        u018(.A(i_2_), .B(i_4_), .Y(men_men_n29_));
  NA3        u019(.A(men_men_n29_), .B(i_6_), .C(i_8_), .Y(men_men_n30_));
  INV        u020(.A(men_men_n30_), .Y(men_men_n31_));
  INV        u021(.A(i_2_), .Y(men_men_n32_));
  NOi21      u022(.An(i_5_), .B(i_0_), .Y(men_men_n33_));
  NOi21      u023(.An(i_6_), .B(i_8_), .Y(men_men_n34_));
  NOi21      u024(.An(i_7_), .B(i_1_), .Y(men_men_n35_));
  NOi21      u025(.An(i_5_), .B(i_6_), .Y(men_men_n36_));
  NOi21      u026(.An(i_0_), .B(i_4_), .Y(men_men_n37_));
  XO2        u027(.A(i_1_), .B(i_3_), .Y(men_men_n38_));
  NOi21      u028(.An(i_7_), .B(i_5_), .Y(men_men_n39_));
  AN3        u029(.A(men_men_n39_), .B(men_men_n38_), .C(men_men_n37_), .Y(men_men_n40_));
  INV        u030(.A(i_1_), .Y(men_men_n41_));
  NOi21      u031(.An(i_3_), .B(i_0_), .Y(men_men_n42_));
  NA2        u032(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA3        u033(.A(i_6_), .B(men_men_n14_), .C(i_7_), .Y(men_men_n44_));
  AOI210     u034(.A0(men_men_n44_), .A1(men_men_n24_), .B0(men_men_n43_), .Y(men_men_n45_));
  NO3        u035(.A(men_men_n45_), .B(men_men_n40_), .C(men_men_n31_), .Y(men_men_n46_));
  NOi21      u036(.An(i_4_), .B(i_0_), .Y(men_men_n47_));
  AOI210     u037(.A0(men_men_n47_), .A1(men_men_n25_), .B0(men_men_n15_), .Y(men_men_n48_));
  NA2        u038(.A(i_1_), .B(men_men_n14_), .Y(men_men_n49_));
  NOi21      u039(.An(i_2_), .B(i_8_), .Y(men_men_n50_));
  NO3        u040(.A(men_men_n50_), .B(men_men_n47_), .C(men_men_n37_), .Y(men_men_n51_));
  NO3        u041(.A(men_men_n51_), .B(men_men_n49_), .C(men_men_n48_), .Y(men_men_n52_));
  INV        u042(.A(men_men_n52_), .Y(men_men_n53_));
  NOi31      u043(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n54_));
  NA2        u044(.A(men_men_n54_), .B(i_0_), .Y(men_men_n55_));
  NOi21      u045(.An(i_4_), .B(i_3_), .Y(men_men_n56_));
  NOi21      u046(.An(i_1_), .B(i_4_), .Y(men_men_n57_));
  OAI210     u047(.A0(men_men_n57_), .A1(men_men_n56_), .B0(men_men_n50_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n58_), .B(men_men_n55_), .Y(men_men_n59_));
  AN2        u049(.A(i_8_), .B(i_7_), .Y(men_men_n60_));
  NA2        u050(.A(men_men_n60_), .B(men_men_n12_), .Y(men_men_n61_));
  NOi21      u051(.An(i_8_), .B(i_7_), .Y(men_men_n62_));
  NA3        u052(.A(men_men_n62_), .B(men_men_n56_), .C(i_6_), .Y(men_men_n63_));
  OAI210     u053(.A0(men_men_n61_), .A1(men_men_n49_), .B0(men_men_n63_), .Y(men_men_n64_));
  AOI220     u054(.A0(men_men_n64_), .A1(men_men_n32_), .B0(men_men_n59_), .B1(men_men_n36_), .Y(men_men_n65_));
  NA4        u055(.A(men_men_n65_), .B(men_men_n53_), .C(men_men_n46_), .D(men_men_n27_), .Y(men_men_n66_));
  NA2        u056(.A(i_8_), .B(i_7_), .Y(men_men_n67_));
  NO3        u057(.A(men_men_n67_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n68_));
  NA2        u058(.A(i_8_), .B(men_men_n23_), .Y(men_men_n69_));
  AOI220     u059(.A0(men_men_n42_), .A1(i_1_), .B0(men_men_n38_), .B1(i_2_), .Y(men_men_n70_));
  NOi21      u060(.An(i_1_), .B(i_2_), .Y(men_men_n71_));
  NO2        u061(.A(men_men_n70_), .B(men_men_n69_), .Y(men_men_n72_));
  OAI210     u062(.A0(men_men_n72_), .A1(men_men_n68_), .B0(men_men_n14_), .Y(men_men_n73_));
  NA3        u063(.A(men_men_n62_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n74_));
  NA3        u064(.A(i_1_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n75_));
  NA2        u065(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  NOi32      u066(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n77_));
  NA2        u067(.A(men_men_n77_), .B(i_3_), .Y(men_men_n78_));
  NA3        u068(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n79_));
  NA2        u069(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NO2        u070(.A(i_0_), .B(i_4_), .Y(men_men_n81_));
  AOI220     u071(.A0(men_men_n81_), .A1(men_men_n80_), .B0(men_men_n76_), .B1(men_men_n56_), .Y(men_men_n82_));
  NA2        u072(.A(men_men_n82_), .B(men_men_n73_), .Y(men_men_n83_));
  NAi21      u073(.An(i_3_), .B(i_6_), .Y(men_men_n84_));
  NA2        u074(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n85_));
  NOi21      u075(.An(i_7_), .B(i_8_), .Y(men_men_n86_));
  NOi31      u076(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n87_));
  AOI210     u077(.A0(men_men_n86_), .A1(men_men_n12_), .B0(men_men_n87_), .Y(men_men_n88_));
  OAI210     u078(.A0(men_men_n88_), .A1(men_men_n11_), .B0(men_men_n85_), .Y(men_men_n89_));
  NA2        u079(.A(men_men_n89_), .B(men_men_n71_), .Y(men_men_n90_));
  NA3        u080(.A(men_men_n25_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n91_));
  NO2        u081(.A(men_men_n22_), .B(men_men_n91_), .Y(men_men_n92_));
  NA3        u082(.A(men_men_n21_), .B(i_5_), .C(i_7_), .Y(men_men_n93_));
  NA2        u083(.A(i_4_), .B(i_5_), .Y(men_men_n94_));
  NA3        u084(.A(men_men_n67_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n95_));
  OAI220     u085(.A0(men_men_n95_), .A1(men_men_n94_), .B0(men_men_n93_), .B1(i_0_), .Y(men_men_n96_));
  NO2        u086(.A(men_men_n96_), .B(men_men_n92_), .Y(men_men_n97_));
  NA3        u087(.A(men_men_n62_), .B(men_men_n32_), .C(i_3_), .Y(men_men_n98_));
  NA2        u088(.A(men_men_n41_), .B(i_6_), .Y(men_men_n99_));
  AOI210     u089(.A0(men_men_n99_), .A1(men_men_n22_), .B0(men_men_n98_), .Y(men_men_n100_));
  NOi21      u090(.An(i_2_), .B(i_1_), .Y(men_men_n101_));
  AN3        u091(.A(men_men_n86_), .B(men_men_n101_), .C(men_men_n47_), .Y(men_men_n102_));
  NAi21      u092(.An(i_6_), .B(i_0_), .Y(men_men_n103_));
  NA3        u093(.A(men_men_n57_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n104_));
  NOi21      u094(.An(i_4_), .B(i_6_), .Y(men_men_n105_));
  NOi21      u095(.An(i_5_), .B(i_3_), .Y(men_men_n106_));
  NA3        u096(.A(men_men_n106_), .B(men_men_n71_), .C(men_men_n105_), .Y(men_men_n107_));
  OAI210     u097(.A0(men_men_n104_), .A1(men_men_n103_), .B0(men_men_n107_), .Y(men_men_n108_));
  NA2        u098(.A(men_men_n71_), .B(men_men_n34_), .Y(men_men_n109_));
  NOi21      u099(.An(men_men_n39_), .B(men_men_n109_), .Y(men_men_n110_));
  NO4        u100(.A(men_men_n110_), .B(men_men_n108_), .C(men_men_n102_), .D(men_men_n100_), .Y(men_men_n111_));
  AOI220     u101(.A0(i_6_), .A1(i_7_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n112_));
  NOi31      u102(.An(men_men_n47_), .B(men_men_n112_), .C(i_2_), .Y(men_men_n113_));
  NA2        u103(.A(men_men_n62_), .B(men_men_n12_), .Y(men_men_n114_));
  NA2        u104(.A(men_men_n34_), .B(men_men_n14_), .Y(men_men_n115_));
  NOi21      u105(.An(i_3_), .B(i_1_), .Y(men_men_n116_));
  NA2        u106(.A(men_men_n116_), .B(i_4_), .Y(men_men_n117_));
  AOI210     u107(.A0(men_men_n115_), .A1(men_men_n114_), .B0(men_men_n117_), .Y(men_men_n118_));
  AOI220     u108(.A0(men_men_n86_), .A1(men_men_n14_), .B0(men_men_n105_), .B1(men_men_n23_), .Y(men_men_n119_));
  NOi31      u109(.An(men_men_n42_), .B(men_men_n119_), .C(men_men_n32_), .Y(men_men_n120_));
  NO3        u110(.A(men_men_n120_), .B(men_men_n118_), .C(men_men_n113_), .Y(men_men_n121_));
  NA4        u111(.A(men_men_n121_), .B(men_men_n111_), .C(men_men_n97_), .D(men_men_n90_), .Y(men_men_n122_));
  NA2        u112(.A(men_men_n50_), .B(men_men_n15_), .Y(men_men_n123_));
  NOi31      u113(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n124_));
  NOi31      u114(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n125_));
  OAI210     u115(.A0(men_men_n125_), .A1(men_men_n124_), .B0(i_7_), .Y(men_men_n126_));
  NA3        u116(.A(men_men_n34_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n127_));
  NA4        u117(.A(men_men_n127_), .B(men_men_n126_), .C(men_men_n123_), .D(men_men_n109_), .Y(men_men_n128_));
  NA2        u118(.A(men_men_n128_), .B(men_men_n37_), .Y(men_men_n129_));
  NA2        u119(.A(men_men_n56_), .B(men_men_n35_), .Y(men_men_n130_));
  AOI210     u120(.A0(men_men_n130_), .A1(men_men_n74_), .B0(men_men_n28_), .Y(men_men_n131_));
  NA4        u121(.A(men_men_n60_), .B(men_men_n101_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n132_));
  NAi31      u122(.An(men_men_n103_), .B(men_men_n86_), .C(men_men_n101_), .Y(men_men_n133_));
  NA3        u123(.A(men_men_n62_), .B(men_men_n54_), .C(i_6_), .Y(men_men_n134_));
  NA3        u124(.A(men_men_n134_), .B(men_men_n133_), .C(men_men_n132_), .Y(men_men_n135_));
  NOi21      u125(.An(i_0_), .B(i_2_), .Y(men_men_n136_));
  NA3        u126(.A(men_men_n136_), .B(men_men_n35_), .C(men_men_n105_), .Y(men_men_n137_));
  NA3        u127(.A(men_men_n47_), .B(men_men_n39_), .C(men_men_n18_), .Y(men_men_n138_));
  NOi32      u128(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n139_));
  NA2        u129(.A(men_men_n139_), .B(men_men_n124_), .Y(men_men_n140_));
  NA3        u130(.A(men_men_n136_), .B(men_men_n56_), .C(men_men_n34_), .Y(men_men_n141_));
  NA4        u131(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n138_), .D(men_men_n137_), .Y(men_men_n142_));
  NA4        u132(.A(men_men_n54_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n143_));
  NA4        u133(.A(men_men_n57_), .B(men_men_n36_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n144_));
  NA3        u134(.A(men_men_n57_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n145_));
  NA3        u135(.A(men_men_n145_), .B(men_men_n144_), .C(men_men_n143_), .Y(men_men_n146_));
  NO4        u136(.A(men_men_n146_), .B(men_men_n142_), .C(men_men_n135_), .D(men_men_n131_), .Y(men_men_n147_));
  NO2        u137(.A(men_men_n123_), .B(men_men_n99_), .Y(men_men_n148_));
  NO4        u138(.A(i_2_), .B(men_men_n21_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n149_));
  NA2        u139(.A(i_2_), .B(i_4_), .Y(men_men_n150_));
  AOI210     u140(.A0(men_men_n103_), .A1(men_men_n84_), .B0(men_men_n150_), .Y(men_men_n151_));
  NO2        u141(.A(i_8_), .B(i_7_), .Y(men_men_n152_));
  OA210      u142(.A0(men_men_n151_), .A1(men_men_n149_), .B0(men_men_n152_), .Y(men_men_n153_));
  NA4        u143(.A(men_men_n116_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n154_));
  NO2        u144(.A(men_men_n154_), .B(i_4_), .Y(men_men_n155_));
  NO3        u145(.A(men_men_n155_), .B(men_men_n153_), .C(men_men_n148_), .Y(men_men_n156_));
  NA2        u146(.A(men_men_n86_), .B(men_men_n12_), .Y(men_men_n157_));
  NA3        u147(.A(i_2_), .B(i_1_), .C(men_men_n14_), .Y(men_men_n158_));
  NA2        u148(.A(men_men_n47_), .B(i_3_), .Y(men_men_n159_));
  AOI210     u149(.A0(men_men_n159_), .A1(men_men_n158_), .B0(men_men_n157_), .Y(men_men_n160_));
  NA3        u150(.A(men_men_n136_), .B(men_men_n62_), .C(men_men_n105_), .Y(men_men_n161_));
  OAI210     u151(.A0(men_men_n98_), .A1(men_men_n28_), .B0(men_men_n161_), .Y(men_men_n162_));
  NA3        u152(.A(men_men_n50_), .B(men_men_n33_), .C(men_men_n15_), .Y(men_men_n163_));
  NOi31      u153(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n164_));
  OAI210     u154(.A0(men_men_n139_), .A1(men_men_n77_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u155(.A(men_men_n165_), .B(men_men_n163_), .Y(men_men_n166_));
  NO3        u156(.A(men_men_n166_), .B(men_men_n162_), .C(men_men_n160_), .Y(men_men_n167_));
  NA4        u157(.A(men_men_n167_), .B(men_men_n156_), .C(men_men_n147_), .D(men_men_n129_), .Y(men_men_n168_));
  OR4        u158(.A(men_men_n168_), .B(men_men_n122_), .C(men_men_n83_), .D(men_men_n66_), .Y(men00));
  INV        u159(.A(i_1_), .Y(men_men_n172_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule