//Benchmark atmr_max1024_476_0.25

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x8), .B(x3), .Y(ori_ori_n26_));
  NA2        o010(.A(x4), .B(x2), .Y(ori_ori_n27_));
  NO3        o011(.A(ori_ori_n27_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n28_));
  NO2        o012(.A(ori_ori_n28_), .B(ori_ori_n24_), .Y(ori_ori_n29_));
  NO2        o013(.A(x4), .B(x3), .Y(ori_ori_n30_));
  INV        o014(.A(ori_ori_n30_), .Y(ori_ori_n31_));
  NOi21      o015(.An(ori_ori_n23_), .B(ori_ori_n29_), .Y(ori00));
  NO2        o016(.A(x1), .B(x0), .Y(ori_ori_n33_));
  INV        o017(.A(x6), .Y(ori_ori_n34_));
  NO2        o018(.A(ori_ori_n34_), .B(ori_ori_n25_), .Y(ori_ori_n35_));
  AN2        o019(.A(x8), .B(x7), .Y(ori_ori_n36_));
  NA2        o020(.A(ori_ori_n35_), .B(ori_ori_n33_), .Y(ori_ori_n37_));
  NA2        o021(.A(x4), .B(x3), .Y(ori_ori_n38_));
  AOI210     o022(.A0(ori_ori_n37_), .A1(ori_ori_n23_), .B0(ori_ori_n38_), .Y(ori_ori_n39_));
  NO2        o023(.A(x2), .B(x0), .Y(ori_ori_n40_));
  INV        o024(.A(x3), .Y(ori_ori_n41_));
  NO2        o025(.A(ori_ori_n41_), .B(ori_ori_n18_), .Y(ori_ori_n42_));
  INV        o026(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n35_), .B(x4), .Y(ori_ori_n44_));
  OAI210     o028(.A0(ori_ori_n44_), .A1(ori_ori_n43_), .B0(ori_ori_n40_), .Y(ori_ori_n45_));
  INV        o029(.A(x4), .Y(ori_ori_n46_));
  NO2        o030(.A(ori_ori_n46_), .B(ori_ori_n17_), .Y(ori_ori_n47_));
  NA2        o031(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n48_));
  OAI210     o032(.A0(ori_ori_n48_), .A1(ori_ori_n20_), .B0(ori_ori_n45_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n50_));
  AOI220     o034(.A0(ori_ori_n50_), .A1(ori_ori_n33_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n51_));
  INV        o035(.A(x2), .Y(ori_ori_n52_));
  NO2        o036(.A(ori_ori_n52_), .B(ori_ori_n17_), .Y(ori_ori_n53_));
  NA2        o037(.A(ori_ori_n41_), .B(ori_ori_n18_), .Y(ori_ori_n54_));
  NA2        o038(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  OAI210     o039(.A0(ori_ori_n51_), .A1(ori_ori_n31_), .B0(ori_ori_n55_), .Y(ori_ori_n56_));
  NO3        o040(.A(ori_ori_n56_), .B(ori_ori_n49_), .C(ori_ori_n39_), .Y(ori01));
  NA2        o041(.A(ori_ori_n41_), .B(x1), .Y(ori_ori_n58_));
  INV        o042(.A(x9), .Y(ori_ori_n59_));
  NO2        o043(.A(ori_ori_n58_), .B(x5), .Y(ori_ori_n60_));
  OAI210     o044(.A0(ori_ori_n42_), .A1(ori_ori_n25_), .B0(ori_ori_n52_), .Y(ori_ori_n61_));
  OAI210     o045(.A0(ori_ori_n54_), .A1(ori_ori_n20_), .B0(ori_ori_n61_), .Y(ori_ori_n62_));
  INV        o046(.A(ori_ori_n62_), .Y(ori_ori_n63_));
  NA2        o047(.A(ori_ori_n63_), .B(x4), .Y(ori_ori_n64_));
  NA2        o048(.A(ori_ori_n46_), .B(x2), .Y(ori_ori_n65_));
  OAI210     o049(.A0(ori_ori_n65_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n66_));
  NA2        o050(.A(x5), .B(x3), .Y(ori_ori_n67_));
  NO2        o051(.A(x8), .B(x6), .Y(ori_ori_n68_));
  NAi21      o052(.An(x4), .B(x3), .Y(ori_ori_n69_));
  INV        o053(.A(ori_ori_n69_), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n70_), .B(ori_ori_n22_), .Y(ori_ori_n71_));
  NO2        o055(.A(x4), .B(x2), .Y(ori_ori_n72_));
  NO2        o056(.A(ori_ori_n71_), .B(ori_ori_n18_), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n73_), .B(ori_ori_n66_), .Y(ori_ori_n74_));
  NA2        o058(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n75_));
  NO2        o059(.A(ori_ori_n75_), .B(ori_ori_n25_), .Y(ori_ori_n76_));
  INV        o060(.A(x8), .Y(ori_ori_n77_));
  NA2        o061(.A(x2), .B(x1), .Y(ori_ori_n78_));
  AOI210     o062(.A0(ori_ori_n54_), .A1(ori_ori_n25_), .B0(ori_ori_n52_), .Y(ori_ori_n79_));
  OAI210     o063(.A0(ori_ori_n43_), .A1(ori_ori_n35_), .B0(ori_ori_n46_), .Y(ori_ori_n80_));
  NO2        o064(.A(ori_ori_n80_), .B(ori_ori_n79_), .Y(ori_ori_n81_));
  NA2        o065(.A(x4), .B(ori_ori_n41_), .Y(ori_ori_n82_));
  NO2        o066(.A(ori_ori_n46_), .B(ori_ori_n52_), .Y(ori_ori_n83_));
  AOI210     o067(.A0(ori_ori_n82_), .A1(ori_ori_n50_), .B0(x1), .Y(ori_ori_n84_));
  NA2        o068(.A(ori_ori_n52_), .B(x1), .Y(ori_ori_n85_));
  OAI210     o069(.A0(ori_ori_n85_), .A1(ori_ori_n38_), .B0(ori_ori_n17_), .Y(ori_ori_n86_));
  NO3        o070(.A(ori_ori_n86_), .B(ori_ori_n84_), .C(ori_ori_n81_), .Y(ori_ori_n87_));
  AO210      o071(.A0(ori_ori_n74_), .A1(ori_ori_n64_), .B0(ori_ori_n87_), .Y(ori02));
  NO2        o072(.A(x3), .B(ori_ori_n52_), .Y(ori_ori_n89_));
  NO2        o073(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n90_));
  NA2        o074(.A(ori_ori_n41_), .B(x0), .Y(ori_ori_n91_));
  OR2        o075(.A(x8), .B(x0), .Y(ori_ori_n92_));
  INV        o076(.A(ori_ori_n92_), .Y(ori_ori_n93_));
  NAi21      o077(.An(x2), .B(x8), .Y(ori_ori_n94_));
  INV        o078(.A(ori_ori_n94_), .Y(ori_ori_n95_));
  NO2        o079(.A(x4), .B(x1), .Y(ori_ori_n96_));
  NA2        o080(.A(ori_ori_n96_), .B(x2), .Y(ori_ori_n97_));
  NOi21      o081(.An(x0), .B(x4), .Y(ori_ori_n98_));
  NO2        o082(.A(ori_ori_n97_), .B(ori_ori_n67_), .Y(ori_ori_n99_));
  NO2        o083(.A(x5), .B(ori_ori_n46_), .Y(ori_ori_n100_));
  NA2        o084(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n101_));
  AOI210     o085(.A0(ori_ori_n101_), .A1(ori_ori_n85_), .B0(ori_ori_n91_), .Y(ori_ori_n102_));
  OAI210     o086(.A0(ori_ori_n102_), .A1(ori_ori_n33_), .B0(ori_ori_n100_), .Y(ori_ori_n103_));
  NO2        o087(.A(x7), .B(x0), .Y(ori_ori_n104_));
  NO2        o088(.A(ori_ori_n72_), .B(ori_ori_n83_), .Y(ori_ori_n105_));
  NO2        o089(.A(ori_ori_n21_), .B(ori_ori_n41_), .Y(ori_ori_n106_));
  NA2        o090(.A(x5), .B(x0), .Y(ori_ori_n107_));
  NO2        o091(.A(ori_ori_n46_), .B(x2), .Y(ori_ori_n108_));
  NA2        o092(.A(ori_ori_n108_), .B(ori_ori_n106_), .Y(ori_ori_n109_));
  NA3        o093(.A(ori_ori_n109_), .B(ori_ori_n103_), .C(ori_ori_n34_), .Y(ori_ori_n110_));
  NO2        o094(.A(ori_ori_n110_), .B(ori_ori_n99_), .Y(ori_ori_n111_));
  NO3        o095(.A(ori_ori_n67_), .B(ori_ori_n65_), .C(ori_ori_n24_), .Y(ori_ori_n112_));
  NO2        o096(.A(ori_ori_n27_), .B(ori_ori_n25_), .Y(ori_ori_n113_));
  NA2        o097(.A(x7), .B(x3), .Y(ori_ori_n114_));
  NO2        o098(.A(ori_ori_n82_), .B(x5), .Y(ori_ori_n115_));
  NOi21      o099(.An(x8), .B(x0), .Y(ori_ori_n116_));
  NO2        o100(.A(ori_ori_n41_), .B(x2), .Y(ori_ori_n117_));
  INV        o101(.A(x7), .Y(ori_ori_n118_));
  NA2        o102(.A(ori_ori_n118_), .B(ori_ori_n18_), .Y(ori_ori_n119_));
  AOI220     o103(.A0(ori_ori_n119_), .A1(ori_ori_n117_), .B0(ori_ori_n89_), .B1(ori_ori_n36_), .Y(ori_ori_n120_));
  NO2        o104(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n121_));
  NO2        o105(.A(ori_ori_n121_), .B(ori_ori_n98_), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n122_), .B(ori_ori_n120_), .Y(ori_ori_n123_));
  AOI210     o107(.A0(ori_ori_n116_), .A1(ori_ori_n115_), .B0(ori_ori_n123_), .Y(ori_ori_n124_));
  OAI210     o108(.A0(ori_ori_n114_), .A1(ori_ori_n48_), .B0(ori_ori_n124_), .Y(ori_ori_n125_));
  NA2        o109(.A(x5), .B(x1), .Y(ori_ori_n126_));
  INV        o110(.A(ori_ori_n126_), .Y(ori_ori_n127_));
  AOI210     o111(.A0(ori_ori_n127_), .A1(ori_ori_n98_), .B0(ori_ori_n34_), .Y(ori_ori_n128_));
  NO2        o112(.A(ori_ori_n59_), .B(ori_ori_n77_), .Y(ori_ori_n129_));
  NAi21      o113(.An(x2), .B(x7), .Y(ori_ori_n130_));
  NO2        o114(.A(ori_ori_n130_), .B(ori_ori_n46_), .Y(ori_ori_n131_));
  NA2        o115(.A(ori_ori_n131_), .B(ori_ori_n60_), .Y(ori_ori_n132_));
  NAi31      o116(.An(ori_ori_n67_), .B(ori_ori_n36_), .C(ori_ori_n33_), .Y(ori_ori_n133_));
  NA3        o117(.A(ori_ori_n133_), .B(ori_ori_n132_), .C(ori_ori_n128_), .Y(ori_ori_n134_));
  NO3        o118(.A(ori_ori_n134_), .B(ori_ori_n125_), .C(ori_ori_n112_), .Y(ori_ori_n135_));
  NO2        o119(.A(ori_ori_n135_), .B(ori_ori_n111_), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n107_), .B(ori_ori_n105_), .Y(ori_ori_n137_));
  NA2        o121(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n138_));
  NA2        o122(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n139_));
  NA3        o123(.A(ori_ori_n139_), .B(ori_ori_n138_), .C(ori_ori_n24_), .Y(ori_ori_n140_));
  AN2        o124(.A(ori_ori_n140_), .B(ori_ori_n108_), .Y(ori_ori_n141_));
  NA2        o125(.A(x8), .B(x0), .Y(ori_ori_n142_));
  NO2        o126(.A(ori_ori_n118_), .B(ori_ori_n25_), .Y(ori_ori_n143_));
  NA2        o127(.A(x2), .B(x0), .Y(ori_ori_n144_));
  NA2        o128(.A(x4), .B(x1), .Y(ori_ori_n145_));
  NAi21      o129(.An(ori_ori_n96_), .B(ori_ori_n145_), .Y(ori_ori_n146_));
  NOi21      o130(.An(ori_ori_n146_), .B(ori_ori_n144_), .Y(ori_ori_n147_));
  NO3        o131(.A(ori_ori_n147_), .B(ori_ori_n141_), .C(ori_ori_n137_), .Y(ori_ori_n148_));
  NO2        o132(.A(ori_ori_n148_), .B(ori_ori_n41_), .Y(ori_ori_n149_));
  NO2        o133(.A(ori_ori_n140_), .B(ori_ori_n65_), .Y(ori_ori_n150_));
  INV        o134(.A(ori_ori_n100_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n85_), .B(ori_ori_n17_), .Y(ori_ori_n152_));
  NO2        o136(.A(ori_ori_n33_), .B(ori_ori_n152_), .Y(ori_ori_n153_));
  NO3        o137(.A(ori_ori_n153_), .B(ori_ori_n151_), .C(x7), .Y(ori_ori_n154_));
  NA3        o138(.A(ori_ori_n146_), .B(ori_ori_n151_), .C(ori_ori_n40_), .Y(ori_ori_n155_));
  OAI210     o139(.A0(ori_ori_n139_), .A1(ori_ori_n105_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NO3        o140(.A(ori_ori_n156_), .B(ori_ori_n154_), .C(ori_ori_n150_), .Y(ori_ori_n157_));
  NO2        o141(.A(ori_ori_n157_), .B(x3), .Y(ori_ori_n158_));
  NO3        o142(.A(ori_ori_n158_), .B(ori_ori_n149_), .C(ori_ori_n136_), .Y(ori03));
  NO2        o143(.A(ori_ori_n46_), .B(x3), .Y(ori_ori_n160_));
  NO2        o144(.A(ori_ori_n52_), .B(x1), .Y(ori_ori_n161_));
  NO2        o145(.A(ori_ori_n67_), .B(x6), .Y(ori_ori_n162_));
  NA2        o146(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n163_));
  NO2        o147(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n164_));
  AN2        o148(.A(ori_ori_n162_), .B(ori_ori_n53_), .Y(ori_ori_n165_));
  INV        o149(.A(ori_ori_n165_), .Y(ori_ori_n166_));
  NA2        o150(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n167_));
  NO2        o151(.A(ori_ori_n167_), .B(ori_ori_n163_), .Y(ori_ori_n168_));
  INV        o152(.A(ori_ori_n163_), .Y(ori_ori_n169_));
  NO2        o153(.A(x3), .B(ori_ori_n144_), .Y(ori_ori_n170_));
  AOI210     o154(.A0(ori_ori_n170_), .A1(ori_ori_n169_), .B0(ori_ori_n168_), .Y(ori_ori_n171_));
  NO3        o155(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n172_));
  NO2        o156(.A(x5), .B(x1), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n167_), .B(ori_ori_n138_), .Y(ori_ori_n174_));
  NO3        o158(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n175_));
  NO2        o159(.A(ori_ori_n175_), .B(ori_ori_n174_), .Y(ori_ori_n176_));
  INV        o160(.A(ori_ori_n176_), .Y(ori_ori_n177_));
  AOI220     o161(.A0(ori_ori_n177_), .A1(ori_ori_n46_), .B0(ori_ori_n172_), .B1(ori_ori_n100_), .Y(ori_ori_n178_));
  NA3        o162(.A(ori_ori_n178_), .B(ori_ori_n171_), .C(ori_ori_n166_), .Y(ori_ori_n179_));
  NO2        o163(.A(ori_ori_n46_), .B(ori_ori_n41_), .Y(ori_ori_n180_));
  NA2        o164(.A(ori_ori_n180_), .B(ori_ori_n19_), .Y(ori_ori_n181_));
  NO2        o165(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n182_));
  NO2        o166(.A(ori_ori_n182_), .B(x6), .Y(ori_ori_n183_));
  NA2        o167(.A(ori_ori_n41_), .B(ori_ori_n52_), .Y(ori_ori_n184_));
  NA2        o168(.A(ori_ori_n108_), .B(ori_ori_n76_), .Y(ori_ori_n185_));
  NA2        o169(.A(x6), .B(ori_ori_n46_), .Y(ori_ori_n186_));
  OAI210     o170(.A0(ori_ori_n93_), .A1(ori_ori_n68_), .B0(x4), .Y(ori_ori_n187_));
  AOI210     o171(.A0(ori_ori_n187_), .A1(ori_ori_n186_), .B0(ori_ori_n67_), .Y(ori_ori_n188_));
  NA2        o172(.A(ori_ori_n100_), .B(x6), .Y(ori_ori_n189_));
  INV        o173(.A(ori_ori_n60_), .Y(ori_ori_n190_));
  NA2        o174(.A(ori_ori_n190_), .B(ori_ori_n189_), .Y(ori_ori_n191_));
  OAI210     o175(.A0(ori_ori_n191_), .A1(ori_ori_n188_), .B0(x2), .Y(ori_ori_n192_));
  NA3        o176(.A(ori_ori_n192_), .B(ori_ori_n185_), .C(x7), .Y(ori_ori_n193_));
  AOI210     o177(.A0(ori_ori_n179_), .A1(x8), .B0(ori_ori_n193_), .Y(ori_ori_n194_));
  NO2        o178(.A(ori_ori_n75_), .B(ori_ori_n25_), .Y(ori_ori_n195_));
  AOI210     o179(.A0(ori_ori_n183_), .A1(ori_ori_n121_), .B0(ori_ori_n195_), .Y(ori_ori_n196_));
  NO2        o180(.A(ori_ori_n196_), .B(x2), .Y(ori_ori_n197_));
  NA2        o181(.A(x2), .B(ori_ori_n60_), .Y(ori_ori_n198_));
  NA2        o182(.A(ori_ori_n41_), .B(ori_ori_n17_), .Y(ori_ori_n199_));
  INV        o183(.A(x6), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n167_), .B(x6), .Y(ori_ori_n201_));
  NAi21      o185(.An(ori_ori_n129_), .B(ori_ori_n201_), .Y(ori_ori_n202_));
  NA3        o186(.A(ori_ori_n202_), .B(ori_ori_n200_), .C(ori_ori_n113_), .Y(ori_ori_n203_));
  NA3        o187(.A(ori_ori_n203_), .B(ori_ori_n198_), .C(ori_ori_n118_), .Y(ori_ori_n204_));
  NA2        o188(.A(x6), .B(x2), .Y(ori_ori_n205_));
  OR2        o189(.A(ori_ori_n162_), .B(ori_ori_n115_), .Y(ori_ori_n206_));
  NA2        o190(.A(x4), .B(x0), .Y(ori_ori_n207_));
  NA2        o191(.A(ori_ori_n206_), .B(ori_ori_n40_), .Y(ori_ori_n208_));
  NO2        o192(.A(ori_ori_n208_), .B(x8), .Y(ori_ori_n209_));
  NA2        o193(.A(ori_ori_n173_), .B(x6), .Y(ori_ori_n210_));
  INV        o194(.A(ori_ori_n142_), .Y(ori_ori_n211_));
  NO2        o195(.A(ori_ori_n210_), .B(ori_ori_n184_), .Y(ori_ori_n212_));
  NO4        o196(.A(ori_ori_n212_), .B(ori_ori_n209_), .C(ori_ori_n204_), .D(ori_ori_n197_), .Y(ori_ori_n213_));
  NA2        o197(.A(ori_ori_n201_), .B(x2), .Y(ori_ori_n214_));
  OAI210     o198(.A0(ori_ori_n211_), .A1(x6), .B0(ori_ori_n42_), .Y(ori_ori_n215_));
  AOI210     o199(.A0(ori_ori_n215_), .A1(ori_ori_n214_), .B0(ori_ori_n151_), .Y(ori_ori_n216_));
  NOi21      o200(.An(ori_ori_n205_), .B(ori_ori_n17_), .Y(ori_ori_n217_));
  NA3        o201(.A(ori_ori_n217_), .B(ori_ori_n173_), .C(ori_ori_n38_), .Y(ori_ori_n218_));
  AOI210     o202(.A0(ori_ori_n34_), .A1(ori_ori_n52_), .B0(x0), .Y(ori_ori_n219_));
  NA3        o203(.A(ori_ori_n219_), .B(ori_ori_n127_), .C(ori_ori_n31_), .Y(ori_ori_n220_));
  NA2        o204(.A(x3), .B(x2), .Y(ori_ori_n221_));
  AOI220     o205(.A0(ori_ori_n221_), .A1(ori_ori_n184_), .B0(ori_ori_n220_), .B1(ori_ori_n218_), .Y(ori_ori_n222_));
  NAi21      o206(.An(x4), .B(x0), .Y(ori_ori_n223_));
  NO3        o207(.A(ori_ori_n223_), .B(ori_ori_n42_), .C(x2), .Y(ori_ori_n224_));
  OAI210     o208(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n224_), .Y(ori_ori_n225_));
  NO2        o209(.A(ori_ori_n219_), .B(ori_ori_n217_), .Y(ori_ori_n226_));
  AOI220     o210(.A0(ori_ori_n226_), .A1(ori_ori_n70_), .B0(ori_ori_n18_), .B1(ori_ori_n30_), .Y(ori_ori_n227_));
  AOI210     o211(.A0(ori_ori_n227_), .A1(ori_ori_n225_), .B0(ori_ori_n25_), .Y(ori_ori_n228_));
  NA3        o212(.A(ori_ori_n34_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n229_));
  NO2        o213(.A(ori_ori_n219_), .B(ori_ori_n217_), .Y(ori_ori_n230_));
  INV        o214(.A(ori_ori_n174_), .Y(ori_ori_n231_));
  NA2        o215(.A(ori_ori_n34_), .B(ori_ori_n41_), .Y(ori_ori_n232_));
  OR2        o216(.A(ori_ori_n232_), .B(ori_ori_n207_), .Y(ori_ori_n233_));
  OAI220     o217(.A0(ori_ori_n233_), .A1(ori_ori_n126_), .B0(ori_ori_n186_), .B1(ori_ori_n231_), .Y(ori_ori_n234_));
  AO210      o218(.A0(ori_ori_n230_), .A1(ori_ori_n115_), .B0(ori_ori_n234_), .Y(ori_ori_n235_));
  NO4        o219(.A(ori_ori_n235_), .B(ori_ori_n228_), .C(ori_ori_n222_), .D(ori_ori_n216_), .Y(ori_ori_n236_));
  OAI210     o220(.A0(ori_ori_n213_), .A1(ori_ori_n194_), .B0(ori_ori_n236_), .Y(ori04));
  NO2        o221(.A(x2), .B(x1), .Y(ori_ori_n238_));
  OAI210     o222(.A0(ori_ori_n199_), .A1(ori_ori_n238_), .B0(ori_ori_n34_), .Y(ori_ori_n239_));
  NO2        o223(.A(ori_ori_n221_), .B(ori_ori_n164_), .Y(ori_ori_n240_));
  NA2        o224(.A(ori_ori_n240_), .B(ori_ori_n77_), .Y(ori_ori_n241_));
  NA2        o225(.A(ori_ori_n241_), .B(x6), .Y(ori_ori_n242_));
  NA2        o226(.A(ori_ori_n242_), .B(ori_ori_n239_), .Y(ori_ori_n243_));
  NO2        o227(.A(x2), .B(ori_ori_n91_), .Y(ori_ori_n244_));
  NO3        o228(.A(ori_ori_n341_), .B(ori_ori_n94_), .C(ori_ori_n18_), .Y(ori_ori_n245_));
  NO2        o229(.A(ori_ori_n245_), .B(ori_ori_n244_), .Y(ori_ori_n246_));
  OAI210     o230(.A0(ori_ori_n92_), .A1(ori_ori_n85_), .B0(ori_ori_n142_), .Y(ori_ori_n247_));
  NA3        o231(.A(ori_ori_n247_), .B(x6), .C(x3), .Y(ori_ori_n248_));
  NOi21      o232(.An(ori_ori_n116_), .B(ori_ori_n101_), .Y(ori_ori_n249_));
  NO2        o233(.A(ori_ori_n344_), .B(ori_ori_n229_), .Y(ori_ori_n250_));
  AOI210     o234(.A0(ori_ori_n249_), .A1(x6), .B0(ori_ori_n250_), .Y(ori_ori_n251_));
  NA2        o235(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n252_));
  OAI210     o236(.A0(ori_ori_n85_), .A1(ori_ori_n17_), .B0(ori_ori_n252_), .Y(ori_ori_n253_));
  NA2        o237(.A(ori_ori_n253_), .B(ori_ori_n68_), .Y(ori_ori_n254_));
  NA4        o238(.A(ori_ori_n254_), .B(ori_ori_n251_), .C(ori_ori_n248_), .D(ori_ori_n246_), .Y(ori_ori_n255_));
  NA2        o239(.A(ori_ori_n172_), .B(ori_ori_n72_), .Y(ori_ori_n256_));
  NA2        o240(.A(ori_ori_n256_), .B(ori_ori_n118_), .Y(ori_ori_n257_));
  AOI210     o241(.A0(ori_ori_n255_), .A1(x4), .B0(ori_ori_n257_), .Y(ori_ori_n258_));
  XO2        o242(.A(x4), .B(x0), .Y(ori_ori_n259_));
  NA2        o243(.A(x4), .B(ori_ori_n78_), .Y(ori_ori_n260_));
  NO2        o244(.A(ori_ori_n260_), .B(x3), .Y(ori_ori_n261_));
  INV        o245(.A(ori_ori_n78_), .Y(ori_ori_n262_));
  NO2        o246(.A(ori_ori_n77_), .B(x4), .Y(ori_ori_n263_));
  AOI220     o247(.A0(ori_ori_n263_), .A1(ori_ori_n42_), .B0(ori_ori_n98_), .B1(ori_ori_n262_), .Y(ori_ori_n264_));
  NA3        o248(.A(ori_ori_n264_), .B(ori_ori_n181_), .C(x6), .Y(ori_ori_n265_));
  OAI220     o249(.A0(ori_ori_n223_), .A1(ori_ori_n75_), .B0(ori_ori_n144_), .B1(ori_ori_n77_), .Y(ori_ori_n266_));
  NA2        o250(.A(ori_ori_n266_), .B(ori_ori_n58_), .Y(ori_ori_n267_));
  NO2        o251(.A(ori_ori_n116_), .B(ori_ori_n69_), .Y(ori_ori_n268_));
  NO2        o252(.A(ori_ori_n33_), .B(x2), .Y(ori_ori_n269_));
  NOi21      o253(.An(ori_ori_n96_), .B(ori_ori_n26_), .Y(ori_ori_n270_));
  AOI210     o254(.A0(ori_ori_n269_), .A1(ori_ori_n268_), .B0(ori_ori_n270_), .Y(ori_ori_n271_));
  OAI210     o255(.A0(ori_ori_n267_), .A1(ori_ori_n59_), .B0(ori_ori_n271_), .Y(ori_ori_n272_));
  OAI220     o256(.A0(ori_ori_n272_), .A1(x6), .B0(ori_ori_n265_), .B1(ori_ori_n261_), .Y(ori_ori_n273_));
  OAI210     o257(.A0(x6), .A1(ori_ori_n46_), .B0(ori_ori_n40_), .Y(ori_ori_n274_));
  OAI210     o258(.A0(ori_ori_n274_), .A1(ori_ori_n77_), .B0(ori_ori_n233_), .Y(ori_ori_n275_));
  AOI210     o259(.A0(ori_ori_n275_), .A1(ori_ori_n18_), .B0(ori_ori_n118_), .Y(ori_ori_n276_));
  AO220      o260(.A0(ori_ori_n276_), .A1(ori_ori_n273_), .B0(ori_ori_n258_), .B1(ori_ori_n243_), .Y(ori_ori_n277_));
  NA2        o261(.A(ori_ori_n269_), .B(x6), .Y(ori_ori_n278_));
  AOI210     o262(.A0(x6), .A1(x1), .B0(ori_ori_n117_), .Y(ori_ori_n279_));
  NA2        o263(.A(ori_ori_n263_), .B(x0), .Y(ori_ori_n280_));
  NA2        o264(.A(ori_ori_n72_), .B(x6), .Y(ori_ori_n281_));
  OAI210     o265(.A0(ori_ori_n280_), .A1(ori_ori_n279_), .B0(ori_ori_n281_), .Y(ori_ori_n282_));
  NA2        o266(.A(ori_ori_n282_), .B(ori_ori_n278_), .Y(ori_ori_n283_));
  NA2        o267(.A(ori_ori_n283_), .B(ori_ori_n277_), .Y(ori_ori_n284_));
  AOI210     o268(.A0(ori_ori_n161_), .A1(x8), .B0(ori_ori_n90_), .Y(ori_ori_n285_));
  NA2        o269(.A(ori_ori_n285_), .B(ori_ori_n252_), .Y(ori_ori_n286_));
  NA3        o270(.A(ori_ori_n286_), .B(ori_ori_n160_), .C(ori_ori_n118_), .Y(ori_ori_n287_));
  OAI210     o271(.A0(ori_ori_n27_), .A1(x1), .B0(ori_ori_n184_), .Y(ori_ori_n288_));
  NA3        o272(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n289_));
  NA2        o273(.A(ori_ori_n180_), .B(x0), .Y(ori_ori_n290_));
  OAI220     o274(.A0(ori_ori_n290_), .A1(x2), .B0(ori_ori_n289_), .B1(ori_ori_n262_), .Y(ori_ori_n291_));
  AOI210     o275(.A0(ori_ori_n288_), .A1(ori_ori_n93_), .B0(ori_ori_n291_), .Y(ori_ori_n292_));
  AOI210     o276(.A0(ori_ori_n292_), .A1(ori_ori_n287_), .B0(ori_ori_n25_), .Y(ori_ori_n293_));
  NA3        o277(.A(ori_ori_n95_), .B(ori_ori_n180_), .C(x0), .Y(ori_ori_n294_));
  NAi31      o278(.An(ori_ori_n48_), .B(ori_ori_n342_), .C(ori_ori_n143_), .Y(ori_ori_n295_));
  NA2        o279(.A(ori_ori_n295_), .B(ori_ori_n294_), .Y(ori_ori_n296_));
  OAI210     o280(.A0(ori_ori_n296_), .A1(ori_ori_n293_), .B0(x6), .Y(ori_ori_n297_));
  OAI210     o281(.A0(ori_ori_n129_), .A1(ori_ori_n46_), .B0(ori_ori_n104_), .Y(ori_ori_n298_));
  NA2        o282(.A(ori_ori_n53_), .B(ori_ori_n36_), .Y(ori_ori_n299_));
  AOI220     o283(.A0(ori_ori_n299_), .A1(ori_ori_n298_), .B0(ori_ori_n38_), .B1(ori_ori_n31_), .Y(ori_ori_n300_));
  NA2        o284(.A(x7), .B(ori_ori_n180_), .Y(ori_ori_n301_));
  INV        o285(.A(x1), .Y(ori_ori_n302_));
  OAI210     o286(.A0(ori_ori_n301_), .A1(x8), .B0(ori_ori_n302_), .Y(ori_ori_n303_));
  NAi31      o287(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n304_));
  OAI210     o288(.A0(ori_ori_n304_), .A1(x4), .B0(ori_ori_n130_), .Y(ori_ori_n305_));
  NA2        o289(.A(ori_ori_n305_), .B(ori_ori_n114_), .Y(ori_ori_n306_));
  NO2        o290(.A(ori_ori_n118_), .B(x0), .Y(ori_ori_n307_));
  AOI220     o291(.A0(ori_ori_n307_), .A1(ori_ori_n343_), .B0(ori_ori_n268_), .B1(ori_ori_n118_), .Y(ori_ori_n308_));
  NA4        o292(.A(ori_ori_n308_), .B(x1), .C(ori_ori_n306_), .D(ori_ori_n48_), .Y(ori_ori_n309_));
  OAI210     o293(.A0(ori_ori_n303_), .A1(ori_ori_n300_), .B0(ori_ori_n309_), .Y(ori_ori_n310_));
  OAI210     o294(.A0(ori_ori_n223_), .A1(ori_ori_n41_), .B0(ori_ori_n259_), .Y(ori_ori_n311_));
  INV        o295(.A(ori_ori_n289_), .Y(ori_ori_n312_));
  AOI220     o296(.A0(ori_ori_n312_), .A1(ori_ori_n77_), .B0(ori_ori_n311_), .B1(ori_ori_n118_), .Y(ori_ori_n313_));
  NO2        o297(.A(ori_ori_n313_), .B(ori_ori_n52_), .Y(ori_ori_n314_));
  INV        o298(.A(ori_ori_n314_), .Y(ori_ori_n315_));
  AOI210     o299(.A0(ori_ori_n315_), .A1(ori_ori_n310_), .B0(ori_ori_n25_), .Y(ori_ori_n316_));
  NA4        o300(.A(ori_ori_n30_), .B(ori_ori_n77_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n317_));
  NO3        o301(.A(ori_ori_n344_), .B(ori_ori_n142_), .C(ori_ori_n38_), .Y(ori_ori_n318_));
  NA2        o302(.A(ori_ori_n318_), .B(x7), .Y(ori_ori_n319_));
  NA2        o303(.A(ori_ori_n319_), .B(ori_ori_n317_), .Y(ori_ori_n320_));
  OAI210     o304(.A0(ori_ori_n320_), .A1(ori_ori_n316_), .B0(ori_ori_n34_), .Y(ori_ori_n321_));
  INV        o305(.A(ori_ori_n307_), .Y(ori_ori_n322_));
  NO4        o306(.A(ori_ori_n322_), .B(ori_ori_n67_), .C(x4), .D(ori_ori_n52_), .Y(ori_ori_n323_));
  NA2        o307(.A(ori_ori_n199_), .B(ori_ori_n21_), .Y(ori_ori_n324_));
  NO2        o308(.A(ori_ori_n126_), .B(ori_ori_n104_), .Y(ori_ori_n325_));
  NA2        o309(.A(ori_ori_n325_), .B(ori_ori_n324_), .Y(ori_ori_n326_));
  AOI210     o310(.A0(ori_ori_n326_), .A1(ori_ori_n133_), .B0(ori_ori_n27_), .Y(ori_ori_n327_));
  NA2        o311(.A(ori_ori_n116_), .B(ori_ori_n161_), .Y(ori_ori_n328_));
  NA2        o312(.A(ori_ori_n328_), .B(ori_ori_n304_), .Y(ori_ori_n329_));
  NA2        o313(.A(ori_ori_n329_), .B(ori_ori_n143_), .Y(ori_ori_n330_));
  NO2        o314(.A(ori_ori_n126_), .B(ori_ori_n41_), .Y(ori_ori_n331_));
  NA2        o315(.A(x3), .B(ori_ori_n52_), .Y(ori_ori_n332_));
  NO2        o316(.A(ori_ori_n119_), .B(ori_ori_n332_), .Y(ori_ori_n333_));
  AOI220     o317(.A0(ori_ori_n333_), .A1(x0), .B0(ori_ori_n331_), .B1(ori_ori_n104_), .Y(ori_ori_n334_));
  AOI210     o318(.A0(ori_ori_n334_), .A1(ori_ori_n330_), .B0(ori_ori_n186_), .Y(ori_ori_n335_));
  NO3        o319(.A(ori_ori_n335_), .B(ori_ori_n327_), .C(ori_ori_n323_), .Y(ori_ori_n336_));
  NA3        o320(.A(ori_ori_n336_), .B(ori_ori_n321_), .C(ori_ori_n297_), .Y(ori_ori_n337_));
  AOI210     o321(.A0(ori_ori_n284_), .A1(ori_ori_n25_), .B0(ori_ori_n337_), .Y(ori05));
  INV        o322(.A(x6), .Y(ori_ori_n341_));
  INV        o323(.A(x1), .Y(ori_ori_n342_));
  INV        o324(.A(x3), .Y(ori_ori_n343_));
  INV        o325(.A(x2), .Y(ori_ori_n344_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  INV        m005(.A(mai_mai_n19_), .Y(mai_mai_n22_));
  NA2        m006(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n23_));
  INV        m007(.A(x5), .Y(mai_mai_n24_));
  NA2        m008(.A(x7), .B(x6), .Y(mai_mai_n25_));
  NA2        m009(.A(x8), .B(x3), .Y(mai_mai_n26_));
  NA2        m010(.A(x4), .B(x2), .Y(mai_mai_n27_));
  INV        m011(.A(mai_mai_n23_), .Y(mai_mai_n28_));
  NO2        m012(.A(x4), .B(x3), .Y(mai_mai_n29_));
  INV        m013(.A(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m014(.An(mai_mai_n22_), .B(mai_mai_n28_), .Y(mai00));
  NO2        m015(.A(x1), .B(x0), .Y(mai_mai_n32_));
  INV        m016(.A(x6), .Y(mai_mai_n33_));
  NO2        m017(.A(mai_mai_n33_), .B(mai_mai_n24_), .Y(mai_mai_n34_));
  NA2        m018(.A(x4), .B(x3), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n22_), .B(mai_mai_n35_), .Y(mai_mai_n36_));
  NO2        m020(.A(x2), .B(x0), .Y(mai_mai_n37_));
  INV        m021(.A(x3), .Y(mai_mai_n38_));
  NO2        m022(.A(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n39_));
  INV        m023(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m024(.A(mai_mai_n34_), .B(x4), .Y(mai_mai_n41_));
  OAI210     m025(.A0(mai_mai_n41_), .A1(mai_mai_n40_), .B0(mai_mai_n37_), .Y(mai_mai_n42_));
  INV        m026(.A(x4), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n44_));
  NA2        m028(.A(mai_mai_n44_), .B(x2), .Y(mai_mai_n45_));
  OAI210     m029(.A0(mai_mai_n45_), .A1(mai_mai_n20_), .B0(mai_mai_n42_), .Y(mai_mai_n46_));
  INV        m030(.A(mai_mai_n32_), .Y(mai_mai_n47_));
  INV        m031(.A(x2), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n50_));
  NA2        m034(.A(mai_mai_n50_), .B(mai_mai_n49_), .Y(mai_mai_n51_));
  OAI210     m035(.A0(mai_mai_n47_), .A1(mai_mai_n30_), .B0(mai_mai_n51_), .Y(mai_mai_n52_));
  NO3        m036(.A(mai_mai_n52_), .B(mai_mai_n46_), .C(mai_mai_n36_), .Y(mai01));
  NA2        m037(.A(x8), .B(x7), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n38_), .B(x1), .Y(mai_mai_n55_));
  INV        m039(.A(x9), .Y(mai_mai_n56_));
  NO2        m040(.A(mai_mai_n56_), .B(mai_mai_n33_), .Y(mai_mai_n57_));
  INV        m041(.A(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m042(.A(mai_mai_n58_), .B(mai_mai_n55_), .Y(mai_mai_n59_));
  NO2        m043(.A(x7), .B(x6), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n61_));
  NO2        m045(.A(x8), .B(x2), .Y(mai_mai_n62_));
  OA210      m046(.A0(mai_mai_n62_), .A1(mai_mai_n61_), .B0(mai_mai_n60_), .Y(mai_mai_n63_));
  OAI210     m047(.A0(mai_mai_n39_), .A1(mai_mai_n24_), .B0(mai_mai_n48_), .Y(mai_mai_n64_));
  OAI210     m048(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n64_), .Y(mai_mai_n65_));
  NAi31      m049(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n66_));
  NO2        m050(.A(mai_mai_n65_), .B(mai_mai_n63_), .Y(mai_mai_n67_));
  OAI210     m051(.A0(mai_mai_n67_), .A1(mai_mai_n59_), .B0(x4), .Y(mai_mai_n68_));
  NA2        m052(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n69_), .A1(mai_mai_n50_), .B0(x0), .Y(mai_mai_n70_));
  NA2        m054(.A(x5), .B(x3), .Y(mai_mai_n71_));
  NO2        m055(.A(x8), .B(x6), .Y(mai_mai_n72_));
  NO3        m056(.A(mai_mai_n71_), .B(mai_mai_n60_), .C(mai_mai_n48_), .Y(mai_mai_n73_));
  NAi21      m057(.An(x4), .B(x3), .Y(mai_mai_n74_));
  INV        m058(.A(mai_mai_n74_), .Y(mai_mai_n75_));
  NO2        m059(.A(x4), .B(x2), .Y(mai_mai_n76_));
  INV        m060(.A(x3), .Y(mai_mai_n77_));
  NO2        m061(.A(mai_mai_n74_), .B(mai_mai_n18_), .Y(mai_mai_n78_));
  NO3        m062(.A(mai_mai_n78_), .B(mai_mai_n73_), .C(mai_mai_n70_), .Y(mai_mai_n79_));
  NO3        m063(.A(mai_mai_n21_), .B(mai_mai_n38_), .C(x1), .Y(mai_mai_n80_));
  NA2        m064(.A(mai_mai_n56_), .B(mai_mai_n43_), .Y(mai_mai_n81_));
  INV        m065(.A(mai_mai_n81_), .Y(mai_mai_n82_));
  OAI210     m066(.A0(mai_mai_n80_), .A1(mai_mai_n61_), .B0(mai_mai_n82_), .Y(mai_mai_n83_));
  NA2        m067(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(mai_mai_n24_), .Y(mai_mai_n85_));
  INV        m069(.A(x8), .Y(mai_mai_n86_));
  NA2        m070(.A(x2), .B(x1), .Y(mai_mai_n87_));
  NO2        m071(.A(x2), .B(mai_mai_n85_), .Y(mai_mai_n88_));
  NO2        m072(.A(mai_mai_n88_), .B(mai_mai_n25_), .Y(mai_mai_n89_));
  AOI210     m073(.A0(mai_mai_n50_), .A1(mai_mai_n24_), .B0(mai_mai_n48_), .Y(mai_mai_n90_));
  NA2        m074(.A(mai_mai_n40_), .B(mai_mai_n43_), .Y(mai_mai_n91_));
  NO3        m075(.A(mai_mai_n91_), .B(mai_mai_n90_), .C(mai_mai_n89_), .Y(mai_mai_n92_));
  NA2        m076(.A(x4), .B(mai_mai_n38_), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n43_), .B(mai_mai_n48_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n93_), .B(x1), .Y(mai_mai_n95_));
  NO2        m079(.A(x3), .B(x2), .Y(mai_mai_n96_));
  NA3        m080(.A(mai_mai_n96_), .B(mai_mai_n25_), .C(mai_mai_n24_), .Y(mai_mai_n97_));
  INV        m081(.A(mai_mai_n97_), .Y(mai_mai_n98_));
  NA2        m082(.A(mai_mai_n48_), .B(x1), .Y(mai_mai_n99_));
  OAI210     m083(.A0(mai_mai_n99_), .A1(mai_mai_n35_), .B0(mai_mai_n17_), .Y(mai_mai_n100_));
  NO4        m084(.A(mai_mai_n100_), .B(mai_mai_n98_), .C(mai_mai_n95_), .D(mai_mai_n92_), .Y(mai_mai_n101_));
  AO220      m085(.A0(mai_mai_n101_), .A1(mai_mai_n83_), .B0(mai_mai_n79_), .B1(mai_mai_n68_), .Y(mai02));
  NO2        m086(.A(x3), .B(mai_mai_n48_), .Y(mai_mai_n103_));
  NO2        m087(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n104_));
  NA2        m088(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n105_));
  NA2        m089(.A(mai_mai_n38_), .B(x0), .Y(mai_mai_n106_));
  OAI210     m090(.A0(mai_mai_n81_), .A1(mai_mai_n105_), .B0(mai_mai_n106_), .Y(mai_mai_n107_));
  AOI220     m091(.A0(mai_mai_n107_), .A1(mai_mai_n104_), .B0(mai_mai_n103_), .B1(x4), .Y(mai_mai_n108_));
  NO3        m092(.A(mai_mai_n108_), .B(x7), .C(x5), .Y(mai_mai_n109_));
  NA2        m093(.A(x9), .B(x2), .Y(mai_mai_n110_));
  OR2        m094(.A(x8), .B(x0), .Y(mai_mai_n111_));
  INV        m095(.A(mai_mai_n111_), .Y(mai_mai_n112_));
  NAi21      m096(.An(x2), .B(x8), .Y(mai_mai_n113_));
  OAI210     m097(.A0(mai_mai_n110_), .A1(x7), .B0(mai_mai_n112_), .Y(mai_mai_n114_));
  NO2        m098(.A(x4), .B(x1), .Y(mai_mai_n115_));
  NA3        m099(.A(mai_mai_n115_), .B(mai_mai_n114_), .C(mai_mai_n54_), .Y(mai_mai_n116_));
  NOi21      m100(.An(x0), .B(x1), .Y(mai_mai_n117_));
  NO3        m101(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n118_));
  NOi21      m102(.An(x0), .B(x4), .Y(mai_mai_n119_));
  NAi21      m103(.An(x8), .B(x7), .Y(mai_mai_n120_));
  NO2        m104(.A(mai_mai_n120_), .B(mai_mai_n56_), .Y(mai_mai_n121_));
  AOI220     m105(.A0(mai_mai_n121_), .A1(mai_mai_n119_), .B0(mai_mai_n118_), .B1(mai_mai_n117_), .Y(mai_mai_n122_));
  AOI210     m106(.A0(mai_mai_n122_), .A1(mai_mai_n116_), .B0(mai_mai_n71_), .Y(mai_mai_n123_));
  NO2        m107(.A(x5), .B(mai_mai_n43_), .Y(mai_mai_n124_));
  NA2        m108(.A(mai_mai_n32_), .B(mai_mai_n124_), .Y(mai_mai_n125_));
  NAi21      m109(.An(x0), .B(x4), .Y(mai_mai_n126_));
  NO2        m110(.A(mai_mai_n126_), .B(x1), .Y(mai_mai_n127_));
  NO2        m111(.A(x7), .B(x0), .Y(mai_mai_n128_));
  NO2        m112(.A(mai_mai_n76_), .B(mai_mai_n94_), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n129_), .B(x3), .Y(mai_mai_n130_));
  OAI210     m114(.A0(mai_mai_n128_), .A1(mai_mai_n127_), .B0(mai_mai_n130_), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n21_), .B(mai_mai_n38_), .Y(mai_mai_n132_));
  NA2        m116(.A(x5), .B(x0), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n134_));
  NA3        m118(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n132_), .Y(mai_mai_n135_));
  NA4        m119(.A(mai_mai_n135_), .B(mai_mai_n131_), .C(mai_mai_n125_), .D(mai_mai_n33_), .Y(mai_mai_n136_));
  NO3        m120(.A(mai_mai_n136_), .B(mai_mai_n123_), .C(mai_mai_n109_), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n27_), .B(mai_mai_n24_), .Y(mai_mai_n138_));
  AOI220     m122(.A0(mai_mai_n117_), .A1(mai_mai_n138_), .B0(mai_mai_n61_), .B1(mai_mai_n17_), .Y(mai_mai_n139_));
  NO3        m123(.A(mai_mai_n139_), .B(mai_mai_n54_), .C(mai_mai_n56_), .Y(mai_mai_n140_));
  NO2        m124(.A(mai_mai_n93_), .B(x5), .Y(mai_mai_n141_));
  NO2        m125(.A(x9), .B(x7), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n38_), .B(x2), .Y(mai_mai_n143_));
  INV        m127(.A(x7), .Y(mai_mai_n144_));
  NA2        m128(.A(x5), .B(x1), .Y(mai_mai_n145_));
  INV        m129(.A(mai_mai_n145_), .Y(mai_mai_n146_));
  AOI210     m130(.A0(mai_mai_n146_), .A1(mai_mai_n119_), .B0(mai_mai_n33_), .Y(mai_mai_n147_));
  NO2        m131(.A(mai_mai_n56_), .B(mai_mai_n86_), .Y(mai_mai_n148_));
  NO3        m132(.A(x2), .B(mai_mai_n148_), .C(mai_mai_n43_), .Y(mai_mai_n149_));
  NA2        m133(.A(mai_mai_n149_), .B(mai_mai_n61_), .Y(mai_mai_n150_));
  NA2        m134(.A(mai_mai_n150_), .B(mai_mai_n147_), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n151_), .B(mai_mai_n140_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n152_), .B(mai_mai_n137_), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n133_), .B(mai_mai_n129_), .Y(mai_mai_n154_));
  NA2        m138(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n155_));
  NA2        m139(.A(mai_mai_n24_), .B(mai_mai_n17_), .Y(mai_mai_n156_));
  NA3        m140(.A(mai_mai_n156_), .B(mai_mai_n155_), .C(mai_mai_n23_), .Y(mai_mai_n157_));
  AN2        m141(.A(mai_mai_n157_), .B(mai_mai_n134_), .Y(mai_mai_n158_));
  NA2        m142(.A(x8), .B(x0), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n144_), .B(mai_mai_n24_), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n117_), .B(x4), .Y(mai_mai_n161_));
  NA2        m145(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  AOI210     m146(.A0(mai_mai_n159_), .A1(x1), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  NA2        m147(.A(x2), .B(x0), .Y(mai_mai_n164_));
  NA2        m148(.A(x4), .B(x1), .Y(mai_mai_n165_));
  NAi21      m149(.An(mai_mai_n115_), .B(mai_mai_n165_), .Y(mai_mai_n166_));
  NOi31      m150(.An(mai_mai_n166_), .B(x5), .C(mai_mai_n164_), .Y(mai_mai_n167_));
  NO4        m151(.A(mai_mai_n167_), .B(mai_mai_n163_), .C(mai_mai_n158_), .D(mai_mai_n154_), .Y(mai_mai_n168_));
  NO2        m152(.A(mai_mai_n168_), .B(mai_mai_n38_), .Y(mai_mai_n169_));
  NO2        m153(.A(mai_mai_n157_), .B(mai_mai_n69_), .Y(mai_mai_n170_));
  INV        m154(.A(mai_mai_n124_), .Y(mai_mai_n171_));
  NO2        m155(.A(mai_mai_n99_), .B(mai_mai_n17_), .Y(mai_mai_n172_));
  NA3        m156(.A(mai_mai_n166_), .B(mai_mai_n171_), .C(mai_mai_n37_), .Y(mai_mai_n173_));
  OAI210     m157(.A0(mai_mai_n156_), .A1(mai_mai_n129_), .B0(mai_mai_n173_), .Y(mai_mai_n174_));
  NO2        m158(.A(mai_mai_n174_), .B(mai_mai_n170_), .Y(mai_mai_n175_));
  NO2        m159(.A(mai_mai_n175_), .B(x3), .Y(mai_mai_n176_));
  NO3        m160(.A(mai_mai_n176_), .B(mai_mai_n169_), .C(mai_mai_n153_), .Y(mai03));
  NO2        m161(.A(mai_mai_n43_), .B(x3), .Y(mai_mai_n178_));
  NO2        m162(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n48_), .B(x1), .Y(mai_mai_n180_));
  OAI210     m164(.A0(mai_mai_n180_), .A1(mai_mai_n24_), .B0(mai_mai_n57_), .Y(mai_mai_n181_));
  OAI220     m165(.A0(mai_mai_n181_), .A1(mai_mai_n17_), .B0(x6), .B1(mai_mai_n99_), .Y(mai_mai_n182_));
  NA2        m166(.A(mai_mai_n182_), .B(mai_mai_n178_), .Y(mai_mai_n183_));
  NO2        m167(.A(mai_mai_n71_), .B(x6), .Y(mai_mai_n184_));
  NA2        m168(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n185_));
  NO2        m169(.A(mai_mai_n185_), .B(x4), .Y(mai_mai_n186_));
  NO2        m170(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n187_));
  AO220      m171(.A0(mai_mai_n187_), .A1(mai_mai_n186_), .B0(mai_mai_n184_), .B1(mai_mai_n49_), .Y(mai_mai_n188_));
  NA2        m172(.A(mai_mai_n188_), .B(mai_mai_n56_), .Y(mai_mai_n189_));
  NA2        m173(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n190_));
  NO2        m174(.A(x5), .B(x1), .Y(mai_mai_n191_));
  AOI220     m175(.A0(mai_mai_n191_), .A1(mai_mai_n17_), .B0(mai_mai_n96_), .B1(x5), .Y(mai_mai_n192_));
  NO2        m176(.A(mai_mai_n190_), .B(mai_mai_n155_), .Y(mai_mai_n193_));
  NO3        m177(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n194_));
  OAI210     m178(.A0(mai_mai_n192_), .A1(mai_mai_n58_), .B0(mai_mai_n398_), .Y(mai_mai_n195_));
  NA2        m179(.A(mai_mai_n195_), .B(mai_mai_n43_), .Y(mai_mai_n196_));
  NA3        m180(.A(mai_mai_n196_), .B(mai_mai_n189_), .C(mai_mai_n183_), .Y(mai_mai_n197_));
  NO2        m181(.A(mai_mai_n43_), .B(mai_mai_n38_), .Y(mai_mai_n198_));
  NO2        m182(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n199_));
  NO2        m183(.A(mai_mai_n76_), .B(mai_mai_n144_), .Y(mai_mai_n200_));
  OR2        m184(.A(mai_mai_n200_), .B(mai_mai_n160_), .Y(mai_mai_n201_));
  NA2        m185(.A(mai_mai_n38_), .B(mai_mai_n48_), .Y(mai_mai_n202_));
  NO3        m186(.A(mai_mai_n165_), .B(mai_mai_n56_), .C(x6), .Y(mai_mai_n203_));
  AOI220     m187(.A0(mai_mai_n203_), .A1(mai_mai_n17_), .B0(mai_mai_n134_), .B1(mai_mai_n85_), .Y(mai_mai_n204_));
  NA2        m188(.A(x6), .B(mai_mai_n43_), .Y(mai_mai_n205_));
  OAI210     m189(.A0(mai_mai_n112_), .A1(mai_mai_n72_), .B0(x4), .Y(mai_mai_n206_));
  AOI210     m190(.A0(mai_mai_n206_), .A1(mai_mai_n205_), .B0(mai_mai_n71_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n56_), .B(x6), .Y(mai_mai_n208_));
  NO2        m192(.A(mai_mai_n145_), .B(mai_mai_n38_), .Y(mai_mai_n209_));
  OAI210     m193(.A0(mai_mai_n209_), .A1(mai_mai_n193_), .B0(mai_mai_n208_), .Y(mai_mai_n210_));
  NA2        m194(.A(mai_mai_n179_), .B(mai_mai_n127_), .Y(mai_mai_n211_));
  OAI210     m195(.A0(mai_mai_n86_), .A1(mai_mai_n33_), .B0(mai_mai_n61_), .Y(mai_mai_n212_));
  NA3        m196(.A(mai_mai_n212_), .B(mai_mai_n211_), .C(mai_mai_n210_), .Y(mai_mai_n213_));
  OAI210     m197(.A0(mai_mai_n213_), .A1(mai_mai_n207_), .B0(x2), .Y(mai_mai_n214_));
  NA3        m198(.A(mai_mai_n214_), .B(mai_mai_n204_), .C(mai_mai_n201_), .Y(mai_mai_n215_));
  AOI210     m199(.A0(mai_mai_n197_), .A1(x8), .B0(mai_mai_n215_), .Y(mai_mai_n216_));
  NO2        m200(.A(mai_mai_n86_), .B(x3), .Y(mai_mai_n217_));
  NA2        m201(.A(mai_mai_n217_), .B(mai_mai_n186_), .Y(mai_mai_n218_));
  NO3        m202(.A(mai_mai_n84_), .B(mai_mai_n72_), .C(mai_mai_n24_), .Y(mai_mai_n219_));
  INV        m203(.A(mai_mai_n219_), .Y(mai_mai_n220_));
  AOI210     m204(.A0(mai_mai_n220_), .A1(mai_mai_n218_), .B0(x2), .Y(mai_mai_n221_));
  NO2        m205(.A(x4), .B(mai_mai_n48_), .Y(mai_mai_n222_));
  AOI220     m206(.A0(mai_mai_n186_), .A1(mai_mai_n172_), .B0(mai_mai_n222_), .B1(mai_mai_n61_), .Y(mai_mai_n223_));
  NA3        m207(.A(mai_mai_n24_), .B(x3), .C(x2), .Y(mai_mai_n224_));
  NO2        m208(.A(mai_mai_n133_), .B(x9), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n38_), .B(mai_mai_n17_), .Y(mai_mai_n226_));
  NA2        m210(.A(mai_mai_n225_), .B(mai_mai_n115_), .Y(mai_mai_n227_));
  NA2        m211(.A(mai_mai_n190_), .B(x6), .Y(mai_mai_n228_));
  NA2        m212(.A(mai_mai_n228_), .B(mai_mai_n138_), .Y(mai_mai_n229_));
  NA4        m213(.A(mai_mai_n229_), .B(mai_mai_n227_), .C(mai_mai_n223_), .D(mai_mai_n144_), .Y(mai_mai_n230_));
  NA2        m214(.A(mai_mai_n179_), .B(mai_mai_n199_), .Y(mai_mai_n231_));
  NO2        m215(.A(x9), .B(x6), .Y(mai_mai_n232_));
  NO2        m216(.A(mai_mai_n133_), .B(mai_mai_n18_), .Y(mai_mai_n233_));
  NAi21      m217(.An(mai_mai_n233_), .B(mai_mai_n224_), .Y(mai_mai_n234_));
  NAi21      m218(.An(x1), .B(x4), .Y(mai_mai_n235_));
  AOI210     m219(.A0(x3), .A1(x2), .B0(mai_mai_n43_), .Y(mai_mai_n236_));
  OAI210     m220(.A0(mai_mai_n133_), .A1(x3), .B0(mai_mai_n236_), .Y(mai_mai_n237_));
  AOI220     m221(.A0(mai_mai_n237_), .A1(mai_mai_n235_), .B0(mai_mai_n234_), .B1(mai_mai_n232_), .Y(mai_mai_n238_));
  NA2        m222(.A(mai_mai_n238_), .B(mai_mai_n231_), .Y(mai_mai_n239_));
  NA2        m223(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n240_));
  NO2        m224(.A(mai_mai_n240_), .B(mai_mai_n231_), .Y(mai_mai_n241_));
  NO3        m225(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n242_));
  INV        m226(.A(mai_mai_n242_), .Y(mai_mai_n243_));
  OAI220     m227(.A0(mai_mai_n243_), .A1(mai_mai_n38_), .B0(mai_mai_n161_), .B1(mai_mai_n41_), .Y(mai_mai_n244_));
  OAI210     m228(.A0(mai_mai_n244_), .A1(mai_mai_n241_), .B0(mai_mai_n239_), .Y(mai_mai_n245_));
  NA2        m229(.A(x9), .B(mai_mai_n38_), .Y(mai_mai_n246_));
  NO2        m230(.A(mai_mai_n246_), .B(mai_mai_n185_), .Y(mai_mai_n247_));
  OR2        m231(.A(mai_mai_n247_), .B(mai_mai_n184_), .Y(mai_mai_n248_));
  NA2        m232(.A(mai_mai_n248_), .B(mai_mai_n37_), .Y(mai_mai_n249_));
  AOI210     m233(.A0(mai_mai_n249_), .A1(mai_mai_n245_), .B0(x8), .Y(mai_mai_n250_));
  NA2        m234(.A(mai_mai_n233_), .B(x6), .Y(mai_mai_n251_));
  NA2        m235(.A(x0), .B(mai_mai_n20_), .Y(mai_mai_n252_));
  AOI210     m236(.A0(mai_mai_n252_), .A1(mai_mai_n251_), .B0(mai_mai_n202_), .Y(mai_mai_n253_));
  NO4        m237(.A(mai_mai_n253_), .B(mai_mai_n250_), .C(mai_mai_n230_), .D(mai_mai_n221_), .Y(mai_mai_n254_));
  NO2        m238(.A(mai_mai_n148_), .B(x1), .Y(mai_mai_n255_));
  NO2        m239(.A(x3), .B(mai_mai_n33_), .Y(mai_mai_n256_));
  NA2        m240(.A(mai_mai_n256_), .B(x2), .Y(mai_mai_n257_));
  OAI210     m241(.A0(x0), .A1(x6), .B0(mai_mai_n39_), .Y(mai_mai_n258_));
  AOI210     m242(.A0(mai_mai_n258_), .A1(mai_mai_n257_), .B0(mai_mai_n171_), .Y(mai_mai_n259_));
  NA3        m243(.A(x0), .B(mai_mai_n191_), .C(mai_mai_n35_), .Y(mai_mai_n260_));
  AOI210     m244(.A0(mai_mai_n33_), .A1(mai_mai_n48_), .B0(x0), .Y(mai_mai_n261_));
  NA3        m245(.A(mai_mai_n261_), .B(mai_mai_n146_), .C(mai_mai_n30_), .Y(mai_mai_n262_));
  NA2        m246(.A(x3), .B(x2), .Y(mai_mai_n263_));
  AOI220     m247(.A0(mai_mai_n263_), .A1(mai_mai_n202_), .B0(mai_mai_n262_), .B1(mai_mai_n260_), .Y(mai_mai_n264_));
  NAi21      m248(.An(x4), .B(x0), .Y(mai_mai_n265_));
  NO3        m249(.A(mai_mai_n265_), .B(mai_mai_n39_), .C(x2), .Y(mai_mai_n266_));
  OAI210     m250(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  OAI220     m251(.A0(mai_mai_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n268_));
  NO2        m252(.A(x9), .B(x8), .Y(mai_mai_n269_));
  NA3        m253(.A(mai_mai_n269_), .B(mai_mai_n33_), .C(mai_mai_n48_), .Y(mai_mai_n270_));
  OAI210     m254(.A0(mai_mai_n261_), .A1(x0), .B0(mai_mai_n270_), .Y(mai_mai_n271_));
  AOI220     m255(.A0(mai_mai_n271_), .A1(mai_mai_n75_), .B0(mai_mai_n268_), .B1(mai_mai_n29_), .Y(mai_mai_n272_));
  AOI210     m256(.A0(mai_mai_n272_), .A1(mai_mai_n267_), .B0(mai_mai_n24_), .Y(mai_mai_n273_));
  NA3        m257(.A(mai_mai_n33_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n274_));
  OAI210     m258(.A0(mai_mai_n261_), .A1(x0), .B0(mai_mai_n274_), .Y(mai_mai_n275_));
  NA2        m259(.A(mai_mai_n33_), .B(mai_mai_n38_), .Y(mai_mai_n276_));
  AN2        m260(.A(mai_mai_n275_), .B(mai_mai_n141_), .Y(mai_mai_n277_));
  NO4        m261(.A(mai_mai_n277_), .B(mai_mai_n273_), .C(mai_mai_n264_), .D(mai_mai_n259_), .Y(mai_mai_n278_));
  OAI210     m262(.A0(mai_mai_n254_), .A1(mai_mai_n216_), .B0(mai_mai_n278_), .Y(mai04));
  OAI210     m263(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n280_));
  NA3        m264(.A(mai_mai_n280_), .B(mai_mai_n242_), .C(mai_mai_n77_), .Y(mai_mai_n281_));
  NO2        m265(.A(x2), .B(x1), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n226_), .A1(mai_mai_n282_), .B0(mai_mai_n33_), .Y(mai_mai_n283_));
  NO2        m267(.A(mai_mai_n282_), .B(mai_mai_n265_), .Y(mai_mai_n284_));
  INV        m268(.A(mai_mai_n105_), .Y(mai_mai_n285_));
  OAI210     m269(.A0(mai_mai_n285_), .A1(mai_mai_n284_), .B0(mai_mai_n217_), .Y(mai_mai_n286_));
  NO2        m270(.A(mai_mai_n240_), .B(mai_mai_n84_), .Y(mai_mai_n287_));
  NO2        m271(.A(mai_mai_n287_), .B(mai_mai_n33_), .Y(mai_mai_n288_));
  NO2        m272(.A(mai_mai_n263_), .B(mai_mai_n187_), .Y(mai_mai_n289_));
  NA2        m273(.A(x9), .B(x0), .Y(mai_mai_n290_));
  AOI210     m274(.A0(mai_mai_n84_), .A1(mai_mai_n69_), .B0(mai_mai_n290_), .Y(mai_mai_n291_));
  OAI210     m275(.A0(mai_mai_n291_), .A1(mai_mai_n289_), .B0(mai_mai_n86_), .Y(mai_mai_n292_));
  NA3        m276(.A(mai_mai_n292_), .B(mai_mai_n288_), .C(mai_mai_n286_), .Y(mai_mai_n293_));
  NA2        m277(.A(mai_mai_n293_), .B(mai_mai_n283_), .Y(mai_mai_n294_));
  AOI210     m278(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n295_));
  OAI220     m279(.A0(mai_mai_n295_), .A1(mai_mai_n276_), .B0(mai_mai_n240_), .B1(mai_mai_n274_), .Y(mai_mai_n296_));
  INV        m280(.A(mai_mai_n296_), .Y(mai_mai_n297_));
  NA2        m281(.A(mai_mai_n287_), .B(mai_mai_n86_), .Y(mai_mai_n298_));
  NA2        m282(.A(mai_mai_n298_), .B(mai_mai_n297_), .Y(mai_mai_n299_));
  OAI210     m283(.A0(mai_mai_n104_), .A1(x3), .B0(mai_mai_n266_), .Y(mai_mai_n300_));
  NA2        m284(.A(mai_mai_n300_), .B(mai_mai_n144_), .Y(mai_mai_n301_));
  AOI210     m285(.A0(mai_mai_n299_), .A1(x4), .B0(mai_mai_n301_), .Y(mai_mai_n302_));
  NA2        m286(.A(mai_mai_n284_), .B(mai_mai_n86_), .Y(mai_mai_n303_));
  NOi21      m287(.An(x4), .B(x0), .Y(mai_mai_n304_));
  XO2        m288(.A(x4), .B(x0), .Y(mai_mai_n305_));
  AOI210     m289(.A0(x2), .A1(x8), .B0(mai_mai_n304_), .Y(mai_mai_n306_));
  AOI210     m290(.A0(mai_mai_n306_), .A1(mai_mai_n303_), .B0(x3), .Y(mai_mai_n307_));
  INV        m291(.A(mai_mai_n87_), .Y(mai_mai_n308_));
  NO2        m292(.A(mai_mai_n86_), .B(x4), .Y(mai_mai_n309_));
  NO3        m293(.A(mai_mai_n305_), .B(mai_mai_n148_), .C(x2), .Y(mai_mai_n310_));
  NO2        m294(.A(mai_mai_n27_), .B(mai_mai_n23_), .Y(mai_mai_n311_));
  NO2        m295(.A(mai_mai_n311_), .B(mai_mai_n310_), .Y(mai_mai_n312_));
  NA2        m296(.A(mai_mai_n312_), .B(x6), .Y(mai_mai_n313_));
  NO2        m297(.A(mai_mai_n38_), .B(x0), .Y(mai_mai_n314_));
  BUFFER     m298(.A(mai_mai_n314_), .Y(mai_mai_n315_));
  AOI220     m299(.A0(mai_mai_n48_), .A1(mai_mai_n315_), .B0(mai_mai_n396_), .B1(mai_mai_n55_), .Y(mai_mai_n316_));
  NO2        m300(.A(mai_mai_n32_), .B(x2), .Y(mai_mai_n317_));
  NOi21      m301(.An(mai_mai_n115_), .B(mai_mai_n26_), .Y(mai_mai_n318_));
  INV        m302(.A(mai_mai_n318_), .Y(mai_mai_n319_));
  OAI210     m303(.A0(mai_mai_n316_), .A1(mai_mai_n56_), .B0(mai_mai_n319_), .Y(mai_mai_n320_));
  OAI220     m304(.A0(mai_mai_n320_), .A1(x6), .B0(mai_mai_n313_), .B1(mai_mai_n307_), .Y(mai_mai_n321_));
  AO220      m305(.A0(x7), .A1(mai_mai_n321_), .B0(mai_mai_n302_), .B1(mai_mai_n294_), .Y(mai_mai_n322_));
  NA2        m306(.A(mai_mai_n317_), .B(x6), .Y(mai_mai_n323_));
  AOI210     m307(.A0(x6), .A1(x1), .B0(mai_mai_n143_), .Y(mai_mai_n324_));
  NA2        m308(.A(mai_mai_n309_), .B(x0), .Y(mai_mai_n325_));
  NA2        m309(.A(mai_mai_n76_), .B(x6), .Y(mai_mai_n326_));
  OAI210     m310(.A0(mai_mai_n325_), .A1(mai_mai_n324_), .B0(mai_mai_n326_), .Y(mai_mai_n327_));
  AOI220     m311(.A0(mai_mai_n327_), .A1(mai_mai_n323_), .B0(mai_mai_n194_), .B1(mai_mai_n44_), .Y(mai_mai_n328_));
  NA3        m312(.A(mai_mai_n328_), .B(mai_mai_n322_), .C(mai_mai_n281_), .Y(mai_mai_n329_));
  NA3        m313(.A(mai_mai_n104_), .B(mai_mai_n178_), .C(mai_mai_n144_), .Y(mai_mai_n330_));
  AO220      m314(.A0(x4), .A1(mai_mai_n142_), .B0(mai_mai_n103_), .B1(x4), .Y(mai_mai_n331_));
  NA3        m315(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n332_));
  NO2        m316(.A(mai_mai_n332_), .B(mai_mai_n308_), .Y(mai_mai_n333_));
  AOI210     m317(.A0(mai_mai_n331_), .A1(mai_mai_n112_), .B0(mai_mai_n333_), .Y(mai_mai_n334_));
  AOI210     m318(.A0(mai_mai_n334_), .A1(mai_mai_n330_), .B0(mai_mai_n24_), .Y(mai_mai_n335_));
  NA3        m319(.A(x8), .B(mai_mai_n198_), .C(x0), .Y(mai_mai_n336_));
  INV        m320(.A(mai_mai_n187_), .Y(mai_mai_n337_));
  NO2        m321(.A(mai_mai_n337_), .B(mai_mai_n24_), .Y(mai_mai_n338_));
  AOI210     m322(.A0(mai_mai_n113_), .A1(mai_mai_n111_), .B0(mai_mai_n37_), .Y(mai_mai_n339_));
  NOi21      m323(.An(mai_mai_n339_), .B(mai_mai_n165_), .Y(mai_mai_n340_));
  OAI210     m324(.A0(mai_mai_n340_), .A1(mai_mai_n338_), .B0(mai_mai_n142_), .Y(mai_mai_n341_));
  NAi31      m325(.An(mai_mai_n45_), .B(mai_mai_n255_), .C(mai_mai_n160_), .Y(mai_mai_n342_));
  NA3        m326(.A(mai_mai_n342_), .B(mai_mai_n341_), .C(mai_mai_n336_), .Y(mai_mai_n343_));
  OAI210     m327(.A0(mai_mai_n343_), .A1(mai_mai_n335_), .B0(x6), .Y(mai_mai_n344_));
  INV        m328(.A(mai_mai_n128_), .Y(mai_mai_n345_));
  AOI210     m329(.A0(mai_mai_n35_), .A1(mai_mai_n30_), .B0(mai_mai_n345_), .Y(mai_mai_n346_));
  AOI220     m330(.A0(mai_mai_n397_), .A1(mai_mai_n198_), .B0(mai_mai_n178_), .B1(mai_mai_n144_), .Y(mai_mai_n347_));
  AOI210     m331(.A0(mai_mai_n121_), .A1(mai_mai_n222_), .B0(x1), .Y(mai_mai_n348_));
  OAI210     m332(.A0(mai_mai_n347_), .A1(x8), .B0(mai_mai_n348_), .Y(mai_mai_n349_));
  NO4        m333(.A(mai_mai_n120_), .B(mai_mai_n265_), .C(x9), .D(x2), .Y(mai_mai_n350_));
  NOi21      m334(.An(mai_mai_n118_), .B(mai_mai_n164_), .Y(mai_mai_n351_));
  NO3        m335(.A(mai_mai_n351_), .B(mai_mai_n350_), .C(mai_mai_n18_), .Y(mai_mai_n352_));
  NO3        m336(.A(x9), .B(mai_mai_n144_), .C(x0), .Y(mai_mai_n353_));
  NA2        m337(.A(mai_mai_n353_), .B(mai_mai_n217_), .Y(mai_mai_n354_));
  NA2        m338(.A(mai_mai_n354_), .B(mai_mai_n352_), .Y(mai_mai_n355_));
  OAI210     m339(.A0(mai_mai_n349_), .A1(mai_mai_n346_), .B0(mai_mai_n355_), .Y(mai_mai_n356_));
  NOi31      m340(.An(mai_mai_n397_), .B(mai_mai_n30_), .C(x8), .Y(mai_mai_n357_));
  INV        m341(.A(mai_mai_n126_), .Y(mai_mai_n358_));
  NO3        m342(.A(mai_mai_n358_), .B(mai_mai_n118_), .C(mai_mai_n38_), .Y(mai_mai_n359_));
  NOi31      m343(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n360_));
  AOI220     m344(.A0(mai_mai_n360_), .A1(mai_mai_n304_), .B0(mai_mai_n119_), .B1(x3), .Y(mai_mai_n361_));
  AOI210     m345(.A0(mai_mai_n235_), .A1(mai_mai_n54_), .B0(mai_mai_n117_), .Y(mai_mai_n362_));
  OAI210     m346(.A0(mai_mai_n362_), .A1(x3), .B0(mai_mai_n361_), .Y(mai_mai_n363_));
  NO3        m347(.A(mai_mai_n363_), .B(mai_mai_n359_), .C(x2), .Y(mai_mai_n364_));
  OAI220     m348(.A0(mai_mai_n305_), .A1(mai_mai_n269_), .B0(mai_mai_n265_), .B1(mai_mai_n38_), .Y(mai_mai_n365_));
  AOI210     m349(.A0(x9), .A1(mai_mai_n43_), .B0(mai_mai_n332_), .Y(mai_mai_n366_));
  AOI220     m350(.A0(mai_mai_n366_), .A1(mai_mai_n86_), .B0(mai_mai_n365_), .B1(mai_mai_n144_), .Y(mai_mai_n367_));
  NO2        m351(.A(mai_mai_n367_), .B(mai_mai_n48_), .Y(mai_mai_n368_));
  NO3        m352(.A(mai_mai_n368_), .B(mai_mai_n364_), .C(mai_mai_n357_), .Y(mai_mai_n369_));
  AOI210     m353(.A0(mai_mai_n369_), .A1(mai_mai_n356_), .B0(mai_mai_n24_), .Y(mai_mai_n370_));
  NO3        m354(.A(mai_mai_n56_), .B(x4), .C(x1), .Y(mai_mai_n371_));
  NO3        m355(.A(mai_mai_n62_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n372_));
  AOI220     m356(.A0(mai_mai_n372_), .A1(mai_mai_n236_), .B0(mai_mai_n371_), .B1(mai_mai_n339_), .Y(mai_mai_n373_));
  NO2        m357(.A(mai_mai_n373_), .B(mai_mai_n96_), .Y(mai_mai_n374_));
  NO3        m358(.A(mai_mai_n240_), .B(mai_mai_n159_), .C(mai_mai_n35_), .Y(mai_mai_n375_));
  OAI210     m359(.A0(mai_mai_n375_), .A1(mai_mai_n374_), .B0(x7), .Y(mai_mai_n376_));
  NA2        m360(.A(mai_mai_n143_), .B(mai_mai_n127_), .Y(mai_mai_n377_));
  NA2        m361(.A(mai_mai_n377_), .B(mai_mai_n376_), .Y(mai_mai_n378_));
  OAI210     m362(.A0(mai_mai_n378_), .A1(mai_mai_n370_), .B0(mai_mai_n33_), .Y(mai_mai_n379_));
  NO2        m363(.A(mai_mai_n353_), .B(mai_mai_n187_), .Y(mai_mai_n380_));
  NO4        m364(.A(mai_mai_n380_), .B(mai_mai_n71_), .C(x4), .D(mai_mai_n48_), .Y(mai_mai_n381_));
  NA2        m365(.A(mai_mai_n314_), .B(mai_mai_n160_), .Y(mai_mai_n382_));
  OAI220     m366(.A0(mai_mai_n246_), .A1(x2), .B0(mai_mai_n145_), .B1(mai_mai_n38_), .Y(mai_mai_n383_));
  AOI210     m367(.A0(x2), .A1(mai_mai_n26_), .B0(mai_mai_n66_), .Y(mai_mai_n384_));
  NO3        m368(.A(mai_mai_n360_), .B(x3), .C(mai_mai_n48_), .Y(mai_mai_n385_));
  NO2        m369(.A(mai_mai_n385_), .B(mai_mai_n384_), .Y(mai_mai_n386_));
  INV        m370(.A(mai_mai_n386_), .Y(mai_mai_n387_));
  AOI220     m371(.A0(mai_mai_n387_), .A1(x0), .B0(mai_mai_n383_), .B1(mai_mai_n128_), .Y(mai_mai_n388_));
  AOI210     m372(.A0(mai_mai_n388_), .A1(mai_mai_n382_), .B0(mai_mai_n205_), .Y(mai_mai_n389_));
  NO3        m373(.A(mai_mai_n99_), .B(mai_mai_n54_), .C(mai_mai_n30_), .Y(mai_mai_n390_));
  NO3        m374(.A(mai_mai_n390_), .B(mai_mai_n389_), .C(mai_mai_n381_), .Y(mai_mai_n391_));
  NA3        m375(.A(mai_mai_n391_), .B(mai_mai_n379_), .C(mai_mai_n344_), .Y(mai_mai_n392_));
  AOI210     m376(.A0(mai_mai_n329_), .A1(mai_mai_n24_), .B0(mai_mai_n392_), .Y(mai05));
  INV        m377(.A(mai_mai_n164_), .Y(mai_mai_n396_));
  INV        m378(.A(x0), .Y(mai_mai_n397_));
  INV        m379(.A(mai_mai_n194_), .Y(mai_mai_n398_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  BUFFER     u005(.A(men_men_n20_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO3        u012(.A(men_men_n28_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  AN2        u021(.A(x8), .B(x7), .Y(men_men_n38_));
  NA3        u022(.A(men_men_n38_), .B(men_men_n37_), .C(men_men_n35_), .Y(men_men_n39_));
  NA2        u023(.A(x4), .B(x3), .Y(men_men_n40_));
  AOI210     u024(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n40_), .Y(men_men_n41_));
  NO2        u025(.A(x2), .B(x0), .Y(men_men_n42_));
  INV        u026(.A(x3), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n44_));
  INV        u028(.A(men_men_n44_), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n37_), .B(x4), .Y(men_men_n46_));
  OAI210     u030(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n42_), .Y(men_men_n47_));
  INV        u031(.A(x4), .Y(men_men_n48_));
  NO2        u032(.A(men_men_n48_), .B(men_men_n17_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(x2), .Y(men_men_n50_));
  OAI210     u034(.A0(men_men_n50_), .A1(men_men_n20_), .B0(men_men_n47_), .Y(men_men_n51_));
  NA2        u035(.A(men_men_n38_), .B(men_men_n37_), .Y(men_men_n52_));
  AOI220     u036(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n53_));
  INV        u037(.A(x2), .Y(men_men_n54_));
  NO2        u038(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n56_));
  NA2        u040(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  OAI210     u041(.A0(men_men_n53_), .A1(men_men_n32_), .B0(men_men_n57_), .Y(men_men_n58_));
  NO3        u042(.A(men_men_n58_), .B(men_men_n51_), .C(men_men_n41_), .Y(men01));
  NA2        u043(.A(x8), .B(x7), .Y(men_men_n60_));
  NA2        u044(.A(men_men_n43_), .B(x1), .Y(men_men_n61_));
  INV        u045(.A(x9), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n62_), .B(men_men_n36_), .Y(men_men_n63_));
  NO2        u047(.A(men_men_n61_), .B(men_men_n60_), .Y(men_men_n64_));
  NO2        u048(.A(x7), .B(x6), .Y(men_men_n65_));
  NO2        u049(.A(men_men_n61_), .B(x5), .Y(men_men_n66_));
  NO2        u050(.A(x8), .B(x2), .Y(men_men_n67_));
  NO2        u051(.A(x2), .B(x1), .Y(men_men_n68_));
  OA210      u052(.A0(men_men_n68_), .A1(men_men_n66_), .B0(men_men_n65_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n56_), .A1(men_men_n20_), .B0(men_men_n70_), .Y(men_men_n71_));
  NAi31      u055(.An(x1), .B(x9), .C(x5), .Y(men_men_n72_));
  OAI220     u056(.A0(men_men_n72_), .A1(men_men_n43_), .B0(men_men_n71_), .B1(men_men_n69_), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n64_), .B0(x4), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n48_), .B(x2), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n56_), .B0(x0), .Y(men_men_n76_));
  NA2        u060(.A(x5), .B(x3), .Y(men_men_n77_));
  NO2        u061(.A(x8), .B(x6), .Y(men_men_n78_));
  NO3        u062(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n54_), .Y(men_men_n79_));
  NAi21      u063(.An(x4), .B(x3), .Y(men_men_n80_));
  INV        u064(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n81_), .B(men_men_n22_), .Y(men_men_n82_));
  NO2        u066(.A(x4), .B(x2), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n83_), .B(x3), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n82_), .C(men_men_n18_), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n79_), .C(men_men_n76_), .Y(men_men_n86_));
  NO3        u070(.A(x6), .B(men_men_n43_), .C(x1), .Y(men_men_n87_));
  NA2        u071(.A(men_men_n87_), .B(men_men_n48_), .Y(men_men_n88_));
  NA2        u072(.A(x3), .B(men_men_n18_), .Y(men_men_n89_));
  NO2        u073(.A(men_men_n89_), .B(men_men_n25_), .Y(men_men_n90_));
  INV        u074(.A(x8), .Y(men_men_n91_));
  NA2        u075(.A(x2), .B(x1), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n91_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n90_), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n26_), .Y(men_men_n95_));
  AOI210     u079(.A0(men_men_n56_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n96_));
  OAI210     u080(.A0(men_men_n45_), .A1(men_men_n37_), .B0(men_men_n48_), .Y(men_men_n97_));
  NO3        u081(.A(men_men_n97_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n98_));
  NA2        u082(.A(x4), .B(men_men_n43_), .Y(men_men_n99_));
  NO2        u083(.A(men_men_n48_), .B(men_men_n54_), .Y(men_men_n100_));
  OAI210     u084(.A0(men_men_n100_), .A1(men_men_n43_), .B0(men_men_n18_), .Y(men_men_n101_));
  AOI210     u085(.A0(men_men_n99_), .A1(men_men_n52_), .B0(men_men_n101_), .Y(men_men_n102_));
  NO2        u086(.A(x3), .B(x2), .Y(men_men_n103_));
  NA2        u087(.A(men_men_n103_), .B(men_men_n25_), .Y(men_men_n104_));
  AOI210     u088(.A0(x8), .A1(x6), .B0(men_men_n104_), .Y(men_men_n105_));
  NA2        u089(.A(men_men_n54_), .B(x1), .Y(men_men_n106_));
  OAI210     u090(.A0(men_men_n106_), .A1(men_men_n40_), .B0(men_men_n17_), .Y(men_men_n107_));
  NO4        u091(.A(men_men_n107_), .B(men_men_n105_), .C(men_men_n102_), .D(men_men_n98_), .Y(men_men_n108_));
  AO220      u092(.A0(men_men_n108_), .A1(men_men_n88_), .B0(men_men_n86_), .B1(men_men_n74_), .Y(men02));
  NO2        u093(.A(x3), .B(men_men_n54_), .Y(men_men_n110_));
  AOI220     u094(.A0(men_men_n54_), .A1(x1), .B0(men_men_n110_), .B1(x4), .Y(men_men_n111_));
  NO3        u095(.A(men_men_n111_), .B(x7), .C(x5), .Y(men_men_n112_));
  NA2        u096(.A(x9), .B(x2), .Y(men_men_n113_));
  OR2        u097(.A(x8), .B(x0), .Y(men_men_n114_));
  NAi21      u098(.An(x2), .B(x8), .Y(men_men_n115_));
  NO2        u099(.A(x4), .B(x1), .Y(men_men_n116_));
  NOi21      u100(.An(x0), .B(x1), .Y(men_men_n117_));
  NO3        u101(.A(x9), .B(x8), .C(x7), .Y(men_men_n118_));
  NOi21      u102(.An(x0), .B(x4), .Y(men_men_n119_));
  NO2        u103(.A(x8), .B(men_men_n62_), .Y(men_men_n120_));
  AOI220     u104(.A0(men_men_n120_), .A1(men_men_n119_), .B0(men_men_n118_), .B1(men_men_n117_), .Y(men_men_n121_));
  NO2        u105(.A(men_men_n121_), .B(men_men_n77_), .Y(men_men_n122_));
  NO2        u106(.A(x5), .B(men_men_n48_), .Y(men_men_n123_));
  NA2        u107(.A(x2), .B(men_men_n18_), .Y(men_men_n124_));
  AOI210     u108(.A0(men_men_n124_), .A1(men_men_n106_), .B0(x3), .Y(men_men_n125_));
  OAI210     u109(.A0(men_men_n125_), .A1(men_men_n35_), .B0(men_men_n123_), .Y(men_men_n126_));
  NAi21      u110(.An(x0), .B(x4), .Y(men_men_n127_));
  NO2        u111(.A(men_men_n127_), .B(x1), .Y(men_men_n128_));
  NO2        u112(.A(x7), .B(x0), .Y(men_men_n129_));
  NO2        u113(.A(men_men_n83_), .B(men_men_n100_), .Y(men_men_n130_));
  NO2        u114(.A(men_men_n130_), .B(x3), .Y(men_men_n131_));
  OAI210     u115(.A0(men_men_n129_), .A1(men_men_n128_), .B0(men_men_n131_), .Y(men_men_n132_));
  NA2        u116(.A(x5), .B(x0), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n48_), .B(x2), .Y(men_men_n134_));
  NA3        u118(.A(men_men_n132_), .B(men_men_n126_), .C(men_men_n36_), .Y(men_men_n135_));
  NO3        u119(.A(men_men_n135_), .B(men_men_n122_), .C(men_men_n112_), .Y(men_men_n136_));
  NO3        u120(.A(men_men_n77_), .B(men_men_n75_), .C(men_men_n24_), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n138_));
  AOI220     u122(.A0(men_men_n117_), .A1(men_men_n138_), .B0(men_men_n66_), .B1(men_men_n17_), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n139_), .B(men_men_n60_), .Y(men_men_n140_));
  NA2        u124(.A(x7), .B(x3), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n99_), .B(x5), .Y(men_men_n142_));
  NO2        u126(.A(x9), .B(x7), .Y(men_men_n143_));
  NOi21      u127(.An(x8), .B(x0), .Y(men_men_n144_));
  OA210      u128(.A0(men_men_n143_), .A1(x1), .B0(men_men_n144_), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n43_), .B(x2), .Y(men_men_n146_));
  INV        u130(.A(x7), .Y(men_men_n147_));
  NA2        u131(.A(men_men_n147_), .B(men_men_n18_), .Y(men_men_n148_));
  AOI220     u132(.A0(men_men_n148_), .A1(men_men_n146_), .B0(men_men_n110_), .B1(men_men_n38_), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n25_), .B(x4), .Y(men_men_n150_));
  NO2        u134(.A(men_men_n150_), .B(men_men_n119_), .Y(men_men_n151_));
  NO2        u135(.A(men_men_n151_), .B(men_men_n149_), .Y(men_men_n152_));
  AOI210     u136(.A0(men_men_n145_), .A1(men_men_n142_), .B0(men_men_n152_), .Y(men_men_n153_));
  OAI210     u137(.A0(men_men_n141_), .A1(men_men_n50_), .B0(men_men_n153_), .Y(men_men_n154_));
  NA2        u138(.A(x5), .B(x1), .Y(men_men_n155_));
  INV        u139(.A(men_men_n155_), .Y(men_men_n156_));
  AOI210     u140(.A0(men_men_n156_), .A1(men_men_n119_), .B0(men_men_n36_), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n62_), .B(men_men_n91_), .Y(men_men_n158_));
  NAi21      u142(.An(x2), .B(x7), .Y(men_men_n159_));
  NAi31      u143(.An(men_men_n77_), .B(men_men_n38_), .C(men_men_n35_), .Y(men_men_n160_));
  NA2        u144(.A(men_men_n160_), .B(men_men_n157_), .Y(men_men_n161_));
  NO4        u145(.A(men_men_n161_), .B(men_men_n154_), .C(men_men_n140_), .D(men_men_n137_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n162_), .B(men_men_n136_), .Y(men_men_n163_));
  NO2        u147(.A(men_men_n133_), .B(men_men_n130_), .Y(men_men_n164_));
  NA2        u148(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n165_));
  NA2        u149(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n166_));
  NA3        u150(.A(men_men_n166_), .B(men_men_n165_), .C(men_men_n24_), .Y(men_men_n167_));
  AN2        u151(.A(men_men_n167_), .B(men_men_n134_), .Y(men_men_n168_));
  NA2        u152(.A(x8), .B(x0), .Y(men_men_n169_));
  NO2        u153(.A(men_men_n147_), .B(men_men_n25_), .Y(men_men_n170_));
  NO2        u154(.A(men_men_n117_), .B(x4), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  AOI210     u156(.A0(men_men_n169_), .A1(men_men_n124_), .B0(men_men_n172_), .Y(men_men_n173_));
  NA2        u157(.A(x2), .B(x0), .Y(men_men_n174_));
  NA2        u158(.A(x4), .B(x1), .Y(men_men_n175_));
  NAi21      u159(.An(men_men_n116_), .B(men_men_n175_), .Y(men_men_n176_));
  NOi31      u160(.An(men_men_n176_), .B(men_men_n150_), .C(men_men_n174_), .Y(men_men_n177_));
  NO4        u161(.A(men_men_n177_), .B(men_men_n173_), .C(men_men_n168_), .D(men_men_n164_), .Y(men_men_n178_));
  NO2        u162(.A(men_men_n178_), .B(men_men_n43_), .Y(men_men_n179_));
  NO2        u163(.A(men_men_n167_), .B(men_men_n75_), .Y(men_men_n180_));
  INV        u164(.A(men_men_n123_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n106_), .B(men_men_n17_), .Y(men_men_n182_));
  AOI210     u166(.A0(men_men_n35_), .A1(men_men_n91_), .B0(men_men_n182_), .Y(men_men_n183_));
  NO3        u167(.A(men_men_n183_), .B(men_men_n181_), .C(x7), .Y(men_men_n184_));
  NA3        u168(.A(men_men_n176_), .B(men_men_n181_), .C(men_men_n42_), .Y(men_men_n185_));
  OAI210     u169(.A0(men_men_n166_), .A1(men_men_n130_), .B0(men_men_n185_), .Y(men_men_n186_));
  NO3        u170(.A(men_men_n186_), .B(men_men_n184_), .C(men_men_n180_), .Y(men_men_n187_));
  NO2        u171(.A(men_men_n187_), .B(x3), .Y(men_men_n188_));
  NO3        u172(.A(men_men_n188_), .B(men_men_n179_), .C(men_men_n163_), .Y(men03));
  NO2        u173(.A(men_men_n48_), .B(x3), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n54_), .B(x1), .Y(men_men_n191_));
  NA2        u175(.A(men_men_n63_), .B(men_men_n190_), .Y(men_men_n192_));
  NA2        u176(.A(x6), .B(men_men_n25_), .Y(men_men_n193_));
  NO2        u177(.A(men_men_n193_), .B(x4), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n18_), .B(x0), .Y(men_men_n195_));
  NA2        u179(.A(x3), .B(men_men_n17_), .Y(men_men_n196_));
  NO2        u180(.A(men_men_n196_), .B(men_men_n193_), .Y(men_men_n197_));
  NA2        u181(.A(x9), .B(men_men_n54_), .Y(men_men_n198_));
  NA2        u182(.A(men_men_n198_), .B(x4), .Y(men_men_n199_));
  NA2        u183(.A(men_men_n193_), .B(men_men_n80_), .Y(men_men_n200_));
  AOI210     u184(.A0(men_men_n25_), .A1(x3), .B0(men_men_n174_), .Y(men_men_n201_));
  AOI220     u185(.A0(men_men_n201_), .A1(men_men_n200_), .B0(men_men_n199_), .B1(men_men_n197_), .Y(men_men_n202_));
  NO2        u186(.A(x5), .B(x1), .Y(men_men_n203_));
  AOI220     u187(.A0(men_men_n203_), .A1(men_men_n17_), .B0(men_men_n103_), .B1(x5), .Y(men_men_n204_));
  NO2        u188(.A(men_men_n196_), .B(men_men_n165_), .Y(men_men_n205_));
  NO2        u189(.A(men_men_n204_), .B(men_men_n36_), .Y(men_men_n206_));
  NA2        u190(.A(men_men_n206_), .B(men_men_n48_), .Y(men_men_n207_));
  NA3        u191(.A(men_men_n207_), .B(men_men_n202_), .C(men_men_n192_), .Y(men_men_n208_));
  NO2        u192(.A(men_men_n48_), .B(men_men_n43_), .Y(men_men_n209_));
  NA2        u193(.A(men_men_n209_), .B(men_men_n19_), .Y(men_men_n210_));
  NO2        u194(.A(x3), .B(men_men_n17_), .Y(men_men_n211_));
  NO2        u195(.A(men_men_n211_), .B(x6), .Y(men_men_n212_));
  NOi21      u196(.An(men_men_n83_), .B(men_men_n212_), .Y(men_men_n213_));
  NA2        u197(.A(men_men_n62_), .B(men_men_n91_), .Y(men_men_n214_));
  NA3        u198(.A(men_men_n214_), .B(men_men_n211_), .C(x6), .Y(men_men_n215_));
  AOI210     u199(.A0(men_men_n215_), .A1(men_men_n213_), .B0(men_men_n147_), .Y(men_men_n216_));
  AO210      u200(.A0(men_men_n216_), .A1(men_men_n210_), .B0(men_men_n170_), .Y(men_men_n217_));
  NA2        u201(.A(men_men_n43_), .B(men_men_n54_), .Y(men_men_n218_));
  INV        u202(.A(men_men_n166_), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n175_), .B(x6), .Y(men_men_n220_));
  AOI220     u204(.A0(men_men_n220_), .A1(men_men_n219_), .B0(men_men_n134_), .B1(men_men_n90_), .Y(men_men_n221_));
  NA2        u205(.A(x6), .B(men_men_n48_), .Y(men_men_n222_));
  NO2        u206(.A(men_men_n155_), .B(men_men_n43_), .Y(men_men_n223_));
  OAI210     u207(.A0(men_men_n223_), .A1(men_men_n205_), .B0(men_men_n401_), .Y(men_men_n224_));
  NA2        u208(.A(x5), .B(men_men_n128_), .Y(men_men_n225_));
  NA3        u209(.A(men_men_n196_), .B(men_men_n123_), .C(x6), .Y(men_men_n226_));
  OAI210     u210(.A0(men_men_n91_), .A1(men_men_n36_), .B0(men_men_n66_), .Y(men_men_n227_));
  NA4        u211(.A(men_men_n227_), .B(men_men_n226_), .C(men_men_n225_), .D(men_men_n224_), .Y(men_men_n228_));
  NA2        u212(.A(men_men_n228_), .B(x2), .Y(men_men_n229_));
  NA3        u213(.A(men_men_n229_), .B(men_men_n221_), .C(men_men_n217_), .Y(men_men_n230_));
  AOI210     u214(.A0(men_men_n208_), .A1(x8), .B0(men_men_n230_), .Y(men_men_n231_));
  INV        u215(.A(men_men_n194_), .Y(men_men_n232_));
  NO3        u216(.A(men_men_n89_), .B(men_men_n78_), .C(men_men_n25_), .Y(men_men_n233_));
  AOI210     u217(.A0(men_men_n212_), .A1(men_men_n150_), .B0(men_men_n233_), .Y(men_men_n234_));
  AOI210     u218(.A0(men_men_n234_), .A1(men_men_n232_), .B0(x2), .Y(men_men_n235_));
  NO2        u219(.A(x4), .B(men_men_n54_), .Y(men_men_n236_));
  AOI220     u220(.A0(men_men_n194_), .A1(men_men_n182_), .B0(men_men_n236_), .B1(men_men_n66_), .Y(men_men_n237_));
  NA2        u221(.A(men_men_n62_), .B(x6), .Y(men_men_n238_));
  NA3        u222(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n239_));
  AOI210     u223(.A0(men_men_n239_), .A1(men_men_n133_), .B0(men_men_n238_), .Y(men_men_n240_));
  NA2        u224(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n241_));
  NO2        u225(.A(men_men_n241_), .B(men_men_n25_), .Y(men_men_n242_));
  OAI210     u226(.A0(men_men_n242_), .A1(men_men_n240_), .B0(men_men_n116_), .Y(men_men_n243_));
  NA2        u227(.A(men_men_n196_), .B(x6), .Y(men_men_n244_));
  NO2        u228(.A(men_men_n196_), .B(x6), .Y(men_men_n245_));
  INV        u229(.A(men_men_n245_), .Y(men_men_n246_));
  NA3        u230(.A(men_men_n246_), .B(men_men_n244_), .C(men_men_n138_), .Y(men_men_n247_));
  NA4        u231(.A(men_men_n247_), .B(men_men_n243_), .C(men_men_n237_), .D(men_men_n147_), .Y(men_men_n248_));
  NA2        u232(.A(x5), .B(men_men_n211_), .Y(men_men_n249_));
  INV        u233(.A(x6), .Y(men_men_n250_));
  NO2        u234(.A(men_men_n133_), .B(men_men_n18_), .Y(men_men_n251_));
  NAi21      u235(.An(men_men_n251_), .B(men_men_n239_), .Y(men_men_n252_));
  NAi21      u236(.An(x1), .B(x4), .Y(men_men_n253_));
  AOI210     u237(.A0(x3), .A1(x2), .B0(men_men_n48_), .Y(men_men_n254_));
  OAI210     u238(.A0(men_men_n133_), .A1(x3), .B0(men_men_n254_), .Y(men_men_n255_));
  AOI220     u239(.A0(men_men_n255_), .A1(men_men_n253_), .B0(men_men_n252_), .B1(men_men_n250_), .Y(men_men_n256_));
  NA2        u240(.A(men_men_n256_), .B(men_men_n249_), .Y(men_men_n257_));
  INV        u241(.A(men_men_n249_), .Y(men_men_n258_));
  NO2        u242(.A(x6), .B(x0), .Y(men_men_n259_));
  NA2        u243(.A(men_men_n106_), .B(men_men_n25_), .Y(men_men_n260_));
  NA2        u244(.A(x6), .B(x2), .Y(men_men_n261_));
  NO2        u245(.A(men_men_n261_), .B(men_men_n165_), .Y(men_men_n262_));
  AOI210     u246(.A0(men_men_n260_), .A1(men_men_n259_), .B0(men_men_n262_), .Y(men_men_n263_));
  OAI220     u247(.A0(men_men_n263_), .A1(men_men_n43_), .B0(men_men_n171_), .B1(men_men_n46_), .Y(men_men_n264_));
  OAI210     u248(.A0(men_men_n264_), .A1(men_men_n258_), .B0(men_men_n257_), .Y(men_men_n265_));
  NA2        u249(.A(x4), .B(x0), .Y(men_men_n266_));
  NO3        u250(.A(men_men_n72_), .B(men_men_n266_), .C(x6), .Y(men_men_n267_));
  INV        u251(.A(men_men_n267_), .Y(men_men_n268_));
  AOI210     u252(.A0(men_men_n268_), .A1(men_men_n265_), .B0(x8), .Y(men_men_n269_));
  INV        u253(.A(men_men_n169_), .Y(men_men_n270_));
  OAI210     u254(.A0(men_men_n270_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n271_));
  AOI210     u255(.A0(men_men_n271_), .A1(men_men_n238_), .B0(men_men_n218_), .Y(men_men_n272_));
  NO4        u256(.A(men_men_n272_), .B(men_men_n269_), .C(men_men_n248_), .D(men_men_n235_), .Y(men_men_n273_));
  NO2        u257(.A(men_men_n158_), .B(x1), .Y(men_men_n274_));
  NO3        u258(.A(men_men_n274_), .B(x3), .C(men_men_n36_), .Y(men_men_n275_));
  OAI210     u259(.A0(men_men_n275_), .A1(men_men_n245_), .B0(x2), .Y(men_men_n276_));
  OAI210     u260(.A0(men_men_n270_), .A1(x6), .B0(men_men_n44_), .Y(men_men_n277_));
  AOI210     u261(.A0(men_men_n277_), .A1(men_men_n276_), .B0(men_men_n181_), .Y(men_men_n278_));
  NOi21      u262(.An(men_men_n261_), .B(men_men_n17_), .Y(men_men_n279_));
  NA3        u263(.A(men_men_n279_), .B(men_men_n203_), .C(men_men_n40_), .Y(men_men_n280_));
  NA3        u264(.A(men_men_n405_), .B(men_men_n156_), .C(men_men_n32_), .Y(men_men_n281_));
  NA2        u265(.A(x3), .B(x2), .Y(men_men_n282_));
  AOI220     u266(.A0(men_men_n282_), .A1(men_men_n218_), .B0(men_men_n281_), .B1(men_men_n280_), .Y(men_men_n283_));
  NAi21      u267(.An(x4), .B(x0), .Y(men_men_n284_));
  NO3        u268(.A(men_men_n284_), .B(men_men_n44_), .C(x2), .Y(men_men_n285_));
  OAI210     u269(.A0(x6), .A1(men_men_n18_), .B0(men_men_n285_), .Y(men_men_n286_));
  OAI220     u270(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n287_));
  NA2        u271(.A(men_men_n36_), .B(men_men_n54_), .Y(men_men_n288_));
  OAI210     u272(.A0(men_men_n405_), .A1(men_men_n279_), .B0(men_men_n288_), .Y(men_men_n289_));
  AOI220     u273(.A0(men_men_n289_), .A1(men_men_n81_), .B0(men_men_n287_), .B1(men_men_n31_), .Y(men_men_n290_));
  AOI210     u274(.A0(men_men_n290_), .A1(men_men_n286_), .B0(men_men_n25_), .Y(men_men_n291_));
  INV        u275(.A(men_men_n205_), .Y(men_men_n292_));
  NA2        u276(.A(men_men_n36_), .B(men_men_n43_), .Y(men_men_n293_));
  OR2        u277(.A(men_men_n293_), .B(men_men_n266_), .Y(men_men_n294_));
  OAI220     u278(.A0(men_men_n294_), .A1(men_men_n155_), .B0(men_men_n222_), .B1(men_men_n292_), .Y(men_men_n295_));
  NO4        u279(.A(men_men_n295_), .B(men_men_n291_), .C(men_men_n283_), .D(men_men_n278_), .Y(men_men_n296_));
  OAI210     u280(.A0(men_men_n273_), .A1(men_men_n231_), .B0(men_men_n296_), .Y(men04));
  NA2        u281(.A(men_men_n259_), .B(men_men_n84_), .Y(men_men_n298_));
  INV        u282(.A(men_men_n284_), .Y(men_men_n299_));
  NA3        u283(.A(men_men_n89_), .B(x6), .C(men_men_n284_), .Y(men_men_n300_));
  NA2        u284(.A(men_men_n300_), .B(x6), .Y(men_men_n301_));
  NO2        u285(.A(men_men_n198_), .B(x3), .Y(men_men_n302_));
  NO3        u286(.A(men_men_n238_), .B(men_men_n115_), .C(men_men_n18_), .Y(men_men_n303_));
  NO2        u287(.A(men_men_n303_), .B(men_men_n302_), .Y(men_men_n304_));
  OAI210     u288(.A0(men_men_n114_), .A1(men_men_n106_), .B0(men_men_n169_), .Y(men_men_n305_));
  NA3        u289(.A(men_men_n305_), .B(x6), .C(x3), .Y(men_men_n306_));
  INV        u290(.A(men_men_n293_), .Y(men_men_n307_));
  AOI210     u291(.A0(men_men_n18_), .A1(men_men_n63_), .B0(men_men_n307_), .Y(men_men_n308_));
  NA4        u292(.A(men_men_n403_), .B(men_men_n308_), .C(men_men_n306_), .D(men_men_n304_), .Y(men_men_n309_));
  OAI210     u293(.A0(x1), .A1(x3), .B0(men_men_n285_), .Y(men_men_n310_));
  NA3        u294(.A(men_men_n214_), .B(x1), .C(men_men_n83_), .Y(men_men_n311_));
  NA3        u295(.A(men_men_n311_), .B(men_men_n310_), .C(men_men_n147_), .Y(men_men_n312_));
  AOI210     u296(.A0(men_men_n309_), .A1(x4), .B0(men_men_n312_), .Y(men_men_n313_));
  NA3        u297(.A(men_men_n299_), .B(men_men_n198_), .C(men_men_n91_), .Y(men_men_n314_));
  XO2        u298(.A(x4), .B(x0), .Y(men_men_n315_));
  OAI210     u299(.A0(men_men_n315_), .A1(men_men_n113_), .B0(men_men_n253_), .Y(men_men_n316_));
  NA2        u300(.A(men_men_n316_), .B(x8), .Y(men_men_n317_));
  AOI210     u301(.A0(men_men_n317_), .A1(men_men_n314_), .B0(x3), .Y(men_men_n318_));
  INV        u302(.A(men_men_n92_), .Y(men_men_n319_));
  AOI220     u303(.A0(x8), .A1(men_men_n44_), .B0(men_men_n119_), .B1(men_men_n319_), .Y(men_men_n320_));
  NO3        u304(.A(men_men_n315_), .B(men_men_n158_), .C(x2), .Y(men_men_n321_));
  NO3        u305(.A(men_men_n214_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n322_));
  NO2        u306(.A(men_men_n322_), .B(men_men_n321_), .Y(men_men_n323_));
  NA4        u307(.A(men_men_n323_), .B(men_men_n320_), .C(men_men_n210_), .D(x6), .Y(men_men_n324_));
  NO2        u308(.A(men_men_n144_), .B(men_men_n106_), .Y(men_men_n325_));
  INV        u309(.A(men_men_n325_), .Y(men_men_n326_));
  NO2        u310(.A(men_men_n144_), .B(men_men_n80_), .Y(men_men_n327_));
  NO2        u311(.A(men_men_n35_), .B(x2), .Y(men_men_n328_));
  NA2        u312(.A(men_men_n328_), .B(men_men_n327_), .Y(men_men_n329_));
  OAI210     u313(.A0(men_men_n326_), .A1(men_men_n62_), .B0(men_men_n329_), .Y(men_men_n330_));
  OAI220     u314(.A0(men_men_n330_), .A1(x6), .B0(men_men_n324_), .B1(men_men_n318_), .Y(men_men_n331_));
  OAI210     u315(.A0(men_men_n63_), .A1(men_men_n48_), .B0(men_men_n42_), .Y(men_men_n332_));
  OAI210     u316(.A0(men_men_n332_), .A1(men_men_n91_), .B0(men_men_n294_), .Y(men_men_n333_));
  AOI210     u317(.A0(men_men_n333_), .A1(men_men_n18_), .B0(men_men_n147_), .Y(men_men_n334_));
  AO220      u318(.A0(men_men_n334_), .A1(men_men_n331_), .B0(men_men_n313_), .B1(men_men_n301_), .Y(men_men_n335_));
  NA2        u319(.A(men_men_n335_), .B(men_men_n298_), .Y(men_men_n336_));
  NA3        u320(.A(x2), .B(men_men_n190_), .C(men_men_n147_), .Y(men_men_n337_));
  NA2        u321(.A(men_men_n209_), .B(x0), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n338_), .B(men_men_n198_), .Y(men_men_n339_));
  INV        u323(.A(men_men_n339_), .Y(men_men_n340_));
  AOI210     u324(.A0(men_men_n340_), .A1(men_men_n337_), .B0(men_men_n25_), .Y(men_men_n341_));
  OAI210     u325(.A0(men_men_n190_), .A1(men_men_n67_), .B0(men_men_n195_), .Y(men_men_n342_));
  NA3        u326(.A(men_men_n191_), .B(men_men_n211_), .C(x8), .Y(men_men_n343_));
  AOI210     u327(.A0(men_men_n343_), .A1(men_men_n342_), .B0(men_men_n25_), .Y(men_men_n344_));
  AOI210     u328(.A0(men_men_n115_), .A1(men_men_n114_), .B0(men_men_n42_), .Y(men_men_n345_));
  NOi31      u329(.An(men_men_n345_), .B(x3), .C(men_men_n175_), .Y(men_men_n346_));
  OAI210     u330(.A0(men_men_n346_), .A1(men_men_n344_), .B0(men_men_n143_), .Y(men_men_n347_));
  INV        u331(.A(men_men_n347_), .Y(men_men_n348_));
  OAI210     u332(.A0(men_men_n348_), .A1(men_men_n341_), .B0(x6), .Y(men_men_n349_));
  AOI210     u333(.A0(men_men_n402_), .A1(x0), .B0(men_men_n32_), .Y(men_men_n350_));
  NA2        u334(.A(men_men_n190_), .B(men_men_n147_), .Y(men_men_n351_));
  AOI210     u335(.A0(men_men_n120_), .A1(men_men_n236_), .B0(x1), .Y(men_men_n352_));
  OAI210     u336(.A0(men_men_n351_), .A1(x8), .B0(men_men_n352_), .Y(men_men_n353_));
  NAi31      u337(.An(x2), .B(x8), .C(x0), .Y(men_men_n354_));
  OAI210     u338(.A0(men_men_n354_), .A1(x4), .B0(men_men_n159_), .Y(men_men_n355_));
  NA3        u339(.A(men_men_n355_), .B(men_men_n141_), .C(x9), .Y(men_men_n356_));
  NO4        u340(.A(x8), .B(men_men_n284_), .C(x9), .D(x2), .Y(men_men_n357_));
  NOi21      u341(.An(men_men_n118_), .B(men_men_n174_), .Y(men_men_n358_));
  NO3        u342(.A(men_men_n358_), .B(men_men_n357_), .C(men_men_n18_), .Y(men_men_n359_));
  NA2        u343(.A(men_men_n327_), .B(men_men_n147_), .Y(men_men_n360_));
  NA4        u344(.A(men_men_n360_), .B(men_men_n359_), .C(men_men_n356_), .D(men_men_n50_), .Y(men_men_n361_));
  OAI210     u345(.A0(men_men_n353_), .A1(men_men_n350_), .B0(men_men_n361_), .Y(men_men_n362_));
  AOI210     u346(.A0(men_men_n38_), .A1(x9), .B0(men_men_n127_), .Y(men_men_n363_));
  NO3        u347(.A(men_men_n363_), .B(men_men_n118_), .C(men_men_n43_), .Y(men_men_n364_));
  AOI210     u348(.A0(men_men_n253_), .A1(men_men_n60_), .B0(men_men_n117_), .Y(men_men_n365_));
  NO2        u349(.A(men_men_n365_), .B(x3), .Y(men_men_n366_));
  NO3        u350(.A(men_men_n366_), .B(men_men_n364_), .C(x2), .Y(men_men_n367_));
  INV        u351(.A(men_men_n367_), .Y(men_men_n368_));
  AOI210     u352(.A0(men_men_n368_), .A1(men_men_n362_), .B0(men_men_n25_), .Y(men_men_n369_));
  NA4        u353(.A(men_men_n31_), .B(men_men_n91_), .C(x2), .D(men_men_n17_), .Y(men_men_n370_));
  NO3        u354(.A(men_men_n67_), .B(men_men_n18_), .C(x0), .Y(men_men_n371_));
  AOI220     u355(.A0(men_men_n371_), .A1(men_men_n254_), .B0(men_men_n404_), .B1(men_men_n345_), .Y(men_men_n372_));
  NO2        u356(.A(men_men_n372_), .B(men_men_n103_), .Y(men_men_n373_));
  NA2        u357(.A(men_men_n373_), .B(x7), .Y(men_men_n374_));
  NA2        u358(.A(men_men_n214_), .B(x7), .Y(men_men_n375_));
  NA3        u359(.A(men_men_n375_), .B(men_men_n146_), .C(men_men_n128_), .Y(men_men_n376_));
  NA3        u360(.A(men_men_n376_), .B(men_men_n374_), .C(men_men_n370_), .Y(men_men_n377_));
  OAI210     u361(.A0(men_men_n377_), .A1(men_men_n369_), .B0(men_men_n36_), .Y(men_men_n378_));
  NA2        u362(.A(men_men_n241_), .B(men_men_n21_), .Y(men_men_n379_));
  NO2        u363(.A(men_men_n155_), .B(men_men_n129_), .Y(men_men_n380_));
  NA2        u364(.A(men_men_n380_), .B(men_men_n379_), .Y(men_men_n381_));
  AOI210     u365(.A0(men_men_n381_), .A1(men_men_n160_), .B0(men_men_n28_), .Y(men_men_n382_));
  AOI220     u366(.A0(x3), .A1(men_men_n91_), .B0(men_men_n144_), .B1(men_men_n191_), .Y(men_men_n383_));
  NA3        u367(.A(men_men_n383_), .B(men_men_n354_), .C(men_men_n89_), .Y(men_men_n384_));
  NA2        u368(.A(men_men_n384_), .B(men_men_n170_), .Y(men_men_n385_));
  NA2        u369(.A(x3), .B(men_men_n54_), .Y(men_men_n386_));
  AOI210     u370(.A0(men_men_n159_), .A1(men_men_n27_), .B0(men_men_n72_), .Y(men_men_n387_));
  OAI210     u371(.A0(men_men_n143_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n388_));
  NO2        u372(.A(x3), .B(men_men_n54_), .Y(men_men_n389_));
  AOI210     u373(.A0(men_men_n389_), .A1(men_men_n388_), .B0(men_men_n387_), .Y(men_men_n390_));
  OAI210     u374(.A0(men_men_n148_), .A1(men_men_n386_), .B0(men_men_n390_), .Y(men_men_n391_));
  AOI220     u375(.A0(men_men_n391_), .A1(x0), .B0(men_men_n67_), .B1(men_men_n129_), .Y(men_men_n392_));
  AOI210     u376(.A0(men_men_n392_), .A1(men_men_n385_), .B0(men_men_n222_), .Y(men_men_n393_));
  NA2        u377(.A(x9), .B(x5), .Y(men_men_n394_));
  NO4        u378(.A(men_men_n106_), .B(men_men_n394_), .C(men_men_n60_), .D(men_men_n32_), .Y(men_men_n395_));
  NO3        u379(.A(men_men_n395_), .B(men_men_n393_), .C(men_men_n382_), .Y(men_men_n396_));
  NA3        u380(.A(men_men_n396_), .B(men_men_n378_), .C(men_men_n349_), .Y(men_men_n397_));
  AOI210     u381(.A0(men_men_n336_), .A1(men_men_n25_), .B0(men_men_n397_), .Y(men05));
  INV        u382(.A(x6), .Y(men_men_n401_));
  INV        u383(.A(men_men_n38_), .Y(men_men_n402_));
  INV        u384(.A(men_men_n78_), .Y(men_men_n403_));
  INV        u385(.A(x4), .Y(men_men_n404_));
  INV        u386(.A(x0), .Y(men_men_n405_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule