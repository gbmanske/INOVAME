// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n132_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1078_, new_new_n1079_,
    new_new_n1080_, new_new_n1081_, new_new_n1082_, new_new_n1083_,
    new_new_n1084_, new_new_n1085_, new_new_n1086_, new_new_n1087_,
    new_new_n1088_, new_new_n1089_, new_new_n1090_, new_new_n1091_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  OAI210     g0006(.A0(new_new_n27_), .A1(new_new_n24_), .B0(i_10_), .Y(new_new_n29_));
  NOi21      g0007(.An(i_11_), .B(i_8_), .Y(new_new_n30_));
  AO210      g0008(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n31_));
  OR2        g0009(.A(new_new_n31_), .B(new_new_n30_), .Y(new_new_n32_));
  NA2        g0010(.A(new_new_n32_), .B(new_new_n29_), .Y(new_new_n33_));
  XO2        g0011(.A(new_new_n33_), .B(new_new_n23_), .Y(new_new_n34_));
  INV        g0012(.A(i_4_), .Y(new_new_n35_));
  INV        g0013(.A(i_10_), .Y(new_new_n36_));
  NAi21      g0014(.An(i_11_), .B(i_9_), .Y(new_new_n37_));
  NO3        g0015(.A(new_new_n37_), .B(i_12_), .C(new_new_n36_), .Y(new_new_n38_));
  NOi21      g0016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g0017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g0018(.A(new_new_n35_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n34_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NA2        g0026(.A(i_7_), .B(new_new_n25_), .Y(new_new_n49_));
  NO2        g0027(.A(new_new_n47_), .B(new_new_n46_), .Y(new_new_n50_));
  NA2        g0028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g0029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g0030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA2        g0031(.A(new_new_n50_), .B(new_new_n45_), .Y(new_new_n54_));
  NA3        g0032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n55_));
  NO2        g0033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g0034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  OAI210     g0035(.A0(new_new_n57_), .A1(new_new_n56_), .B0(new_new_n55_), .Y(new_new_n58_));
  NA2        g0036(.A(new_new_n58_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g0037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g0038(.A(i_1_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA2        g0040(.A(i_1_), .B(i_10_), .Y(new_new_n63_));
  NO2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NAi21      g0042(.An(new_new_n64_), .B(new_new_n59_), .Y(new_new_n65_));
  NA2        g0043(.A(new_new_n49_), .B(i_2_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_6_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(new_new_n25_), .Y(new_new_n68_));
  INV        g0046(.A(i_0_), .Y(new_new_n69_));
  NAi21      g0047(.An(i_5_), .B(i_10_), .Y(new_new_n70_));
  NA2        g0048(.A(i_5_), .B(i_9_), .Y(new_new_n71_));
  AOI210     g0049(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n69_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n68_), .Y(new_new_n73_));
  OAI210     g0051(.A0(new_new_n72_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n74_));
  NA2        g0052(.A(i_12_), .B(i_5_), .Y(new_new_n75_));
  NA2        g0053(.A(i_2_), .B(i_8_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n56_), .Y(new_new_n77_));
  NO2        g0055(.A(i_3_), .B(i_9_), .Y(new_new_n78_));
  NO2        g0056(.A(i_3_), .B(i_7_), .Y(new_new_n79_));
  NO3        g0057(.A(new_new_n79_), .B(new_new_n78_), .C(new_new_n61_), .Y(new_new_n80_));
  INV        g0058(.A(i_6_), .Y(new_new_n81_));
  OR4        g0059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n82_));
  INV        g0060(.A(new_new_n82_), .Y(new_new_n83_));
  NO2        g0061(.A(i_2_), .B(i_7_), .Y(new_new_n84_));
  OAI210     g0062(.A0(new_new_n80_), .A1(new_new_n77_), .B0(i_2_), .Y(new_new_n85_));
  NAi21      g0063(.An(i_6_), .B(i_10_), .Y(new_new_n86_));
  NA2        g0064(.A(i_6_), .B(i_9_), .Y(new_new_n87_));
  NA2        g0065(.A(i_2_), .B(i_6_), .Y(new_new_n88_));
  AOI210     g0066(.A0(new_new_n87_), .A1(new_new_n85_), .B0(new_new_n75_), .Y(new_new_n89_));
  AN3        g0067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n90_));
  NAi21      g0068(.An(i_6_), .B(i_11_), .Y(new_new_n91_));
  NO2        g0069(.A(i_5_), .B(i_8_), .Y(new_new_n92_));
  NOi21      g0070(.An(new_new_n92_), .B(new_new_n91_), .Y(new_new_n93_));
  AOI220     g0071(.A0(new_new_n93_), .A1(new_new_n60_), .B0(new_new_n90_), .B1(new_new_n31_), .Y(new_new_n94_));
  INV        g0072(.A(i_7_), .Y(new_new_n95_));
  NA2        g0073(.A(new_new_n46_), .B(new_new_n95_), .Y(new_new_n96_));
  NO2        g0074(.A(i_0_), .B(i_5_), .Y(new_new_n97_));
  NO2        g0075(.A(new_new_n97_), .B(new_new_n81_), .Y(new_new_n98_));
  NA2        g0076(.A(i_12_), .B(i_3_), .Y(new_new_n99_));
  INV        g0077(.A(new_new_n99_), .Y(new_new_n100_));
  NA3        g0078(.A(new_new_n100_), .B(new_new_n98_), .C(new_new_n96_), .Y(new_new_n101_));
  NAi21      g0079(.An(i_7_), .B(i_11_), .Y(new_new_n102_));
  NO3        g0080(.A(new_new_n102_), .B(new_new_n86_), .C(new_new_n51_), .Y(new_new_n103_));
  AN2        g0081(.A(i_2_), .B(i_10_), .Y(new_new_n104_));
  NO2        g0082(.A(new_new_n104_), .B(i_7_), .Y(new_new_n105_));
  OR2        g0083(.A(new_new_n75_), .B(new_new_n56_), .Y(new_new_n106_));
  NO2        g0084(.A(i_8_), .B(new_new_n95_), .Y(new_new_n107_));
  NO3        g0085(.A(new_new_n107_), .B(new_new_n106_), .C(new_new_n105_), .Y(new_new_n108_));
  NA2        g0086(.A(i_12_), .B(i_7_), .Y(new_new_n109_));
  NO2        g0087(.A(new_new_n61_), .B(new_new_n26_), .Y(new_new_n110_));
  INV        g0088(.A(new_new_n110_), .Y(new_new_n111_));
  NA2        g0089(.A(i_11_), .B(i_12_), .Y(new_new_n112_));
  OAI210     g0090(.A0(new_new_n111_), .A1(new_new_n109_), .B0(new_new_n112_), .Y(new_new_n113_));
  NO2        g0091(.A(new_new_n113_), .B(new_new_n108_), .Y(new_new_n114_));
  NAi41      g0092(.An(new_new_n103_), .B(new_new_n114_), .C(new_new_n101_), .D(new_new_n94_), .Y(new_new_n115_));
  NOi21      g0093(.An(i_1_), .B(i_5_), .Y(new_new_n116_));
  NA2        g0094(.A(new_new_n116_), .B(i_11_), .Y(new_new_n117_));
  NA2        g0095(.A(new_new_n95_), .B(new_new_n36_), .Y(new_new_n118_));
  NA2        g0096(.A(i_7_), .B(new_new_n25_), .Y(new_new_n119_));
  NA2        g0097(.A(new_new_n119_), .B(new_new_n118_), .Y(new_new_n120_));
  NO2        g0098(.A(new_new_n120_), .B(new_new_n46_), .Y(new_new_n121_));
  NAi21      g0099(.An(i_3_), .B(i_8_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(new_new_n60_), .Y(new_new_n123_));
  INV        g0101(.A(new_new_n121_), .Y(new_new_n124_));
  NO2        g0102(.A(i_1_), .B(new_new_n81_), .Y(new_new_n125_));
  NO2        g0103(.A(i_6_), .B(i_5_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(i_3_), .Y(new_new_n127_));
  AO210      g0105(.A0(new_new_n127_), .A1(new_new_n47_), .B0(new_new_n125_), .Y(new_new_n128_));
  OAI220     g0106(.A0(new_new_n128_), .A1(new_new_n102_), .B0(new_new_n124_), .B1(new_new_n117_), .Y(new_new_n129_));
  NO3        g0107(.A(new_new_n129_), .B(new_new_n115_), .C(new_new_n89_), .Y(new_new_n130_));
  NA3        g0108(.A(new_new_n130_), .B(new_new_n74_), .C(new_new_n54_), .Y(men2));
  NO2        g0109(.A(new_new_n61_), .B(new_new_n36_), .Y(new_new_n132_));
  NA3        g0110(.A(new_new_n73_), .B(new_new_n66_), .C(new_new_n29_), .Y(men0));
  AN2        g0111(.A(i_8_), .B(i_7_), .Y(new_new_n134_));
  NA2        g0112(.A(new_new_n134_), .B(i_6_), .Y(new_new_n135_));
  NO2        g0113(.A(i_12_), .B(i_13_), .Y(new_new_n136_));
  NAi21      g0114(.An(i_5_), .B(i_11_), .Y(new_new_n137_));
  NOi21      g0115(.An(new_new_n136_), .B(new_new_n137_), .Y(new_new_n138_));
  NO2        g0116(.A(i_0_), .B(i_1_), .Y(new_new_n139_));
  NA2        g0117(.A(i_2_), .B(i_3_), .Y(new_new_n140_));
  NO2        g0118(.A(new_new_n140_), .B(i_4_), .Y(new_new_n141_));
  NA3        g0119(.A(new_new_n141_), .B(new_new_n139_), .C(new_new_n138_), .Y(new_new_n142_));
  OR2        g0120(.A(new_new_n142_), .B(new_new_n25_), .Y(new_new_n143_));
  AN2        g0121(.A(new_new_n136_), .B(new_new_n78_), .Y(new_new_n144_));
  NO2        g0122(.A(new_new_n144_), .B(new_new_n27_), .Y(new_new_n145_));
  NA2        g0123(.A(i_1_), .B(i_5_), .Y(new_new_n146_));
  NO2        g0124(.A(new_new_n69_), .B(new_new_n46_), .Y(new_new_n147_));
  NA2        g0125(.A(new_new_n147_), .B(new_new_n35_), .Y(new_new_n148_));
  NO3        g0126(.A(new_new_n148_), .B(new_new_n146_), .C(new_new_n145_), .Y(new_new_n149_));
  OR2        g0127(.A(i_0_), .B(i_1_), .Y(new_new_n150_));
  NO3        g0128(.A(new_new_n150_), .B(new_new_n75_), .C(i_13_), .Y(new_new_n151_));
  NAi32      g0129(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n152_));
  NAi21      g0130(.An(new_new_n152_), .B(new_new_n151_), .Y(new_new_n153_));
  NOi21      g0131(.An(i_4_), .B(i_10_), .Y(new_new_n154_));
  NA2        g0132(.A(new_new_n154_), .B(new_new_n39_), .Y(new_new_n155_));
  NO2        g0133(.A(i_3_), .B(i_5_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n69_), .B(i_2_), .C(i_1_), .Y(new_new_n157_));
  NA2        g0135(.A(new_new_n157_), .B(new_new_n156_), .Y(new_new_n158_));
  OAI210     g0136(.A0(new_new_n158_), .A1(new_new_n155_), .B0(new_new_n153_), .Y(new_new_n159_));
  NO2        g0137(.A(new_new_n159_), .B(new_new_n149_), .Y(new_new_n160_));
  AOI210     g0138(.A0(new_new_n160_), .A1(new_new_n143_), .B0(new_new_n135_), .Y(new_new_n161_));
  NA3        g0139(.A(new_new_n69_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n162_));
  NA2        g0140(.A(i_3_), .B(new_new_n48_), .Y(new_new_n163_));
  NOi21      g0141(.An(i_4_), .B(i_9_), .Y(new_new_n164_));
  NOi21      g0142(.An(i_11_), .B(i_13_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OR2        g0144(.A(new_new_n166_), .B(new_new_n163_), .Y(new_new_n167_));
  NO2        g0145(.A(i_4_), .B(i_5_), .Y(new_new_n168_));
  NAi21      g0146(.An(i_12_), .B(i_11_), .Y(new_new_n169_));
  NO2        g0147(.A(new_new_n169_), .B(i_13_), .Y(new_new_n170_));
  NA3        g0148(.A(new_new_n170_), .B(new_new_n168_), .C(new_new_n78_), .Y(new_new_n171_));
  AOI210     g0149(.A0(new_new_n171_), .A1(new_new_n167_), .B0(new_new_n162_), .Y(new_new_n172_));
  NO2        g0150(.A(new_new_n69_), .B(new_new_n61_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n173_), .B(new_new_n46_), .Y(new_new_n174_));
  NA2        g0152(.A(new_new_n35_), .B(i_5_), .Y(new_new_n175_));
  NAi31      g0153(.An(new_new_n175_), .B(new_new_n144_), .C(i_11_), .Y(new_new_n176_));
  NA2        g0154(.A(i_3_), .B(i_5_), .Y(new_new_n177_));
  OR2        g0155(.A(new_new_n177_), .B(new_new_n166_), .Y(new_new_n178_));
  AOI210     g0156(.A0(new_new_n178_), .A1(new_new_n176_), .B0(new_new_n174_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n69_), .B(i_5_), .Y(new_new_n180_));
  NO2        g0158(.A(i_13_), .B(i_10_), .Y(new_new_n181_));
  NA3        g0159(.A(new_new_n181_), .B(new_new_n180_), .C(new_new_n44_), .Y(new_new_n182_));
  NO2        g0160(.A(i_2_), .B(i_1_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n183_), .B(i_3_), .Y(new_new_n184_));
  NAi21      g0162(.An(i_4_), .B(i_12_), .Y(new_new_n185_));
  NO3        g0163(.A(new_new_n185_), .B(new_new_n184_), .C(new_new_n182_), .Y(new_new_n186_));
  NO3        g0164(.A(new_new_n186_), .B(new_new_n179_), .C(new_new_n172_), .Y(new_new_n187_));
  INV        g0165(.A(i_8_), .Y(new_new_n188_));
  NO2        g0166(.A(new_new_n188_), .B(i_7_), .Y(new_new_n189_));
  NA2        g0167(.A(new_new_n189_), .B(i_6_), .Y(new_new_n190_));
  NO3        g0168(.A(i_3_), .B(new_new_n81_), .C(new_new_n48_), .Y(new_new_n191_));
  NA2        g0169(.A(new_new_n191_), .B(new_new_n107_), .Y(new_new_n192_));
  NO3        g0170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n193_));
  NA3        g0171(.A(new_new_n193_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n194_));
  NO3        g0172(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n195_));
  OAI210     g0173(.A0(new_new_n90_), .A1(i_12_), .B0(new_new_n195_), .Y(new_new_n196_));
  AOI210     g0174(.A0(new_new_n196_), .A1(new_new_n194_), .B0(new_new_n192_), .Y(new_new_n197_));
  NO2        g0175(.A(i_3_), .B(i_8_), .Y(new_new_n198_));
  NO3        g0176(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n199_));
  NA3        g0177(.A(new_new_n199_), .B(new_new_n198_), .C(new_new_n39_), .Y(new_new_n200_));
  NO2        g0178(.A(new_new_n97_), .B(new_new_n56_), .Y(new_new_n201_));
  NO2        g0179(.A(i_13_), .B(i_9_), .Y(new_new_n202_));
  NAi21      g0180(.An(i_12_), .B(i_3_), .Y(new_new_n203_));
  OR2        g0181(.A(new_new_n203_), .B(new_new_n1081_), .Y(new_new_n204_));
  NO2        g0182(.A(new_new_n44_), .B(i_5_), .Y(new_new_n205_));
  NO3        g0183(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n206_));
  NA3        g0184(.A(new_new_n206_), .B(new_new_n205_), .C(i_10_), .Y(new_new_n207_));
  OAI220     g0185(.A0(new_new_n207_), .A1(new_new_n204_), .B0(new_new_n97_), .B1(new_new_n200_), .Y(new_new_n208_));
  AOI210     g0186(.A0(new_new_n208_), .A1(i_7_), .B0(new_new_n197_), .Y(new_new_n209_));
  OAI220     g0187(.A0(new_new_n209_), .A1(i_4_), .B0(new_new_n190_), .B1(new_new_n187_), .Y(new_new_n210_));
  NAi21      g0188(.An(i_12_), .B(i_7_), .Y(new_new_n211_));
  NA3        g0189(.A(i_13_), .B(new_new_n188_), .C(i_10_), .Y(new_new_n212_));
  NO2        g0190(.A(new_new_n212_), .B(new_new_n211_), .Y(new_new_n213_));
  NA2        g0191(.A(i_0_), .B(i_5_), .Y(new_new_n214_));
  NA2        g0192(.A(new_new_n214_), .B(new_new_n98_), .Y(new_new_n215_));
  OAI220     g0193(.A0(new_new_n215_), .A1(new_new_n184_), .B0(new_new_n174_), .B1(new_new_n127_), .Y(new_new_n216_));
  NAi31      g0194(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n35_), .B(i_13_), .Y(new_new_n218_));
  NO2        g0196(.A(new_new_n69_), .B(new_new_n26_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n46_), .B(new_new_n61_), .Y(new_new_n220_));
  NA3        g0198(.A(new_new_n220_), .B(new_new_n219_), .C(new_new_n218_), .Y(new_new_n221_));
  INV        g0199(.A(i_13_), .Y(new_new_n222_));
  NO2        g0200(.A(i_12_), .B(new_new_n222_), .Y(new_new_n223_));
  NA3        g0201(.A(new_new_n223_), .B(new_new_n193_), .C(new_new_n191_), .Y(new_new_n224_));
  OAI210     g0202(.A0(new_new_n221_), .A1(new_new_n217_), .B0(new_new_n224_), .Y(new_new_n225_));
  AOI220     g0203(.A0(new_new_n225_), .A1(new_new_n134_), .B0(new_new_n216_), .B1(new_new_n213_), .Y(new_new_n226_));
  NO2        g0204(.A(i_12_), .B(new_new_n36_), .Y(new_new_n227_));
  NO2        g0205(.A(new_new_n177_), .B(i_4_), .Y(new_new_n228_));
  NA2        g0206(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n229_));
  OR2        g0207(.A(i_8_), .B(i_7_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n230_), .B(new_new_n81_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n51_), .B(i_1_), .Y(new_new_n232_));
  NA2        g0210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  INV        g0211(.A(i_12_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n44_), .B(new_new_n234_), .Y(new_new_n235_));
  NO3        g0213(.A(new_new_n35_), .B(i_8_), .C(i_10_), .Y(new_new_n236_));
  NA2        g0214(.A(i_2_), .B(i_1_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n233_), .B(new_new_n229_), .Y(new_new_n238_));
  NO3        g0216(.A(i_11_), .B(i_7_), .C(new_new_n36_), .Y(new_new_n239_));
  NAi21      g0217(.An(i_4_), .B(i_3_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n240_), .B(new_new_n71_), .Y(new_new_n241_));
  NO2        g0219(.A(i_0_), .B(i_6_), .Y(new_new_n242_));
  NOi41      g0220(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n243_));
  NA2        g0221(.A(new_new_n243_), .B(new_new_n242_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n237_), .B(new_new_n177_), .Y(new_new_n245_));
  NAi21      g0223(.An(new_new_n244_), .B(new_new_n245_), .Y(new_new_n246_));
  INV        g0224(.A(new_new_n246_), .Y(new_new_n247_));
  AOI220     g0225(.A0(new_new_n247_), .A1(new_new_n39_), .B0(new_new_n238_), .B1(new_new_n202_), .Y(new_new_n248_));
  NO2        g0226(.A(i_11_), .B(new_new_n222_), .Y(new_new_n249_));
  NOi21      g0227(.An(i_1_), .B(i_6_), .Y(new_new_n250_));
  NAi21      g0228(.An(i_3_), .B(i_7_), .Y(new_new_n251_));
  NA2        g0229(.A(new_new_n234_), .B(i_9_), .Y(new_new_n252_));
  OR4        g0230(.A(new_new_n252_), .B(new_new_n251_), .C(new_new_n250_), .D(new_new_n180_), .Y(new_new_n253_));
  NO2        g0231(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n254_));
  NO2        g0232(.A(i_12_), .B(i_3_), .Y(new_new_n255_));
  NA2        g0233(.A(new_new_n69_), .B(i_5_), .Y(new_new_n256_));
  NA2        g0234(.A(i_3_), .B(i_9_), .Y(new_new_n257_));
  NAi21      g0235(.An(i_7_), .B(i_10_), .Y(new_new_n258_));
  NO2        g0236(.A(new_new_n258_), .B(new_new_n257_), .Y(new_new_n259_));
  NA3        g0237(.A(new_new_n259_), .B(new_new_n256_), .C(new_new_n62_), .Y(new_new_n260_));
  NA2        g0238(.A(new_new_n260_), .B(new_new_n253_), .Y(new_new_n261_));
  NA3        g0239(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n262_));
  INV        g0240(.A(new_new_n135_), .Y(new_new_n263_));
  NA2        g0241(.A(new_new_n234_), .B(i_13_), .Y(new_new_n264_));
  NO2        g0242(.A(new_new_n264_), .B(new_new_n71_), .Y(new_new_n265_));
  AOI220     g0243(.A0(new_new_n265_), .A1(new_new_n263_), .B0(new_new_n261_), .B1(new_new_n249_), .Y(new_new_n266_));
  NO2        g0244(.A(new_new_n230_), .B(new_new_n36_), .Y(new_new_n267_));
  NA2        g0245(.A(i_12_), .B(i_6_), .Y(new_new_n268_));
  OR2        g0246(.A(i_13_), .B(i_9_), .Y(new_new_n269_));
  NO3        g0247(.A(new_new_n269_), .B(new_new_n268_), .C(new_new_n48_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n240_), .B(i_2_), .Y(new_new_n271_));
  NA3        g0249(.A(new_new_n271_), .B(new_new_n270_), .C(new_new_n44_), .Y(new_new_n272_));
  NA2        g0250(.A(new_new_n249_), .B(i_9_), .Y(new_new_n273_));
  OAI210     g0251(.A0(new_new_n69_), .A1(new_new_n273_), .B0(new_new_n272_), .Y(new_new_n274_));
  NO3        g0252(.A(i_11_), .B(new_new_n222_), .C(new_new_n25_), .Y(new_new_n275_));
  NO2        g0253(.A(new_new_n251_), .B(i_8_), .Y(new_new_n276_));
  NO2        g0254(.A(i_6_), .B(new_new_n48_), .Y(new_new_n277_));
  NA3        g0255(.A(new_new_n277_), .B(new_new_n276_), .C(new_new_n275_), .Y(new_new_n278_));
  NO3        g0256(.A(new_new_n26_), .B(new_new_n81_), .C(i_5_), .Y(new_new_n279_));
  NA3        g0257(.A(new_new_n279_), .B(new_new_n267_), .C(new_new_n223_), .Y(new_new_n280_));
  AOI210     g0258(.A0(new_new_n280_), .A1(new_new_n278_), .B0(new_new_n69_), .Y(new_new_n281_));
  AOI210     g0259(.A0(new_new_n274_), .A1(new_new_n267_), .B0(new_new_n281_), .Y(new_new_n282_));
  NA4        g0260(.A(new_new_n282_), .B(new_new_n266_), .C(new_new_n248_), .D(new_new_n226_), .Y(new_new_n283_));
  NO3        g0261(.A(i_12_), .B(new_new_n222_), .C(new_new_n36_), .Y(new_new_n284_));
  INV        g0262(.A(new_new_n284_), .Y(new_new_n285_));
  NOi21      g0263(.An(new_new_n156_), .B(new_new_n81_), .Y(new_new_n286_));
  NO3        g0264(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n287_));
  AOI220     g0265(.A0(new_new_n287_), .A1(new_new_n191_), .B0(new_new_n286_), .B1(new_new_n232_), .Y(new_new_n288_));
  NO2        g0266(.A(new_new_n288_), .B(i_7_), .Y(new_new_n289_));
  NO3        g0267(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n237_), .B(i_0_), .Y(new_new_n291_));
  AOI220     g0269(.A0(new_new_n291_), .A1(new_new_n189_), .B0(new_new_n290_), .B1(new_new_n134_), .Y(new_new_n292_));
  NA2        g0270(.A(new_new_n277_), .B(new_new_n26_), .Y(new_new_n293_));
  NO2        g0271(.A(new_new_n293_), .B(new_new_n292_), .Y(new_new_n294_));
  NA2        g0272(.A(i_0_), .B(i_1_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n295_), .B(i_2_), .Y(new_new_n296_));
  NO2        g0274(.A(new_new_n57_), .B(i_6_), .Y(new_new_n297_));
  NA3        g0275(.A(new_new_n297_), .B(new_new_n296_), .C(new_new_n156_), .Y(new_new_n298_));
  OAI210     g0276(.A0(new_new_n158_), .A1(new_new_n135_), .B0(new_new_n298_), .Y(new_new_n299_));
  NO3        g0277(.A(new_new_n299_), .B(new_new_n294_), .C(new_new_n289_), .Y(new_new_n300_));
  NO2        g0278(.A(i_3_), .B(i_10_), .Y(new_new_n301_));
  NA3        g0279(.A(new_new_n301_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n302_));
  NO2        g0280(.A(i_2_), .B(new_new_n95_), .Y(new_new_n303_));
  NO2        g0281(.A(i_4_), .B(i_8_), .Y(new_new_n304_));
  NOi21      g0282(.An(new_new_n214_), .B(new_new_n97_), .Y(new_new_n305_));
  NA3        g0283(.A(new_new_n305_), .B(new_new_n304_), .C(new_new_n303_), .Y(new_new_n306_));
  AN2        g0284(.A(i_3_), .B(i_10_), .Y(new_new_n307_));
  NA4        g0285(.A(new_new_n307_), .B(new_new_n193_), .C(new_new_n170_), .D(new_new_n168_), .Y(new_new_n308_));
  NO2        g0286(.A(i_5_), .B(new_new_n36_), .Y(new_new_n309_));
  NO2        g0287(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n310_));
  OR2        g0288(.A(new_new_n306_), .B(new_new_n302_), .Y(new_new_n311_));
  OAI220     g0289(.A0(new_new_n311_), .A1(i_6_), .B0(new_new_n300_), .B1(new_new_n285_), .Y(new_new_n312_));
  NO4        g0290(.A(new_new_n312_), .B(new_new_n283_), .C(new_new_n210_), .D(new_new_n161_), .Y(new_new_n313_));
  NO3        g0291(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n314_));
  NO2        g0292(.A(new_new_n57_), .B(new_new_n81_), .Y(new_new_n315_));
  NA2        g0293(.A(new_new_n291_), .B(new_new_n315_), .Y(new_new_n316_));
  NO3        g0294(.A(i_6_), .B(new_new_n188_), .C(i_7_), .Y(new_new_n317_));
  AOI210     g0295(.A0(new_new_n1084_), .A1(new_new_n316_), .B0(new_new_n163_), .Y(new_new_n318_));
  NO2        g0296(.A(i_2_), .B(i_3_), .Y(new_new_n319_));
  OR2        g0297(.A(i_0_), .B(i_5_), .Y(new_new_n320_));
  NA2        g0298(.A(new_new_n214_), .B(new_new_n320_), .Y(new_new_n321_));
  NA4        g0299(.A(new_new_n321_), .B(new_new_n231_), .C(new_new_n319_), .D(i_1_), .Y(new_new_n322_));
  NA3        g0300(.A(new_new_n291_), .B(new_new_n286_), .C(new_new_n107_), .Y(new_new_n323_));
  NAi21      g0301(.An(i_8_), .B(i_7_), .Y(new_new_n324_));
  NO2        g0302(.A(new_new_n324_), .B(i_6_), .Y(new_new_n325_));
  NO2        g0303(.A(new_new_n150_), .B(new_new_n46_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n326_), .B(new_new_n325_), .C(new_new_n156_), .Y(new_new_n327_));
  NA3        g0305(.A(new_new_n327_), .B(new_new_n323_), .C(new_new_n322_), .Y(new_new_n328_));
  OAI210     g0306(.A0(new_new_n328_), .A1(new_new_n318_), .B0(i_4_), .Y(new_new_n329_));
  NO2        g0307(.A(i_12_), .B(i_10_), .Y(new_new_n330_));
  NOi21      g0308(.An(i_5_), .B(i_0_), .Y(new_new_n331_));
  AOI210     g0309(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n95_), .Y(new_new_n332_));
  NO4        g0310(.A(new_new_n332_), .B(i_4_), .C(new_new_n331_), .D(new_new_n122_), .Y(new_new_n333_));
  NA4        g0311(.A(new_new_n79_), .B(new_new_n35_), .C(new_new_n81_), .D(i_8_), .Y(new_new_n334_));
  NA2        g0312(.A(new_new_n333_), .B(new_new_n330_), .Y(new_new_n335_));
  NO2        g0313(.A(i_6_), .B(i_8_), .Y(new_new_n336_));
  NOi21      g0314(.An(i_0_), .B(i_2_), .Y(new_new_n337_));
  AN2        g0315(.A(new_new_n337_), .B(new_new_n336_), .Y(new_new_n338_));
  NO2        g0316(.A(i_1_), .B(i_7_), .Y(new_new_n339_));
  AO220      g0317(.A0(new_new_n339_), .A1(new_new_n338_), .B0(new_new_n325_), .B1(new_new_n232_), .Y(new_new_n340_));
  NA2        g0318(.A(new_new_n340_), .B(new_new_n41_), .Y(new_new_n341_));
  NA3        g0319(.A(new_new_n341_), .B(new_new_n335_), .C(new_new_n329_), .Y(new_new_n342_));
  NO3        g0320(.A(new_new_n230_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n343_));
  NO3        g0321(.A(new_new_n324_), .B(i_2_), .C(i_1_), .Y(new_new_n344_));
  OAI210     g0322(.A0(new_new_n344_), .A1(new_new_n343_), .B0(i_6_), .Y(new_new_n345_));
  NA3        g0323(.A(new_new_n250_), .B(new_new_n303_), .C(new_new_n188_), .Y(new_new_n346_));
  NA2        g0324(.A(new_new_n346_), .B(new_new_n345_), .Y(new_new_n347_));
  NOi21      g0325(.An(new_new_n146_), .B(new_new_n98_), .Y(new_new_n348_));
  NO2        g0326(.A(new_new_n348_), .B(new_new_n119_), .Y(new_new_n349_));
  OAI210     g0327(.A0(new_new_n349_), .A1(new_new_n347_), .B0(i_3_), .Y(new_new_n350_));
  INV        g0328(.A(new_new_n79_), .Y(new_new_n351_));
  NO2        g0329(.A(new_new_n295_), .B(new_new_n76_), .Y(new_new_n352_));
  NA2        g0330(.A(new_new_n352_), .B(new_new_n126_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n88_), .B(new_new_n188_), .Y(new_new_n354_));
  NA3        g0332(.A(new_new_n305_), .B(new_new_n354_), .C(new_new_n61_), .Y(new_new_n355_));
  AOI210     g0333(.A0(new_new_n355_), .A1(new_new_n353_), .B0(new_new_n351_), .Y(new_new_n356_));
  NO2        g0334(.A(new_new_n188_), .B(i_9_), .Y(new_new_n357_));
  NA2        g0335(.A(new_new_n357_), .B(new_new_n201_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n358_), .B(new_new_n46_), .Y(new_new_n359_));
  NO3        g0337(.A(new_new_n359_), .B(new_new_n356_), .C(new_new_n294_), .Y(new_new_n360_));
  AOI210     g0338(.A0(new_new_n360_), .A1(new_new_n350_), .B0(new_new_n155_), .Y(new_new_n361_));
  AOI210     g0339(.A0(new_new_n342_), .A1(new_new_n314_), .B0(new_new_n361_), .Y(new_new_n362_));
  NOi32      g0340(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n363_));
  INV        g0341(.A(new_new_n363_), .Y(new_new_n364_));
  NAi21      g0342(.An(i_0_), .B(i_6_), .Y(new_new_n365_));
  NAi21      g0343(.An(i_1_), .B(i_5_), .Y(new_new_n366_));
  NA2        g0344(.A(new_new_n366_), .B(new_new_n365_), .Y(new_new_n367_));
  NA2        g0345(.A(new_new_n367_), .B(new_new_n25_), .Y(new_new_n368_));
  OAI210     g0346(.A0(new_new_n368_), .A1(new_new_n152_), .B0(new_new_n244_), .Y(new_new_n369_));
  NAi41      g0347(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n370_));
  OAI220     g0348(.A0(new_new_n370_), .A1(new_new_n366_), .B0(new_new_n217_), .B1(new_new_n152_), .Y(new_new_n371_));
  AOI210     g0349(.A0(new_new_n370_), .A1(new_new_n152_), .B0(new_new_n150_), .Y(new_new_n372_));
  NOi32      g0350(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n373_));
  NAi21      g0351(.An(i_6_), .B(i_1_), .Y(new_new_n374_));
  NA3        g0352(.A(new_new_n374_), .B(new_new_n373_), .C(new_new_n46_), .Y(new_new_n375_));
  NO2        g0353(.A(new_new_n375_), .B(i_0_), .Y(new_new_n376_));
  OR3        g0354(.A(new_new_n376_), .B(new_new_n372_), .C(new_new_n371_), .Y(new_new_n377_));
  NO2        g0355(.A(i_1_), .B(new_new_n95_), .Y(new_new_n378_));
  NAi21      g0356(.An(i_3_), .B(i_4_), .Y(new_new_n379_));
  NO2        g0357(.A(new_new_n379_), .B(i_9_), .Y(new_new_n380_));
  AN2        g0358(.A(i_6_), .B(i_7_), .Y(new_new_n381_));
  OAI210     g0359(.A0(new_new_n381_), .A1(new_new_n378_), .B0(new_new_n380_), .Y(new_new_n382_));
  NA2        g0360(.A(i_2_), .B(i_7_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n379_), .B(i_10_), .Y(new_new_n384_));
  NA3        g0362(.A(new_new_n384_), .B(new_new_n383_), .C(new_new_n242_), .Y(new_new_n385_));
  AOI210     g0363(.A0(new_new_n385_), .A1(new_new_n382_), .B0(new_new_n180_), .Y(new_new_n386_));
  AOI210     g0364(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n387_));
  OAI210     g0365(.A0(new_new_n387_), .A1(new_new_n183_), .B0(new_new_n384_), .Y(new_new_n388_));
  AOI220     g0366(.A0(new_new_n384_), .A1(new_new_n339_), .B0(new_new_n236_), .B1(new_new_n183_), .Y(new_new_n389_));
  AOI210     g0367(.A0(new_new_n389_), .A1(new_new_n388_), .B0(i_5_), .Y(new_new_n390_));
  NO4        g0368(.A(new_new_n390_), .B(new_new_n386_), .C(new_new_n377_), .D(new_new_n369_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(new_new_n364_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n393_));
  AN2        g0371(.A(i_12_), .B(i_5_), .Y(new_new_n394_));
  NO2        g0372(.A(i_4_), .B(new_new_n26_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n395_), .B(new_new_n394_), .Y(new_new_n396_));
  NO2        g0374(.A(i_11_), .B(i_6_), .Y(new_new_n397_));
  NA3        g0375(.A(new_new_n397_), .B(new_new_n326_), .C(new_new_n222_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n398_), .B(new_new_n396_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n240_), .B(i_5_), .Y(new_new_n400_));
  NO2        g0378(.A(i_5_), .B(i_10_), .Y(new_new_n401_));
  AOI220     g0379(.A0(new_new_n401_), .A1(new_new_n271_), .B0(new_new_n400_), .B1(new_new_n193_), .Y(new_new_n402_));
  NA2        g0380(.A(new_new_n136_), .B(new_new_n45_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(new_new_n402_), .Y(new_new_n404_));
  OAI210     g0382(.A0(new_new_n404_), .A1(new_new_n399_), .B0(new_new_n393_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n36_), .B(new_new_n25_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n142_), .B(new_new_n81_), .Y(new_new_n407_));
  OAI210     g0385(.A0(new_new_n407_), .A1(new_new_n399_), .B0(new_new_n406_), .Y(new_new_n408_));
  NO3        g0386(.A(new_new_n81_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n409_));
  NO2        g0387(.A(i_3_), .B(new_new_n95_), .Y(new_new_n410_));
  NO2        g0388(.A(i_11_), .B(i_12_), .Y(new_new_n411_));
  NA2        g0389(.A(new_new_n401_), .B(new_new_n234_), .Y(new_new_n412_));
  NA3        g0390(.A(new_new_n107_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n413_));
  OAI220     g0391(.A0(new_new_n413_), .A1(new_new_n217_), .B0(new_new_n412_), .B1(new_new_n334_), .Y(new_new_n414_));
  NAi21      g0392(.An(i_13_), .B(i_0_), .Y(new_new_n415_));
  INV        g0393(.A(new_new_n415_), .Y(new_new_n416_));
  NA2        g0394(.A(new_new_n414_), .B(new_new_n416_), .Y(new_new_n417_));
  NA3        g0395(.A(new_new_n417_), .B(new_new_n408_), .C(new_new_n405_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n44_), .B(new_new_n222_), .Y(new_new_n419_));
  NO3        g0397(.A(i_1_), .B(i_12_), .C(new_new_n81_), .Y(new_new_n420_));
  NO2        g0398(.A(i_0_), .B(i_11_), .Y(new_new_n421_));
  NOi21      g0399(.An(i_2_), .B(i_12_), .Y(new_new_n422_));
  NA2        g0400(.A(new_new_n422_), .B(i_6_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n423_), .B(new_new_n1078_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n134_), .B(i_9_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n425_), .B(i_4_), .Y(new_new_n426_));
  NA2        g0404(.A(new_new_n424_), .B(new_new_n426_), .Y(new_new_n427_));
  NAi21      g0405(.An(i_9_), .B(i_4_), .Y(new_new_n428_));
  OR2        g0406(.A(i_13_), .B(i_10_), .Y(new_new_n429_));
  NO3        g0407(.A(new_new_n429_), .B(new_new_n112_), .C(new_new_n428_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n166_), .B(new_new_n118_), .Y(new_new_n431_));
  OR2        g0409(.A(new_new_n212_), .B(new_new_n211_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n95_), .B(new_new_n25_), .Y(new_new_n433_));
  NA2        g0411(.A(new_new_n284_), .B(new_new_n433_), .Y(new_new_n434_));
  NA2        g0412(.A(new_new_n277_), .B(new_new_n206_), .Y(new_new_n435_));
  OAI220     g0413(.A0(new_new_n435_), .A1(new_new_n432_), .B0(new_new_n434_), .B1(new_new_n348_), .Y(new_new_n436_));
  INV        g0414(.A(new_new_n436_), .Y(new_new_n437_));
  AOI210     g0415(.A0(new_new_n437_), .A1(new_new_n427_), .B0(new_new_n26_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n323_), .B(new_new_n322_), .Y(new_new_n439_));
  AOI220     g0417(.A0(new_new_n297_), .A1(new_new_n287_), .B0(new_new_n291_), .B1(new_new_n315_), .Y(new_new_n440_));
  NO2        g0418(.A(new_new_n440_), .B(new_new_n163_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n177_), .B(new_new_n81_), .Y(new_new_n442_));
  AOI220     g0420(.A0(new_new_n442_), .A1(new_new_n296_), .B0(new_new_n279_), .B1(new_new_n206_), .Y(new_new_n443_));
  NO2        g0421(.A(new_new_n443_), .B(i_7_), .Y(new_new_n444_));
  NO3        g0422(.A(new_new_n444_), .B(new_new_n441_), .C(new_new_n439_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n191_), .B(new_new_n90_), .Y(new_new_n446_));
  NA3        g0424(.A(new_new_n326_), .B(new_new_n156_), .C(new_new_n81_), .Y(new_new_n447_));
  AOI210     g0425(.A0(new_new_n447_), .A1(new_new_n446_), .B0(new_new_n324_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n188_), .B(i_10_), .Y(new_new_n449_));
  NA3        g0427(.A(new_new_n256_), .B(new_new_n62_), .C(i_2_), .Y(new_new_n450_));
  NA2        g0428(.A(new_new_n297_), .B(new_new_n232_), .Y(new_new_n451_));
  OAI220     g0429(.A0(new_new_n451_), .A1(new_new_n177_), .B0(new_new_n450_), .B1(new_new_n449_), .Y(new_new_n452_));
  NO2        g0430(.A(i_3_), .B(new_new_n48_), .Y(new_new_n453_));
  NA3        g0431(.A(new_new_n339_), .B(new_new_n338_), .C(new_new_n453_), .Y(new_new_n454_));
  NA2        g0432(.A(new_new_n317_), .B(new_new_n321_), .Y(new_new_n455_));
  OAI210     g0433(.A0(new_new_n455_), .A1(new_new_n184_), .B0(new_new_n454_), .Y(new_new_n456_));
  NO3        g0434(.A(new_new_n456_), .B(new_new_n452_), .C(new_new_n448_), .Y(new_new_n457_));
  AOI210     g0435(.A0(new_new_n457_), .A1(new_new_n445_), .B0(new_new_n273_), .Y(new_new_n458_));
  NO4        g0436(.A(new_new_n458_), .B(new_new_n438_), .C(new_new_n418_), .D(new_new_n392_), .Y(new_new_n459_));
  NO2        g0437(.A(new_new_n61_), .B(i_4_), .Y(new_new_n460_));
  NO2        g0438(.A(new_new_n69_), .B(i_13_), .Y(new_new_n461_));
  NA3        g0439(.A(new_new_n461_), .B(new_new_n460_), .C(i_2_), .Y(new_new_n462_));
  NO2        g0440(.A(i_10_), .B(i_9_), .Y(new_new_n463_));
  NAi21      g0441(.An(i_12_), .B(i_8_), .Y(new_new_n464_));
  NO2        g0442(.A(new_new_n464_), .B(i_3_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n465_), .B(new_new_n463_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n1086_), .B(new_new_n98_), .Y(new_new_n467_));
  OAI220     g0445(.A0(new_new_n467_), .A1(new_new_n200_), .B0(new_new_n466_), .B1(new_new_n462_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n310_), .B(i_0_), .Y(new_new_n469_));
  NO3        g0447(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n470_));
  NA2        g0448(.A(new_new_n268_), .B(new_new_n91_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n471_), .B(new_new_n470_), .Y(new_new_n472_));
  NA2        g0450(.A(i_8_), .B(i_9_), .Y(new_new_n473_));
  AOI210     g0451(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n474_));
  OR2        g0452(.A(new_new_n474_), .B(new_new_n473_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n284_), .B(new_new_n201_), .Y(new_new_n476_));
  OAI220     g0454(.A0(new_new_n476_), .A1(new_new_n475_), .B0(new_new_n472_), .B1(new_new_n469_), .Y(new_new_n477_));
  NA2        g0455(.A(new_new_n249_), .B(new_new_n309_), .Y(new_new_n478_));
  NO3        g0456(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n479_));
  INV        g0457(.A(new_new_n479_), .Y(new_new_n480_));
  NA3        g0458(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n481_));
  NA4        g0459(.A(new_new_n137_), .B(new_new_n110_), .C(new_new_n75_), .D(new_new_n23_), .Y(new_new_n482_));
  OAI220     g0460(.A0(new_new_n482_), .A1(new_new_n481_), .B0(new_new_n480_), .B1(new_new_n478_), .Y(new_new_n483_));
  NO3        g0461(.A(new_new_n483_), .B(new_new_n477_), .C(new_new_n468_), .Y(new_new_n484_));
  NA2        g0462(.A(new_new_n296_), .B(new_new_n102_), .Y(new_new_n485_));
  OR2        g0463(.A(new_new_n485_), .B(new_new_n1081_), .Y(new_new_n486_));
  OA210      g0464(.A0(new_new_n358_), .A1(new_new_n95_), .B0(new_new_n298_), .Y(new_new_n487_));
  OA220      g0465(.A0(new_new_n487_), .A1(new_new_n155_), .B0(new_new_n486_), .B1(new_new_n229_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n90_), .B(i_13_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n442_), .B(new_new_n393_), .Y(new_new_n490_));
  NO2        g0468(.A(i_2_), .B(i_13_), .Y(new_new_n491_));
  NO2        g0469(.A(new_new_n490_), .B(new_new_n489_), .Y(new_new_n492_));
  NO3        g0470(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n493_));
  NO2        g0471(.A(i_6_), .B(i_7_), .Y(new_new_n494_));
  NA2        g0472(.A(new_new_n494_), .B(new_new_n493_), .Y(new_new_n495_));
  OR2        g0473(.A(i_11_), .B(i_8_), .Y(new_new_n496_));
  NOi21      g0474(.An(i_2_), .B(i_7_), .Y(new_new_n497_));
  NAi31      g0475(.An(new_new_n496_), .B(new_new_n497_), .C(new_new_n1080_), .Y(new_new_n498_));
  NO2        g0476(.A(new_new_n429_), .B(i_6_), .Y(new_new_n499_));
  NA3        g0477(.A(new_new_n499_), .B(new_new_n460_), .C(new_new_n71_), .Y(new_new_n500_));
  NO2        g0478(.A(new_new_n500_), .B(new_new_n498_), .Y(new_new_n501_));
  NO2        g0479(.A(i_6_), .B(i_10_), .Y(new_new_n502_));
  NA3        g0480(.A(new_new_n243_), .B(new_new_n165_), .C(new_new_n126_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n504_));
  NO2        g0482(.A(new_new_n150_), .B(i_3_), .Y(new_new_n505_));
  NAi31      g0483(.An(new_new_n504_), .B(new_new_n505_), .C(new_new_n223_), .Y(new_new_n506_));
  NA3        g0484(.A(new_new_n406_), .B(new_new_n173_), .C(new_new_n141_), .Y(new_new_n507_));
  NA3        g0485(.A(new_new_n507_), .B(new_new_n506_), .C(new_new_n503_), .Y(new_new_n508_));
  NO3        g0486(.A(new_new_n508_), .B(new_new_n501_), .C(new_new_n492_), .Y(new_new_n509_));
  NA2        g0487(.A(new_new_n479_), .B(new_new_n401_), .Y(new_new_n510_));
  NO2        g0488(.A(new_new_n510_), .B(new_new_n221_), .Y(new_new_n511_));
  NAi21      g0489(.An(new_new_n212_), .B(new_new_n411_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n339_), .B(new_new_n214_), .Y(new_new_n513_));
  NO2        g0491(.A(new_new_n26_), .B(i_5_), .Y(new_new_n514_));
  NO2        g0492(.A(i_0_), .B(new_new_n81_), .Y(new_new_n515_));
  NA3        g0493(.A(new_new_n515_), .B(new_new_n514_), .C(new_new_n134_), .Y(new_new_n516_));
  OR3        g0494(.A(i_4_), .B(new_new_n37_), .C(new_new_n46_), .Y(new_new_n517_));
  OAI220     g0495(.A0(new_new_n517_), .A1(new_new_n516_), .B0(new_new_n513_), .B1(new_new_n512_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n27_), .B(i_10_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n314_), .B(new_new_n236_), .Y(new_new_n520_));
  OAI220     g0498(.A0(new_new_n520_), .A1(new_new_n450_), .B0(new_new_n519_), .B1(new_new_n489_), .Y(new_new_n521_));
  NA4        g0499(.A(new_new_n307_), .B(new_new_n220_), .C(new_new_n69_), .D(new_new_n234_), .Y(new_new_n522_));
  NO2        g0500(.A(new_new_n522_), .B(new_new_n495_), .Y(new_new_n523_));
  NO4        g0501(.A(new_new_n523_), .B(new_new_n521_), .C(new_new_n518_), .D(new_new_n511_), .Y(new_new_n524_));
  NA4        g0502(.A(new_new_n524_), .B(new_new_n509_), .C(new_new_n488_), .D(new_new_n484_), .Y(new_new_n525_));
  NA3        g0503(.A(new_new_n307_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n526_));
  OAI210     g0504(.A0(new_new_n302_), .A1(new_new_n175_), .B0(new_new_n526_), .Y(new_new_n527_));
  AN2        g0505(.A(new_new_n287_), .B(new_new_n231_), .Y(new_new_n528_));
  NA2        g0506(.A(new_new_n528_), .B(new_new_n527_), .Y(new_new_n529_));
  NA2        g0507(.A(new_new_n117_), .B(new_new_n106_), .Y(new_new_n530_));
  AO220      g0508(.A0(new_new_n530_), .A1(new_new_n470_), .B0(new_new_n430_), .B1(i_6_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n314_), .B(new_new_n157_), .Y(new_new_n532_));
  OAI210     g0510(.A0(new_new_n532_), .A1(new_new_n229_), .B0(new_new_n308_), .Y(new_new_n533_));
  AOI220     g0511(.A0(new_new_n533_), .A1(new_new_n325_), .B0(new_new_n531_), .B1(new_new_n310_), .Y(new_new_n534_));
  NA4        g0512(.A(new_new_n461_), .B(new_new_n460_), .C(new_new_n198_), .D(i_2_), .Y(new_new_n535_));
  INV        g0513(.A(new_new_n535_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n394_), .B(new_new_n222_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n363_), .B(new_new_n69_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n381_), .B(new_new_n373_), .Y(new_new_n539_));
  AO210      g0517(.A0(new_new_n538_), .A1(new_new_n537_), .B0(new_new_n539_), .Y(new_new_n540_));
  NO2        g0518(.A(new_new_n35_), .B(i_8_), .Y(new_new_n541_));
  NAi41      g0519(.An(new_new_n538_), .B(new_new_n502_), .C(new_new_n541_), .D(new_new_n46_), .Y(new_new_n542_));
  AOI210     g0520(.A0(new_new_n38_), .A1(i_13_), .B0(new_new_n430_), .Y(new_new_n543_));
  NA3        g0521(.A(new_new_n543_), .B(new_new_n542_), .C(new_new_n540_), .Y(new_new_n544_));
  AOI210     g0522(.A0(new_new_n536_), .A1(new_new_n199_), .B0(new_new_n544_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n256_), .B(new_new_n62_), .Y(new_new_n546_));
  OAI210     g0524(.A0(i_8_), .A1(new_new_n546_), .B0(new_new_n128_), .Y(new_new_n547_));
  AOI210     g0525(.A0(new_new_n189_), .A1(i_9_), .B0(new_new_n267_), .Y(new_new_n548_));
  NO2        g0526(.A(new_new_n548_), .B(new_new_n194_), .Y(new_new_n549_));
  OR2        g0527(.A(new_new_n177_), .B(i_4_), .Y(new_new_n550_));
  NO2        g0528(.A(new_new_n550_), .B(new_new_n81_), .Y(new_new_n551_));
  AOI220     g0529(.A0(new_new_n551_), .A1(new_new_n549_), .B0(new_new_n547_), .B1(new_new_n431_), .Y(new_new_n552_));
  NA4        g0530(.A(new_new_n552_), .B(new_new_n545_), .C(new_new_n534_), .D(new_new_n529_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n400_), .B(new_new_n296_), .Y(new_new_n554_));
  OAI210     g0532(.A0(new_new_n396_), .A1(new_new_n162_), .B0(new_new_n554_), .Y(new_new_n555_));
  NO2        g0533(.A(i_12_), .B(new_new_n188_), .Y(new_new_n556_));
  NA2        g0534(.A(new_new_n556_), .B(new_new_n222_), .Y(new_new_n557_));
  NA3        g0535(.A(new_new_n502_), .B(new_new_n168_), .C(new_new_n27_), .Y(new_new_n558_));
  NO3        g0536(.A(new_new_n558_), .B(new_new_n557_), .C(new_new_n485_), .Y(new_new_n559_));
  NOi31      g0537(.An(new_new_n317_), .B(new_new_n429_), .C(new_new_n37_), .Y(new_new_n560_));
  OAI210     g0538(.A0(new_new_n560_), .A1(new_new_n559_), .B0(new_new_n555_), .Y(new_new_n561_));
  NO2        g0539(.A(i_8_), .B(i_7_), .Y(new_new_n562_));
  OAI210     g0540(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n563_), .B(new_new_n220_), .Y(new_new_n564_));
  AOI220     g0542(.A0(new_new_n326_), .A1(new_new_n39_), .B0(new_new_n232_), .B1(new_new_n202_), .Y(new_new_n565_));
  OAI220     g0543(.A0(new_new_n565_), .A1(new_new_n550_), .B0(new_new_n564_), .B1(new_new_n240_), .Y(new_new_n566_));
  NA2        g0544(.A(new_new_n44_), .B(i_10_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n567_), .B(i_6_), .Y(new_new_n568_));
  NA3        g0546(.A(new_new_n568_), .B(new_new_n566_), .C(new_new_n562_), .Y(new_new_n569_));
  AOI220     g0547(.A0(new_new_n442_), .A1(new_new_n326_), .B0(new_new_n245_), .B1(new_new_n242_), .Y(new_new_n570_));
  OAI220     g0548(.A0(new_new_n570_), .A1(new_new_n264_), .B0(new_new_n489_), .B1(new_new_n127_), .Y(new_new_n571_));
  NA2        g0549(.A(new_new_n571_), .B(new_new_n267_), .Y(new_new_n572_));
  NOi31      g0550(.An(new_new_n291_), .B(new_new_n302_), .C(new_new_n175_), .Y(new_new_n573_));
  NA3        g0551(.A(new_new_n307_), .B(new_new_n168_), .C(new_new_n90_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n218_), .B(new_new_n44_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n150_), .B(i_5_), .Y(new_new_n576_));
  NA3        g0554(.A(new_new_n576_), .B(new_new_n419_), .C(new_new_n319_), .Y(new_new_n577_));
  OAI210     g0555(.A0(new_new_n577_), .A1(new_new_n575_), .B0(new_new_n574_), .Y(new_new_n578_));
  OAI210     g0556(.A0(new_new_n578_), .A1(new_new_n573_), .B0(new_new_n479_), .Y(new_new_n579_));
  NA4        g0557(.A(new_new_n579_), .B(new_new_n572_), .C(new_new_n569_), .D(new_new_n561_), .Y(new_new_n580_));
  NA2        g0558(.A(new_new_n284_), .B(new_new_n79_), .Y(new_new_n581_));
  AOI210     g0559(.A0(i_11_), .A1(new_new_n353_), .B0(new_new_n581_), .Y(new_new_n582_));
  NA2        g0560(.A(new_new_n297_), .B(new_new_n287_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n583_), .B(new_new_n167_), .Y(new_new_n584_));
  NA2        g0562(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n585_));
  NA2        g0563(.A(new_new_n463_), .B(new_new_n218_), .Y(new_new_n586_));
  NO2        g0564(.A(new_new_n585_), .B(new_new_n586_), .Y(new_new_n587_));
  NA2        g0565(.A(i_0_), .B(new_new_n48_), .Y(new_new_n588_));
  NA3        g0566(.A(new_new_n556_), .B(new_new_n275_), .C(new_new_n588_), .Y(new_new_n589_));
  NO2        g0567(.A(new_new_n1085_), .B(new_new_n589_), .Y(new_new_n590_));
  NO4        g0568(.A(new_new_n590_), .B(new_new_n587_), .C(new_new_n584_), .D(new_new_n582_), .Y(new_new_n591_));
  NO4        g0569(.A(new_new_n250_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n592_));
  NO3        g0570(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n230_), .B(new_new_n35_), .Y(new_new_n594_));
  AN2        g0572(.A(new_new_n594_), .B(new_new_n593_), .Y(new_new_n595_));
  AN2        g0573(.A(new_new_n592_), .B(new_new_n363_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n429_), .B(i_1_), .Y(new_new_n597_));
  NOi31      g0575(.An(new_new_n597_), .B(new_new_n471_), .C(new_new_n69_), .Y(new_new_n598_));
  AN3        g0576(.A(new_new_n598_), .B(new_new_n426_), .C(i_2_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n440_), .B(new_new_n171_), .Y(new_new_n600_));
  NO3        g0578(.A(new_new_n600_), .B(new_new_n599_), .C(new_new_n596_), .Y(new_new_n601_));
  NOi21      g0579(.An(i_10_), .B(i_6_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n81_), .B(new_new_n25_), .Y(new_new_n603_));
  AOI220     g0581(.A0(new_new_n284_), .A1(new_new_n603_), .B0(new_new_n275_), .B1(new_new_n602_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n604_), .B(new_new_n469_), .Y(new_new_n605_));
  NA2        g0583(.A(new_new_n317_), .B(new_new_n157_), .Y(new_new_n606_));
  AOI220     g0584(.A0(new_new_n606_), .A1(new_new_n451_), .B0(new_new_n178_), .B1(new_new_n176_), .Y(new_new_n607_));
  NO2        g0585(.A(new_new_n193_), .B(new_new_n36_), .Y(new_new_n608_));
  NOi31      g0586(.An(new_new_n138_), .B(new_new_n608_), .C(new_new_n334_), .Y(new_new_n609_));
  NO3        g0587(.A(new_new_n609_), .B(new_new_n607_), .C(new_new_n605_), .Y(new_new_n610_));
  NO2        g0588(.A(new_new_n538_), .B(new_new_n389_), .Y(new_new_n611_));
  INV        g0589(.A(new_new_n319_), .Y(new_new_n612_));
  NO2        g0590(.A(i_12_), .B(new_new_n81_), .Y(new_new_n613_));
  NA3        g0591(.A(new_new_n613_), .B(new_new_n275_), .C(new_new_n588_), .Y(new_new_n614_));
  NA3        g0592(.A(new_new_n397_), .B(new_new_n284_), .C(new_new_n214_), .Y(new_new_n615_));
  AOI210     g0593(.A0(new_new_n615_), .A1(new_new_n614_), .B0(new_new_n612_), .Y(new_new_n616_));
  NA2        g0594(.A(new_new_n168_), .B(i_0_), .Y(new_new_n617_));
  NO3        g0595(.A(new_new_n617_), .B(new_new_n345_), .C(new_new_n302_), .Y(new_new_n618_));
  OR2        g0596(.A(i_2_), .B(i_5_), .Y(new_new_n619_));
  BUFFER     g0597(.A(new_new_n619_), .Y(new_new_n620_));
  AOI210     g0598(.A0(new_new_n383_), .A1(new_new_n242_), .B0(new_new_n193_), .Y(new_new_n621_));
  AOI210     g0599(.A0(new_new_n621_), .A1(new_new_n620_), .B0(new_new_n512_), .Y(new_new_n622_));
  NO4        g0600(.A(new_new_n622_), .B(new_new_n618_), .C(new_new_n616_), .D(new_new_n611_), .Y(new_new_n623_));
  NA4        g0601(.A(new_new_n623_), .B(new_new_n610_), .C(new_new_n601_), .D(new_new_n591_), .Y(new_new_n624_));
  NO4        g0602(.A(new_new_n624_), .B(new_new_n580_), .C(new_new_n553_), .D(new_new_n525_), .Y(new_new_n625_));
  NA4        g0603(.A(new_new_n625_), .B(new_new_n459_), .C(new_new_n362_), .D(new_new_n313_), .Y(men7));
  NO2        g0604(.A(new_new_n88_), .B(new_new_n52_), .Y(new_new_n627_));
  NO2        g0605(.A(new_new_n102_), .B(new_new_n86_), .Y(new_new_n628_));
  NA2        g0606(.A(new_new_n395_), .B(new_new_n628_), .Y(new_new_n629_));
  NA2        g0607(.A(new_new_n502_), .B(new_new_n79_), .Y(new_new_n630_));
  OAI210     g0608(.A0(new_new_n1082_), .A1(new_new_n630_), .B0(new_new_n629_), .Y(new_new_n631_));
  NA3        g0609(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n632_));
  NA2        g0610(.A(i_12_), .B(i_8_), .Y(new_new_n633_));
  AOI210     g0611(.A0(new_new_n633_), .A1(new_new_n99_), .B0(new_new_n632_), .Y(new_new_n634_));
  NA2        g0612(.A(i_2_), .B(new_new_n81_), .Y(new_new_n635_));
  OAI210     g0613(.A0(new_new_n84_), .A1(new_new_n198_), .B0(new_new_n199_), .Y(new_new_n636_));
  NO2        g0614(.A(i_7_), .B(new_new_n36_), .Y(new_new_n637_));
  NA2        g0615(.A(i_4_), .B(i_8_), .Y(new_new_n638_));
  NO2        g0616(.A(new_new_n307_), .B(new_new_n637_), .Y(new_new_n639_));
  OAI220     g0617(.A0(new_new_n639_), .A1(new_new_n635_), .B0(new_new_n636_), .B1(i_13_), .Y(new_new_n640_));
  NO4        g0618(.A(new_new_n640_), .B(new_new_n634_), .C(new_new_n631_), .D(new_new_n627_), .Y(new_new_n641_));
  AOI210     g0619(.A0(new_new_n122_), .A1(new_new_n60_), .B0(i_10_), .Y(new_new_n642_));
  AOI210     g0620(.A0(new_new_n642_), .A1(new_new_n234_), .B0(new_new_n154_), .Y(new_new_n643_));
  OR2        g0621(.A(i_6_), .B(i_10_), .Y(new_new_n644_));
  NO2        g0622(.A(new_new_n644_), .B(new_new_n23_), .Y(new_new_n645_));
  OR3        g0623(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n646_));
  NO2        g0624(.A(new_new_n646_), .B(i_8_), .Y(new_new_n647_));
  INV        g0625(.A(new_new_n195_), .Y(new_new_n648_));
  OA220      g0626(.A0(new_new_n646_), .A1(new_new_n612_), .B0(new_new_n643_), .B1(new_new_n269_), .Y(new_new_n649_));
  AOI210     g0627(.A0(new_new_n649_), .A1(new_new_n641_), .B0(new_new_n61_), .Y(new_new_n650_));
  NOi21      g0628(.An(i_11_), .B(i_7_), .Y(new_new_n651_));
  AO210      g0629(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n652_), .B(new_new_n651_), .Y(new_new_n653_));
  NA3        g0631(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n654_));
  NAi21      g0632(.An(new_new_n654_), .B(i_11_), .Y(new_new_n655_));
  NO2        g0633(.A(new_new_n655_), .B(new_new_n61_), .Y(new_new_n656_));
  NA2        g0634(.A(new_new_n83_), .B(new_new_n61_), .Y(new_new_n657_));
  AO210      g0635(.A0(new_new_n657_), .A1(new_new_n389_), .B0(new_new_n40_), .Y(new_new_n658_));
  NO3        g0636(.A(new_new_n258_), .B(new_new_n203_), .C(i_8_), .Y(new_new_n659_));
  OAI210     g0637(.A0(new_new_n659_), .A1(new_new_n223_), .B0(new_new_n61_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n422_), .B(new_new_n30_), .Y(new_new_n661_));
  OR2        g0639(.A(new_new_n203_), .B(new_new_n102_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(new_new_n661_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n61_), .B(i_9_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n664_), .B(i_4_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n665_), .B(new_new_n663_), .Y(new_new_n666_));
  NO2        g0644(.A(i_1_), .B(i_12_), .Y(new_new_n667_));
  NA2        g0645(.A(new_new_n667_), .B(new_new_n104_), .Y(new_new_n668_));
  NA4        g0646(.A(new_new_n668_), .B(new_new_n666_), .C(new_new_n660_), .D(new_new_n658_), .Y(new_new_n669_));
  OAI210     g0647(.A0(new_new_n669_), .A1(new_new_n656_), .B0(i_6_), .Y(new_new_n670_));
  OAI210     g0648(.A0(new_new_n654_), .A1(new_new_n102_), .B0(new_new_n481_), .Y(new_new_n671_));
  NA2        g0649(.A(new_new_n671_), .B(new_new_n613_), .Y(new_new_n672_));
  NO2        g0650(.A(i_6_), .B(i_11_), .Y(new_new_n673_));
  NA2        g0651(.A(new_new_n672_), .B(new_new_n472_), .Y(new_new_n674_));
  NO4        g0652(.A(new_new_n211_), .B(new_new_n122_), .C(i_13_), .D(new_new_n81_), .Y(new_new_n675_));
  INV        g0653(.A(new_new_n675_), .Y(new_new_n676_));
  NA2        g0654(.A(new_new_n234_), .B(i_6_), .Y(new_new_n677_));
  NO3        g0655(.A(new_new_n644_), .B(new_new_n230_), .C(new_new_n23_), .Y(new_new_n678_));
  AOI210     g0656(.A0(i_1_), .A1(new_new_n259_), .B0(new_new_n678_), .Y(new_new_n679_));
  OAI210     g0657(.A0(new_new_n679_), .A1(new_new_n44_), .B0(new_new_n676_), .Y(new_new_n680_));
  NA3        g0658(.A(new_new_n562_), .B(i_11_), .C(new_new_n35_), .Y(new_new_n681_));
  NA3        g0659(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n46_), .B(i_1_), .Y(new_new_n683_));
  NA3        g0661(.A(new_new_n683_), .B(new_new_n268_), .C(new_new_n44_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n684_), .B(new_new_n682_), .Y(new_new_n685_));
  NA3        g0663(.A(new_new_n664_), .B(new_new_n319_), .C(i_6_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n686_), .B(new_new_n23_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n683_), .B(new_new_n268_), .Y(new_new_n688_));
  NO2        g0666(.A(i_11_), .B(new_new_n36_), .Y(new_new_n689_));
  NA2        g0667(.A(new_new_n689_), .B(new_new_n24_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n690_), .B(new_new_n688_), .Y(new_new_n691_));
  OR3        g0669(.A(new_new_n691_), .B(new_new_n687_), .C(new_new_n685_), .Y(new_new_n692_));
  NO3        g0670(.A(new_new_n692_), .B(new_new_n680_), .C(new_new_n674_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n234_), .B(new_new_n95_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n694_), .B(new_new_n651_), .Y(new_new_n695_));
  NA2        g0673(.A(new_new_n695_), .B(i_1_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n696_), .B(new_new_n646_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n428_), .B(new_new_n81_), .Y(new_new_n698_));
  NA2        g0676(.A(new_new_n697_), .B(new_new_n46_), .Y(new_new_n699_));
  NA2        g0677(.A(i_3_), .B(new_new_n188_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n230_), .B(new_new_n44_), .Y(new_new_n701_));
  NO3        g0679(.A(new_new_n701_), .B(new_new_n310_), .C(new_new_n235_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n112_), .B(new_new_n36_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n81_), .B(i_9_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n704_), .B(new_new_n61_), .Y(new_new_n705_));
  NO2        g0683(.A(new_new_n705_), .B(new_new_n667_), .Y(new_new_n706_));
  NO4        g0684(.A(new_new_n706_), .B(new_new_n1088_), .C(new_new_n702_), .D(i_4_), .Y(new_new_n707_));
  NA2        g0685(.A(i_1_), .B(i_3_), .Y(new_new_n708_));
  NO2        g0686(.A(new_new_n473_), .B(new_new_n88_), .Y(new_new_n709_));
  AOI210     g0687(.A0(new_new_n701_), .A1(new_new_n602_), .B0(new_new_n709_), .Y(new_new_n710_));
  NO2        g0688(.A(new_new_n710_), .B(new_new_n708_), .Y(new_new_n711_));
  NO2        g0689(.A(new_new_n711_), .B(new_new_n707_), .Y(new_new_n712_));
  NA4        g0690(.A(new_new_n712_), .B(new_new_n699_), .C(new_new_n693_), .D(new_new_n670_), .Y(new_new_n713_));
  NO3        g0691(.A(new_new_n496_), .B(i_3_), .C(i_7_), .Y(new_new_n714_));
  NOi21      g0692(.An(new_new_n714_), .B(i_10_), .Y(new_new_n715_));
  OA210      g0693(.A0(new_new_n715_), .A1(new_new_n243_), .B0(new_new_n81_), .Y(new_new_n716_));
  NA2        g0694(.A(new_new_n381_), .B(new_new_n380_), .Y(new_new_n717_));
  NA3        g0695(.A(new_new_n502_), .B(new_new_n541_), .C(new_new_n46_), .Y(new_new_n718_));
  NO3        g0696(.A(new_new_n497_), .B(new_new_n638_), .C(new_new_n81_), .Y(new_new_n719_));
  NA2        g0697(.A(new_new_n719_), .B(new_new_n25_), .Y(new_new_n720_));
  NA3        g0698(.A(new_new_n154_), .B(new_new_n79_), .C(new_new_n81_), .Y(new_new_n721_));
  NA4        g0699(.A(new_new_n721_), .B(new_new_n720_), .C(new_new_n718_), .D(new_new_n717_), .Y(new_new_n722_));
  OAI210     g0700(.A0(new_new_n722_), .A1(new_new_n716_), .B0(i_1_), .Y(new_new_n723_));
  NO2        g0701(.A(new_new_n686_), .B(new_new_n464_), .Y(new_new_n724_));
  INV        g0702(.A(new_new_n724_), .Y(new_new_n725_));
  AOI210     g0703(.A0(new_new_n725_), .A1(new_new_n723_), .B0(i_13_), .Y(new_new_n726_));
  OR2        g0704(.A(i_11_), .B(i_7_), .Y(new_new_n727_));
  NA3        g0705(.A(new_new_n727_), .B(new_new_n100_), .C(new_new_n132_), .Y(new_new_n728_));
  AOI220     g0706(.A0(new_new_n491_), .A1(new_new_n154_), .B0(new_new_n1086_), .B1(new_new_n132_), .Y(new_new_n729_));
  OAI210     g0707(.A0(new_new_n729_), .A1(new_new_n44_), .B0(new_new_n728_), .Y(new_new_n730_));
  NO2        g0708(.A(new_new_n497_), .B(new_new_n24_), .Y(new_new_n731_));
  AOI220     g0709(.A0(new_new_n731_), .A1(new_new_n698_), .B0(new_new_n243_), .B1(new_new_n125_), .Y(new_new_n732_));
  NO2        g0710(.A(new_new_n732_), .B(new_new_n40_), .Y(new_new_n733_));
  AOI210     g0711(.A0(new_new_n730_), .A1(new_new_n336_), .B0(new_new_n733_), .Y(new_new_n734_));
  NA2        g0712(.A(i_7_), .B(new_new_n68_), .Y(new_new_n735_));
  NO2        g0713(.A(new_new_n735_), .B(new_new_n240_), .Y(new_new_n736_));
  AOI210     g0714(.A0(new_new_n464_), .A1(new_new_n35_), .B0(i_13_), .Y(new_new_n737_));
  NOi31      g0715(.An(new_new_n737_), .B(new_new_n630_), .C(new_new_n44_), .Y(new_new_n738_));
  NO2        g0716(.A(new_new_n682_), .B(new_new_n109_), .Y(new_new_n739_));
  INV        g0717(.A(new_new_n739_), .Y(new_new_n740_));
  NO2        g0718(.A(new_new_n740_), .B(new_new_n67_), .Y(new_new_n741_));
  NO3        g0719(.A(new_new_n67_), .B(new_new_n31_), .C(new_new_n95_), .Y(new_new_n742_));
  NA2        g0720(.A(new_new_n26_), .B(new_new_n188_), .Y(new_new_n743_));
  NA2        g0721(.A(new_new_n743_), .B(i_7_), .Y(new_new_n744_));
  NO3        g0722(.A(new_new_n497_), .B(new_new_n234_), .C(new_new_n81_), .Y(new_new_n745_));
  AOI210     g0723(.A0(new_new_n745_), .A1(new_new_n744_), .B0(new_new_n742_), .Y(new_new_n746_));
  NA2        g0724(.A(new_new_n397_), .B(new_new_n683_), .Y(new_new_n747_));
  OAI220     g0725(.A0(new_new_n747_), .A1(new_new_n633_), .B0(new_new_n746_), .B1(new_new_n648_), .Y(new_new_n748_));
  NO4        g0726(.A(new_new_n748_), .B(new_new_n741_), .C(new_new_n738_), .D(new_new_n736_), .Y(new_new_n749_));
  OR2        g0727(.A(i_11_), .B(i_6_), .Y(new_new_n750_));
  NA3        g0728(.A(i_12_), .B(new_new_n743_), .C(i_7_), .Y(new_new_n751_));
  NO2        g0729(.A(new_new_n751_), .B(new_new_n750_), .Y(new_new_n752_));
  NA2        g0730(.A(new_new_n673_), .B(i_13_), .Y(new_new_n753_));
  NA2        g0731(.A(new_new_n96_), .B(new_new_n743_), .Y(new_new_n754_));
  NAi21      g0732(.An(i_11_), .B(i_12_), .Y(new_new_n755_));
  NOi41      g0733(.An(new_new_n105_), .B(new_new_n755_), .C(i_13_), .D(new_new_n81_), .Y(new_new_n756_));
  NO3        g0734(.A(new_new_n497_), .B(new_new_n613_), .C(new_new_n638_), .Y(new_new_n757_));
  AOI220     g0735(.A0(new_new_n757_), .A1(new_new_n314_), .B0(new_new_n756_), .B1(new_new_n754_), .Y(new_new_n758_));
  NA2        g0736(.A(new_new_n758_), .B(new_new_n753_), .Y(new_new_n759_));
  OAI210     g0737(.A0(new_new_n759_), .A1(new_new_n752_), .B0(new_new_n61_), .Y(new_new_n760_));
  NO2        g0738(.A(i_2_), .B(i_12_), .Y(new_new_n761_));
  NA2        g0739(.A(new_new_n378_), .B(new_new_n761_), .Y(new_new_n762_));
  OAI210     g0740(.A0(i_8_), .A1(new_new_n380_), .B0(new_new_n378_), .Y(new_new_n763_));
  NO2        g0741(.A(new_new_n122_), .B(i_2_), .Y(new_new_n764_));
  NA2        g0742(.A(new_new_n764_), .B(new_new_n667_), .Y(new_new_n765_));
  NA3        g0743(.A(new_new_n765_), .B(new_new_n763_), .C(new_new_n762_), .Y(new_new_n766_));
  NA3        g0744(.A(new_new_n766_), .B(new_new_n45_), .C(new_new_n222_), .Y(new_new_n767_));
  NA4        g0745(.A(new_new_n767_), .B(new_new_n760_), .C(new_new_n749_), .D(new_new_n734_), .Y(new_new_n768_));
  OR4        g0746(.A(new_new_n768_), .B(new_new_n726_), .C(new_new_n713_), .D(new_new_n650_), .Y(men5));
  AOI210     g0747(.A0(new_new_n695_), .A1(new_new_n271_), .B0(new_new_n431_), .Y(new_new_n770_));
  NA3        g0748(.A(new_new_n24_), .B(new_new_n761_), .C(new_new_n102_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n771_), .B(new_new_n770_), .Y(new_new_n772_));
  NO3        g0750(.A(i_11_), .B(new_new_n234_), .C(i_13_), .Y(new_new_n773_));
  NO2        g0751(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n774_));
  NA2        g0752(.A(i_12_), .B(i_8_), .Y(new_new_n775_));
  INV        g0753(.A(new_new_n463_), .Y(new_new_n776_));
  INV        g0754(.A(new_new_n772_), .Y(new_new_n777_));
  INV        g0755(.A(new_new_n165_), .Y(new_new_n778_));
  NO2        g0756(.A(new_new_n473_), .B(new_new_n26_), .Y(new_new_n779_));
  NO2        g0757(.A(new_new_n779_), .B(new_new_n433_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n780_), .B(i_2_), .Y(new_new_n781_));
  INV        g0759(.A(new_new_n781_), .Y(new_new_n782_));
  AOI210     g0760(.A0(new_new_n32_), .A1(new_new_n35_), .B0(new_new_n429_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(new_new_n782_), .Y(new_new_n784_));
  NO2        g0762(.A(new_new_n185_), .B(new_new_n120_), .Y(new_new_n785_));
  OAI210     g0763(.A0(new_new_n785_), .A1(new_new_n774_), .B0(i_2_), .Y(new_new_n786_));
  NO3        g0764(.A(new_new_n652_), .B(new_new_n37_), .C(new_new_n26_), .Y(new_new_n787_));
  AOI210     g0765(.A0(new_new_n165_), .A1(new_new_n84_), .B0(new_new_n787_), .Y(new_new_n788_));
  AOI210     g0766(.A0(new_new_n788_), .A1(new_new_n786_), .B0(new_new_n188_), .Y(new_new_n789_));
  AN2        g0767(.A(new_new_n121_), .B(i_13_), .Y(new_new_n790_));
  NA2        g0768(.A(new_new_n195_), .B(new_new_n198_), .Y(new_new_n791_));
  NA2        g0769(.A(new_new_n144_), .B(i_8_), .Y(new_new_n792_));
  AOI210     g0770(.A0(new_new_n792_), .A1(new_new_n791_), .B0(new_new_n383_), .Y(new_new_n793_));
  NA3        g0771(.A(new_new_n307_), .B(new_new_n119_), .C(new_new_n42_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n794_), .B(new_new_n46_), .Y(new_new_n795_));
  NO4        g0773(.A(new_new_n795_), .B(new_new_n793_), .C(new_new_n790_), .D(new_new_n789_), .Y(new_new_n796_));
  NO2        g0774(.A(new_new_n60_), .B(i_12_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n121_), .Y(new_new_n798_));
  NO2        g0776(.A(new_new_n798_), .B(i_8_), .Y(new_new_n799_));
  AOI220     g0777(.A0(new_new_n799_), .A1(new_new_n35_), .B0(new_new_n276_), .B1(new_new_n46_), .Y(new_new_n800_));
  NA4        g0778(.A(new_new_n800_), .B(new_new_n796_), .C(new_new_n784_), .D(new_new_n777_), .Y(men6));
  NA4        g0779(.A(new_new_n401_), .B(new_new_n1089_), .C(new_new_n67_), .D(new_new_n95_), .Y(new_new_n802_));
  INV        g0780(.A(new_new_n802_), .Y(new_new_n803_));
  NO2        g0781(.A(new_new_n217_), .B(new_new_n504_), .Y(new_new_n804_));
  NO2        g0782(.A(i_11_), .B(i_9_), .Y(new_new_n805_));
  NO2        g0783(.A(new_new_n803_), .B(new_new_n331_), .Y(new_new_n806_));
  OR2        g0784(.A(new_new_n806_), .B(i_12_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n384_), .B(new_new_n339_), .Y(new_new_n808_));
  NA2        g0786(.A(new_new_n715_), .B(new_new_n67_), .Y(new_new_n809_));
  NA3        g0787(.A(new_new_n657_), .B(new_new_n809_), .C(new_new_n808_), .Y(new_new_n810_));
  INV        g0788(.A(new_new_n192_), .Y(new_new_n811_));
  AOI220     g0789(.A0(new_new_n811_), .A1(new_new_n805_), .B0(new_new_n810_), .B1(new_new_n69_), .Y(new_new_n812_));
  INV        g0790(.A(new_new_n330_), .Y(new_new_n813_));
  INV        g0791(.A(new_new_n125_), .Y(new_new_n814_));
  NO2        g0792(.A(new_new_n814_), .B(new_new_n813_), .Y(new_new_n815_));
  NO3        g0793(.A(new_new_n250_), .B(new_new_n126_), .C(i_9_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n816_), .B(new_new_n797_), .Y(new_new_n817_));
  AOI210     g0795(.A0(new_new_n817_), .A1(new_new_n539_), .B0(new_new_n180_), .Y(new_new_n818_));
  NO2        g0796(.A(new_new_n31_), .B(i_11_), .Y(new_new_n819_));
  NA3        g0797(.A(new_new_n819_), .B(new_new_n494_), .C(new_new_n401_), .Y(new_new_n820_));
  NAi32      g0798(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n821_));
  AOI210     g0799(.A0(new_new_n750_), .A1(new_new_n82_), .B0(new_new_n821_), .Y(new_new_n822_));
  OAI210     g0800(.A0(new_new_n714_), .A1(new_new_n594_), .B0(new_new_n593_), .Y(new_new_n823_));
  NAi31      g0801(.An(new_new_n822_), .B(new_new_n823_), .C(new_new_n820_), .Y(new_new_n824_));
  OR3        g0802(.A(new_new_n824_), .B(new_new_n818_), .C(new_new_n815_), .Y(new_new_n825_));
  NO2        g0803(.A(new_new_n727_), .B(i_2_), .Y(new_new_n826_));
  NA2        g0804(.A(new_new_n48_), .B(new_new_n36_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n1083_), .B(new_new_n826_), .Y(new_new_n828_));
  AO220      g0806(.A0(new_new_n367_), .A1(new_new_n357_), .B0(new_new_n409_), .B1(i_8_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n829_), .B(new_new_n255_), .Y(new_new_n830_));
  OR2        g0808(.A(new_new_n653_), .B(new_new_n465_), .Y(new_new_n831_));
  NA3        g0809(.A(new_new_n831_), .B(new_new_n139_), .C(new_new_n66_), .Y(new_new_n832_));
  AO210      g0810(.A0(new_new_n510_), .A1(new_new_n776_), .B0(new_new_n35_), .Y(new_new_n833_));
  NA4        g0811(.A(new_new_n833_), .B(new_new_n832_), .C(new_new_n830_), .D(new_new_n828_), .Y(new_new_n834_));
  OAI210     g0812(.A0(i_6_), .A1(i_11_), .B0(new_new_n82_), .Y(new_new_n835_));
  AOI220     g0813(.A0(new_new_n835_), .A1(new_new_n593_), .B0(new_new_n804_), .B1(new_new_n744_), .Y(new_new_n836_));
  NA3        g0814(.A(new_new_n383_), .B(new_new_n236_), .C(new_new_n139_), .Y(new_new_n837_));
  NA3        g0815(.A(new_new_n837_), .B(new_new_n836_), .C(new_new_n636_), .Y(new_new_n838_));
  AO210      g0816(.A0(new_new_n541_), .A1(new_new_n46_), .B0(new_new_n83_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n839_), .B(new_new_n502_), .Y(new_new_n840_));
  INV        g0818(.A(new_new_n592_), .Y(new_new_n841_));
  NO2        g0819(.A(new_new_n644_), .B(new_new_n96_), .Y(new_new_n842_));
  OAI210     g0820(.A0(new_new_n842_), .A1(new_new_n106_), .B0(new_new_n421_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n242_), .B(new_new_n46_), .Y(new_new_n844_));
  INV        g0822(.A(new_new_n620_), .Y(new_new_n845_));
  NA3        g0823(.A(new_new_n845_), .B(new_new_n330_), .C(i_7_), .Y(new_new_n846_));
  NA4        g0824(.A(new_new_n846_), .B(new_new_n843_), .C(new_new_n841_), .D(new_new_n840_), .Y(new_new_n847_));
  NO4        g0825(.A(new_new_n847_), .B(new_new_n838_), .C(new_new_n834_), .D(new_new_n825_), .Y(new_new_n848_));
  NA4        g0826(.A(new_new_n848_), .B(new_new_n812_), .C(new_new_n807_), .D(new_new_n391_), .Y(men3));
  NA2        g0827(.A(i_12_), .B(i_10_), .Y(new_new_n850_));
  NA2        g0828(.A(i_6_), .B(i_7_), .Y(new_new_n851_));
  NO2        g0829(.A(new_new_n851_), .B(i_0_), .Y(new_new_n852_));
  NO2        g0830(.A(i_11_), .B(new_new_n234_), .Y(new_new_n853_));
  OAI210     g0831(.A0(new_new_n852_), .A1(new_new_n291_), .B0(new_new_n853_), .Y(new_new_n854_));
  NO2        g0832(.A(new_new_n854_), .B(new_new_n188_), .Y(new_new_n855_));
  NO3        g0833(.A(new_new_n469_), .B(new_new_n86_), .C(new_new_n44_), .Y(new_new_n856_));
  OA210      g0834(.A0(new_new_n856_), .A1(new_new_n855_), .B0(new_new_n168_), .Y(new_new_n857_));
  NA3        g0835(.A(new_new_n837_), .B(new_new_n636_), .C(new_new_n382_), .Y(new_new_n858_));
  NA2        g0836(.A(new_new_n858_), .B(new_new_n39_), .Y(new_new_n859_));
  NOi21      g0837(.An(new_new_n90_), .B(new_new_n780_), .Y(new_new_n860_));
  NO3        g0838(.A(new_new_n662_), .B(new_new_n473_), .C(new_new_n125_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n422_), .B(new_new_n45_), .Y(new_new_n862_));
  NO3        g0840(.A(new_new_n53_), .B(new_new_n861_), .C(new_new_n860_), .Y(new_new_n863_));
  AOI210     g0841(.A0(new_new_n863_), .A1(new_new_n859_), .B0(new_new_n48_), .Y(new_new_n864_));
  NA2        g0842(.A(new_new_n180_), .B(new_new_n602_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n737_), .B(new_new_n704_), .Y(new_new_n866_));
  NA2        g0844(.A(new_new_n337_), .B(new_new_n453_), .Y(new_new_n867_));
  OAI220     g0845(.A0(new_new_n867_), .A1(new_new_n866_), .B0(new_new_n865_), .B1(new_new_n61_), .Y(new_new_n868_));
  NOi21      g0846(.An(i_5_), .B(i_9_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n869_), .B(new_new_n461_), .Y(new_new_n870_));
  INV        g0848(.A(new_new_n719_), .Y(new_new_n871_));
  NO3        g0849(.A(new_new_n425_), .B(new_new_n268_), .C(new_new_n69_), .Y(new_new_n872_));
  NO2        g0850(.A(new_new_n169_), .B(new_new_n140_), .Y(new_new_n873_));
  AOI210     g0851(.A0(new_new_n873_), .A1(new_new_n242_), .B0(new_new_n872_), .Y(new_new_n874_));
  OAI220     g0852(.A0(new_new_n874_), .A1(new_new_n175_), .B0(new_new_n871_), .B1(new_new_n870_), .Y(new_new_n875_));
  NO4        g0853(.A(new_new_n875_), .B(new_new_n868_), .C(new_new_n864_), .D(new_new_n857_), .Y(new_new_n876_));
  NA2        g0854(.A(new_new_n180_), .B(new_new_n24_), .Y(new_new_n877_));
  NO2        g0855(.A(new_new_n703_), .B(new_new_n628_), .Y(new_new_n878_));
  NO2        g0856(.A(new_new_n878_), .B(new_new_n877_), .Y(new_new_n879_));
  NA2        g0857(.A(new_new_n314_), .B(new_new_n123_), .Y(new_new_n880_));
  NAi21      g0858(.An(new_new_n155_), .B(new_new_n453_), .Y(new_new_n881_));
  OAI220     g0859(.A0(new_new_n881_), .A1(new_new_n844_), .B0(new_new_n880_), .B1(new_new_n412_), .Y(new_new_n882_));
  NO2        g0860(.A(new_new_n882_), .B(new_new_n879_), .Y(new_new_n883_));
  NO2        g0861(.A(new_new_n401_), .B(new_new_n295_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n884_), .B(new_new_n739_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n603_), .B(i_0_), .Y(new_new_n886_));
  NO3        g0864(.A(new_new_n886_), .B(new_new_n396_), .C(new_new_n84_), .Y(new_new_n887_));
  NO3        g0865(.A(new_new_n619_), .B(new_new_n211_), .C(new_new_n429_), .Y(new_new_n888_));
  AOI210     g0866(.A0(new_new_n888_), .A1(i_11_), .B0(new_new_n887_), .Y(new_new_n889_));
  INV        g0867(.A(new_new_n494_), .Y(new_new_n890_));
  AN2        g0868(.A(new_new_n90_), .B(new_new_n241_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n773_), .B(new_new_n331_), .Y(new_new_n892_));
  AOI210     g0870(.A0(new_new_n502_), .A1(new_new_n84_), .B0(new_new_n56_), .Y(new_new_n893_));
  OAI220     g0871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n690_), .B1(new_new_n564_), .Y(new_new_n894_));
  NO2        g0872(.A(new_new_n252_), .B(new_new_n146_), .Y(new_new_n895_));
  NA2        g0873(.A(i_0_), .B(i_10_), .Y(new_new_n896_));
  OAI210     g0874(.A0(new_new_n896_), .A1(new_new_n81_), .B0(new_new_n567_), .Y(new_new_n897_));
  NO4        g0875(.A(new_new_n109_), .B(new_new_n56_), .C(new_new_n700_), .D(i_5_), .Y(new_new_n898_));
  AO220      g0876(.A0(new_new_n898_), .A1(new_new_n897_), .B0(new_new_n895_), .B1(i_6_), .Y(new_new_n899_));
  AOI220     g0877(.A0(new_new_n337_), .A1(new_new_n92_), .B0(new_new_n180_), .B1(new_new_n79_), .Y(new_new_n900_));
  NA2        g0878(.A(new_new_n597_), .B(i_4_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n183_), .B(new_new_n198_), .Y(new_new_n902_));
  OAI220     g0880(.A0(new_new_n902_), .A1(new_new_n892_), .B0(new_new_n901_), .B1(new_new_n900_), .Y(new_new_n903_));
  NO4        g0881(.A(new_new_n903_), .B(new_new_n899_), .C(new_new_n894_), .D(new_new_n891_), .Y(new_new_n904_));
  NA4        g0882(.A(new_new_n904_), .B(new_new_n889_), .C(new_new_n885_), .D(new_new_n883_), .Y(new_new_n905_));
  NO2        g0883(.A(new_new_n97_), .B(new_new_n36_), .Y(new_new_n906_));
  NA2        g0884(.A(i_11_), .B(i_9_), .Y(new_new_n907_));
  NO3        g0885(.A(i_12_), .B(new_new_n907_), .C(new_new_n635_), .Y(new_new_n908_));
  AN2        g0886(.A(new_new_n908_), .B(new_new_n906_), .Y(new_new_n909_));
  NO2        g0887(.A(new_new_n48_), .B(i_7_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n406_), .B(new_new_n173_), .Y(new_new_n911_));
  NAi41      g0889(.An(new_new_n265_), .B(new_new_n911_), .C(new_new_n478_), .D(new_new_n153_), .Y(new_new_n912_));
  NO2        g0890(.A(new_new_n907_), .B(new_new_n69_), .Y(new_new_n913_));
  NO2        g0891(.A(new_new_n169_), .B(i_0_), .Y(new_new_n914_));
  INV        g0892(.A(new_new_n914_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n494_), .B(new_new_n228_), .Y(new_new_n916_));
  AOI210     g0894(.A0(new_new_n381_), .A1(new_new_n41_), .B0(new_new_n420_), .Y(new_new_n917_));
  OAI220     g0895(.A0(new_new_n917_), .A1(new_new_n870_), .B0(new_new_n916_), .B1(new_new_n915_), .Y(new_new_n918_));
  NO3        g0896(.A(new_new_n918_), .B(new_new_n912_), .C(new_new_n909_), .Y(new_new_n919_));
  AOI210     g0897(.A0(new_new_n464_), .A1(new_new_n35_), .B0(i_3_), .Y(new_new_n920_));
  NA2        g0898(.A(new_new_n165_), .B(new_new_n97_), .Y(new_new_n921_));
  NOi32      g0899(.An(new_new_n920_), .Bn(new_new_n183_), .C(new_new_n921_), .Y(new_new_n922_));
  AOI210     g0900(.A0(new_new_n637_), .A1(new_new_n331_), .B0(new_new_n241_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n923_), .B(new_new_n862_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n924_), .B(new_new_n922_), .Y(new_new_n925_));
  NOi21      g0903(.An(i_7_), .B(i_5_), .Y(new_new_n926_));
  NOi31      g0904(.An(new_new_n926_), .B(i_0_), .C(new_new_n755_), .Y(new_new_n927_));
  NA3        g0905(.A(new_new_n927_), .B(new_new_n395_), .C(i_6_), .Y(new_new_n928_));
  OA210      g0906(.A0(new_new_n921_), .A1(new_new_n539_), .B0(new_new_n928_), .Y(new_new_n929_));
  NO3        g0907(.A(new_new_n415_), .B(new_new_n370_), .C(new_new_n366_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n262_), .B(new_new_n320_), .Y(new_new_n931_));
  NO2        g0909(.A(new_new_n755_), .B(new_new_n257_), .Y(new_new_n932_));
  AOI210     g0910(.A0(new_new_n932_), .A1(new_new_n931_), .B0(new_new_n930_), .Y(new_new_n933_));
  NA4        g0911(.A(new_new_n933_), .B(new_new_n929_), .C(new_new_n925_), .D(new_new_n919_), .Y(new_new_n934_));
  NO2        g0912(.A(new_new_n877_), .B(new_new_n237_), .Y(new_new_n935_));
  AN2        g0913(.A(new_new_n336_), .B(new_new_n331_), .Y(new_new_n936_));
  AN2        g0914(.A(new_new_n936_), .B(new_new_n873_), .Y(new_new_n937_));
  OAI210     g0915(.A0(new_new_n937_), .A1(new_new_n935_), .B0(i_10_), .Y(new_new_n938_));
  NO2        g0916(.A(new_new_n850_), .B(new_new_n319_), .Y(new_new_n939_));
  OA210      g0917(.A0(new_new_n494_), .A1(new_new_n220_), .B0(new_new_n493_), .Y(new_new_n940_));
  NA2        g0918(.A(new_new_n939_), .B(new_new_n913_), .Y(new_new_n941_));
  NA3        g0919(.A(new_new_n493_), .B(new_new_n422_), .C(new_new_n45_), .Y(new_new_n942_));
  OAI210     g0920(.A0(new_new_n881_), .A1(new_new_n890_), .B0(new_new_n942_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n255_), .B(new_new_n46_), .Y(new_new_n944_));
  NA2        g0922(.A(new_new_n913_), .B(new_new_n307_), .Y(new_new_n945_));
  OAI210     g0923(.A0(new_new_n944_), .A1(new_new_n182_), .B0(new_new_n945_), .Y(new_new_n946_));
  AOI220     g0924(.A0(new_new_n946_), .A1(new_new_n494_), .B0(new_new_n943_), .B1(new_new_n69_), .Y(new_new_n947_));
  NA3        g0925(.A(new_new_n827_), .B(new_new_n393_), .C(i_6_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n88_), .B(new_new_n44_), .Y(new_new_n949_));
  NO2        g0927(.A(new_new_n71_), .B(new_new_n775_), .Y(new_new_n950_));
  AOI220     g0928(.A0(new_new_n950_), .A1(new_new_n949_), .B0(new_new_n168_), .B1(new_new_n628_), .Y(new_new_n951_));
  AOI210     g0929(.A0(new_new_n951_), .A1(new_new_n948_), .B0(new_new_n47_), .Y(new_new_n952_));
  NO3        g0930(.A(new_new_n619_), .B(new_new_n365_), .C(new_new_n24_), .Y(new_new_n953_));
  AOI210     g0931(.A0(new_new_n731_), .A1(new_new_n576_), .B0(new_new_n953_), .Y(new_new_n954_));
  NAi21      g0932(.An(i_9_), .B(i_5_), .Y(new_new_n955_));
  NO2        g0933(.A(new_new_n955_), .B(new_new_n415_), .Y(new_new_n956_));
  NO2        g0934(.A(new_new_n632_), .B(new_new_n99_), .Y(new_new_n957_));
  AOI220     g0935(.A0(new_new_n957_), .A1(i_0_), .B0(new_new_n956_), .B1(new_new_n653_), .Y(new_new_n958_));
  OAI220     g0936(.A0(new_new_n958_), .A1(new_new_n81_), .B0(new_new_n954_), .B1(new_new_n166_), .Y(new_new_n959_));
  NO3        g0937(.A(new_new_n959_), .B(new_new_n952_), .C(new_new_n544_), .Y(new_new_n960_));
  NA4        g0938(.A(new_new_n960_), .B(new_new_n947_), .C(new_new_n941_), .D(new_new_n938_), .Y(new_new_n961_));
  NO3        g0939(.A(new_new_n961_), .B(new_new_n934_), .C(new_new_n905_), .Y(new_new_n962_));
  NO2        g0940(.A(i_0_), .B(new_new_n755_), .Y(new_new_n963_));
  NA2        g0941(.A(new_new_n69_), .B(new_new_n44_), .Y(new_new_n964_));
  NO3        g0942(.A(new_new_n99_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n965_));
  AO220      g0943(.A0(new_new_n965_), .A1(new_new_n69_), .B0(new_new_n963_), .B1(new_new_n168_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n717_), .B(new_new_n921_), .Y(new_new_n967_));
  AOI210     g0945(.A0(new_new_n966_), .A1(new_new_n354_), .B0(new_new_n967_), .Y(new_new_n968_));
  NA2        g0946(.A(new_new_n764_), .B(new_new_n138_), .Y(new_new_n969_));
  INV        g0947(.A(new_new_n969_), .Y(new_new_n970_));
  NA2        g0948(.A(new_new_n970_), .B(new_new_n704_), .Y(new_new_n971_));
  NO2        g0949(.A(new_new_n823_), .B(new_new_n415_), .Y(new_new_n972_));
  NA3        g0950(.A(new_new_n852_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n973_));
  AOI210     g0951(.A0(new_new_n973_), .A1(new_new_n516_), .B0(new_new_n1091_), .Y(new_new_n974_));
  NO2        g0952(.A(new_new_n974_), .B(new_new_n972_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n975_), .B(new_new_n971_), .C(new_new_n968_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n936_), .B(new_new_n383_), .Y(new_new_n977_));
  AOI210     g0955(.A0(new_new_n302_), .A1(new_new_n155_), .B0(new_new_n977_), .Y(new_new_n978_));
  NA3        g0956(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n910_), .B(new_new_n505_), .Y(new_new_n980_));
  AOI210     g0958(.A0(new_new_n979_), .A1(new_new_n155_), .B0(new_new_n980_), .Y(new_new_n981_));
  NO2        g0959(.A(new_new_n981_), .B(new_new_n978_), .Y(new_new_n982_));
  NO3        g0960(.A(new_new_n896_), .B(new_new_n869_), .C(new_new_n185_), .Y(new_new_n983_));
  NA2        g0961(.A(new_new_n983_), .B(i_11_), .Y(new_new_n984_));
  INV        g0962(.A(new_new_n214_), .Y(new_new_n985_));
  OAI220     g0963(.A0(new_new_n557_), .A1(new_new_n1090_), .B0(new_new_n677_), .B1(new_new_n648_), .Y(new_new_n986_));
  NA3        g0964(.A(new_new_n986_), .B(new_new_n410_), .C(new_new_n985_), .Y(new_new_n987_));
  NA3        g0965(.A(new_new_n987_), .B(new_new_n984_), .C(new_new_n982_), .Y(new_new_n988_));
  NO2        g0966(.A(new_new_n240_), .B(new_new_n88_), .Y(new_new_n989_));
  NA2        g0967(.A(new_new_n989_), .B(new_new_n963_), .Y(new_new_n990_));
  AOI220     g0968(.A0(new_new_n926_), .A1(new_new_n505_), .B0(new_new_n852_), .B1(new_new_n156_), .Y(new_new_n991_));
  NA2        g0969(.A(new_new_n357_), .B(new_new_n170_), .Y(new_new_n992_));
  OA220      g0970(.A0(new_new_n992_), .A1(new_new_n991_), .B0(new_new_n990_), .B1(i_5_), .Y(new_new_n993_));
  AOI210     g0971(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n169_), .Y(new_new_n994_));
  NA2        g0972(.A(new_new_n994_), .B(new_new_n940_), .Y(new_new_n995_));
  NA3        g0973(.A(new_new_n645_), .B(new_new_n180_), .C(new_new_n79_), .Y(new_new_n996_));
  NA2        g0974(.A(new_new_n996_), .B(new_new_n574_), .Y(new_new_n997_));
  NO3        g0975(.A(new_new_n862_), .B(new_new_n52_), .C(new_new_n48_), .Y(new_new_n998_));
  NO3        g0976(.A(new_new_n1079_), .B(new_new_n998_), .C(new_new_n997_), .Y(new_new_n999_));
  NA3        g0977(.A(new_new_n401_), .B(new_new_n165_), .C(new_new_n164_), .Y(new_new_n1000_));
  NA3        g0978(.A(new_new_n910_), .B(new_new_n291_), .C(new_new_n227_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n1001_), .B(new_new_n1000_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n401_), .B(new_new_n338_), .C(new_new_n218_), .Y(new_new_n1003_));
  INV        g0981(.A(new_new_n1003_), .Y(new_new_n1004_));
  NOi31      g0982(.An(new_new_n400_), .B(new_new_n964_), .C(new_new_n237_), .Y(new_new_n1005_));
  NO3        g0983(.A(new_new_n907_), .B(new_new_n214_), .C(new_new_n185_), .Y(new_new_n1006_));
  NO4        g0984(.A(new_new_n1006_), .B(new_new_n1005_), .C(new_new_n1004_), .D(new_new_n1002_), .Y(new_new_n1007_));
  NA4        g0985(.A(new_new_n1007_), .B(new_new_n999_), .C(new_new_n995_), .D(new_new_n993_), .Y(new_new_n1008_));
  INV        g0986(.A(new_new_n647_), .Y(new_new_n1009_));
  NO3        g0987(.A(new_new_n1009_), .B(new_new_n588_), .C(new_new_n351_), .Y(new_new_n1010_));
  NA3        g0988(.A(new_new_n853_), .B(new_new_n104_), .C(new_new_n119_), .Y(new_new_n1011_));
  INV        g0989(.A(new_new_n1011_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n1012_), .A1(new_new_n1087_), .B0(new_new_n1010_), .Y(new_new_n1013_));
  NA3        g0991(.A(new_new_n307_), .B(i_5_), .C(new_new_n188_), .Y(new_new_n1014_));
  NAi31      g0992(.An(new_new_n239_), .B(new_new_n1014_), .C(new_new_n240_), .Y(new_new_n1015_));
  NO4        g0993(.A(new_new_n237_), .B(new_new_n205_), .C(i_0_), .D(i_12_), .Y(new_new_n1016_));
  AOI220     g0994(.A0(new_new_n1016_), .A1(new_new_n1015_), .B0(new_new_n803_), .B1(new_new_n170_), .Y(new_new_n1017_));
  AN2        g0995(.A(new_new_n896_), .B(new_new_n146_), .Y(new_new_n1018_));
  NO4        g0996(.A(new_new_n1018_), .B(i_12_), .C(new_new_n681_), .D(new_new_n125_), .Y(new_new_n1019_));
  NA2        g0997(.A(new_new_n1019_), .B(new_new_n214_), .Y(new_new_n1020_));
  NA3        g0998(.A(new_new_n92_), .B(new_new_n602_), .C(i_11_), .Y(new_new_n1021_));
  NO2        g0999(.A(new_new_n1021_), .B(new_new_n148_), .Y(new_new_n1022_));
  NA2        g1000(.A(new_new_n926_), .B(new_new_n491_), .Y(new_new_n1023_));
  OAI220     g1001(.A0(i_7_), .A1(new_new_n1014_), .B0(new_new_n1023_), .B1(new_new_n705_), .Y(new_new_n1024_));
  AOI210     g1002(.A0(new_new_n1024_), .A1(new_new_n914_), .B0(new_new_n1022_), .Y(new_new_n1025_));
  NA4        g1003(.A(new_new_n1025_), .B(new_new_n1020_), .C(new_new_n1017_), .D(new_new_n1013_), .Y(new_new_n1026_));
  NO4        g1004(.A(new_new_n1026_), .B(new_new_n1008_), .C(new_new_n988_), .D(new_new_n976_), .Y(new_new_n1027_));
  OAI210     g1005(.A0(new_new_n826_), .A1(new_new_n819_), .B0(new_new_n36_), .Y(new_new_n1028_));
  NA3        g1006(.A(new_new_n920_), .B(new_new_n378_), .C(i_5_), .Y(new_new_n1029_));
  NA3        g1007(.A(new_new_n1029_), .B(new_new_n1028_), .C(new_new_n643_), .Y(new_new_n1030_));
  NA2        g1008(.A(new_new_n1030_), .B(new_new_n202_), .Y(new_new_n1031_));
  AN2        g1009(.A(new_new_n727_), .B(new_new_n379_), .Y(new_new_n1032_));
  NA2        g1010(.A(new_new_n181_), .B(new_new_n183_), .Y(new_new_n1033_));
  AO210      g1011(.A0(new_new_n1032_), .A1(new_new_n32_), .B0(new_new_n1033_), .Y(new_new_n1034_));
  OAI210     g1012(.A0(new_new_n647_), .A1(new_new_n645_), .B0(new_new_n319_), .Y(new_new_n1035_));
  NAi31      g1013(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1036_));
  INV        g1014(.A(new_new_n1036_), .Y(new_new_n1037_));
  NO2        g1015(.A(new_new_n1037_), .B(new_new_n678_), .Y(new_new_n1038_));
  NA3        g1016(.A(new_new_n1038_), .B(new_new_n1035_), .C(new_new_n1034_), .Y(new_new_n1039_));
  NO2        g1017(.A(new_new_n481_), .B(new_new_n268_), .Y(new_new_n1040_));
  NO4        g1018(.A(new_new_n230_), .B(new_new_n137_), .C(new_new_n708_), .D(new_new_n36_), .Y(new_new_n1041_));
  NO3        g1019(.A(new_new_n1041_), .B(new_new_n1040_), .C(new_new_n888_), .Y(new_new_n1042_));
  OAI210     g1020(.A0(new_new_n1021_), .A1(new_new_n140_), .B0(new_new_n1042_), .Y(new_new_n1043_));
  AOI210     g1021(.A0(new_new_n1039_), .A1(new_new_n48_), .B0(new_new_n1043_), .Y(new_new_n1044_));
  AOI210     g1022(.A0(new_new_n1044_), .A1(new_new_n1031_), .B0(new_new_n69_), .Y(new_new_n1045_));
  NO2        g1023(.A(new_new_n595_), .B(new_new_n390_), .Y(new_new_n1046_));
  NO2        g1024(.A(new_new_n1046_), .B(new_new_n778_), .Y(new_new_n1047_));
  OAI210     g1025(.A0(new_new_n75_), .A1(new_new_n52_), .B0(new_new_n102_), .Y(new_new_n1048_));
  NA2        g1026(.A(new_new_n1048_), .B(new_new_n72_), .Y(new_new_n1049_));
  AOI210     g1027(.A0(new_new_n994_), .A1(new_new_n910_), .B0(new_new_n927_), .Y(new_new_n1050_));
  AOI210     g1028(.A0(new_new_n1050_), .A1(new_new_n1049_), .B0(new_new_n708_), .Y(new_new_n1051_));
  NA2        g1029(.A(new_new_n262_), .B(new_new_n55_), .Y(new_new_n1052_));
  AOI220     g1030(.A0(new_new_n1052_), .A1(new_new_n72_), .B0(new_new_n352_), .B1(new_new_n254_), .Y(new_new_n1053_));
  NO2        g1031(.A(new_new_n1053_), .B(new_new_n234_), .Y(new_new_n1054_));
  NA3        g1032(.A(new_new_n90_), .B(new_new_n309_), .C(new_new_n30_), .Y(new_new_n1055_));
  INV        g1033(.A(new_new_n1055_), .Y(new_new_n1056_));
  NO3        g1034(.A(new_new_n1056_), .B(new_new_n1054_), .C(new_new_n1051_), .Y(new_new_n1057_));
  OAI210     g1035(.A0(new_new_n270_), .A1(new_new_n151_), .B0(new_new_n84_), .Y(new_new_n1058_));
  NA3        g1036(.A(new_new_n779_), .B(new_new_n291_), .C(new_new_n75_), .Y(new_new_n1059_));
  AOI210     g1037(.A0(new_new_n1059_), .A1(new_new_n1058_), .B0(i_11_), .Y(new_new_n1060_));
  NA2        g1038(.A(new_new_n638_), .B(new_new_n211_), .Y(new_new_n1061_));
  OAI210     g1039(.A0(new_new_n1061_), .A1(new_new_n920_), .B0(new_new_n202_), .Y(new_new_n1062_));
  NA2        g1040(.A(new_new_n157_), .B(i_5_), .Y(new_new_n1063_));
  AOI210     g1041(.A0(new_new_n1062_), .A1(new_new_n791_), .B0(new_new_n1063_), .Y(new_new_n1064_));
  NO3        g1042(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n1065_));
  OAI210     g1043(.A0(new_new_n931_), .A1(new_new_n309_), .B0(new_new_n1065_), .Y(new_new_n1066_));
  NO2        g1044(.A(new_new_n1066_), .B(new_new_n755_), .Y(new_new_n1067_));
  NO4        g1045(.A(new_new_n955_), .B(new_new_n496_), .C(new_new_n251_), .D(new_new_n250_), .Y(new_new_n1068_));
  NO2        g1046(.A(new_new_n1068_), .B(new_new_n592_), .Y(new_new_n1069_));
  NO2        g1047(.A(new_new_n822_), .B(new_new_n371_), .Y(new_new_n1070_));
  AOI210     g1048(.A0(new_new_n1070_), .A1(new_new_n1069_), .B0(new_new_n40_), .Y(new_new_n1071_));
  NO4        g1049(.A(new_new_n1071_), .B(new_new_n1067_), .C(new_new_n1064_), .D(new_new_n1060_), .Y(new_new_n1072_));
  OAI210     g1050(.A0(new_new_n1057_), .A1(i_4_), .B0(new_new_n1072_), .Y(new_new_n1073_));
  NO3        g1051(.A(new_new_n1073_), .B(new_new_n1047_), .C(new_new_n1045_), .Y(new_new_n1074_));
  NA4        g1052(.A(new_new_n1074_), .B(new_new_n1027_), .C(new_new_n962_), .D(new_new_n876_), .Y(men4));
  INV        g1053(.A(i_5_), .Y(new_new_n1078_));
  INV        g1054(.A(new_new_n503_), .Y(new_new_n1079_));
  INV        g1055(.A(i_3_), .Y(new_new_n1080_));
  INV        g1056(.A(i_6_), .Y(new_new_n1081_));
  INV        g1057(.A(new_new_n136_), .Y(new_new_n1082_));
  INV        g1058(.A(new_new_n827_), .Y(new_new_n1083_));
  INV        g1059(.A(new_new_n193_), .Y(new_new_n1084_));
  INV        g1060(.A(new_new_n374_), .Y(new_new_n1085_));
  INV        g1061(.A(i_4_), .Y(new_new_n1086_));
  INV        g1062(.A(i_5_), .Y(new_new_n1087_));
  INV        g1063(.A(i_6_), .Y(new_new_n1088_));
  INV        g1064(.A(i_3_), .Y(new_new_n1089_));
  INV        g1065(.A(i_6_), .Y(new_new_n1090_));
  INV        g1066(.A(i_9_), .Y(new_new_n1091_));
endmodule


