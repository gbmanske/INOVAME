// Benchmark "top" written by ABC on Fri Jun 21 17:49:24 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n137_, new_new_n138_, new_new_n139_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1039_,
    new_new_n1040_, new_new_n1041_, new_new_n1042_, new_new_n1043_,
    new_new_n1044_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g0016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g0017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g0018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g0028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g0029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g0032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(new_new_n65_), .B(new_new_n61_), .Y(new_new_n66_));
  NA2        g0044(.A(new_new_n50_), .B(i_2_), .Y(new_new_n67_));
  NA2        g0045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g0046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g0047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g0048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g0049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g0050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g0051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  INV        g0052(.A(new_new_n74_), .Y(new_new_n75_));
  OAI210     g0053(.A0(new_new_n75_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g0054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NA2        g0055(.A(i_2_), .B(i_8_), .Y(new_new_n78_));
  NO2        g0056(.A(new_new_n78_), .B(new_new_n58_), .Y(new_new_n79_));
  NO2        g0057(.A(i_3_), .B(i_9_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_7_), .Y(new_new_n81_));
  INV        g0059(.A(i_6_), .Y(new_new_n82_));
  OR4        g0060(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n83_));
  INV        g0061(.A(new_new_n83_), .Y(new_new_n84_));
  NO2        g0062(.A(i_2_), .B(i_7_), .Y(new_new_n85_));
  INV        g0063(.A(new_new_n79_), .Y(new_new_n86_));
  NAi21      g0064(.An(i_6_), .B(i_10_), .Y(new_new_n87_));
  NA2        g0065(.A(i_6_), .B(i_9_), .Y(new_new_n88_));
  AOI210     g0066(.A0(new_new_n88_), .A1(new_new_n87_), .B0(new_new_n63_), .Y(new_new_n89_));
  NA2        g0067(.A(i_2_), .B(i_6_), .Y(new_new_n90_));
  NO3        g0068(.A(new_new_n90_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n91_));
  NO2        g0069(.A(new_new_n91_), .B(new_new_n89_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n92_), .A1(new_new_n86_), .B0(new_new_n77_), .Y(new_new_n93_));
  AN3        g0071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n94_));
  NAi21      g0072(.An(i_6_), .B(i_11_), .Y(new_new_n95_));
  NO2        g0073(.A(i_5_), .B(i_8_), .Y(new_new_n96_));
  NOi21      g0074(.An(new_new_n96_), .B(new_new_n95_), .Y(new_new_n97_));
  AOI220     g0075(.A0(new_new_n97_), .A1(new_new_n62_), .B0(new_new_n94_), .B1(new_new_n32_), .Y(new_new_n98_));
  INV        g0076(.A(i_7_), .Y(new_new_n99_));
  NA2        g0077(.A(new_new_n46_), .B(new_new_n99_), .Y(new_new_n100_));
  NO2        g0078(.A(i_0_), .B(i_5_), .Y(new_new_n101_));
  NO2        g0079(.A(new_new_n101_), .B(new_new_n82_), .Y(new_new_n102_));
  NA2        g0080(.A(i_12_), .B(i_3_), .Y(new_new_n103_));
  INV        g0081(.A(new_new_n103_), .Y(new_new_n104_));
  NA3        g0082(.A(new_new_n104_), .B(new_new_n102_), .C(new_new_n100_), .Y(new_new_n105_));
  NAi21      g0083(.An(i_7_), .B(i_11_), .Y(new_new_n106_));
  NO3        g0084(.A(new_new_n106_), .B(new_new_n87_), .C(new_new_n53_), .Y(new_new_n107_));
  AN2        g0085(.A(i_2_), .B(i_10_), .Y(new_new_n108_));
  NO2        g0086(.A(new_new_n108_), .B(i_7_), .Y(new_new_n109_));
  OR2        g0087(.A(new_new_n77_), .B(new_new_n58_), .Y(new_new_n110_));
  NO2        g0088(.A(i_8_), .B(new_new_n99_), .Y(new_new_n111_));
  NO3        g0089(.A(new_new_n111_), .B(new_new_n110_), .C(new_new_n109_), .Y(new_new_n112_));
  NA2        g0090(.A(i_12_), .B(i_7_), .Y(new_new_n113_));
  NO2        g0091(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n114_));
  NA2        g0092(.A(new_new_n114_), .B(i_0_), .Y(new_new_n115_));
  NA2        g0093(.A(i_11_), .B(i_12_), .Y(new_new_n116_));
  OAI210     g0094(.A0(new_new_n115_), .A1(new_new_n113_), .B0(new_new_n116_), .Y(new_new_n117_));
  NO2        g0095(.A(new_new_n117_), .B(new_new_n112_), .Y(new_new_n118_));
  NAi41      g0096(.An(new_new_n107_), .B(new_new_n118_), .C(new_new_n105_), .D(new_new_n98_), .Y(new_new_n119_));
  NOi21      g0097(.An(i_1_), .B(i_5_), .Y(new_new_n120_));
  NA2        g0098(.A(new_new_n120_), .B(i_11_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n122_));
  NA2        g0100(.A(i_7_), .B(new_new_n25_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n123_), .B(new_new_n122_), .Y(new_new_n124_));
  NO2        g0102(.A(new_new_n124_), .B(new_new_n46_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n88_), .B(new_new_n87_), .Y(new_new_n126_));
  NAi21      g0104(.An(i_3_), .B(i_8_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n127_), .B(new_new_n62_), .Y(new_new_n128_));
  NOi21      g0106(.An(new_new_n128_), .B(new_new_n126_), .Y(new_new_n129_));
  NO2        g0107(.A(i_1_), .B(new_new_n82_), .Y(new_new_n130_));
  NO2        g0108(.A(i_6_), .B(i_5_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n131_), .B(i_3_), .Y(new_new_n132_));
  AO210      g0110(.A0(new_new_n132_), .A1(new_new_n47_), .B0(new_new_n130_), .Y(new_new_n133_));
  OAI220     g0111(.A0(new_new_n133_), .A1(new_new_n106_), .B0(new_new_n129_), .B1(new_new_n121_), .Y(new_new_n134_));
  NO3        g0112(.A(new_new_n134_), .B(new_new_n119_), .C(new_new_n93_), .Y(new_new_n135_));
  NA3        g0113(.A(new_new_n135_), .B(new_new_n76_), .C(new_new_n56_), .Y(men2));
  NO2        g0114(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n137_));
  NA2        g0115(.A(i_6_), .B(new_new_n25_), .Y(new_new_n138_));
  NA2        g0116(.A(new_new_n138_), .B(new_new_n137_), .Y(new_new_n139_));
  NA4        g0117(.A(new_new_n139_), .B(new_new_n74_), .C(new_new_n67_), .D(new_new_n30_), .Y(men0));
  AN2        g0118(.A(i_8_), .B(i_7_), .Y(new_new_n141_));
  NA2        g0119(.A(new_new_n141_), .B(i_6_), .Y(new_new_n142_));
  NO2        g0120(.A(i_12_), .B(i_13_), .Y(new_new_n143_));
  NAi21      g0121(.An(i_5_), .B(i_11_), .Y(new_new_n144_));
  NOi21      g0122(.An(new_new_n143_), .B(new_new_n144_), .Y(new_new_n145_));
  NO2        g0123(.A(i_0_), .B(i_1_), .Y(new_new_n146_));
  NA2        g0124(.A(i_2_), .B(i_3_), .Y(new_new_n147_));
  NO2        g0125(.A(new_new_n147_), .B(i_4_), .Y(new_new_n148_));
  NA3        g0126(.A(new_new_n148_), .B(new_new_n146_), .C(new_new_n145_), .Y(new_new_n149_));
  OR2        g0127(.A(new_new_n149_), .B(new_new_n25_), .Y(new_new_n150_));
  AN2        g0128(.A(new_new_n143_), .B(new_new_n80_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(new_new_n27_), .Y(new_new_n152_));
  NA2        g0130(.A(i_1_), .B(i_5_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n70_), .B(new_new_n46_), .Y(new_new_n154_));
  NA2        g0132(.A(new_new_n154_), .B(new_new_n36_), .Y(new_new_n155_));
  NO3        g0133(.A(new_new_n155_), .B(new_new_n153_), .C(new_new_n152_), .Y(new_new_n156_));
  OR2        g0134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n77_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g0137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g0138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g0139(.A(new_new_n161_), .B(new_new_n39_), .Y(new_new_n162_));
  NO2        g0140(.A(i_3_), .B(i_5_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n70_), .B(i_2_), .C(i_1_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  OAI210     g0143(.A0(new_new_n165_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n166_));
  NO2        g0144(.A(new_new_n166_), .B(new_new_n156_), .Y(new_new_n167_));
  AOI210     g0145(.A0(new_new_n167_), .A1(new_new_n150_), .B0(new_new_n142_), .Y(new_new_n168_));
  NA3        g0146(.A(new_new_n70_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n169_));
  NOi21      g0147(.An(i_4_), .B(i_9_), .Y(new_new_n170_));
  NOi21      g0148(.An(i_11_), .B(i_13_), .Y(new_new_n171_));
  NA2        g0149(.A(new_new_n171_), .B(new_new_n170_), .Y(new_new_n172_));
  NO2        g0150(.A(i_4_), .B(i_5_), .Y(new_new_n173_));
  NAi21      g0151(.An(i_12_), .B(i_11_), .Y(new_new_n174_));
  NO2        g0152(.A(new_new_n174_), .B(i_13_), .Y(new_new_n175_));
  NA3        g0153(.A(new_new_n175_), .B(new_new_n173_), .C(new_new_n80_), .Y(new_new_n176_));
  AOI210     g0154(.A0(new_new_n176_), .A1(new_new_n172_), .B0(new_new_n169_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n70_), .B(new_new_n63_), .Y(new_new_n178_));
  NA2        g0156(.A(new_new_n36_), .B(i_5_), .Y(new_new_n179_));
  NAi31      g0157(.An(new_new_n179_), .B(new_new_n151_), .C(i_11_), .Y(new_new_n180_));
  NA2        g0158(.A(i_3_), .B(i_5_), .Y(new_new_n181_));
  OR2        g0159(.A(new_new_n181_), .B(new_new_n172_), .Y(new_new_n182_));
  AOI210     g0160(.A0(new_new_n182_), .A1(new_new_n180_), .B0(i_2_), .Y(new_new_n183_));
  NO2        g0161(.A(new_new_n70_), .B(i_5_), .Y(new_new_n184_));
  NO2        g0162(.A(i_13_), .B(i_10_), .Y(new_new_n185_));
  NA3        g0163(.A(new_new_n185_), .B(new_new_n184_), .C(new_new_n44_), .Y(new_new_n186_));
  NO2        g0164(.A(i_2_), .B(i_1_), .Y(new_new_n187_));
  NA2        g0165(.A(new_new_n187_), .B(i_3_), .Y(new_new_n188_));
  NAi21      g0166(.An(i_4_), .B(i_12_), .Y(new_new_n189_));
  NO4        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n186_), .D(new_new_n25_), .Y(new_new_n190_));
  NO3        g0168(.A(new_new_n190_), .B(new_new_n183_), .C(new_new_n177_), .Y(new_new_n191_));
  INV        g0169(.A(i_8_), .Y(new_new_n192_));
  NO2        g0170(.A(new_new_n192_), .B(i_7_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_6_), .Y(new_new_n194_));
  NO3        g0172(.A(i_3_), .B(new_new_n82_), .C(new_new_n48_), .Y(new_new_n195_));
  NA2        g0173(.A(new_new_n195_), .B(new_new_n111_), .Y(new_new_n196_));
  NO3        g0174(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n197_));
  NA3        g0175(.A(new_new_n197_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n198_));
  NO3        g0176(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n199_));
  OAI210     g0177(.A0(new_new_n94_), .A1(i_12_), .B0(new_new_n199_), .Y(new_new_n200_));
  AOI210     g0178(.A0(new_new_n200_), .A1(new_new_n198_), .B0(new_new_n196_), .Y(new_new_n201_));
  NO2        g0179(.A(i_3_), .B(i_8_), .Y(new_new_n202_));
  NO3        g0180(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n203_));
  NA3        g0181(.A(new_new_n203_), .B(new_new_n202_), .C(new_new_n39_), .Y(new_new_n204_));
  NO2        g0182(.A(new_new_n101_), .B(new_new_n58_), .Y(new_new_n205_));
  INV        g0183(.A(new_new_n205_), .Y(new_new_n206_));
  NO2        g0184(.A(i_13_), .B(i_9_), .Y(new_new_n207_));
  NAi21      g0185(.An(i_12_), .B(i_3_), .Y(new_new_n208_));
  NO2        g0186(.A(new_new_n44_), .B(i_5_), .Y(new_new_n209_));
  NO3        g0187(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n210_));
  NA2        g0188(.A(new_new_n210_), .B(i_10_), .Y(new_new_n211_));
  OAI220     g0189(.A0(new_new_n211_), .A1(new_new_n208_), .B0(new_new_n206_), .B1(new_new_n204_), .Y(new_new_n212_));
  AOI210     g0190(.A0(new_new_n212_), .A1(i_7_), .B0(new_new_n201_), .Y(new_new_n213_));
  OAI220     g0191(.A0(new_new_n213_), .A1(i_4_), .B0(new_new_n194_), .B1(new_new_n191_), .Y(new_new_n214_));
  NAi21      g0192(.An(i_12_), .B(i_7_), .Y(new_new_n215_));
  NA3        g0193(.A(i_13_), .B(new_new_n192_), .C(i_10_), .Y(new_new_n216_));
  NO2        g0194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NA2        g0195(.A(i_0_), .B(i_5_), .Y(new_new_n218_));
  NA2        g0196(.A(new_new_n218_), .B(new_new_n102_), .Y(new_new_n219_));
  OAI220     g0197(.A0(new_new_n219_), .A1(new_new_n188_), .B0(i_2_), .B1(new_new_n132_), .Y(new_new_n220_));
  NAi31      g0198(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n36_), .B(i_13_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n70_), .B(new_new_n26_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n224_));
  NA3        g0202(.A(new_new_n224_), .B(new_new_n223_), .C(new_new_n222_), .Y(new_new_n225_));
  INV        g0203(.A(i_13_), .Y(new_new_n226_));
  NO2        g0204(.A(i_12_), .B(new_new_n226_), .Y(new_new_n227_));
  NA3        g0205(.A(new_new_n227_), .B(new_new_n197_), .C(new_new_n195_), .Y(new_new_n228_));
  OAI210     g0206(.A0(new_new_n225_), .A1(new_new_n221_), .B0(new_new_n228_), .Y(new_new_n229_));
  AOI220     g0207(.A0(new_new_n229_), .A1(new_new_n141_), .B0(new_new_n220_), .B1(new_new_n217_), .Y(new_new_n230_));
  NO2        g0208(.A(i_12_), .B(new_new_n37_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n181_), .B(i_4_), .Y(new_new_n232_));
  NA2        g0210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  OR2        g0211(.A(i_8_), .B(i_7_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n234_), .B(new_new_n82_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n53_), .B(i_1_), .Y(new_new_n236_));
  NA2        g0214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  INV        g0215(.A(i_12_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n44_), .B(new_new_n238_), .Y(new_new_n239_));
  NO3        g0217(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n240_));
  NA2        g0218(.A(i_2_), .B(i_1_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n237_), .B(new_new_n233_), .Y(new_new_n242_));
  NO3        g0220(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n243_));
  NAi21      g0221(.An(i_4_), .B(i_3_), .Y(new_new_n244_));
  NO2        g0222(.A(i_0_), .B(i_6_), .Y(new_new_n245_));
  NOi41      g0223(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n246_));
  NA2        g0224(.A(new_new_n246_), .B(new_new_n245_), .Y(new_new_n247_));
  NO2        g0225(.A(new_new_n241_), .B(new_new_n181_), .Y(new_new_n248_));
  NAi21      g0226(.An(new_new_n247_), .B(new_new_n248_), .Y(new_new_n249_));
  INV        g0227(.A(new_new_n249_), .Y(new_new_n250_));
  NO2        g0228(.A(new_new_n250_), .B(new_new_n242_), .Y(new_new_n251_));
  NO2        g0229(.A(i_11_), .B(new_new_n226_), .Y(new_new_n252_));
  NOi21      g0230(.An(i_1_), .B(i_6_), .Y(new_new_n253_));
  NAi21      g0231(.An(i_3_), .B(i_7_), .Y(new_new_n254_));
  NA2        g0232(.A(new_new_n238_), .B(i_9_), .Y(new_new_n255_));
  OR4        g0233(.A(new_new_n255_), .B(new_new_n254_), .C(new_new_n253_), .D(new_new_n184_), .Y(new_new_n256_));
  NO2        g0234(.A(i_12_), .B(i_3_), .Y(new_new_n257_));
  NA2        g0235(.A(new_new_n70_), .B(i_5_), .Y(new_new_n258_));
  NA2        g0236(.A(i_3_), .B(i_9_), .Y(new_new_n259_));
  NAi21      g0237(.An(i_7_), .B(i_10_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n260_), .B(new_new_n259_), .Y(new_new_n261_));
  NA3        g0239(.A(new_new_n261_), .B(new_new_n258_), .C(new_new_n64_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n262_), .B(new_new_n256_), .Y(new_new_n263_));
  NA3        g0241(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n264_));
  INV        g0242(.A(new_new_n142_), .Y(new_new_n265_));
  NA2        g0243(.A(new_new_n238_), .B(i_13_), .Y(new_new_n266_));
  NO2        g0244(.A(new_new_n266_), .B(new_new_n72_), .Y(new_new_n267_));
  AOI220     g0245(.A0(new_new_n267_), .A1(new_new_n265_), .B0(new_new_n263_), .B1(new_new_n252_), .Y(new_new_n268_));
  NO2        g0246(.A(new_new_n234_), .B(new_new_n37_), .Y(new_new_n269_));
  NA2        g0247(.A(i_12_), .B(i_6_), .Y(new_new_n270_));
  OR2        g0248(.A(i_13_), .B(i_9_), .Y(new_new_n271_));
  NO3        g0249(.A(new_new_n271_), .B(new_new_n270_), .C(new_new_n48_), .Y(new_new_n272_));
  NO2        g0250(.A(new_new_n244_), .B(i_2_), .Y(new_new_n273_));
  NA3        g0251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n44_), .Y(new_new_n274_));
  NA2        g0252(.A(new_new_n252_), .B(i_9_), .Y(new_new_n275_));
  OAI210     g0253(.A0(new_new_n70_), .A1(new_new_n275_), .B0(new_new_n274_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n154_), .B(new_new_n63_), .Y(new_new_n277_));
  NO3        g0255(.A(i_11_), .B(new_new_n226_), .C(new_new_n25_), .Y(new_new_n278_));
  NO2        g0256(.A(new_new_n254_), .B(i_8_), .Y(new_new_n279_));
  NO2        g0257(.A(i_6_), .B(new_new_n48_), .Y(new_new_n280_));
  NA3        g0258(.A(new_new_n280_), .B(new_new_n279_), .C(new_new_n278_), .Y(new_new_n281_));
  NA3        g0259(.A(i_6_), .B(new_new_n269_), .C(new_new_n227_), .Y(new_new_n282_));
  AOI210     g0260(.A0(new_new_n282_), .A1(new_new_n281_), .B0(new_new_n277_), .Y(new_new_n283_));
  AOI210     g0261(.A0(new_new_n276_), .A1(new_new_n269_), .B0(new_new_n283_), .Y(new_new_n284_));
  NA4        g0262(.A(new_new_n284_), .B(new_new_n268_), .C(new_new_n251_), .D(new_new_n230_), .Y(new_new_n285_));
  NO3        g0263(.A(i_12_), .B(new_new_n226_), .C(new_new_n37_), .Y(new_new_n286_));
  INV        g0264(.A(new_new_n286_), .Y(new_new_n287_));
  NA2        g0265(.A(i_8_), .B(new_new_n99_), .Y(new_new_n288_));
  NOi21      g0266(.An(new_new_n163_), .B(new_new_n82_), .Y(new_new_n289_));
  NO3        g0267(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n290_));
  AOI220     g0268(.A0(new_new_n290_), .A1(new_new_n195_), .B0(new_new_n289_), .B1(new_new_n236_), .Y(new_new_n291_));
  NO2        g0269(.A(new_new_n291_), .B(new_new_n288_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n241_), .B(i_0_), .Y(new_new_n293_));
  AOI220     g0271(.A0(new_new_n293_), .A1(new_new_n193_), .B0(i_1_), .B1(new_new_n141_), .Y(new_new_n294_));
  NA2        g0272(.A(new_new_n280_), .B(new_new_n26_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n295_), .B(new_new_n294_), .Y(new_new_n296_));
  NA2        g0274(.A(i_0_), .B(i_1_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(i_2_), .Y(new_new_n298_));
  NO2        g0276(.A(new_new_n59_), .B(i_6_), .Y(new_new_n299_));
  NA3        g0277(.A(new_new_n299_), .B(new_new_n298_), .C(new_new_n163_), .Y(new_new_n300_));
  OAI210     g0278(.A0(new_new_n165_), .A1(new_new_n142_), .B0(new_new_n300_), .Y(new_new_n301_));
  NO3        g0279(.A(new_new_n301_), .B(new_new_n296_), .C(new_new_n292_), .Y(new_new_n302_));
  NO2        g0280(.A(i_3_), .B(i_10_), .Y(new_new_n303_));
  NA3        g0281(.A(new_new_n303_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n304_));
  NO2        g0282(.A(i_2_), .B(new_new_n99_), .Y(new_new_n305_));
  NA2        g0283(.A(i_1_), .B(new_new_n36_), .Y(new_new_n306_));
  NOi21      g0284(.An(new_new_n218_), .B(new_new_n101_), .Y(new_new_n307_));
  NA3        g0285(.A(new_new_n307_), .B(i_1_), .C(new_new_n305_), .Y(new_new_n308_));
  AN2        g0286(.A(i_3_), .B(i_10_), .Y(new_new_n309_));
  NA3        g0287(.A(new_new_n309_), .B(new_new_n175_), .C(new_new_n173_), .Y(new_new_n310_));
  NO2        g0288(.A(i_5_), .B(new_new_n37_), .Y(new_new_n311_));
  NO2        g0289(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n312_));
  OR2        g0290(.A(new_new_n308_), .B(new_new_n304_), .Y(new_new_n313_));
  OAI220     g0291(.A0(new_new_n313_), .A1(i_6_), .B0(new_new_n302_), .B1(new_new_n287_), .Y(new_new_n314_));
  NO4        g0292(.A(new_new_n314_), .B(new_new_n285_), .C(new_new_n214_), .D(new_new_n168_), .Y(new_new_n315_));
  NO3        g0293(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n316_));
  NO2        g0294(.A(new_new_n59_), .B(new_new_n82_), .Y(new_new_n317_));
  NA2        g0295(.A(new_new_n293_), .B(new_new_n317_), .Y(new_new_n318_));
  NO3        g0296(.A(i_6_), .B(new_new_n192_), .C(i_7_), .Y(new_new_n319_));
  NA2        g0297(.A(new_new_n319_), .B(new_new_n197_), .Y(new_new_n320_));
  AOI210     g0298(.A0(new_new_n320_), .A1(new_new_n318_), .B0(i_5_), .Y(new_new_n321_));
  NO2        g0299(.A(i_2_), .B(i_3_), .Y(new_new_n322_));
  OR2        g0300(.A(i_0_), .B(i_5_), .Y(new_new_n323_));
  NA2        g0301(.A(new_new_n218_), .B(new_new_n323_), .Y(new_new_n324_));
  NA4        g0302(.A(new_new_n324_), .B(new_new_n235_), .C(new_new_n322_), .D(i_1_), .Y(new_new_n325_));
  NA3        g0303(.A(new_new_n293_), .B(new_new_n289_), .C(new_new_n111_), .Y(new_new_n326_));
  NAi21      g0304(.An(i_8_), .B(i_7_), .Y(new_new_n327_));
  NO2        g0305(.A(new_new_n327_), .B(i_6_), .Y(new_new_n328_));
  NO2        g0306(.A(new_new_n157_), .B(new_new_n46_), .Y(new_new_n329_));
  NA3        g0307(.A(new_new_n329_), .B(new_new_n328_), .C(new_new_n163_), .Y(new_new_n330_));
  NA3        g0308(.A(new_new_n330_), .B(new_new_n326_), .C(new_new_n325_), .Y(new_new_n331_));
  OAI210     g0309(.A0(new_new_n331_), .A1(new_new_n321_), .B0(i_4_), .Y(new_new_n332_));
  NO2        g0310(.A(i_12_), .B(i_10_), .Y(new_new_n333_));
  NOi21      g0311(.An(i_5_), .B(i_0_), .Y(new_new_n334_));
  AOI210     g0312(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n99_), .Y(new_new_n335_));
  NO3        g0313(.A(new_new_n335_), .B(new_new_n306_), .C(new_new_n127_), .Y(new_new_n336_));
  NA4        g0314(.A(new_new_n81_), .B(new_new_n36_), .C(new_new_n82_), .D(i_8_), .Y(new_new_n337_));
  NA2        g0315(.A(new_new_n336_), .B(new_new_n333_), .Y(new_new_n338_));
  NO2        g0316(.A(i_6_), .B(i_8_), .Y(new_new_n339_));
  NOi21      g0317(.An(i_0_), .B(i_2_), .Y(new_new_n340_));
  AN2        g0318(.A(new_new_n340_), .B(new_new_n339_), .Y(new_new_n341_));
  NO2        g0319(.A(i_1_), .B(i_7_), .Y(new_new_n342_));
  AO220      g0320(.A0(new_new_n342_), .A1(new_new_n341_), .B0(new_new_n328_), .B1(new_new_n236_), .Y(new_new_n343_));
  NA3        g0321(.A(new_new_n343_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n344_));
  NA3        g0322(.A(new_new_n344_), .B(new_new_n338_), .C(new_new_n332_), .Y(new_new_n345_));
  NO2        g0323(.A(i_8_), .B(new_new_n324_), .Y(new_new_n346_));
  NO2        g0324(.A(new_new_n101_), .B(new_new_n123_), .Y(new_new_n347_));
  OAI210     g0325(.A0(new_new_n347_), .A1(new_new_n346_), .B0(i_3_), .Y(new_new_n348_));
  NO2        g0326(.A(new_new_n297_), .B(new_new_n78_), .Y(new_new_n349_));
  NA2        g0327(.A(new_new_n349_), .B(new_new_n131_), .Y(new_new_n350_));
  NO2        g0328(.A(new_new_n90_), .B(new_new_n192_), .Y(new_new_n351_));
  NA3        g0329(.A(new_new_n307_), .B(new_new_n351_), .C(new_new_n63_), .Y(new_new_n352_));
  AOI210     g0330(.A0(new_new_n352_), .A1(new_new_n350_), .B0(i_7_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n192_), .B(i_9_), .Y(new_new_n354_));
  NA2        g0332(.A(new_new_n354_), .B(new_new_n205_), .Y(new_new_n355_));
  NO2        g0333(.A(new_new_n353_), .B(new_new_n296_), .Y(new_new_n356_));
  AOI210     g0334(.A0(new_new_n356_), .A1(new_new_n348_), .B0(new_new_n162_), .Y(new_new_n357_));
  AOI210     g0335(.A0(new_new_n345_), .A1(new_new_n316_), .B0(new_new_n357_), .Y(new_new_n358_));
  NOi32      g0336(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n359_));
  INV        g0337(.A(new_new_n359_), .Y(new_new_n360_));
  NAi21      g0338(.An(i_0_), .B(i_6_), .Y(new_new_n361_));
  NAi21      g0339(.An(i_1_), .B(i_5_), .Y(new_new_n362_));
  NA2        g0340(.A(new_new_n362_), .B(new_new_n361_), .Y(new_new_n363_));
  NA2        g0341(.A(new_new_n363_), .B(new_new_n25_), .Y(new_new_n364_));
  OAI210     g0342(.A0(new_new_n364_), .A1(new_new_n159_), .B0(new_new_n247_), .Y(new_new_n365_));
  NAi41      g0343(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n366_));
  OAI220     g0344(.A0(new_new_n366_), .A1(new_new_n362_), .B0(new_new_n221_), .B1(new_new_n159_), .Y(new_new_n367_));
  AOI210     g0345(.A0(new_new_n366_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n368_));
  NOi32      g0346(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n369_));
  NA2        g0347(.A(new_new_n369_), .B(new_new_n46_), .Y(new_new_n370_));
  NO2        g0348(.A(new_new_n370_), .B(i_0_), .Y(new_new_n371_));
  OR3        g0349(.A(new_new_n371_), .B(new_new_n368_), .C(new_new_n367_), .Y(new_new_n372_));
  NO2        g0350(.A(i_1_), .B(new_new_n99_), .Y(new_new_n373_));
  NAi21      g0351(.An(i_3_), .B(i_4_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n374_), .B(i_9_), .Y(new_new_n375_));
  AN2        g0353(.A(i_6_), .B(i_7_), .Y(new_new_n376_));
  OAI210     g0354(.A0(new_new_n376_), .A1(new_new_n373_), .B0(new_new_n375_), .Y(new_new_n377_));
  NA2        g0355(.A(i_2_), .B(i_7_), .Y(new_new_n378_));
  NO2        g0356(.A(new_new_n374_), .B(i_10_), .Y(new_new_n379_));
  NA3        g0357(.A(new_new_n379_), .B(new_new_n378_), .C(new_new_n245_), .Y(new_new_n380_));
  AOI210     g0358(.A0(new_new_n380_), .A1(new_new_n377_), .B0(new_new_n184_), .Y(new_new_n381_));
  AOI220     g0359(.A0(new_new_n379_), .A1(new_new_n342_), .B0(new_new_n240_), .B1(new_new_n187_), .Y(new_new_n382_));
  NO3        g0360(.A(new_new_n381_), .B(new_new_n372_), .C(new_new_n365_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n383_), .B(new_new_n360_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n385_));
  AN2        g0363(.A(i_12_), .B(i_5_), .Y(new_new_n386_));
  NO2        g0364(.A(i_4_), .B(new_new_n26_), .Y(new_new_n387_));
  NA2        g0365(.A(new_new_n387_), .B(new_new_n386_), .Y(new_new_n388_));
  NO2        g0366(.A(i_11_), .B(i_6_), .Y(new_new_n389_));
  NA3        g0367(.A(new_new_n389_), .B(new_new_n329_), .C(new_new_n226_), .Y(new_new_n390_));
  NO2        g0368(.A(new_new_n390_), .B(new_new_n388_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n244_), .B(i_5_), .Y(new_new_n392_));
  NO2        g0370(.A(i_5_), .B(i_10_), .Y(new_new_n393_));
  NA2        g0371(.A(new_new_n143_), .B(new_new_n45_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n394_), .B(new_new_n244_), .Y(new_new_n395_));
  OAI210     g0373(.A0(new_new_n395_), .A1(new_new_n391_), .B0(new_new_n385_), .Y(new_new_n396_));
  NO2        g0374(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n397_));
  INV        g0375(.A(new_new_n149_), .Y(new_new_n398_));
  OAI210     g0376(.A0(new_new_n398_), .A1(new_new_n391_), .B0(new_new_n397_), .Y(new_new_n399_));
  NO2        g0377(.A(i_3_), .B(new_new_n99_), .Y(new_new_n400_));
  NA2        g0378(.A(new_new_n303_), .B(new_new_n72_), .Y(new_new_n401_));
  NO2        g0379(.A(i_11_), .B(i_12_), .Y(new_new_n402_));
  NA2        g0380(.A(new_new_n402_), .B(new_new_n36_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n401_), .B(new_new_n403_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n393_), .B(new_new_n238_), .Y(new_new_n405_));
  NA3        g0383(.A(new_new_n111_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n406_), .B(new_new_n221_), .Y(new_new_n407_));
  NAi21      g0385(.An(i_13_), .B(i_0_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n408_), .B(new_new_n241_), .Y(new_new_n409_));
  OAI210     g0387(.A0(new_new_n407_), .A1(new_new_n404_), .B0(new_new_n409_), .Y(new_new_n410_));
  NA3        g0388(.A(new_new_n410_), .B(new_new_n399_), .C(new_new_n396_), .Y(new_new_n411_));
  NO3        g0389(.A(i_1_), .B(i_12_), .C(new_new_n82_), .Y(new_new_n412_));
  NO2        g0390(.A(i_0_), .B(i_11_), .Y(new_new_n413_));
  AN2        g0391(.A(i_1_), .B(i_6_), .Y(new_new_n414_));
  NOi21      g0392(.An(i_2_), .B(i_12_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n415_), .B(new_new_n414_), .Y(new_new_n416_));
  INV        g0394(.A(new_new_n416_), .Y(new_new_n417_));
  NA2        g0395(.A(new_new_n141_), .B(i_9_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n418_), .B(i_4_), .Y(new_new_n419_));
  NA2        g0397(.A(new_new_n417_), .B(new_new_n419_), .Y(new_new_n420_));
  OR2        g0398(.A(i_13_), .B(i_10_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n172_), .B(new_new_n122_), .Y(new_new_n422_));
  OR2        g0400(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n99_), .B(new_new_n25_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n286_), .B(new_new_n424_), .Y(new_new_n425_));
  INV        g0403(.A(new_new_n210_), .Y(new_new_n426_));
  OAI220     g0404(.A0(new_new_n426_), .A1(new_new_n423_), .B0(new_new_n425_), .B1(new_new_n101_), .Y(new_new_n427_));
  INV        g0405(.A(new_new_n427_), .Y(new_new_n428_));
  AOI210     g0406(.A0(new_new_n428_), .A1(new_new_n420_), .B0(new_new_n26_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n326_), .B(new_new_n325_), .Y(new_new_n430_));
  AOI220     g0408(.A0(new_new_n299_), .A1(new_new_n290_), .B0(new_new_n293_), .B1(new_new_n317_), .Y(new_new_n431_));
  NO2        g0409(.A(new_new_n431_), .B(i_5_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n181_), .B(new_new_n82_), .Y(new_new_n433_));
  AOI220     g0411(.A0(new_new_n433_), .A1(new_new_n298_), .B0(i_6_), .B1(new_new_n210_), .Y(new_new_n434_));
  NO2        g0412(.A(new_new_n434_), .B(new_new_n288_), .Y(new_new_n435_));
  NO3        g0413(.A(new_new_n435_), .B(new_new_n432_), .C(new_new_n430_), .Y(new_new_n436_));
  NA2        g0414(.A(new_new_n195_), .B(new_new_n94_), .Y(new_new_n437_));
  NA3        g0415(.A(new_new_n329_), .B(new_new_n163_), .C(new_new_n82_), .Y(new_new_n438_));
  AOI210     g0416(.A0(new_new_n438_), .A1(new_new_n437_), .B0(new_new_n327_), .Y(new_new_n439_));
  NA3        g0417(.A(new_new_n258_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n440_));
  NA2        g0418(.A(new_new_n299_), .B(new_new_n236_), .Y(new_new_n441_));
  OAI220     g0419(.A0(new_new_n441_), .A1(new_new_n181_), .B0(new_new_n440_), .B1(new_new_n1043_), .Y(new_new_n442_));
  NO2        g0420(.A(i_3_), .B(new_new_n48_), .Y(new_new_n443_));
  NA3        g0421(.A(new_new_n342_), .B(new_new_n341_), .C(new_new_n443_), .Y(new_new_n444_));
  NA2        g0422(.A(new_new_n319_), .B(new_new_n324_), .Y(new_new_n445_));
  OAI210     g0423(.A0(new_new_n445_), .A1(new_new_n188_), .B0(new_new_n444_), .Y(new_new_n446_));
  NO3        g0424(.A(new_new_n446_), .B(new_new_n442_), .C(new_new_n439_), .Y(new_new_n447_));
  AOI210     g0425(.A0(new_new_n447_), .A1(new_new_n436_), .B0(new_new_n275_), .Y(new_new_n448_));
  NO4        g0426(.A(new_new_n448_), .B(new_new_n429_), .C(new_new_n411_), .D(new_new_n384_), .Y(new_new_n449_));
  NO2        g0427(.A(new_new_n63_), .B(i_4_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n70_), .B(i_13_), .Y(new_new_n451_));
  NO2        g0429(.A(i_10_), .B(i_9_), .Y(new_new_n452_));
  NAi21      g0430(.An(i_12_), .B(i_8_), .Y(new_new_n453_));
  NO2        g0431(.A(new_new_n453_), .B(i_3_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n46_), .B(i_4_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n455_), .B(new_new_n102_), .Y(new_new_n456_));
  NO2        g0434(.A(new_new_n456_), .B(new_new_n204_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n312_), .B(i_0_), .Y(new_new_n458_));
  NO3        g0436(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n270_), .B(new_new_n95_), .Y(new_new_n460_));
  NA2        g0438(.A(new_new_n460_), .B(new_new_n459_), .Y(new_new_n461_));
  NA2        g0439(.A(i_8_), .B(i_9_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n461_), .B(new_new_n458_), .Y(new_new_n463_));
  NO3        g0441(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n464_));
  NA3        g0442(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n465_));
  NO2        g0443(.A(new_new_n463_), .B(new_new_n457_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n298_), .B(new_new_n106_), .Y(new_new_n467_));
  OA220      g0445(.A0(new_new_n355_), .A1(new_new_n162_), .B0(new_new_n467_), .B1(new_new_n233_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n94_), .B(i_13_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n433_), .B(new_new_n385_), .Y(new_new_n470_));
  NO2        g0448(.A(i_2_), .B(i_13_), .Y(new_new_n471_));
  NA3        g0449(.A(new_new_n471_), .B(new_new_n161_), .C(new_new_n97_), .Y(new_new_n472_));
  OAI220     g0450(.A0(new_new_n472_), .A1(new_new_n238_), .B0(new_new_n470_), .B1(new_new_n469_), .Y(new_new_n473_));
  NO3        g0451(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n474_));
  NO2        g0452(.A(i_6_), .B(i_7_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n475_), .B(new_new_n474_), .Y(new_new_n476_));
  NO2        g0454(.A(i_11_), .B(i_1_), .Y(new_new_n477_));
  OR2        g0455(.A(i_11_), .B(i_8_), .Y(new_new_n478_));
  NOi21      g0456(.An(i_2_), .B(i_7_), .Y(new_new_n479_));
  NAi31      g0457(.An(new_new_n478_), .B(new_new_n479_), .C(i_0_), .Y(new_new_n480_));
  NO2        g0458(.A(new_new_n421_), .B(i_6_), .Y(new_new_n481_));
  NA3        g0459(.A(new_new_n481_), .B(new_new_n450_), .C(new_new_n72_), .Y(new_new_n482_));
  NO2        g0460(.A(new_new_n482_), .B(new_new_n480_), .Y(new_new_n483_));
  NO2        g0461(.A(i_3_), .B(new_new_n192_), .Y(new_new_n484_));
  NO2        g0462(.A(i_6_), .B(i_10_), .Y(new_new_n485_));
  NA4        g0463(.A(new_new_n485_), .B(new_new_n316_), .C(new_new_n484_), .D(new_new_n238_), .Y(new_new_n486_));
  NO2        g0464(.A(new_new_n486_), .B(new_new_n155_), .Y(new_new_n487_));
  NA3        g0465(.A(new_new_n246_), .B(new_new_n171_), .C(new_new_n131_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n489_));
  NO2        g0467(.A(new_new_n157_), .B(i_3_), .Y(new_new_n490_));
  NAi31      g0468(.An(new_new_n489_), .B(new_new_n490_), .C(new_new_n227_), .Y(new_new_n491_));
  NA3        g0469(.A(new_new_n397_), .B(new_new_n178_), .C(new_new_n148_), .Y(new_new_n492_));
  NA3        g0470(.A(new_new_n492_), .B(new_new_n491_), .C(new_new_n488_), .Y(new_new_n493_));
  NO4        g0471(.A(new_new_n493_), .B(new_new_n487_), .C(new_new_n483_), .D(new_new_n473_), .Y(new_new_n494_));
  NA2        g0472(.A(new_new_n459_), .B(new_new_n386_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n464_), .B(new_new_n393_), .Y(new_new_n496_));
  NO2        g0474(.A(new_new_n496_), .B(new_new_n225_), .Y(new_new_n497_));
  NAi21      g0475(.An(new_new_n216_), .B(new_new_n402_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n342_), .B(new_new_n218_), .Y(new_new_n499_));
  NO2        g0477(.A(new_new_n26_), .B(i_5_), .Y(new_new_n500_));
  NO2        g0478(.A(i_0_), .B(new_new_n82_), .Y(new_new_n501_));
  NA3        g0479(.A(new_new_n501_), .B(new_new_n500_), .C(new_new_n141_), .Y(new_new_n502_));
  OAI220     g0480(.A0(new_new_n38_), .A1(new_new_n502_), .B0(new_new_n499_), .B1(new_new_n498_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n316_), .B(new_new_n240_), .Y(new_new_n504_));
  NO2        g0482(.A(new_new_n504_), .B(new_new_n440_), .Y(new_new_n505_));
  NA4        g0483(.A(new_new_n309_), .B(new_new_n224_), .C(new_new_n70_), .D(new_new_n238_), .Y(new_new_n506_));
  NO2        g0484(.A(new_new_n506_), .B(new_new_n476_), .Y(new_new_n507_));
  NO4        g0485(.A(new_new_n507_), .B(new_new_n505_), .C(new_new_n503_), .D(new_new_n497_), .Y(new_new_n508_));
  NA4        g0486(.A(new_new_n508_), .B(new_new_n494_), .C(new_new_n468_), .D(new_new_n466_), .Y(new_new_n509_));
  NA3        g0487(.A(new_new_n309_), .B(new_new_n175_), .C(new_new_n173_), .Y(new_new_n510_));
  OAI210     g0488(.A0(new_new_n304_), .A1(new_new_n179_), .B0(new_new_n510_), .Y(new_new_n511_));
  AN2        g0489(.A(new_new_n290_), .B(new_new_n235_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n512_), .B(new_new_n511_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n121_), .B(new_new_n110_), .Y(new_new_n514_));
  AN2        g0492(.A(new_new_n514_), .B(new_new_n459_), .Y(new_new_n515_));
  OAI210     g0493(.A0(i_2_), .A1(new_new_n233_), .B0(new_new_n310_), .Y(new_new_n516_));
  AOI220     g0494(.A0(new_new_n516_), .A1(new_new_n328_), .B0(new_new_n515_), .B1(new_new_n312_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n386_), .B(new_new_n226_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n359_), .B(new_new_n70_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n376_), .B(new_new_n369_), .Y(new_new_n520_));
  AO210      g0498(.A0(new_new_n519_), .A1(new_new_n518_), .B0(new_new_n520_), .Y(new_new_n521_));
  NO2        g0499(.A(new_new_n36_), .B(i_8_), .Y(new_new_n522_));
  INV        g0500(.A(new_new_n521_), .Y(new_new_n523_));
  OAI210     g0501(.A0(i_8_), .A1(new_new_n63_), .B0(new_new_n133_), .Y(new_new_n524_));
  AOI210     g0502(.A0(new_new_n193_), .A1(i_9_), .B0(new_new_n269_), .Y(new_new_n525_));
  NO2        g0503(.A(new_new_n525_), .B(new_new_n198_), .Y(new_new_n526_));
  AOI220     g0504(.A0(i_6_), .A1(new_new_n526_), .B0(new_new_n524_), .B1(new_new_n422_), .Y(new_new_n527_));
  NA4        g0505(.A(new_new_n527_), .B(new_new_n521_), .C(new_new_n517_), .D(new_new_n513_), .Y(new_new_n528_));
  NA2        g0506(.A(new_new_n392_), .B(new_new_n298_), .Y(new_new_n529_));
  NA2        g0507(.A(new_new_n169_), .B(new_new_n529_), .Y(new_new_n530_));
  NO2        g0508(.A(i_12_), .B(new_new_n192_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n531_), .B(new_new_n226_), .Y(new_new_n532_));
  NO3        g0510(.A(i_10_), .B(new_new_n532_), .C(new_new_n467_), .Y(new_new_n533_));
  NOi31      g0511(.An(new_new_n319_), .B(new_new_n421_), .C(new_new_n38_), .Y(new_new_n534_));
  OAI210     g0512(.A0(new_new_n534_), .A1(new_new_n533_), .B0(new_new_n530_), .Y(new_new_n535_));
  NO2        g0513(.A(i_8_), .B(i_7_), .Y(new_new_n536_));
  OAI210     g0514(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n537_), .B(new_new_n224_), .Y(new_new_n538_));
  AOI220     g0516(.A0(new_new_n329_), .A1(new_new_n39_), .B0(new_new_n236_), .B1(new_new_n207_), .Y(new_new_n539_));
  OAI220     g0517(.A0(new_new_n539_), .A1(new_new_n181_), .B0(new_new_n538_), .B1(new_new_n244_), .Y(new_new_n540_));
  NA2        g0518(.A(new_new_n44_), .B(i_10_), .Y(new_new_n541_));
  NO2        g0519(.A(new_new_n541_), .B(i_6_), .Y(new_new_n542_));
  NA3        g0520(.A(new_new_n542_), .B(new_new_n540_), .C(new_new_n536_), .Y(new_new_n543_));
  AOI220     g0521(.A0(new_new_n433_), .A1(new_new_n329_), .B0(new_new_n248_), .B1(new_new_n245_), .Y(new_new_n544_));
  OAI220     g0522(.A0(new_new_n544_), .A1(new_new_n266_), .B0(new_new_n469_), .B1(new_new_n132_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n545_), .B(new_new_n269_), .Y(new_new_n546_));
  NOi31      g0524(.An(new_new_n293_), .B(new_new_n304_), .C(new_new_n179_), .Y(new_new_n547_));
  NA3        g0525(.A(new_new_n309_), .B(new_new_n173_), .C(new_new_n94_), .Y(new_new_n548_));
  NO2        g0526(.A(new_new_n157_), .B(i_5_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n549_), .B(new_new_n322_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n550_), .B(new_new_n548_), .Y(new_new_n551_));
  OAI210     g0529(.A0(new_new_n551_), .A1(new_new_n547_), .B0(new_new_n464_), .Y(new_new_n552_));
  NA4        g0530(.A(new_new_n552_), .B(new_new_n546_), .C(new_new_n543_), .D(new_new_n535_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n286_), .B(new_new_n81_), .Y(new_new_n554_));
  NO2        g0532(.A(new_new_n350_), .B(new_new_n554_), .Y(new_new_n555_));
  NA2        g0533(.A(new_new_n299_), .B(new_new_n290_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n556_), .B(new_new_n172_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n558_));
  NA2        g0536(.A(new_new_n452_), .B(new_new_n222_), .Y(new_new_n559_));
  NO2        g0537(.A(new_new_n558_), .B(new_new_n559_), .Y(new_new_n560_));
  NA3        g0538(.A(new_new_n531_), .B(new_new_n278_), .C(i_5_), .Y(new_new_n561_));
  NO2        g0539(.A(i_1_), .B(new_new_n561_), .Y(new_new_n562_));
  NO4        g0540(.A(new_new_n562_), .B(new_new_n560_), .C(new_new_n557_), .D(new_new_n555_), .Y(new_new_n563_));
  NO4        g0541(.A(new_new_n253_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n564_));
  NO3        g0542(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n234_), .B(new_new_n36_), .Y(new_new_n566_));
  AN2        g0544(.A(new_new_n566_), .B(new_new_n565_), .Y(new_new_n567_));
  AN2        g0545(.A(new_new_n567_), .B(new_new_n359_), .Y(new_new_n568_));
  NO2        g0546(.A(new_new_n421_), .B(i_1_), .Y(new_new_n569_));
  NOi31      g0547(.An(new_new_n569_), .B(new_new_n460_), .C(new_new_n70_), .Y(new_new_n570_));
  AN3        g0548(.A(new_new_n570_), .B(new_new_n419_), .C(new_new_n500_), .Y(new_new_n571_));
  NO2        g0549(.A(new_new_n431_), .B(new_new_n176_), .Y(new_new_n572_));
  NO3        g0550(.A(new_new_n572_), .B(new_new_n571_), .C(new_new_n568_), .Y(new_new_n573_));
  NOi21      g0551(.An(i_10_), .B(i_6_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n82_), .B(new_new_n25_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n113_), .B(new_new_n23_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n319_), .B(new_new_n164_), .Y(new_new_n577_));
  AOI220     g0555(.A0(new_new_n577_), .A1(new_new_n441_), .B0(new_new_n182_), .B1(new_new_n180_), .Y(new_new_n578_));
  NOi21      g0556(.An(new_new_n145_), .B(new_new_n337_), .Y(new_new_n579_));
  NO2        g0557(.A(new_new_n579_), .B(new_new_n578_), .Y(new_new_n580_));
  NO2        g0558(.A(new_new_n519_), .B(new_new_n382_), .Y(new_new_n581_));
  INV        g0559(.A(new_new_n322_), .Y(new_new_n582_));
  NO2        g0560(.A(i_12_), .B(new_new_n82_), .Y(new_new_n583_));
  NA3        g0561(.A(new_new_n583_), .B(new_new_n278_), .C(i_5_), .Y(new_new_n584_));
  NA3        g0562(.A(new_new_n389_), .B(new_new_n286_), .C(new_new_n218_), .Y(new_new_n585_));
  AOI210     g0563(.A0(new_new_n585_), .A1(new_new_n584_), .B0(new_new_n582_), .Y(new_new_n586_));
  NA2        g0564(.A(new_new_n173_), .B(i_0_), .Y(new_new_n587_));
  NO3        g0565(.A(new_new_n587_), .B(new_new_n1042_), .C(new_new_n304_), .Y(new_new_n588_));
  OR2        g0566(.A(i_2_), .B(i_5_), .Y(new_new_n589_));
  OR2        g0567(.A(new_new_n589_), .B(new_new_n414_), .Y(new_new_n590_));
  AOI210     g0568(.A0(new_new_n378_), .A1(new_new_n245_), .B0(new_new_n197_), .Y(new_new_n591_));
  AOI210     g0569(.A0(new_new_n591_), .A1(new_new_n590_), .B0(new_new_n498_), .Y(new_new_n592_));
  NO4        g0570(.A(new_new_n592_), .B(new_new_n588_), .C(new_new_n586_), .D(new_new_n581_), .Y(new_new_n593_));
  NA4        g0571(.A(new_new_n593_), .B(new_new_n580_), .C(new_new_n573_), .D(new_new_n563_), .Y(new_new_n594_));
  NO4        g0572(.A(new_new_n594_), .B(new_new_n553_), .C(new_new_n528_), .D(new_new_n509_), .Y(new_new_n595_));
  NA4        g0573(.A(new_new_n595_), .B(new_new_n449_), .C(new_new_n358_), .D(new_new_n315_), .Y(men7));
  NO2        g0574(.A(new_new_n90_), .B(new_new_n54_), .Y(new_new_n597_));
  NO2        g0575(.A(new_new_n106_), .B(new_new_n87_), .Y(new_new_n598_));
  NA2        g0576(.A(new_new_n387_), .B(new_new_n598_), .Y(new_new_n599_));
  NA2        g0577(.A(new_new_n485_), .B(new_new_n81_), .Y(new_new_n600_));
  NA2        g0578(.A(i_11_), .B(new_new_n192_), .Y(new_new_n601_));
  NA2        g0579(.A(new_new_n143_), .B(new_new_n601_), .Y(new_new_n602_));
  OAI210     g0580(.A0(new_new_n602_), .A1(new_new_n600_), .B0(new_new_n599_), .Y(new_new_n603_));
  NA3        g0581(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n238_), .B(i_4_), .Y(new_new_n605_));
  NA2        g0583(.A(i_2_), .B(new_new_n82_), .Y(new_new_n606_));
  OAI210     g0584(.A0(new_new_n85_), .A1(new_new_n202_), .B0(new_new_n203_), .Y(new_new_n607_));
  NO2        g0585(.A(i_7_), .B(new_new_n37_), .Y(new_new_n608_));
  NA2        g0586(.A(i_4_), .B(i_8_), .Y(new_new_n609_));
  AOI210     g0587(.A0(new_new_n609_), .A1(new_new_n309_), .B0(new_new_n608_), .Y(new_new_n610_));
  OAI220     g0588(.A0(new_new_n610_), .A1(new_new_n606_), .B0(new_new_n607_), .B1(i_13_), .Y(new_new_n611_));
  NO3        g0589(.A(new_new_n611_), .B(new_new_n603_), .C(new_new_n597_), .Y(new_new_n612_));
  INV        g0590(.A(new_new_n161_), .Y(new_new_n613_));
  OR2        g0591(.A(i_6_), .B(i_10_), .Y(new_new_n614_));
  NO2        g0592(.A(new_new_n614_), .B(new_new_n23_), .Y(new_new_n615_));
  OR3        g0593(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n616_));
  NO3        g0594(.A(new_new_n616_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n617_));
  INV        g0595(.A(new_new_n199_), .Y(new_new_n618_));
  NO2        g0596(.A(new_new_n617_), .B(new_new_n615_), .Y(new_new_n619_));
  OA220      g0597(.A0(new_new_n619_), .A1(new_new_n582_), .B0(new_new_n613_), .B1(new_new_n271_), .Y(new_new_n620_));
  AOI210     g0598(.A0(new_new_n620_), .A1(new_new_n612_), .B0(new_new_n63_), .Y(new_new_n621_));
  NOi21      g0599(.An(i_11_), .B(i_7_), .Y(new_new_n622_));
  AO210      g0600(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n623_));
  NO2        g0601(.A(new_new_n623_), .B(new_new_n622_), .Y(new_new_n624_));
  NA3        g0602(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n625_));
  NAi21      g0603(.An(new_new_n625_), .B(i_11_), .Y(new_new_n626_));
  NO2        g0604(.A(new_new_n626_), .B(new_new_n63_), .Y(new_new_n627_));
  NA2        g0605(.A(new_new_n84_), .B(new_new_n63_), .Y(new_new_n628_));
  AO210      g0606(.A0(new_new_n628_), .A1(new_new_n382_), .B0(new_new_n40_), .Y(new_new_n629_));
  NA2        g0607(.A(new_new_n227_), .B(new_new_n63_), .Y(new_new_n630_));
  NA2        g0608(.A(new_new_n415_), .B(new_new_n31_), .Y(new_new_n631_));
  OR2        g0609(.A(new_new_n208_), .B(new_new_n106_), .Y(new_new_n632_));
  NA2        g0610(.A(new_new_n632_), .B(new_new_n631_), .Y(new_new_n633_));
  NO2        g0611(.A(new_new_n63_), .B(i_9_), .Y(new_new_n634_));
  NA2        g0612(.A(new_new_n63_), .B(new_new_n633_), .Y(new_new_n635_));
  NO2        g0613(.A(i_1_), .B(i_12_), .Y(new_new_n636_));
  NA3        g0614(.A(new_new_n635_), .B(new_new_n630_), .C(new_new_n629_), .Y(new_new_n637_));
  OAI210     g0615(.A0(new_new_n637_), .A1(new_new_n627_), .B0(i_6_), .Y(new_new_n638_));
  NO2        g0616(.A(i_6_), .B(i_11_), .Y(new_new_n639_));
  INV        g0617(.A(new_new_n461_), .Y(new_new_n640_));
  NO4        g0618(.A(new_new_n215_), .B(new_new_n127_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n641_));
  NA2        g0619(.A(new_new_n641_), .B(new_new_n634_), .Y(new_new_n642_));
  NO3        g0620(.A(new_new_n614_), .B(new_new_n234_), .C(new_new_n23_), .Y(new_new_n643_));
  AOI210     g0621(.A0(i_1_), .A1(new_new_n261_), .B0(new_new_n643_), .Y(new_new_n644_));
  OAI210     g0622(.A0(new_new_n644_), .A1(new_new_n44_), .B0(new_new_n642_), .Y(new_new_n645_));
  NA3        g0623(.A(new_new_n536_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n646_));
  NA2        g0624(.A(new_new_n137_), .B(i_9_), .Y(new_new_n647_));
  NA3        g0625(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n46_), .B(i_1_), .Y(new_new_n649_));
  NA3        g0627(.A(new_new_n649_), .B(new_new_n270_), .C(new_new_n44_), .Y(new_new_n650_));
  OAI220     g0628(.A0(new_new_n650_), .A1(new_new_n648_), .B0(new_new_n647_), .B1(new_new_n1039_), .Y(new_new_n651_));
  NA3        g0629(.A(new_new_n634_), .B(new_new_n322_), .C(i_6_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n652_), .B(new_new_n23_), .Y(new_new_n653_));
  AOI210     g0631(.A0(new_new_n477_), .A1(new_new_n424_), .B0(new_new_n243_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n654_), .B(new_new_n606_), .Y(new_new_n655_));
  NAi21      g0633(.An(new_new_n646_), .B(new_new_n89_), .Y(new_new_n656_));
  NA2        g0634(.A(new_new_n649_), .B(new_new_n270_), .Y(new_new_n657_));
  NO2        g0635(.A(i_11_), .B(new_new_n37_), .Y(new_new_n658_));
  NA2        g0636(.A(new_new_n658_), .B(new_new_n24_), .Y(new_new_n659_));
  OAI210     g0637(.A0(new_new_n659_), .A1(new_new_n657_), .B0(new_new_n656_), .Y(new_new_n660_));
  OR4        g0638(.A(new_new_n660_), .B(new_new_n655_), .C(new_new_n653_), .D(new_new_n651_), .Y(new_new_n661_));
  NO3        g0639(.A(new_new_n661_), .B(new_new_n645_), .C(new_new_n640_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n238_), .B(new_new_n99_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n663_), .B(new_new_n622_), .Y(new_new_n664_));
  NA2        g0642(.A(new_new_n664_), .B(i_1_), .Y(new_new_n665_));
  NO2        g0643(.A(new_new_n665_), .B(new_new_n616_), .Y(new_new_n666_));
  NA2        g0644(.A(new_new_n666_), .B(new_new_n46_), .Y(new_new_n667_));
  NA2        g0645(.A(i_3_), .B(new_new_n192_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n668_), .B(new_new_n113_), .Y(new_new_n669_));
  AN2        g0647(.A(new_new_n669_), .B(new_new_n542_), .Y(new_new_n670_));
  NO2        g0648(.A(new_new_n234_), .B(new_new_n44_), .Y(new_new_n671_));
  NO3        g0649(.A(new_new_n671_), .B(new_new_n312_), .C(new_new_n239_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n116_), .B(new_new_n37_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n673_), .B(i_6_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n82_), .B(i_9_), .Y(new_new_n675_));
  NO2        g0653(.A(new_new_n675_), .B(new_new_n63_), .Y(new_new_n676_));
  NO2        g0654(.A(new_new_n676_), .B(new_new_n636_), .Y(new_new_n677_));
  NO4        g0655(.A(new_new_n677_), .B(new_new_n674_), .C(new_new_n672_), .D(i_4_), .Y(new_new_n678_));
  NA2        g0656(.A(i_1_), .B(i_3_), .Y(new_new_n679_));
  NO2        g0657(.A(new_new_n462_), .B(new_new_n90_), .Y(new_new_n680_));
  AOI210     g0658(.A0(new_new_n671_), .A1(new_new_n574_), .B0(new_new_n680_), .Y(new_new_n681_));
  NO2        g0659(.A(new_new_n681_), .B(new_new_n679_), .Y(new_new_n682_));
  NO3        g0660(.A(new_new_n682_), .B(new_new_n678_), .C(new_new_n670_), .Y(new_new_n683_));
  NA4        g0661(.A(new_new_n683_), .B(new_new_n667_), .C(new_new_n662_), .D(new_new_n638_), .Y(new_new_n684_));
  NO3        g0662(.A(new_new_n478_), .B(i_3_), .C(i_7_), .Y(new_new_n685_));
  NOi21      g0663(.An(new_new_n685_), .B(i_10_), .Y(new_new_n686_));
  OA210      g0664(.A0(new_new_n686_), .A1(new_new_n246_), .B0(new_new_n82_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n688_));
  NA3        g0666(.A(new_new_n485_), .B(new_new_n522_), .C(new_new_n46_), .Y(new_new_n689_));
  NO3        g0667(.A(new_new_n479_), .B(new_new_n609_), .C(new_new_n82_), .Y(new_new_n690_));
  NA2        g0668(.A(new_new_n690_), .B(new_new_n25_), .Y(new_new_n691_));
  NA3        g0669(.A(new_new_n161_), .B(new_new_n81_), .C(new_new_n82_), .Y(new_new_n692_));
  NA4        g0670(.A(new_new_n692_), .B(new_new_n691_), .C(new_new_n689_), .D(new_new_n688_), .Y(new_new_n693_));
  OAI210     g0671(.A0(new_new_n693_), .A1(new_new_n687_), .B0(i_1_), .Y(new_new_n694_));
  AOI210     g0672(.A0(new_new_n270_), .A1(new_new_n95_), .B0(i_1_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n374_), .B(i_2_), .Y(new_new_n696_));
  NA2        g0674(.A(new_new_n696_), .B(new_new_n695_), .Y(new_new_n697_));
  OAI210     g0675(.A0(new_new_n652_), .A1(new_new_n453_), .B0(new_new_n697_), .Y(new_new_n698_));
  INV        g0676(.A(new_new_n698_), .Y(new_new_n699_));
  AOI210     g0677(.A0(new_new_n699_), .A1(new_new_n694_), .B0(i_13_), .Y(new_new_n700_));
  OR2        g0678(.A(i_11_), .B(i_7_), .Y(new_new_n701_));
  NA3        g0679(.A(new_new_n701_), .B(new_new_n104_), .C(new_new_n137_), .Y(new_new_n702_));
  AOI220     g0680(.A0(new_new_n471_), .A1(new_new_n161_), .B0(new_new_n455_), .B1(new_new_n137_), .Y(new_new_n703_));
  OAI210     g0681(.A0(new_new_n703_), .A1(new_new_n44_), .B0(new_new_n702_), .Y(new_new_n704_));
  NA2        g0682(.A(new_new_n246_), .B(new_new_n130_), .Y(new_new_n705_));
  NO2        g0683(.A(new_new_n705_), .B(new_new_n40_), .Y(new_new_n706_));
  AOI210     g0684(.A0(new_new_n704_), .A1(new_new_n339_), .B0(new_new_n706_), .Y(new_new_n707_));
  AOI220     g0685(.A0(i_7_), .A1(new_new_n69_), .B0(new_new_n389_), .B1(new_new_n649_), .Y(new_new_n708_));
  NO2        g0686(.A(new_new_n708_), .B(new_new_n244_), .Y(new_new_n709_));
  AOI210     g0687(.A0(new_new_n453_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n710_));
  NA2        g0688(.A(new_new_n126_), .B(i_13_), .Y(new_new_n711_));
  NO2        g0689(.A(new_new_n648_), .B(new_new_n113_), .Y(new_new_n712_));
  INV        g0690(.A(new_new_n712_), .Y(new_new_n713_));
  OAI220     g0691(.A0(new_new_n713_), .A1(new_new_n68_), .B0(new_new_n711_), .B1(new_new_n695_), .Y(new_new_n714_));
  NO3        g0692(.A(new_new_n68_), .B(new_new_n32_), .C(new_new_n99_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n26_), .B(new_new_n192_), .Y(new_new_n716_));
  NA2        g0694(.A(new_new_n716_), .B(i_7_), .Y(new_new_n717_));
  NO3        g0695(.A(new_new_n479_), .B(new_new_n238_), .C(new_new_n82_), .Y(new_new_n718_));
  AOI210     g0696(.A0(new_new_n718_), .A1(new_new_n717_), .B0(new_new_n715_), .Y(new_new_n719_));
  NO2        g0697(.A(new_new_n719_), .B(new_new_n618_), .Y(new_new_n720_));
  NO3        g0698(.A(new_new_n720_), .B(new_new_n714_), .C(new_new_n709_), .Y(new_new_n721_));
  OR2        g0699(.A(i_11_), .B(i_6_), .Y(new_new_n722_));
  NA3        g0700(.A(new_new_n605_), .B(new_new_n716_), .C(i_7_), .Y(new_new_n723_));
  AOI210     g0701(.A0(new_new_n723_), .A1(new_new_n713_), .B0(new_new_n722_), .Y(new_new_n724_));
  NA2        g0702(.A(new_new_n639_), .B(i_13_), .Y(new_new_n725_));
  NAi21      g0703(.An(i_11_), .B(i_12_), .Y(new_new_n726_));
  NOi41      g0704(.An(new_new_n109_), .B(new_new_n726_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n727_));
  NO3        g0705(.A(new_new_n479_), .B(new_new_n583_), .C(new_new_n609_), .Y(new_new_n728_));
  AOI220     g0706(.A0(new_new_n728_), .A1(new_new_n316_), .B0(new_new_n727_), .B1(new_new_n192_), .Y(new_new_n729_));
  NA2        g0707(.A(new_new_n729_), .B(new_new_n725_), .Y(new_new_n730_));
  OAI210     g0708(.A0(new_new_n730_), .A1(new_new_n724_), .B0(new_new_n63_), .Y(new_new_n731_));
  NA2        g0709(.A(i_8_), .B(new_new_n25_), .Y(new_new_n732_));
  NO3        g0710(.A(new_new_n732_), .B(new_new_n387_), .C(new_new_n605_), .Y(new_new_n733_));
  OAI210     g0711(.A0(new_new_n733_), .A1(new_new_n375_), .B0(new_new_n373_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n127_), .B(i_2_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n735_), .B(new_new_n636_), .Y(new_new_n736_));
  NA2        g0714(.A(new_new_n736_), .B(new_new_n734_), .Y(new_new_n737_));
  NA3        g0715(.A(new_new_n737_), .B(new_new_n45_), .C(new_new_n226_), .Y(new_new_n738_));
  NA4        g0716(.A(new_new_n738_), .B(new_new_n731_), .C(new_new_n721_), .D(new_new_n707_), .Y(new_new_n739_));
  OR4        g0717(.A(new_new_n739_), .B(new_new_n700_), .C(new_new_n684_), .D(new_new_n621_), .Y(men5));
  AOI210     g0718(.A0(new_new_n664_), .A1(new_new_n273_), .B0(new_new_n422_), .Y(new_new_n741_));
  NO3        g0719(.A(i_11_), .B(new_new_n238_), .C(i_13_), .Y(new_new_n742_));
  NO2        g0720(.A(new_new_n123_), .B(new_new_n23_), .Y(new_new_n743_));
  NA2        g0721(.A(i_12_), .B(i_8_), .Y(new_new_n744_));
  OAI210     g0722(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n744_), .Y(new_new_n745_));
  INV        g0723(.A(new_new_n452_), .Y(new_new_n746_));
  AOI220     g0724(.A0(new_new_n322_), .A1(new_new_n576_), .B0(new_new_n745_), .B1(new_new_n743_), .Y(new_new_n747_));
  INV        g0725(.A(new_new_n747_), .Y(new_new_n748_));
  NO2        g0726(.A(new_new_n748_), .B(new_new_n1041_), .Y(new_new_n749_));
  INV        g0727(.A(new_new_n171_), .Y(new_new_n750_));
  INV        g0728(.A(new_new_n246_), .Y(new_new_n751_));
  OAI210     g0729(.A0(new_new_n696_), .A1(new_new_n454_), .B0(new_new_n109_), .Y(new_new_n752_));
  AOI210     g0730(.A0(new_new_n752_), .A1(new_new_n751_), .B0(new_new_n750_), .Y(new_new_n753_));
  NO2        g0731(.A(new_new_n462_), .B(new_new_n26_), .Y(new_new_n754_));
  NO2        g0732(.A(new_new_n754_), .B(new_new_n424_), .Y(new_new_n755_));
  NA2        g0733(.A(new_new_n755_), .B(i_2_), .Y(new_new_n756_));
  INV        g0734(.A(new_new_n756_), .Y(new_new_n757_));
  AOI210     g0735(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n421_), .Y(new_new_n758_));
  AOI210     g0736(.A0(new_new_n758_), .A1(new_new_n757_), .B0(new_new_n753_), .Y(new_new_n759_));
  NO2        g0737(.A(new_new_n189_), .B(new_new_n124_), .Y(new_new_n760_));
  OAI210     g0738(.A0(new_new_n760_), .A1(new_new_n743_), .B0(i_2_), .Y(new_new_n761_));
  NO2        g0739(.A(new_new_n761_), .B(new_new_n192_), .Y(new_new_n762_));
  OA210      g0740(.A0(new_new_n624_), .A1(new_new_n125_), .B0(i_13_), .Y(new_new_n763_));
  NA2        g0741(.A(new_new_n199_), .B(new_new_n202_), .Y(new_new_n764_));
  NA2        g0742(.A(new_new_n151_), .B(new_new_n601_), .Y(new_new_n765_));
  AOI210     g0743(.A0(new_new_n765_), .A1(new_new_n764_), .B0(new_new_n378_), .Y(new_new_n766_));
  AOI210     g0744(.A0(new_new_n208_), .A1(new_new_n147_), .B0(new_new_n522_), .Y(new_new_n767_));
  NA2        g0745(.A(new_new_n767_), .B(new_new_n424_), .Y(new_new_n768_));
  NO2        g0746(.A(new_new_n100_), .B(new_new_n44_), .Y(new_new_n769_));
  INV        g0747(.A(new_new_n305_), .Y(new_new_n770_));
  NA4        g0748(.A(new_new_n770_), .B(new_new_n309_), .C(new_new_n123_), .D(new_new_n42_), .Y(new_new_n771_));
  OAI210     g0749(.A0(new_new_n771_), .A1(new_new_n769_), .B0(new_new_n768_), .Y(new_new_n772_));
  NO4        g0750(.A(new_new_n772_), .B(new_new_n766_), .C(new_new_n763_), .D(new_new_n762_), .Y(new_new_n773_));
  NA2        g0751(.A(new_new_n576_), .B(new_new_n28_), .Y(new_new_n774_));
  NA2        g0752(.A(new_new_n742_), .B(new_new_n279_), .Y(new_new_n775_));
  NA2        g0753(.A(new_new_n775_), .B(new_new_n774_), .Y(new_new_n776_));
  NO2        g0754(.A(new_new_n62_), .B(i_12_), .Y(new_new_n777_));
  NO2        g0755(.A(new_new_n777_), .B(new_new_n125_), .Y(new_new_n778_));
  NO2        g0756(.A(new_new_n778_), .B(new_new_n601_), .Y(new_new_n779_));
  AOI220     g0757(.A0(new_new_n779_), .A1(new_new_n36_), .B0(new_new_n776_), .B1(new_new_n46_), .Y(new_new_n780_));
  NA4        g0758(.A(new_new_n780_), .B(new_new_n773_), .C(new_new_n759_), .D(new_new_n749_), .Y(men6));
  NA2        g0759(.A(new_new_n1044_), .B(new_new_n735_), .Y(new_new_n782_));
  NA4        g0760(.A(new_new_n393_), .B(new_new_n484_), .C(new_new_n68_), .D(new_new_n99_), .Y(new_new_n783_));
  INV        g0761(.A(new_new_n783_), .Y(new_new_n784_));
  NO2        g0762(.A(new_new_n221_), .B(new_new_n489_), .Y(new_new_n785_));
  NO2        g0763(.A(i_11_), .B(i_9_), .Y(new_new_n786_));
  NO2        g0764(.A(new_new_n784_), .B(new_new_n334_), .Y(new_new_n787_));
  AO210      g0765(.A0(new_new_n787_), .A1(new_new_n782_), .B0(i_12_), .Y(new_new_n788_));
  NA2        g0766(.A(new_new_n379_), .B(new_new_n342_), .Y(new_new_n789_));
  NA2        g0767(.A(new_new_n583_), .B(new_new_n63_), .Y(new_new_n790_));
  NA2        g0768(.A(new_new_n686_), .B(new_new_n68_), .Y(new_new_n791_));
  NA4        g0769(.A(new_new_n628_), .B(new_new_n791_), .C(new_new_n790_), .D(new_new_n789_), .Y(new_new_n792_));
  INV        g0770(.A(new_new_n196_), .Y(new_new_n793_));
  AOI220     g0771(.A0(new_new_n793_), .A1(new_new_n786_), .B0(new_new_n792_), .B1(new_new_n70_), .Y(new_new_n794_));
  INV        g0772(.A(new_new_n333_), .Y(new_new_n795_));
  NA2        g0773(.A(new_new_n72_), .B(new_new_n130_), .Y(new_new_n796_));
  NO2        g0774(.A(new_new_n796_), .B(new_new_n795_), .Y(new_new_n797_));
  NA2        g0775(.A(new_new_n1040_), .B(new_new_n777_), .Y(new_new_n798_));
  AOI210     g0776(.A0(new_new_n798_), .A1(new_new_n520_), .B0(new_new_n184_), .Y(new_new_n799_));
  INV        g0777(.A(i_11_), .Y(new_new_n800_));
  NA3        g0778(.A(new_new_n800_), .B(new_new_n475_), .C(new_new_n393_), .Y(new_new_n801_));
  NAi32      g0779(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n802_));
  AOI210     g0780(.A0(new_new_n722_), .A1(new_new_n83_), .B0(new_new_n802_), .Y(new_new_n803_));
  OAI210     g0781(.A0(new_new_n685_), .A1(new_new_n566_), .B0(new_new_n565_), .Y(new_new_n804_));
  NAi31      g0782(.An(new_new_n803_), .B(new_new_n804_), .C(new_new_n801_), .Y(new_new_n805_));
  OR3        g0783(.A(new_new_n805_), .B(new_new_n799_), .C(new_new_n797_), .Y(new_new_n806_));
  NA3        g0784(.A(new_new_n354_), .B(new_new_n257_), .C(i_7_), .Y(new_new_n807_));
  NA3        g0785(.A(new_new_n454_), .B(new_new_n146_), .C(new_new_n67_), .Y(new_new_n808_));
  OR2        g0786(.A(new_new_n746_), .B(new_new_n36_), .Y(new_new_n809_));
  NA3        g0787(.A(new_new_n809_), .B(new_new_n808_), .C(new_new_n807_), .Y(new_new_n810_));
  OAI210     g0788(.A0(i_6_), .A1(i_11_), .B0(new_new_n83_), .Y(new_new_n811_));
  AOI220     g0789(.A0(new_new_n811_), .A1(new_new_n565_), .B0(new_new_n785_), .B1(new_new_n717_), .Y(new_new_n812_));
  NA3        g0790(.A(new_new_n378_), .B(new_new_n240_), .C(new_new_n146_), .Y(new_new_n813_));
  NA3        g0791(.A(new_new_n813_), .B(new_new_n812_), .C(new_new_n607_), .Y(new_new_n814_));
  AO210      g0792(.A0(new_new_n522_), .A1(new_new_n46_), .B0(new_new_n84_), .Y(new_new_n815_));
  NA3        g0793(.A(new_new_n815_), .B(new_new_n485_), .C(new_new_n218_), .Y(new_new_n816_));
  INV        g0794(.A(new_new_n564_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n614_), .B(new_new_n100_), .Y(new_new_n818_));
  OAI210     g0796(.A0(new_new_n818_), .A1(new_new_n110_), .B0(new_new_n413_), .Y(new_new_n819_));
  INV        g0797(.A(new_new_n590_), .Y(new_new_n820_));
  NA3        g0798(.A(new_new_n820_), .B(new_new_n333_), .C(i_7_), .Y(new_new_n821_));
  NA4        g0799(.A(new_new_n821_), .B(new_new_n819_), .C(new_new_n817_), .D(new_new_n816_), .Y(new_new_n822_));
  NO4        g0800(.A(new_new_n822_), .B(new_new_n814_), .C(new_new_n810_), .D(new_new_n806_), .Y(new_new_n823_));
  NA4        g0801(.A(new_new_n823_), .B(new_new_n794_), .C(new_new_n788_), .D(new_new_n383_), .Y(men3));
  NA2        g0802(.A(i_12_), .B(i_10_), .Y(new_new_n825_));
  NA2        g0803(.A(i_6_), .B(i_7_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n826_), .B(i_0_), .Y(new_new_n827_));
  NO2        g0805(.A(i_11_), .B(new_new_n238_), .Y(new_new_n828_));
  OAI210     g0806(.A0(new_new_n827_), .A1(new_new_n293_), .B0(new_new_n828_), .Y(new_new_n829_));
  NO2        g0807(.A(new_new_n829_), .B(new_new_n192_), .Y(new_new_n830_));
  NO3        g0808(.A(new_new_n458_), .B(new_new_n87_), .C(new_new_n44_), .Y(new_new_n831_));
  OA210      g0809(.A0(new_new_n831_), .A1(new_new_n830_), .B0(new_new_n173_), .Y(new_new_n832_));
  NA3        g0810(.A(new_new_n813_), .B(new_new_n607_), .C(new_new_n377_), .Y(new_new_n833_));
  NA2        g0811(.A(new_new_n833_), .B(new_new_n39_), .Y(new_new_n834_));
  NO2        g0812(.A(new_new_n632_), .B(new_new_n462_), .Y(new_new_n835_));
  NA2        g0813(.A(new_new_n415_), .B(new_new_n45_), .Y(new_new_n836_));
  AN2        g0814(.A(new_new_n460_), .B(new_new_n55_), .Y(new_new_n837_));
  NO2        g0815(.A(new_new_n837_), .B(new_new_n835_), .Y(new_new_n838_));
  AOI210     g0816(.A0(new_new_n838_), .A1(new_new_n834_), .B0(new_new_n48_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n184_), .B(new_new_n574_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n710_), .B(new_new_n675_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n340_), .B(new_new_n443_), .Y(new_new_n842_));
  OAI220     g0820(.A0(new_new_n842_), .A1(new_new_n841_), .B0(new_new_n840_), .B1(new_new_n63_), .Y(new_new_n843_));
  NOi21      g0821(.An(i_5_), .B(i_9_), .Y(new_new_n844_));
  NA2        g0822(.A(new_new_n844_), .B(new_new_n451_), .Y(new_new_n845_));
  AOI210     g0823(.A0(new_new_n270_), .A1(new_new_n477_), .B0(new_new_n690_), .Y(new_new_n846_));
  NO2        g0824(.A(new_new_n174_), .B(new_new_n147_), .Y(new_new_n847_));
  NA2        g0825(.A(new_new_n847_), .B(new_new_n245_), .Y(new_new_n848_));
  OAI220     g0826(.A0(new_new_n848_), .A1(new_new_n179_), .B0(new_new_n846_), .B1(new_new_n845_), .Y(new_new_n849_));
  NO4        g0827(.A(new_new_n849_), .B(new_new_n843_), .C(new_new_n839_), .D(new_new_n832_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n184_), .B(new_new_n24_), .Y(new_new_n851_));
  NO2        g0829(.A(new_new_n673_), .B(new_new_n598_), .Y(new_new_n852_));
  NO2        g0830(.A(new_new_n852_), .B(new_new_n851_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n316_), .B(new_new_n128_), .Y(new_new_n854_));
  NAi21      g0832(.An(new_new_n162_), .B(new_new_n443_), .Y(new_new_n855_));
  NO2        g0833(.A(new_new_n854_), .B(new_new_n405_), .Y(new_new_n856_));
  NO2        g0834(.A(new_new_n856_), .B(new_new_n853_), .Y(new_new_n857_));
  NA2        g0835(.A(new_new_n575_), .B(i_0_), .Y(new_new_n858_));
  NO3        g0836(.A(new_new_n858_), .B(new_new_n388_), .C(new_new_n85_), .Y(new_new_n859_));
  NO4        g0837(.A(new_new_n589_), .B(new_new_n215_), .C(new_new_n421_), .D(new_new_n414_), .Y(new_new_n860_));
  AOI210     g0838(.A0(new_new_n860_), .A1(i_11_), .B0(new_new_n859_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n742_), .B(new_new_n334_), .Y(new_new_n862_));
  AOI210     g0840(.A0(new_new_n485_), .A1(new_new_n85_), .B0(new_new_n58_), .Y(new_new_n863_));
  OAI220     g0841(.A0(new_new_n863_), .A1(new_new_n862_), .B0(new_new_n659_), .B1(new_new_n538_), .Y(new_new_n864_));
  NA2        g0842(.A(i_0_), .B(i_10_), .Y(new_new_n865_));
  OAI210     g0843(.A0(new_new_n865_), .A1(new_new_n82_), .B0(new_new_n541_), .Y(new_new_n866_));
  NO4        g0844(.A(new_new_n113_), .B(new_new_n58_), .C(new_new_n668_), .D(i_5_), .Y(new_new_n867_));
  AN2        g0845(.A(new_new_n867_), .B(new_new_n866_), .Y(new_new_n868_));
  AOI220     g0846(.A0(new_new_n340_), .A1(new_new_n96_), .B0(new_new_n184_), .B1(new_new_n81_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n569_), .B(i_4_), .Y(new_new_n870_));
  NA2        g0848(.A(new_new_n187_), .B(new_new_n202_), .Y(new_new_n871_));
  OAI220     g0849(.A0(new_new_n871_), .A1(new_new_n862_), .B0(new_new_n870_), .B1(new_new_n869_), .Y(new_new_n872_));
  NO3        g0850(.A(new_new_n872_), .B(new_new_n868_), .C(new_new_n864_), .Y(new_new_n873_));
  NA3        g0851(.A(new_new_n873_), .B(new_new_n861_), .C(new_new_n857_), .Y(new_new_n874_));
  NO2        g0852(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n875_));
  NA2        g0853(.A(i_11_), .B(i_9_), .Y(new_new_n876_));
  NO3        g0854(.A(i_12_), .B(new_new_n876_), .C(new_new_n606_), .Y(new_new_n877_));
  AN2        g0855(.A(new_new_n877_), .B(new_new_n875_), .Y(new_new_n878_));
  NA2        g0856(.A(new_new_n397_), .B(new_new_n178_), .Y(new_new_n879_));
  NA2        g0857(.A(new_new_n879_), .B(new_new_n160_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n876_), .B(new_new_n70_), .Y(new_new_n881_));
  NO2        g0859(.A(new_new_n174_), .B(i_0_), .Y(new_new_n882_));
  INV        g0860(.A(new_new_n882_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n475_), .B(new_new_n232_), .Y(new_new_n884_));
  AOI210     g0862(.A0(new_new_n376_), .A1(new_new_n41_), .B0(new_new_n412_), .Y(new_new_n885_));
  OAI220     g0863(.A0(new_new_n885_), .A1(new_new_n845_), .B0(new_new_n884_), .B1(new_new_n883_), .Y(new_new_n886_));
  NO3        g0864(.A(new_new_n886_), .B(new_new_n880_), .C(new_new_n878_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n658_), .B(new_new_n120_), .Y(new_new_n888_));
  NO2        g0866(.A(i_6_), .B(new_new_n888_), .Y(new_new_n889_));
  AOI210     g0867(.A0(new_new_n453_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n890_));
  NA2        g0868(.A(new_new_n171_), .B(new_new_n101_), .Y(new_new_n891_));
  NOi32      g0869(.An(new_new_n890_), .Bn(new_new_n187_), .C(new_new_n891_), .Y(new_new_n892_));
  NA2        g0870(.A(new_new_n608_), .B(new_new_n334_), .Y(new_new_n893_));
  NO2        g0871(.A(new_new_n893_), .B(new_new_n836_), .Y(new_new_n894_));
  NO3        g0872(.A(new_new_n894_), .B(new_new_n892_), .C(new_new_n889_), .Y(new_new_n895_));
  NOi21      g0873(.An(i_7_), .B(i_5_), .Y(new_new_n896_));
  NOi31      g0874(.An(new_new_n896_), .B(i_0_), .C(new_new_n726_), .Y(new_new_n897_));
  NA3        g0875(.A(new_new_n897_), .B(new_new_n387_), .C(i_6_), .Y(new_new_n898_));
  OA210      g0876(.A0(new_new_n891_), .A1(new_new_n520_), .B0(new_new_n898_), .Y(new_new_n899_));
  NO3        g0877(.A(new_new_n408_), .B(new_new_n366_), .C(new_new_n362_), .Y(new_new_n900_));
  NO2        g0878(.A(new_new_n264_), .B(new_new_n323_), .Y(new_new_n901_));
  NO2        g0879(.A(new_new_n726_), .B(new_new_n259_), .Y(new_new_n902_));
  AOI210     g0880(.A0(new_new_n902_), .A1(new_new_n901_), .B0(new_new_n900_), .Y(new_new_n903_));
  NA4        g0881(.A(new_new_n903_), .B(new_new_n899_), .C(new_new_n895_), .D(new_new_n887_), .Y(new_new_n904_));
  NO2        g0882(.A(new_new_n851_), .B(new_new_n241_), .Y(new_new_n905_));
  AN2        g0883(.A(new_new_n339_), .B(new_new_n334_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n905_), .B(i_10_), .Y(new_new_n907_));
  NO2        g0885(.A(new_new_n825_), .B(new_new_n322_), .Y(new_new_n908_));
  OA210      g0886(.A0(new_new_n475_), .A1(new_new_n224_), .B0(new_new_n474_), .Y(new_new_n909_));
  NA2        g0887(.A(new_new_n908_), .B(new_new_n881_), .Y(new_new_n910_));
  NA3        g0888(.A(new_new_n474_), .B(new_new_n415_), .C(new_new_n45_), .Y(new_new_n911_));
  OAI210     g0889(.A0(new_new_n855_), .A1(i_6_), .B0(new_new_n911_), .Y(new_new_n912_));
  NA2        g0890(.A(new_new_n881_), .B(new_new_n309_), .Y(new_new_n913_));
  NA2        g0891(.A(new_new_n186_), .B(new_new_n913_), .Y(new_new_n914_));
  AOI220     g0892(.A0(new_new_n914_), .A1(new_new_n475_), .B0(new_new_n912_), .B1(new_new_n70_), .Y(new_new_n915_));
  NO2        g0893(.A(new_new_n72_), .B(new_new_n744_), .Y(new_new_n916_));
  AOI210     g0894(.A0(new_new_n173_), .A1(new_new_n598_), .B0(new_new_n916_), .Y(new_new_n917_));
  NO2        g0895(.A(new_new_n917_), .B(new_new_n47_), .Y(new_new_n918_));
  NO3        g0896(.A(new_new_n589_), .B(new_new_n361_), .C(new_new_n24_), .Y(new_new_n919_));
  INV        g0897(.A(new_new_n919_), .Y(new_new_n920_));
  NAi21      g0898(.An(i_9_), .B(i_5_), .Y(new_new_n921_));
  NO2        g0899(.A(new_new_n921_), .B(new_new_n408_), .Y(new_new_n922_));
  NO2        g0900(.A(new_new_n604_), .B(new_new_n103_), .Y(new_new_n923_));
  AOI220     g0901(.A0(new_new_n923_), .A1(i_0_), .B0(new_new_n922_), .B1(new_new_n624_), .Y(new_new_n924_));
  OAI220     g0902(.A0(new_new_n924_), .A1(new_new_n82_), .B0(new_new_n920_), .B1(new_new_n172_), .Y(new_new_n925_));
  NO3        g0903(.A(new_new_n925_), .B(new_new_n918_), .C(new_new_n523_), .Y(new_new_n926_));
  NA4        g0904(.A(new_new_n926_), .B(new_new_n915_), .C(new_new_n910_), .D(new_new_n907_), .Y(new_new_n927_));
  NO3        g0905(.A(new_new_n927_), .B(new_new_n904_), .C(new_new_n874_), .Y(new_new_n928_));
  NO2        g0906(.A(i_0_), .B(new_new_n726_), .Y(new_new_n929_));
  NA2        g0907(.A(new_new_n70_), .B(new_new_n44_), .Y(new_new_n930_));
  NA2        g0908(.A(new_new_n865_), .B(new_new_n930_), .Y(new_new_n931_));
  NO2        g0909(.A(i_5_), .B(new_new_n25_), .Y(new_new_n932_));
  AO220      g0910(.A0(new_new_n932_), .A1(new_new_n931_), .B0(new_new_n929_), .B1(new_new_n173_), .Y(new_new_n933_));
  AOI210     g0911(.A0(new_new_n790_), .A1(new_new_n688_), .B0(new_new_n891_), .Y(new_new_n934_));
  AOI210     g0912(.A0(new_new_n933_), .A1(new_new_n351_), .B0(new_new_n934_), .Y(new_new_n935_));
  NA2        g0913(.A(new_new_n735_), .B(new_new_n145_), .Y(new_new_n936_));
  INV        g0914(.A(new_new_n936_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n937_), .B(new_new_n675_), .Y(new_new_n938_));
  NO2        g0916(.A(new_new_n804_), .B(new_new_n408_), .Y(new_new_n939_));
  NA3        g0917(.A(new_new_n827_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n940_));
  NA2        g0918(.A(new_new_n828_), .B(i_9_), .Y(new_new_n941_));
  AOI210     g0919(.A0(new_new_n940_), .A1(new_new_n502_), .B0(new_new_n941_), .Y(new_new_n942_));
  OAI210     g0920(.A0(new_new_n245_), .A1(i_9_), .B0(new_new_n231_), .Y(new_new_n943_));
  AOI210     g0921(.A0(new_new_n943_), .A1(new_new_n858_), .B0(new_new_n153_), .Y(new_new_n944_));
  NO3        g0922(.A(new_new_n944_), .B(new_new_n942_), .C(new_new_n939_), .Y(new_new_n945_));
  NA3        g0923(.A(new_new_n945_), .B(new_new_n938_), .C(new_new_n935_), .Y(new_new_n946_));
  NA2        g0924(.A(new_new_n906_), .B(new_new_n378_), .Y(new_new_n947_));
  AOI210     g0925(.A0(new_new_n304_), .A1(new_new_n162_), .B0(new_new_n947_), .Y(new_new_n948_));
  NA3        g0926(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n949_));
  NA2        g0927(.A(i_5_), .B(new_new_n490_), .Y(new_new_n950_));
  AOI210     g0928(.A0(new_new_n949_), .A1(new_new_n162_), .B0(new_new_n950_), .Y(new_new_n951_));
  NO2        g0929(.A(new_new_n951_), .B(new_new_n948_), .Y(new_new_n952_));
  NO3        g0930(.A(new_new_n865_), .B(new_new_n844_), .C(new_new_n189_), .Y(new_new_n953_));
  AOI220     g0931(.A0(new_new_n953_), .A1(i_11_), .B0(new_new_n570_), .B1(new_new_n72_), .Y(new_new_n954_));
  NO3        g0932(.A(new_new_n209_), .B(new_new_n386_), .C(i_0_), .Y(new_new_n955_));
  OAI210     g0933(.A0(new_new_n955_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n956_));
  OAI220     g0934(.A0(new_new_n532_), .A1(new_new_n138_), .B0(i_12_), .B1(new_new_n618_), .Y(new_new_n957_));
  NA3        g0935(.A(new_new_n957_), .B(new_new_n400_), .C(i_0_), .Y(new_new_n958_));
  NA4        g0936(.A(new_new_n958_), .B(new_new_n956_), .C(new_new_n954_), .D(new_new_n952_), .Y(new_new_n959_));
  NO2        g0937(.A(new_new_n244_), .B(new_new_n90_), .Y(new_new_n960_));
  AOI210     g0938(.A0(new_new_n960_), .A1(new_new_n929_), .B0(new_new_n107_), .Y(new_new_n961_));
  AOI220     g0939(.A0(new_new_n896_), .A1(new_new_n490_), .B0(new_new_n827_), .B1(new_new_n163_), .Y(new_new_n962_));
  NA2        g0940(.A(new_new_n354_), .B(new_new_n175_), .Y(new_new_n963_));
  OA220      g0941(.A0(new_new_n963_), .A1(new_new_n962_), .B0(new_new_n961_), .B1(i_5_), .Y(new_new_n964_));
  AOI210     g0942(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n174_), .Y(new_new_n965_));
  NA2        g0943(.A(new_new_n965_), .B(new_new_n909_), .Y(new_new_n966_));
  NA3        g0944(.A(new_new_n495_), .B(new_new_n488_), .C(new_new_n472_), .Y(new_new_n967_));
  INV        g0945(.A(new_new_n967_), .Y(new_new_n968_));
  NA3        g0946(.A(new_new_n393_), .B(new_new_n171_), .C(new_new_n170_), .Y(new_new_n969_));
  NA3        g0947(.A(i_5_), .B(new_new_n293_), .C(new_new_n231_), .Y(new_new_n970_));
  NA2        g0948(.A(new_new_n970_), .B(new_new_n969_), .Y(new_new_n971_));
  NA3        g0949(.A(new_new_n393_), .B(new_new_n341_), .C(new_new_n222_), .Y(new_new_n972_));
  INV        g0950(.A(new_new_n972_), .Y(new_new_n973_));
  NOi31      g0951(.An(new_new_n392_), .B(new_new_n930_), .C(new_new_n241_), .Y(new_new_n974_));
  NO3        g0952(.A(new_new_n974_), .B(new_new_n973_), .C(new_new_n971_), .Y(new_new_n975_));
  NA4        g0953(.A(new_new_n975_), .B(new_new_n968_), .C(new_new_n966_), .D(new_new_n964_), .Y(new_new_n976_));
  NO2        g0954(.A(new_new_n82_), .B(i_5_), .Y(new_new_n977_));
  NA3        g0955(.A(new_new_n828_), .B(new_new_n108_), .C(new_new_n123_), .Y(new_new_n978_));
  INV        g0956(.A(new_new_n978_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n979_), .B(new_new_n977_), .Y(new_new_n980_));
  NA3        g0958(.A(new_new_n309_), .B(i_5_), .C(new_new_n192_), .Y(new_new_n981_));
  NO3        g0959(.A(new_new_n241_), .B(i_0_), .C(i_12_), .Y(new_new_n982_));
  AOI220     g0960(.A0(new_new_n982_), .A1(new_new_n243_), .B0(new_new_n784_), .B1(new_new_n175_), .Y(new_new_n983_));
  AN2        g0961(.A(new_new_n865_), .B(new_new_n153_), .Y(new_new_n984_));
  NO3        g0962(.A(new_new_n984_), .B(i_12_), .C(new_new_n646_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n985_), .B(new_new_n218_), .Y(new_new_n986_));
  NA3        g0964(.A(new_new_n96_), .B(new_new_n574_), .C(i_11_), .Y(new_new_n987_));
  NO2        g0965(.A(new_new_n987_), .B(new_new_n155_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n896_), .B(new_new_n471_), .Y(new_new_n989_));
  INV        g0967(.A(new_new_n64_), .Y(new_new_n990_));
  OAI220     g0968(.A0(new_new_n990_), .A1(new_new_n981_), .B0(new_new_n989_), .B1(new_new_n676_), .Y(new_new_n991_));
  AOI210     g0969(.A0(new_new_n991_), .A1(new_new_n882_), .B0(new_new_n988_), .Y(new_new_n992_));
  NA4        g0970(.A(new_new_n992_), .B(new_new_n986_), .C(new_new_n983_), .D(new_new_n980_), .Y(new_new_n993_));
  NO4        g0971(.A(new_new_n993_), .B(new_new_n976_), .C(new_new_n959_), .D(new_new_n946_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n890_), .B(new_new_n373_), .C(i_5_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n995_), .B(new_new_n613_), .Y(new_new_n996_));
  NA2        g0974(.A(new_new_n996_), .B(new_new_n207_), .Y(new_new_n997_));
  AN2        g0975(.A(new_new_n701_), .B(new_new_n374_), .Y(new_new_n998_));
  NA2        g0976(.A(new_new_n185_), .B(new_new_n187_), .Y(new_new_n999_));
  AO210      g0977(.A0(new_new_n998_), .A1(new_new_n33_), .B0(new_new_n999_), .Y(new_new_n1000_));
  OAI210     g0978(.A0(new_new_n617_), .A1(new_new_n615_), .B0(new_new_n322_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n1001_), .B(new_new_n1000_), .Y(new_new_n1002_));
  NO2        g0980(.A(new_new_n465_), .B(new_new_n270_), .Y(new_new_n1003_));
  NO4        g0981(.A(new_new_n234_), .B(new_new_n144_), .C(new_new_n679_), .D(new_new_n37_), .Y(new_new_n1004_));
  NO3        g0982(.A(new_new_n1004_), .B(new_new_n1003_), .C(new_new_n860_), .Y(new_new_n1005_));
  OAI210     g0983(.A0(new_new_n987_), .A1(new_new_n147_), .B0(new_new_n1005_), .Y(new_new_n1006_));
  AOI210     g0984(.A0(new_new_n1002_), .A1(new_new_n48_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  AOI210     g0985(.A0(new_new_n1007_), .A1(new_new_n997_), .B0(new_new_n70_), .Y(new_new_n1008_));
  INV        g0986(.A(new_new_n567_), .Y(new_new_n1009_));
  NO2        g0987(.A(new_new_n1009_), .B(new_new_n750_), .Y(new_new_n1010_));
  INV        g0988(.A(new_new_n73_), .Y(new_new_n1011_));
  AOI210     g0989(.A0(new_new_n965_), .A1(i_5_), .B0(new_new_n897_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n1012_), .A1(new_new_n1011_), .B0(new_new_n679_), .Y(new_new_n1013_));
  NA2        g0991(.A(i_8_), .B(new_new_n73_), .Y(new_new_n1014_));
  NO2        g0992(.A(new_new_n1014_), .B(new_new_n238_), .Y(new_new_n1015_));
  NA3        g0993(.A(new_new_n94_), .B(new_new_n311_), .C(new_new_n31_), .Y(new_new_n1016_));
  INV        g0994(.A(new_new_n1016_), .Y(new_new_n1017_));
  NO3        g0995(.A(new_new_n1017_), .B(new_new_n1015_), .C(new_new_n1013_), .Y(new_new_n1018_));
  OAI210     g0996(.A0(new_new_n272_), .A1(new_new_n158_), .B0(new_new_n85_), .Y(new_new_n1019_));
  NA3        g0997(.A(new_new_n754_), .B(new_new_n293_), .C(new_new_n77_), .Y(new_new_n1020_));
  AOI210     g0998(.A0(new_new_n1020_), .A1(new_new_n1019_), .B0(i_11_), .Y(new_new_n1021_));
  NA2        g0999(.A(new_new_n609_), .B(new_new_n215_), .Y(new_new_n1022_));
  OAI210     g1000(.A0(new_new_n1022_), .A1(new_new_n890_), .B0(new_new_n207_), .Y(new_new_n1023_));
  NA2        g1001(.A(new_new_n164_), .B(i_5_), .Y(new_new_n1024_));
  AOI210     g1002(.A0(new_new_n1023_), .A1(new_new_n764_), .B0(new_new_n1024_), .Y(new_new_n1025_));
  NO3        g1003(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1026_));
  OAI210     g1004(.A0(new_new_n901_), .A1(new_new_n311_), .B0(new_new_n1026_), .Y(new_new_n1027_));
  NO2        g1005(.A(new_new_n1027_), .B(new_new_n726_), .Y(new_new_n1028_));
  NO4        g1006(.A(new_new_n921_), .B(new_new_n478_), .C(new_new_n254_), .D(new_new_n253_), .Y(new_new_n1029_));
  NO2        g1007(.A(new_new_n1029_), .B(new_new_n564_), .Y(new_new_n1030_));
  INV        g1008(.A(new_new_n367_), .Y(new_new_n1031_));
  AOI210     g1009(.A0(new_new_n1031_), .A1(new_new_n1030_), .B0(new_new_n40_), .Y(new_new_n1032_));
  NO4        g1010(.A(new_new_n1032_), .B(new_new_n1028_), .C(new_new_n1025_), .D(new_new_n1021_), .Y(new_new_n1033_));
  OAI210     g1011(.A0(new_new_n1018_), .A1(i_4_), .B0(new_new_n1033_), .Y(new_new_n1034_));
  NO3        g1012(.A(new_new_n1034_), .B(new_new_n1010_), .C(new_new_n1008_), .Y(new_new_n1035_));
  NA4        g1013(.A(new_new_n1035_), .B(new_new_n994_), .C(new_new_n928_), .D(new_new_n850_), .Y(men4));
  INV        g1014(.A(i_2_), .Y(new_new_n1039_));
  INV        g1015(.A(i_9_), .Y(new_new_n1040_));
  INV        g1016(.A(new_new_n741_), .Y(new_new_n1041_));
  INV        g1017(.A(i_6_), .Y(new_new_n1042_));
  INV        g1018(.A(i_10_), .Y(new_new_n1043_));
  INV        g1019(.A(i_9_), .Y(new_new_n1044_));
endmodule


