//Benchmark atmr_misex3_1774_0.25

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1397_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  INV        o000(.A(d), .Y(ori_ori_n29_));
  NA3        o001(.A(e), .B(ori_ori_n29_), .C(b), .Y(ori_ori_n30_));
  NOi32      o002(.An(i), .Bn(o), .C(h), .Y(ori_ori_n31_));
  NA2        o003(.A(ori_ori_n31_), .B(m), .Y(ori_ori_n32_));
  NOi32      o004(.An(j), .Bn(o), .C(k), .Y(ori_ori_n33_));
  INV        o005(.A(i), .Y(ori_ori_n34_));
  AN2        o006(.A(h), .B(o), .Y(ori_ori_n35_));
  NAi21      o007(.An(n), .B(m), .Y(ori_ori_n36_));
  NOi32      o008(.An(k), .Bn(h), .C(l), .Y(ori_ori_n37_));
  NOi32      o009(.An(k), .Bn(h), .C(o), .Y(ori_ori_n38_));
  INV        o010(.A(ori_ori_n38_), .Y(ori_ori_n39_));
  NO2        o011(.A(ori_ori_n39_), .B(ori_ori_n36_), .Y(ori_ori_n40_));
  INV        o012(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  AOI210     o013(.A0(ori_ori_n41_), .A1(ori_ori_n32_), .B0(ori_ori_n30_), .Y(ori_ori_n42_));
  INV        o014(.A(c), .Y(ori_ori_n43_));
  INV        o015(.A(d), .Y(ori_ori_n44_));
  NAi21      o016(.An(i), .B(h), .Y(ori_ori_n45_));
  NAi31      o017(.An(e), .B(d), .C(b), .Y(ori_ori_n46_));
  NAi31      o018(.An(l), .B(m), .C(k), .Y(ori_ori_n47_));
  NAi41      o019(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n48_));
  INV        o020(.A(m), .Y(ori_ori_n49_));
  NOi21      o021(.An(k), .B(l), .Y(ori_ori_n50_));
  NA2        o022(.A(ori_ori_n50_), .B(ori_ori_n49_), .Y(ori_ori_n51_));
  AN4        o023(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n52_));
  NOi21      o024(.An(h), .B(f), .Y(ori_ori_n53_));
  NA2        o025(.A(ori_ori_n53_), .B(ori_ori_n52_), .Y(ori_ori_n54_));
  NAi32      o026(.An(m), .Bn(k), .C(j), .Y(ori_ori_n55_));
  NOi32      o027(.An(h), .Bn(o), .C(f), .Y(ori_ori_n56_));
  OR2        o028(.A(ori_ori_n54_), .B(ori_ori_n51_), .Y(ori_ori_n57_));
  INV        o029(.A(ori_ori_n57_), .Y(ori_ori_n58_));
  INV        o030(.A(n), .Y(ori_ori_n59_));
  NOi32      o031(.An(e), .Bn(b), .C(d), .Y(ori_ori_n60_));
  INV        o032(.A(ori_ori_n60_), .Y(ori_ori_n61_));
  INV        o033(.A(j), .Y(ori_ori_n62_));
  AN3        o034(.A(m), .B(k), .C(i), .Y(ori_ori_n63_));
  NA3        o035(.A(ori_ori_n63_), .B(ori_ori_n62_), .C(o), .Y(ori_ori_n64_));
  NO2        o036(.A(ori_ori_n64_), .B(f), .Y(ori_ori_n65_));
  NAi32      o037(.An(o), .Bn(f), .C(h), .Y(ori_ori_n66_));
  NAi31      o038(.An(j), .B(m), .C(l), .Y(ori_ori_n67_));
  NO2        o039(.A(ori_ori_n67_), .B(ori_ori_n66_), .Y(ori_ori_n68_));
  NA2        o040(.A(m), .B(l), .Y(ori_ori_n69_));
  NAi31      o041(.An(k), .B(j), .C(o), .Y(ori_ori_n70_));
  NO3        o042(.A(ori_ori_n70_), .B(ori_ori_n69_), .C(f), .Y(ori_ori_n71_));
  NAi41      o043(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n72_));
  AN2        o044(.A(e), .B(b), .Y(ori_ori_n73_));
  NOi31      o045(.An(c), .B(h), .C(f), .Y(ori_ori_n74_));
  NA2        o046(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  NO2        o047(.A(ori_ori_n75_), .B(ori_ori_n72_), .Y(ori_ori_n76_));
  NOi21      o048(.An(i), .B(h), .Y(ori_ori_n77_));
  INV        o049(.A(a), .Y(ori_ori_n78_));
  NA2        o050(.A(ori_ori_n73_), .B(ori_ori_n78_), .Y(ori_ori_n79_));
  INV        o051(.A(l), .Y(ori_ori_n80_));
  NOi21      o052(.An(m), .B(n), .Y(ori_ori_n81_));
  AN2        o053(.A(k), .B(h), .Y(ori_ori_n82_));
  INV        o054(.A(b), .Y(ori_ori_n83_));
  NA2        o055(.A(l), .B(j), .Y(ori_ori_n84_));
  AN2        o056(.A(k), .B(i), .Y(ori_ori_n85_));
  NA2        o057(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n86_));
  INV        o058(.A(ori_ori_n76_), .Y(ori_ori_n87_));
  OAI210     o059(.A0(ori_ori_n932_), .A1(ori_ori_n61_), .B0(ori_ori_n87_), .Y(ori_ori_n88_));
  NOi31      o060(.An(k), .B(m), .C(j), .Y(ori_ori_n89_));
  NA3        o061(.A(ori_ori_n89_), .B(ori_ori_n53_), .C(ori_ori_n52_), .Y(ori_ori_n90_));
  NOi31      o062(.An(k), .B(m), .C(i), .Y(ori_ori_n91_));
  INV        o063(.A(ori_ori_n90_), .Y(ori_ori_n92_));
  NOi32      o064(.An(f), .Bn(b), .C(e), .Y(ori_ori_n93_));
  NAi21      o065(.An(o), .B(h), .Y(ori_ori_n94_));
  NAi21      o066(.An(m), .B(n), .Y(ori_ori_n95_));
  NO3        o067(.A(j), .B(ori_ori_n95_), .C(ori_ori_n94_), .Y(ori_ori_n96_));
  NAi41      o068(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n97_));
  NAi31      o069(.An(j), .B(k), .C(h), .Y(ori_ori_n98_));
  NA2        o070(.A(ori_ori_n96_), .B(ori_ori_n93_), .Y(ori_ori_n99_));
  INV        o071(.A(ori_ori_n95_), .Y(ori_ori_n100_));
  AN2        o072(.A(k), .B(j), .Y(ori_ori_n101_));
  NAi21      o073(.An(c), .B(b), .Y(ori_ori_n102_));
  NA2        o074(.A(f), .B(d), .Y(ori_ori_n103_));
  NO4        o075(.A(ori_ori_n103_), .B(ori_ori_n102_), .C(ori_ori_n101_), .D(ori_ori_n94_), .Y(ori_ori_n104_));
  NA2        o076(.A(h), .B(c), .Y(ori_ori_n105_));
  NAi31      o077(.An(f), .B(e), .C(b), .Y(ori_ori_n106_));
  NA2        o078(.A(ori_ori_n104_), .B(ori_ori_n100_), .Y(ori_ori_n107_));
  NA2        o079(.A(d), .B(b), .Y(ori_ori_n108_));
  INV        o080(.A(ori_ori_n108_), .Y(ori_ori_n109_));
  NA2        o081(.A(b), .B(a), .Y(ori_ori_n110_));
  NAi21      o082(.An(e), .B(o), .Y(ori_ori_n111_));
  NAi21      o083(.An(c), .B(d), .Y(ori_ori_n112_));
  NAi31      o084(.An(l), .B(k), .C(h), .Y(ori_ori_n113_));
  NO2        o085(.A(ori_ori_n95_), .B(ori_ori_n113_), .Y(ori_ori_n114_));
  NA2        o086(.A(ori_ori_n114_), .B(ori_ori_n109_), .Y(ori_ori_n115_));
  NAi31      o087(.An(ori_ori_n92_), .B(ori_ori_n107_), .C(ori_ori_n99_), .Y(ori_ori_n116_));
  NAi31      o088(.An(e), .B(f), .C(b), .Y(ori_ori_n117_));
  INV        o089(.A(ori_ori_n117_), .Y(ori_ori_n118_));
  NOi21      o090(.An(h), .B(i), .Y(ori_ori_n119_));
  NOi21      o091(.An(k), .B(m), .Y(ori_ori_n120_));
  NA3        o092(.A(ori_ori_n120_), .B(ori_ori_n119_), .C(n), .Y(ori_ori_n121_));
  NOi21      o093(.An(ori_ori_n118_), .B(ori_ori_n121_), .Y(ori_ori_n122_));
  NOi21      o094(.An(h), .B(o), .Y(ori_ori_n123_));
  NAi31      o095(.An(d), .B(f), .C(c), .Y(ori_ori_n124_));
  NAi31      o096(.An(e), .B(f), .C(c), .Y(ori_ori_n125_));
  NA2        o097(.A(ori_ori_n125_), .B(ori_ori_n124_), .Y(ori_ori_n126_));
  NA2        o098(.A(j), .B(h), .Y(ori_ori_n127_));
  OR3        o099(.A(n), .B(m), .C(k), .Y(ori_ori_n128_));
  NO2        o100(.A(ori_ori_n128_), .B(ori_ori_n127_), .Y(ori_ori_n129_));
  NAi32      o101(.An(m), .Bn(k), .C(n), .Y(ori_ori_n130_));
  NO2        o102(.A(ori_ori_n130_), .B(ori_ori_n127_), .Y(ori_ori_n131_));
  AOI220     o103(.A0(ori_ori_n131_), .A1(ori_ori_n118_), .B0(ori_ori_n129_), .B1(ori_ori_n126_), .Y(ori_ori_n132_));
  NO2        o104(.A(n), .B(m), .Y(ori_ori_n133_));
  NA2        o105(.A(ori_ori_n133_), .B(ori_ori_n37_), .Y(ori_ori_n134_));
  NAi21      o106(.An(f), .B(e), .Y(ori_ori_n135_));
  NA2        o107(.A(d), .B(c), .Y(ori_ori_n136_));
  NO2        o108(.A(ori_ori_n136_), .B(ori_ori_n135_), .Y(ori_ori_n137_));
  NOi21      o109(.An(ori_ori_n137_), .B(ori_ori_n134_), .Y(ori_ori_n138_));
  NAi31      o110(.An(m), .B(n), .C(b), .Y(ori_ori_n139_));
  NA2        o111(.A(k), .B(i), .Y(ori_ori_n140_));
  NAi21      o112(.An(h), .B(f), .Y(ori_ori_n141_));
  NO2        o113(.A(ori_ori_n141_), .B(ori_ori_n140_), .Y(ori_ori_n142_));
  NO2        o114(.A(ori_ori_n139_), .B(ori_ori_n112_), .Y(ori_ori_n143_));
  NA2        o115(.A(ori_ori_n143_), .B(ori_ori_n142_), .Y(ori_ori_n144_));
  NOi32      o116(.An(f), .Bn(c), .C(d), .Y(ori_ori_n145_));
  NOi32      o117(.An(f), .Bn(c), .C(e), .Y(ori_ori_n146_));
  NO2        o118(.A(ori_ori_n146_), .B(ori_ori_n145_), .Y(ori_ori_n147_));
  NO3        o119(.A(n), .B(m), .C(j), .Y(ori_ori_n148_));
  NA2        o120(.A(ori_ori_n148_), .B(ori_ori_n82_), .Y(ori_ori_n149_));
  AO210      o121(.A0(ori_ori_n149_), .A1(ori_ori_n134_), .B0(ori_ori_n147_), .Y(ori_ori_n150_));
  NAi41      o122(.An(ori_ori_n138_), .B(ori_ori_n150_), .C(ori_ori_n144_), .D(ori_ori_n132_), .Y(ori_ori_n151_));
  OR3        o123(.A(ori_ori_n151_), .B(ori_ori_n122_), .C(ori_ori_n116_), .Y(ori_ori_n152_));
  NO4        o124(.A(ori_ori_n152_), .B(ori_ori_n88_), .C(ori_ori_n58_), .D(ori_ori_n42_), .Y(ori_ori_n153_));
  INV        o125(.A(m), .Y(ori_ori_n154_));
  NAi31      o126(.An(n), .B(h), .C(o), .Y(ori_ori_n155_));
  NO2        o127(.A(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NOi32      o128(.An(m), .Bn(k), .C(l), .Y(ori_ori_n157_));
  NA3        o129(.A(ori_ori_n157_), .B(ori_ori_n62_), .C(o), .Y(ori_ori_n158_));
  NO2        o130(.A(ori_ori_n158_), .B(n), .Y(ori_ori_n159_));
  NOi21      o131(.An(k), .B(j), .Y(ori_ori_n160_));
  NA4        o132(.A(ori_ori_n160_), .B(ori_ori_n81_), .C(i), .D(o), .Y(ori_ori_n161_));
  INV        o133(.A(ori_ori_n161_), .Y(ori_ori_n162_));
  NO3        o134(.A(ori_ori_n162_), .B(ori_ori_n159_), .C(ori_ori_n156_), .Y(ori_ori_n163_));
  NAi41      o135(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n164_));
  INV        o136(.A(ori_ori_n164_), .Y(ori_ori_n165_));
  INV        o137(.A(f), .Y(ori_ori_n166_));
  INV        o138(.A(o), .Y(ori_ori_n167_));
  NOi31      o139(.An(i), .B(j), .C(h), .Y(ori_ori_n168_));
  NOi21      o140(.An(l), .B(m), .Y(ori_ori_n169_));
  NA2        o141(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  NO3        o142(.A(ori_ori_n170_), .B(ori_ori_n167_), .C(ori_ori_n166_), .Y(ori_ori_n171_));
  NA2        o143(.A(ori_ori_n171_), .B(ori_ori_n165_), .Y(ori_ori_n172_));
  OAI210     o144(.A0(ori_ori_n163_), .A1(ori_ori_n30_), .B0(ori_ori_n172_), .Y(ori_ori_n173_));
  NOi21      o145(.An(n), .B(m), .Y(ori_ori_n174_));
  OR2        o146(.A(ori_ori_n55_), .B(ori_ori_n54_), .Y(ori_ori_n175_));
  NAi21      o147(.An(j), .B(h), .Y(ori_ori_n176_));
  XN2        o148(.A(i), .B(h), .Y(ori_ori_n177_));
  NA2        o149(.A(ori_ori_n177_), .B(ori_ori_n176_), .Y(ori_ori_n178_));
  NOi31      o150(.An(k), .B(n), .C(m), .Y(ori_ori_n179_));
  NAi31      o151(.An(f), .B(e), .C(c), .Y(ori_ori_n180_));
  NA3        o152(.A(e), .B(c), .C(b), .Y(ori_ori_n181_));
  NAi32      o153(.An(m), .Bn(i), .C(k), .Y(ori_ori_n182_));
  INV        o154(.A(k), .Y(ori_ori_n183_));
  NAi21      o155(.An(n), .B(a), .Y(ori_ori_n184_));
  NO2        o156(.A(ori_ori_n184_), .B(ori_ori_n108_), .Y(ori_ori_n185_));
  NAi41      o157(.An(o), .B(m), .C(k), .D(h), .Y(ori_ori_n186_));
  NO2        o158(.A(ori_ori_n186_), .B(e), .Y(ori_ori_n187_));
  OR2        o159(.A(h), .B(o), .Y(ori_ori_n188_));
  NO2        o160(.A(ori_ori_n188_), .B(ori_ori_n72_), .Y(ori_ori_n189_));
  NA2        o161(.A(ori_ori_n189_), .B(ori_ori_n93_), .Y(ori_ori_n190_));
  NAi41      o162(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n191_));
  NO2        o163(.A(ori_ori_n191_), .B(ori_ori_n166_), .Y(ori_ori_n192_));
  NA2        o164(.A(ori_ori_n120_), .B(ori_ori_n77_), .Y(ori_ori_n193_));
  NAi21      o165(.An(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n194_));
  NAi21      o166(.An(h), .B(i), .Y(ori_ori_n195_));
  NA2        o167(.A(ori_ori_n133_), .B(k), .Y(ori_ori_n196_));
  NO2        o168(.A(ori_ori_n196_), .B(ori_ori_n195_), .Y(ori_ori_n197_));
  NA2        o169(.A(ori_ori_n197_), .B(ori_ori_n145_), .Y(ori_ori_n198_));
  NA3        o170(.A(ori_ori_n198_), .B(ori_ori_n194_), .C(ori_ori_n190_), .Y(ori_ori_n199_));
  NOi21      o171(.An(o), .B(e), .Y(ori_ori_n200_));
  NO2        o172(.A(ori_ori_n48_), .B(ori_ori_n49_), .Y(ori_ori_n201_));
  NA2        o173(.A(ori_ori_n201_), .B(ori_ori_n200_), .Y(ori_ori_n202_));
  NOi32      o174(.An(l), .Bn(j), .C(i), .Y(ori_ori_n203_));
  AOI210     o175(.A0(ori_ori_n50_), .A1(ori_ori_n62_), .B0(ori_ori_n203_), .Y(ori_ori_n204_));
  NAi21      o176(.An(f), .B(o), .Y(ori_ori_n205_));
  NO2        o177(.A(ori_ori_n205_), .B(ori_ori_n46_), .Y(ori_ori_n206_));
  NO2        o178(.A(ori_ori_n204_), .B(ori_ori_n202_), .Y(ori_ori_n207_));
  NOi41      o179(.An(ori_ori_n175_), .B(ori_ori_n207_), .C(ori_ori_n199_), .D(ori_ori_n173_), .Y(ori_ori_n208_));
  NA3        o180(.A(ori_ori_n44_), .B(c), .C(b), .Y(ori_ori_n209_));
  NO2        o181(.A(ori_ori_n193_), .B(ori_ori_n205_), .Y(ori_ori_n210_));
  NA3        o182(.A(ori_ori_n120_), .B(ori_ori_n119_), .C(ori_ori_n59_), .Y(ori_ori_n211_));
  NO2        o183(.A(ori_ori_n211_), .B(ori_ori_n147_), .Y(ori_ori_n212_));
  INV        o184(.A(ori_ori_n212_), .Y(ori_ori_n213_));
  NA3        o185(.A(e), .B(c), .C(b), .Y(ori_ori_n214_));
  NAi31      o186(.An(h), .B(l), .C(i), .Y(ori_ori_n215_));
  INV        o187(.A(ori_ori_n215_), .Y(ori_ori_n216_));
  NOi21      o188(.An(ori_ori_n216_), .B(ori_ori_n36_), .Y(ori_ori_n217_));
  NA2        o189(.A(ori_ori_n206_), .B(ori_ori_n217_), .Y(ori_ori_n218_));
  NAi32      o190(.An(j), .Bn(h), .C(i), .Y(ori_ori_n219_));
  NAi21      o191(.An(m), .B(l), .Y(ori_ori_n220_));
  NA2        o192(.A(h), .B(o), .Y(ori_ori_n221_));
  NA2        o193(.A(ori_ori_n218_), .B(ori_ori_n213_), .Y(ori_ori_n222_));
  NO2        o194(.A(ori_ori_n106_), .B(d), .Y(ori_ori_n223_));
  NO2        o195(.A(ori_ori_n75_), .B(ori_ori_n72_), .Y(ori_ori_n224_));
  NAi32      o196(.An(n), .Bn(m), .C(l), .Y(ori_ori_n225_));
  NO2        o197(.A(ori_ori_n225_), .B(ori_ori_n219_), .Y(ori_ori_n226_));
  NA2        o198(.A(ori_ori_n226_), .B(ori_ori_n137_), .Y(ori_ori_n227_));
  NAi31      o199(.An(k), .B(l), .C(j), .Y(ori_ori_n228_));
  INV        o200(.A(ori_ori_n227_), .Y(ori_ori_n229_));
  NO2        o201(.A(ori_ori_n229_), .B(ori_ori_n222_), .Y(ori_ori_n230_));
  NA2        o202(.A(ori_ori_n197_), .B(ori_ori_n146_), .Y(ori_ori_n231_));
  NAi21      o203(.An(m), .B(k), .Y(ori_ori_n232_));
  NO2        o204(.A(ori_ori_n177_), .B(ori_ori_n232_), .Y(ori_ori_n233_));
  NAi41      o205(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n234_));
  NO2        o206(.A(ori_ori_n234_), .B(ori_ori_n111_), .Y(ori_ori_n235_));
  NA2        o207(.A(ori_ori_n235_), .B(ori_ori_n233_), .Y(ori_ori_n236_));
  NA2        o208(.A(e), .B(c), .Y(ori_ori_n237_));
  NO3        o209(.A(ori_ori_n237_), .B(n), .C(d), .Y(ori_ori_n238_));
  NOi21      o210(.An(f), .B(h), .Y(ori_ori_n239_));
  NA2        o211(.A(ori_ori_n239_), .B(ori_ori_n85_), .Y(ori_ori_n240_));
  NO2        o212(.A(ori_ori_n240_), .B(ori_ori_n167_), .Y(ori_ori_n241_));
  NAi31      o213(.An(d), .B(e), .C(b), .Y(ori_ori_n242_));
  NO2        o214(.A(ori_ori_n95_), .B(ori_ori_n242_), .Y(ori_ori_n243_));
  NA2        o215(.A(ori_ori_n243_), .B(ori_ori_n241_), .Y(ori_ori_n244_));
  NA3        o216(.A(ori_ori_n244_), .B(ori_ori_n236_), .C(ori_ori_n231_), .Y(ori_ori_n245_));
  NO4        o217(.A(ori_ori_n234_), .B(ori_ori_n55_), .C(e), .D(ori_ori_n167_), .Y(ori_ori_n246_));
  NOi31      o218(.An(l), .B(n), .C(m), .Y(ori_ori_n247_));
  NA2        o219(.A(ori_ori_n247_), .B(ori_ori_n168_), .Y(ori_ori_n248_));
  NO2        o220(.A(ori_ori_n248_), .B(ori_ori_n147_), .Y(ori_ori_n249_));
  OR2        o221(.A(ori_ori_n249_), .B(ori_ori_n246_), .Y(ori_ori_n250_));
  NAi32      o222(.An(m), .Bn(j), .C(k), .Y(ori_ori_n251_));
  NAi41      o223(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n252_));
  NA2        o224(.A(ori_ori_n164_), .B(ori_ori_n252_), .Y(ori_ori_n253_));
  NOi31      o225(.An(j), .B(m), .C(k), .Y(ori_ori_n254_));
  NO2        o226(.A(ori_ori_n89_), .B(ori_ori_n254_), .Y(ori_ori_n255_));
  AN3        o227(.A(h), .B(o), .C(f), .Y(ori_ori_n256_));
  NAi31      o228(.An(ori_ori_n255_), .B(ori_ori_n256_), .C(ori_ori_n253_), .Y(ori_ori_n257_));
  NO2        o229(.A(ori_ori_n220_), .B(ori_ori_n219_), .Y(ori_ori_n258_));
  NO2        o230(.A(ori_ori_n170_), .B(o), .Y(ori_ori_n259_));
  NO2        o231(.A(ori_ori_n117_), .B(ori_ori_n59_), .Y(ori_ori_n260_));
  AOI220     o232(.A0(ori_ori_n260_), .A1(ori_ori_n259_), .B0(ori_ori_n192_), .B1(ori_ori_n258_), .Y(ori_ori_n261_));
  NA2        o233(.A(ori_ori_n261_), .B(ori_ori_n257_), .Y(ori_ori_n262_));
  NA3        o234(.A(h), .B(o), .C(f), .Y(ori_ori_n263_));
  NO2        o235(.A(ori_ori_n263_), .B(ori_ori_n51_), .Y(ori_ori_n264_));
  NA2        o236(.A(b), .B(ori_ori_n264_), .Y(ori_ori_n265_));
  NA2        o237(.A(o), .B(ori_ori_n81_), .Y(ori_ori_n266_));
  AO210      o238(.A0(ori_ori_n79_), .A1(ori_ori_n30_), .B0(ori_ori_n266_), .Y(ori_ori_n267_));
  NOi32      o239(.An(e), .Bn(b), .C(a), .Y(ori_ori_n268_));
  AN2        o240(.A(l), .B(j), .Y(ori_ori_n269_));
  NO2        o241(.A(ori_ori_n232_), .B(ori_ori_n269_), .Y(ori_ori_n270_));
  NO3        o242(.A(ori_ori_n234_), .B(e), .C(ori_ori_n167_), .Y(ori_ori_n271_));
  NA2        o243(.A(ori_ori_n161_), .B(ori_ori_n32_), .Y(ori_ori_n272_));
  AOI220     o244(.A0(ori_ori_n272_), .A1(ori_ori_n268_), .B0(ori_ori_n271_), .B1(ori_ori_n270_), .Y(ori_ori_n273_));
  NA4        o245(.A(ori_ori_n157_), .B(ori_ori_n62_), .C(o), .D(ori_ori_n166_), .Y(ori_ori_n274_));
  NA2        o246(.A(ori_ori_n38_), .B(ori_ori_n81_), .Y(ori_ori_n275_));
  NA3        o247(.A(ori_ori_n273_), .B(ori_ori_n267_), .C(ori_ori_n265_), .Y(ori_ori_n276_));
  NO4        o248(.A(ori_ori_n276_), .B(ori_ori_n262_), .C(ori_ori_n250_), .D(ori_ori_n245_), .Y(ori_ori_n277_));
  NA4        o249(.A(ori_ori_n277_), .B(ori_ori_n230_), .C(ori_ori_n208_), .D(ori_ori_n153_), .Y(ori10));
  NA3        o250(.A(m), .B(k), .C(i), .Y(ori_ori_n279_));
  NOi21      o251(.An(e), .B(f), .Y(ori_ori_n280_));
  INV        o252(.A(n), .Y(ori_ori_n281_));
  NAi31      o253(.An(b), .B(f), .C(c), .Y(ori_ori_n282_));
  INV        o254(.A(ori_ori_n282_), .Y(ori_ori_n283_));
  NOi32      o255(.An(k), .Bn(h), .C(j), .Y(ori_ori_n284_));
  NA2        o256(.A(ori_ori_n284_), .B(ori_ori_n174_), .Y(ori_ori_n285_));
  NA2        o257(.A(ori_ori_n121_), .B(ori_ori_n285_), .Y(ori_ori_n286_));
  NA2        o258(.A(ori_ori_n286_), .B(ori_ori_n283_), .Y(ori_ori_n287_));
  AN2        o259(.A(j), .B(h), .Y(ori_ori_n288_));
  NO3        o260(.A(n), .B(m), .C(k), .Y(ori_ori_n289_));
  NA2        o261(.A(ori_ori_n289_), .B(ori_ori_n288_), .Y(ori_ori_n290_));
  NO3        o262(.A(ori_ori_n290_), .B(ori_ori_n112_), .C(ori_ori_n166_), .Y(ori_ori_n291_));
  OR2        o263(.A(m), .B(k), .Y(ori_ori_n292_));
  NO2        o264(.A(ori_ori_n127_), .B(ori_ori_n292_), .Y(ori_ori_n293_));
  NA4        o265(.A(n), .B(f), .C(c), .D(ori_ori_n83_), .Y(ori_ori_n294_));
  NOi21      o266(.An(ori_ori_n293_), .B(ori_ori_n294_), .Y(ori_ori_n295_));
  NOi32      o267(.An(d), .Bn(a), .C(c), .Y(ori_ori_n296_));
  NA2        o268(.A(ori_ori_n296_), .B(ori_ori_n135_), .Y(ori_ori_n297_));
  NAi21      o269(.An(i), .B(o), .Y(ori_ori_n298_));
  NAi31      o270(.An(k), .B(m), .C(j), .Y(ori_ori_n299_));
  NO3        o271(.A(ori_ori_n299_), .B(ori_ori_n298_), .C(n), .Y(ori_ori_n300_));
  NOi21      o272(.An(ori_ori_n300_), .B(ori_ori_n297_), .Y(ori_ori_n301_));
  NO3        o273(.A(ori_ori_n301_), .B(ori_ori_n295_), .C(ori_ori_n291_), .Y(ori_ori_n302_));
  NO2        o274(.A(ori_ori_n294_), .B(ori_ori_n220_), .Y(ori_ori_n303_));
  NOi32      o275(.An(f), .Bn(d), .C(c), .Y(ori_ori_n304_));
  AOI220     o276(.A0(ori_ori_n304_), .A1(ori_ori_n226_), .B0(ori_ori_n303_), .B1(ori_ori_n168_), .Y(ori_ori_n305_));
  NA3        o277(.A(ori_ori_n305_), .B(ori_ori_n302_), .C(ori_ori_n287_), .Y(ori_ori_n306_));
  INV        o278(.A(e), .Y(ori_ori_n307_));
  NO2        o279(.A(ori_ori_n64_), .B(ori_ori_n307_), .Y(ori_ori_n308_));
  NOi21      o280(.An(o), .B(h), .Y(ori_ori_n309_));
  AN3        o281(.A(m), .B(l), .C(i), .Y(ori_ori_n310_));
  AN3        o282(.A(h), .B(o), .C(e), .Y(ori_ori_n311_));
  NO2        o283(.A(ori_ori_n64_), .B(n), .Y(ori_ori_n312_));
  NAi31      o284(.An(b), .B(c), .C(a), .Y(ori_ori_n313_));
  NO2        o285(.A(ori_ori_n313_), .B(n), .Y(ori_ori_n314_));
  NA2        o286(.A(ori_ori_n38_), .B(m), .Y(ori_ori_n315_));
  INV        o287(.A(ori_ori_n315_), .Y(ori_ori_n316_));
  NA2        o288(.A(ori_ori_n316_), .B(ori_ori_n314_), .Y(ori_ori_n317_));
  INV        o289(.A(ori_ori_n317_), .Y(ori_ori_n318_));
  NO3        o290(.A(ori_ori_n318_), .B(ori_ori_n312_), .C(ori_ori_n306_), .Y(ori_ori_n319_));
  NA2        o291(.A(i), .B(o), .Y(ori_ori_n320_));
  NOi21      o292(.An(a), .B(n), .Y(ori_ori_n321_));
  NOi21      o293(.An(d), .B(c), .Y(ori_ori_n322_));
  NA2        o294(.A(ori_ori_n322_), .B(ori_ori_n321_), .Y(ori_ori_n323_));
  NA3        o295(.A(i), .B(o), .C(f), .Y(ori_ori_n324_));
  OR2        o296(.A(ori_ori_n324_), .B(ori_ori_n47_), .Y(ori_ori_n325_));
  NA3        o297(.A(ori_ori_n310_), .B(ori_ori_n309_), .C(ori_ori_n135_), .Y(ori_ori_n326_));
  AOI210     o298(.A0(ori_ori_n326_), .A1(ori_ori_n325_), .B0(ori_ori_n323_), .Y(ori_ori_n327_));
  INV        o299(.A(ori_ori_n327_), .Y(ori_ori_n328_));
  OR2        o300(.A(n), .B(m), .Y(ori_ori_n329_));
  NO2        o301(.A(ori_ori_n329_), .B(ori_ori_n113_), .Y(ori_ori_n330_));
  INV        o302(.A(ori_ori_n136_), .Y(ori_ori_n331_));
  OAI210     o303(.A0(ori_ori_n330_), .A1(ori_ori_n129_), .B0(ori_ori_n331_), .Y(ori_ori_n332_));
  INV        o304(.A(ori_ori_n275_), .Y(ori_ori_n333_));
  NO2        o305(.A(ori_ori_n313_), .B(ori_ori_n36_), .Y(ori_ori_n334_));
  NAi21      o306(.An(k), .B(j), .Y(ori_ori_n335_));
  NA2        o307(.A(ori_ori_n195_), .B(ori_ori_n335_), .Y(ori_ori_n336_));
  NA3        o308(.A(ori_ori_n336_), .B(l), .C(ori_ori_n334_), .Y(ori_ori_n337_));
  NAi21      o309(.An(e), .B(d), .Y(ori_ori_n338_));
  INV        o310(.A(ori_ori_n338_), .Y(ori_ori_n339_));
  NO2        o311(.A(ori_ori_n196_), .B(ori_ori_n166_), .Y(ori_ori_n340_));
  NA3        o312(.A(ori_ori_n340_), .B(ori_ori_n339_), .C(ori_ori_n178_), .Y(ori_ori_n341_));
  NA3        o313(.A(ori_ori_n341_), .B(ori_ori_n337_), .C(ori_ori_n332_), .Y(ori_ori_n342_));
  NO2        o314(.A(ori_ori_n248_), .B(ori_ori_n166_), .Y(ori_ori_n343_));
  NA2        o315(.A(ori_ori_n343_), .B(ori_ori_n339_), .Y(ori_ori_n344_));
  NOi31      o316(.An(n), .B(m), .C(k), .Y(ori_ori_n345_));
  AOI220     o317(.A0(ori_ori_n345_), .A1(ori_ori_n288_), .B0(ori_ori_n174_), .B1(ori_ori_n37_), .Y(ori_ori_n346_));
  NAi31      o318(.An(o), .B(f), .C(c), .Y(ori_ori_n347_));
  NA2        o319(.A(ori_ori_n344_), .B(ori_ori_n227_), .Y(ori_ori_n348_));
  NOi41      o320(.An(ori_ori_n328_), .B(ori_ori_n348_), .C(ori_ori_n342_), .D(ori_ori_n207_), .Y(ori_ori_n349_));
  NOi32      o321(.An(c), .Bn(a), .C(b), .Y(ori_ori_n350_));
  NA2        o322(.A(ori_ori_n350_), .B(ori_ori_n81_), .Y(ori_ori_n351_));
  AN2        o323(.A(e), .B(d), .Y(ori_ori_n352_));
  NO2        o324(.A(ori_ori_n94_), .B(ori_ori_n351_), .Y(ori_ori_n353_));
  NO2        o325(.A(n), .B(ori_ori_n158_), .Y(ori_ori_n354_));
  NO4        o326(.A(ori_ori_n141_), .B(ori_ori_n72_), .C(ori_ori_n43_), .D(b), .Y(ori_ori_n355_));
  NA2        o327(.A(ori_ori_n283_), .B(ori_ori_n114_), .Y(ori_ori_n356_));
  NA2        o328(.A(l), .B(k), .Y(ori_ori_n357_));
  NA3        o329(.A(ori_ori_n357_), .B(j), .C(ori_ori_n174_), .Y(ori_ori_n358_));
  AOI210     o330(.A0(ori_ori_n182_), .A1(ori_ori_n251_), .B0(ori_ori_n59_), .Y(ori_ori_n359_));
  NOi21      o331(.An(ori_ori_n358_), .B(ori_ori_n359_), .Y(ori_ori_n360_));
  OR3        o332(.A(ori_ori_n360_), .B(ori_ori_n105_), .C(ori_ori_n97_), .Y(ori_ori_n361_));
  INV        o333(.A(ori_ori_n90_), .Y(ori_ori_n362_));
  NA3        o334(.A(ori_ori_n90_), .B(ori_ori_n361_), .C(ori_ori_n356_), .Y(ori_ori_n363_));
  NO4        o335(.A(ori_ori_n363_), .B(ori_ori_n355_), .C(ori_ori_n159_), .D(ori_ori_n353_), .Y(ori_ori_n364_));
  INV        o336(.A(e), .Y(ori_ori_n365_));
  NO2        o337(.A(ori_ori_n141_), .B(ori_ori_n43_), .Y(ori_ori_n366_));
  NAi31      o338(.An(j), .B(l), .C(i), .Y(ori_ori_n367_));
  OAI210     o339(.A0(ori_ori_n367_), .A1(ori_ori_n95_), .B0(ori_ori_n72_), .Y(ori_ori_n368_));
  NA3        o340(.A(ori_ori_n368_), .B(ori_ori_n366_), .C(ori_ori_n365_), .Y(ori_ori_n369_));
  NO2        o341(.A(ori_ori_n297_), .B(ori_ori_n275_), .Y(ori_ori_n370_));
  NO2        o342(.A(ori_ori_n138_), .B(ori_ori_n224_), .Y(ori_ori_n371_));
  NA3        o343(.A(ori_ori_n371_), .B(ori_ori_n369_), .C(ori_ori_n175_), .Y(ori_ori_n372_));
  OAI210     o344(.A0(ori_ori_n91_), .A1(ori_ori_n89_), .B0(n), .Y(ori_ori_n373_));
  NO2        o345(.A(ori_ori_n373_), .B(ori_ori_n94_), .Y(ori_ori_n374_));
  XO2        o346(.A(i), .B(h), .Y(ori_ori_n375_));
  NA3        o347(.A(ori_ori_n375_), .B(ori_ori_n120_), .C(n), .Y(ori_ori_n376_));
  NA3        o348(.A(ori_ori_n376_), .B(ori_ori_n346_), .C(ori_ori_n285_), .Y(ori_ori_n377_));
  NOi32      o349(.An(ori_ori_n377_), .Bn(ori_ori_n936_), .C(ori_ori_n209_), .Y(ori_ori_n378_));
  NAi31      o350(.An(c), .B(f), .C(d), .Y(ori_ori_n379_));
  BUFFER     o351(.A(ori_ori_n57_), .Y(ori_ori_n380_));
  NA2        o352(.A(ori_ori_n179_), .B(ori_ori_n77_), .Y(ori_ori_n381_));
  NO2        o353(.A(ori_ori_n134_), .B(ori_ori_n379_), .Y(ori_ori_n382_));
  INV        o354(.A(ori_ori_n382_), .Y(ori_ori_n383_));
  AN2        o355(.A(ori_ori_n217_), .B(ori_ori_n206_), .Y(ori_ori_n384_));
  NAi31      o356(.An(ori_ori_n384_), .B(ori_ori_n383_), .C(ori_ori_n380_), .Y(ori_ori_n385_));
  NO3        o357(.A(ori_ori_n385_), .B(ori_ori_n378_), .C(ori_ori_n372_), .Y(ori_ori_n386_));
  NA4        o358(.A(ori_ori_n386_), .B(ori_ori_n364_), .C(ori_ori_n349_), .D(ori_ori_n319_), .Y(ori11));
  NO2        o359(.A(ori_ori_n48_), .B(f), .Y(ori_ori_n388_));
  NA2        o360(.A(j), .B(o), .Y(ori_ori_n389_));
  NAi31      o361(.An(i), .B(m), .C(l), .Y(ori_ori_n390_));
  NA3        o362(.A(m), .B(k), .C(j), .Y(ori_ori_n391_));
  OAI220     o363(.A0(ori_ori_n391_), .A1(ori_ori_n94_), .B0(ori_ori_n390_), .B1(ori_ori_n389_), .Y(ori_ori_n392_));
  NA2        o364(.A(ori_ori_n392_), .B(ori_ori_n388_), .Y(ori_ori_n393_));
  NOi32      o365(.An(e), .Bn(b), .C(f), .Y(ori_ori_n394_));
  NA2        o366(.A(ori_ori_n35_), .B(j), .Y(ori_ori_n395_));
  NAi31      o367(.An(d), .B(e), .C(a), .Y(ori_ori_n396_));
  NO2        o368(.A(ori_ori_n396_), .B(n), .Y(ori_ori_n397_));
  NA2        o369(.A(j), .B(i), .Y(ori_ori_n398_));
  NO3        o370(.A(n), .B(d), .C(ori_ori_n83_), .Y(ori_ori_n399_));
  OR2        o371(.A(n), .B(c), .Y(ori_ori_n400_));
  NO2        o372(.A(ori_ori_n400_), .B(ori_ori_n110_), .Y(ori_ori_n401_));
  NA2        o373(.A(ori_ori_n392_), .B(f), .Y(ori_ori_n402_));
  NO2        o374(.A(ori_ori_n402_), .B(n), .Y(ori_ori_n403_));
  INV        o375(.A(ori_ori_n403_), .Y(ori_ori_n404_));
  NA2        o376(.A(ori_ori_n101_), .B(ori_ori_n31_), .Y(ori_ori_n405_));
  OAI220     o377(.A0(ori_ori_n405_), .A1(m), .B0(ori_ori_n395_), .B1(ori_ori_n182_), .Y(ori_ori_n406_));
  NOi41      o378(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n407_));
  NAi32      o379(.An(e), .Bn(b), .C(c), .Y(ori_ori_n408_));
  OR2        o380(.A(ori_ori_n408_), .B(ori_ori_n59_), .Y(ori_ori_n409_));
  AN2        o381(.A(ori_ori_n252_), .B(ori_ori_n234_), .Y(ori_ori_n410_));
  NA2        o382(.A(ori_ori_n410_), .B(ori_ori_n409_), .Y(ori_ori_n411_));
  OA210      o383(.A0(ori_ori_n411_), .A1(ori_ori_n407_), .B0(ori_ori_n406_), .Y(ori_ori_n412_));
  OAI220     o384(.A0(ori_ori_n299_), .A1(ori_ori_n298_), .B0(ori_ori_n390_), .B1(ori_ori_n389_), .Y(ori_ori_n413_));
  NAi21      o385(.An(d), .B(b), .Y(ori_ori_n414_));
  NO2        o386(.A(ori_ori_n414_), .B(ori_ori_n36_), .Y(ori_ori_n415_));
  NA2        o387(.A(h), .B(f), .Y(ori_ori_n416_));
  NO2        o388(.A(ori_ori_n416_), .B(ori_ori_n70_), .Y(ori_ori_n417_));
  NO3        o389(.A(ori_ori_n130_), .B(ori_ori_n127_), .C(o), .Y(ori_ori_n418_));
  AOI220     o390(.A0(ori_ori_n418_), .A1(b), .B0(ori_ori_n417_), .B1(ori_ori_n415_), .Y(ori_ori_n419_));
  INV        o391(.A(ori_ori_n419_), .Y(ori_ori_n420_));
  AN3        o392(.A(j), .B(h), .C(o), .Y(ori_ori_n421_));
  NO2        o393(.A(ori_ori_n108_), .B(c), .Y(ori_ori_n422_));
  NA3        o394(.A(ori_ori_n422_), .B(ori_ori_n421_), .C(ori_ori_n345_), .Y(ori_ori_n423_));
  NA3        o395(.A(f), .B(d), .C(b), .Y(ori_ori_n424_));
  INV        o396(.A(ori_ori_n423_), .Y(ori_ori_n425_));
  NO3        o397(.A(ori_ori_n425_), .B(ori_ori_n420_), .C(ori_ori_n412_), .Y(ori_ori_n426_));
  AN3        o398(.A(ori_ori_n426_), .B(ori_ori_n404_), .C(ori_ori_n393_), .Y(ori_ori_n427_));
  INV        o399(.A(k), .Y(ori_ori_n428_));
  NA4        o400(.A(ori_ori_n296_), .B(ori_ori_n309_), .C(ori_ori_n135_), .D(ori_ori_n81_), .Y(ori_ori_n429_));
  NAi41      o401(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n430_));
  OAI210     o402(.A0(ori_ori_n396_), .A1(n), .B0(ori_ori_n430_), .Y(ori_ori_n431_));
  NA2        o403(.A(ori_ori_n431_), .B(m), .Y(ori_ori_n432_));
  NAi31      o404(.An(h), .B(o), .C(f), .Y(ori_ori_n433_));
  NO3        o405(.A(f), .B(ori_ori_n48_), .C(ori_ori_n49_), .Y(ori_ori_n434_));
  NAi21      o406(.An(ori_ori_n434_), .B(ori_ori_n429_), .Y(ori_ori_n435_));
  NAi31      o407(.An(f), .B(h), .C(o), .Y(ori_ori_n436_));
  NO2        o408(.A(n), .B(c), .Y(ori_ori_n437_));
  NA3        o409(.A(ori_ori_n437_), .B(b), .C(m), .Y(ori_ori_n438_));
  NOi32      o410(.An(e), .Bn(a), .C(d), .Y(ori_ori_n439_));
  AOI210     o411(.A0(b), .A1(d), .B0(ori_ori_n439_), .Y(ori_ori_n440_));
  NA2        o412(.A(ori_ori_n435_), .B(i), .Y(ori_ori_n441_));
  NO3        o413(.A(ori_ori_n232_), .B(ori_ori_n45_), .C(n), .Y(ori_ori_n442_));
  NA3        o414(.A(ori_ori_n379_), .B(ori_ori_n125_), .C(ori_ori_n124_), .Y(ori_ori_n443_));
  NA2        o415(.A(ori_ori_n347_), .B(ori_ori_n180_), .Y(ori_ori_n444_));
  NA2        o416(.A(ori_ori_n443_), .B(ori_ori_n442_), .Y(ori_ori_n445_));
  NO2        o417(.A(ori_ori_n445_), .B(ori_ori_n62_), .Y(ori_ori_n446_));
  NA3        o418(.A(ori_ori_n407_), .B(ori_ori_n254_), .C(ori_ori_n35_), .Y(ori_ori_n447_));
  NOi32      o419(.An(e), .Bn(c), .C(f), .Y(ori_ori_n448_));
  NOi21      o420(.An(f), .B(o), .Y(ori_ori_n449_));
  NO2        o421(.A(ori_ori_n449_), .B(ori_ori_n164_), .Y(ori_ori_n450_));
  AOI220     o422(.A0(ori_ori_n450_), .A1(ori_ori_n293_), .B0(ori_ori_n448_), .B1(ori_ori_n129_), .Y(ori_ori_n451_));
  NA3        o423(.A(ori_ori_n451_), .B(ori_ori_n447_), .C(ori_ori_n132_), .Y(ori_ori_n452_));
  NOi21      o424(.An(j), .B(l), .Y(ori_ori_n453_));
  NO2        o425(.A(k), .B(ori_ori_n205_), .Y(ori_ori_n454_));
  NA2        o426(.A(ori_ori_n454_), .B(ori_ori_n453_), .Y(ori_ori_n455_));
  OR2        o427(.A(ori_ori_n455_), .B(ori_ori_n432_), .Y(ori_ori_n456_));
  NO2        o428(.A(ori_ori_n228_), .B(ori_ori_n436_), .Y(ori_ori_n457_));
  NO2        o429(.A(ori_ori_n396_), .B(ori_ori_n36_), .Y(ori_ori_n458_));
  NA2        o430(.A(ori_ori_n458_), .B(ori_ori_n457_), .Y(ori_ori_n459_));
  NA2        o431(.A(ori_ori_n459_), .B(ori_ori_n456_), .Y(ori_ori_n460_));
  NA2        o432(.A(ori_ori_n77_), .B(m), .Y(ori_ori_n461_));
  NO2        o433(.A(ori_ori_n395_), .B(ori_ori_n130_), .Y(ori_ori_n462_));
  NA3        o434(.A(ori_ori_n408_), .B(ori_ori_n209_), .C(ori_ori_n106_), .Y(ori_ori_n463_));
  NA2        o435(.A(ori_ori_n375_), .B(ori_ori_n120_), .Y(ori_ori_n464_));
  NO3        o436(.A(ori_ori_n294_), .B(ori_ori_n464_), .C(ori_ori_n62_), .Y(ori_ori_n465_));
  AOI210     o437(.A0(ori_ori_n463_), .A1(ori_ori_n462_), .B0(ori_ori_n465_), .Y(ori_ori_n466_));
  AN3        o438(.A(f), .B(d), .C(b), .Y(ori_ori_n467_));
  OAI210     o439(.A0(ori_ori_n467_), .A1(ori_ori_n93_), .B0(n), .Y(ori_ori_n468_));
  NA2        o440(.A(ori_ori_n375_), .B(ori_ori_n120_), .Y(ori_ori_n469_));
  AOI210     o441(.A0(ori_ori_n468_), .A1(ori_ori_n181_), .B0(ori_ori_n469_), .Y(ori_ori_n470_));
  NAi31      o442(.An(m), .B(n), .C(k), .Y(ori_ori_n471_));
  OR2        o443(.A(ori_ori_n97_), .B(ori_ori_n45_), .Y(ori_ori_n472_));
  NA2        o444(.A(ori_ori_n470_), .B(j), .Y(ori_ori_n473_));
  NA2        o445(.A(ori_ori_n473_), .B(ori_ori_n466_), .Y(ori_ori_n474_));
  NO4        o446(.A(ori_ori_n474_), .B(ori_ori_n460_), .C(ori_ori_n452_), .D(ori_ori_n446_), .Y(ori_ori_n475_));
  NA2        o447(.A(ori_ori_n281_), .B(ori_ori_n123_), .Y(ori_ori_n476_));
  NAi31      o448(.An(o), .B(h), .C(f), .Y(ori_ori_n477_));
  OA210      o449(.A0(ori_ori_n396_), .A1(n), .B0(ori_ori_n430_), .Y(ori_ori_n478_));
  NO2        o450(.A(ori_ori_n476_), .B(ori_ori_n391_), .Y(ori_ori_n479_));
  OR2        o451(.A(ori_ori_n48_), .B(ori_ori_n49_), .Y(ori_ori_n480_));
  OR2        o452(.A(ori_ori_n455_), .B(ori_ori_n480_), .Y(ori_ori_n481_));
  AN2        o453(.A(h), .B(f), .Y(ori_ori_n482_));
  NA2        o454(.A(ori_ori_n482_), .B(ori_ori_n33_), .Y(ori_ori_n483_));
  NO2        o455(.A(ori_ori_n483_), .B(ori_ori_n351_), .Y(ori_ori_n484_));
  AOI210     o456(.A0(ori_ori_n414_), .A1(ori_ori_n313_), .B0(ori_ori_n36_), .Y(ori_ori_n485_));
  AOI210     o457(.A0(ori_ori_n935_), .A1(ori_ori_n485_), .B0(ori_ori_n484_), .Y(ori_ori_n486_));
  NA2        o458(.A(ori_ori_n486_), .B(ori_ori_n481_), .Y(ori_ori_n487_));
  NO2        o459(.A(ori_ori_n195_), .B(f), .Y(ori_ori_n488_));
  NO2        o460(.A(ori_ori_n449_), .B(ori_ori_n45_), .Y(ori_ori_n489_));
  NO3        o461(.A(ori_ori_n489_), .B(ori_ori_n488_), .C(ori_ori_n31_), .Y(ori_ori_n490_));
  NA2        o462(.A(ori_ori_n243_), .B(ori_ori_n101_), .Y(ori_ori_n491_));
  NA2        o463(.A(ori_ori_n268_), .B(ori_ori_n81_), .Y(ori_ori_n492_));
  OR2        o464(.A(ori_ori_n492_), .B(ori_ori_n405_), .Y(ori_ori_n493_));
  OAI210     o465(.A0(ori_ori_n491_), .A1(ori_ori_n490_), .B0(ori_ori_n493_), .Y(ori_ori_n494_));
  NO3        o466(.A(ori_ori_n304_), .B(ori_ori_n146_), .C(ori_ori_n145_), .Y(ori_ori_n495_));
  NA2        o467(.A(ori_ori_n495_), .B(ori_ori_n180_), .Y(ori_ori_n496_));
  NA3        o468(.A(ori_ori_n496_), .B(ori_ori_n197_), .C(j), .Y(ori_ori_n497_));
  NO3        o469(.A(ori_ori_n347_), .B(ori_ori_n127_), .C(i), .Y(ori_ori_n498_));
  NA2        o470(.A(ori_ori_n350_), .B(ori_ori_n59_), .Y(ori_ori_n499_));
  NO3        o471(.A(ori_ori_n391_), .B(ori_ori_n499_), .C(ori_ori_n94_), .Y(ori_ori_n500_));
  INV        o472(.A(ori_ori_n500_), .Y(ori_ori_n501_));
  NA3        o473(.A(ori_ori_n501_), .B(ori_ori_n497_), .C(ori_ori_n302_), .Y(ori_ori_n502_));
  NO4        o474(.A(ori_ori_n502_), .B(ori_ori_n494_), .C(ori_ori_n487_), .D(ori_ori_n479_), .Y(ori_ori_n503_));
  NA4        o475(.A(ori_ori_n503_), .B(ori_ori_n475_), .C(ori_ori_n441_), .D(ori_ori_n427_), .Y(ori08));
  NO2        o476(.A(k), .B(h), .Y(ori_ori_n505_));
  AO210      o477(.A0(ori_ori_n195_), .A1(ori_ori_n335_), .B0(ori_ori_n505_), .Y(ori_ori_n506_));
  NO2        o478(.A(ori_ori_n506_), .B(ori_ori_n220_), .Y(ori_ori_n507_));
  INV        o479(.A(ori_ori_n448_), .Y(ori_ori_n508_));
  NO3        o480(.A(ori_ori_n279_), .B(ori_ori_n80_), .C(ori_ori_n167_), .Y(ori_ori_n509_));
  NA2        o481(.A(ori_ori_n509_), .B(e), .Y(ori_ori_n510_));
  AOI210     o482(.A0(ori_ori_n424_), .A1(ori_ori_n117_), .B0(ori_ori_n59_), .Y(ori_ori_n511_));
  NA3        o483(.A(ori_ori_n169_), .B(ori_ori_n34_), .C(h), .Y(ori_ori_n512_));
  AN2        o484(.A(l), .B(k), .Y(ori_ori_n513_));
  NA3        o485(.A(ori_ori_n513_), .B(ori_ori_n77_), .C(ori_ori_n49_), .Y(ori_ori_n514_));
  OAI210     o486(.A0(ori_ori_n512_), .A1(o), .B0(ori_ori_n514_), .Y(ori_ori_n515_));
  NA2        o487(.A(ori_ori_n515_), .B(ori_ori_n511_), .Y(ori_ori_n516_));
  NA3        o488(.A(ori_ori_n516_), .B(ori_ori_n510_), .C(ori_ori_n261_), .Y(ori_ori_n517_));
  AN2        o489(.A(ori_ori_n397_), .B(ori_ori_n71_), .Y(ori_ori_n518_));
  NO4        o490(.A(ori_ori_n127_), .B(ori_ori_n292_), .C(ori_ori_n80_), .D(o), .Y(ori_ori_n519_));
  NA2        o491(.A(ori_ori_n450_), .B(ori_ori_n258_), .Y(ori_ori_n520_));
  INV        o492(.A(ori_ori_n520_), .Y(ori_ori_n521_));
  NA2        o493(.A(ori_ori_n408_), .B(ori_ori_n472_), .Y(ori_ori_n522_));
  NO2        o494(.A(ori_ori_n357_), .B(ori_ori_n95_), .Y(ori_ori_n523_));
  NA2        o495(.A(ori_ori_n523_), .B(ori_ori_n522_), .Y(ori_ori_n524_));
  NO3        o496(.A(ori_ori_n232_), .B(ori_ori_n94_), .C(j), .Y(ori_ori_n525_));
  NAi21      o497(.An(ori_ori_n525_), .B(ori_ori_n514_), .Y(ori_ori_n526_));
  AOI220     o498(.A0(i), .A1(ori_ori_n303_), .B0(ori_ori_n526_), .B1(ori_ori_n52_), .Y(ori_ori_n527_));
  NA2        o499(.A(ori_ori_n524_), .B(ori_ori_n527_), .Y(ori_ori_n528_));
  NA3        o500(.A(ori_ori_n496_), .B(ori_ori_n247_), .C(ori_ori_n284_), .Y(ori_ori_n529_));
  NA3        o501(.A(m), .B(l), .C(k), .Y(ori_ori_n530_));
  INV        o502(.A(ori_ori_n529_), .Y(ori_ori_n531_));
  NO4        o503(.A(ori_ori_n531_), .B(ori_ori_n528_), .C(ori_ori_n521_), .D(ori_ori_n517_), .Y(ori_ori_n532_));
  NA2        o504(.A(ori_ori_n450_), .B(ori_ori_n293_), .Y(ori_ori_n533_));
  NO3        o505(.A(ori_ori_n297_), .B(ori_ori_n389_), .C(h), .Y(ori_ori_n534_));
  AOI210     o506(.A0(ori_ori_n534_), .A1(ori_ori_n81_), .B0(ori_ori_n370_), .Y(ori_ori_n535_));
  NA2        o507(.A(ori_ori_n535_), .B(ori_ori_n533_), .Y(ori_ori_n536_));
  INV        o508(.A(ori_ori_n513_), .Y(ori_ori_n537_));
  NO4        o509(.A(ori_ori_n495_), .B(ori_ori_n127_), .C(n), .D(i), .Y(ori_ori_n538_));
  BUFFER     o510(.A(h), .Y(ori_ori_n539_));
  NO2        o511(.A(ori_ori_n538_), .B(ori_ori_n498_), .Y(ori_ori_n540_));
  NO2        o512(.A(ori_ori_n540_), .B(ori_ori_n537_), .Y(ori_ori_n541_));
  AOI210     o513(.A0(ori_ori_n536_), .A1(l), .B0(ori_ori_n541_), .Y(ori_ori_n542_));
  NA2        o514(.A(ori_ori_n56_), .B(l), .Y(ori_ori_n543_));
  OR2        o515(.A(ori_ori_n543_), .B(ori_ori_n432_), .Y(ori_ori_n544_));
  NO3        o516(.A(ori_ori_n400_), .B(ori_ori_n110_), .C(ori_ori_n49_), .Y(ori_ori_n545_));
  AOI210     o517(.A0(ori_ori_n394_), .A1(n), .B0(ori_ori_n407_), .Y(ori_ori_n546_));
  NA2        o518(.A(ori_ori_n546_), .B(ori_ori_n410_), .Y(ori_ori_n547_));
  NO3        o519(.A(ori_ori_n127_), .B(ori_ori_n292_), .C(ori_ori_n80_), .Y(ori_ori_n548_));
  AOI220     o520(.A0(ori_ori_n548_), .A1(ori_ori_n192_), .B0(ori_ori_n444_), .B1(ori_ori_n226_), .Y(ori_ori_n549_));
  NAi31      o521(.An(ori_ori_n440_), .B(ori_ori_n68_), .C(ori_ori_n59_), .Y(ori_ori_n550_));
  NA2        o522(.A(ori_ori_n550_), .B(ori_ori_n549_), .Y(ori_ori_n551_));
  NO2        o523(.A(ori_ori_n220_), .B(ori_ori_n98_), .Y(ori_ori_n552_));
  AOI220     o524(.A0(ori_ori_n552_), .A1(ori_ori_n450_), .B0(ori_ori_n525_), .B1(ori_ori_n511_), .Y(ori_ori_n553_));
  NO2        o525(.A(ori_ori_n530_), .B(ori_ori_n66_), .Y(ori_ori_n554_));
  NA2        o526(.A(ori_ori_n554_), .B(ori_ori_n431_), .Y(ori_ori_n555_));
  NO2        o527(.A(ori_ori_n433_), .B(ori_ori_n84_), .Y(ori_ori_n556_));
  NA2        o528(.A(ori_ori_n556_), .B(ori_ori_n485_), .Y(ori_ori_n557_));
  NA3        o529(.A(ori_ori_n557_), .B(ori_ori_n555_), .C(ori_ori_n553_), .Y(ori_ori_n558_));
  OR2        o530(.A(ori_ori_n558_), .B(ori_ori_n551_), .Y(ori_ori_n559_));
  NA3        o531(.A(ori_ori_n546_), .B(ori_ori_n410_), .C(ori_ori_n409_), .Y(ori_ori_n560_));
  NA4        o532(.A(ori_ori_n560_), .B(ori_ori_n169_), .C(ori_ori_n335_), .D(ori_ori_n31_), .Y(ori_ori_n561_));
  NO2        o533(.A(ori_ori_n357_), .B(ori_ori_n320_), .Y(ori_ori_n562_));
  NA2        o534(.A(ori_ori_n562_), .B(ori_ori_n201_), .Y(ori_ori_n563_));
  NA2        o535(.A(ori_ori_n563_), .B(ori_ori_n561_), .Y(ori_ori_n564_));
  BUFFER     o536(.A(ori_ori_n554_), .Y(ori_ori_n565_));
  NA2        o537(.A(ori_ori_n565_), .B(ori_ori_n185_), .Y(ori_ori_n566_));
  NO2        o538(.A(ori_ori_n478_), .B(ori_ori_n49_), .Y(ori_ori_n567_));
  AOI210     o539(.A0(ori_ori_n562_), .A1(ori_ori_n567_), .B0(ori_ori_n249_), .Y(ori_ori_n568_));
  NO2        o540(.A(ori_ori_n530_), .B(ori_ori_n477_), .Y(ori_ori_n569_));
  NA2        o541(.A(ori_ori_n59_), .B(ori_ori_n569_), .Y(ori_ori_n570_));
  NA3        o542(.A(ori_ori_n570_), .B(ori_ori_n568_), .C(ori_ori_n566_), .Y(ori_ori_n571_));
  NOi41      o543(.An(ori_ori_n544_), .B(ori_ori_n571_), .C(ori_ori_n564_), .D(ori_ori_n559_), .Y(ori_ori_n572_));
  NO3        o544(.A(ori_ori_n255_), .B(ori_ori_n221_), .C(ori_ori_n80_), .Y(ori_ori_n573_));
  NA2        o545(.A(ori_ori_n573_), .B(ori_ori_n547_), .Y(ori_ori_n574_));
  NA2        o546(.A(ori_ori_n574_), .B(ori_ori_n305_), .Y(ori_ori_n575_));
  BUFFER     o547(.A(ori_ori_n477_), .Y(ori_ori_n576_));
  NO2        o548(.A(ori_ori_n408_), .B(ori_ori_n59_), .Y(ori_ori_n577_));
  NA2        o549(.A(ori_ori_n573_), .B(ori_ori_n577_), .Y(ori_ori_n578_));
  OAI210     o550(.A0(ori_ori_n512_), .A1(ori_ori_n294_), .B0(ori_ori_n578_), .Y(ori_ori_n579_));
  NO2        o551(.A(ori_ori_n495_), .B(n), .Y(ori_ori_n580_));
  NA2        o552(.A(ori_ori_n580_), .B(ori_ori_n507_), .Y(ori_ori_n581_));
  NO2        o553(.A(ori_ori_n237_), .B(ori_ori_n184_), .Y(ori_ori_n582_));
  OAI210     o554(.A0(ori_ori_n71_), .A1(ori_ori_n68_), .B0(ori_ori_n582_), .Y(ori_ori_n583_));
  INV        o555(.A(ori_ori_n583_), .Y(ori_ori_n584_));
  NA2        o556(.A(ori_ori_n519_), .B(ori_ori_n260_), .Y(ori_ori_n585_));
  NA2        o557(.A(ori_ori_n434_), .B(ori_ori_n269_), .Y(ori_ori_n586_));
  AN2        o558(.A(ori_ori_n586_), .B(ori_ori_n585_), .Y(ori_ori_n587_));
  NAi31      o559(.An(ori_ori_n584_), .B(ori_ori_n587_), .C(ori_ori_n581_), .Y(ori_ori_n588_));
  NO3        o560(.A(ori_ori_n588_), .B(ori_ori_n579_), .C(ori_ori_n575_), .Y(ori_ori_n589_));
  NA4        o561(.A(ori_ori_n589_), .B(ori_ori_n572_), .C(ori_ori_n542_), .D(ori_ori_n532_), .Y(ori09));
  NA3        o562(.A(m), .B(l), .C(i), .Y(ori_ori_n591_));
  INV        o563(.A(ori_ori_n252_), .Y(ori_ori_n592_));
  NO2        o564(.A(ori_ori_n91_), .B(ori_ori_n89_), .Y(ori_ori_n593_));
  NOi31      o565(.An(k), .B(m), .C(l), .Y(ori_ori_n594_));
  NO2        o566(.A(ori_ori_n254_), .B(ori_ori_n594_), .Y(ori_ori_n595_));
  AOI210     o567(.A0(ori_ori_n595_), .A1(ori_ori_n593_), .B0(ori_ori_n436_), .Y(ori_ori_n596_));
  NA2        o568(.A(ori_ori_n596_), .B(ori_ori_n592_), .Y(ori_ori_n597_));
  NA2        o569(.A(ori_ori_n506_), .B(ori_ori_n98_), .Y(ori_ori_n598_));
  NA3        o570(.A(ori_ori_n598_), .B(ori_ori_n143_), .C(e), .Y(ori_ori_n599_));
  NA4        o571(.A(ori_ori_n599_), .B(ori_ori_n597_), .C(ori_ori_n451_), .D(ori_ori_n57_), .Y(ori_ori_n600_));
  NO2        o572(.A(f), .B(ori_ori_n367_), .Y(ori_ori_n601_));
  NA2        o573(.A(ori_ori_n601_), .B(ori_ori_n143_), .Y(ori_ori_n602_));
  NA2        o574(.A(f), .B(m), .Y(ori_ori_n603_));
  NO2        o575(.A(ori_ori_n603_), .B(ori_ori_n39_), .Y(ori_ori_n604_));
  NOi32      o576(.An(o), .Bn(f), .C(d), .Y(ori_ori_n605_));
  NA4        o577(.A(ori_ori_n605_), .B(ori_ori_n437_), .C(b), .D(m), .Y(ori_ori_n606_));
  INV        o578(.A(ori_ori_n606_), .Y(ori_ori_n607_));
  AOI210     o579(.A0(ori_ori_n604_), .A1(ori_ori_n401_), .B0(ori_ori_n607_), .Y(ori_ori_n608_));
  NA3        o580(.A(ori_ori_n228_), .B(ori_ori_n204_), .C(ori_ori_n86_), .Y(ori_ori_n609_));
  NA3        o581(.A(a), .B(f), .C(ori_ori_n59_), .Y(ori_ori_n610_));
  NO3        o582(.A(ori_ori_n610_), .B(ori_ori_n49_), .C(ori_ori_n167_), .Y(ori_ori_n611_));
  NA2        o583(.A(ori_ori_n609_), .B(ori_ori_n611_), .Y(ori_ori_n612_));
  NAi41      o584(.An(ori_ori_n362_), .B(ori_ori_n612_), .C(ori_ori_n608_), .D(ori_ori_n602_), .Y(ori_ori_n613_));
  NO4        o585(.A(ori_ori_n449_), .B(ori_ori_n95_), .C(ori_ori_n242_), .D(ori_ori_n113_), .Y(ori_ori_n614_));
  NO2        o586(.A(ori_ori_n471_), .B(ori_ori_n242_), .Y(ori_ori_n615_));
  AN2        o587(.A(ori_ori_n615_), .B(ori_ori_n488_), .Y(ori_ori_n616_));
  NO2        o588(.A(ori_ori_n616_), .B(ori_ori_n614_), .Y(ori_ori_n617_));
  NOi21      o589(.An(ori_ori_n175_), .B(ori_ori_n224_), .Y(ori_ori_n618_));
  NA2        o590(.A(c), .B(ori_ori_n83_), .Y(ori_ori_n619_));
  NO2        o591(.A(ori_ori_n619_), .B(ori_ori_n307_), .Y(ori_ori_n620_));
  NA3        o592(.A(ori_ori_n620_), .B(ori_ori_n377_), .C(f), .Y(ori_ori_n621_));
  OR2        o593(.A(ori_ori_n477_), .B(n), .Y(ori_ori_n622_));
  NA3        o594(.A(ori_ori_n621_), .B(ori_ori_n618_), .C(ori_ori_n617_), .Y(ori_ori_n623_));
  NO3        o595(.A(ori_ori_n623_), .B(ori_ori_n613_), .C(ori_ori_n600_), .Y(ori_ori_n624_));
  NO2        o596(.A(ori_ori_n98_), .B(ori_ori_n95_), .Y(ori_ori_n625_));
  NO2        o597(.A(ori_ori_n180_), .B(ori_ori_n176_), .Y(ori_ori_n626_));
  AOI220     o598(.A0(ori_ori_n626_), .A1(ori_ori_n179_), .B0(ori_ori_n223_), .B1(ori_ori_n625_), .Y(ori_ori_n627_));
  INV        o599(.A(ori_ori_n627_), .Y(ori_ori_n628_));
  NA2        o600(.A(e), .B(d), .Y(ori_ori_n629_));
  OAI220     o601(.A0(ori_ori_n629_), .A1(c), .B0(ori_ori_n237_), .B1(d), .Y(ori_ori_n630_));
  NA3        o602(.A(ori_ori_n630_), .B(ori_ori_n340_), .C(ori_ori_n375_), .Y(ori_ori_n631_));
  NA2        o603(.A(ori_ori_n450_), .B(ori_ori_n258_), .Y(ori_ori_n632_));
  NA3        o604(.A(k), .B(ori_ori_n60_), .C(ori_ori_n31_), .Y(ori_ori_n633_));
  NA3        o605(.A(ori_ori_n633_), .B(ori_ori_n632_), .C(ori_ori_n631_), .Y(ori_ori_n634_));
  NO2        o606(.A(ori_ori_n634_), .B(ori_ori_n628_), .Y(ori_ori_n635_));
  OR2        o607(.A(ori_ori_n508_), .B(ori_ori_n170_), .Y(ori_ori_n636_));
  OAI220     o608(.A0(ori_ori_n449_), .A1(ori_ori_n45_), .B0(ori_ori_n221_), .B1(j), .Y(ori_ori_n637_));
  NA2        o609(.A(ori_ori_n637_), .B(ori_ori_n615_), .Y(ori_ori_n638_));
  INV        o610(.A(ori_ori_n638_), .Y(ori_ori_n639_));
  INV        o611(.A(ori_ori_n606_), .Y(ori_ori_n640_));
  BUFFER     o612(.A(ori_ori_n640_), .Y(ori_ori_n641_));
  NO2        o613(.A(ori_ori_n641_), .B(ori_ori_n639_), .Y(ori_ori_n642_));
  AO220      o614(.A0(ori_ori_n340_), .A1(ori_ori_n539_), .B0(ori_ori_n129_), .B1(f), .Y(ori_ori_n643_));
  OAI210     o615(.A0(ori_ori_n643_), .A1(ori_ori_n343_), .B0(ori_ori_n630_), .Y(ori_ori_n644_));
  NO2        o616(.A(ori_ori_n324_), .B(ori_ori_n47_), .Y(ori_ori_n645_));
  AN3        o617(.A(ori_ori_n644_), .B(ori_ori_n642_), .C(ori_ori_n636_), .Y(ori_ori_n646_));
  NA3        o618(.A(ori_ori_n646_), .B(ori_ori_n635_), .C(ori_ori_n624_), .Y(ori12));
  NO2        o619(.A(ori_ori_n338_), .B(c), .Y(ori_ori_n648_));
  NO4        o620(.A(ori_ori_n329_), .B(ori_ori_n195_), .C(ori_ori_n428_), .D(ori_ori_n167_), .Y(ori_ori_n649_));
  NA2        o621(.A(ori_ori_n649_), .B(ori_ori_n648_), .Y(ori_ori_n650_));
  NA2        o622(.A(ori_ori_n401_), .B(ori_ori_n645_), .Y(ori_ori_n651_));
  NO2        o623(.A(ori_ori_n338_), .B(ori_ori_n83_), .Y(ori_ori_n652_));
  NO2        o624(.A(ori_ori_n593_), .B(ori_ori_n263_), .Y(ori_ori_n653_));
  NO2        o625(.A(ori_ori_n477_), .B(ori_ori_n279_), .Y(ori_ori_n654_));
  AOI220     o626(.A0(ori_ori_n654_), .A1(ori_ori_n399_), .B0(ori_ori_n653_), .B1(ori_ori_n652_), .Y(ori_ori_n655_));
  NA4        o627(.A(ori_ori_n655_), .B(ori_ori_n651_), .C(ori_ori_n650_), .D(ori_ori_n328_), .Y(ori_ori_n656_));
  AOI210     o628(.A0(ori_ori_n182_), .A1(ori_ori_n251_), .B0(ori_ori_n155_), .Y(ori_ori_n657_));
  AOI210     o629(.A0(ori_ori_n248_), .A1(ori_ori_n290_), .B0(ori_ori_n167_), .Y(ori_ori_n658_));
  NA2        o630(.A(ori_ori_n658_), .B(ori_ori_n304_), .Y(ori_ori_n659_));
  NO2        o631(.A(ori_ori_n461_), .B(ori_ori_n205_), .Y(ori_ori_n660_));
  NO2        o632(.A(ori_ori_n433_), .B(ori_ori_n591_), .Y(ori_ori_n661_));
  NO2        o633(.A(ori_ori_n112_), .B(ori_ori_n184_), .Y(ori_ori_n662_));
  NA2        o634(.A(ori_ori_n662_), .B(ori_ori_n187_), .Y(ori_ori_n663_));
  NA2        o635(.A(ori_ori_n663_), .B(ori_ori_n659_), .Y(ori_ori_n664_));
  OR2        o636(.A(ori_ori_n238_), .B(ori_ori_n652_), .Y(ori_ori_n665_));
  NA2        o637(.A(ori_ori_n665_), .B(ori_ori_n264_), .Y(ori_ori_n666_));
  NO3        o638(.A(ori_ori_n95_), .B(ori_ori_n113_), .C(ori_ori_n167_), .Y(ori_ori_n667_));
  NA2        o639(.A(ori_ori_n667_), .B(ori_ori_n394_), .Y(ori_ori_n668_));
  NA3        o640(.A(ori_ori_n330_), .B(ori_ori_n322_), .C(ori_ori_n135_), .Y(ori_ori_n669_));
  NA3        o641(.A(ori_ori_n669_), .B(ori_ori_n668_), .C(ori_ori_n666_), .Y(ori_ori_n670_));
  NO3        o642(.A(ori_ori_n670_), .B(ori_ori_n664_), .C(ori_ori_n656_), .Y(ori_ori_n671_));
  NA2        o643(.A(ori_ori_n408_), .B(ori_ori_n106_), .Y(ori_ori_n672_));
  NOi21      o644(.An(ori_ori_n31_), .B(ori_ori_n471_), .Y(ori_ori_n673_));
  NA2        o645(.A(ori_ori_n673_), .B(ori_ori_n672_), .Y(ori_ori_n674_));
  INV        o646(.A(ori_ori_n674_), .Y(ori_ori_n675_));
  INV        o647(.A(ori_ori_n236_), .Y(ori_ori_n676_));
  NO2        o648(.A(ori_ori_n373_), .B(ori_ori_n221_), .Y(ori_ori_n677_));
  INV        o649(.A(ori_ori_n677_), .Y(ori_ori_n678_));
  NO2        o650(.A(ori_ori_n678_), .B(ori_ori_n106_), .Y(ori_ori_n679_));
  INV        o651(.A(ori_ori_n273_), .Y(ori_ori_n680_));
  NO4        o652(.A(ori_ori_n680_), .B(ori_ori_n679_), .C(ori_ori_n676_), .D(ori_ori_n675_), .Y(ori_ori_n681_));
  NA2        o653(.A(ori_ori_n258_), .B(o), .Y(ori_ori_n682_));
  NA2        o654(.A(ori_ori_n123_), .B(i), .Y(ori_ori_n683_));
  NA2        o655(.A(ori_ori_n35_), .B(i), .Y(ori_ori_n684_));
  NO2        o656(.A(ori_ori_n106_), .B(ori_ori_n59_), .Y(ori_ori_n685_));
  OR2        o657(.A(ori_ori_n685_), .B(ori_ori_n407_), .Y(ori_ori_n686_));
  NA2        o658(.A(ori_ori_n408_), .B(ori_ori_n282_), .Y(ori_ori_n687_));
  AOI210     o659(.A0(ori_ori_n687_), .A1(n), .B0(ori_ori_n686_), .Y(ori_ori_n688_));
  NO2        o660(.A(ori_ori_n688_), .B(ori_ori_n682_), .Y(ori_ori_n689_));
  NO2        o661(.A(ori_ori_n477_), .B(ori_ori_n367_), .Y(ori_ori_n690_));
  NA3        o662(.A(ori_ori_n256_), .B(ori_ori_n453_), .C(i), .Y(ori_ori_n691_));
  OAI210     o663(.A0(ori_ori_n324_), .A1(ori_ori_n228_), .B0(ori_ori_n691_), .Y(ori_ori_n692_));
  OAI220     o664(.A0(ori_ori_n692_), .A1(ori_ori_n690_), .B0(ori_ori_n485_), .B1(ori_ori_n545_), .Y(ori_ori_n693_));
  NA2        o665(.A(ori_ori_n439_), .B(ori_ori_n81_), .Y(ori_ori_n694_));
  OR3        o666(.A(ori_ori_n228_), .B(ori_ori_n320_), .C(f), .Y(ori_ori_n695_));
  NA3        o667(.A(ori_ori_n453_), .B(ori_ori_n56_), .C(i), .Y(ori_ori_n696_));
  OA220      o668(.A0(ori_ori_n696_), .A1(ori_ori_n694_), .B0(ori_ori_n695_), .B1(ori_ori_n432_), .Y(ori_ori_n697_));
  NA3        o669(.A(ori_ori_n239_), .B(ori_ori_n85_), .C(o), .Y(ori_ori_n698_));
  AOI210     o670(.A0(ori_ori_n483_), .A1(ori_ori_n698_), .B0(m), .Y(ori_ori_n699_));
  OAI210     o671(.A0(ori_ori_n699_), .A1(ori_ori_n653_), .B0(ori_ori_n238_), .Y(ori_ori_n700_));
  INV        o672(.A(ori_ori_n696_), .Y(ori_ori_n701_));
  NA2        o673(.A(ori_ori_n701_), .B(ori_ori_n201_), .Y(ori_ori_n702_));
  NA4        o674(.A(ori_ori_n702_), .B(ori_ori_n700_), .C(ori_ori_n697_), .D(ori_ori_n693_), .Y(ori_ori_n703_));
  NO2        o675(.A(ori_ori_n279_), .B(ori_ori_n66_), .Y(ori_ori_n704_));
  OAI210     o676(.A0(ori_ori_n704_), .A1(ori_ori_n660_), .B0(ori_ori_n185_), .Y(ori_ori_n705_));
  NO2        o677(.A(ori_ori_n346_), .B(ori_ori_n167_), .Y(ori_ori_n706_));
  AOI220     o678(.A0(ori_ori_n706_), .A1(ori_ori_n283_), .B0(ori_ori_n665_), .B1(ori_ori_n171_), .Y(ori_ori_n707_));
  AOI220     o679(.A0(ori_ori_n654_), .A1(ori_ori_n662_), .B0(ori_ori_n431_), .B1(ori_ori_n65_), .Y(ori_ori_n708_));
  NA3        o680(.A(ori_ori_n708_), .B(ori_ori_n707_), .C(ori_ori_n705_), .Y(ori_ori_n709_));
  NA2        o681(.A(ori_ori_n661_), .B(ori_ori_n399_), .Y(ori_ori_n710_));
  NA2        o682(.A(ori_ori_n699_), .B(ori_ori_n652_), .Y(ori_ori_n711_));
  NA2        o683(.A(ori_ori_n462_), .B(ori_ori_n394_), .Y(ori_ori_n712_));
  NA3        o684(.A(ori_ori_n712_), .B(ori_ori_n711_), .C(ori_ori_n710_), .Y(ori_ori_n713_));
  NO4        o685(.A(ori_ori_n713_), .B(ori_ori_n709_), .C(ori_ori_n703_), .D(ori_ori_n689_), .Y(ori_ori_n714_));
  NAi31      o686(.An(ori_ori_n102_), .B(ori_ori_n311_), .C(n), .Y(ori_ori_n715_));
  NO3        o687(.A(ori_ori_n89_), .B(ori_ori_n254_), .C(ori_ori_n594_), .Y(ori_ori_n716_));
  NO2        o688(.A(ori_ori_n716_), .B(ori_ori_n715_), .Y(ori_ori_n717_));
  NO3        o689(.A(h), .B(ori_ori_n102_), .C(ori_ori_n307_), .Y(ori_ori_n718_));
  AOI210     o690(.A0(ori_ori_n718_), .A1(ori_ori_n368_), .B0(ori_ori_n717_), .Y(ori_ori_n719_));
  INV        o691(.A(ori_ori_n719_), .Y(ori_ori_n720_));
  NA2        o692(.A(ori_ori_n180_), .B(ori_ori_n125_), .Y(ori_ori_n721_));
  NO3        o693(.A(ori_ori_n226_), .B(ori_ori_n330_), .C(ori_ori_n129_), .Y(ori_ori_n722_));
  NOi31      o694(.An(ori_ori_n721_), .B(ori_ori_n722_), .C(ori_ori_n167_), .Y(ori_ori_n723_));
  NAi21      o695(.An(ori_ori_n408_), .B(ori_ori_n706_), .Y(ori_ori_n724_));
  NA2        o696(.A(ori_ori_n355_), .B(o), .Y(ori_ori_n725_));
  NA2        o697(.A(ori_ori_n725_), .B(ori_ori_n724_), .Y(ori_ori_n726_));
  NA2        o698(.A(ori_ori_n657_), .B(ori_ori_n648_), .Y(ori_ori_n727_));
  OAI220     o699(.A0(ori_ori_n654_), .A1(ori_ori_n661_), .B0(ori_ori_n401_), .B1(ori_ori_n314_), .Y(ori_ori_n728_));
  NA3        o700(.A(ori_ori_n728_), .B(ori_ori_n727_), .C(ori_ori_n447_), .Y(ori_ori_n729_));
  NA3        o701(.A(ori_ori_n687_), .B(ori_ori_n359_), .C(ori_ori_n35_), .Y(ori_ori_n730_));
  INV        o702(.A(ori_ori_n246_), .Y(ori_ori_n731_));
  NA2        o703(.A(ori_ori_n731_), .B(ori_ori_n730_), .Y(ori_ori_n732_));
  OR2        o704(.A(ori_ori_n732_), .B(ori_ori_n729_), .Y(ori_ori_n733_));
  NO4        o705(.A(ori_ori_n733_), .B(ori_ori_n726_), .C(ori_ori_n723_), .D(ori_ori_n720_), .Y(ori_ori_n734_));
  NA4        o706(.A(ori_ori_n734_), .B(ori_ori_n714_), .C(ori_ori_n681_), .D(ori_ori_n671_), .Y(ori13));
  AN2        o707(.A(d), .B(c), .Y(ori_ori_n736_));
  NA2        o708(.A(ori_ori_n736_), .B(ori_ori_n83_), .Y(ori_ori_n737_));
  NAi32      o709(.An(f), .Bn(e), .C(c), .Y(ori_ori_n738_));
  NA3        o710(.A(k), .B(j), .C(i), .Y(ori_ori_n739_));
  NO2        o711(.A(f), .B(c), .Y(ori_ori_n740_));
  NOi21      o712(.An(ori_ori_n740_), .B(ori_ori_n329_), .Y(ori_ori_n741_));
  OR2        o713(.A(m), .B(i), .Y(ori_ori_n742_));
  AN3        o714(.A(o), .B(f), .C(c), .Y(ori_ori_n743_));
  NA3        o715(.A(l), .B(k), .C(j), .Y(ori_ori_n744_));
  NA2        o716(.A(i), .B(h), .Y(ori_ori_n745_));
  NO3        o717(.A(ori_ori_n745_), .B(ori_ori_n744_), .C(ori_ori_n95_), .Y(ori_ori_n746_));
  NO3        o718(.A(ori_ori_n103_), .B(ori_ori_n214_), .C(ori_ori_n167_), .Y(ori_ori_n747_));
  NA2        o719(.A(c), .B(b), .Y(ori_ori_n748_));
  NO2        o720(.A(ori_ori_n390_), .B(ori_ori_n436_), .Y(ori_ori_n749_));
  NA4        o721(.A(ori_ori_n63_), .B(ori_ori_n62_), .C(o), .D(ori_ori_n166_), .Y(ori_ori_n750_));
  NA4        o722(.A(ori_ori_n421_), .B(m), .C(ori_ori_n80_), .D(ori_ori_n166_), .Y(ori_ori_n751_));
  NA3        o723(.A(ori_ori_n751_), .B(ori_ori_n274_), .C(ori_ori_n750_), .Y(ori_ori_n752_));
  NO2        o724(.A(ori_ori_n752_), .B(ori_ori_n749_), .Y(ori_ori_n753_));
  OAI220     o725(.A0(ori_ori_n576_), .A1(ori_ori_n499_), .B0(ori_ori_n753_), .B1(ori_ori_n430_), .Y(ori_ori_n754_));
  NOi31      o726(.An(m), .B(n), .C(f), .Y(ori_ori_n755_));
  NA2        o727(.A(ori_ori_n755_), .B(ori_ori_n38_), .Y(ori_ori_n756_));
  OAI220     o728(.A0(ori_ori_n934_), .A1(ori_ori_n756_), .B0(ori_ori_n622_), .B1(ori_ori_n313_), .Y(ori_ori_n757_));
  NO3        o729(.A(ori_ori_n757_), .B(ori_ori_n754_), .C(ori_ori_n584_), .Y(ori_ori_n758_));
  NA2        o730(.A(c), .B(b), .Y(ori_ori_n759_));
  NO2        o731(.A(a), .B(ori_ori_n759_), .Y(ori_ori_n760_));
  OAI210     o732(.A0(ori_ori_n308_), .A1(ori_ori_n604_), .B0(ori_ori_n760_), .Y(ori_ori_n761_));
  NA3        o733(.A(ori_ori_n314_), .B(ori_ori_n413_), .C(f), .Y(ori_ori_n762_));
  INV        o734(.A(ori_ori_n762_), .Y(ori_ori_n763_));
  NA2        o735(.A(ori_ori_n204_), .B(ori_ori_n86_), .Y(ori_ori_n764_));
  OAI210     o736(.A0(ori_ori_n764_), .A1(ori_ori_n216_), .B0(o), .Y(ori_ori_n765_));
  NO2        o737(.A(f), .B(ori_ori_n748_), .Y(ori_ori_n766_));
  INV        o738(.A(ori_ori_n766_), .Y(ori_ori_n767_));
  NO2        o739(.A(ori_ori_n765_), .B(ori_ori_n767_), .Y(ori_ori_n768_));
  AOI210     o740(.A0(ori_ori_n768_), .A1(ori_ori_n81_), .B0(ori_ori_n763_), .Y(ori_ori_n769_));
  NA2        o741(.A(ori_ori_n333_), .B(ori_ori_n766_), .Y(ori_ori_n770_));
  NA4        o742(.A(ori_ori_n770_), .B(ori_ori_n769_), .C(ori_ori_n761_), .D(ori_ori_n758_), .Y(ori00));
  NA2        o743(.A(ori_ori_n377_), .B(f), .Y(ori_ori_n772_));
  NA2        o744(.A(ori_ori_n716_), .B(ori_ori_n464_), .Y(ori_ori_n773_));
  NA3        o745(.A(ori_ori_n773_), .B(ori_ori_n200_), .C(n), .Y(ori_ori_n774_));
  AOI210     o746(.A0(ori_ori_n774_), .A1(ori_ori_n772_), .B0(ori_ori_n737_), .Y(ori_ori_n775_));
  NO2        o747(.A(ori_ori_n775_), .B(ori_ori_n518_), .Y(ori_ori_n776_));
  NA2        o748(.A(d), .B(b), .Y(ori_ori_n777_));
  NO4        o749(.A(ori_ori_n360_), .B(ori_ori_n937_), .C(ori_ori_n759_), .D(ori_ori_n44_), .Y(ori_ori_n778_));
  NA3        o750(.A(ori_ori_n284_), .B(ori_ori_n174_), .C(o), .Y(ori_ori_n779_));
  OR2        o751(.A(ori_ori_n779_), .B(ori_ori_n777_), .Y(ori_ori_n780_));
  NO2        o752(.A(h), .B(o), .Y(ori_ori_n781_));
  NA4        o753(.A(ori_ori_n368_), .B(ori_ori_n352_), .C(ori_ori_n781_), .D(b), .Y(ori_ori_n782_));
  AOI220     o754(.A0(ori_ori_n233_), .A1(ori_ori_n192_), .B0(ori_ori_n131_), .B1(ori_ori_n109_), .Y(ori_ori_n783_));
  NA3        o755(.A(ori_ori_n783_), .B(ori_ori_n782_), .C(ori_ori_n780_), .Y(ori_ori_n784_));
  NO3        o756(.A(ori_ori_n784_), .B(ori_ori_n778_), .C(ori_ori_n207_), .Y(ori_ori_n785_));
  NA2        o757(.A(ori_ori_n192_), .B(ori_ori_n258_), .Y(ori_ori_n786_));
  NA2        o758(.A(ori_ori_n786_), .B(ori_ori_n115_), .Y(ori_ori_n787_));
  NO2        o759(.A(ori_ori_n186_), .B(ori_ori_n135_), .Y(ori_ori_n788_));
  NA2        o760(.A(ori_ori_n788_), .B(ori_ori_n314_), .Y(ori_ori_n789_));
  INV        o761(.A(ori_ori_n789_), .Y(ori_ori_n790_));
  NO3        o762(.A(ori_ori_n790_), .B(ori_ori_n787_), .C(ori_ori_n384_), .Y(ori_ori_n791_));
  AN2        o763(.A(ori_ori_n791_), .B(ori_ori_n785_), .Y(ori_ori_n792_));
  NA3        o764(.A(ori_ori_n755_), .B(ori_ori_n439_), .C(h), .Y(ori_ori_n793_));
  INV        o765(.A(ori_ori_n793_), .Y(ori_ori_n794_));
  NA2        o766(.A(ori_ori_n752_), .B(ori_ori_n397_), .Y(ori_ori_n795_));
  NA4        o767(.A(ori_ori_n467_), .B(ori_ori_n160_), .C(ori_ori_n174_), .D(ori_ori_n123_), .Y(ori_ori_n796_));
  NA2        o768(.A(ori_ori_n796_), .B(ori_ori_n795_), .Y(ori_ori_n797_));
  NO2        o769(.A(ori_ori_n170_), .B(ori_ori_n167_), .Y(ori_ori_n798_));
  NA2        o770(.A(n), .B(e), .Y(ori_ori_n799_));
  NO2        o771(.A(ori_ori_n799_), .B(ori_ori_n108_), .Y(ori_ori_n800_));
  AOI220     o772(.A0(ori_ori_n800_), .A1(ori_ori_n210_), .B0(ori_ori_n592_), .B1(ori_ori_n798_), .Y(ori_ori_n801_));
  OAI210     o773(.A0(ori_ori_n123_), .A1(o), .B0(ori_ori_n334_), .Y(ori_ori_n802_));
  NA2        o774(.A(ori_ori_n802_), .B(ori_ori_n801_), .Y(ori_ori_n803_));
  NA2        o775(.A(ori_ori_n800_), .B(ori_ori_n596_), .Y(ori_ori_n804_));
  AOI220     o776(.A0(ori_ori_n673_), .A1(ori_ori_n422_), .B0(ori_ori_n467_), .B1(ori_ori_n189_), .Y(ori_ori_n805_));
  NA3        o777(.A(ori_ori_n805_), .B(ori_ori_n804_), .C(ori_ori_n608_), .Y(ori_ori_n806_));
  NO4        o778(.A(ori_ori_n806_), .B(ori_ori_n803_), .C(ori_ori_n797_), .D(ori_ori_n794_), .Y(ori_ori_n807_));
  NA3        o779(.A(ori_ori_n807_), .B(ori_ori_n792_), .C(ori_ori_n776_), .Y(ori01));
  NO2        o780(.A(ori_ori_n354_), .B(ori_ori_n212_), .Y(ori_ori_n809_));
  NA2        o781(.A(ori_ori_n295_), .B(i), .Y(ori_ori_n810_));
  NA3        o782(.A(ori_ori_n810_), .B(ori_ori_n809_), .C(ori_ori_n727_), .Y(ori_ori_n811_));
  NA2        o783(.A(ori_ori_n34_), .B(f), .Y(ori_ori_n812_));
  NA2        o784(.A(ori_ori_n513_), .B(o), .Y(ori_ori_n813_));
  NO2        o785(.A(ori_ori_n813_), .B(ori_ori_n812_), .Y(ori_ori_n814_));
  INV        o786(.A(ori_ori_n85_), .Y(ori_ori_n815_));
  OA220      o787(.A0(ori_ori_n815_), .A1(ori_ori_n429_), .B0(ori_ori_n478_), .B1(ori_ori_n274_), .Y(ori_ori_n816_));
  NAi41      o788(.An(ori_ori_n122_), .B(ori_ori_n816_), .C(ori_ori_n796_), .D(ori_ori_n627_), .Y(ori_ori_n817_));
  INV        o789(.A(ori_ori_n484_), .Y(ori_ori_n818_));
  NA3        o790(.A(ori_ori_n513_), .B(o), .C(ori_ori_n166_), .Y(ori_ori_n819_));
  OR2        o791(.A(ori_ori_n149_), .B(ori_ori_n147_), .Y(ori_ori_n820_));
  NA2        o792(.A(ori_ori_n820_), .B(ori_ori_n818_), .Y(ori_ori_n821_));
  NO4        o793(.A(ori_ori_n821_), .B(ori_ori_n817_), .C(ori_ori_n677_), .D(ori_ori_n811_), .Y(ori_ori_n822_));
  NA2        o794(.A(ori_ori_n434_), .B(ori_ori_n85_), .Y(ori_ori_n823_));
  INV        o795(.A(ori_ori_n823_), .Y(ori_ori_n824_));
  OAI210     o796(.A0(ori_ori_n814_), .A1(ori_ori_n241_), .B0(ori_ori_n485_), .Y(ori_ori_n825_));
  INV        o797(.A(ori_ori_n825_), .Y(ori_ori_n826_));
  NO2        o798(.A(ori_ori_n826_), .B(ori_ori_n824_), .Y(ori_ori_n827_));
  NO2        o799(.A(n), .B(ori_ori_n158_), .Y(ori_ori_n828_));
  AOI210     o800(.A0(ori_ori_n374_), .A1(b), .B0(ori_ori_n828_), .Y(ori_ori_n829_));
  OR3        o801(.A(ori_ori_n813_), .B(ori_ori_n438_), .C(ori_ori_n812_), .Y(ori_ori_n830_));
  NO2        o802(.A(ori_ori_n819_), .B(ori_ori_n694_), .Y(ori_ori_n831_));
  NO2        o803(.A(ori_ori_n161_), .B(ori_ori_n79_), .Y(ori_ori_n832_));
  NO2        o804(.A(ori_ori_n832_), .B(ori_ori_n831_), .Y(ori_ori_n833_));
  NA4        o805(.A(ori_ori_n833_), .B(ori_ori_n830_), .C(ori_ori_n829_), .D(ori_ori_n544_), .Y(ori_ori_n834_));
  NO2        o806(.A(ori_ori_n683_), .B(ori_ori_n181_), .Y(ori_ori_n835_));
  NO2        o807(.A(ori_ori_n684_), .B(ori_ori_n410_), .Y(ori_ori_n836_));
  OAI210     o808(.A0(ori_ori_n836_), .A1(ori_ori_n835_), .B0(ori_ori_n254_), .Y(ori_ori_n837_));
  NA2        o809(.A(ori_ori_n417_), .B(ori_ori_n415_), .Y(ori_ori_n838_));
  NO3        o810(.A(ori_ori_n55_), .B(ori_ori_n221_), .C(ori_ori_n34_), .Y(ori_ori_n839_));
  NA2        o811(.A(ori_ori_n839_), .B(ori_ori_n407_), .Y(ori_ori_n840_));
  NA3        o812(.A(ori_ori_n840_), .B(ori_ori_n838_), .C(ori_ori_n481_), .Y(ori_ori_n841_));
  NO2        o813(.A(ori_ori_n274_), .B(ori_ori_n48_), .Y(ori_ori_n842_));
  INV        o814(.A(ori_ori_n842_), .Y(ori_ori_n843_));
  NA2        o815(.A(ori_ori_n839_), .B(ori_ori_n577_), .Y(ori_ori_n844_));
  NA3        o816(.A(ori_ori_n844_), .B(ori_ori_n843_), .C(ori_ori_n287_), .Y(ori_ori_n845_));
  NOi41      o817(.An(ori_ori_n837_), .B(ori_ori_n845_), .C(ori_ori_n841_), .D(ori_ori_n834_), .Y(ori_ori_n846_));
  NO2        o818(.A(ori_ori_n94_), .B(ori_ori_n34_), .Y(ori_ori_n847_));
  AO220      o819(.A0(i), .A1(ori_ori_n450_), .B0(ori_ori_n847_), .B1(ori_ori_n511_), .Y(ori_ori_n848_));
  NA2        o820(.A(ori_ori_n848_), .B(ori_ori_n254_), .Y(ori_ori_n849_));
  INV        o821(.A(ori_ori_n97_), .Y(ori_ori_n850_));
  NO3        o822(.A(ori_ori_n745_), .B(ori_ori_n130_), .C(ori_ori_n62_), .Y(ori_ori_n851_));
  AOI220     o823(.A0(ori_ori_n851_), .A1(ori_ori_n850_), .B0(ori_ori_n839_), .B1(ori_ori_n685_), .Y(ori_ori_n852_));
  NA2        o824(.A(ori_ori_n852_), .B(ori_ori_n849_), .Y(ori_ori_n853_));
  NO2        o825(.A(ori_ori_n444_), .B(ori_ori_n443_), .Y(ori_ori_n854_));
  NO4        o826(.A(ori_ori_n745_), .B(ori_ori_n854_), .C(ori_ori_n128_), .D(ori_ori_n62_), .Y(ori_ori_n855_));
  NO3        o827(.A(ori_ori_n855_), .B(ori_ori_n853_), .C(ori_ori_n460_), .Y(ori_ori_n856_));
  NA4        o828(.A(ori_ori_n856_), .B(ori_ori_n846_), .C(ori_ori_n827_), .D(ori_ori_n822_), .Y(ori06));
  NO2        o829(.A(ori_ori_n176_), .B(ori_ori_n72_), .Y(ori_ori_n858_));
  OAI210     o830(.A0(ori_ori_n858_), .A1(ori_ori_n851_), .B0(ori_ori_n283_), .Y(ori_ori_n859_));
  NA2        o831(.A(ori_ori_n859_), .B(ori_ori_n837_), .Y(ori_ori_n860_));
  NO3        o832(.A(ori_ori_n860_), .B(ori_ori_n841_), .C(ori_ori_n199_), .Y(ori_ori_n861_));
  NA2        o833(.A(i), .B(ori_ori_n686_), .Y(ori_ori_n862_));
  AOI210     o834(.A0(i), .A1(ori_ori_n411_), .B0(ori_ori_n848_), .Y(ori_ori_n863_));
  AOI210     o835(.A0(ori_ori_n863_), .A1(ori_ori_n862_), .B0(ori_ori_n251_), .Y(ori_ori_n864_));
  INV        o836(.A(ori_ori_n64_), .Y(ori_ori_n865_));
  NA2        o837(.A(ori_ori_n865_), .B(ori_ori_n268_), .Y(ori_ori_n866_));
  NO2        o838(.A(ori_ori_n381_), .B(ori_ori_n125_), .Y(ori_ori_n867_));
  NO2        o839(.A(ori_ori_n440_), .B(ori_ori_n756_), .Y(ori_ori_n868_));
  INV        o840(.A(ori_ori_n633_), .Y(ori_ori_n869_));
  NO3        o841(.A(ori_ori_n869_), .B(ori_ori_n868_), .C(ori_ori_n867_), .Y(ori_ori_n870_));
  NA2        o842(.A(ori_ori_n870_), .B(ori_ori_n866_), .Y(ori_ori_n871_));
  AN2        o843(.A(ori_ori_n673_), .B(ori_ori_n463_), .Y(ori_ori_n872_));
  NO3        o844(.A(ori_ori_n872_), .B(ori_ori_n871_), .C(ori_ori_n864_), .Y(ori_ori_n873_));
  NO3        o845(.A(ori_ori_n188_), .B(ori_ori_n72_), .C(ori_ori_n214_), .Y(ori_ori_n874_));
  INV        o846(.A(k), .Y(ori_ori_n875_));
  NO3        o847(.A(ori_ori_n875_), .B(ori_ori_n436_), .C(j), .Y(ori_ori_n876_));
  NOi21      o848(.An(ori_ori_n876_), .B(ori_ori_n480_), .Y(ori_ori_n877_));
  NO3        o849(.A(ori_ori_n877_), .B(ori_ori_n874_), .C(ori_ori_n757_), .Y(ori_ori_n878_));
  NA2        o850(.A(ori_ori_n878_), .B(ori_ori_n805_), .Y(ori_ori_n879_));
  NA2        o851(.A(ori_ori_n417_), .B(ori_ori_n334_), .Y(ori_ori_n880_));
  NA2        o852(.A(ori_ori_n876_), .B(ori_ori_n567_), .Y(ori_ori_n881_));
  NA2        o853(.A(ori_ori_n881_), .B(ori_ori_n880_), .Y(ori_ori_n882_));
  AN2        o854(.A(ori_ori_n649_), .B(ori_ori_n648_), .Y(ori_ori_n883_));
  NO4        o855(.A(ori_ori_n883_), .B(ori_ori_n616_), .C(ori_ori_n370_), .D(ori_ori_n355_), .Y(ori_ori_n884_));
  NA2        o856(.A(ori_ori_n884_), .B(ori_ori_n844_), .Y(ori_ori_n885_));
  NAi21      o857(.An(j), .B(i), .Y(ori_ori_n886_));
  NO4        o858(.A(ori_ori_n854_), .B(ori_ori_n886_), .C(ori_ori_n329_), .D(ori_ori_n183_), .Y(ori_ori_n887_));
  NO4        o859(.A(ori_ori_n887_), .B(ori_ori_n885_), .C(ori_ori_n882_), .D(ori_ori_n879_), .Y(ori_ori_n888_));
  NA4        o860(.A(ori_ori_n888_), .B(ori_ori_n873_), .C(ori_ori_n861_), .D(ori_ori_n856_), .Y(ori07));
  NOi31      o861(.An(n), .B(m), .C(b), .Y(ori_ori_n890_));
  NO3        o862(.A(ori_ori_n95_), .B(ori_ori_n335_), .C(h), .Y(ori_ori_n891_));
  NO2        o863(.A(ori_ori_n738_), .B(ori_ori_n329_), .Y(ori_ori_n892_));
  INV        o864(.A(ori_ori_n892_), .Y(ori_ori_n893_));
  NO2        o865(.A(ori_ori_n739_), .B(ori_ori_n225_), .Y(ori_ori_n894_));
  INV        o866(.A(ori_ori_n893_), .Y(ori_ori_n895_));
  INV        o867(.A(ori_ori_n895_), .Y(ori_ori_n896_));
  NO3        o868(.A(ori_ori_n329_), .B(d), .C(c), .Y(ori_ori_n897_));
  NA2        o869(.A(ori_ori_n743_), .B(ori_ori_n352_), .Y(ori_ori_n898_));
  NO2        o870(.A(ori_ori_n898_), .B(ori_ori_n329_), .Y(ori_ori_n899_));
  INV        o871(.A(ori_ori_n899_), .Y(ori_ori_n900_));
  NA2        o872(.A(ori_ori_n890_), .B(ori_ori_n280_), .Y(ori_ori_n901_));
  INV        o873(.A(ori_ori_n901_), .Y(ori_ori_n902_));
  INV        o874(.A(ori_ori_n746_), .Y(ori_ori_n903_));
  NAi21      o875(.An(ori_ori_n902_), .B(ori_ori_n903_), .Y(ori_ori_n904_));
  NO4        o876(.A(ori_ori_n95_), .B(o), .C(f), .D(e), .Y(ori_ori_n905_));
  INV        o877(.A(ori_ori_n904_), .Y(ori_ori_n906_));
  NA3        o878(.A(ori_ori_n906_), .B(ori_ori_n900_), .C(ori_ori_n896_), .Y(ori_ori_n907_));
  NO2        o879(.A(ori_ori_n292_), .B(j), .Y(ori_ori_n908_));
  NA2        o880(.A(ori_ori_n741_), .B(ori_ori_n111_), .Y(ori_ori_n909_));
  INV        o881(.A(ori_ori_n909_), .Y(ori_ori_n910_));
  NA2        o882(.A(ori_ori_n908_), .B(ori_ori_n119_), .Y(ori_ori_n911_));
  INV        o883(.A(ori_ori_n911_), .Y(ori_ori_n912_));
  NO2        o884(.A(ori_ori_n912_), .B(ori_ori_n910_), .Y(ori_ori_n913_));
  NO2        o885(.A(ori_ori_n176_), .B(ori_ori_n130_), .Y(ori_ori_n914_));
  NO2        o886(.A(ori_ori_n742_), .B(h), .Y(ori_ori_n915_));
  NO2        o887(.A(ori_ori_n886_), .B(ori_ori_n128_), .Y(ori_ori_n916_));
  NA2        o888(.A(h), .B(ori_ori_n916_), .Y(ori_ori_n917_));
  INV        o889(.A(ori_ori_n917_), .Y(ori_ori_n918_));
  NO3        o890(.A(ori_ori_n918_), .B(ori_ori_n81_), .C(ori_ori_n915_), .Y(ori_ori_n919_));
  NA3        o891(.A(ori_ori_n919_), .B(ori_ori_n933_), .C(ori_ori_n913_), .Y(ori_ori_n920_));
  NA2        o892(.A(h), .B(ori_ori_n894_), .Y(ori_ori_n921_));
  OAI210     o893(.A0(ori_ori_n905_), .A1(ori_ori_n890_), .B0(ori_ori_n619_), .Y(ori_ori_n922_));
  NA2        o894(.A(ori_ori_n922_), .B(ori_ori_n921_), .Y(ori_ori_n923_));
  INV        o895(.A(ori_ori_n923_), .Y(ori_ori_n924_));
  OR2        o896(.A(h), .B(ori_ori_n398_), .Y(ori_ori_n925_));
  NO2        o897(.A(ori_ori_n925_), .B(ori_ori_n128_), .Y(ori_ori_n926_));
  NO3        o898(.A(ori_ori_n747_), .B(ori_ori_n926_), .C(ori_ori_n897_), .Y(ori_ori_n927_));
  NA2        o899(.A(ori_ori_n927_), .B(ori_ori_n924_), .Y(ori_ori_n928_));
  OR4        o900(.A(ori_ori_n891_), .B(ori_ori_n928_), .C(ori_ori_n920_), .D(ori_ori_n907_), .Y(ori04));
  INV        o901(.A(ori_ori_n68_), .Y(ori_ori_n932_));
  INV        o902(.A(ori_ori_n914_), .Y(ori_ori_n933_));
  INV        o903(.A(e), .Y(ori_ori_n934_));
  INV        o904(.A(ori_ori_n433_), .Y(ori_ori_n935_));
  INV        o905(.A(e), .Y(ori_ori_n936_));
  INV        o906(.A(h), .Y(ori_ori_n937_));
  ZERO       o907(.Y(ori02));
  ZERO       o908(.Y(ori03));
  ZERO       o909(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA2        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(m), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(m), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(m), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(m), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(m), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO4        m0025(.A(mai_mai_n53_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NAi21      m0031(.An(i), .B(h), .Y(mai_mai_n60_));
  NAi31      m0032(.An(i), .B(l), .C(j), .Y(mai_mai_n61_));
  NO2        m0033(.A(mai_mai_n60_), .B(mai_mai_n44_), .Y(mai_mai_n62_));
  NA2        m0034(.A(mai_mai_n62_), .B(mai_mai_n58_), .Y(mai_mai_n63_));
  NAi41      m0035(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n64_));
  NA2        m0036(.A(m), .B(f), .Y(mai_mai_n65_));
  NO2        m0037(.A(mai_mai_n65_), .B(mai_mai_n64_), .Y(mai_mai_n66_));
  NAi21      m0038(.An(i), .B(j), .Y(mai_mai_n67_));
  NAi32      m0039(.An(n), .Bn(k), .C(m), .Y(mai_mai_n68_));
  NAi31      m0040(.An(l), .B(m), .C(k), .Y(mai_mai_n69_));
  NAi21      m0041(.An(e), .B(h), .Y(mai_mai_n70_));
  NAi41      m0042(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n71_));
  INV        m0043(.A(m), .Y(mai_mai_n72_));
  NOi21      m0044(.An(k), .B(l), .Y(mai_mai_n73_));
  AN4        m0045(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n74_));
  NOi31      m0046(.An(h), .B(m), .C(f), .Y(mai_mai_n75_));
  NA2        m0047(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n76_));
  NAi32      m0048(.An(m), .Bn(k), .C(j), .Y(mai_mai_n77_));
  NOi32      m0049(.An(h), .Bn(m), .C(f), .Y(mai_mai_n78_));
  NA2        m0050(.A(mai_mai_n78_), .B(mai_mai_n74_), .Y(mai_mai_n79_));
  OA220      m0051(.A0(mai_mai_n79_), .A1(mai_mai_n77_), .B0(mai_mai_n76_), .B1(l), .Y(mai_mai_n80_));
  NA2        m0052(.A(mai_mai_n80_), .B(mai_mai_n63_), .Y(mai_mai_n81_));
  INV        m0053(.A(n), .Y(mai_mai_n82_));
  NOi32      m0054(.An(e), .Bn(b), .C(d), .Y(mai_mai_n83_));
  NA2        m0055(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n84_));
  INV        m0056(.A(j), .Y(mai_mai_n85_));
  AN3        m0057(.A(m), .B(k), .C(i), .Y(mai_mai_n86_));
  NA3        m0058(.A(mai_mai_n86_), .B(mai_mai_n85_), .C(m), .Y(mai_mai_n87_));
  NAi32      m0059(.An(m), .Bn(f), .C(h), .Y(mai_mai_n88_));
  NAi31      m0060(.An(j), .B(m), .C(l), .Y(mai_mai_n89_));
  NAi31      m0061(.An(k), .B(j), .C(m), .Y(mai_mai_n90_));
  NO2        m0062(.A(mai_mai_n90_), .B(f), .Y(mai_mai_n91_));
  AN2        m0063(.A(j), .B(m), .Y(mai_mai_n92_));
  NOi32      m0064(.An(m), .Bn(l), .C(i), .Y(mai_mai_n93_));
  NOi21      m0065(.An(m), .B(i), .Y(mai_mai_n94_));
  NOi32      m0066(.An(m), .Bn(j), .C(k), .Y(mai_mai_n95_));
  AOI220     m0067(.A0(mai_mai_n95_), .A1(mai_mai_n94_), .B0(mai_mai_n93_), .B1(mai_mai_n92_), .Y(mai_mai_n96_));
  NO2        m0068(.A(mai_mai_n96_), .B(f), .Y(mai_mai_n97_));
  NAi41      m0069(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n98_));
  AN2        m0070(.A(e), .B(b), .Y(mai_mai_n99_));
  NOi31      m0071(.An(c), .B(h), .C(f), .Y(mai_mai_n100_));
  NA2        m0072(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  NOi21      m0073(.An(i), .B(h), .Y(mai_mai_n102_));
  NA3        m0074(.A(mai_mai_n102_), .B(m), .C(mai_mai_n36_), .Y(mai_mai_n103_));
  INV        m0075(.A(a), .Y(mai_mai_n104_));
  NA2        m0076(.A(mai_mai_n99_), .B(mai_mai_n104_), .Y(mai_mai_n105_));
  INV        m0077(.A(l), .Y(mai_mai_n106_));
  NOi21      m0078(.An(m), .B(n), .Y(mai_mai_n107_));
  AN2        m0079(.A(k), .B(h), .Y(mai_mai_n108_));
  NO2        m0080(.A(mai_mai_n103_), .B(mai_mai_n84_), .Y(mai_mai_n109_));
  INV        m0081(.A(b), .Y(mai_mai_n110_));
  NA2        m0082(.A(l), .B(j), .Y(mai_mai_n111_));
  AN2        m0083(.A(k), .B(i), .Y(mai_mai_n112_));
  NA2        m0084(.A(mai_mai_n112_), .B(mai_mai_n111_), .Y(mai_mai_n113_));
  NA2        m0085(.A(m), .B(e), .Y(mai_mai_n114_));
  NOi32      m0086(.An(c), .Bn(a), .C(d), .Y(mai_mai_n115_));
  NA2        m0087(.A(mai_mai_n115_), .B(mai_mai_n107_), .Y(mai_mai_n116_));
  NO3        m0088(.A(mai_mai_n116_), .B(mai_mai_n114_), .C(mai_mai_n113_), .Y(mai_mai_n117_));
  NO2        m0089(.A(mai_mai_n117_), .B(mai_mai_n109_), .Y(mai_mai_n118_));
  OAI210     m0090(.A0(mai_mai_n96_), .A1(mai_mai_n84_), .B0(mai_mai_n118_), .Y(mai_mai_n119_));
  NOi31      m0091(.An(k), .B(m), .C(j), .Y(mai_mai_n120_));
  NOi31      m0092(.An(k), .B(m), .C(i), .Y(mai_mai_n121_));
  NA3        m0093(.A(mai_mai_n121_), .B(mai_mai_n78_), .C(mai_mai_n74_), .Y(mai_mai_n122_));
  INV        m0094(.A(mai_mai_n122_), .Y(mai_mai_n123_));
  NOi32      m0095(.An(f), .Bn(b), .C(e), .Y(mai_mai_n124_));
  NAi21      m0096(.An(m), .B(h), .Y(mai_mai_n125_));
  NAi21      m0097(.An(m), .B(n), .Y(mai_mai_n126_));
  NAi21      m0098(.An(j), .B(k), .Y(mai_mai_n127_));
  NO3        m0099(.A(mai_mai_n127_), .B(mai_mai_n126_), .C(mai_mai_n125_), .Y(mai_mai_n128_));
  NAi41      m0100(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n129_));
  NAi31      m0101(.An(j), .B(k), .C(h), .Y(mai_mai_n130_));
  NO3        m0102(.A(mai_mai_n130_), .B(mai_mai_n129_), .C(mai_mai_n126_), .Y(mai_mai_n131_));
  AOI210     m0103(.A0(mai_mai_n128_), .A1(mai_mai_n124_), .B0(mai_mai_n131_), .Y(mai_mai_n132_));
  NO2        m0104(.A(k), .B(j), .Y(mai_mai_n133_));
  AN2        m0105(.A(k), .B(j), .Y(mai_mai_n134_));
  NA2        m0106(.A(f), .B(d), .Y(mai_mai_n135_));
  NAi31      m0107(.An(f), .B(e), .C(b), .Y(mai_mai_n136_));
  NA2        m0108(.A(d), .B(b), .Y(mai_mai_n137_));
  NAi21      m0109(.An(e), .B(f), .Y(mai_mai_n138_));
  NO2        m0110(.A(mai_mai_n138_), .B(mai_mai_n137_), .Y(mai_mai_n139_));
  NA2        m0111(.A(b), .B(a), .Y(mai_mai_n140_));
  NAi21      m0112(.An(c), .B(d), .Y(mai_mai_n141_));
  NAi21      m0113(.An(mai_mai_n123_), .B(mai_mai_n132_), .Y(mai_mai_n142_));
  NAi31      m0114(.An(e), .B(f), .C(b), .Y(mai_mai_n143_));
  NOi21      m0115(.An(h), .B(i), .Y(mai_mai_n144_));
  NOi21      m0116(.An(k), .B(m), .Y(mai_mai_n145_));
  NA3        m0117(.A(mai_mai_n145_), .B(mai_mai_n144_), .C(n), .Y(mai_mai_n146_));
  NOi21      m0118(.An(h), .B(m), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n135_), .B(c), .Y(mai_mai_n148_));
  NA2        m0120(.A(mai_mai_n148_), .B(mai_mai_n147_), .Y(mai_mai_n149_));
  NAi31      m0121(.An(l), .B(j), .C(h), .Y(mai_mai_n150_));
  NO2        m0122(.A(mai_mai_n150_), .B(mai_mai_n49_), .Y(mai_mai_n151_));
  NA2        m0123(.A(mai_mai_n151_), .B(mai_mai_n66_), .Y(mai_mai_n152_));
  NOi32      m0124(.An(n), .Bn(k), .C(m), .Y(mai_mai_n153_));
  NA2        m0125(.A(l), .B(i), .Y(mai_mai_n154_));
  NA2        m0126(.A(mai_mai_n154_), .B(mai_mai_n153_), .Y(mai_mai_n155_));
  OAI210     m0127(.A0(mai_mai_n155_), .A1(mai_mai_n149_), .B0(mai_mai_n152_), .Y(mai_mai_n156_));
  NAi31      m0128(.An(e), .B(f), .C(c), .Y(mai_mai_n157_));
  NA2        m0129(.A(j), .B(h), .Y(mai_mai_n158_));
  OR3        m0130(.A(n), .B(m), .C(k), .Y(mai_mai_n159_));
  NAi32      m0131(.An(m), .Bn(k), .C(n), .Y(mai_mai_n160_));
  NO2        m0132(.A(n), .B(m), .Y(mai_mai_n161_));
  NA2        m0133(.A(mai_mai_n161_), .B(mai_mai_n50_), .Y(mai_mai_n162_));
  NAi21      m0134(.An(f), .B(e), .Y(mai_mai_n163_));
  NA2        m0135(.A(d), .B(c), .Y(mai_mai_n164_));
  NO2        m0136(.A(mai_mai_n164_), .B(mai_mai_n163_), .Y(mai_mai_n165_));
  NOi21      m0137(.An(mai_mai_n165_), .B(mai_mai_n162_), .Y(mai_mai_n166_));
  NAi21      m0138(.An(d), .B(c), .Y(mai_mai_n167_));
  NAi31      m0139(.An(m), .B(n), .C(b), .Y(mai_mai_n168_));
  NA2        m0140(.A(k), .B(i), .Y(mai_mai_n169_));
  NAi21      m0141(.An(h), .B(f), .Y(mai_mai_n170_));
  NO2        m0142(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n171_));
  NO2        m0143(.A(mai_mai_n168_), .B(mai_mai_n141_), .Y(mai_mai_n172_));
  NA2        m0144(.A(mai_mai_n172_), .B(mai_mai_n171_), .Y(mai_mai_n173_));
  NOi32      m0145(.An(f), .Bn(c), .C(e), .Y(mai_mai_n174_));
  NO3        m0146(.A(n), .B(m), .C(j), .Y(mai_mai_n175_));
  NA2        m0147(.A(mai_mai_n175_), .B(mai_mai_n108_), .Y(mai_mai_n176_));
  NAi21      m0148(.An(mai_mai_n166_), .B(mai_mai_n173_), .Y(mai_mai_n177_));
  OR3        m0149(.A(mai_mai_n177_), .B(mai_mai_n156_), .C(mai_mai_n142_), .Y(mai_mai_n178_));
  NO4        m0150(.A(mai_mai_n178_), .B(mai_mai_n119_), .C(mai_mai_n81_), .D(mai_mai_n55_), .Y(mai_mai_n179_));
  NA3        m0151(.A(m), .B(mai_mai_n106_), .C(j), .Y(mai_mai_n180_));
  NAi31      m0152(.An(n), .B(h), .C(m), .Y(mai_mai_n181_));
  NO2        m0153(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  NOi32      m0154(.An(m), .Bn(k), .C(l), .Y(mai_mai_n183_));
  NA3        m0155(.A(mai_mai_n183_), .B(mai_mai_n85_), .C(m), .Y(mai_mai_n184_));
  NO2        m0156(.A(mai_mai_n184_), .B(n), .Y(mai_mai_n185_));
  AN2        m0157(.A(i), .B(m), .Y(mai_mai_n186_));
  NA3        m0158(.A(mai_mai_n73_), .B(mai_mai_n186_), .C(mai_mai_n107_), .Y(mai_mai_n187_));
  INV        m0159(.A(mai_mai_n187_), .Y(mai_mai_n188_));
  NAi31      m0160(.An(d), .B(n), .C(e), .Y(mai_mai_n189_));
  INV        m0161(.A(mai_mai_n189_), .Y(mai_mai_n190_));
  INV        m0162(.A(f), .Y(mai_mai_n191_));
  INV        m0163(.A(m), .Y(mai_mai_n192_));
  NOi31      m0164(.An(i), .B(j), .C(h), .Y(mai_mai_n193_));
  NOi21      m0165(.An(l), .B(m), .Y(mai_mai_n194_));
  NA2        m0166(.A(mai_mai_n194_), .B(mai_mai_n193_), .Y(mai_mai_n195_));
  NO2        m0167(.A(mai_mai_n187_), .B(mai_mai_n32_), .Y(mai_mai_n196_));
  NOi21      m0168(.An(n), .B(m), .Y(mai_mai_n197_));
  NOi32      m0169(.An(l), .Bn(i), .C(j), .Y(mai_mai_n198_));
  NA2        m0170(.A(mai_mai_n198_), .B(mai_mai_n197_), .Y(mai_mai_n199_));
  OA220      m0171(.A0(mai_mai_n199_), .A1(mai_mai_n101_), .B0(mai_mai_n77_), .B1(mai_mai_n76_), .Y(mai_mai_n200_));
  NAi21      m0172(.An(j), .B(h), .Y(mai_mai_n201_));
  XN2        m0173(.A(i), .B(h), .Y(mai_mai_n202_));
  NA2        m0174(.A(mai_mai_n202_), .B(mai_mai_n201_), .Y(mai_mai_n203_));
  NOi31      m0175(.An(k), .B(n), .C(m), .Y(mai_mai_n204_));
  NOi31      m0176(.An(mai_mai_n204_), .B(mai_mai_n164_), .C(mai_mai_n163_), .Y(mai_mai_n205_));
  NA2        m0177(.A(mai_mai_n205_), .B(mai_mai_n203_), .Y(mai_mai_n206_));
  NAi31      m0178(.An(f), .B(e), .C(c), .Y(mai_mai_n207_));
  NO3        m0179(.A(mai_mai_n207_), .B(mai_mai_n159_), .C(mai_mai_n158_), .Y(mai_mai_n208_));
  NA4        m0180(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n209_));
  NAi32      m0181(.An(m), .Bn(i), .C(k), .Y(mai_mai_n210_));
  NO3        m0182(.A(mai_mai_n210_), .B(mai_mai_n88_), .C(mai_mai_n209_), .Y(mai_mai_n211_));
  NO2        m0183(.A(mai_mai_n211_), .B(mai_mai_n208_), .Y(mai_mai_n212_));
  NAi21      m0184(.An(n), .B(a), .Y(mai_mai_n213_));
  NO2        m0185(.A(mai_mai_n213_), .B(mai_mai_n137_), .Y(mai_mai_n214_));
  NAi41      m0186(.An(m), .B(m), .C(k), .D(h), .Y(mai_mai_n215_));
  NO2        m0187(.A(mai_mai_n215_), .B(e), .Y(mai_mai_n216_));
  NO2        m0188(.A(mai_mai_n138_), .B(mai_mai_n90_), .Y(mai_mai_n217_));
  OAI210     m0189(.A0(mai_mai_n217_), .A1(mai_mai_n216_), .B0(mai_mai_n214_), .Y(mai_mai_n218_));
  AN4        m0190(.A(mai_mai_n218_), .B(mai_mai_n212_), .C(mai_mai_n206_), .D(mai_mai_n200_), .Y(mai_mai_n219_));
  OR2        m0191(.A(h), .B(m), .Y(mai_mai_n220_));
  NO2        m0192(.A(mai_mai_n220_), .B(mai_mai_n98_), .Y(mai_mai_n221_));
  NA2        m0193(.A(mai_mai_n221_), .B(mai_mai_n124_), .Y(mai_mai_n222_));
  NA2        m0194(.A(mai_mai_n145_), .B(mai_mai_n102_), .Y(mai_mai_n223_));
  NO2        m0195(.A(n), .B(a), .Y(mai_mai_n224_));
  NAi31      m0196(.An(mai_mai_n215_), .B(mai_mai_n224_), .C(mai_mai_n99_), .Y(mai_mai_n225_));
  NAi21      m0197(.An(h), .B(i), .Y(mai_mai_n226_));
  NA2        m0198(.A(mai_mai_n161_), .B(k), .Y(mai_mai_n227_));
  NO2        m0199(.A(mai_mai_n227_), .B(mai_mai_n226_), .Y(mai_mai_n228_));
  NA2        m0200(.A(mai_mai_n225_), .B(mai_mai_n222_), .Y(mai_mai_n229_));
  NOi21      m0201(.An(m), .B(e), .Y(mai_mai_n230_));
  NO2        m0202(.A(mai_mai_n71_), .B(mai_mai_n72_), .Y(mai_mai_n231_));
  NA2        m0203(.A(mai_mai_n231_), .B(mai_mai_n230_), .Y(mai_mai_n232_));
  NOi32      m0204(.An(l), .Bn(j), .C(i), .Y(mai_mai_n233_));
  AOI210     m0205(.A0(mai_mai_n73_), .A1(mai_mai_n85_), .B0(mai_mai_n233_), .Y(mai_mai_n234_));
  NO2        m0206(.A(mai_mai_n226_), .B(mai_mai_n44_), .Y(mai_mai_n235_));
  NAi21      m0207(.An(f), .B(m), .Y(mai_mai_n236_));
  NO2        m0208(.A(mai_mai_n236_), .B(mai_mai_n64_), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n68_), .B(mai_mai_n111_), .Y(mai_mai_n238_));
  AOI220     m0210(.A0(mai_mai_n238_), .A1(mai_mai_n237_), .B0(mai_mai_n235_), .B1(mai_mai_n66_), .Y(mai_mai_n239_));
  OAI210     m0211(.A0(mai_mai_n234_), .A1(mai_mai_n232_), .B0(mai_mai_n239_), .Y(mai_mai_n240_));
  NO3        m0212(.A(mai_mai_n127_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n241_));
  NOi41      m0213(.An(mai_mai_n219_), .B(mai_mai_n240_), .C(mai_mai_n229_), .D(mai_mai_n196_), .Y(mai_mai_n242_));
  NO4        m0214(.A(mai_mai_n182_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n243_));
  NO2        m0215(.A(mai_mai_n243_), .B(mai_mai_n105_), .Y(mai_mai_n244_));
  NAi21      m0216(.An(h), .B(m), .Y(mai_mai_n245_));
  OR4        m0217(.A(mai_mai_n245_), .B(mai_mai_n1281_), .C(mai_mai_n199_), .D(e), .Y(mai_mai_n246_));
  NO2        m0218(.A(mai_mai_n223_), .B(mai_mai_n236_), .Y(mai_mai_n247_));
  NA2        m0219(.A(mai_mai_n247_), .B(mai_mai_n74_), .Y(mai_mai_n248_));
  NAi31      m0220(.An(m), .B(k), .C(h), .Y(mai_mai_n249_));
  NO3        m0221(.A(mai_mai_n126_), .B(mai_mai_n249_), .C(l), .Y(mai_mai_n250_));
  NAi31      m0222(.An(e), .B(d), .C(a), .Y(mai_mai_n251_));
  NA2        m0223(.A(mai_mai_n250_), .B(mai_mai_n124_), .Y(mai_mai_n252_));
  NA3        m0224(.A(mai_mai_n252_), .B(mai_mai_n248_), .C(mai_mai_n246_), .Y(mai_mai_n253_));
  NA3        m0225(.A(mai_mai_n145_), .B(mai_mai_n144_), .C(mai_mai_n82_), .Y(mai_mai_n254_));
  NA3        m0226(.A(e), .B(c), .C(b), .Y(mai_mai_n255_));
  NAi32      m0227(.An(k), .Bn(i), .C(j), .Y(mai_mai_n256_));
  NA2        m0228(.A(mai_mai_n256_), .B(mai_mai_n150_), .Y(mai_mai_n257_));
  NOi21      m0229(.An(mai_mai_n257_), .B(mai_mai_n49_), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n237_), .B(mai_mai_n258_), .Y(mai_mai_n259_));
  NAi21      m0231(.An(l), .B(k), .Y(mai_mai_n260_));
  NO2        m0232(.A(mai_mai_n260_), .B(mai_mai_n49_), .Y(mai_mai_n261_));
  NOi21      m0233(.An(l), .B(j), .Y(mai_mai_n262_));
  NA2        m0234(.A(mai_mai_n147_), .B(mai_mai_n262_), .Y(mai_mai_n263_));
  NA2        m0235(.A(mai_mai_n112_), .B(m), .Y(mai_mai_n264_));
  OR3        m0236(.A(mai_mai_n71_), .B(mai_mai_n72_), .C(e), .Y(mai_mai_n265_));
  AOI210     m0237(.A0(mai_mai_n264_), .A1(mai_mai_n263_), .B0(mai_mai_n265_), .Y(mai_mai_n266_));
  INV        m0238(.A(mai_mai_n266_), .Y(mai_mai_n267_));
  NAi32      m0239(.An(j), .Bn(h), .C(i), .Y(mai_mai_n268_));
  NAi21      m0240(.An(m), .B(l), .Y(mai_mai_n269_));
  NO3        m0241(.A(mai_mai_n269_), .B(mai_mai_n268_), .C(mai_mai_n82_), .Y(mai_mai_n270_));
  NA2        m0242(.A(h), .B(m), .Y(mai_mai_n271_));
  NA2        m0243(.A(mai_mai_n153_), .B(mai_mai_n45_), .Y(mai_mai_n272_));
  NO2        m0244(.A(mai_mai_n272_), .B(mai_mai_n271_), .Y(mai_mai_n273_));
  OAI210     m0245(.A0(mai_mai_n273_), .A1(mai_mai_n270_), .B0(mai_mai_n148_), .Y(mai_mai_n274_));
  NA3        m0246(.A(mai_mai_n274_), .B(mai_mai_n267_), .C(mai_mai_n259_), .Y(mai_mai_n275_));
  NO2        m0247(.A(mai_mai_n136_), .B(d), .Y(mai_mai_n276_));
  NA2        m0248(.A(mai_mai_n276_), .B(mai_mai_n53_), .Y(mai_mai_n277_));
  NO2        m0249(.A(mai_mai_n101_), .B(mai_mai_n98_), .Y(mai_mai_n278_));
  NAi32      m0250(.An(n), .Bn(m), .C(l), .Y(mai_mai_n279_));
  NO2        m0251(.A(mai_mai_n279_), .B(mai_mai_n268_), .Y(mai_mai_n280_));
  NA2        m0252(.A(mai_mai_n280_), .B(mai_mai_n165_), .Y(mai_mai_n281_));
  NO2        m0253(.A(mai_mai_n116_), .B(mai_mai_n110_), .Y(mai_mai_n282_));
  NAi31      m0254(.An(k), .B(l), .C(j), .Y(mai_mai_n283_));
  OAI210     m0255(.A0(mai_mai_n260_), .A1(j), .B0(mai_mai_n283_), .Y(mai_mai_n284_));
  NOi21      m0256(.An(mai_mai_n284_), .B(mai_mai_n114_), .Y(mai_mai_n285_));
  NA2        m0257(.A(mai_mai_n285_), .B(mai_mai_n282_), .Y(mai_mai_n286_));
  NA3        m0258(.A(mai_mai_n286_), .B(mai_mai_n281_), .C(mai_mai_n277_), .Y(mai_mai_n287_));
  NO4        m0259(.A(mai_mai_n287_), .B(mai_mai_n275_), .C(mai_mai_n253_), .D(mai_mai_n244_), .Y(mai_mai_n288_));
  NA2        m0260(.A(mai_mai_n228_), .B(mai_mai_n174_), .Y(mai_mai_n289_));
  NAi21      m0261(.An(m), .B(k), .Y(mai_mai_n290_));
  NAi41      m0262(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n291_));
  NAi31      m0263(.An(i), .B(l), .C(h), .Y(mai_mai_n292_));
  NO3        m0264(.A(mai_mai_n292_), .B(mai_mai_n71_), .C(mai_mai_n72_), .Y(mai_mai_n293_));
  NA2        m0265(.A(f), .B(mai_mai_n112_), .Y(mai_mai_n294_));
  NO2        m0266(.A(mai_mai_n294_), .B(mai_mai_n192_), .Y(mai_mai_n295_));
  NAi31      m0267(.An(d), .B(e), .C(b), .Y(mai_mai_n296_));
  NO2        m0268(.A(mai_mai_n126_), .B(mai_mai_n296_), .Y(mai_mai_n297_));
  NA2        m0269(.A(mai_mai_n297_), .B(mai_mai_n295_), .Y(mai_mai_n298_));
  NAi31      m0270(.An(mai_mai_n293_), .B(mai_mai_n298_), .C(mai_mai_n289_), .Y(mai_mai_n299_));
  NO4        m0271(.A(mai_mai_n291_), .B(mai_mai_n77_), .C(mai_mai_n70_), .D(mai_mai_n192_), .Y(mai_mai_n300_));
  NA2        m0272(.A(mai_mai_n224_), .B(mai_mai_n99_), .Y(mai_mai_n301_));
  OR2        m0273(.A(mai_mai_n301_), .B(mai_mai_n184_), .Y(mai_mai_n302_));
  NOi31      m0274(.An(l), .B(n), .C(m), .Y(mai_mai_n303_));
  NAi21      m0275(.An(mai_mai_n300_), .B(mai_mai_n302_), .Y(mai_mai_n304_));
  NAi32      m0276(.An(m), .Bn(j), .C(k), .Y(mai_mai_n305_));
  NAi41      m0277(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n189_), .B(mai_mai_n306_), .Y(mai_mai_n307_));
  NOi31      m0279(.An(j), .B(m), .C(k), .Y(mai_mai_n308_));
  NO2        m0280(.A(mai_mai_n120_), .B(mai_mai_n308_), .Y(mai_mai_n309_));
  AN3        m0281(.A(h), .B(m), .C(f), .Y(mai_mai_n310_));
  NAi31      m0282(.An(mai_mai_n309_), .B(mai_mai_n310_), .C(mai_mai_n307_), .Y(mai_mai_n311_));
  NOi32      m0283(.An(m), .Bn(j), .C(l), .Y(mai_mai_n312_));
  NO2        m0284(.A(mai_mai_n312_), .B(mai_mai_n93_), .Y(mai_mai_n313_));
  NO2        m0285(.A(mai_mai_n195_), .B(m), .Y(mai_mai_n314_));
  INV        m0286(.A(mai_mai_n210_), .Y(mai_mai_n315_));
  NA3        m0287(.A(mai_mai_n315_), .B(mai_mai_n310_), .C(mai_mai_n190_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n316_), .B(mai_mai_n311_), .Y(mai_mai_n317_));
  NA3        m0289(.A(h), .B(m), .C(f), .Y(mai_mai_n318_));
  NA2        m0290(.A(mai_mai_n147_), .B(e), .Y(mai_mai_n319_));
  INV        m0291(.A(mai_mai_n319_), .Y(mai_mai_n320_));
  NA2        m0292(.A(mai_mai_n320_), .B(mai_mai_n282_), .Y(mai_mai_n321_));
  NOi32      m0293(.An(j), .Bn(m), .C(i), .Y(mai_mai_n322_));
  NA3        m0294(.A(mai_mai_n322_), .B(mai_mai_n260_), .C(mai_mai_n107_), .Y(mai_mai_n323_));
  NOi32      m0295(.An(e), .Bn(b), .C(a), .Y(mai_mai_n324_));
  NO3        m0296(.A(mai_mai_n291_), .B(mai_mai_n70_), .C(mai_mai_n192_), .Y(mai_mai_n325_));
  NA2        m0297(.A(mai_mai_n187_), .B(mai_mai_n35_), .Y(mai_mai_n326_));
  AOI220     m0298(.A0(mai_mai_n326_), .A1(mai_mai_n324_), .B0(mai_mai_n325_), .B1(k), .Y(mai_mai_n327_));
  NO2        m0299(.A(mai_mai_n296_), .B(n), .Y(mai_mai_n328_));
  NA2        m0300(.A(mai_mai_n186_), .B(k), .Y(mai_mai_n329_));
  NA3        m0301(.A(m), .B(mai_mai_n106_), .C(mai_mai_n191_), .Y(mai_mai_n330_));
  NA4        m0302(.A(mai_mai_n183_), .B(mai_mai_n85_), .C(m), .D(mai_mai_n191_), .Y(mai_mai_n331_));
  OAI210     m0303(.A0(mai_mai_n330_), .A1(mai_mai_n329_), .B0(mai_mai_n331_), .Y(mai_mai_n332_));
  NAi41      m0304(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n333_));
  NA2        m0305(.A(mai_mai_n51_), .B(mai_mai_n107_), .Y(mai_mai_n334_));
  NA2        m0306(.A(mai_mai_n332_), .B(mai_mai_n328_), .Y(mai_mai_n335_));
  NA3        m0307(.A(mai_mai_n335_), .B(mai_mai_n327_), .C(mai_mai_n321_), .Y(mai_mai_n336_));
  NO4        m0308(.A(mai_mai_n336_), .B(mai_mai_n317_), .C(mai_mai_n304_), .D(mai_mai_n299_), .Y(mai_mai_n337_));
  NA4        m0309(.A(mai_mai_n337_), .B(mai_mai_n288_), .C(mai_mai_n242_), .D(mai_mai_n179_), .Y(mai10));
  NA3        m0310(.A(m), .B(k), .C(i), .Y(mai_mai_n339_));
  NO3        m0311(.A(mai_mai_n339_), .B(j), .C(mai_mai_n192_), .Y(mai_mai_n340_));
  NOi21      m0312(.An(e), .B(f), .Y(mai_mai_n341_));
  NO4        m0313(.A(mai_mai_n141_), .B(mai_mai_n341_), .C(n), .D(mai_mai_n104_), .Y(mai_mai_n342_));
  NA2        m0314(.A(h), .B(mai_mai_n197_), .Y(mai_mai_n343_));
  NA2        m0315(.A(mai_mai_n342_), .B(mai_mai_n340_), .Y(mai_mai_n344_));
  NO3        m0316(.A(n), .B(m), .C(k), .Y(mai_mai_n345_));
  NA2        m0317(.A(mai_mai_n345_), .B(h), .Y(mai_mai_n346_));
  NO3        m0318(.A(mai_mai_n346_), .B(mai_mai_n141_), .C(mai_mai_n191_), .Y(mai_mai_n347_));
  OR2        m0319(.A(m), .B(k), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n158_), .B(mai_mai_n348_), .Y(mai_mai_n349_));
  NA4        m0321(.A(n), .B(f), .C(c), .D(mai_mai_n110_), .Y(mai_mai_n350_));
  NOi32      m0322(.An(d), .Bn(a), .C(c), .Y(mai_mai_n351_));
  NA2        m0323(.A(mai_mai_n351_), .B(mai_mai_n163_), .Y(mai_mai_n352_));
  NAi21      m0324(.An(i), .B(m), .Y(mai_mai_n353_));
  NAi31      m0325(.An(k), .B(m), .C(j), .Y(mai_mai_n354_));
  NO3        m0326(.A(mai_mai_n354_), .B(mai_mai_n353_), .C(n), .Y(mai_mai_n355_));
  INV        m0327(.A(mai_mai_n347_), .Y(mai_mai_n356_));
  NOi32      m0328(.An(f), .Bn(d), .C(c), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n356_), .B(mai_mai_n344_), .Y(mai_mai_n358_));
  NO2        m0330(.A(mai_mai_n59_), .B(mai_mai_n110_), .Y(mai_mai_n359_));
  NA2        m0331(.A(mai_mai_n224_), .B(mai_mai_n359_), .Y(mai_mai_n360_));
  INV        m0332(.A(e), .Y(mai_mai_n361_));
  NA2        m0333(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n362_));
  OAI220     m0334(.A0(mai_mai_n362_), .A1(mai_mai_n180_), .B0(mai_mai_n184_), .B1(mai_mai_n361_), .Y(mai_mai_n363_));
  AN2        m0335(.A(m), .B(e), .Y(mai_mai_n364_));
  NA3        m0336(.A(mai_mai_n364_), .B(mai_mai_n183_), .C(i), .Y(mai_mai_n365_));
  INV        m0337(.A(mai_mai_n365_), .Y(mai_mai_n366_));
  NO2        m0338(.A(mai_mai_n96_), .B(mai_mai_n361_), .Y(mai_mai_n367_));
  NO3        m0339(.A(mai_mai_n367_), .B(mai_mai_n366_), .C(mai_mai_n363_), .Y(mai_mai_n368_));
  NOi32      m0340(.An(h), .Bn(e), .C(m), .Y(mai_mai_n369_));
  NA3        m0341(.A(mai_mai_n369_), .B(mai_mai_n262_), .C(m), .Y(mai_mai_n370_));
  NOi21      m0342(.An(m), .B(h), .Y(mai_mai_n371_));
  AN3        m0343(.A(m), .B(l), .C(i), .Y(mai_mai_n372_));
  NA3        m0344(.A(mai_mai_n372_), .B(mai_mai_n371_), .C(e), .Y(mai_mai_n373_));
  AN3        m0345(.A(h), .B(m), .C(e), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n374_), .B(mai_mai_n93_), .Y(mai_mai_n375_));
  AN3        m0347(.A(mai_mai_n375_), .B(mai_mai_n373_), .C(mai_mai_n370_), .Y(mai_mai_n376_));
  AOI210     m0348(.A0(mai_mai_n376_), .A1(mai_mai_n368_), .B0(mai_mai_n360_), .Y(mai_mai_n377_));
  NA3        m0349(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n378_));
  NO2        m0350(.A(mai_mai_n378_), .B(mai_mai_n360_), .Y(mai_mai_n379_));
  NA3        m0351(.A(mai_mai_n351_), .B(mai_mai_n163_), .C(mai_mai_n82_), .Y(mai_mai_n380_));
  NAi31      m0352(.An(b), .B(c), .C(a), .Y(mai_mai_n381_));
  NO2        m0353(.A(mai_mai_n381_), .B(n), .Y(mai_mai_n382_));
  OAI210     m0354(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n383_));
  NO2        m0355(.A(mai_mai_n383_), .B(mai_mai_n138_), .Y(mai_mai_n384_));
  NA2        m0356(.A(mai_mai_n384_), .B(mai_mai_n382_), .Y(mai_mai_n385_));
  INV        m0357(.A(mai_mai_n385_), .Y(mai_mai_n386_));
  NO4        m0358(.A(mai_mai_n386_), .B(mai_mai_n379_), .C(mai_mai_n377_), .D(mai_mai_n358_), .Y(mai_mai_n387_));
  NA2        m0359(.A(i), .B(m), .Y(mai_mai_n388_));
  NO3        m0360(.A(mai_mai_n251_), .B(mai_mai_n388_), .C(c), .Y(mai_mai_n389_));
  NA2        m0361(.A(d), .B(a), .Y(mai_mai_n390_));
  NA3        m0362(.A(i), .B(m), .C(f), .Y(mai_mai_n391_));
  OR2        m0363(.A(mai_mai_n391_), .B(mai_mai_n69_), .Y(mai_mai_n392_));
  NA2        m0364(.A(mai_mai_n389_), .B(mai_mai_n261_), .Y(mai_mai_n393_));
  OR2        m0365(.A(n), .B(m), .Y(mai_mai_n394_));
  INV        m0366(.A(mai_mai_n334_), .Y(mai_mai_n395_));
  NA2        m0367(.A(mai_mai_n395_), .B(mai_mai_n324_), .Y(mai_mai_n396_));
  NAi21      m0368(.An(k), .B(j), .Y(mai_mai_n397_));
  NAi21      m0369(.An(e), .B(d), .Y(mai_mai_n398_));
  INV        m0370(.A(mai_mai_n398_), .Y(mai_mai_n399_));
  NO2        m0371(.A(mai_mai_n227_), .B(mai_mai_n191_), .Y(mai_mai_n400_));
  NA3        m0372(.A(mai_mai_n400_), .B(mai_mai_n399_), .C(mai_mai_n203_), .Y(mai_mai_n401_));
  NA2        m0373(.A(mai_mai_n401_), .B(mai_mai_n396_), .Y(mai_mai_n402_));
  NOi31      m0374(.An(n), .B(m), .C(k), .Y(mai_mai_n403_));
  NAi31      m0375(.An(m), .B(f), .C(c), .Y(mai_mai_n404_));
  INV        m0376(.A(mai_mai_n281_), .Y(mai_mai_n405_));
  NOi41      m0377(.An(mai_mai_n393_), .B(mai_mai_n405_), .C(mai_mai_n402_), .D(mai_mai_n240_), .Y(mai_mai_n406_));
  NOi32      m0378(.An(c), .Bn(a), .C(b), .Y(mai_mai_n407_));
  NA2        m0379(.A(mai_mai_n407_), .B(mai_mai_n107_), .Y(mai_mai_n408_));
  INV        m0380(.A(mai_mai_n249_), .Y(mai_mai_n409_));
  AN2        m0381(.A(e), .B(d), .Y(mai_mai_n410_));
  NA2        m0382(.A(mai_mai_n410_), .B(mai_mai_n409_), .Y(mai_mai_n411_));
  NO2        m0383(.A(mai_mai_n125_), .B(mai_mai_n41_), .Y(mai_mai_n412_));
  NO2        m0384(.A(mai_mai_n65_), .B(e), .Y(mai_mai_n413_));
  NOi31      m0385(.An(j), .B(k), .C(i), .Y(mai_mai_n414_));
  NOi21      m0386(.An(mai_mai_n150_), .B(mai_mai_n414_), .Y(mai_mai_n415_));
  NA4        m0387(.A(mai_mai_n292_), .B(mai_mai_n415_), .C(mai_mai_n234_), .D(mai_mai_n113_), .Y(mai_mai_n416_));
  NA2        m0388(.A(mai_mai_n416_), .B(mai_mai_n413_), .Y(mai_mai_n417_));
  AOI210     m0389(.A0(mai_mai_n417_), .A1(mai_mai_n411_), .B0(mai_mai_n408_), .Y(mai_mai_n418_));
  NO2        m0390(.A(mai_mai_n188_), .B(mai_mai_n185_), .Y(mai_mai_n419_));
  NOi21      m0391(.An(a), .B(b), .Y(mai_mai_n420_));
  NA3        m0392(.A(e), .B(d), .C(c), .Y(mai_mai_n421_));
  NAi21      m0393(.An(mai_mai_n421_), .B(mai_mai_n420_), .Y(mai_mai_n422_));
  NO2        m0394(.A(mai_mai_n380_), .B(mai_mai_n184_), .Y(mai_mai_n423_));
  NOi21      m0395(.An(mai_mai_n422_), .B(mai_mai_n423_), .Y(mai_mai_n424_));
  AOI210     m0396(.A0(mai_mai_n243_), .A1(mai_mai_n419_), .B0(mai_mai_n424_), .Y(mai_mai_n425_));
  NO4        m0397(.A(mai_mai_n170_), .B(mai_mai_n98_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n426_));
  OR2        m0398(.A(k), .B(j), .Y(mai_mai_n427_));
  INV        m0399(.A(mai_mai_n122_), .Y(mai_mai_n428_));
  NA2        m0400(.A(mai_mai_n351_), .B(mai_mai_n107_), .Y(mai_mai_n429_));
  NO4        m0401(.A(mai_mai_n429_), .B(mai_mai_n90_), .C(mai_mai_n106_), .D(e), .Y(mai_mai_n430_));
  NO3        m0402(.A(mai_mai_n380_), .B(mai_mai_n89_), .C(mai_mai_n125_), .Y(mai_mai_n431_));
  NO4        m0403(.A(mai_mai_n431_), .B(mai_mai_n430_), .C(mai_mai_n428_), .D(mai_mai_n293_), .Y(mai_mai_n432_));
  INV        m0404(.A(mai_mai_n432_), .Y(mai_mai_n433_));
  NO4        m0405(.A(mai_mai_n433_), .B(mai_mai_n426_), .C(mai_mai_n425_), .D(mai_mai_n418_), .Y(mai_mai_n434_));
  NOi21      m0406(.An(d), .B(e), .Y(mai_mai_n435_));
  NO3        m0407(.A(mai_mai_n352_), .B(mai_mai_n313_), .C(mai_mai_n181_), .Y(mai_mai_n436_));
  NO2        m0408(.A(mai_mai_n352_), .B(mai_mai_n334_), .Y(mai_mai_n437_));
  NO4        m0409(.A(mai_mai_n437_), .B(mai_mai_n436_), .C(mai_mai_n166_), .D(mai_mai_n278_), .Y(mai_mai_n438_));
  NA2        m0410(.A(mai_mai_n438_), .B(mai_mai_n219_), .Y(mai_mai_n439_));
  OAI210     m0411(.A0(mai_mai_n121_), .A1(mai_mai_n120_), .B0(n), .Y(mai_mai_n440_));
  NO2        m0412(.A(mai_mai_n440_), .B(mai_mai_n125_), .Y(mai_mai_n441_));
  OA210      m0413(.A0(mai_mai_n221_), .A1(mai_mai_n441_), .B0(mai_mai_n174_), .Y(mai_mai_n442_));
  XO2        m0414(.A(i), .B(h), .Y(mai_mai_n443_));
  NA3        m0415(.A(mai_mai_n443_), .B(mai_mai_n145_), .C(n), .Y(mai_mai_n444_));
  NAi31      m0416(.An(mai_mai_n270_), .B(mai_mai_n444_), .C(mai_mai_n343_), .Y(mai_mai_n445_));
  NOi32      m0417(.An(mai_mai_n445_), .Bn(mai_mai_n413_), .C(mai_mai_n1281_), .Y(mai_mai_n446_));
  NAi31      m0418(.An(c), .B(f), .C(d), .Y(mai_mai_n447_));
  AOI210     m0419(.A0(mai_mai_n254_), .A1(mai_mai_n176_), .B0(mai_mai_n447_), .Y(mai_mai_n448_));
  NOi21      m0420(.An(mai_mai_n80_), .B(mai_mai_n448_), .Y(mai_mai_n449_));
  NA3        m0421(.A(mai_mai_n342_), .B(mai_mai_n93_), .C(mai_mai_n92_), .Y(mai_mai_n450_));
  NA2        m0422(.A(mai_mai_n204_), .B(mai_mai_n102_), .Y(mai_mai_n451_));
  NO2        m0423(.A(mai_mai_n451_), .B(mai_mai_n447_), .Y(mai_mai_n452_));
  AOI210     m0424(.A0(mai_mai_n323_), .A1(mai_mai_n35_), .B0(mai_mai_n422_), .Y(mai_mai_n453_));
  NOi31      m0425(.An(mai_mai_n450_), .B(mai_mai_n453_), .C(mai_mai_n452_), .Y(mai_mai_n454_));
  AO220      m0426(.A0(mai_mai_n258_), .A1(mai_mai_n237_), .B0(mai_mai_n151_), .B1(mai_mai_n66_), .Y(mai_mai_n455_));
  NA3        m0427(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n456_));
  NO2        m0428(.A(mai_mai_n456_), .B(mai_mai_n390_), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n457_), .B(mai_mai_n266_), .Y(mai_mai_n458_));
  NAi41      m0430(.An(mai_mai_n455_), .B(mai_mai_n458_), .C(mai_mai_n454_), .D(mai_mai_n449_), .Y(mai_mai_n459_));
  NO4        m0431(.A(mai_mai_n459_), .B(mai_mai_n446_), .C(mai_mai_n442_), .D(mai_mai_n439_), .Y(mai_mai_n460_));
  NA4        m0432(.A(mai_mai_n460_), .B(mai_mai_n434_), .C(mai_mai_n406_), .D(mai_mai_n387_), .Y(mai11));
  NO2        m0433(.A(mai_mai_n71_), .B(f), .Y(mai_mai_n462_));
  NA2        m0434(.A(j), .B(m), .Y(mai_mai_n463_));
  NAi31      m0435(.An(i), .B(m), .C(l), .Y(mai_mai_n464_));
  NA3        m0436(.A(m), .B(k), .C(j), .Y(mai_mai_n465_));
  OAI220     m0437(.A0(mai_mai_n465_), .A1(mai_mai_n125_), .B0(mai_mai_n464_), .B1(mai_mai_n463_), .Y(mai_mai_n466_));
  NA2        m0438(.A(mai_mai_n466_), .B(mai_mai_n462_), .Y(mai_mai_n467_));
  NOi32      m0439(.An(e), .Bn(b), .C(f), .Y(mai_mai_n468_));
  NA2        m0440(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n469_));
  NO2        m0441(.A(mai_mai_n469_), .B(mai_mai_n272_), .Y(mai_mai_n470_));
  NAi31      m0442(.An(d), .B(e), .C(a), .Y(mai_mai_n471_));
  NO2        m0443(.A(mai_mai_n471_), .B(n), .Y(mai_mai_n472_));
  AOI220     m0444(.A0(mai_mai_n472_), .A1(mai_mai_n97_), .B0(mai_mai_n470_), .B1(mai_mai_n468_), .Y(mai_mai_n473_));
  NAi41      m0445(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n474_));
  AN2        m0446(.A(mai_mai_n474_), .B(mai_mai_n333_), .Y(mai_mai_n475_));
  AOI210     m0447(.A0(mai_mai_n475_), .A1(mai_mai_n352_), .B0(mai_mai_n245_), .Y(mai_mai_n476_));
  NA2        m0448(.A(j), .B(i), .Y(mai_mai_n477_));
  NAi31      m0449(.An(n), .B(m), .C(k), .Y(mai_mai_n478_));
  NO3        m0450(.A(mai_mai_n478_), .B(mai_mai_n477_), .C(mai_mai_n106_), .Y(mai_mai_n479_));
  NO4        m0451(.A(n), .B(d), .C(mai_mai_n110_), .D(a), .Y(mai_mai_n480_));
  OR2        m0452(.A(n), .B(c), .Y(mai_mai_n481_));
  NO2        m0453(.A(mai_mai_n481_), .B(mai_mai_n140_), .Y(mai_mai_n482_));
  NO2        m0454(.A(mai_mai_n482_), .B(mai_mai_n480_), .Y(mai_mai_n483_));
  NOi32      m0455(.An(m), .Bn(f), .C(i), .Y(mai_mai_n484_));
  AOI220     m0456(.A0(mai_mai_n484_), .A1(mai_mai_n95_), .B0(mai_mai_n466_), .B1(f), .Y(mai_mai_n485_));
  NO2        m0457(.A(mai_mai_n249_), .B(mai_mai_n49_), .Y(mai_mai_n486_));
  NO2        m0458(.A(mai_mai_n485_), .B(mai_mai_n483_), .Y(mai_mai_n487_));
  AOI210     m0459(.A0(mai_mai_n479_), .A1(mai_mai_n476_), .B0(mai_mai_n487_), .Y(mai_mai_n488_));
  NA2        m0460(.A(mai_mai_n134_), .B(mai_mai_n34_), .Y(mai_mai_n489_));
  OAI220     m0461(.A0(mai_mai_n489_), .A1(m), .B0(mai_mai_n469_), .B1(mai_mai_n210_), .Y(mai_mai_n490_));
  NOi41      m0462(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n491_));
  AN2        m0463(.A(mai_mai_n306_), .B(mai_mai_n291_), .Y(mai_mai_n492_));
  AN2        m0464(.A(mai_mai_n491_), .B(mai_mai_n490_), .Y(mai_mai_n493_));
  OAI220     m0465(.A0(mai_mai_n354_), .A1(mai_mai_n353_), .B0(mai_mai_n464_), .B1(mai_mai_n463_), .Y(mai_mai_n494_));
  NAi31      m0466(.An(d), .B(c), .C(a), .Y(mai_mai_n495_));
  NO2        m0467(.A(mai_mai_n495_), .B(n), .Y(mai_mai_n496_));
  NA3        m0468(.A(mai_mai_n496_), .B(mai_mai_n494_), .C(e), .Y(mai_mai_n497_));
  NO3        m0469(.A(mai_mai_n61_), .B(mai_mai_n49_), .C(mai_mai_n192_), .Y(mai_mai_n498_));
  NO2        m0470(.A(mai_mai_n207_), .B(mai_mai_n104_), .Y(mai_mai_n499_));
  OAI210     m0471(.A0(mai_mai_n498_), .A1(mai_mai_n355_), .B0(mai_mai_n499_), .Y(mai_mai_n500_));
  NA2        m0472(.A(mai_mai_n500_), .B(mai_mai_n497_), .Y(mai_mai_n501_));
  NO2        m0473(.A(mai_mai_n251_), .B(n), .Y(mai_mai_n502_));
  NO2        m0474(.A(mai_mai_n382_), .B(mai_mai_n502_), .Y(mai_mai_n503_));
  NA2        m0475(.A(mai_mai_n494_), .B(f), .Y(mai_mai_n504_));
  NAi32      m0476(.An(d), .Bn(a), .C(b), .Y(mai_mai_n505_));
  NA2        m0477(.A(h), .B(f), .Y(mai_mai_n506_));
  NO2        m0478(.A(mai_mai_n506_), .B(mai_mai_n90_), .Y(mai_mai_n507_));
  NO3        m0479(.A(mai_mai_n160_), .B(mai_mai_n158_), .C(m), .Y(mai_mai_n508_));
  NA2        m0480(.A(mai_mai_n508_), .B(mai_mai_n58_), .Y(mai_mai_n509_));
  OAI210     m0481(.A0(mai_mai_n504_), .A1(mai_mai_n503_), .B0(mai_mai_n509_), .Y(mai_mai_n510_));
  AN3        m0482(.A(j), .B(h), .C(m), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n137_), .B(c), .Y(mai_mai_n512_));
  NA3        m0484(.A(mai_mai_n512_), .B(mai_mai_n511_), .C(mai_mai_n403_), .Y(mai_mai_n513_));
  NA3        m0485(.A(f), .B(d), .C(b), .Y(mai_mai_n514_));
  INV        m0486(.A(mai_mai_n513_), .Y(mai_mai_n515_));
  NO4        m0487(.A(mai_mai_n515_), .B(mai_mai_n510_), .C(mai_mai_n501_), .D(mai_mai_n493_), .Y(mai_mai_n516_));
  AN4        m0488(.A(mai_mai_n516_), .B(mai_mai_n488_), .C(mai_mai_n473_), .D(mai_mai_n467_), .Y(mai_mai_n517_));
  INV        m0489(.A(k), .Y(mai_mai_n518_));
  NA3        m0490(.A(l), .B(mai_mai_n518_), .C(i), .Y(mai_mai_n519_));
  INV        m0491(.A(mai_mai_n519_), .Y(mai_mai_n520_));
  NAi32      m0492(.An(h), .Bn(f), .C(m), .Y(mai_mai_n521_));
  NAi41      m0493(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n522_));
  OAI210     m0494(.A0(mai_mai_n471_), .A1(n), .B0(mai_mai_n522_), .Y(mai_mai_n523_));
  NA2        m0495(.A(mai_mai_n523_), .B(m), .Y(mai_mai_n524_));
  NAi31      m0496(.An(h), .B(m), .C(f), .Y(mai_mai_n525_));
  OR3        m0497(.A(mai_mai_n525_), .B(mai_mai_n251_), .C(mai_mai_n49_), .Y(mai_mai_n526_));
  NA4        m0498(.A(mai_mai_n371_), .B(mai_mai_n115_), .C(mai_mai_n107_), .D(e), .Y(mai_mai_n527_));
  AN2        m0499(.A(mai_mai_n527_), .B(mai_mai_n526_), .Y(mai_mai_n528_));
  OA210      m0500(.A0(mai_mai_n524_), .A1(mai_mai_n521_), .B0(mai_mai_n528_), .Y(mai_mai_n529_));
  INV        m0501(.A(mai_mai_n529_), .Y(mai_mai_n530_));
  NAi31      m0502(.An(f), .B(h), .C(m), .Y(mai_mai_n531_));
  NO4        m0503(.A(mai_mai_n283_), .B(mai_mai_n531_), .C(mai_mai_n71_), .D(mai_mai_n72_), .Y(mai_mai_n532_));
  NOi32      m0504(.An(b), .Bn(a), .C(c), .Y(mai_mai_n533_));
  NOi41      m0505(.An(mai_mai_n533_), .B(mai_mai_n318_), .C(mai_mai_n68_), .D(mai_mai_n111_), .Y(mai_mai_n534_));
  OR2        m0506(.A(mai_mai_n534_), .B(mai_mai_n532_), .Y(mai_mai_n535_));
  NOi32      m0507(.An(d), .Bn(a), .C(e), .Y(mai_mai_n536_));
  NA2        m0508(.A(mai_mai_n536_), .B(mai_mai_n107_), .Y(mai_mai_n537_));
  NO2        m0509(.A(n), .B(c), .Y(mai_mai_n538_));
  NA3        m0510(.A(mai_mai_n538_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n539_));
  NOi32      m0511(.An(e), .Bn(a), .C(d), .Y(mai_mai_n540_));
  AOI210     m0512(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n540_), .Y(mai_mai_n541_));
  NO2        m0513(.A(mai_mai_n541_), .B(mai_mai_n489_), .Y(mai_mai_n542_));
  AOI210     m0514(.A0(mai_mai_n542_), .A1(mai_mai_n107_), .B0(mai_mai_n535_), .Y(mai_mai_n543_));
  INV        m0515(.A(mai_mai_n543_), .Y(mai_mai_n544_));
  AOI210     m0516(.A0(mai_mai_n530_), .A1(mai_mai_n520_), .B0(mai_mai_n544_), .Y(mai_mai_n545_));
  NO3        m0517(.A(mai_mai_n290_), .B(mai_mai_n60_), .C(n), .Y(mai_mai_n546_));
  INV        m0518(.A(mai_mai_n207_), .Y(mai_mai_n547_));
  NA2        m0519(.A(mai_mai_n73_), .B(mai_mai_n107_), .Y(mai_mai_n548_));
  NO2        m0520(.A(mai_mai_n548_), .B(mai_mai_n45_), .Y(mai_mai_n549_));
  AOI220     m0521(.A0(mai_mai_n549_), .A1(mai_mai_n476_), .B0(mai_mai_n547_), .B1(mai_mai_n546_), .Y(mai_mai_n550_));
  NO2        m0522(.A(mai_mai_n550_), .B(mai_mai_n85_), .Y(mai_mai_n551_));
  NOi32      m0523(.An(e), .Bn(c), .C(f), .Y(mai_mai_n552_));
  NOi21      m0524(.An(f), .B(m), .Y(mai_mai_n553_));
  AOI210     m0525(.A0(mai_mai_n475_), .A1(mai_mai_n352_), .B0(mai_mai_n271_), .Y(mai_mai_n554_));
  NA2        m0526(.A(mai_mai_n554_), .B(mai_mai_n238_), .Y(mai_mai_n555_));
  NOi31      m0527(.An(m), .B(n), .C(k), .Y(mai_mai_n556_));
  NA2        m0528(.A(j), .B(mai_mai_n556_), .Y(mai_mai_n557_));
  AOI210     m0529(.A0(mai_mai_n352_), .A1(mai_mai_n333_), .B0(mai_mai_n271_), .Y(mai_mai_n558_));
  NAi21      m0530(.An(mai_mai_n557_), .B(mai_mai_n558_), .Y(mai_mai_n559_));
  NO2        m0531(.A(mai_mai_n251_), .B(mai_mai_n49_), .Y(mai_mai_n560_));
  NO2        m0532(.A(mai_mai_n471_), .B(mai_mai_n49_), .Y(mai_mai_n561_));
  NA2        m0533(.A(mai_mai_n560_), .B(mai_mai_n507_), .Y(mai_mai_n562_));
  NA3        m0534(.A(mai_mai_n562_), .B(mai_mai_n559_), .C(mai_mai_n555_), .Y(mai_mai_n563_));
  NA2        m0535(.A(mai_mai_n102_), .B(mai_mai_n36_), .Y(mai_mai_n564_));
  NO2        m0536(.A(k), .B(mai_mai_n192_), .Y(mai_mai_n565_));
  NO2        m0537(.A(mai_mai_n468_), .B(mai_mai_n324_), .Y(mai_mai_n566_));
  NO2        m0538(.A(mai_mai_n566_), .B(n), .Y(mai_mai_n567_));
  NAi31      m0539(.An(mai_mai_n564_), .B(mai_mai_n567_), .C(mai_mai_n565_), .Y(mai_mai_n568_));
  NO2        m0540(.A(mai_mai_n469_), .B(mai_mai_n160_), .Y(mai_mai_n569_));
  AN3        m0541(.A(f), .B(d), .C(b), .Y(mai_mai_n570_));
  NA3        m0542(.A(mai_mai_n443_), .B(mai_mai_n145_), .C(mai_mai_n192_), .Y(mai_mai_n571_));
  AOI210     m0543(.A0(mai_mai_n1282_), .A1(mai_mai_n209_), .B0(mai_mai_n571_), .Y(mai_mai_n572_));
  NAi31      m0544(.An(m), .B(n), .C(k), .Y(mai_mai_n573_));
  INV        m0545(.A(mai_mai_n225_), .Y(mai_mai_n574_));
  OAI210     m0546(.A0(mai_mai_n574_), .A1(mai_mai_n572_), .B0(j), .Y(mai_mai_n575_));
  NA2        m0547(.A(mai_mai_n575_), .B(mai_mai_n568_), .Y(mai_mai_n576_));
  NO3        m0548(.A(mai_mai_n576_), .B(mai_mai_n563_), .C(mai_mai_n551_), .Y(mai_mai_n577_));
  NAi31      m0549(.An(m), .B(h), .C(f), .Y(mai_mai_n578_));
  OR3        m0550(.A(mai_mai_n578_), .B(mai_mai_n251_), .C(n), .Y(mai_mai_n579_));
  OA210      m0551(.A0(mai_mai_n471_), .A1(n), .B0(mai_mai_n522_), .Y(mai_mai_n580_));
  NA3        m0552(.A(mai_mai_n369_), .B(mai_mai_n115_), .C(mai_mai_n82_), .Y(mai_mai_n581_));
  OAI210     m0553(.A0(mai_mai_n580_), .A1(mai_mai_n88_), .B0(mai_mai_n581_), .Y(mai_mai_n582_));
  NOi21      m0554(.An(mai_mai_n579_), .B(mai_mai_n582_), .Y(mai_mai_n583_));
  NO2        m0555(.A(mai_mai_n583_), .B(mai_mai_n465_), .Y(mai_mai_n584_));
  NO3        m0556(.A(m), .B(mai_mai_n191_), .C(mai_mai_n56_), .Y(mai_mai_n585_));
  NAi21      m0557(.An(h), .B(j), .Y(mai_mai_n586_));
  NO2        m0558(.A(mai_mai_n451_), .B(mai_mai_n85_), .Y(mai_mai_n587_));
  OAI210     m0559(.A0(mai_mai_n587_), .A1(mai_mai_n349_), .B0(mai_mai_n585_), .Y(mai_mai_n588_));
  BUFFER     m0560(.A(mai_mai_n71_), .Y(mai_mai_n589_));
  NA3        m0561(.A(mai_mai_n462_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n590_));
  NA2        m0562(.A(mai_mai_n95_), .B(mai_mai_n46_), .Y(mai_mai_n591_));
  NO2        m0563(.A(mai_mai_n591_), .B(mai_mai_n301_), .Y(mai_mai_n592_));
  AOI210     m0564(.A0(mai_mai_n505_), .A1(mai_mai_n381_), .B0(mai_mai_n49_), .Y(mai_mai_n593_));
  OAI220     m0565(.A0(mai_mai_n525_), .A1(mai_mai_n519_), .B0(mai_mai_n294_), .B1(mai_mai_n463_), .Y(mai_mai_n594_));
  AOI210     m0566(.A0(mai_mai_n594_), .A1(mai_mai_n593_), .B0(mai_mai_n592_), .Y(mai_mai_n595_));
  NA3        m0567(.A(mai_mai_n595_), .B(mai_mai_n590_), .C(mai_mai_n588_), .Y(mai_mai_n596_));
  NO2        m0568(.A(mai_mai_n226_), .B(f), .Y(mai_mai_n597_));
  NA2        m0569(.A(mai_mai_n297_), .B(mai_mai_n134_), .Y(mai_mai_n598_));
  NA2        m0570(.A(mai_mai_n126_), .B(mai_mai_n49_), .Y(mai_mai_n599_));
  AOI220     m0571(.A0(mai_mai_n599_), .A1(mai_mai_n468_), .B0(mai_mai_n324_), .B1(mai_mai_n107_), .Y(mai_mai_n600_));
  OA220      m0572(.A0(mai_mai_n600_), .A1(mai_mai_n489_), .B0(mai_mai_n323_), .B1(mai_mai_n105_), .Y(mai_mai_n601_));
  NA2        m0573(.A(mai_mai_n598_), .B(mai_mai_n601_), .Y(mai_mai_n602_));
  NA2        m0574(.A(mai_mai_n407_), .B(mai_mai_n82_), .Y(mai_mai_n603_));
  NO4        m0575(.A(mai_mai_n465_), .B(mai_mai_n603_), .C(mai_mai_n125_), .D(mai_mai_n191_), .Y(mai_mai_n604_));
  INV        m0576(.A(mai_mai_n604_), .Y(mai_mai_n605_));
  NA3        m0577(.A(mai_mai_n605_), .B(mai_mai_n450_), .C(mai_mai_n356_), .Y(mai_mai_n606_));
  NO4        m0578(.A(mai_mai_n606_), .B(mai_mai_n602_), .C(mai_mai_n596_), .D(mai_mai_n584_), .Y(mai_mai_n607_));
  NA4        m0579(.A(mai_mai_n607_), .B(mai_mai_n577_), .C(mai_mai_n545_), .D(mai_mai_n517_), .Y(mai08));
  NO2        m0580(.A(k), .B(h), .Y(mai_mai_n609_));
  AO210      m0581(.A0(mai_mai_n226_), .A1(mai_mai_n397_), .B0(mai_mai_n609_), .Y(mai_mai_n610_));
  NO2        m0582(.A(mai_mai_n610_), .B(mai_mai_n269_), .Y(mai_mai_n611_));
  NA2        m0583(.A(mai_mai_n552_), .B(mai_mai_n82_), .Y(mai_mai_n612_));
  NA2        m0584(.A(mai_mai_n612_), .B(mai_mai_n404_), .Y(mai_mai_n613_));
  AOI210     m0585(.A0(mai_mai_n613_), .A1(mai_mai_n611_), .B0(mai_mai_n431_), .Y(mai_mai_n614_));
  NA2        m0586(.A(mai_mai_n82_), .B(mai_mai_n104_), .Y(mai_mai_n615_));
  NO2        m0587(.A(mai_mai_n615_), .B(mai_mai_n57_), .Y(mai_mai_n616_));
  NA2        m0588(.A(mai_mai_n514_), .B(mai_mai_n209_), .Y(mai_mai_n617_));
  NA2        m0589(.A(mai_mai_n617_), .B(mai_mai_n314_), .Y(mai_mai_n618_));
  NA2        m0590(.A(mai_mai_n514_), .B(mai_mai_n143_), .Y(mai_mai_n619_));
  NA4        m0591(.A(mai_mai_n194_), .B(mai_mai_n134_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n620_));
  AN2        m0592(.A(l), .B(k), .Y(mai_mai_n621_));
  NA4        m0593(.A(mai_mai_n621_), .B(mai_mai_n102_), .C(mai_mai_n72_), .D(mai_mai_n192_), .Y(mai_mai_n622_));
  OAI210     m0594(.A0(mai_mai_n620_), .A1(m), .B0(mai_mai_n622_), .Y(mai_mai_n623_));
  NA2        m0595(.A(mai_mai_n623_), .B(mai_mai_n619_), .Y(mai_mai_n624_));
  NA3        m0596(.A(mai_mai_n624_), .B(mai_mai_n618_), .C(mai_mai_n614_), .Y(mai_mai_n625_));
  NO4        m0597(.A(mai_mai_n158_), .B(mai_mai_n348_), .C(mai_mai_n106_), .D(m), .Y(mai_mai_n626_));
  AOI210     m0598(.A0(mai_mai_n626_), .A1(mai_mai_n617_), .B0(mai_mai_n457_), .Y(mai_mai_n627_));
  NO2        m0599(.A(mai_mai_n38_), .B(mai_mai_n191_), .Y(mai_mai_n628_));
  INV        m0600(.A(mai_mai_n627_), .Y(mai_mai_n629_));
  NA2        m0601(.A(mai_mai_n324_), .B(mai_mai_n43_), .Y(mai_mai_n630_));
  NA2        m0602(.A(mai_mai_n621_), .B(mai_mai_n197_), .Y(mai_mai_n631_));
  NO2        m0603(.A(mai_mai_n631_), .B(mai_mai_n296_), .Y(mai_mai_n632_));
  AOI210     m0604(.A0(mai_mai_n632_), .A1(mai_mai_n597_), .B0(mai_mai_n430_), .Y(mai_mai_n633_));
  NA3        m0605(.A(m), .B(l), .C(k), .Y(mai_mai_n634_));
  AOI210     m0606(.A0(mai_mai_n581_), .A1(mai_mai_n579_), .B0(mai_mai_n634_), .Y(mai_mai_n635_));
  NO2        m0607(.A(mai_mai_n474_), .B(mai_mai_n245_), .Y(mai_mai_n636_));
  NOi21      m0608(.An(mai_mai_n636_), .B(n), .Y(mai_mai_n637_));
  NA4        m0609(.A(mai_mai_n107_), .B(l), .C(k), .D(mai_mai_n85_), .Y(mai_mai_n638_));
  NA3        m0610(.A(mai_mai_n115_), .B(mai_mai_n364_), .C(i), .Y(mai_mai_n639_));
  NO2        m0611(.A(mai_mai_n639_), .B(mai_mai_n638_), .Y(mai_mai_n640_));
  NO3        m0612(.A(mai_mai_n640_), .B(mai_mai_n637_), .C(mai_mai_n635_), .Y(mai_mai_n641_));
  NA3        m0613(.A(mai_mai_n641_), .B(mai_mai_n633_), .C(mai_mai_n630_), .Y(mai_mai_n642_));
  NO3        m0614(.A(mai_mai_n642_), .B(mai_mai_n629_), .C(mai_mai_n625_), .Y(mai_mai_n643_));
  NOi31      m0615(.An(m), .B(h), .C(f), .Y(mai_mai_n644_));
  NA2        m0616(.A(mai_mai_n561_), .B(mai_mai_n644_), .Y(mai_mai_n645_));
  INV        m0617(.A(mai_mai_n225_), .Y(mai_mai_n646_));
  NA2        m0618(.A(mai_mai_n621_), .B(mai_mai_n72_), .Y(mai_mai_n647_));
  NOi21      m0619(.An(h), .B(j), .Y(mai_mai_n648_));
  NA2        m0620(.A(mai_mai_n648_), .B(f), .Y(mai_mai_n649_));
  NO2        m0621(.A(mai_mai_n649_), .B(e), .Y(mai_mai_n650_));
  INV        m0622(.A(mai_mai_n650_), .Y(mai_mai_n651_));
  OAI210     m0623(.A0(mai_mai_n651_), .A1(mai_mai_n647_), .B0(mai_mai_n528_), .Y(mai_mai_n652_));
  NO2        m0624(.A(mai_mai_n646_), .B(mai_mai_n652_), .Y(mai_mai_n653_));
  NO2        m0625(.A(j), .B(i), .Y(mai_mai_n654_));
  NA2        m0626(.A(mai_mai_n654_), .B(mai_mai_n33_), .Y(mai_mai_n655_));
  NA2        m0627(.A(mai_mai_n374_), .B(mai_mai_n115_), .Y(mai_mai_n656_));
  OR2        m0628(.A(mai_mai_n656_), .B(mai_mai_n655_), .Y(mai_mai_n657_));
  NO3        m0629(.A(mai_mai_n141_), .B(mai_mai_n49_), .C(mai_mai_n104_), .Y(mai_mai_n658_));
  NO3        m0630(.A(mai_mai_n481_), .B(mai_mai_n140_), .C(mai_mai_n72_), .Y(mai_mai_n659_));
  NO2        m0631(.A(mai_mai_n391_), .B(j), .Y(mai_mai_n660_));
  OAI210     m0632(.A0(mai_mai_n659_), .A1(mai_mai_n658_), .B0(mai_mai_n660_), .Y(mai_mai_n661_));
  NA2        m0633(.A(mai_mai_n645_), .B(mai_mai_n661_), .Y(mai_mai_n662_));
  NA2        m0634(.A(k), .B(j), .Y(mai_mai_n663_));
  NO3        m0635(.A(mai_mai_n269_), .B(mai_mai_n663_), .C(mai_mai_n40_), .Y(mai_mai_n664_));
  AOI210     m0636(.A0(mai_mai_n468_), .A1(n), .B0(mai_mai_n491_), .Y(mai_mai_n665_));
  NA2        m0637(.A(mai_mai_n665_), .B(mai_mai_n492_), .Y(mai_mai_n666_));
  AN3        m0638(.A(mai_mai_n666_), .B(mai_mai_n664_), .C(mai_mai_n94_), .Y(mai_mai_n667_));
  NO2        m0639(.A(mai_mai_n269_), .B(mai_mai_n130_), .Y(mai_mai_n668_));
  NO2        m0640(.A(mai_mai_n634_), .B(mai_mai_n88_), .Y(mai_mai_n669_));
  NA2        m0641(.A(mai_mai_n669_), .B(mai_mai_n523_), .Y(mai_mai_n670_));
  NO2        m0642(.A(mai_mai_n525_), .B(mai_mai_n111_), .Y(mai_mai_n671_));
  OAI210     m0643(.A0(mai_mai_n671_), .A1(mai_mai_n660_), .B0(mai_mai_n593_), .Y(mai_mai_n672_));
  NA2        m0644(.A(mai_mai_n672_), .B(mai_mai_n670_), .Y(mai_mai_n673_));
  OR3        m0645(.A(mai_mai_n673_), .B(mai_mai_n667_), .C(mai_mai_n662_), .Y(mai_mai_n674_));
  OAI220     m0646(.A0(mai_mai_n620_), .A1(mai_mai_n612_), .B0(mai_mai_n301_), .B1(mai_mai_n38_), .Y(mai_mai_n675_));
  INV        m0647(.A(mai_mai_n675_), .Y(mai_mai_n676_));
  NA3        m0648(.A(mai_mai_n484_), .B(mai_mai_n262_), .C(h), .Y(mai_mai_n677_));
  NOi21      m0649(.An(mai_mai_n593_), .B(mai_mai_n677_), .Y(mai_mai_n678_));
  NO2        m0650(.A(mai_mai_n89_), .B(mai_mai_n47_), .Y(mai_mai_n679_));
  NO2        m0651(.A(mai_mai_n677_), .B(mai_mai_n539_), .Y(mai_mai_n680_));
  AOI210     m0652(.A0(mai_mai_n679_), .A1(mai_mai_n567_), .B0(mai_mai_n680_), .Y(mai_mai_n681_));
  NAi31      m0653(.An(mai_mai_n678_), .B(mai_mai_n681_), .C(mai_mai_n676_), .Y(mai_mai_n682_));
  OR2        m0654(.A(mai_mai_n669_), .B(mai_mai_n91_), .Y(mai_mai_n683_));
  AOI220     m0655(.A0(mai_mai_n683_), .A1(mai_mai_n214_), .B0(mai_mai_n660_), .B1(mai_mai_n560_), .Y(mai_mai_n684_));
  OAI210     m0656(.A0(mai_mai_n634_), .A1(mai_mai_n578_), .B0(mai_mai_n456_), .Y(mai_mai_n685_));
  NA3        m0657(.A(mai_mai_n224_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n686_));
  AOI220     m0658(.A0(mai_mai_n538_), .A1(mai_mai_n29_), .B0(mai_mai_n407_), .B1(mai_mai_n82_), .Y(mai_mai_n687_));
  NA2        m0659(.A(mai_mai_n687_), .B(mai_mai_n686_), .Y(mai_mai_n688_));
  NO2        m0660(.A(mai_mai_n677_), .B(mai_mai_n429_), .Y(mai_mai_n689_));
  AOI210     m0661(.A0(mai_mai_n688_), .A1(mai_mai_n685_), .B0(mai_mai_n689_), .Y(mai_mai_n690_));
  NA2        m0662(.A(mai_mai_n690_), .B(mai_mai_n684_), .Y(mai_mai_n691_));
  NOi41      m0663(.An(mai_mai_n657_), .B(mai_mai_n691_), .C(mai_mai_n682_), .D(mai_mai_n674_), .Y(mai_mai_n692_));
  OR3        m0664(.A(mai_mai_n620_), .B(mai_mai_n209_), .C(m), .Y(mai_mai_n693_));
  NO3        m0665(.A(mai_mai_n309_), .B(mai_mai_n271_), .C(mai_mai_n106_), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n694_), .B(mai_mai_n666_), .Y(mai_mai_n695_));
  INV        m0667(.A(mai_mai_n46_), .Y(mai_mai_n696_));
  NO3        m0668(.A(mai_mai_n696_), .B(mai_mai_n655_), .C(mai_mai_n251_), .Y(mai_mai_n697_));
  NO2        m0669(.A(mai_mai_n463_), .B(h), .Y(mai_mai_n698_));
  AOI210     m0670(.A0(mai_mai_n698_), .A1(mai_mai_n616_), .B0(mai_mai_n697_), .Y(mai_mai_n699_));
  NA3        m0671(.A(mai_mai_n699_), .B(mai_mai_n695_), .C(mai_mai_n693_), .Y(mai_mai_n700_));
  OR2        m0672(.A(mai_mai_n578_), .B(mai_mai_n89_), .Y(mai_mai_n701_));
  NOi31      m0673(.An(b), .B(d), .C(a), .Y(mai_mai_n702_));
  NO2        m0674(.A(mai_mai_n702_), .B(mai_mai_n536_), .Y(mai_mai_n703_));
  NO2        m0675(.A(mai_mai_n703_), .B(n), .Y(mai_mai_n704_));
  NOi21      m0676(.An(mai_mai_n687_), .B(mai_mai_n704_), .Y(mai_mai_n705_));
  NO2        m0677(.A(mai_mai_n705_), .B(mai_mai_n701_), .Y(mai_mai_n706_));
  NO2        m0678(.A(mai_mai_n296_), .B(mai_mai_n111_), .Y(mai_mai_n707_));
  NOi21      m0679(.An(mai_mai_n707_), .B(mai_mai_n146_), .Y(mai_mai_n708_));
  INV        m0680(.A(mai_mai_n708_), .Y(mai_mai_n709_));
  OAI210     m0681(.A0(mai_mai_n620_), .A1(mai_mai_n350_), .B0(mai_mai_n709_), .Y(mai_mai_n710_));
  NA2        m0682(.A(mai_mai_n668_), .B(mai_mai_n585_), .Y(mai_mai_n711_));
  INV        m0683(.A(mai_mai_n213_), .Y(mai_mai_n712_));
  NA2        m0684(.A(mai_mai_n115_), .B(mai_mai_n82_), .Y(mai_mai_n713_));
  AOI210     m0685(.A0(mai_mai_n378_), .A1(mai_mai_n370_), .B0(mai_mai_n713_), .Y(mai_mai_n714_));
  NA2        m0686(.A(mai_mai_n632_), .B(mai_mai_n34_), .Y(mai_mai_n715_));
  NAi21      m0687(.An(mai_mai_n638_), .B(mai_mai_n389_), .Y(mai_mai_n716_));
  NO2        m0688(.A(mai_mai_n245_), .B(i), .Y(mai_mai_n717_));
  NAi41      m0689(.An(mai_mai_n714_), .B(mai_mai_n716_), .C(mai_mai_n715_), .D(mai_mai_n711_), .Y(mai_mai_n718_));
  NO4        m0690(.A(mai_mai_n718_), .B(mai_mai_n710_), .C(mai_mai_n706_), .D(mai_mai_n700_), .Y(mai_mai_n719_));
  NA4        m0691(.A(mai_mai_n719_), .B(mai_mai_n692_), .C(mai_mai_n653_), .D(mai_mai_n643_), .Y(mai09));
  INV        m0692(.A(mai_mai_n116_), .Y(mai_mai_n721_));
  NA2        m0693(.A(f), .B(e), .Y(mai_mai_n722_));
  NO2        m0694(.A(mai_mai_n202_), .B(mai_mai_n106_), .Y(mai_mai_n723_));
  NA2        m0695(.A(mai_mai_n723_), .B(m), .Y(mai_mai_n724_));
  NA4        m0696(.A(mai_mai_n283_), .B(mai_mai_n415_), .C(mai_mai_n234_), .D(mai_mai_n113_), .Y(mai_mai_n725_));
  AOI210     m0697(.A0(mai_mai_n725_), .A1(m), .B0(mai_mai_n412_), .Y(mai_mai_n726_));
  AOI210     m0698(.A0(mai_mai_n726_), .A1(mai_mai_n724_), .B0(mai_mai_n722_), .Y(mai_mai_n727_));
  NA2        m0699(.A(mai_mai_n727_), .B(mai_mai_n721_), .Y(mai_mai_n728_));
  NO2        m0700(.A(mai_mai_n184_), .B(mai_mai_n191_), .Y(mai_mai_n729_));
  NA3        m0701(.A(m), .B(l), .C(i), .Y(mai_mai_n730_));
  OAI220     m0702(.A0(mai_mai_n525_), .A1(mai_mai_n730_), .B0(mai_mai_n318_), .B1(mai_mai_n464_), .Y(mai_mai_n731_));
  NA4        m0703(.A(mai_mai_n86_), .B(mai_mai_n85_), .C(m), .D(f), .Y(mai_mai_n732_));
  NAi31      m0704(.An(mai_mai_n731_), .B(mai_mai_n732_), .C(mai_mai_n392_), .Y(mai_mai_n733_));
  OR2        m0705(.A(mai_mai_n733_), .B(mai_mai_n729_), .Y(mai_mai_n734_));
  NA3        m0706(.A(mai_mai_n701_), .B(mai_mai_n504_), .C(mai_mai_n456_), .Y(mai_mai_n735_));
  OA210      m0707(.A0(mai_mai_n735_), .A1(mai_mai_n734_), .B0(mai_mai_n704_), .Y(mai_mai_n736_));
  INV        m0708(.A(mai_mai_n306_), .Y(mai_mai_n737_));
  NO2        m0709(.A(mai_mai_n121_), .B(mai_mai_n120_), .Y(mai_mai_n738_));
  NA2        m0710(.A(mai_mai_n686_), .B(mai_mai_n301_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n310_), .B(mai_mai_n312_), .Y(mai_mai_n740_));
  OAI210     m0712(.A0(mai_mai_n184_), .A1(mai_mai_n191_), .B0(mai_mai_n740_), .Y(mai_mai_n741_));
  NA2        m0713(.A(mai_mai_n741_), .B(mai_mai_n739_), .Y(mai_mai_n742_));
  NA2        m0714(.A(mai_mai_n154_), .B(mai_mai_n108_), .Y(mai_mai_n743_));
  NA2        m0715(.A(mai_mai_n743_), .B(mai_mai_n610_), .Y(mai_mai_n744_));
  NA3        m0716(.A(mai_mai_n744_), .B(mai_mai_n172_), .C(mai_mai_n31_), .Y(mai_mai_n745_));
  NA3        m0717(.A(mai_mai_n745_), .B(mai_mai_n742_), .C(mai_mai_n80_), .Y(mai_mai_n746_));
  NO2        m0718(.A(mai_mai_n521_), .B(j), .Y(mai_mai_n747_));
  NOi21      m0719(.An(f), .B(d), .Y(mai_mai_n748_));
  NA2        m0720(.A(mai_mai_n748_), .B(m), .Y(mai_mai_n749_));
  NO2        m0721(.A(mai_mai_n749_), .B(mai_mai_n52_), .Y(mai_mai_n750_));
  NOi32      m0722(.An(m), .Bn(f), .C(d), .Y(mai_mai_n751_));
  NA4        m0723(.A(mai_mai_n751_), .B(mai_mai_n538_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n752_));
  NA2        m0724(.A(mai_mai_n750_), .B(mai_mai_n482_), .Y(mai_mai_n753_));
  NA3        m0725(.A(mai_mai_n420_), .B(d), .C(mai_mai_n82_), .Y(mai_mai_n754_));
  NO3        m0726(.A(mai_mai_n754_), .B(mai_mai_n72_), .C(mai_mai_n192_), .Y(mai_mai_n755_));
  NO2        m0727(.A(mai_mai_n256_), .B(mai_mai_n56_), .Y(mai_mai_n756_));
  NAi21      m0728(.An(mai_mai_n428_), .B(mai_mai_n753_), .Y(mai_mai_n757_));
  NO2        m0729(.A(mai_mai_n573_), .B(mai_mai_n296_), .Y(mai_mai_n758_));
  AN2        m0730(.A(mai_mai_n758_), .B(mai_mai_n597_), .Y(mai_mai_n759_));
  NO2        m0731(.A(mai_mai_n759_), .B(mai_mai_n211_), .Y(mai_mai_n760_));
  NA2        m0732(.A(mai_mai_n536_), .B(mai_mai_n82_), .Y(mai_mai_n761_));
  NO2        m0733(.A(mai_mai_n740_), .B(mai_mai_n761_), .Y(mai_mai_n762_));
  NA3        m0734(.A(mai_mai_n145_), .B(mai_mai_n102_), .C(m), .Y(mai_mai_n763_));
  OAI220     m0735(.A0(mai_mai_n754_), .A1(mai_mai_n383_), .B0(mai_mai_n306_), .B1(mai_mai_n763_), .Y(mai_mai_n764_));
  NOi41      m0736(.An(mai_mai_n200_), .B(mai_mai_n764_), .C(mai_mai_n762_), .D(mai_mai_n278_), .Y(mai_mai_n765_));
  NA2        m0737(.A(c), .B(mai_mai_n110_), .Y(mai_mai_n766_));
  INV        m0738(.A(mai_mai_n766_), .Y(mai_mai_n767_));
  NA3        m0739(.A(mai_mai_n767_), .B(mai_mai_n445_), .C(f), .Y(mai_mai_n768_));
  OR2        m0740(.A(mai_mai_n578_), .B(mai_mai_n478_), .Y(mai_mai_n769_));
  INV        m0741(.A(mai_mai_n769_), .Y(mai_mai_n770_));
  NA2        m0742(.A(mai_mai_n703_), .B(mai_mai_n105_), .Y(mai_mai_n771_));
  NA2        m0743(.A(mai_mai_n771_), .B(mai_mai_n770_), .Y(mai_mai_n772_));
  NA4        m0744(.A(mai_mai_n772_), .B(mai_mai_n768_), .C(mai_mai_n765_), .D(mai_mai_n760_), .Y(mai_mai_n773_));
  NO4        m0745(.A(mai_mai_n773_), .B(mai_mai_n757_), .C(mai_mai_n746_), .D(mai_mai_n736_), .Y(mai_mai_n774_));
  OR2        m0746(.A(mai_mai_n754_), .B(mai_mai_n72_), .Y(mai_mai_n775_));
  NA2        m0747(.A(mai_mai_n723_), .B(m), .Y(mai_mai_n776_));
  AOI210     m0748(.A0(mai_mai_n776_), .A1(mai_mai_n263_), .B0(mai_mai_n775_), .Y(mai_mai_n777_));
  NO2        m0749(.A(mai_mai_n301_), .B(mai_mai_n732_), .Y(mai_mai_n778_));
  NO2        m0750(.A(mai_mai_n383_), .B(mai_mai_n722_), .Y(mai_mai_n779_));
  NA2        m0751(.A(mai_mai_n779_), .B(mai_mai_n496_), .Y(mai_mai_n780_));
  INV        m0752(.A(mai_mai_n780_), .Y(mai_mai_n781_));
  NA2        m0753(.A(e), .B(d), .Y(mai_mai_n782_));
  AOI210     m0754(.A0(mai_mai_n451_), .A1(mai_mai_n162_), .B0(mai_mai_n207_), .Y(mai_mai_n783_));
  INV        m0755(.A(mai_mai_n783_), .Y(mai_mai_n784_));
  NA2        m0756(.A(mai_mai_n256_), .B(mai_mai_n150_), .Y(mai_mai_n785_));
  NA2        m0757(.A(mai_mai_n755_), .B(mai_mai_n785_), .Y(mai_mai_n786_));
  NA3        m0758(.A(mai_mai_n153_), .B(mai_mai_n83_), .C(mai_mai_n34_), .Y(mai_mai_n787_));
  NA3        m0759(.A(mai_mai_n787_), .B(mai_mai_n786_), .C(mai_mai_n784_), .Y(mai_mai_n788_));
  NO4        m0760(.A(mai_mai_n788_), .B(mai_mai_n781_), .C(mai_mai_n778_), .D(mai_mai_n777_), .Y(mai_mai_n789_));
  NA2        m0761(.A(mai_mai_n737_), .B(mai_mai_n31_), .Y(mai_mai_n790_));
  OR2        m0762(.A(mai_mai_n790_), .B(mai_mai_n195_), .Y(mai_mai_n791_));
  NO2        m0763(.A(mai_mai_n553_), .B(mai_mai_n60_), .Y(mai_mai_n792_));
  AOI220     m0764(.A0(mai_mai_n792_), .A1(mai_mai_n758_), .B0(mai_mai_n546_), .B1(mai_mai_n552_), .Y(mai_mai_n793_));
  INV        m0765(.A(mai_mai_n793_), .Y(mai_mai_n794_));
  OAI210     m0766(.A0(mai_mai_n723_), .A1(mai_mai_n785_), .B0(mai_mai_n751_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n795_), .B(mai_mai_n539_), .Y(mai_mai_n796_));
  AOI210     m0768(.A0(mai_mai_n112_), .A1(mai_mai_n111_), .B0(mai_mai_n233_), .Y(mai_mai_n797_));
  AN2        m0769(.A(mai_mai_n739_), .B(mai_mai_n731_), .Y(mai_mai_n798_));
  NOi31      m0770(.An(mai_mai_n482_), .B(mai_mai_n749_), .C(mai_mai_n263_), .Y(mai_mai_n799_));
  NO4        m0771(.A(mai_mai_n799_), .B(mai_mai_n798_), .C(mai_mai_n796_), .D(mai_mai_n794_), .Y(mai_mai_n800_));
  NO2        m0772(.A(mai_mai_n391_), .B(mai_mai_n69_), .Y(mai_mai_n801_));
  OAI210     m0773(.A0(mai_mai_n735_), .A1(mai_mai_n801_), .B0(mai_mai_n616_), .Y(mai_mai_n802_));
  AN3        m0774(.A(mai_mai_n802_), .B(mai_mai_n800_), .C(mai_mai_n791_), .Y(mai_mai_n803_));
  NA4        m0775(.A(mai_mai_n803_), .B(mai_mai_n789_), .C(mai_mai_n774_), .D(mai_mai_n728_), .Y(mai12));
  NO2        m0776(.A(mai_mai_n398_), .B(c), .Y(mai_mai_n805_));
  NO4        m0777(.A(mai_mai_n394_), .B(mai_mai_n226_), .C(mai_mai_n518_), .D(mai_mai_n192_), .Y(mai_mai_n806_));
  NA2        m0778(.A(mai_mai_n806_), .B(mai_mai_n805_), .Y(mai_mai_n807_));
  INV        m0779(.A(mai_mai_n398_), .Y(mai_mai_n808_));
  NO2        m0780(.A(mai_mai_n738_), .B(mai_mai_n318_), .Y(mai_mai_n809_));
  NO2        m0781(.A(mai_mai_n578_), .B(mai_mai_n339_), .Y(mai_mai_n810_));
  AOI220     m0782(.A0(mai_mai_n810_), .A1(mai_mai_n480_), .B0(mai_mai_n809_), .B1(mai_mai_n808_), .Y(mai_mai_n811_));
  NA3        m0783(.A(mai_mai_n811_), .B(mai_mai_n807_), .C(mai_mai_n393_), .Y(mai_mai_n812_));
  AOI210     m0784(.A0(mai_mai_n210_), .A1(mai_mai_n305_), .B0(mai_mai_n181_), .Y(mai_mai_n813_));
  OR2        m0785(.A(mai_mai_n813_), .B(mai_mai_n806_), .Y(mai_mai_n814_));
  NO2        m0786(.A(mai_mai_n346_), .B(mai_mai_n192_), .Y(mai_mai_n815_));
  OAI210     m0787(.A0(mai_mai_n815_), .A1(mai_mai_n814_), .B0(mai_mai_n357_), .Y(mai_mai_n816_));
  NO2        m0788(.A(mai_mai_n564_), .B(mai_mai_n236_), .Y(mai_mai_n817_));
  NO2        m0789(.A(mai_mai_n525_), .B(mai_mai_n730_), .Y(mai_mai_n818_));
  AOI220     m0790(.A0(mai_mai_n818_), .A1(mai_mai_n502_), .B0(mai_mai_n712_), .B1(mai_mai_n817_), .Y(mai_mai_n819_));
  INV        m0791(.A(mai_mai_n213_), .Y(mai_mai_n820_));
  NA2        m0792(.A(mai_mai_n819_), .B(mai_mai_n816_), .Y(mai_mai_n821_));
  NO3        m0793(.A(mai_mai_n583_), .B(mai_mai_n89_), .C(mai_mai_n45_), .Y(mai_mai_n822_));
  NO3        m0794(.A(mai_mai_n822_), .B(mai_mai_n821_), .C(mai_mai_n812_), .Y(mai_mai_n823_));
  NO2        m0795(.A(mai_mai_n330_), .B(mai_mai_n329_), .Y(mai_mai_n824_));
  NA2        m0796(.A(mai_mai_n522_), .B(mai_mai_n71_), .Y(mai_mai_n825_));
  INV        m0797(.A(mai_mai_n136_), .Y(mai_mai_n826_));
  NOi21      m0798(.An(mai_mai_n34_), .B(mai_mai_n573_), .Y(mai_mai_n827_));
  AOI220     m0799(.A0(mai_mai_n827_), .A1(mai_mai_n826_), .B0(mai_mai_n825_), .B1(mai_mai_n824_), .Y(mai_mai_n828_));
  NA2        m0800(.A(mai_mai_n225_), .B(mai_mai_n828_), .Y(mai_mai_n829_));
  NO3        m0801(.A(mai_mai_n713_), .B(mai_mai_n87_), .C(mai_mai_n361_), .Y(mai_mai_n830_));
  NO2        m0802(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n831_));
  NO2        m0803(.A(mai_mai_n440_), .B(mai_mai_n271_), .Y(mai_mai_n832_));
  INV        m0804(.A(mai_mai_n832_), .Y(mai_mai_n833_));
  NO2        m0805(.A(mai_mai_n833_), .B(mai_mai_n136_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n556_), .B(j), .Y(mai_mai_n835_));
  INV        m0807(.A(mai_mai_n327_), .Y(mai_mai_n836_));
  NO4        m0808(.A(mai_mai_n836_), .B(mai_mai_n834_), .C(mai_mai_n830_), .D(mai_mai_n829_), .Y(mai_mai_n837_));
  NA2        m0809(.A(mai_mai_n147_), .B(i), .Y(mai_mai_n838_));
  NA2        m0810(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n839_));
  OAI220     m0811(.A0(mai_mai_n839_), .A1(mai_mai_n180_), .B0(mai_mai_n838_), .B1(mai_mai_n89_), .Y(mai_mai_n840_));
  AOI210     m0812(.A0(mai_mai_n372_), .A1(mai_mai_n37_), .B0(mai_mai_n840_), .Y(mai_mai_n841_));
  NO2        m0813(.A(mai_mai_n841_), .B(mai_mai_n301_), .Y(mai_mai_n842_));
  NA3        m0814(.A(mai_mai_n310_), .B(j), .C(i), .Y(mai_mai_n843_));
  NA2        m0815(.A(mai_mai_n540_), .B(mai_mai_n107_), .Y(mai_mai_n844_));
  NA2        m0816(.A(mai_mai_n603_), .B(mai_mai_n761_), .Y(mai_mai_n845_));
  NA2        m0817(.A(mai_mai_n732_), .B(mai_mai_n392_), .Y(mai_mai_n846_));
  NA2        m0818(.A(mai_mai_n198_), .B(mai_mai_n75_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n847_), .B(mai_mai_n283_), .Y(mai_mai_n848_));
  AOI220     m0820(.A0(mai_mai_n848_), .A1(mai_mai_n231_), .B0(mai_mai_n846_), .B1(mai_mai_n845_), .Y(mai_mai_n849_));
  INV        m0821(.A(mai_mai_n849_), .Y(mai_mai_n850_));
  NO2        m0822(.A(mai_mai_n339_), .B(mai_mai_n88_), .Y(mai_mai_n851_));
  NA2        m0823(.A(mai_mai_n851_), .B(mai_mai_n214_), .Y(mai_mai_n852_));
  NA2        m0824(.A(mai_mai_n582_), .B(mai_mai_n86_), .Y(mai_mai_n853_));
  NA2        m0825(.A(mai_mai_n853_), .B(mai_mai_n852_), .Y(mai_mai_n854_));
  OAI210     m0826(.A0(mai_mai_n846_), .A1(mai_mai_n818_), .B0(mai_mai_n480_), .Y(mai_mai_n855_));
  AOI210     m0827(.A0(mai_mai_n373_), .A1(mai_mai_n365_), .B0(mai_mai_n713_), .Y(mai_mai_n856_));
  OAI210     m0828(.A0(mai_mai_n330_), .A1(mai_mai_n329_), .B0(mai_mai_n103_), .Y(mai_mai_n857_));
  AOI210     m0829(.A0(mai_mai_n857_), .A1(mai_mai_n472_), .B0(mai_mai_n856_), .Y(mai_mai_n858_));
  NO3        m0830(.A(mai_mai_n1279_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n859_));
  AOI220     m0831(.A0(mai_mai_n859_), .A1(mai_mai_n554_), .B0(mai_mai_n569_), .B1(mai_mai_n468_), .Y(mai_mai_n860_));
  NA3        m0832(.A(mai_mai_n860_), .B(mai_mai_n858_), .C(mai_mai_n855_), .Y(mai_mai_n861_));
  NO4        m0833(.A(mai_mai_n861_), .B(mai_mai_n854_), .C(mai_mai_n850_), .D(mai_mai_n842_), .Y(mai_mai_n862_));
  NAi31      m0834(.An(c), .B(mai_mai_n374_), .C(n), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n431_), .B(i), .Y(mai_mai_n864_));
  INV        m0836(.A(mai_mai_n864_), .Y(mai_mai_n865_));
  NA2        m0837(.A(mai_mai_n207_), .B(mai_mai_n157_), .Y(mai_mai_n866_));
  NA2        m0838(.A(mai_mai_n426_), .B(m), .Y(mai_mai_n867_));
  INV        m0839(.A(mai_mai_n867_), .Y(mai_mai_n868_));
  OAI220     m0840(.A0(mai_mai_n863_), .A1(mai_mai_n210_), .B0(mai_mai_n843_), .B1(mai_mai_n537_), .Y(mai_mai_n869_));
  NO2        m0841(.A(mai_mai_n579_), .B(mai_mai_n339_), .Y(mai_mai_n870_));
  NA2        m0842(.A(mai_mai_n813_), .B(mai_mai_n805_), .Y(mai_mai_n871_));
  NO3        m0843(.A(mai_mai_n481_), .B(mai_mai_n140_), .C(mai_mai_n191_), .Y(mai_mai_n872_));
  OAI210     m0844(.A0(mai_mai_n872_), .A1(mai_mai_n462_), .B0(mai_mai_n340_), .Y(mai_mai_n873_));
  OAI220     m0845(.A0(mai_mai_n810_), .A1(mai_mai_n818_), .B0(mai_mai_n482_), .B1(mai_mai_n382_), .Y(mai_mai_n874_));
  NA3        m0846(.A(mai_mai_n874_), .B(mai_mai_n873_), .C(mai_mai_n871_), .Y(mai_mai_n875_));
  OAI210     m0847(.A0(mai_mai_n813_), .A1(mai_mai_n806_), .B0(mai_mai_n866_), .Y(mai_mai_n876_));
  AOI210     m0848(.A0(mai_mai_n342_), .A1(mai_mai_n340_), .B0(mai_mai_n300_), .Y(mai_mai_n877_));
  NA3        m0849(.A(mai_mai_n877_), .B(mai_mai_n876_), .C(mai_mai_n246_), .Y(mai_mai_n878_));
  OR4        m0850(.A(mai_mai_n878_), .B(mai_mai_n875_), .C(mai_mai_n870_), .D(mai_mai_n869_), .Y(mai_mai_n879_));
  NO3        m0851(.A(mai_mai_n879_), .B(mai_mai_n868_), .C(mai_mai_n865_), .Y(mai_mai_n880_));
  NA4        m0852(.A(mai_mai_n880_), .B(mai_mai_n862_), .C(mai_mai_n837_), .D(mai_mai_n823_), .Y(mai13));
  NA3        m0853(.A(mai_mai_n224_), .B(b), .C(m), .Y(mai_mai_n882_));
  NA2        m0854(.A(mai_mai_n435_), .B(f), .Y(mai_mai_n883_));
  NO3        m0855(.A(mai_mai_n883_), .B(mai_mai_n882_), .C(mai_mai_n519_), .Y(mai_mai_n884_));
  NAi32      m0856(.An(d), .Bn(c), .C(e), .Y(mai_mai_n885_));
  NO3        m0857(.A(mai_mai_n885_), .B(mai_mai_n525_), .C(mai_mai_n279_), .Y(mai_mai_n886_));
  NA2        m0858(.A(mai_mai_n586_), .B(mai_mai_n201_), .Y(mai_mai_n887_));
  NA2        m0859(.A(c), .B(mai_mai_n110_), .Y(mai_mai_n888_));
  NO3        m0860(.A(mai_mai_n888_), .B(mai_mai_n160_), .C(mai_mai_n154_), .Y(mai_mai_n889_));
  NA2        m0861(.A(mai_mai_n435_), .B(c), .Y(mai_mai_n890_));
  NO3        m0862(.A(mai_mai_n521_), .B(mai_mai_n890_), .C(mai_mai_n279_), .Y(mai_mai_n891_));
  AO210      m0863(.A0(mai_mai_n889_), .A1(mai_mai_n887_), .B0(mai_mai_n891_), .Y(mai_mai_n892_));
  OR3        m0864(.A(mai_mai_n892_), .B(mai_mai_n886_), .C(mai_mai_n884_), .Y(mai_mai_n893_));
  NAi32      m0865(.An(f), .Bn(e), .C(c), .Y(mai_mai_n894_));
  OR3        m0866(.A(mai_mai_n201_), .B(mai_mai_n160_), .C(mai_mai_n154_), .Y(mai_mai_n895_));
  NO2        m0867(.A(mai_mai_n895_), .B(mai_mai_n894_), .Y(mai_mai_n896_));
  NO2        m0868(.A(mai_mai_n890_), .B(mai_mai_n279_), .Y(mai_mai_n897_));
  NO2        m0869(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n898_));
  NA2        m0870(.A(m), .B(mai_mai_n898_), .Y(mai_mai_n899_));
  NOi21      m0871(.An(mai_mai_n897_), .B(mai_mai_n899_), .Y(mai_mai_n900_));
  NO2        m0872(.A(mai_mai_n663_), .B(mai_mai_n106_), .Y(mai_mai_n901_));
  NOi41      m0873(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n902_));
  NA2        m0874(.A(mai_mai_n902_), .B(mai_mai_n901_), .Y(mai_mai_n903_));
  NO2        m0875(.A(mai_mai_n903_), .B(mai_mai_n894_), .Y(mai_mai_n904_));
  NA3        m0876(.A(k), .B(j), .C(i), .Y(mai_mai_n905_));
  NO3        m0877(.A(mai_mai_n905_), .B(mai_mai_n279_), .C(mai_mai_n88_), .Y(mai_mai_n906_));
  BUFFER     m0878(.A(mai_mai_n906_), .Y(mai_mai_n907_));
  OR4        m0879(.A(mai_mai_n907_), .B(mai_mai_n904_), .C(mai_mai_n900_), .D(mai_mai_n896_), .Y(mai_mai_n908_));
  NA3        m0880(.A(mai_mai_n410_), .B(mai_mai_n303_), .C(mai_mai_n56_), .Y(mai_mai_n909_));
  NO2        m0881(.A(mai_mai_n909_), .B(mai_mai_n899_), .Y(mai_mai_n910_));
  NO2        m0882(.A(mai_mai_n909_), .B(mai_mai_n521_), .Y(mai_mai_n911_));
  NO2        m0883(.A(f), .B(c), .Y(mai_mai_n912_));
  NOi21      m0884(.An(mai_mai_n912_), .B(mai_mai_n394_), .Y(mai_mai_n913_));
  NA2        m0885(.A(mai_mai_n913_), .B(mai_mai_n59_), .Y(mai_mai_n914_));
  NO3        m0886(.A(k), .B(mai_mai_n220_), .C(l), .Y(mai_mai_n915_));
  NOi31      m0887(.An(mai_mai_n915_), .B(mai_mai_n914_), .C(j), .Y(mai_mai_n916_));
  OR3        m0888(.A(mai_mai_n916_), .B(mai_mai_n911_), .C(mai_mai_n910_), .Y(mai_mai_n917_));
  OR3        m0889(.A(mai_mai_n917_), .B(mai_mai_n908_), .C(mai_mai_n893_), .Y(mai02));
  OR2        m0890(.A(l), .B(k), .Y(mai_mai_n919_));
  OR3        m0891(.A(n), .B(m), .C(i), .Y(mai_mai_n920_));
  NO4        m0892(.A(mai_mai_n920_), .B(h), .C(mai_mai_n919_), .D(e), .Y(mai_mai_n921_));
  NO2        m0893(.A(mai_mai_n906_), .B(mai_mai_n886_), .Y(mai_mai_n922_));
  AN3        m0894(.A(m), .B(f), .C(c), .Y(mai_mai_n923_));
  NA2        m0895(.A(mai_mai_n923_), .B(mai_mai_n410_), .Y(mai_mai_n924_));
  OR2        m0896(.A(mai_mai_n905_), .B(mai_mai_n279_), .Y(mai_mai_n925_));
  OR2        m0897(.A(mai_mai_n925_), .B(mai_mai_n924_), .Y(mai_mai_n926_));
  NO2        m0898(.A(mai_mai_n909_), .B(mai_mai_n521_), .Y(mai_mai_n927_));
  NO2        m0899(.A(mai_mai_n927_), .B(mai_mai_n896_), .Y(mai_mai_n928_));
  NA3        m0900(.A(l), .B(k), .C(j), .Y(mai_mai_n929_));
  NA2        m0901(.A(i), .B(h), .Y(mai_mai_n930_));
  NO3        m0902(.A(mai_mai_n930_), .B(mai_mai_n929_), .C(mai_mai_n126_), .Y(mai_mai_n931_));
  NO3        m0903(.A(mai_mai_n135_), .B(mai_mai_n255_), .C(mai_mai_n192_), .Y(mai_mai_n932_));
  AOI210     m0904(.A0(mai_mai_n932_), .A1(mai_mai_n931_), .B0(mai_mai_n900_), .Y(mai_mai_n933_));
  NA3        m0905(.A(c), .B(b), .C(a), .Y(mai_mai_n934_));
  NO3        m0906(.A(mai_mai_n934_), .B(mai_mai_n782_), .C(mai_mai_n191_), .Y(mai_mai_n935_));
  NO3        m0907(.A(mai_mai_n271_), .B(mai_mai_n49_), .C(mai_mai_n106_), .Y(mai_mai_n936_));
  AOI210     m0908(.A0(mai_mai_n936_), .A1(mai_mai_n935_), .B0(mai_mai_n910_), .Y(mai_mai_n937_));
  AN4        m0909(.A(mai_mai_n937_), .B(mai_mai_n933_), .C(mai_mai_n928_), .D(mai_mai_n926_), .Y(mai_mai_n938_));
  INV        m0910(.A(mai_mai_n888_), .Y(mai_mai_n939_));
  NA2        m0911(.A(mai_mai_n903_), .B(mai_mai_n895_), .Y(mai_mai_n940_));
  AOI210     m0912(.A0(mai_mai_n940_), .A1(mai_mai_n939_), .B0(mai_mai_n884_), .Y(mai_mai_n941_));
  NAi41      m0913(.An(mai_mai_n921_), .B(mai_mai_n941_), .C(mai_mai_n938_), .D(mai_mai_n922_), .Y(mai03));
  INV        m0914(.A(mai_mai_n857_), .Y(mai_mai_n943_));
  NO3        m0915(.A(mai_mai_n741_), .B(mai_mai_n733_), .C(mai_mai_n628_), .Y(mai_mai_n944_));
  OAI220     m0916(.A0(mai_mai_n944_), .A1(mai_mai_n603_), .B0(mai_mai_n943_), .B1(mai_mai_n522_), .Y(mai_mai_n945_));
  NOi31      m0917(.An(i), .B(k), .C(j), .Y(mai_mai_n946_));
  NA4        m0918(.A(mai_mai_n946_), .B(e), .C(mai_mai_n310_), .D(mai_mai_n303_), .Y(mai_mai_n947_));
  OAI210     m0919(.A0(mai_mai_n713_), .A1(mai_mai_n375_), .B0(mai_mai_n947_), .Y(mai_mai_n948_));
  NOi31      m0920(.An(m), .B(n), .C(f), .Y(mai_mai_n949_));
  NA2        m0921(.A(mai_mai_n949_), .B(mai_mai_n51_), .Y(mai_mai_n950_));
  AN2        m0922(.A(e), .B(c), .Y(mai_mai_n951_));
  NA2        m0923(.A(mai_mai_n951_), .B(a), .Y(mai_mai_n952_));
  OAI220     m0924(.A0(mai_mai_n952_), .A1(mai_mai_n950_), .B0(mai_mai_n769_), .B1(mai_mai_n381_), .Y(mai_mai_n953_));
  NA2        m0925(.A(mai_mai_n443_), .B(l), .Y(mai_mai_n954_));
  NOi31      m0926(.An(mai_mai_n751_), .B(mai_mai_n882_), .C(mai_mai_n954_), .Y(mai_mai_n955_));
  NO4        m0927(.A(mai_mai_n955_), .B(mai_mai_n953_), .C(mai_mai_n948_), .D(mai_mai_n856_), .Y(mai_mai_n956_));
  INV        m0928(.A(mai_mai_n255_), .Y(mai_mai_n957_));
  INV        m0929(.A(mai_mai_n886_), .Y(mai_mai_n958_));
  NO2        m0930(.A(mai_mai_n85_), .B(m), .Y(mai_mai_n959_));
  AOI210     m0931(.A0(mai_mai_n959_), .A1(i), .B0(mai_mai_n915_), .Y(mai_mai_n960_));
  OR2        m0932(.A(mai_mai_n960_), .B(mai_mai_n914_), .Y(mai_mai_n961_));
  NA3        m0933(.A(mai_mai_n961_), .B(mai_mai_n958_), .C(mai_mai_n956_), .Y(mai_mai_n962_));
  NO4        m0934(.A(mai_mai_n962_), .B(mai_mai_n945_), .C(mai_mai_n714_), .D(mai_mai_n501_), .Y(mai_mai_n963_));
  NA2        m0935(.A(c), .B(b), .Y(mai_mai_n964_));
  NO2        m0936(.A(mai_mai_n615_), .B(mai_mai_n964_), .Y(mai_mai_n965_));
  OAI210     m0937(.A0(mai_mai_n749_), .A1(mai_mai_n726_), .B0(mai_mai_n368_), .Y(mai_mai_n966_));
  OAI210     m0938(.A0(mai_mai_n966_), .A1(mai_mai_n750_), .B0(mai_mai_n965_), .Y(mai_mai_n967_));
  NAi21      m0939(.An(mai_mai_n376_), .B(mai_mai_n965_), .Y(mai_mai_n968_));
  OAI210     m0940(.A0(mai_mai_n486_), .A1(mai_mai_n39_), .B0(mai_mai_n957_), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n969_), .B(mai_mai_n968_), .Y(mai_mai_n970_));
  INV        m0942(.A(mai_mai_n234_), .Y(mai_mai_n971_));
  OAI210     m0943(.A0(mai_mai_n971_), .A1(mai_mai_n257_), .B0(m), .Y(mai_mai_n972_));
  NAi21      m0944(.An(f), .B(d), .Y(mai_mai_n973_));
  NO2        m0945(.A(mai_mai_n973_), .B(mai_mai_n934_), .Y(mai_mai_n974_));
  INV        m0946(.A(mai_mai_n974_), .Y(mai_mai_n975_));
  AOI210     m0947(.A0(mai_mai_n972_), .A1(mai_mai_n263_), .B0(mai_mai_n975_), .Y(mai_mai_n976_));
  AOI210     m0948(.A0(mai_mai_n976_), .A1(mai_mai_n107_), .B0(mai_mai_n970_), .Y(mai_mai_n977_));
  INV        m0949(.A(mai_mai_n412_), .Y(mai_mai_n978_));
  NO2        m0950(.A(mai_mai_n164_), .B(mai_mai_n213_), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n979_), .B(m), .Y(mai_mai_n980_));
  NA3        m0952(.A(mai_mai_n797_), .B(mai_mai_n954_), .C(mai_mai_n415_), .Y(mai_mai_n981_));
  OAI210     m0953(.A0(mai_mai_n981_), .A1(mai_mai_n284_), .B0(mai_mai_n413_), .Y(mai_mai_n982_));
  AOI210     m0954(.A0(mai_mai_n982_), .A1(mai_mai_n978_), .B0(mai_mai_n980_), .Y(mai_mai_n983_));
  NA2        m0955(.A(mai_mai_n496_), .B(mai_mai_n363_), .Y(mai_mai_n984_));
  NA2        m0956(.A(mai_mai_n144_), .B(mai_mai_n33_), .Y(mai_mai_n985_));
  AOI210     m0957(.A0(mai_mai_n835_), .A1(mai_mai_n985_), .B0(mai_mai_n192_), .Y(mai_mai_n986_));
  OAI210     m0958(.A0(mai_mai_n986_), .A1(mai_mai_n395_), .B0(mai_mai_n974_), .Y(mai_mai_n987_));
  AOI210     m0959(.A0(mai_mai_n979_), .A1(mai_mai_n384_), .B0(mai_mai_n830_), .Y(mai_mai_n988_));
  NA3        m0960(.A(mai_mai_n988_), .B(mai_mai_n987_), .C(mai_mai_n984_), .Y(mai_mai_n989_));
  NO2        m0961(.A(mai_mai_n989_), .B(mai_mai_n983_), .Y(mai_mai_n990_));
  NA4        m0962(.A(mai_mai_n990_), .B(mai_mai_n977_), .C(mai_mai_n967_), .D(mai_mai_n963_), .Y(mai00));
  AOI210     m0963(.A0(mai_mai_n270_), .A1(mai_mai_n192_), .B0(mai_mai_n250_), .Y(mai_mai_n992_));
  NO2        m0964(.A(mai_mai_n992_), .B(mai_mai_n514_), .Y(mai_mai_n993_));
  AOI210     m0965(.A0(mai_mai_n779_), .A1(mai_mai_n820_), .B0(mai_mai_n948_), .Y(mai_mai_n994_));
  NO2        m0966(.A(mai_mai_n927_), .B(mai_mai_n830_), .Y(mai_mai_n995_));
  NA3        m0967(.A(mai_mai_n995_), .B(mai_mai_n994_), .C(mai_mai_n858_), .Y(mai_mai_n996_));
  NA2        m0968(.A(mai_mai_n445_), .B(f), .Y(mai_mai_n997_));
  NO2        m0969(.A(mai_mai_n997_), .B(mai_mai_n888_), .Y(mai_mai_n998_));
  NO4        m0970(.A(mai_mai_n998_), .B(mai_mai_n996_), .C(mai_mai_n993_), .D(mai_mai_n908_), .Y(mai_mai_n999_));
  NA2        m0971(.A(mai_mai_n153_), .B(mai_mai_n46_), .Y(mai_mai_n1000_));
  NA3        m0972(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1001_));
  NOi31      m0973(.An(n), .B(m), .C(i), .Y(mai_mai_n1002_));
  NA3        m0974(.A(mai_mai_n1002_), .B(mai_mai_n570_), .C(mai_mai_n51_), .Y(mai_mai_n1003_));
  OAI210     m0975(.A0(mai_mai_n1001_), .A1(mai_mai_n1000_), .B0(mai_mai_n1003_), .Y(mai_mai_n1004_));
  INV        m0976(.A(mai_mai_n513_), .Y(mai_mai_n1005_));
  NO3        m0977(.A(mai_mai_n1005_), .B(mai_mai_n1004_), .C(mai_mai_n799_), .Y(mai_mai_n1006_));
  NO4        m0978(.A(m), .B(mai_mai_n319_), .C(mai_mai_n964_), .D(mai_mai_n59_), .Y(mai_mai_n1007_));
  OR2        m0979(.A(mai_mai_n343_), .B(mai_mai_n129_), .Y(mai_mai_n1008_));
  NO2        m0980(.A(h), .B(m), .Y(mai_mai_n1009_));
  INV        m0981(.A(mai_mai_n1008_), .Y(mai_mai_n1010_));
  NO3        m0982(.A(mai_mai_n1010_), .B(mai_mai_n1007_), .C(mai_mai_n240_), .Y(mai_mai_n1011_));
  NO2        m0983(.A(mai_mai_n215_), .B(mai_mai_n163_), .Y(mai_mai_n1012_));
  NA2        m0984(.A(mai_mai_n1012_), .B(mai_mai_n382_), .Y(mai_mai_n1013_));
  NA3        m0985(.A(mai_mai_n161_), .B(mai_mai_n106_), .C(m), .Y(mai_mai_n1014_));
  NOi21      m0986(.An(mai_mai_n756_), .B(mai_mai_n1014_), .Y(mai_mai_n1015_));
  NAi31      m0987(.An(mai_mai_n168_), .B(mai_mai_n747_), .C(mai_mai_n410_), .Y(mai_mai_n1016_));
  NAi31      m0988(.An(mai_mai_n1015_), .B(mai_mai_n1016_), .C(mai_mai_n1013_), .Y(mai_mai_n1017_));
  INV        m0989(.A(mai_mai_n921_), .Y(mai_mai_n1018_));
  NAi21      m0990(.An(mai_mai_n891_), .B(mai_mai_n1018_), .Y(mai_mai_n1019_));
  NO4        m0991(.A(mai_mai_n1019_), .B(mai_mai_n1017_), .C(mai_mai_n293_), .D(mai_mai_n455_), .Y(mai_mai_n1020_));
  AN3        m0992(.A(mai_mai_n1020_), .B(mai_mai_n1011_), .C(mai_mai_n1006_), .Y(mai_mai_n1021_));
  NA2        m0993(.A(mai_mai_n472_), .B(mai_mai_n97_), .Y(mai_mai_n1022_));
  NA3        m0994(.A(mai_mai_n949_), .B(mai_mai_n540_), .C(mai_mai_n409_), .Y(mai_mai_n1023_));
  NA4        m0995(.A(mai_mai_n1023_), .B(mai_mai_n497_), .C(mai_mai_n1022_), .D(mai_mai_n218_), .Y(mai_mai_n1024_));
  OAI210     m0996(.A0(mai_mai_n408_), .A1(mai_mai_n114_), .B0(mai_mai_n752_), .Y(mai_mai_n1025_));
  AOI220     m0997(.A0(mai_mai_n1025_), .A1(mai_mai_n981_), .B0(mai_mai_n496_), .B1(mai_mai_n363_), .Y(mai_mai_n1026_));
  OR3        m0998(.A(mai_mai_n888_), .B(mai_mai_n199_), .C(e), .Y(mai_mai_n1027_));
  INV        m0999(.A(mai_mai_n137_), .Y(mai_mai_n1028_));
  NA2        m1000(.A(mai_mai_n1028_), .B(mai_mai_n247_), .Y(mai_mai_n1029_));
  NA3        m1001(.A(mai_mai_n1029_), .B(mai_mai_n1027_), .C(mai_mai_n1026_), .Y(mai_mai_n1030_));
  INV        m1002(.A(mai_mai_n714_), .Y(mai_mai_n1031_));
  AOI220     m1003(.A0(mai_mai_n827_), .A1(mai_mai_n512_), .B0(mai_mai_n570_), .B1(mai_mai_n221_), .Y(mai_mai_n1032_));
  NO2        m1004(.A(mai_mai_n67_), .B(h), .Y(mai_mai_n1033_));
  NO2        m1005(.A(mai_mai_n888_), .B(mai_mai_n631_), .Y(mai_mai_n1034_));
  NO2        m1006(.A(mai_mai_n919_), .B(mai_mai_n126_), .Y(mai_mai_n1035_));
  AN2        m1007(.A(mai_mai_n1035_), .B(mai_mai_n932_), .Y(mai_mai_n1036_));
  OAI210     m1008(.A0(mai_mai_n1036_), .A1(mai_mai_n1034_), .B0(mai_mai_n1033_), .Y(mai_mai_n1037_));
  NA4        m1009(.A(mai_mai_n1037_), .B(mai_mai_n1032_), .C(mai_mai_n1031_), .D(mai_mai_n753_), .Y(mai_mai_n1038_));
  NO4        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1030_), .C(mai_mai_n266_), .D(mai_mai_n1024_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n727_), .B(mai_mai_n658_), .Y(mai_mai_n1040_));
  NA4        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1039_), .C(mai_mai_n1021_), .D(mai_mai_n999_), .Y(mai01));
  AN2        m1013(.A(mai_mai_n873_), .B(mai_mai_n871_), .Y(mai_mai_n1042_));
  NO3        m1014(.A(mai_mai_n697_), .B(mai_mai_n689_), .C(mai_mai_n423_), .Y(mai_mai_n1043_));
  NA2        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1042_), .Y(mai_mai_n1044_));
  NA2        m1016(.A(mai_mai_n793_), .B(mai_mai_n302_), .Y(mai_mai_n1045_));
  NA2        m1017(.A(mai_mai_n621_), .B(mai_mai_n92_), .Y(mai_mai_n1046_));
  NO2        m1018(.A(mai_mai_n1046_), .B(mai_mai_n1280_), .Y(mai_mai_n1047_));
  INV        m1019(.A(mai_mai_n112_), .Y(mai_mai_n1048_));
  NO3        m1020(.A(mai_mai_n678_), .B(mai_mai_n592_), .C(mai_mai_n448_), .Y(mai_mai_n1049_));
  NA3        m1021(.A(mai_mai_n621_), .B(mai_mai_n92_), .C(mai_mai_n45_), .Y(mai_mai_n1050_));
  OR2        m1022(.A(mai_mai_n1050_), .B(mai_mai_n589_), .Y(mai_mai_n1051_));
  NA3        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1049_), .C(mai_mai_n132_), .Y(mai_mai_n1052_));
  NO3        m1024(.A(mai_mai_n1052_), .B(mai_mai_n1045_), .C(mai_mai_n1044_), .Y(mai_mai_n1053_));
  NA2        m1025(.A(mai_mai_n273_), .B(mai_mai_n468_), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n475_), .B(mai_mai_n352_), .Y(mai_mai_n1055_));
  NOi21      m1027(.An(mai_mai_n498_), .B(mai_mai_n518_), .Y(mai_mai_n1056_));
  NA2        m1028(.A(mai_mai_n1056_), .B(mai_mai_n1055_), .Y(mai_mai_n1057_));
  AOI210     m1029(.A0(mai_mai_n184_), .A1(mai_mai_n87_), .B0(mai_mai_n191_), .Y(mai_mai_n1058_));
  OAI210     m1030(.A0(mai_mai_n704_), .A1(mai_mai_n382_), .B0(mai_mai_n1058_), .Y(mai_mai_n1059_));
  AN3        m1031(.A(m), .B(l), .C(k), .Y(mai_mai_n1060_));
  OAI210     m1032(.A0(mai_mai_n322_), .A1(mai_mai_n34_), .B0(mai_mai_n1060_), .Y(mai_mai_n1061_));
  NA2        m1033(.A(mai_mai_n183_), .B(mai_mai_n34_), .Y(mai_mai_n1062_));
  AO210      m1034(.A0(mai_mai_n1062_), .A1(mai_mai_n1061_), .B0(mai_mai_n301_), .Y(mai_mai_n1063_));
  NA4        m1035(.A(mai_mai_n1063_), .B(mai_mai_n1059_), .C(mai_mai_n1057_), .D(mai_mai_n1054_), .Y(mai_mai_n1064_));
  INV        m1036(.A(mai_mai_n535_), .Y(mai_mai_n1065_));
  OAI210     m1037(.A0(mai_mai_n1048_), .A1(mai_mai_n529_), .B0(mai_mai_n1065_), .Y(mai_mai_n1066_));
  NA2        m1038(.A(mai_mai_n254_), .B(mai_mai_n176_), .Y(mai_mai_n1067_));
  NA2        m1039(.A(mai_mai_n1067_), .B(mai_mai_n585_), .Y(mai_mai_n1068_));
  NO3        m1040(.A(mai_mai_n713_), .B(mai_mai_n184_), .C(mai_mai_n361_), .Y(mai_mai_n1069_));
  NO2        m1041(.A(mai_mai_n1069_), .B(mai_mai_n830_), .Y(mai_mai_n1070_));
  OAI210     m1042(.A0(mai_mai_n1047_), .A1(mai_mai_n295_), .B0(mai_mai_n593_), .Y(mai_mai_n1071_));
  NA4        m1043(.A(mai_mai_n1071_), .B(mai_mai_n1070_), .C(mai_mai_n1068_), .D(mai_mai_n681_), .Y(mai_mai_n1072_));
  NO3        m1044(.A(mai_mai_n1072_), .B(mai_mai_n1066_), .C(mai_mai_n1064_), .Y(mai_mai_n1073_));
  NA2        m1045(.A(mai_mai_n441_), .B(mai_mai_n58_), .Y(mai_mai_n1074_));
  NO2        m1046(.A(mai_mai_n1050_), .B(mai_mai_n844_), .Y(mai_mai_n1075_));
  NO2        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1004_), .Y(mai_mai_n1076_));
  NA3        m1048(.A(mai_mai_n1076_), .B(mai_mai_n1074_), .C(mai_mai_n657_), .Y(mai_mai_n1077_));
  NO2        m1049(.A(mai_mai_n838_), .B(mai_mai_n209_), .Y(mai_mai_n1078_));
  NO2        m1050(.A(mai_mai_n839_), .B(mai_mai_n492_), .Y(mai_mai_n1079_));
  OAI210     m1051(.A0(mai_mai_n1079_), .A1(mai_mai_n1078_), .B0(mai_mai_n308_), .Y(mai_mai_n1080_));
  NO2        m1052(.A(mai_mai_n331_), .B(mai_mai_n71_), .Y(mai_mai_n1081_));
  INV        m1053(.A(mai_mai_n1081_), .Y(mai_mai_n1082_));
  NA2        m1054(.A(mai_mai_n1082_), .B(mai_mai_n344_), .Y(mai_mai_n1083_));
  NOi31      m1055(.An(mai_mai_n1080_), .B(mai_mai_n1083_), .C(mai_mai_n1077_), .Y(mai_mai_n1084_));
  INV        m1056(.A(mai_mai_n563_), .Y(mai_mai_n1085_));
  NA4        m1057(.A(mai_mai_n1085_), .B(mai_mai_n1084_), .C(mai_mai_n1073_), .D(mai_mai_n1053_), .Y(mai06));
  NO2        m1058(.A(mai_mai_n362_), .B(mai_mai_n495_), .Y(mai_mai_n1087_));
  INV        m1059(.A(mai_mai_n638_), .Y(mai_mai_n1088_));
  OAI210     m1060(.A0(mai_mai_n1088_), .A1(mai_mai_n241_), .B0(mai_mai_n1087_), .Y(mai_mai_n1089_));
  NO3        m1061(.A(mai_mai_n533_), .B(mai_mai_n702_), .C(mai_mai_n536_), .Y(mai_mai_n1090_));
  BUFFER     m1062(.A(mai_mai_n769_), .Y(mai_mai_n1091_));
  NA3        m1063(.A(mai_mai_n1091_), .B(mai_mai_n1089_), .C(mai_mai_n1080_), .Y(mai_mai_n1092_));
  NO2        m1064(.A(mai_mai_n1092_), .B(mai_mai_n229_), .Y(mai_mai_n1093_));
  INV        m1065(.A(mai_mai_n1078_), .Y(mai_mai_n1094_));
  NO2        m1066(.A(mai_mai_n1094_), .B(mai_mai_n305_), .Y(mai_mai_n1095_));
  INV        m1067(.A(mai_mai_n591_), .Y(mai_mai_n1096_));
  NA2        m1068(.A(mai_mai_n1096_), .B(mai_mai_n567_), .Y(mai_mai_n1097_));
  NO2        m1069(.A(mai_mai_n451_), .B(mai_mai_n157_), .Y(mai_mai_n1098_));
  NOi21      m1070(.An(mai_mai_n131_), .B(mai_mai_n45_), .Y(mai_mai_n1099_));
  NO2        m1071(.A(mai_mai_n541_), .B(mai_mai_n950_), .Y(mai_mai_n1100_));
  OAI210     m1072(.A0(mai_mai_n404_), .A1(mai_mai_n223_), .B0(mai_mai_n787_), .Y(mai_mai_n1101_));
  NO4        m1073(.A(mai_mai_n1101_), .B(mai_mai_n1100_), .C(mai_mai_n1099_), .D(mai_mai_n1098_), .Y(mai_mai_n1102_));
  OR2        m1074(.A(mai_mai_n534_), .B(mai_mai_n532_), .Y(mai_mai_n1103_));
  INV        m1075(.A(mai_mai_n1103_), .Y(mai_mai_n1104_));
  NA3        m1076(.A(mai_mai_n1104_), .B(mai_mai_n1102_), .C(mai_mai_n1097_), .Y(mai_mai_n1105_));
  NO2        m1077(.A(mai_mai_n1105_), .B(mai_mai_n1095_), .Y(mai_mai_n1106_));
  OAI220     m1078(.A0(mai_mai_n638_), .A1(mai_mai_n47_), .B0(mai_mai_n201_), .B1(mai_mai_n548_), .Y(mai_mai_n1107_));
  OAI210     m1079(.A0(mai_mai_n251_), .A1(c), .B0(mai_mai_n566_), .Y(mai_mai_n1108_));
  AOI220     m1080(.A0(mai_mai_n1108_), .A1(mai_mai_n1107_), .B0(mai_mai_n46_), .B1(mai_mai_n241_), .Y(mai_mai_n1109_));
  OAI220     m1081(.A0(mai_mai_n612_), .A1(mai_mai_n223_), .B0(mai_mai_n447_), .B1(mai_mai_n451_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(mai_mai_n1110_), .B(mai_mai_n953_), .Y(mai_mai_n1111_));
  NAi31      m1083(.An(mai_mai_n649_), .B(mai_mai_n82_), .C(mai_mai_n183_), .Y(mai_mai_n1112_));
  NA4        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1111_), .C(mai_mai_n1109_), .D(mai_mai_n1032_), .Y(mai_mai_n1113_));
  NOi31      m1085(.An(mai_mai_n1090_), .B(mai_mai_n407_), .C(mai_mai_n351_), .Y(mai_mai_n1114_));
  OR3        m1086(.A(mai_mai_n1114_), .B(mai_mai_n677_), .C(mai_mai_n478_), .Y(mai_mai_n1115_));
  INV        m1087(.A(mai_mai_n1115_), .Y(mai_mai_n1116_));
  AN2        m1088(.A(mai_mai_n806_), .B(mai_mai_n805_), .Y(mai_mai_n1117_));
  NO4        m1089(.A(mai_mai_n1117_), .B(mai_mai_n759_), .C(mai_mai_n437_), .D(mai_mai_n426_), .Y(mai_mai_n1118_));
  INV        m1090(.A(mai_mai_n1118_), .Y(mai_mai_n1119_));
  NAi21      m1091(.An(j), .B(i), .Y(mai_mai_n1120_));
  NO3        m1092(.A(mai_mai_n1119_), .B(mai_mai_n1116_), .C(mai_mai_n1113_), .Y(mai_mai_n1121_));
  NA4        m1093(.A(mai_mai_n1121_), .B(mai_mai_n1106_), .C(mai_mai_n1093_), .D(mai_mai_n1085_), .Y(mai07));
  NA4        m1094(.A(mai_mai_n161_), .B(mai_mai_n102_), .C(j), .D(f), .Y(mai_mai_n1123_));
  NAi32      m1095(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1124_));
  NO3        m1096(.A(mai_mai_n1124_), .B(m), .C(f), .Y(mai_mai_n1125_));
  OAI210     m1097(.A0(mai_mai_n292_), .A1(mai_mai_n427_), .B0(mai_mai_n1125_), .Y(mai_mai_n1126_));
  NAi21      m1098(.An(f), .B(c), .Y(mai_mai_n1127_));
  OR2        m1099(.A(e), .B(d), .Y(mai_mai_n1128_));
  NOi31      m1100(.An(n), .B(m), .C(b), .Y(mai_mai_n1129_));
  NO3        m1101(.A(mai_mai_n126_), .B(mai_mai_n397_), .C(h), .Y(mai_mai_n1130_));
  NA2        m1102(.A(mai_mai_n1126_), .B(mai_mai_n1123_), .Y(mai_mai_n1131_));
  NA2        m1103(.A(mai_mai_n85_), .B(mai_mai_n45_), .Y(mai_mai_n1132_));
  NO2        m1104(.A(mai_mai_n894_), .B(mai_mai_n394_), .Y(mai_mai_n1133_));
  NA3        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1132_), .C(mai_mai_n192_), .Y(mai_mai_n1134_));
  NO2        m1106(.A(mai_mai_n905_), .B(mai_mai_n279_), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n479_), .B(mai_mai_n78_), .Y(mai_mai_n1136_));
  NA2        m1108(.A(mai_mai_n1033_), .B(mai_mai_n261_), .Y(mai_mai_n1137_));
  NA3        m1109(.A(mai_mai_n1137_), .B(mai_mai_n1136_), .C(mai_mai_n1134_), .Y(mai_mai_n1138_));
  NO2        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1131_), .Y(mai_mai_n1139_));
  NO3        m1111(.A(e), .B(d), .C(c), .Y(mai_mai_n1140_));
  NA2        m1112(.A(mai_mai_n1276_), .B(mai_mai_n1140_), .Y(mai_mai_n1141_));
  NO2        m1113(.A(mai_mai_n1141_), .B(mai_mai_n192_), .Y(mai_mai_n1142_));
  NA3        m1114(.A(mai_mai_n609_), .B(mai_mai_n599_), .C(mai_mai_n106_), .Y(mai_mai_n1143_));
  NO2        m1115(.A(mai_mai_n1143_), .B(mai_mai_n45_), .Y(mai_mai_n1144_));
  NO2        m1116(.A(l), .B(k), .Y(mai_mai_n1145_));
  NOi41      m1117(.An(mai_mai_n484_), .B(mai_mai_n1145_), .C(mai_mai_n421_), .D(mai_mai_n394_), .Y(mai_mai_n1146_));
  NO3        m1118(.A(mai_mai_n394_), .B(d), .C(c), .Y(mai_mai_n1147_));
  NO3        m1119(.A(mai_mai_n1146_), .B(mai_mai_n1144_), .C(mai_mai_n1142_), .Y(mai_mai_n1148_));
  NO2        m1120(.A(k), .B(l), .Y(mai_mai_n1149_));
  NO2        m1121(.A(m), .B(c), .Y(mai_mai_n1150_));
  NA2        m1122(.A(mai_mai_n1150_), .B(mai_mai_n169_), .Y(mai_mai_n1151_));
  NO2        m1123(.A(mai_mai_n1151_), .B(mai_mai_n1149_), .Y(mai_mai_n1152_));
  NA2        m1124(.A(mai_mai_n1152_), .B(mai_mai_n161_), .Y(mai_mai_n1153_));
  NO2        m1125(.A(mai_mai_n398_), .B(a), .Y(mai_mai_n1154_));
  NA3        m1126(.A(mai_mai_n1154_), .B(mai_mai_n1278_), .C(mai_mai_n107_), .Y(mai_mai_n1155_));
  NO2        m1127(.A(i), .B(h), .Y(mai_mai_n1156_));
  NA2        m1128(.A(mai_mai_n1156_), .B(mai_mai_n197_), .Y(mai_mai_n1157_));
  AOI210     m1129(.A0(mai_mai_n230_), .A1(mai_mai_n110_), .B0(mai_mai_n468_), .Y(mai_mai_n1158_));
  NO2        m1130(.A(mai_mai_n1158_), .B(mai_mai_n1157_), .Y(mai_mai_n1159_));
  NO2        m1131(.A(mai_mai_n655_), .B(mai_mai_n170_), .Y(mai_mai_n1160_));
  NOi31      m1132(.An(m), .B(n), .C(b), .Y(mai_mai_n1161_));
  NOi31      m1133(.An(f), .B(d), .C(c), .Y(mai_mai_n1162_));
  NA2        m1134(.A(mai_mai_n1162_), .B(mai_mai_n1161_), .Y(mai_mai_n1163_));
  INV        m1135(.A(mai_mai_n1163_), .Y(mai_mai_n1164_));
  NO3        m1136(.A(mai_mai_n1164_), .B(mai_mai_n1160_), .C(mai_mai_n1159_), .Y(mai_mai_n1165_));
  NA2        m1137(.A(mai_mai_n923_), .B(mai_mai_n410_), .Y(mai_mai_n1166_));
  NO4        m1138(.A(mai_mai_n1166_), .B(mai_mai_n901_), .C(mai_mai_n394_), .D(mai_mai_n45_), .Y(mai_mai_n1167_));
  OAI210     m1139(.A0(mai_mai_n164_), .A1(mai_mai_n463_), .B0(mai_mai_n902_), .Y(mai_mai_n1168_));
  INV        m1140(.A(mai_mai_n1168_), .Y(mai_mai_n1169_));
  NO2        m1141(.A(mai_mai_n1169_), .B(mai_mai_n1167_), .Y(mai_mai_n1170_));
  AN4        m1142(.A(mai_mai_n1170_), .B(mai_mai_n1165_), .C(mai_mai_n1155_), .D(mai_mai_n1153_), .Y(mai_mai_n1171_));
  NA2        m1143(.A(mai_mai_n1129_), .B(mai_mai_n341_), .Y(mai_mai_n1172_));
  NO2        m1144(.A(mai_mai_n1172_), .B(mai_mai_n887_), .Y(mai_mai_n1173_));
  NA2        m1145(.A(mai_mai_n931_), .B(mai_mai_n1166_), .Y(mai_mai_n1174_));
  NAi21      m1146(.An(mai_mai_n1173_), .B(mai_mai_n1174_), .Y(mai_mai_n1175_));
  NO4        m1147(.A(mai_mai_n126_), .B(m), .C(f), .D(e), .Y(mai_mai_n1176_));
  INV        m1148(.A(mai_mai_n262_), .Y(mai_mai_n1177_));
  NA2        m1149(.A(mai_mai_n175_), .B(mai_mai_n94_), .Y(mai_mai_n1178_));
  OR2        m1150(.A(e), .B(a), .Y(mai_mai_n1179_));
  OR3        m1151(.A(mai_mai_n478_), .B(mai_mai_n477_), .C(mai_mai_n106_), .Y(mai_mai_n1180_));
  NA2        m1152(.A(mai_mai_n949_), .B(mai_mai_n361_), .Y(mai_mai_n1181_));
  INV        m1153(.A(mai_mai_n1175_), .Y(mai_mai_n1182_));
  NA4        m1154(.A(mai_mai_n1182_), .B(mai_mai_n1171_), .C(mai_mai_n1148_), .D(mai_mai_n1139_), .Y(mai_mai_n1183_));
  NA2        m1155(.A(mai_mai_n341_), .B(mai_mai_n56_), .Y(mai_mai_n1184_));
  NA2        m1156(.A(mai_mai_n193_), .B(mai_mai_n161_), .Y(mai_mai_n1185_));
  AOI210     m1157(.A0(mai_mai_n1185_), .A1(mai_mai_n1014_), .B0(mai_mai_n1184_), .Y(mai_mai_n1186_));
  NO2        m1158(.A(mai_mai_n348_), .B(j), .Y(mai_mai_n1187_));
  NA3        m1159(.A(m), .B(mai_mai_n1187_), .C(mai_mai_n144_), .Y(mai_mai_n1188_));
  NO2        m1160(.A(mai_mai_n1178_), .B(mai_mai_n894_), .Y(mai_mai_n1189_));
  OAI210     m1161(.A0(n), .A1(mai_mai_n912_), .B0(mai_mai_n49_), .Y(mai_mai_n1190_));
  AOI220     m1162(.A0(mai_mai_n1190_), .A1(mai_mai_n1009_), .B0(mai_mai_n717_), .B1(mai_mai_n175_), .Y(mai_mai_n1191_));
  INV        m1163(.A(mai_mai_n1191_), .Y(mai_mai_n1192_));
  OAI220     m1164(.A0(mai_mai_n586_), .A1(m), .B0(mai_mai_n201_), .B1(c), .Y(mai_mai_n1193_));
  INV        m1165(.A(mai_mai_n1193_), .Y(mai_mai_n1194_));
  NO2        m1166(.A(mai_mai_n201_), .B(k), .Y(mai_mai_n1195_));
  NO2        m1167(.A(mai_mai_n1194_), .B(mai_mai_n160_), .Y(mai_mai_n1196_));
  NO3        m1168(.A(mai_mai_n1180_), .B(mai_mai_n410_), .C(mai_mai_n318_), .Y(mai_mai_n1197_));
  NO4        m1169(.A(mai_mai_n1197_), .B(mai_mai_n1196_), .C(mai_mai_n1192_), .D(mai_mai_n1189_), .Y(mai_mai_n1198_));
  NO3        m1170(.A(mai_mai_n934_), .B(mai_mai_n1128_), .C(mai_mai_n49_), .Y(mai_mai_n1199_));
  NO2        m1171(.A(mai_mai_n920_), .B(h), .Y(mai_mai_n1200_));
  NO2        m1172(.A(mai_mai_n1120_), .B(mai_mai_n159_), .Y(mai_mai_n1201_));
  NOi21      m1173(.An(d), .B(f), .Y(mai_mai_n1202_));
  NO2        m1174(.A(mai_mai_n1162_), .B(mai_mai_n1202_), .Y(mai_mai_n1203_));
  NA2        m1175(.A(mai_mai_n1203_), .B(mai_mai_n1201_), .Y(mai_mai_n1204_));
  NO2        m1176(.A(mai_mai_n1128_), .B(f), .Y(mai_mai_n1205_));
  NA4        m1177(.A(mai_mai_n1204_), .B(mai_mai_n1198_), .C(mai_mai_n1188_), .D(mai_mai_n1277_), .Y(mai_mai_n1206_));
  NO3        m1178(.A(mai_mai_n923_), .B(mai_mai_n912_), .C(mai_mai_n40_), .Y(mai_mai_n1207_));
  NO2        m1179(.A(mai_mai_n410_), .B(mai_mai_n271_), .Y(mai_mai_n1208_));
  OAI210     m1180(.A0(mai_mai_n1208_), .A1(mai_mai_n1207_), .B0(mai_mai_n1135_), .Y(mai_mai_n1209_));
  OAI210     m1181(.A0(mai_mai_n1176_), .A1(mai_mai_n1129_), .B0(mai_mai_n766_), .Y(mai_mai_n1210_));
  NO2        m1182(.A(mai_mai_n885_), .B(mai_mai_n126_), .Y(mai_mai_n1211_));
  NA2        m1183(.A(mai_mai_n1211_), .B(mai_mai_n553_), .Y(mai_mai_n1212_));
  NA3        m1184(.A(mai_mai_n1212_), .B(mai_mai_n1210_), .C(mai_mai_n1209_), .Y(mai_mai_n1213_));
  NA2        m1185(.A(mai_mai_n1150_), .B(mai_mai_n1202_), .Y(mai_mai_n1214_));
  NO2        m1186(.A(mai_mai_n1214_), .B(m), .Y(mai_mai_n1215_));
  NO2        m1187(.A(mai_mai_n141_), .B(mai_mai_n163_), .Y(mai_mai_n1216_));
  OAI210     m1188(.A0(mai_mai_n1216_), .A1(mai_mai_n104_), .B0(mai_mai_n1161_), .Y(mai_mai_n1217_));
  INV        m1189(.A(mai_mai_n1217_), .Y(mai_mai_n1218_));
  NO3        m1190(.A(mai_mai_n1218_), .B(mai_mai_n1215_), .C(mai_mai_n1213_), .Y(mai_mai_n1219_));
  NO2        m1191(.A(mai_mai_n1127_), .B(e), .Y(mai_mai_n1220_));
  NA2        m1192(.A(mai_mai_n1220_), .B(mai_mai_n359_), .Y(mai_mai_n1221_));
  OR3        m1193(.A(mai_mai_n1195_), .B(mai_mai_n1033_), .C(mai_mai_n126_), .Y(mai_mai_n1222_));
  NO2        m1194(.A(mai_mai_n1222_), .B(mai_mai_n1221_), .Y(mai_mai_n1223_));
  INV        m1195(.A(mai_mai_n1223_), .Y(mai_mai_n1224_));
  NO2        m1196(.A(mai_mai_n163_), .B(c), .Y(mai_mai_n1225_));
  OAI210     m1197(.A0(mai_mai_n1225_), .A1(mai_mai_n1220_), .B0(mai_mai_n161_), .Y(mai_mai_n1226_));
  AOI220     m1198(.A0(mai_mai_n1226_), .A1(mai_mai_n914_), .B0(mai_mai_n469_), .B1(mai_mai_n329_), .Y(mai_mai_n1227_));
  NA2        m1199(.A(mai_mai_n477_), .B(m), .Y(mai_mai_n1228_));
  AOI210     m1200(.A0(mai_mai_n1228_), .A1(mai_mai_n1147_), .B0(mai_mai_n1199_), .Y(mai_mai_n1229_));
  NO2        m1201(.A(mai_mai_n1179_), .B(f), .Y(mai_mai_n1230_));
  AOI210     m1202(.A0(mai_mai_n959_), .A1(a), .B0(mai_mai_n1230_), .Y(mai_mai_n1231_));
  OAI220     m1203(.A0(mai_mai_n1231_), .A1(mai_mai_n68_), .B0(mai_mai_n1229_), .B1(mai_mai_n191_), .Y(mai_mai_n1232_));
  AOI210     m1204(.A0(mai_mai_n782_), .A1(mai_mai_n371_), .B0(mai_mai_n100_), .Y(mai_mai_n1233_));
  NA2        m1205(.A(mai_mai_n1230_), .B(mai_mai_n1132_), .Y(mai_mai_n1234_));
  OAI220     m1206(.A0(mai_mai_n1234_), .A1(mai_mai_n49_), .B0(mai_mai_n1233_), .B1(mai_mai_n159_), .Y(mai_mai_n1235_));
  NA4        m1207(.A(mai_mai_n932_), .B(mai_mai_n929_), .C(mai_mai_n197_), .D(mai_mai_n67_), .Y(mai_mai_n1236_));
  NA2        m1208(.A(mai_mai_n1130_), .B(mai_mai_n164_), .Y(mai_mai_n1237_));
  NO2        m1209(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1238_));
  OAI210     m1210(.A0(mai_mai_n1179_), .A1(mai_mai_n748_), .B0(mai_mai_n427_), .Y(mai_mai_n1239_));
  OAI210     m1211(.A0(mai_mai_n1239_), .A1(mai_mai_n935_), .B0(mai_mai_n1238_), .Y(mai_mai_n1240_));
  NA3        m1212(.A(mai_mai_n1240_), .B(mai_mai_n1237_), .C(mai_mai_n1236_), .Y(mai_mai_n1241_));
  NO4        m1213(.A(mai_mai_n1241_), .B(mai_mai_n1235_), .C(mai_mai_n1232_), .D(mai_mai_n1227_), .Y(mai_mai_n1242_));
  NA3        m1214(.A(mai_mai_n1242_), .B(mai_mai_n1224_), .C(mai_mai_n1219_), .Y(mai_mai_n1243_));
  NA3        m1215(.A(mai_mai_n831_), .B(mai_mai_n133_), .C(mai_mai_n46_), .Y(mai_mai_n1244_));
  AOI210     m1216(.A0(mai_mai_n139_), .A1(c), .B0(mai_mai_n1244_), .Y(mai_mai_n1245_));
  INV        m1217(.A(mai_mai_n167_), .Y(mai_mai_n1246_));
  NA2        m1218(.A(mai_mai_n1246_), .B(mai_mai_n1200_), .Y(mai_mai_n1247_));
  AO210      m1219(.A0(mai_mai_n127_), .A1(l), .B0(mai_mai_n1172_), .Y(mai_mai_n1248_));
  NO2        m1220(.A(mai_mai_n70_), .B(c), .Y(mai_mai_n1249_));
  NA2        m1221(.A(mai_mai_n1201_), .B(mai_mai_n1249_), .Y(mai_mai_n1250_));
  NA3        m1222(.A(mai_mai_n1250_), .B(mai_mai_n1248_), .C(mai_mai_n1247_), .Y(mai_mai_n1251_));
  NO2        m1223(.A(mai_mai_n1251_), .B(mai_mai_n1245_), .Y(mai_mai_n1252_));
  NO4        m1224(.A(mai_mai_n201_), .B(mai_mai_n168_), .C(mai_mai_n230_), .D(k), .Y(mai_mai_n1253_));
  NOi21      m1225(.An(mai_mai_n1130_), .B(e), .Y(mai_mai_n1254_));
  NO2        m1226(.A(mai_mai_n1254_), .B(mai_mai_n1253_), .Y(mai_mai_n1255_));
  AN2        m1227(.A(mai_mai_n932_), .B(mai_mai_n919_), .Y(mai_mai_n1256_));
  NA2        m1228(.A(mai_mai_n898_), .B(mai_mai_n145_), .Y(mai_mai_n1257_));
  NOi31      m1229(.An(mai_mai_n30_), .B(mai_mai_n1257_), .C(n), .Y(mai_mai_n1258_));
  AOI210     m1230(.A0(mai_mai_n1256_), .A1(mai_mai_n1002_), .B0(mai_mai_n1258_), .Y(mai_mai_n1259_));
  NA2        m1231(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1260_));
  NO2        m1232(.A(mai_mai_n1181_), .B(mai_mai_n1260_), .Y(mai_mai_n1261_));
  INV        m1233(.A(mai_mai_n1261_), .Y(mai_mai_n1262_));
  NA4        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1259_), .C(mai_mai_n1255_), .D(mai_mai_n1252_), .Y(mai_mai_n1263_));
  OR4        m1235(.A(mai_mai_n1263_), .B(mai_mai_n1243_), .C(mai_mai_n1206_), .D(mai_mai_n1183_), .Y(mai04));
  NOi31      m1236(.An(mai_mai_n1176_), .B(mai_mai_n1177_), .C(mai_mai_n888_), .Y(mai_mai_n1265_));
  NA2        m1237(.A(mai_mai_n1205_), .B(mai_mai_n717_), .Y(mai_mai_n1266_));
  NO2        m1238(.A(mai_mai_n1266_), .B(mai_mai_n882_), .Y(mai_mai_n1267_));
  OR3        m1239(.A(mai_mai_n1267_), .B(mai_mai_n1265_), .C(mai_mai_n904_), .Y(mai_mai_n1268_));
  NO2        m1240(.A(mai_mai_n1132_), .B(mai_mai_n88_), .Y(mai_mai_n1269_));
  AOI210     m1241(.A0(mai_mai_n1269_), .A1(mai_mai_n897_), .B0(mai_mai_n1015_), .Y(mai_mai_n1270_));
  NA2        m1242(.A(mai_mai_n1270_), .B(mai_mai_n1037_), .Y(mai_mai_n1271_));
  NO4        m1243(.A(mai_mai_n1271_), .B(mai_mai_n1268_), .C(mai_mai_n911_), .D(mai_mai_n893_), .Y(mai_mai_n1272_));
  NA4        m1244(.A(mai_mai_n1272_), .B(mai_mai_n961_), .C(mai_mai_n947_), .D(mai_mai_n938_), .Y(mai05));
  INV        m1245(.A(m), .Y(mai_mai_n1276_));
  INV        m1246(.A(mai_mai_n1186_), .Y(mai_mai_n1277_));
  INV        m1247(.A(i), .Y(mai_mai_n1278_));
  INV        m1248(.A(j), .Y(mai_mai_n1279_));
  INV        m1249(.A(f), .Y(mai_mai_n1280_));
  INV        m1250(.A(c), .Y(mai_mai_n1281_));
  INV        m1251(.A(f), .Y(mai_mai_n1282_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(u), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(u), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(u), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(u), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(u), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n43_), .B(men_men_n39_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n32_), .Y(men_men_n53_));
  INV        u0025(.A(c), .Y(men_men_n54_));
  NA2        u0026(.A(e), .B(b), .Y(men_men_n55_));
  INV        u0027(.A(d), .Y(men_men_n56_));
  NA2        u0028(.A(u), .B(men_men_n56_), .Y(men_men_n57_));
  NAi21      u0029(.An(i), .B(h), .Y(men_men_n58_));
  NAi31      u0030(.An(i), .B(l), .C(j), .Y(men_men_n59_));
  NO2        u0031(.A(men_men_n58_), .B(men_men_n44_), .Y(men_men_n60_));
  NAi31      u0032(.An(men_men_n57_), .B(men_men_n60_), .C(b), .Y(men_men_n61_));
  NAi41      u0033(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n62_));
  NA2        u0034(.A(u), .B(f), .Y(men_men_n63_));
  NO2        u0035(.A(men_men_n63_), .B(men_men_n62_), .Y(men_men_n64_));
  NAi21      u0036(.An(i), .B(j), .Y(men_men_n65_));
  NAi32      u0037(.An(n), .Bn(k), .C(m), .Y(men_men_n66_));
  NAi31      u0038(.An(l), .B(m), .C(k), .Y(men_men_n67_));
  NAi41      u0039(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n68_));
  INV        u0040(.A(m), .Y(men_men_n69_));
  NOi21      u0041(.An(k), .B(l), .Y(men_men_n70_));
  NA2        u0042(.A(men_men_n70_), .B(men_men_n69_), .Y(men_men_n71_));
  NOi32      u0043(.An(h), .Bn(u), .C(f), .Y(men_men_n72_));
  INV        u0044(.A(men_men_n61_), .Y(men_men_n73_));
  INV        u0045(.A(n), .Y(men_men_n74_));
  NOi32      u0046(.An(e), .Bn(b), .C(d), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  INV        u0048(.A(j), .Y(men_men_n77_));
  AN3        u0049(.A(m), .B(k), .C(i), .Y(men_men_n78_));
  NA3        u0050(.A(men_men_n78_), .B(men_men_n77_), .C(u), .Y(men_men_n79_));
  NO2        u0051(.A(men_men_n79_), .B(f), .Y(men_men_n80_));
  NAi32      u0052(.An(u), .Bn(f), .C(h), .Y(men_men_n81_));
  NAi31      u0053(.An(j), .B(m), .C(l), .Y(men_men_n82_));
  NO2        u0054(.A(men_men_n82_), .B(men_men_n81_), .Y(men_men_n83_));
  NA2        u0055(.A(m), .B(l), .Y(men_men_n84_));
  NAi31      u0056(.An(k), .B(j), .C(u), .Y(men_men_n85_));
  NO3        u0057(.A(men_men_n85_), .B(men_men_n84_), .C(f), .Y(men_men_n86_));
  AN2        u0058(.A(j), .B(u), .Y(men_men_n87_));
  NOi32      u0059(.An(m), .Bn(l), .C(i), .Y(men_men_n88_));
  NOi21      u0060(.An(u), .B(i), .Y(men_men_n89_));
  NOi32      u0061(.An(m), .Bn(j), .C(k), .Y(men_men_n90_));
  AOI220     u0062(.A0(men_men_n90_), .A1(men_men_n89_), .B0(men_men_n88_), .B1(men_men_n87_), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NO4        u0064(.A(men_men_n92_), .B(men_men_n86_), .C(men_men_n83_), .D(men_men_n80_), .Y(men_men_n93_));
  NAi41      u0065(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n94_));
  AN2        u0066(.A(e), .B(b), .Y(men_men_n95_));
  NA2        u0067(.A(c), .B(men_men_n95_), .Y(men_men_n96_));
  NO3        u0068(.A(men_men_n96_), .B(men_men_n94_), .C(u), .Y(men_men_n97_));
  NOi21      u0069(.An(u), .B(f), .Y(men_men_n98_));
  NOi21      u0070(.An(i), .B(h), .Y(men_men_n99_));
  NA3        u0071(.A(men_men_n99_), .B(men_men_n98_), .C(men_men_n36_), .Y(men_men_n100_));
  INV        u0072(.A(a), .Y(men_men_n101_));
  NA2        u0073(.A(men_men_n95_), .B(men_men_n101_), .Y(men_men_n102_));
  INV        u0074(.A(l), .Y(men_men_n103_));
  NOi21      u0075(.An(m), .B(n), .Y(men_men_n104_));
  AN2        u0076(.A(k), .B(h), .Y(men_men_n105_));
  NO2        u0077(.A(men_men_n100_), .B(men_men_n76_), .Y(men_men_n106_));
  INV        u0078(.A(b), .Y(men_men_n107_));
  NA2        u0079(.A(l), .B(j), .Y(men_men_n108_));
  AN2        u0080(.A(k), .B(i), .Y(men_men_n109_));
  NA2        u0081(.A(men_men_n109_), .B(men_men_n108_), .Y(men_men_n110_));
  NA2        u0082(.A(u), .B(e), .Y(men_men_n111_));
  NOi32      u0083(.An(c), .Bn(a), .C(d), .Y(men_men_n112_));
  NA2        u0084(.A(men_men_n112_), .B(men_men_n104_), .Y(men_men_n113_));
  NO3        u0085(.A(men_men_n113_), .B(men_men_n110_), .C(men_men_n107_), .Y(men_men_n114_));
  NO3        u0086(.A(men_men_n114_), .B(men_men_n106_), .C(men_men_n97_), .Y(men_men_n115_));
  OAI210     u0087(.A0(men_men_n93_), .A1(men_men_n76_), .B0(men_men_n115_), .Y(men_men_n116_));
  NOi31      u0088(.An(k), .B(m), .C(j), .Y(men_men_n117_));
  NOi31      u0089(.An(k), .B(m), .C(i), .Y(men_men_n118_));
  NA3        u0090(.A(men_men_n118_), .B(men_men_n72_), .C(e), .Y(men_men_n119_));
  INV        u0091(.A(men_men_n119_), .Y(men_men_n120_));
  NAi21      u0092(.An(u), .B(h), .Y(men_men_n121_));
  NAi21      u0093(.An(m), .B(n), .Y(men_men_n122_));
  NAi41      u0094(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n123_));
  NAi31      u0095(.An(j), .B(k), .C(h), .Y(men_men_n124_));
  NO3        u0096(.A(men_men_n124_), .B(men_men_n123_), .C(men_men_n122_), .Y(men_men_n125_));
  INV        u0097(.A(men_men_n125_), .Y(men_men_n126_));
  NO2        u0098(.A(k), .B(j), .Y(men_men_n127_));
  NO2        u0099(.A(men_men_n127_), .B(men_men_n122_), .Y(men_men_n128_));
  AN2        u0100(.A(k), .B(j), .Y(men_men_n129_));
  NAi21      u0101(.An(c), .B(b), .Y(men_men_n130_));
  NA2        u0102(.A(f), .B(d), .Y(men_men_n131_));
  NO3        u0103(.A(men_men_n131_), .B(men_men_n130_), .C(men_men_n121_), .Y(men_men_n132_));
  NAi31      u0104(.An(f), .B(e), .C(b), .Y(men_men_n133_));
  NA2        u0105(.A(men_men_n132_), .B(men_men_n128_), .Y(men_men_n134_));
  NA2        u0106(.A(d), .B(b), .Y(men_men_n135_));
  NAi21      u0107(.An(e), .B(f), .Y(men_men_n136_));
  NO2        u0108(.A(men_men_n136_), .B(men_men_n135_), .Y(men_men_n137_));
  NA2        u0109(.A(b), .B(a), .Y(men_men_n138_));
  NAi21      u0110(.An(e), .B(u), .Y(men_men_n139_));
  NAi21      u0111(.An(c), .B(d), .Y(men_men_n140_));
  NAi31      u0112(.An(l), .B(k), .C(h), .Y(men_men_n141_));
  NO2        u0113(.A(men_men_n122_), .B(men_men_n141_), .Y(men_men_n142_));
  NA2        u0114(.A(men_men_n142_), .B(men_men_n137_), .Y(men_men_n143_));
  NAi41      u0115(.An(men_men_n120_), .B(men_men_n143_), .C(men_men_n134_), .D(men_men_n126_), .Y(men_men_n144_));
  NAi31      u0116(.An(e), .B(f), .C(b), .Y(men_men_n145_));
  NOi21      u0117(.An(u), .B(d), .Y(men_men_n146_));
  NO2        u0118(.A(men_men_n146_), .B(men_men_n145_), .Y(men_men_n147_));
  NOi21      u0119(.An(h), .B(i), .Y(men_men_n148_));
  NOi21      u0120(.An(k), .B(m), .Y(men_men_n149_));
  NA3        u0121(.A(men_men_n149_), .B(men_men_n148_), .C(n), .Y(men_men_n150_));
  NOi21      u0122(.An(men_men_n147_), .B(men_men_n150_), .Y(men_men_n151_));
  NOi21      u0123(.An(h), .B(u), .Y(men_men_n152_));
  NO2        u0124(.A(men_men_n131_), .B(men_men_n130_), .Y(men_men_n153_));
  NAi31      u0125(.An(l), .B(j), .C(h), .Y(men_men_n154_));
  NO2        u0126(.A(men_men_n154_), .B(men_men_n49_), .Y(men_men_n155_));
  NA2        u0127(.A(men_men_n155_), .B(men_men_n64_), .Y(men_men_n156_));
  NOi32      u0128(.An(n), .Bn(k), .C(m), .Y(men_men_n157_));
  NA2        u0129(.A(l), .B(i), .Y(men_men_n158_));
  INV        u0130(.A(men_men_n156_), .Y(men_men_n159_));
  NAi31      u0131(.An(d), .B(f), .C(c), .Y(men_men_n160_));
  NAi31      u0132(.An(e), .B(f), .C(c), .Y(men_men_n161_));
  NA2        u0133(.A(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  NA2        u0134(.A(j), .B(h), .Y(men_men_n163_));
  OR3        u0135(.A(n), .B(m), .C(k), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  NAi32      u0137(.An(m), .Bn(k), .C(n), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n166_), .B(men_men_n163_), .Y(men_men_n167_));
  AOI220     u0139(.A0(men_men_n167_), .A1(men_men_n147_), .B0(men_men_n165_), .B1(men_men_n162_), .Y(men_men_n168_));
  NO2        u0140(.A(n), .B(m), .Y(men_men_n169_));
  NA2        u0141(.A(men_men_n169_), .B(men_men_n50_), .Y(men_men_n170_));
  NAi21      u0142(.An(f), .B(e), .Y(men_men_n171_));
  NA2        u0143(.A(d), .B(c), .Y(men_men_n172_));
  NAi31      u0144(.An(m), .B(n), .C(b), .Y(men_men_n173_));
  NAi21      u0145(.An(h), .B(f), .Y(men_men_n174_));
  INV        u0146(.A(men_men_n173_), .Y(men_men_n175_));
  NOi32      u0147(.An(f), .Bn(c), .C(d), .Y(men_men_n176_));
  NOi32      u0148(.An(f), .Bn(c), .C(e), .Y(men_men_n177_));
  NO2        u0149(.A(men_men_n177_), .B(men_men_n176_), .Y(men_men_n178_));
  NO3        u0150(.A(n), .B(m), .C(j), .Y(men_men_n179_));
  NA2        u0151(.A(men_men_n179_), .B(men_men_n105_), .Y(men_men_n180_));
  AO210      u0152(.A0(men_men_n180_), .A1(men_men_n170_), .B0(men_men_n178_), .Y(men_men_n181_));
  NA2        u0153(.A(men_men_n181_), .B(men_men_n168_), .Y(men_men_n182_));
  OR4        u0154(.A(men_men_n182_), .B(men_men_n159_), .C(men_men_n151_), .D(men_men_n144_), .Y(men_men_n183_));
  NO4        u0155(.A(men_men_n183_), .B(men_men_n116_), .C(men_men_n73_), .D(men_men_n53_), .Y(men_men_n184_));
  NA3        u0156(.A(m), .B(men_men_n103_), .C(j), .Y(men_men_n185_));
  NAi31      u0157(.An(n), .B(h), .C(u), .Y(men_men_n186_));
  NO2        u0158(.A(men_men_n186_), .B(men_men_n185_), .Y(men_men_n187_));
  NOi32      u0159(.An(m), .Bn(k), .C(l), .Y(men_men_n188_));
  NA3        u0160(.A(men_men_n188_), .B(men_men_n77_), .C(u), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(n), .Y(men_men_n190_));
  NOi21      u0162(.An(k), .B(j), .Y(men_men_n191_));
  NA4        u0163(.A(men_men_n191_), .B(men_men_n104_), .C(i), .D(u), .Y(men_men_n192_));
  NA3        u0164(.A(men_men_n70_), .B(i), .C(men_men_n104_), .Y(men_men_n193_));
  NA2        u0165(.A(men_men_n193_), .B(men_men_n192_), .Y(men_men_n194_));
  NO3        u0166(.A(men_men_n194_), .B(men_men_n190_), .C(men_men_n187_), .Y(men_men_n195_));
  NAi41      u0167(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n196_));
  INV        u0168(.A(men_men_n196_), .Y(men_men_n197_));
  INV        u0169(.A(f), .Y(men_men_n198_));
  INV        u0170(.A(u), .Y(men_men_n199_));
  NOi31      u0171(.An(i), .B(j), .C(h), .Y(men_men_n200_));
  NOi21      u0172(.An(l), .B(m), .Y(men_men_n201_));
  NA2        u0173(.A(men_men_n201_), .B(men_men_n200_), .Y(men_men_n202_));
  NO3        u0174(.A(men_men_n202_), .B(men_men_n199_), .C(men_men_n198_), .Y(men_men_n203_));
  NA2        u0175(.A(men_men_n203_), .B(men_men_n197_), .Y(men_men_n204_));
  OAI210     u0176(.A0(men_men_n195_), .A1(men_men_n32_), .B0(men_men_n204_), .Y(men_men_n205_));
  NOi21      u0177(.An(n), .B(m), .Y(men_men_n206_));
  NOi32      u0178(.An(l), .Bn(i), .C(j), .Y(men_men_n207_));
  NA2        u0179(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  OR2        u0180(.A(men_men_n208_), .B(men_men_n96_), .Y(men_men_n209_));
  NAi21      u0181(.An(j), .B(h), .Y(men_men_n210_));
  XN2        u0182(.A(i), .B(h), .Y(men_men_n211_));
  NOi31      u0183(.An(k), .B(n), .C(m), .Y(men_men_n212_));
  NOi31      u0184(.An(men_men_n212_), .B(men_men_n172_), .C(men_men_n171_), .Y(men_men_n213_));
  INV        u0185(.A(men_men_n213_), .Y(men_men_n214_));
  NAi31      u0186(.An(f), .B(e), .C(c), .Y(men_men_n215_));
  NO4        u0187(.A(men_men_n215_), .B(men_men_n164_), .C(men_men_n163_), .D(men_men_n56_), .Y(men_men_n216_));
  NA4        u0188(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n217_));
  NAi32      u0189(.An(m), .Bn(i), .C(k), .Y(men_men_n218_));
  NO3        u0190(.A(men_men_n218_), .B(men_men_n81_), .C(men_men_n217_), .Y(men_men_n219_));
  INV        u0191(.A(k), .Y(men_men_n220_));
  NO2        u0192(.A(men_men_n219_), .B(men_men_n216_), .Y(men_men_n221_));
  NAi21      u0193(.An(n), .B(a), .Y(men_men_n222_));
  NO2        u0194(.A(men_men_n222_), .B(men_men_n135_), .Y(men_men_n223_));
  NAi41      u0195(.An(u), .B(m), .C(k), .D(h), .Y(men_men_n224_));
  NO2        u0196(.A(men_men_n224_), .B(e), .Y(men_men_n225_));
  NO3        u0197(.A(men_men_n136_), .B(men_men_n85_), .C(men_men_n84_), .Y(men_men_n226_));
  OAI210     u0198(.A0(men_men_n226_), .A1(men_men_n225_), .B0(men_men_n223_), .Y(men_men_n227_));
  AN4        u0199(.A(men_men_n227_), .B(men_men_n221_), .C(men_men_n214_), .D(men_men_n209_), .Y(men_men_n228_));
  NAi41      u0200(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n229_));
  NO2        u0201(.A(men_men_n229_), .B(men_men_n198_), .Y(men_men_n230_));
  NA2        u0202(.A(men_men_n149_), .B(men_men_n99_), .Y(men_men_n231_));
  NAi21      u0203(.An(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  NO2        u0204(.A(n), .B(a), .Y(men_men_n233_));
  NAi31      u0205(.An(men_men_n224_), .B(men_men_n233_), .C(men_men_n95_), .Y(men_men_n234_));
  AN2        u0206(.A(men_men_n234_), .B(men_men_n232_), .Y(men_men_n235_));
  NAi21      u0207(.An(h), .B(i), .Y(men_men_n236_));
  NA2        u0208(.A(men_men_n169_), .B(k), .Y(men_men_n237_));
  NO2        u0209(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  NA2        u0210(.A(men_men_n238_), .B(men_men_n176_), .Y(men_men_n239_));
  NA2        u0211(.A(men_men_n239_), .B(men_men_n235_), .Y(men_men_n240_));
  NO2        u0212(.A(men_men_n68_), .B(men_men_n69_), .Y(men_men_n241_));
  NOi32      u0213(.An(l), .Bn(j), .C(i), .Y(men_men_n242_));
  NO2        u0214(.A(men_men_n236_), .B(men_men_n44_), .Y(men_men_n243_));
  NAi21      u0215(.An(f), .B(u), .Y(men_men_n244_));
  NO2        u0216(.A(men_men_n244_), .B(men_men_n62_), .Y(men_men_n245_));
  NO2        u0217(.A(men_men_n66_), .B(men_men_n108_), .Y(men_men_n246_));
  AOI220     u0218(.A0(men_men_n246_), .A1(men_men_n245_), .B0(men_men_n243_), .B1(men_men_n64_), .Y(men_men_n247_));
  INV        u0219(.A(men_men_n247_), .Y(men_men_n248_));
  NO3        u0220(.A(j), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n249_));
  NOi41      u0221(.An(men_men_n228_), .B(men_men_n248_), .C(men_men_n240_), .D(men_men_n205_), .Y(men_men_n250_));
  NO4        u0222(.A(men_men_n187_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n251_));
  NO2        u0223(.A(men_men_n251_), .B(men_men_n102_), .Y(men_men_n252_));
  NA3        u0224(.A(men_men_n56_), .B(c), .C(b), .Y(men_men_n253_));
  NAi21      u0225(.An(h), .B(u), .Y(men_men_n254_));
  OR3        u0226(.A(men_men_n254_), .B(men_men_n253_), .C(men_men_n208_), .Y(men_men_n255_));
  NAi31      u0227(.An(u), .B(k), .C(h), .Y(men_men_n256_));
  NO3        u0228(.A(men_men_n122_), .B(men_men_n256_), .C(l), .Y(men_men_n257_));
  NAi31      u0229(.An(e), .B(d), .C(a), .Y(men_men_n258_));
  NA2        u0230(.A(men_men_n257_), .B(b), .Y(men_men_n259_));
  NA2        u0231(.A(men_men_n259_), .B(men_men_n255_), .Y(men_men_n260_));
  NA4        u0232(.A(men_men_n149_), .B(men_men_n72_), .C(e), .D(men_men_n108_), .Y(men_men_n261_));
  NA3        u0233(.A(men_men_n149_), .B(men_men_n148_), .C(men_men_n74_), .Y(men_men_n262_));
  NO2        u0234(.A(men_men_n262_), .B(men_men_n178_), .Y(men_men_n263_));
  NOi21      u0235(.An(men_men_n261_), .B(men_men_n263_), .Y(men_men_n264_));
  NA3        u0236(.A(e), .B(c), .C(b), .Y(men_men_n265_));
  NO2        u0237(.A(men_men_n57_), .B(men_men_n265_), .Y(men_men_n266_));
  NAi32      u0238(.An(k), .Bn(i), .C(j), .Y(men_men_n267_));
  NAi31      u0239(.An(h), .B(l), .C(i), .Y(men_men_n268_));
  NA3        u0240(.A(men_men_n268_), .B(men_men_n267_), .C(men_men_n154_), .Y(men_men_n269_));
  NOi21      u0241(.An(men_men_n269_), .B(men_men_n49_), .Y(men_men_n270_));
  OAI210     u0242(.A0(men_men_n245_), .A1(men_men_n266_), .B0(men_men_n270_), .Y(men_men_n271_));
  NAi21      u0243(.An(l), .B(k), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n272_), .B(men_men_n49_), .Y(men_men_n273_));
  NOi21      u0245(.An(l), .B(j), .Y(men_men_n274_));
  NA2        u0246(.A(men_men_n152_), .B(men_men_n274_), .Y(men_men_n275_));
  NA3        u0247(.A(men_men_n109_), .B(men_men_n108_), .C(u), .Y(men_men_n276_));
  OR3        u0248(.A(men_men_n68_), .B(men_men_n69_), .C(e), .Y(men_men_n277_));
  AOI210     u0249(.A0(men_men_n276_), .A1(men_men_n275_), .B0(men_men_n277_), .Y(men_men_n278_));
  INV        u0250(.A(men_men_n278_), .Y(men_men_n279_));
  NAi32      u0251(.An(j), .Bn(h), .C(i), .Y(men_men_n280_));
  NAi21      u0252(.An(m), .B(l), .Y(men_men_n281_));
  NO3        u0253(.A(men_men_n281_), .B(men_men_n280_), .C(men_men_n74_), .Y(men_men_n282_));
  NA2        u0254(.A(h), .B(u), .Y(men_men_n283_));
  NA2        u0255(.A(men_men_n157_), .B(men_men_n45_), .Y(men_men_n284_));
  NO2        u0256(.A(men_men_n284_), .B(men_men_n283_), .Y(men_men_n285_));
  OAI210     u0257(.A0(men_men_n285_), .A1(men_men_n282_), .B0(men_men_n153_), .Y(men_men_n286_));
  NA4        u0258(.A(men_men_n286_), .B(men_men_n279_), .C(men_men_n271_), .D(men_men_n264_), .Y(men_men_n287_));
  NO2        u0259(.A(men_men_n133_), .B(d), .Y(men_men_n288_));
  NAi32      u0260(.An(n), .Bn(m), .C(l), .Y(men_men_n289_));
  NO2        u0261(.A(men_men_n289_), .B(men_men_n280_), .Y(men_men_n290_));
  NO2        u0262(.A(men_men_n113_), .B(men_men_n107_), .Y(men_men_n291_));
  NAi31      u0263(.An(k), .B(l), .C(j), .Y(men_men_n292_));
  OAI210     u0264(.A0(men_men_n272_), .A1(j), .B0(men_men_n292_), .Y(men_men_n293_));
  NOi21      u0265(.An(men_men_n293_), .B(men_men_n111_), .Y(men_men_n294_));
  NA2        u0266(.A(men_men_n294_), .B(men_men_n291_), .Y(men_men_n295_));
  INV        u0267(.A(men_men_n295_), .Y(men_men_n296_));
  NO4        u0268(.A(men_men_n296_), .B(men_men_n287_), .C(men_men_n260_), .D(men_men_n252_), .Y(men_men_n297_));
  NAi21      u0269(.An(m), .B(k), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n211_), .B(men_men_n298_), .Y(men_men_n299_));
  NAi41      u0271(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n300_));
  INV        u0272(.A(men_men_n300_), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n301_), .B(men_men_n299_), .Y(men_men_n302_));
  NO4        u0274(.A(i), .B(men_men_n139_), .C(men_men_n68_), .D(men_men_n69_), .Y(men_men_n303_));
  NA2        u0275(.A(e), .B(c), .Y(men_men_n304_));
  NO3        u0276(.A(men_men_n304_), .B(n), .C(d), .Y(men_men_n305_));
  NAi31      u0277(.An(d), .B(e), .C(b), .Y(men_men_n306_));
  NAi21      u0278(.An(men_men_n303_), .B(men_men_n302_), .Y(men_men_n307_));
  NA2        u0279(.A(men_men_n233_), .B(men_men_n95_), .Y(men_men_n308_));
  OR2        u0280(.A(men_men_n308_), .B(men_men_n189_), .Y(men_men_n309_));
  NOi31      u0281(.An(l), .B(n), .C(m), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n310_), .B(men_men_n200_), .Y(men_men_n311_));
  NO2        u0283(.A(men_men_n311_), .B(men_men_n178_), .Y(men_men_n312_));
  NAi21      u0284(.An(men_men_n312_), .B(men_men_n309_), .Y(men_men_n313_));
  NAi32      u0285(.An(m), .Bn(j), .C(k), .Y(men_men_n314_));
  NAi41      u0286(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n315_));
  NOi31      u0287(.An(j), .B(m), .C(k), .Y(men_men_n316_));
  NO2        u0288(.A(men_men_n117_), .B(men_men_n316_), .Y(men_men_n317_));
  AN3        u0289(.A(h), .B(u), .C(f), .Y(men_men_n318_));
  NOi32      u0290(.An(m), .Bn(j), .C(l), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n319_), .B(men_men_n88_), .Y(men_men_n320_));
  NAi32      u0292(.An(men_men_n320_), .Bn(men_men_n186_), .C(men_men_n288_), .Y(men_men_n321_));
  NO2        u0293(.A(men_men_n281_), .B(men_men_n280_), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n202_), .B(u), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n145_), .B(men_men_n74_), .Y(men_men_n324_));
  AOI220     u0296(.A0(men_men_n324_), .A1(men_men_n323_), .B0(men_men_n230_), .B1(men_men_n322_), .Y(men_men_n325_));
  INV        u0297(.A(men_men_n218_), .Y(men_men_n326_));
  NA3        u0298(.A(men_men_n326_), .B(men_men_n318_), .C(men_men_n197_), .Y(men_men_n327_));
  NA3        u0299(.A(men_men_n327_), .B(men_men_n325_), .C(men_men_n321_), .Y(men_men_n328_));
  NA3        u0300(.A(h), .B(u), .C(f), .Y(men_men_n329_));
  NO2        u0301(.A(men_men_n329_), .B(men_men_n71_), .Y(men_men_n330_));
  NA2        u0302(.A(men_men_n315_), .B(men_men_n196_), .Y(men_men_n331_));
  NA2        u0303(.A(men_men_n152_), .B(e), .Y(men_men_n332_));
  NO2        u0304(.A(men_men_n332_), .B(men_men_n41_), .Y(men_men_n333_));
  AOI220     u0305(.A0(men_men_n333_), .A1(men_men_n291_), .B0(men_men_n331_), .B1(men_men_n330_), .Y(men_men_n334_));
  NOi32      u0306(.An(j), .Bn(u), .C(i), .Y(men_men_n335_));
  NA3        u0307(.A(men_men_n335_), .B(men_men_n272_), .C(men_men_n104_), .Y(men_men_n336_));
  AO210      u0308(.A0(men_men_n102_), .A1(men_men_n32_), .B0(men_men_n336_), .Y(men_men_n337_));
  NOi32      u0309(.An(e), .Bn(b), .C(a), .Y(men_men_n338_));
  AN2        u0310(.A(l), .B(j), .Y(men_men_n339_));
  NA3        u0311(.A(men_men_n193_), .B(men_men_n192_), .C(men_men_n35_), .Y(men_men_n340_));
  NA2        u0312(.A(men_men_n340_), .B(men_men_n338_), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n306_), .B(n), .Y(men_men_n342_));
  NA2        u0314(.A(i), .B(k), .Y(men_men_n343_));
  NA3        u0315(.A(m), .B(men_men_n103_), .C(men_men_n198_), .Y(men_men_n344_));
  NA4        u0316(.A(men_men_n188_), .B(men_men_n77_), .C(u), .D(men_men_n198_), .Y(men_men_n345_));
  OAI210     u0317(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n345_), .Y(men_men_n346_));
  NAi41      u0318(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n347_));
  NA2        u0319(.A(men_men_n51_), .B(men_men_n104_), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n348_), .B(men_men_n347_), .Y(men_men_n349_));
  AOI220     u0321(.A0(men_men_n349_), .A1(b), .B0(men_men_n346_), .B1(men_men_n342_), .Y(men_men_n350_));
  NA4        u0322(.A(men_men_n350_), .B(men_men_n341_), .C(men_men_n337_), .D(men_men_n334_), .Y(men_men_n351_));
  NO4        u0323(.A(men_men_n351_), .B(men_men_n328_), .C(men_men_n313_), .D(men_men_n307_), .Y(men_men_n352_));
  NA4        u0324(.A(men_men_n352_), .B(men_men_n297_), .C(men_men_n250_), .D(men_men_n184_), .Y(men10));
  NA3        u0325(.A(m), .B(k), .C(i), .Y(men_men_n354_));
  NO3        u0326(.A(men_men_n354_), .B(j), .C(men_men_n199_), .Y(men_men_n355_));
  NOi21      u0327(.An(e), .B(f), .Y(men_men_n356_));
  NO4        u0328(.A(men_men_n140_), .B(men_men_n356_), .C(n), .D(men_men_n101_), .Y(men_men_n357_));
  NAi31      u0329(.An(b), .B(f), .C(c), .Y(men_men_n358_));
  INV        u0330(.A(men_men_n358_), .Y(men_men_n359_));
  NOi32      u0331(.An(k), .Bn(h), .C(j), .Y(men_men_n360_));
  NA2        u0332(.A(men_men_n360_), .B(men_men_n206_), .Y(men_men_n361_));
  NA2        u0333(.A(men_men_n150_), .B(men_men_n361_), .Y(men_men_n362_));
  AOI220     u0334(.A0(men_men_n362_), .A1(men_men_n359_), .B0(men_men_n357_), .B1(men_men_n355_), .Y(men_men_n363_));
  AN2        u0335(.A(j), .B(h), .Y(men_men_n364_));
  OR2        u0336(.A(m), .B(k), .Y(men_men_n365_));
  NO2        u0337(.A(men_men_n163_), .B(men_men_n365_), .Y(men_men_n366_));
  NA4        u0338(.A(n), .B(f), .C(c), .D(men_men_n107_), .Y(men_men_n367_));
  NOi21      u0339(.An(men_men_n366_), .B(men_men_n367_), .Y(men_men_n368_));
  NOi32      u0340(.An(d), .Bn(a), .C(c), .Y(men_men_n369_));
  NA2        u0341(.A(men_men_n369_), .B(men_men_n171_), .Y(men_men_n370_));
  NAi21      u0342(.An(i), .B(u), .Y(men_men_n371_));
  NAi31      u0343(.An(k), .B(m), .C(j), .Y(men_men_n372_));
  NO3        u0344(.A(men_men_n372_), .B(men_men_n371_), .C(n), .Y(men_men_n373_));
  NOi21      u0345(.An(men_men_n373_), .B(men_men_n370_), .Y(men_men_n374_));
  NO2        u0346(.A(men_men_n374_), .B(men_men_n368_), .Y(men_men_n375_));
  NO2        u0347(.A(men_men_n367_), .B(men_men_n281_), .Y(men_men_n376_));
  NOi32      u0348(.An(f), .Bn(d), .C(c), .Y(men_men_n377_));
  AOI220     u0349(.A0(men_men_n377_), .A1(men_men_n290_), .B0(men_men_n376_), .B1(men_men_n200_), .Y(men_men_n378_));
  NA2        u0350(.A(men_men_n375_), .B(men_men_n363_), .Y(men_men_n379_));
  NO2        u0351(.A(men_men_n56_), .B(men_men_n107_), .Y(men_men_n380_));
  NA2        u0352(.A(men_men_n233_), .B(men_men_n380_), .Y(men_men_n381_));
  INV        u0353(.A(e), .Y(men_men_n382_));
  NA2        u0354(.A(men_men_n46_), .B(e), .Y(men_men_n383_));
  OAI220     u0355(.A0(men_men_n383_), .A1(men_men_n185_), .B0(men_men_n189_), .B1(men_men_n382_), .Y(men_men_n384_));
  AN2        u0356(.A(u), .B(e), .Y(men_men_n385_));
  NA3        u0357(.A(men_men_n385_), .B(men_men_n188_), .C(i), .Y(men_men_n386_));
  OAI210     u0358(.A0(men_men_n79_), .A1(men_men_n382_), .B0(men_men_n386_), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n91_), .B(men_men_n382_), .Y(men_men_n388_));
  NO3        u0360(.A(men_men_n388_), .B(men_men_n387_), .C(men_men_n384_), .Y(men_men_n389_));
  NOi32      u0361(.An(h), .Bn(e), .C(u), .Y(men_men_n390_));
  NA3        u0362(.A(men_men_n390_), .B(men_men_n274_), .C(m), .Y(men_men_n391_));
  NOi21      u0363(.An(u), .B(h), .Y(men_men_n392_));
  AN3        u0364(.A(m), .B(l), .C(i), .Y(men_men_n393_));
  NA3        u0365(.A(men_men_n393_), .B(men_men_n392_), .C(e), .Y(men_men_n394_));
  AN3        u0366(.A(h), .B(u), .C(e), .Y(men_men_n395_));
  NA2        u0367(.A(men_men_n395_), .B(men_men_n88_), .Y(men_men_n396_));
  AN3        u0368(.A(men_men_n396_), .B(men_men_n394_), .C(men_men_n391_), .Y(men_men_n397_));
  AOI210     u0369(.A0(men_men_n397_), .A1(men_men_n389_), .B0(men_men_n381_), .Y(men_men_n398_));
  NA3        u0370(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n399_));
  NO2        u0371(.A(men_men_n399_), .B(men_men_n381_), .Y(men_men_n400_));
  NA3        u0372(.A(men_men_n369_), .B(men_men_n171_), .C(men_men_n74_), .Y(men_men_n401_));
  NAi31      u0373(.An(b), .B(c), .C(a), .Y(men_men_n402_));
  NO2        u0374(.A(men_men_n402_), .B(n), .Y(men_men_n403_));
  OAI210     u0375(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n404_));
  NO2        u0376(.A(men_men_n404_), .B(men_men_n136_), .Y(men_men_n405_));
  NO3        u0377(.A(men_men_n400_), .B(men_men_n398_), .C(men_men_n379_), .Y(men_men_n406_));
  NA2        u0378(.A(i), .B(u), .Y(men_men_n407_));
  NO3        u0379(.A(men_men_n258_), .B(men_men_n407_), .C(c), .Y(men_men_n408_));
  NOi21      u0380(.An(a), .B(n), .Y(men_men_n409_));
  NOi21      u0381(.An(d), .B(c), .Y(men_men_n410_));
  NA2        u0382(.A(men_men_n410_), .B(men_men_n409_), .Y(men_men_n411_));
  NA3        u0383(.A(i), .B(u), .C(f), .Y(men_men_n412_));
  OR2        u0384(.A(men_men_n412_), .B(men_men_n67_), .Y(men_men_n413_));
  NA3        u0385(.A(men_men_n393_), .B(men_men_n392_), .C(men_men_n171_), .Y(men_men_n414_));
  AOI210     u0386(.A0(men_men_n414_), .A1(men_men_n413_), .B0(men_men_n411_), .Y(men_men_n415_));
  AOI210     u0387(.A0(men_men_n408_), .A1(men_men_n273_), .B0(men_men_n415_), .Y(men_men_n416_));
  OR2        u0388(.A(n), .B(m), .Y(men_men_n417_));
  NO2        u0389(.A(men_men_n417_), .B(men_men_n141_), .Y(men_men_n418_));
  NO2        u0390(.A(men_men_n172_), .B(men_men_n136_), .Y(men_men_n419_));
  OAI210     u0391(.A0(men_men_n418_), .A1(men_men_n165_), .B0(men_men_n419_), .Y(men_men_n420_));
  INV        u0392(.A(men_men_n348_), .Y(men_men_n421_));
  NA3        u0393(.A(men_men_n421_), .B(men_men_n338_), .C(d), .Y(men_men_n422_));
  NO2        u0394(.A(men_men_n402_), .B(men_men_n49_), .Y(men_men_n423_));
  NAi21      u0395(.An(k), .B(j), .Y(men_men_n424_));
  NAi21      u0396(.An(e), .B(d), .Y(men_men_n425_));
  NO2        u0397(.A(men_men_n237_), .B(men_men_n198_), .Y(men_men_n426_));
  NA2        u0398(.A(men_men_n422_), .B(men_men_n420_), .Y(men_men_n427_));
  INV        u0399(.A(men_men_n311_), .Y(men_men_n428_));
  NA2        u0400(.A(men_men_n428_), .B(d), .Y(men_men_n429_));
  NOi31      u0401(.An(n), .B(m), .C(k), .Y(men_men_n430_));
  AOI220     u0402(.A0(men_men_n430_), .A1(men_men_n364_), .B0(men_men_n206_), .B1(men_men_n50_), .Y(men_men_n431_));
  NAi31      u0403(.An(u), .B(f), .C(c), .Y(men_men_n432_));
  OR2        u0404(.A(men_men_n432_), .B(men_men_n431_), .Y(men_men_n433_));
  NA2        u0405(.A(men_men_n433_), .B(men_men_n429_), .Y(men_men_n434_));
  NOi41      u0406(.An(men_men_n416_), .B(men_men_n434_), .C(men_men_n427_), .D(men_men_n248_), .Y(men_men_n435_));
  NOi32      u0407(.An(c), .Bn(a), .C(b), .Y(men_men_n436_));
  NA2        u0408(.A(men_men_n436_), .B(men_men_n104_), .Y(men_men_n437_));
  AN2        u0409(.A(e), .B(d), .Y(men_men_n438_));
  INV        u0410(.A(men_men_n136_), .Y(men_men_n439_));
  NO2        u0411(.A(men_men_n121_), .B(men_men_n41_), .Y(men_men_n440_));
  NO2        u0412(.A(men_men_n63_), .B(e), .Y(men_men_n441_));
  NOi31      u0413(.An(j), .B(k), .C(i), .Y(men_men_n442_));
  NOi21      u0414(.An(men_men_n154_), .B(men_men_n442_), .Y(men_men_n443_));
  AOI210     u0415(.A0(men_men_n440_), .A1(men_men_n439_), .B0(men_men_n441_), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n444_), .B(men_men_n437_), .Y(men_men_n445_));
  NO2        u0417(.A(men_men_n194_), .B(men_men_n190_), .Y(men_men_n446_));
  NOi21      u0418(.An(a), .B(b), .Y(men_men_n447_));
  NA3        u0419(.A(e), .B(d), .C(c), .Y(men_men_n448_));
  NAi21      u0420(.An(men_men_n448_), .B(men_men_n447_), .Y(men_men_n449_));
  AOI210     u0421(.A0(men_men_n251_), .A1(men_men_n446_), .B0(men_men_n449_), .Y(men_men_n450_));
  NA2        u0422(.A(men_men_n359_), .B(men_men_n142_), .Y(men_men_n451_));
  OR2        u0423(.A(k), .B(j), .Y(men_men_n452_));
  NA2        u0424(.A(l), .B(k), .Y(men_men_n453_));
  AOI210     u0425(.A0(men_men_n218_), .A1(men_men_n314_), .B0(men_men_n74_), .Y(men_men_n454_));
  NA2        u0426(.A(men_men_n261_), .B(men_men_n119_), .Y(men_men_n455_));
  NA2        u0427(.A(men_men_n369_), .B(men_men_n104_), .Y(men_men_n456_));
  NO4        u0428(.A(men_men_n456_), .B(men_men_n85_), .C(men_men_n103_), .D(e), .Y(men_men_n457_));
  NO3        u0429(.A(men_men_n401_), .B(men_men_n82_), .C(men_men_n121_), .Y(men_men_n458_));
  NO4        u0430(.A(men_men_n458_), .B(men_men_n457_), .C(men_men_n455_), .D(men_men_n303_), .Y(men_men_n459_));
  NA2        u0431(.A(men_men_n459_), .B(men_men_n451_), .Y(men_men_n460_));
  NO3        u0432(.A(men_men_n460_), .B(men_men_n450_), .C(men_men_n445_), .Y(men_men_n461_));
  NO2        u0433(.A(men_men_n174_), .B(men_men_n54_), .Y(men_men_n462_));
  NAi31      u0434(.An(j), .B(l), .C(i), .Y(men_men_n463_));
  OAI210     u0435(.A0(men_men_n463_), .A1(men_men_n122_), .B0(men_men_n94_), .Y(men_men_n464_));
  NA2        u0436(.A(men_men_n464_), .B(men_men_n462_), .Y(men_men_n465_));
  NO3        u0437(.A(men_men_n370_), .B(men_men_n320_), .C(men_men_n186_), .Y(men_men_n466_));
  NO2        u0438(.A(men_men_n370_), .B(men_men_n348_), .Y(men_men_n467_));
  NO2        u0439(.A(men_men_n467_), .B(men_men_n466_), .Y(men_men_n468_));
  NA3        u0440(.A(men_men_n468_), .B(men_men_n465_), .C(men_men_n228_), .Y(men_men_n469_));
  OAI210     u0441(.A0(men_men_n118_), .A1(men_men_n117_), .B0(n), .Y(men_men_n470_));
  NO2        u0442(.A(men_men_n470_), .B(men_men_n121_), .Y(men_men_n471_));
  AN2        u0443(.A(men_men_n471_), .B(men_men_n177_), .Y(men_men_n472_));
  XO2        u0444(.A(i), .B(h), .Y(men_men_n473_));
  NAi31      u0445(.An(c), .B(f), .C(d), .Y(men_men_n474_));
  AOI210     u0446(.A0(men_men_n262_), .A1(men_men_n180_), .B0(men_men_n474_), .Y(men_men_n475_));
  INV        u0447(.A(men_men_n475_), .Y(men_men_n476_));
  NA3        u0448(.A(men_men_n357_), .B(men_men_n88_), .C(men_men_n87_), .Y(men_men_n477_));
  NA2        u0449(.A(men_men_n212_), .B(men_men_n99_), .Y(men_men_n478_));
  AOI210     u0450(.A0(men_men_n478_), .A1(men_men_n170_), .B0(men_men_n474_), .Y(men_men_n479_));
  AOI210     u0451(.A0(men_men_n336_), .A1(men_men_n35_), .B0(men_men_n449_), .Y(men_men_n480_));
  NOi31      u0452(.An(men_men_n477_), .B(men_men_n480_), .C(men_men_n479_), .Y(men_men_n481_));
  AO220      u0453(.A0(men_men_n270_), .A1(men_men_n245_), .B0(men_men_n155_), .B1(men_men_n64_), .Y(men_men_n482_));
  NA3        u0454(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n483_));
  NO2        u0455(.A(men_men_n483_), .B(men_men_n411_), .Y(men_men_n484_));
  NO2        u0456(.A(men_men_n484_), .B(men_men_n278_), .Y(men_men_n485_));
  NAi41      u0457(.An(men_men_n482_), .B(men_men_n485_), .C(men_men_n481_), .D(men_men_n476_), .Y(men_men_n486_));
  NO3        u0458(.A(men_men_n486_), .B(men_men_n472_), .C(men_men_n469_), .Y(men_men_n487_));
  NA4        u0459(.A(men_men_n487_), .B(men_men_n461_), .C(men_men_n435_), .D(men_men_n406_), .Y(men11));
  NO2        u0460(.A(men_men_n68_), .B(f), .Y(men_men_n489_));
  NA2        u0461(.A(j), .B(u), .Y(men_men_n490_));
  NAi31      u0462(.An(i), .B(m), .C(l), .Y(men_men_n491_));
  NA3        u0463(.A(m), .B(k), .C(j), .Y(men_men_n492_));
  NOi32      u0464(.An(e), .Bn(b), .C(f), .Y(men_men_n493_));
  NA2        u0465(.A(men_men_n242_), .B(men_men_n104_), .Y(men_men_n494_));
  NA2        u0466(.A(men_men_n46_), .B(j), .Y(men_men_n495_));
  NO2        u0467(.A(men_men_n495_), .B(men_men_n284_), .Y(men_men_n496_));
  NAi31      u0468(.An(d), .B(e), .C(a), .Y(men_men_n497_));
  NO2        u0469(.A(men_men_n497_), .B(n), .Y(men_men_n498_));
  AOI220     u0470(.A0(men_men_n498_), .A1(men_men_n92_), .B0(men_men_n496_), .B1(men_men_n493_), .Y(men_men_n499_));
  NAi41      u0471(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n500_));
  AN2        u0472(.A(men_men_n500_), .B(men_men_n347_), .Y(men_men_n501_));
  AOI210     u0473(.A0(men_men_n501_), .A1(men_men_n370_), .B0(men_men_n254_), .Y(men_men_n502_));
  NA2        u0474(.A(j), .B(i), .Y(men_men_n503_));
  NAi31      u0475(.An(n), .B(m), .C(k), .Y(men_men_n504_));
  NO3        u0476(.A(men_men_n504_), .B(men_men_n503_), .C(men_men_n103_), .Y(men_men_n505_));
  NO4        u0477(.A(n), .B(d), .C(men_men_n107_), .D(a), .Y(men_men_n506_));
  OR2        u0478(.A(n), .B(c), .Y(men_men_n507_));
  NO2        u0479(.A(men_men_n507_), .B(men_men_n138_), .Y(men_men_n508_));
  NO2        u0480(.A(men_men_n508_), .B(men_men_n506_), .Y(men_men_n509_));
  NOi32      u0481(.An(u), .Bn(f), .C(i), .Y(men_men_n510_));
  NA2        u0482(.A(men_men_n510_), .B(men_men_n90_), .Y(men_men_n511_));
  NO2        u0483(.A(men_men_n511_), .B(men_men_n509_), .Y(men_men_n512_));
  AOI210     u0484(.A0(men_men_n505_), .A1(men_men_n502_), .B0(men_men_n512_), .Y(men_men_n513_));
  NA2        u0485(.A(men_men_n129_), .B(men_men_n34_), .Y(men_men_n514_));
  OAI220     u0486(.A0(men_men_n514_), .A1(m), .B0(men_men_n495_), .B1(men_men_n218_), .Y(men_men_n515_));
  NOi41      u0487(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n516_));
  NAi32      u0488(.An(e), .Bn(b), .C(c), .Y(men_men_n517_));
  AN2        u0489(.A(men_men_n315_), .B(men_men_n300_), .Y(men_men_n518_));
  NA2        u0490(.A(men_men_n518_), .B(men_men_n517_), .Y(men_men_n519_));
  AN2        u0491(.A(men_men_n519_), .B(men_men_n515_), .Y(men_men_n520_));
  OAI220     u0492(.A0(men_men_n372_), .A1(men_men_n371_), .B0(men_men_n491_), .B1(men_men_n490_), .Y(men_men_n521_));
  NAi31      u0493(.An(d), .B(c), .C(a), .Y(men_men_n522_));
  NO2        u0494(.A(men_men_n522_), .B(n), .Y(men_men_n523_));
  NA3        u0495(.A(men_men_n523_), .B(men_men_n521_), .C(e), .Y(men_men_n524_));
  NO3        u0496(.A(men_men_n59_), .B(men_men_n49_), .C(men_men_n199_), .Y(men_men_n525_));
  NO2        u0497(.A(men_men_n215_), .B(men_men_n101_), .Y(men_men_n526_));
  OAI210     u0498(.A0(men_men_n525_), .A1(men_men_n373_), .B0(men_men_n526_), .Y(men_men_n527_));
  NA2        u0499(.A(men_men_n527_), .B(men_men_n524_), .Y(men_men_n528_));
  NO2        u0500(.A(men_men_n258_), .B(n), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n403_), .B(men_men_n529_), .Y(men_men_n530_));
  NA2        u0502(.A(men_men_n521_), .B(f), .Y(men_men_n531_));
  NAi32      u0503(.An(d), .Bn(a), .C(b), .Y(men_men_n532_));
  NO2        u0504(.A(men_men_n532_), .B(men_men_n49_), .Y(men_men_n533_));
  NA2        u0505(.A(h), .B(f), .Y(men_men_n534_));
  NO2        u0506(.A(men_men_n534_), .B(men_men_n85_), .Y(men_men_n535_));
  NA2        u0507(.A(men_men_n535_), .B(men_men_n533_), .Y(men_men_n536_));
  OAI210     u0508(.A0(men_men_n531_), .A1(men_men_n530_), .B0(men_men_n536_), .Y(men_men_n537_));
  AN3        u0509(.A(j), .B(h), .C(u), .Y(men_men_n538_));
  NO2        u0510(.A(men_men_n135_), .B(c), .Y(men_men_n539_));
  NA3        u0511(.A(f), .B(d), .C(b), .Y(men_men_n540_));
  NO4        u0512(.A(men_men_n540_), .B(men_men_n166_), .C(men_men_n163_), .D(u), .Y(men_men_n541_));
  NO4        u0513(.A(men_men_n541_), .B(men_men_n537_), .C(men_men_n528_), .D(men_men_n520_), .Y(men_men_n542_));
  AN3        u0514(.A(men_men_n542_), .B(men_men_n513_), .C(men_men_n499_), .Y(men_men_n543_));
  INV        u0515(.A(k), .Y(men_men_n544_));
  NA3        u0516(.A(l), .B(men_men_n544_), .C(i), .Y(men_men_n545_));
  INV        u0517(.A(men_men_n545_), .Y(men_men_n546_));
  NA4        u0518(.A(men_men_n369_), .B(men_men_n392_), .C(men_men_n171_), .D(men_men_n104_), .Y(men_men_n547_));
  NAi32      u0519(.An(h), .Bn(f), .C(u), .Y(men_men_n548_));
  NAi41      u0520(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n549_));
  OAI210     u0521(.A0(men_men_n497_), .A1(n), .B0(men_men_n549_), .Y(men_men_n550_));
  NA2        u0522(.A(men_men_n550_), .B(m), .Y(men_men_n551_));
  NAi31      u0523(.An(h), .B(u), .C(f), .Y(men_men_n552_));
  OR3        u0524(.A(men_men_n552_), .B(men_men_n258_), .C(men_men_n49_), .Y(men_men_n553_));
  NA4        u0525(.A(men_men_n392_), .B(men_men_n112_), .C(men_men_n104_), .D(e), .Y(men_men_n554_));
  AN2        u0526(.A(men_men_n554_), .B(men_men_n553_), .Y(men_men_n555_));
  OA210      u0527(.A0(men_men_n551_), .A1(men_men_n548_), .B0(men_men_n555_), .Y(men_men_n556_));
  NO3        u0528(.A(men_men_n548_), .B(men_men_n68_), .C(men_men_n69_), .Y(men_men_n557_));
  NO4        u0529(.A(men_men_n552_), .B(men_men_n507_), .C(men_men_n138_), .D(men_men_n69_), .Y(men_men_n558_));
  OR2        u0530(.A(men_men_n558_), .B(men_men_n557_), .Y(men_men_n559_));
  NAi31      u0531(.An(men_men_n559_), .B(men_men_n556_), .C(men_men_n547_), .Y(men_men_n560_));
  NAi31      u0532(.An(f), .B(h), .C(u), .Y(men_men_n561_));
  NO3        u0533(.A(men_men_n292_), .B(men_men_n561_), .C(men_men_n68_), .Y(men_men_n562_));
  NOi32      u0534(.An(b), .Bn(a), .C(c), .Y(men_men_n563_));
  NOi41      u0535(.An(men_men_n563_), .B(men_men_n329_), .C(men_men_n66_), .D(men_men_n108_), .Y(men_men_n564_));
  OR2        u0536(.A(men_men_n564_), .B(men_men_n562_), .Y(men_men_n565_));
  NOi32      u0537(.An(d), .Bn(a), .C(e), .Y(men_men_n566_));
  NA2        u0538(.A(men_men_n566_), .B(men_men_n104_), .Y(men_men_n567_));
  NO2        u0539(.A(n), .B(c), .Y(men_men_n568_));
  NA3        u0540(.A(men_men_n568_), .B(men_men_n29_), .C(m), .Y(men_men_n569_));
  NAi32      u0541(.An(n), .Bn(f), .C(m), .Y(men_men_n570_));
  NA3        u0542(.A(men_men_n570_), .B(men_men_n569_), .C(men_men_n567_), .Y(men_men_n571_));
  AOI210     u0543(.A0(men_men_n29_), .A1(d), .B0(e), .Y(men_men_n572_));
  AOI210     u0544(.A0(men_men_n572_), .A1(men_men_n198_), .B0(men_men_n514_), .Y(men_men_n573_));
  AOI210     u0545(.A0(men_men_n573_), .A1(men_men_n571_), .B0(men_men_n565_), .Y(men_men_n574_));
  INV        u0546(.A(men_men_n574_), .Y(men_men_n575_));
  AOI210     u0547(.A0(men_men_n560_), .A1(men_men_n546_), .B0(men_men_n575_), .Y(men_men_n576_));
  NO3        u0548(.A(men_men_n298_), .B(men_men_n58_), .C(n), .Y(men_men_n577_));
  NA3        u0549(.A(men_men_n474_), .B(men_men_n161_), .C(men_men_n160_), .Y(men_men_n578_));
  NA2        u0550(.A(men_men_n432_), .B(men_men_n215_), .Y(men_men_n579_));
  OR2        u0551(.A(men_men_n579_), .B(men_men_n578_), .Y(men_men_n580_));
  NA2        u0552(.A(men_men_n70_), .B(men_men_n104_), .Y(men_men_n581_));
  NO2        u0553(.A(men_men_n581_), .B(men_men_n45_), .Y(men_men_n582_));
  AOI220     u0554(.A0(men_men_n582_), .A1(men_men_n502_), .B0(men_men_n580_), .B1(men_men_n577_), .Y(men_men_n583_));
  NO2        u0555(.A(men_men_n583_), .B(men_men_n77_), .Y(men_men_n584_));
  NA3        u0556(.A(men_men_n516_), .B(men_men_n316_), .C(men_men_n46_), .Y(men_men_n585_));
  NOi32      u0557(.An(e), .Bn(c), .C(f), .Y(men_men_n586_));
  NOi21      u0558(.An(f), .B(u), .Y(men_men_n587_));
  NO2        u0559(.A(men_men_n587_), .B(men_men_n196_), .Y(men_men_n588_));
  AOI220     u0560(.A0(men_men_n588_), .A1(men_men_n366_), .B0(men_men_n586_), .B1(men_men_n165_), .Y(men_men_n589_));
  NA3        u0561(.A(men_men_n589_), .B(men_men_n585_), .C(men_men_n168_), .Y(men_men_n590_));
  AOI210     u0562(.A0(men_men_n501_), .A1(men_men_n370_), .B0(men_men_n283_), .Y(men_men_n591_));
  NA2        u0563(.A(men_men_n591_), .B(men_men_n246_), .Y(men_men_n592_));
  NOi21      u0564(.An(j), .B(l), .Y(men_men_n593_));
  NAi21      u0565(.An(k), .B(h), .Y(men_men_n594_));
  NO2        u0566(.A(men_men_n594_), .B(men_men_n244_), .Y(men_men_n595_));
  NA2        u0567(.A(men_men_n595_), .B(men_men_n593_), .Y(men_men_n596_));
  OR2        u0568(.A(men_men_n596_), .B(men_men_n551_), .Y(men_men_n597_));
  NOi31      u0569(.An(m), .B(n), .C(k), .Y(men_men_n598_));
  NA2        u0570(.A(men_men_n593_), .B(men_men_n598_), .Y(men_men_n599_));
  AOI210     u0571(.A0(men_men_n370_), .A1(men_men_n347_), .B0(men_men_n283_), .Y(men_men_n600_));
  NAi21      u0572(.An(men_men_n599_), .B(men_men_n600_), .Y(men_men_n601_));
  NO2        u0573(.A(men_men_n258_), .B(men_men_n49_), .Y(men_men_n602_));
  NO2        u0574(.A(men_men_n292_), .B(men_men_n561_), .Y(men_men_n603_));
  NO2        u0575(.A(men_men_n497_), .B(men_men_n49_), .Y(men_men_n604_));
  AOI220     u0576(.A0(men_men_n604_), .A1(men_men_n603_), .B0(men_men_n602_), .B1(men_men_n535_), .Y(men_men_n605_));
  NA4        u0577(.A(men_men_n605_), .B(men_men_n601_), .C(men_men_n597_), .D(men_men_n592_), .Y(men_men_n606_));
  NA2        u0578(.A(men_men_n99_), .B(men_men_n36_), .Y(men_men_n607_));
  NO2        u0579(.A(k), .B(men_men_n199_), .Y(men_men_n608_));
  NO2        u0580(.A(men_men_n493_), .B(men_men_n338_), .Y(men_men_n609_));
  NO2        u0581(.A(men_men_n609_), .B(n), .Y(men_men_n610_));
  NAi31      u0582(.An(men_men_n607_), .B(men_men_n610_), .C(men_men_n608_), .Y(men_men_n611_));
  NO2        u0583(.A(men_men_n495_), .B(men_men_n166_), .Y(men_men_n612_));
  NA2        u0584(.A(men_men_n473_), .B(men_men_n149_), .Y(men_men_n613_));
  NO3        u0585(.A(men_men_n367_), .B(men_men_n613_), .C(men_men_n77_), .Y(men_men_n614_));
  AOI210     u0586(.A0(c), .A1(men_men_n612_), .B0(men_men_n614_), .Y(men_men_n615_));
  AN3        u0587(.A(f), .B(d), .C(b), .Y(men_men_n616_));
  NAi31      u0588(.An(m), .B(n), .C(k), .Y(men_men_n617_));
  OAI210     u0589(.A0(men_men_n123_), .A1(men_men_n617_), .B0(men_men_n234_), .Y(men_men_n618_));
  NA2        u0590(.A(men_men_n618_), .B(j), .Y(men_men_n619_));
  NA3        u0591(.A(men_men_n619_), .B(men_men_n615_), .C(men_men_n611_), .Y(men_men_n620_));
  NO4        u0592(.A(men_men_n620_), .B(men_men_n606_), .C(men_men_n590_), .D(men_men_n584_), .Y(men_men_n621_));
  NA2        u0593(.A(men_men_n357_), .B(men_men_n152_), .Y(men_men_n622_));
  NAi31      u0594(.An(u), .B(h), .C(f), .Y(men_men_n623_));
  OR3        u0595(.A(men_men_n623_), .B(men_men_n258_), .C(n), .Y(men_men_n624_));
  OA210      u0596(.A0(men_men_n497_), .A1(n), .B0(men_men_n549_), .Y(men_men_n625_));
  NA3        u0597(.A(men_men_n390_), .B(men_men_n112_), .C(men_men_n74_), .Y(men_men_n626_));
  OAI210     u0598(.A0(men_men_n625_), .A1(men_men_n81_), .B0(men_men_n626_), .Y(men_men_n627_));
  NOi21      u0599(.An(men_men_n624_), .B(men_men_n627_), .Y(men_men_n628_));
  AOI210     u0600(.A0(men_men_n628_), .A1(men_men_n622_), .B0(men_men_n492_), .Y(men_men_n629_));
  NO3        u0601(.A(u), .B(men_men_n198_), .C(men_men_n54_), .Y(men_men_n630_));
  NO2        u0602(.A(men_men_n478_), .B(men_men_n77_), .Y(men_men_n631_));
  OAI210     u0603(.A0(men_men_n631_), .A1(men_men_n366_), .B0(men_men_n630_), .Y(men_men_n632_));
  NA2        u0604(.A(men_men_n563_), .B(men_men_n318_), .Y(men_men_n633_));
  OA220      u0605(.A0(men_men_n599_), .A1(men_men_n633_), .B0(men_men_n596_), .B1(men_men_n68_), .Y(men_men_n634_));
  NA3        u0606(.A(men_men_n489_), .B(men_men_n90_), .C(men_men_n89_), .Y(men_men_n635_));
  NA2        u0607(.A(h), .B(men_men_n37_), .Y(men_men_n636_));
  NA2        u0608(.A(men_men_n90_), .B(men_men_n46_), .Y(men_men_n637_));
  OAI220     u0609(.A0(men_men_n637_), .A1(men_men_n308_), .B0(men_men_n636_), .B1(men_men_n437_), .Y(men_men_n638_));
  AOI210     u0610(.A0(men_men_n532_), .A1(men_men_n402_), .B0(men_men_n49_), .Y(men_men_n639_));
  INV        u0611(.A(men_men_n638_), .Y(men_men_n640_));
  NA4        u0612(.A(men_men_n640_), .B(men_men_n635_), .C(men_men_n634_), .D(men_men_n632_), .Y(men_men_n641_));
  OR2        u0613(.A(men_men_n336_), .B(men_men_n102_), .Y(men_men_n642_));
  INV        u0614(.A(men_men_n642_), .Y(men_men_n643_));
  NO3        u0615(.A(men_men_n377_), .B(men_men_n177_), .C(men_men_n176_), .Y(men_men_n644_));
  NA2        u0616(.A(men_men_n644_), .B(men_men_n215_), .Y(men_men_n645_));
  NA3        u0617(.A(men_men_n645_), .B(men_men_n238_), .C(j), .Y(men_men_n646_));
  NO3        u0618(.A(men_men_n432_), .B(men_men_n163_), .C(i), .Y(men_men_n647_));
  NA2        u0619(.A(men_men_n436_), .B(men_men_n74_), .Y(men_men_n648_));
  NA3        u0620(.A(men_men_n646_), .B(men_men_n477_), .C(men_men_n375_), .Y(men_men_n649_));
  NO4        u0621(.A(men_men_n649_), .B(men_men_n643_), .C(men_men_n641_), .D(men_men_n629_), .Y(men_men_n650_));
  NA4        u0622(.A(men_men_n650_), .B(men_men_n621_), .C(men_men_n576_), .D(men_men_n543_), .Y(men08));
  NO2        u0623(.A(k), .B(h), .Y(men_men_n652_));
  AO210      u0624(.A0(men_men_n236_), .A1(men_men_n424_), .B0(men_men_n652_), .Y(men_men_n653_));
  NO2        u0625(.A(men_men_n653_), .B(men_men_n281_), .Y(men_men_n654_));
  NA2        u0626(.A(men_men_n586_), .B(men_men_n74_), .Y(men_men_n655_));
  NA2        u0627(.A(men_men_n655_), .B(men_men_n432_), .Y(men_men_n656_));
  AOI210     u0628(.A0(men_men_n656_), .A1(men_men_n654_), .B0(men_men_n458_), .Y(men_men_n657_));
  NA2        u0629(.A(men_men_n74_), .B(men_men_n101_), .Y(men_men_n658_));
  NO2        u0630(.A(men_men_n658_), .B(men_men_n55_), .Y(men_men_n659_));
  NO4        u0631(.A(men_men_n354_), .B(men_men_n103_), .C(j), .D(men_men_n199_), .Y(men_men_n660_));
  NA2        u0632(.A(men_men_n540_), .B(men_men_n217_), .Y(men_men_n661_));
  AOI220     u0633(.A0(men_men_n661_), .A1(men_men_n323_), .B0(men_men_n660_), .B1(men_men_n659_), .Y(men_men_n662_));
  AOI210     u0634(.A0(men_men_n540_), .A1(men_men_n145_), .B0(men_men_n74_), .Y(men_men_n663_));
  NA4        u0635(.A(men_men_n201_), .B(men_men_n129_), .C(men_men_n45_), .D(h), .Y(men_men_n664_));
  AN2        u0636(.A(l), .B(k), .Y(men_men_n665_));
  NA4        u0637(.A(men_men_n665_), .B(men_men_n99_), .C(men_men_n69_), .D(men_men_n199_), .Y(men_men_n666_));
  NA3        u0638(.A(men_men_n662_), .B(men_men_n657_), .C(men_men_n325_), .Y(men_men_n667_));
  AN2        u0639(.A(men_men_n498_), .B(men_men_n86_), .Y(men_men_n668_));
  NO4        u0640(.A(men_men_n163_), .B(men_men_n365_), .C(men_men_n103_), .D(u), .Y(men_men_n669_));
  AOI210     u0641(.A0(men_men_n669_), .A1(men_men_n661_), .B0(men_men_n484_), .Y(men_men_n670_));
  NO2        u0642(.A(men_men_n38_), .B(men_men_n198_), .Y(men_men_n671_));
  AOI220     u0643(.A0(men_men_n588_), .A1(men_men_n322_), .B0(men_men_n671_), .B1(men_men_n529_), .Y(men_men_n672_));
  NAi31      u0644(.An(men_men_n668_), .B(men_men_n672_), .C(men_men_n670_), .Y(men_men_n673_));
  NO2        u0645(.A(men_men_n501_), .B(men_men_n35_), .Y(men_men_n674_));
  OAI210     u0646(.A0(men_men_n517_), .A1(men_men_n47_), .B0(men_men_n123_), .Y(men_men_n675_));
  NO2        u0647(.A(men_men_n453_), .B(men_men_n122_), .Y(men_men_n676_));
  AOI210     u0648(.A0(men_men_n676_), .A1(men_men_n675_), .B0(men_men_n674_), .Y(men_men_n677_));
  NO3        u0649(.A(men_men_n298_), .B(men_men_n121_), .C(men_men_n41_), .Y(men_men_n678_));
  NAi21      u0650(.An(men_men_n678_), .B(men_men_n666_), .Y(men_men_n679_));
  NA2        u0651(.A(men_men_n653_), .B(men_men_n124_), .Y(men_men_n680_));
  AOI220     u0652(.A0(men_men_n680_), .A1(men_men_n376_), .B0(men_men_n679_), .B1(e), .Y(men_men_n681_));
  OAI210     u0653(.A0(men_men_n677_), .A1(men_men_n77_), .B0(men_men_n681_), .Y(men_men_n682_));
  NA2        u0654(.A(men_men_n338_), .B(men_men_n43_), .Y(men_men_n683_));
  NA3        u0655(.A(men_men_n645_), .B(men_men_n310_), .C(men_men_n360_), .Y(men_men_n684_));
  NA2        u0656(.A(men_men_n665_), .B(men_men_n206_), .Y(men_men_n685_));
  NO2        u0657(.A(men_men_n685_), .B(men_men_n306_), .Y(men_men_n686_));
  AOI210     u0658(.A0(men_men_n686_), .A1(i), .B0(men_men_n457_), .Y(men_men_n687_));
  NA3        u0659(.A(m), .B(l), .C(k), .Y(men_men_n688_));
  AOI210     u0660(.A0(men_men_n626_), .A1(men_men_n624_), .B0(men_men_n688_), .Y(men_men_n689_));
  NO2        u0661(.A(men_men_n500_), .B(men_men_n254_), .Y(men_men_n690_));
  NOi21      u0662(.An(men_men_n690_), .B(men_men_n494_), .Y(men_men_n691_));
  NA4        u0663(.A(men_men_n104_), .B(l), .C(k), .D(men_men_n77_), .Y(men_men_n692_));
  NA3        u0664(.A(men_men_n112_), .B(men_men_n385_), .C(i), .Y(men_men_n693_));
  NO2        u0665(.A(men_men_n693_), .B(men_men_n692_), .Y(men_men_n694_));
  NO3        u0666(.A(men_men_n694_), .B(men_men_n691_), .C(men_men_n689_), .Y(men_men_n695_));
  NA4        u0667(.A(men_men_n695_), .B(men_men_n687_), .C(men_men_n684_), .D(men_men_n683_), .Y(men_men_n696_));
  NO4        u0668(.A(men_men_n696_), .B(men_men_n682_), .C(men_men_n673_), .D(men_men_n667_), .Y(men_men_n697_));
  NA2        u0669(.A(men_men_n588_), .B(men_men_n366_), .Y(men_men_n698_));
  NOi31      u0670(.An(u), .B(h), .C(f), .Y(men_men_n699_));
  NA2        u0671(.A(men_men_n604_), .B(men_men_n699_), .Y(men_men_n700_));
  AO210      u0672(.A0(men_men_n700_), .A1(men_men_n553_), .B0(men_men_n503_), .Y(men_men_n701_));
  NO3        u0673(.A(men_men_n370_), .B(men_men_n490_), .C(h), .Y(men_men_n702_));
  AOI210     u0674(.A0(men_men_n702_), .A1(men_men_n104_), .B0(men_men_n467_), .Y(men_men_n703_));
  NA4        u0675(.A(men_men_n703_), .B(men_men_n701_), .C(men_men_n698_), .D(men_men_n235_), .Y(men_men_n704_));
  NA2        u0676(.A(men_men_n665_), .B(men_men_n69_), .Y(men_men_n705_));
  NO3        u0677(.A(men_men_n644_), .B(men_men_n163_), .C(i), .Y(men_men_n706_));
  NOi21      u0678(.An(h), .B(j), .Y(men_men_n707_));
  NA2        u0679(.A(men_men_n707_), .B(f), .Y(men_men_n708_));
  NO2        u0680(.A(men_men_n708_), .B(men_men_n229_), .Y(men_men_n709_));
  NO3        u0681(.A(men_men_n709_), .B(men_men_n706_), .C(men_men_n647_), .Y(men_men_n710_));
  OAI220     u0682(.A0(men_men_n710_), .A1(men_men_n705_), .B0(men_men_n555_), .B1(men_men_n59_), .Y(men_men_n711_));
  AOI210     u0683(.A0(men_men_n704_), .A1(l), .B0(men_men_n711_), .Y(men_men_n712_));
  NO2        u0684(.A(j), .B(i), .Y(men_men_n713_));
  NA3        u0685(.A(men_men_n713_), .B(men_men_n72_), .C(l), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n713_), .B(men_men_n33_), .Y(men_men_n715_));
  NA2        u0687(.A(men_men_n395_), .B(men_men_n112_), .Y(men_men_n716_));
  OA220      u0688(.A0(men_men_n716_), .A1(men_men_n715_), .B0(men_men_n714_), .B1(men_men_n551_), .Y(men_men_n717_));
  NO3        u0689(.A(men_men_n140_), .B(men_men_n49_), .C(men_men_n101_), .Y(men_men_n718_));
  NO3        u0690(.A(men_men_n507_), .B(men_men_n138_), .C(men_men_n69_), .Y(men_men_n719_));
  NO3        u0691(.A(men_men_n453_), .B(men_men_n412_), .C(j), .Y(men_men_n720_));
  OAI210     u0692(.A0(men_men_n719_), .A1(men_men_n718_), .B0(men_men_n720_), .Y(men_men_n721_));
  OAI210     u0693(.A0(men_men_n700_), .A1(men_men_n59_), .B0(men_men_n721_), .Y(men_men_n722_));
  NO2        u0694(.A(men_men_n281_), .B(men_men_n40_), .Y(men_men_n723_));
  AOI210     u0695(.A0(men_men_n493_), .A1(n), .B0(men_men_n516_), .Y(men_men_n724_));
  NA2        u0696(.A(men_men_n724_), .B(men_men_n518_), .Y(men_men_n725_));
  AN3        u0697(.A(men_men_n725_), .B(men_men_n723_), .C(men_men_n89_), .Y(men_men_n726_));
  NO3        u0698(.A(men_men_n163_), .B(men_men_n365_), .C(men_men_n103_), .Y(men_men_n727_));
  AOI220     u0699(.A0(men_men_n727_), .A1(men_men_n230_), .B0(men_men_n579_), .B1(men_men_n290_), .Y(men_men_n728_));
  NAi31      u0700(.An(men_men_n572_), .B(men_men_n83_), .C(men_men_n74_), .Y(men_men_n729_));
  NA2        u0701(.A(men_men_n729_), .B(men_men_n728_), .Y(men_men_n730_));
  NO2        u0702(.A(men_men_n281_), .B(men_men_n124_), .Y(men_men_n731_));
  AOI220     u0703(.A0(men_men_n731_), .A1(men_men_n588_), .B0(men_men_n678_), .B1(men_men_n663_), .Y(men_men_n732_));
  NA2        u0704(.A(men_men_n720_), .B(men_men_n639_), .Y(men_men_n733_));
  NA2        u0705(.A(men_men_n733_), .B(men_men_n732_), .Y(men_men_n734_));
  OR4        u0706(.A(men_men_n734_), .B(men_men_n730_), .C(men_men_n726_), .D(men_men_n722_), .Y(men_men_n735_));
  NA3        u0707(.A(men_men_n724_), .B(men_men_n518_), .C(men_men_n517_), .Y(men_men_n736_));
  NA4        u0708(.A(men_men_n736_), .B(men_men_n201_), .C(men_men_n424_), .D(men_men_n34_), .Y(men_men_n737_));
  NO4        u0709(.A(men_men_n453_), .B(men_men_n407_), .C(j), .D(f), .Y(men_men_n738_));
  OAI220     u0710(.A0(men_men_n664_), .A1(men_men_n655_), .B0(men_men_n308_), .B1(men_men_n38_), .Y(men_men_n739_));
  AOI210     u0711(.A0(men_men_n738_), .A1(men_men_n241_), .B0(men_men_n739_), .Y(men_men_n740_));
  NA3        u0712(.A(men_men_n510_), .B(men_men_n274_), .C(h), .Y(men_men_n741_));
  NOi21      u0713(.An(men_men_n639_), .B(men_men_n741_), .Y(men_men_n742_));
  NO2        u0714(.A(men_men_n82_), .B(men_men_n47_), .Y(men_men_n743_));
  OAI220     u0715(.A0(men_men_n741_), .A1(men_men_n569_), .B0(men_men_n714_), .B1(men_men_n68_), .Y(men_men_n744_));
  AOI210     u0716(.A0(men_men_n743_), .A1(men_men_n610_), .B0(men_men_n744_), .Y(men_men_n745_));
  NAi41      u0717(.An(men_men_n742_), .B(men_men_n745_), .C(men_men_n740_), .D(men_men_n737_), .Y(men_men_n746_));
  AOI220     u0718(.A0(men_men_n86_), .A1(men_men_n223_), .B0(men_men_n720_), .B1(men_men_n602_), .Y(men_men_n747_));
  NO2        u0719(.A(men_men_n625_), .B(men_men_n69_), .Y(men_men_n748_));
  AOI210     u0720(.A0(men_men_n738_), .A1(men_men_n748_), .B0(men_men_n312_), .Y(men_men_n749_));
  INV        u0721(.A(men_men_n483_), .Y(men_men_n750_));
  NA3        u0722(.A(men_men_n233_), .B(men_men_n56_), .C(b), .Y(men_men_n751_));
  AOI220     u0723(.A0(men_men_n568_), .A1(men_men_n29_), .B0(men_men_n436_), .B1(men_men_n74_), .Y(men_men_n752_));
  NA2        u0724(.A(men_men_n752_), .B(men_men_n751_), .Y(men_men_n753_));
  NO2        u0725(.A(men_men_n741_), .B(men_men_n456_), .Y(men_men_n754_));
  AOI210     u0726(.A0(men_men_n753_), .A1(men_men_n750_), .B0(men_men_n754_), .Y(men_men_n755_));
  NA3        u0727(.A(men_men_n755_), .B(men_men_n749_), .C(men_men_n747_), .Y(men_men_n756_));
  NOi41      u0728(.An(men_men_n717_), .B(men_men_n756_), .C(men_men_n746_), .D(men_men_n735_), .Y(men_men_n757_));
  OR2        u0729(.A(men_men_n664_), .B(men_men_n217_), .Y(men_men_n758_));
  NO3        u0730(.A(men_men_n317_), .B(men_men_n283_), .C(men_men_n103_), .Y(men_men_n759_));
  NA2        u0731(.A(men_men_n46_), .B(men_men_n54_), .Y(men_men_n760_));
  NO3        u0732(.A(men_men_n760_), .B(men_men_n715_), .C(men_men_n258_), .Y(men_men_n761_));
  NO3        u0733(.A(men_men_n490_), .B(men_men_n84_), .C(h), .Y(men_men_n762_));
  AOI210     u0734(.A0(men_men_n762_), .A1(men_men_n659_), .B0(men_men_n761_), .Y(men_men_n763_));
  NA3        u0735(.A(men_men_n763_), .B(men_men_n758_), .C(men_men_n378_), .Y(men_men_n764_));
  OR2        u0736(.A(men_men_n623_), .B(men_men_n82_), .Y(men_men_n765_));
  NOi31      u0737(.An(b), .B(d), .C(a), .Y(men_men_n766_));
  NO2        u0738(.A(men_men_n766_), .B(men_men_n566_), .Y(men_men_n767_));
  NO2        u0739(.A(men_men_n767_), .B(n), .Y(men_men_n768_));
  NOi21      u0740(.An(men_men_n752_), .B(men_men_n768_), .Y(men_men_n769_));
  OAI220     u0741(.A0(men_men_n769_), .A1(men_men_n765_), .B0(men_men_n741_), .B1(men_men_n567_), .Y(men_men_n770_));
  INV        u0742(.A(men_men_n517_), .Y(men_men_n771_));
  NO3        u0743(.A(men_men_n587_), .B(men_men_n306_), .C(men_men_n108_), .Y(men_men_n772_));
  NOi21      u0744(.An(men_men_n772_), .B(men_men_n150_), .Y(men_men_n773_));
  AOI210     u0745(.A0(men_men_n759_), .A1(men_men_n771_), .B0(men_men_n773_), .Y(men_men_n774_));
  INV        u0746(.A(men_men_n774_), .Y(men_men_n775_));
  NO2        u0747(.A(men_men_n644_), .B(n), .Y(men_men_n776_));
  NA2        u0748(.A(men_men_n776_), .B(men_men_n654_), .Y(men_men_n777_));
  NO2        u0749(.A(men_men_n304_), .B(men_men_n222_), .Y(men_men_n778_));
  OAI210     u0750(.A0(men_men_n86_), .A1(men_men_n83_), .B0(men_men_n778_), .Y(men_men_n779_));
  NA2        u0751(.A(men_men_n112_), .B(men_men_n74_), .Y(men_men_n780_));
  AOI210     u0752(.A0(men_men_n399_), .A1(men_men_n391_), .B0(men_men_n780_), .Y(men_men_n781_));
  NAi21      u0753(.An(men_men_n781_), .B(men_men_n779_), .Y(men_men_n782_));
  NA2        u0754(.A(men_men_n686_), .B(men_men_n34_), .Y(men_men_n783_));
  NAi21      u0755(.An(men_men_n692_), .B(men_men_n408_), .Y(men_men_n784_));
  NA2        u0756(.A(men_men_n669_), .B(men_men_n324_), .Y(men_men_n785_));
  OAI210     u0757(.A0(men_men_n558_), .A1(men_men_n557_), .B0(men_men_n339_), .Y(men_men_n786_));
  AN3        u0758(.A(men_men_n786_), .B(men_men_n785_), .C(men_men_n784_), .Y(men_men_n787_));
  NAi41      u0759(.An(men_men_n782_), .B(men_men_n787_), .C(men_men_n783_), .D(men_men_n777_), .Y(men_men_n788_));
  NO4        u0760(.A(men_men_n788_), .B(men_men_n775_), .C(men_men_n770_), .D(men_men_n764_), .Y(men_men_n789_));
  NA4        u0761(.A(men_men_n789_), .B(men_men_n757_), .C(men_men_n712_), .D(men_men_n697_), .Y(men09));
  INV        u0762(.A(men_men_n113_), .Y(men_men_n791_));
  NA2        u0763(.A(f), .B(e), .Y(men_men_n792_));
  NO2        u0764(.A(men_men_n211_), .B(men_men_n103_), .Y(men_men_n793_));
  NO2        u0765(.A(u), .B(men_men_n440_), .Y(men_men_n794_));
  NO2        u0766(.A(men_men_n794_), .B(men_men_n792_), .Y(men_men_n795_));
  NA2        u0767(.A(men_men_n418_), .B(e), .Y(men_men_n796_));
  NO2        u0768(.A(men_men_n796_), .B(men_men_n474_), .Y(men_men_n797_));
  AOI210     u0769(.A0(men_men_n795_), .A1(men_men_n791_), .B0(men_men_n797_), .Y(men_men_n798_));
  NO2        u0770(.A(men_men_n189_), .B(men_men_n198_), .Y(men_men_n799_));
  NA3        u0771(.A(m), .B(l), .C(i), .Y(men_men_n800_));
  OAI220     u0772(.A0(men_men_n552_), .A1(men_men_n800_), .B0(men_men_n329_), .B1(men_men_n491_), .Y(men_men_n801_));
  NA4        u0773(.A(men_men_n78_), .B(men_men_n77_), .C(u), .D(f), .Y(men_men_n802_));
  NAi31      u0774(.An(men_men_n801_), .B(men_men_n802_), .C(men_men_n413_), .Y(men_men_n803_));
  OR2        u0775(.A(men_men_n803_), .B(men_men_n799_), .Y(men_men_n804_));
  NA3        u0776(.A(men_men_n765_), .B(men_men_n531_), .C(men_men_n483_), .Y(men_men_n805_));
  OA210      u0777(.A0(men_men_n805_), .A1(men_men_n804_), .B0(men_men_n768_), .Y(men_men_n806_));
  INV        u0778(.A(men_men_n315_), .Y(men_men_n807_));
  NO2        u0779(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n808_));
  NOi31      u0780(.An(k), .B(m), .C(l), .Y(men_men_n809_));
  NO2        u0781(.A(men_men_n316_), .B(men_men_n809_), .Y(men_men_n810_));
  AOI210     u0782(.A0(men_men_n810_), .A1(men_men_n808_), .B0(men_men_n561_), .Y(men_men_n811_));
  NA2        u0783(.A(men_men_n751_), .B(men_men_n308_), .Y(men_men_n812_));
  NA2        u0784(.A(men_men_n318_), .B(men_men_n319_), .Y(men_men_n813_));
  OAI210     u0785(.A0(men_men_n189_), .A1(men_men_n198_), .B0(men_men_n813_), .Y(men_men_n814_));
  AOI220     u0786(.A0(men_men_n814_), .A1(men_men_n812_), .B0(men_men_n811_), .B1(men_men_n807_), .Y(men_men_n815_));
  NA3        u0787(.A(men_men_n105_), .B(men_men_n175_), .C(men_men_n31_), .Y(men_men_n816_));
  NA3        u0788(.A(men_men_n816_), .B(men_men_n815_), .C(men_men_n589_), .Y(men_men_n817_));
  NO2        u0789(.A(men_men_n548_), .B(men_men_n463_), .Y(men_men_n818_));
  NA2        u0790(.A(men_men_n818_), .B(men_men_n175_), .Y(men_men_n819_));
  NOi21      u0791(.An(f), .B(d), .Y(men_men_n820_));
  NA2        u0792(.A(men_men_n820_), .B(m), .Y(men_men_n821_));
  NOi32      u0793(.An(u), .Bn(f), .C(d), .Y(men_men_n822_));
  NA4        u0794(.A(men_men_n822_), .B(men_men_n568_), .C(men_men_n29_), .D(m), .Y(men_men_n823_));
  NOi21      u0795(.An(men_men_n293_), .B(men_men_n823_), .Y(men_men_n824_));
  INV        u0796(.A(men_men_n824_), .Y(men_men_n825_));
  AN2        u0797(.A(f), .B(d), .Y(men_men_n826_));
  NA3        u0798(.A(men_men_n447_), .B(men_men_n826_), .C(men_men_n74_), .Y(men_men_n827_));
  NO3        u0799(.A(men_men_n827_), .B(men_men_n69_), .C(men_men_n199_), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n267_), .B(men_men_n54_), .Y(men_men_n829_));
  INV        u0801(.A(men_men_n828_), .Y(men_men_n830_));
  NAi41      u0802(.An(men_men_n455_), .B(men_men_n830_), .C(men_men_n825_), .D(men_men_n819_), .Y(men_men_n831_));
  NO3        u0803(.A(men_men_n122_), .B(men_men_n306_), .C(men_men_n141_), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n617_), .B(men_men_n306_), .Y(men_men_n833_));
  NO2        u0805(.A(men_men_n832_), .B(men_men_n219_), .Y(men_men_n834_));
  NA2        u0806(.A(men_men_n566_), .B(men_men_n74_), .Y(men_men_n835_));
  NO2        u0807(.A(men_men_n813_), .B(men_men_n835_), .Y(men_men_n836_));
  NA3        u0808(.A(men_men_n149_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n837_));
  OAI220     u0809(.A0(men_men_n827_), .A1(men_men_n404_), .B0(men_men_n315_), .B1(men_men_n837_), .Y(men_men_n838_));
  NOi31      u0810(.An(men_men_n209_), .B(men_men_n838_), .C(men_men_n836_), .Y(men_men_n839_));
  NA3        u0811(.A(e), .B(men_men_n282_), .C(f), .Y(men_men_n840_));
  OR2        u0812(.A(men_men_n623_), .B(men_men_n504_), .Y(men_men_n841_));
  INV        u0813(.A(men_men_n841_), .Y(men_men_n842_));
  NA2        u0814(.A(men_men_n767_), .B(men_men_n102_), .Y(men_men_n843_));
  NA2        u0815(.A(men_men_n843_), .B(men_men_n842_), .Y(men_men_n844_));
  NA4        u0816(.A(men_men_n844_), .B(men_men_n840_), .C(men_men_n839_), .D(men_men_n834_), .Y(men_men_n845_));
  NO4        u0817(.A(men_men_n845_), .B(men_men_n831_), .C(men_men_n817_), .D(men_men_n806_), .Y(men_men_n846_));
  BUFFER     u0818(.A(men_men_n827_), .Y(men_men_n847_));
  NO2        u0819(.A(men_men_n275_), .B(men_men_n847_), .Y(men_men_n848_));
  NO2        u0820(.A(men_men_n308_), .B(men_men_n802_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n124_), .B(men_men_n122_), .Y(men_men_n850_));
  NO2        u0822(.A(men_men_n215_), .B(men_men_n210_), .Y(men_men_n851_));
  AOI220     u0823(.A0(men_men_n851_), .A1(men_men_n212_), .B0(men_men_n288_), .B1(men_men_n850_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n404_), .B(men_men_n792_), .Y(men_men_n853_));
  NA2        u0825(.A(men_men_n853_), .B(men_men_n523_), .Y(men_men_n854_));
  NA2        u0826(.A(men_men_n854_), .B(men_men_n852_), .Y(men_men_n855_));
  NA2        u0827(.A(e), .B(d), .Y(men_men_n856_));
  OAI220     u0828(.A0(men_men_n856_), .A1(c), .B0(men_men_n304_), .B1(d), .Y(men_men_n857_));
  NA3        u0829(.A(men_men_n857_), .B(men_men_n426_), .C(men_men_n473_), .Y(men_men_n858_));
  AOI210     u0830(.A0(men_men_n478_), .A1(men_men_n170_), .B0(men_men_n215_), .Y(men_men_n859_));
  AOI210     u0831(.A0(men_men_n588_), .A1(men_men_n322_), .B0(men_men_n859_), .Y(men_men_n860_));
  NA2        u0832(.A(men_men_n267_), .B(men_men_n154_), .Y(men_men_n861_));
  NA2        u0833(.A(men_men_n860_), .B(men_men_n858_), .Y(men_men_n862_));
  NO4        u0834(.A(men_men_n862_), .B(men_men_n855_), .C(men_men_n849_), .D(men_men_n848_), .Y(men_men_n863_));
  NA2        u0835(.A(men_men_n807_), .B(men_men_n31_), .Y(men_men_n864_));
  AO210      u0836(.A0(men_men_n864_), .A1(men_men_n655_), .B0(men_men_n202_), .Y(men_men_n865_));
  AOI220     u0837(.A0(u), .A1(men_men_n833_), .B0(men_men_n577_), .B1(men_men_n586_), .Y(men_men_n866_));
  OAI210     u0838(.A0(men_men_n796_), .A1(men_men_n160_), .B0(men_men_n866_), .Y(men_men_n867_));
  OAI210     u0839(.A0(men_men_n793_), .A1(men_men_n861_), .B0(men_men_n822_), .Y(men_men_n868_));
  NO2        u0840(.A(men_men_n868_), .B(men_men_n569_), .Y(men_men_n869_));
  AOI210     u0841(.A0(men_men_n109_), .A1(men_men_n108_), .B0(men_men_n242_), .Y(men_men_n870_));
  NO2        u0842(.A(men_men_n870_), .B(men_men_n823_), .Y(men_men_n871_));
  AO210      u0843(.A0(men_men_n812_), .A1(men_men_n801_), .B0(men_men_n871_), .Y(men_men_n872_));
  NOi31      u0844(.An(men_men_n508_), .B(men_men_n821_), .C(men_men_n275_), .Y(men_men_n873_));
  NO4        u0845(.A(men_men_n873_), .B(men_men_n872_), .C(men_men_n869_), .D(men_men_n867_), .Y(men_men_n874_));
  AO210      u0846(.A0(men_men_n426_), .A1(men_men_n707_), .B0(men_men_n165_), .Y(men_men_n875_));
  OAI210     u0847(.A0(men_men_n875_), .A1(men_men_n428_), .B0(men_men_n857_), .Y(men_men_n876_));
  NO2        u0848(.A(men_men_n412_), .B(men_men_n67_), .Y(men_men_n877_));
  OAI210     u0849(.A0(men_men_n805_), .A1(men_men_n877_), .B0(men_men_n659_), .Y(men_men_n878_));
  AN4        u0850(.A(men_men_n878_), .B(men_men_n876_), .C(men_men_n874_), .D(men_men_n865_), .Y(men_men_n879_));
  NA4        u0851(.A(men_men_n879_), .B(men_men_n863_), .C(men_men_n846_), .D(men_men_n798_), .Y(men12));
  NO4        u0852(.A(men_men_n417_), .B(men_men_n236_), .C(men_men_n544_), .D(men_men_n199_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n508_), .B(men_men_n877_), .Y(men_men_n882_));
  NO2        u0854(.A(men_men_n425_), .B(men_men_n107_), .Y(men_men_n883_));
  NO2        u0855(.A(men_men_n623_), .B(men_men_n354_), .Y(men_men_n884_));
  NA2        u0856(.A(men_men_n882_), .B(men_men_n416_), .Y(men_men_n885_));
  AOI210     u0857(.A0(men_men_n218_), .A1(men_men_n314_), .B0(men_men_n186_), .Y(men_men_n886_));
  OR2        u0858(.A(men_men_n886_), .B(men_men_n881_), .Y(men_men_n887_));
  NA2        u0859(.A(men_men_n887_), .B(men_men_n377_), .Y(men_men_n888_));
  NO2        u0860(.A(men_men_n607_), .B(men_men_n244_), .Y(men_men_n889_));
  NO2        u0861(.A(men_men_n552_), .B(men_men_n800_), .Y(men_men_n890_));
  AOI220     u0862(.A0(men_men_n890_), .A1(men_men_n529_), .B0(men_men_n778_), .B1(men_men_n889_), .Y(men_men_n891_));
  NO2        u0863(.A(men_men_n140_), .B(men_men_n222_), .Y(men_men_n892_));
  NA3        u0864(.A(men_men_n892_), .B(men_men_n225_), .C(i), .Y(men_men_n893_));
  NA3        u0865(.A(men_men_n893_), .B(men_men_n891_), .C(men_men_n888_), .Y(men_men_n894_));
  NO3        u0866(.A(men_men_n122_), .B(men_men_n141_), .C(men_men_n199_), .Y(men_men_n895_));
  NA2        u0867(.A(men_men_n895_), .B(men_men_n493_), .Y(men_men_n896_));
  NA3        u0868(.A(men_men_n418_), .B(men_men_n410_), .C(u), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n897_), .B(men_men_n896_), .Y(men_men_n898_));
  NO3        u0870(.A(men_men_n628_), .B(men_men_n82_), .C(men_men_n45_), .Y(men_men_n899_));
  NO4        u0871(.A(men_men_n899_), .B(men_men_n898_), .C(men_men_n894_), .D(men_men_n885_), .Y(men_men_n900_));
  NO2        u0872(.A(men_men_n344_), .B(men_men_n343_), .Y(men_men_n901_));
  NA2        u0873(.A(men_men_n549_), .B(men_men_n68_), .Y(men_men_n902_));
  INV        u0874(.A(men_men_n517_), .Y(men_men_n903_));
  NOi21      u0875(.An(men_men_n34_), .B(men_men_n617_), .Y(men_men_n904_));
  AOI220     u0876(.A0(men_men_n904_), .A1(men_men_n903_), .B0(men_men_n902_), .B1(men_men_n901_), .Y(men_men_n905_));
  OAI210     u0877(.A0(men_men_n234_), .A1(men_men_n45_), .B0(men_men_n905_), .Y(men_men_n906_));
  NA2        u0878(.A(men_men_n408_), .B(men_men_n246_), .Y(men_men_n907_));
  NO3        u0879(.A(men_men_n780_), .B(men_men_n79_), .C(men_men_n382_), .Y(men_men_n908_));
  NAi31      u0880(.An(men_men_n908_), .B(men_men_n907_), .C(men_men_n302_), .Y(men_men_n909_));
  NO2        u0881(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n910_));
  NO2        u0882(.A(men_men_n470_), .B(men_men_n283_), .Y(men_men_n911_));
  NA2        u0883(.A(men_men_n598_), .B(men_men_n339_), .Y(men_men_n912_));
  OAI210     u0884(.A0(men_men_n693_), .A1(men_men_n912_), .B0(men_men_n341_), .Y(men_men_n913_));
  NO3        u0885(.A(men_men_n913_), .B(men_men_n909_), .C(men_men_n906_), .Y(men_men_n914_));
  NA2        u0886(.A(men_men_n322_), .B(u), .Y(men_men_n915_));
  NA2        u0887(.A(men_men_n152_), .B(i), .Y(men_men_n916_));
  NA2        u0888(.A(men_men_n46_), .B(i), .Y(men_men_n917_));
  OAI220     u0889(.A0(men_men_n917_), .A1(men_men_n185_), .B0(men_men_n916_), .B1(men_men_n82_), .Y(men_men_n918_));
  AOI210     u0890(.A0(men_men_n393_), .A1(men_men_n37_), .B0(men_men_n918_), .Y(men_men_n919_));
  OR2        u0891(.A(e), .B(men_men_n516_), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n517_), .B(men_men_n358_), .Y(men_men_n921_));
  NO2        u0893(.A(men_men_n921_), .B(men_men_n920_), .Y(men_men_n922_));
  OAI220     u0894(.A0(men_men_n922_), .A1(men_men_n915_), .B0(men_men_n919_), .B1(men_men_n308_), .Y(men_men_n923_));
  NO2        u0895(.A(men_men_n623_), .B(men_men_n463_), .Y(men_men_n924_));
  NA3        u0896(.A(men_men_n318_), .B(men_men_n593_), .C(i), .Y(men_men_n925_));
  OAI210     u0897(.A0(men_men_n412_), .A1(men_men_n292_), .B0(men_men_n925_), .Y(men_men_n926_));
  OAI220     u0898(.A0(men_men_n926_), .A1(men_men_n924_), .B0(men_men_n639_), .B1(men_men_n719_), .Y(men_men_n927_));
  NA2        u0899(.A(e), .B(men_men_n104_), .Y(men_men_n928_));
  OR3        u0900(.A(men_men_n292_), .B(men_men_n407_), .C(f), .Y(men_men_n929_));
  NA3        u0901(.A(men_men_n593_), .B(men_men_n72_), .C(i), .Y(men_men_n930_));
  OA220      u0902(.A0(men_men_n930_), .A1(men_men_n928_), .B0(men_men_n929_), .B1(men_men_n551_), .Y(men_men_n931_));
  NA3        u0903(.A(f), .B(men_men_n109_), .C(u), .Y(men_men_n932_));
  AOI210     u0904(.A0(men_men_n636_), .A1(men_men_n932_), .B0(m), .Y(men_men_n933_));
  OAI210     u0905(.A0(men_men_n933_), .A1(men_men_n118_), .B0(men_men_n305_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n648_), .B(men_men_n835_), .Y(men_men_n935_));
  NA2        u0907(.A(men_men_n802_), .B(men_men_n413_), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n207_), .B(h), .Y(men_men_n937_));
  NA3        u0909(.A(men_men_n937_), .B(men_men_n930_), .C(men_men_n929_), .Y(men_men_n938_));
  AOI220     u0910(.A0(men_men_n938_), .A1(men_men_n241_), .B0(men_men_n936_), .B1(men_men_n935_), .Y(men_men_n939_));
  NA4        u0911(.A(men_men_n939_), .B(men_men_n934_), .C(men_men_n931_), .D(men_men_n927_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n889_), .B(men_men_n223_), .Y(men_men_n941_));
  NA2        u0913(.A(men_men_n627_), .B(men_men_n78_), .Y(men_men_n942_));
  NO2        u0914(.A(men_men_n431_), .B(men_men_n199_), .Y(men_men_n943_));
  AOI210     u0915(.A0(men_men_n943_), .A1(men_men_n359_), .B0(men_men_n203_), .Y(men_men_n944_));
  AOI220     u0916(.A0(men_men_n884_), .A1(men_men_n892_), .B0(men_men_n550_), .B1(men_men_n80_), .Y(men_men_n945_));
  NA4        u0917(.A(men_men_n945_), .B(men_men_n944_), .C(men_men_n942_), .D(men_men_n941_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n936_), .B(men_men_n506_), .Y(men_men_n947_));
  AOI210     u0919(.A0(men_men_n394_), .A1(men_men_n386_), .B0(men_men_n780_), .Y(men_men_n948_));
  OAI210     u0920(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n100_), .Y(men_men_n949_));
  AOI210     u0921(.A0(men_men_n949_), .A1(men_men_n498_), .B0(men_men_n948_), .Y(men_men_n950_));
  NA2        u0922(.A(men_men_n933_), .B(men_men_n883_), .Y(men_men_n951_));
  NO3        u0923(.A(l), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n952_), .B(men_men_n591_), .Y(men_men_n953_));
  NA4        u0925(.A(men_men_n953_), .B(men_men_n951_), .C(men_men_n950_), .D(men_men_n947_), .Y(men_men_n954_));
  NO4        u0926(.A(men_men_n954_), .B(men_men_n946_), .C(men_men_n940_), .D(men_men_n923_), .Y(men_men_n955_));
  NAi31      u0927(.An(men_men_n130_), .B(men_men_n395_), .C(n), .Y(men_men_n956_));
  NO3        u0928(.A(men_men_n117_), .B(men_men_n316_), .C(men_men_n809_), .Y(men_men_n957_));
  NO2        u0929(.A(men_men_n957_), .B(men_men_n956_), .Y(men_men_n958_));
  NO2        u0930(.A(men_men_n254_), .B(men_men_n130_), .Y(men_men_n959_));
  AOI210     u0931(.A0(men_men_n959_), .A1(men_men_n464_), .B0(men_men_n958_), .Y(men_men_n960_));
  NA2        u0932(.A(men_men_n458_), .B(i), .Y(men_men_n961_));
  NA2        u0933(.A(men_men_n961_), .B(men_men_n960_), .Y(men_men_n962_));
  NA2        u0934(.A(men_men_n215_), .B(men_men_n161_), .Y(men_men_n963_));
  NO3        u0935(.A(men_men_n290_), .B(men_men_n418_), .C(men_men_n165_), .Y(men_men_n964_));
  NOi31      u0936(.An(men_men_n963_), .B(men_men_n964_), .C(men_men_n199_), .Y(men_men_n965_));
  NAi21      u0937(.An(men_men_n517_), .B(men_men_n943_), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n411_), .B(men_men_n835_), .Y(men_men_n967_));
  NO2        u0939(.A(men_men_n412_), .B(men_men_n292_), .Y(men_men_n968_));
  NA2        u0940(.A(men_men_n968_), .B(men_men_n967_), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n969_), .B(men_men_n966_), .Y(men_men_n970_));
  OAI220     u0942(.A0(men_men_n956_), .A1(men_men_n218_), .B0(men_men_n925_), .B1(men_men_n567_), .Y(men_men_n971_));
  NO2        u0943(.A(men_men_n624_), .B(men_men_n354_), .Y(men_men_n972_));
  NO3        u0944(.A(men_men_n507_), .B(men_men_n138_), .C(men_men_n198_), .Y(men_men_n973_));
  OAI210     u0945(.A0(men_men_n973_), .A1(men_men_n489_), .B0(men_men_n355_), .Y(men_men_n974_));
  NA2        u0946(.A(men_men_n974_), .B(men_men_n585_), .Y(men_men_n975_));
  OAI210     u0947(.A0(men_men_n886_), .A1(men_men_n881_), .B0(men_men_n963_), .Y(men_men_n976_));
  NA3        u0948(.A(men_men_n921_), .B(men_men_n454_), .C(men_men_n46_), .Y(men_men_n977_));
  NA2        u0949(.A(men_men_n357_), .B(men_men_n355_), .Y(men_men_n978_));
  NA4        u0950(.A(men_men_n978_), .B(men_men_n977_), .C(men_men_n976_), .D(men_men_n255_), .Y(men_men_n979_));
  OR4        u0951(.A(men_men_n979_), .B(men_men_n975_), .C(men_men_n972_), .D(men_men_n971_), .Y(men_men_n980_));
  NO4        u0952(.A(men_men_n980_), .B(men_men_n970_), .C(men_men_n965_), .D(men_men_n962_), .Y(men_men_n981_));
  NA4        u0953(.A(men_men_n981_), .B(men_men_n955_), .C(men_men_n914_), .D(men_men_n900_), .Y(men13));
  NA2        u0954(.A(men_men_n46_), .B(men_men_n77_), .Y(men_men_n983_));
  NA3        u0955(.A(men_men_n233_), .B(c), .C(m), .Y(men_men_n984_));
  NO3        u0956(.A(men_men_n984_), .B(men_men_n983_), .C(men_men_n545_), .Y(men_men_n985_));
  NA2        u0957(.A(men_men_n246_), .B(c), .Y(men_men_n986_));
  NO3        u0958(.A(men_men_n986_), .B(men_men_n916_), .C(a), .Y(men_men_n987_));
  NA2        u0959(.A(men_men_n129_), .B(men_men_n45_), .Y(men_men_n988_));
  NO4        u0960(.A(men_men_n988_), .B(c), .C(men_men_n552_), .D(men_men_n289_), .Y(men_men_n989_));
  NA2        u0961(.A(men_men_n385_), .B(men_men_n198_), .Y(men_men_n990_));
  AN2        u0962(.A(d), .B(c), .Y(men_men_n991_));
  NA2        u0963(.A(men_men_n991_), .B(men_men_n107_), .Y(men_men_n992_));
  NO3        u0964(.A(men_men_n992_), .B(men_men_n990_), .C(men_men_n166_), .Y(men_men_n993_));
  NA2        u0965(.A(d), .B(c), .Y(men_men_n994_));
  NO4        u0966(.A(men_men_n988_), .B(men_men_n548_), .C(men_men_n994_), .D(men_men_n289_), .Y(men_men_n995_));
  OR2        u0967(.A(men_men_n993_), .B(men_men_n995_), .Y(men_men_n996_));
  OR4        u0968(.A(men_men_n996_), .B(men_men_n989_), .C(men_men_n987_), .D(men_men_n985_), .Y(men_men_n997_));
  NO2        u0969(.A(f), .B(men_men_n135_), .Y(men_men_n998_));
  NA2        u0970(.A(men_men_n998_), .B(u), .Y(men_men_n999_));
  OR2        u0971(.A(men_men_n210_), .B(men_men_n166_), .Y(men_men_n1000_));
  NO2        u0972(.A(men_men_n1000_), .B(men_men_n999_), .Y(men_men_n1001_));
  NO2        u0973(.A(men_men_n994_), .B(men_men_n289_), .Y(men_men_n1002_));
  INV        u0974(.A(men_men_n595_), .Y(men_men_n1003_));
  NOi21      u0975(.An(men_men_n1002_), .B(men_men_n1003_), .Y(men_men_n1004_));
  NOi41      u0976(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1005_));
  NA2        u0977(.A(men_men_n1005_), .B(j), .Y(men_men_n1006_));
  NO2        u0978(.A(men_men_n1006_), .B(men_men_n999_), .Y(men_men_n1007_));
  OR3        u0979(.A(e), .B(d), .C(c), .Y(men_men_n1008_));
  NA3        u0980(.A(k), .B(j), .C(i), .Y(men_men_n1009_));
  NO3        u0981(.A(men_men_n1009_), .B(men_men_n289_), .C(men_men_n81_), .Y(men_men_n1010_));
  NOi21      u0982(.An(men_men_n1010_), .B(men_men_n1008_), .Y(men_men_n1011_));
  OR4        u0983(.A(men_men_n1011_), .B(men_men_n1007_), .C(men_men_n1004_), .D(men_men_n1001_), .Y(men_men_n1012_));
  NA2        u0984(.A(men_men_n438_), .B(men_men_n310_), .Y(men_men_n1013_));
  NO2        u0985(.A(men_men_n1013_), .B(men_men_n1003_), .Y(men_men_n1014_));
  NO4        u0986(.A(men_men_n1013_), .B(men_men_n548_), .C(men_men_n424_), .D(men_men_n45_), .Y(men_men_n1015_));
  NO2        u0987(.A(f), .B(c), .Y(men_men_n1016_));
  NOi21      u0988(.An(men_men_n1016_), .B(men_men_n417_), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n1017_), .B(men_men_n56_), .Y(men_men_n1018_));
  NO3        u0990(.A(i), .B(h), .C(l), .Y(men_men_n1019_));
  NOi21      u0991(.An(men_men_n1019_), .B(men_men_n1018_), .Y(men_men_n1020_));
  OR3        u0992(.A(men_men_n1020_), .B(men_men_n1015_), .C(men_men_n1014_), .Y(men_men_n1021_));
  OR3        u0993(.A(men_men_n1021_), .B(men_men_n1012_), .C(men_men_n997_), .Y(men02));
  OR3        u0994(.A(h), .B(u), .C(f), .Y(men_men_n1023_));
  OR3        u0995(.A(n), .B(m), .C(i), .Y(men_men_n1024_));
  NO4        u0996(.A(men_men_n1024_), .B(men_men_n1023_), .C(l), .D(men_men_n1008_), .Y(men_men_n1025_));
  NOi31      u0997(.An(e), .B(d), .C(c), .Y(men_men_n1026_));
  AOI210     u0998(.A0(men_men_n1010_), .A1(men_men_n1026_), .B0(men_men_n989_), .Y(men_men_n1027_));
  NA3        u0999(.A(u), .B(men_men_n438_), .C(h), .Y(men_men_n1028_));
  OR2        u1000(.A(men_men_n1009_), .B(men_men_n1028_), .Y(men_men_n1029_));
  NO3        u1001(.A(men_men_n1013_), .B(men_men_n988_), .C(men_men_n548_), .Y(men_men_n1030_));
  NO2        u1002(.A(men_men_n1030_), .B(men_men_n1001_), .Y(men_men_n1031_));
  NA2        u1003(.A(i), .B(h), .Y(men_men_n1032_));
  INV        u1004(.A(men_men_n1004_), .Y(men_men_n1033_));
  NA3        u1005(.A(c), .B(b), .C(a), .Y(men_men_n1034_));
  NO3        u1006(.A(men_men_n1034_), .B(men_men_n856_), .C(men_men_n198_), .Y(men_men_n1035_));
  INV        u1007(.A(men_men_n1014_), .Y(men_men_n1036_));
  AN4        u1008(.A(men_men_n1036_), .B(men_men_n1033_), .C(men_men_n1031_), .D(men_men_n1029_), .Y(men_men_n1037_));
  NO2        u1009(.A(men_men_n992_), .B(men_men_n990_), .Y(men_men_n1038_));
  NA2        u1010(.A(men_men_n1006_), .B(men_men_n1000_), .Y(men_men_n1039_));
  AOI210     u1011(.A0(men_men_n1039_), .A1(men_men_n1038_), .B0(men_men_n985_), .Y(men_men_n1040_));
  NAi41      u1012(.An(men_men_n1025_), .B(men_men_n1040_), .C(men_men_n1037_), .D(men_men_n1027_), .Y(men03));
  NO2        u1013(.A(men_men_n491_), .B(men_men_n561_), .Y(men_men_n1042_));
  NA4        u1014(.A(men_men_n78_), .B(men_men_n77_), .C(u), .D(men_men_n198_), .Y(men_men_n1043_));
  NA4        u1015(.A(men_men_n538_), .B(m), .C(men_men_n103_), .D(men_men_n198_), .Y(men_men_n1044_));
  NA3        u1016(.A(men_men_n1044_), .B(men_men_n345_), .C(men_men_n1043_), .Y(men_men_n1045_));
  NO3        u1017(.A(men_men_n1045_), .B(men_men_n1042_), .C(men_men_n949_), .Y(men_men_n1046_));
  NOi41      u1018(.An(men_men_n765_), .B(men_men_n814_), .C(men_men_n803_), .D(men_men_n671_), .Y(men_men_n1047_));
  OAI220     u1019(.A0(men_men_n1047_), .A1(men_men_n648_), .B0(men_men_n1046_), .B1(men_men_n549_), .Y(men_men_n1048_));
  NA4        u1020(.A(i), .B(men_men_n1026_), .C(men_men_n318_), .D(men_men_n310_), .Y(men_men_n1049_));
  OAI210     u1021(.A0(men_men_n780_), .A1(men_men_n396_), .B0(men_men_n1049_), .Y(men_men_n1050_));
  NOi31      u1022(.An(m), .B(n), .C(f), .Y(men_men_n1051_));
  AN2        u1023(.A(e), .B(c), .Y(men_men_n1052_));
  NA2        u1024(.A(men_men_n473_), .B(l), .Y(men_men_n1053_));
  NO2        u1025(.A(men_men_n1050_), .B(men_men_n948_), .Y(men_men_n1054_));
  NO2        u1026(.A(men_men_n265_), .B(a), .Y(men_men_n1055_));
  INV        u1027(.A(men_men_n989_), .Y(men_men_n1056_));
  NO2        u1028(.A(men_men_n1032_), .B(men_men_n453_), .Y(men_men_n1057_));
  NO2        u1029(.A(men_men_n77_), .B(u), .Y(men_men_n1058_));
  NO2        u1030(.A(men_men_n1057_), .B(men_men_n1019_), .Y(men_men_n1059_));
  OR2        u1031(.A(men_men_n1059_), .B(men_men_n1018_), .Y(men_men_n1060_));
  NA3        u1032(.A(men_men_n1060_), .B(men_men_n1056_), .C(men_men_n1054_), .Y(men_men_n1061_));
  NO4        u1033(.A(men_men_n1061_), .B(men_men_n1048_), .C(men_men_n782_), .D(men_men_n528_), .Y(men_men_n1062_));
  NA2        u1034(.A(c), .B(b), .Y(men_men_n1063_));
  NO2        u1035(.A(men_men_n658_), .B(men_men_n1063_), .Y(men_men_n1064_));
  OAI210     u1036(.A0(men_men_n821_), .A1(men_men_n794_), .B0(men_men_n389_), .Y(men_men_n1065_));
  NA2        u1037(.A(men_men_n1065_), .B(men_men_n1064_), .Y(men_men_n1066_));
  NAi21      u1038(.An(men_men_n397_), .B(men_men_n1064_), .Y(men_men_n1067_));
  NA3        u1039(.A(men_men_n403_), .B(men_men_n521_), .C(f), .Y(men_men_n1068_));
  NA2        u1040(.A(men_men_n39_), .B(men_men_n1055_), .Y(men_men_n1069_));
  NA3        u1041(.A(men_men_n1069_), .B(men_men_n1068_), .C(men_men_n1067_), .Y(men_men_n1070_));
  OAI210     u1042(.A0(men_men_n109_), .A1(men_men_n269_), .B0(u), .Y(men_men_n1071_));
  NAi21      u1043(.An(f), .B(d), .Y(men_men_n1072_));
  NO2        u1044(.A(men_men_n1072_), .B(men_men_n1034_), .Y(men_men_n1073_));
  INV        u1045(.A(men_men_n1073_), .Y(men_men_n1074_));
  NO2        u1046(.A(men_men_n1071_), .B(men_men_n1074_), .Y(men_men_n1075_));
  AOI210     u1047(.A0(men_men_n1075_), .A1(men_men_n104_), .B0(men_men_n1070_), .Y(men_men_n1076_));
  NA2        u1048(.A(men_men_n440_), .B(men_men_n439_), .Y(men_men_n1077_));
  NO2        u1049(.A(men_men_n172_), .B(men_men_n222_), .Y(men_men_n1078_));
  NA2        u1050(.A(men_men_n1078_), .B(m), .Y(men_men_n1079_));
  NA3        u1051(.A(men_men_n870_), .B(men_men_n1053_), .C(men_men_n443_), .Y(men_men_n1080_));
  INV        u1052(.A(men_men_n441_), .Y(men_men_n1081_));
  AOI210     u1053(.A0(men_men_n1081_), .A1(men_men_n1077_), .B0(men_men_n1079_), .Y(men_men_n1082_));
  NA2        u1054(.A(men_men_n523_), .B(men_men_n384_), .Y(men_men_n1083_));
  NA2        u1055(.A(men_men_n33_), .B(men_men_n1073_), .Y(men_men_n1084_));
  NO2        u1056(.A(men_men_n348_), .B(men_men_n347_), .Y(men_men_n1085_));
  AOI210     u1057(.A0(men_men_n1078_), .A1(men_men_n405_), .B0(men_men_n908_), .Y(men_men_n1086_));
  NAi41      u1058(.An(men_men_n1085_), .B(men_men_n1086_), .C(men_men_n1084_), .D(men_men_n1083_), .Y(men_men_n1087_));
  NO2        u1059(.A(men_men_n1087_), .B(men_men_n1082_), .Y(men_men_n1088_));
  NA4        u1060(.A(men_men_n1088_), .B(men_men_n1076_), .C(men_men_n1066_), .D(men_men_n1062_), .Y(men00));
  NO2        u1061(.A(men_men_n282_), .B(men_men_n257_), .Y(men_men_n1090_));
  NO2        u1062(.A(men_men_n1090_), .B(men_men_n540_), .Y(men_men_n1091_));
  AOI210     u1063(.A0(men_men_n853_), .A1(men_men_n892_), .B0(men_men_n1050_), .Y(men_men_n1092_));
  NO3        u1064(.A(men_men_n1030_), .B(men_men_n908_), .C(men_men_n668_), .Y(men_men_n1093_));
  NA3        u1065(.A(men_men_n1093_), .B(men_men_n1092_), .C(men_men_n950_), .Y(men_men_n1094_));
  NA2        u1066(.A(men_men_n282_), .B(f), .Y(men_men_n1095_));
  OAI210     u1067(.A0(men_men_n957_), .A1(men_men_n40_), .B0(men_men_n613_), .Y(men_men_n1096_));
  NA3        u1068(.A(men_men_n1096_), .B(u), .C(n), .Y(men_men_n1097_));
  AOI210     u1069(.A0(men_men_n1097_), .A1(men_men_n1095_), .B0(men_men_n992_), .Y(men_men_n1098_));
  NO4        u1070(.A(men_men_n1098_), .B(men_men_n1094_), .C(men_men_n1091_), .D(men_men_n1012_), .Y(men_men_n1099_));
  NA3        u1071(.A(men_men_n157_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1100_));
  NA3        u1072(.A(d), .B(men_men_n54_), .C(b), .Y(men_men_n1101_));
  NOi31      u1073(.An(n), .B(m), .C(i), .Y(men_men_n1102_));
  NA3        u1074(.A(men_men_n1102_), .B(men_men_n616_), .C(men_men_n51_), .Y(men_men_n1103_));
  OAI210     u1075(.A0(men_men_n1101_), .A1(men_men_n1100_), .B0(men_men_n1103_), .Y(men_men_n1104_));
  NO3        u1076(.A(men_men_n1104_), .B(men_men_n1085_), .C(men_men_n873_), .Y(men_men_n1105_));
  NA3        u1077(.A(men_men_n360_), .B(men_men_n206_), .C(u), .Y(men_men_n1106_));
  OR2        u1078(.A(men_men_n361_), .B(men_men_n123_), .Y(men_men_n1107_));
  NO2        u1079(.A(h), .B(u), .Y(men_men_n1108_));
  NA4        u1080(.A(men_men_n464_), .B(men_men_n438_), .C(men_men_n1108_), .D(c), .Y(men_men_n1109_));
  OAI220     u1081(.A0(men_men_n491_), .A1(men_men_n561_), .B0(men_men_n82_), .B1(men_men_n81_), .Y(men_men_n1110_));
  AOI220     u1082(.A0(men_men_n1110_), .A1(men_men_n498_), .B0(men_men_n895_), .B1(men_men_n539_), .Y(men_men_n1111_));
  AOI220     u1083(.A0(men_men_n299_), .A1(men_men_n230_), .B0(men_men_n167_), .B1(men_men_n137_), .Y(men_men_n1112_));
  NA4        u1084(.A(men_men_n1112_), .B(men_men_n1111_), .C(men_men_n1109_), .D(men_men_n1107_), .Y(men_men_n1113_));
  NO2        u1085(.A(men_men_n1113_), .B(men_men_n248_), .Y(men_men_n1114_));
  INV        u1086(.A(men_men_n303_), .Y(men_men_n1115_));
  INV        u1087(.A(men_men_n541_), .Y(men_men_n1116_));
  NA3        u1088(.A(men_men_n1116_), .B(men_men_n1115_), .C(men_men_n143_), .Y(men_men_n1117_));
  NA3        u1089(.A(men_men_n438_), .B(men_men_n40_), .C(f), .Y(men_men_n1118_));
  NOi21      u1090(.An(men_men_n829_), .B(men_men_n1118_), .Y(men_men_n1119_));
  NAi31      u1091(.An(men_men_n173_), .B(men_men_n818_), .C(men_men_n438_), .Y(men_men_n1120_));
  NAi21      u1092(.An(men_men_n1119_), .B(men_men_n1120_), .Y(men_men_n1121_));
  NO2        u1093(.A(men_men_n256_), .B(men_men_n69_), .Y(men_men_n1122_));
  NO3        u1094(.A(men_men_n402_), .B(men_men_n792_), .C(n), .Y(men_men_n1123_));
  AOI210     u1095(.A0(men_men_n1123_), .A1(men_men_n1122_), .B0(men_men_n1025_), .Y(men_men_n1124_));
  NAi21      u1096(.An(men_men_n995_), .B(men_men_n1124_), .Y(men_men_n1125_));
  NO4        u1097(.A(men_men_n1125_), .B(men_men_n1121_), .C(men_men_n1117_), .D(men_men_n482_), .Y(men_men_n1126_));
  AN3        u1098(.A(men_men_n1126_), .B(men_men_n1114_), .C(men_men_n1105_), .Y(men_men_n1127_));
  NA2        u1099(.A(men_men_n498_), .B(men_men_n92_), .Y(men_men_n1128_));
  NA3        u1100(.A(men_men_n524_), .B(men_men_n1128_), .C(men_men_n227_), .Y(men_men_n1129_));
  NA2        u1101(.A(men_men_n1045_), .B(men_men_n498_), .Y(men_men_n1130_));
  NA4        u1102(.A(men_men_n616_), .B(men_men_n191_), .C(men_men_n206_), .D(men_men_n152_), .Y(men_men_n1131_));
  NA3        u1103(.A(men_men_n1131_), .B(men_men_n1130_), .C(men_men_n279_), .Y(men_men_n1132_));
  OAI210     u1104(.A0(men_men_n437_), .A1(men_men_n111_), .B0(men_men_n823_), .Y(men_men_n1133_));
  AOI220     u1105(.A0(men_men_n1133_), .A1(men_men_n1080_), .B0(men_men_n523_), .B1(men_men_n384_), .Y(men_men_n1134_));
  OR3        u1106(.A(men_men_n992_), .B(men_men_n254_), .C(men_men_n208_), .Y(men_men_n1135_));
  NO2        u1107(.A(men_men_n202_), .B(men_men_n199_), .Y(men_men_n1136_));
  NA2        u1108(.A(n), .B(e), .Y(men_men_n1137_));
  NO2        u1109(.A(men_men_n1137_), .B(men_men_n135_), .Y(men_men_n1138_));
  NA2        u1110(.A(men_men_n807_), .B(men_men_n1136_), .Y(men_men_n1139_));
  OAI210     u1111(.A0(men_men_n333_), .A1(men_men_n294_), .B0(men_men_n423_), .Y(men_men_n1140_));
  NA4        u1112(.A(men_men_n1140_), .B(men_men_n1139_), .C(men_men_n1135_), .D(men_men_n1134_), .Y(men_men_n1141_));
  AOI210     u1113(.A0(men_men_n1138_), .A1(men_men_n811_), .B0(men_men_n781_), .Y(men_men_n1142_));
  NO2        u1114(.A(men_men_n65_), .B(h), .Y(men_men_n1143_));
  NO3        u1115(.A(men_men_n992_), .B(men_men_n990_), .C(men_men_n685_), .Y(men_men_n1144_));
  INV        u1116(.A(men_men_n1144_), .Y(men_men_n1145_));
  NA3        u1117(.A(men_men_n1145_), .B(men_men_n1142_), .C(men_men_n825_), .Y(men_men_n1146_));
  NO4        u1118(.A(men_men_n1146_), .B(men_men_n1141_), .C(men_men_n1132_), .D(men_men_n1129_), .Y(men_men_n1147_));
  NA2        u1119(.A(men_men_n795_), .B(men_men_n718_), .Y(men_men_n1148_));
  NA4        u1120(.A(men_men_n1148_), .B(men_men_n1147_), .C(men_men_n1127_), .D(men_men_n1099_), .Y(men01));
  NO3        u1121(.A(men_men_n761_), .B(men_men_n754_), .C(men_men_n263_), .Y(men_men_n1150_));
  NA2        u1122(.A(men_men_n1150_), .B(men_men_n974_), .Y(men_men_n1151_));
  NA2        u1123(.A(men_men_n550_), .B(men_men_n80_), .Y(men_men_n1152_));
  NA2        u1124(.A(men_men_n517_), .B(men_men_n253_), .Y(men_men_n1153_));
  NA2        u1125(.A(men_men_n911_), .B(men_men_n1153_), .Y(men_men_n1154_));
  NA4        u1126(.A(men_men_n1154_), .B(men_men_n1152_), .C(men_men_n866_), .D(men_men_n309_), .Y(men_men_n1155_));
  NA2        u1127(.A(men_men_n665_), .B(men_men_n87_), .Y(men_men_n1156_));
  NO2        u1128(.A(men_men_n1156_), .B(i), .Y(men_men_n1157_));
  OAI210     u1129(.A0(men_men_n741_), .A1(men_men_n567_), .B0(men_men_n1131_), .Y(men_men_n1158_));
  AOI210     u1130(.A0(men_men_n1157_), .A1(men_men_n602_), .B0(men_men_n1158_), .Y(men_men_n1159_));
  INV        u1131(.A(men_men_n109_), .Y(men_men_n1160_));
  OA220      u1132(.A0(men_men_n1160_), .A1(men_men_n547_), .B0(men_men_n625_), .B1(men_men_n345_), .Y(men_men_n1161_));
  NAi41      u1133(.An(men_men_n151_), .B(men_men_n1161_), .C(men_men_n1159_), .D(men_men_n852_), .Y(men_men_n1162_));
  NO3        u1134(.A(men_men_n742_), .B(men_men_n638_), .C(men_men_n475_), .Y(men_men_n1163_));
  OR2        u1135(.A(men_men_n180_), .B(men_men_n178_), .Y(men_men_n1164_));
  NA3        u1136(.A(men_men_n1164_), .B(men_men_n1163_), .C(men_men_n126_), .Y(men_men_n1165_));
  NO4        u1137(.A(men_men_n1165_), .B(men_men_n1162_), .C(men_men_n1155_), .D(men_men_n1151_), .Y(men_men_n1166_));
  NA2        u1138(.A(men_men_n1106_), .B(men_men_n192_), .Y(men_men_n1167_));
  OAI210     u1139(.A0(men_men_n1167_), .A1(men_men_n285_), .B0(men_men_n493_), .Y(men_men_n1168_));
  NA2        u1140(.A(men_men_n501_), .B(men_men_n370_), .Y(men_men_n1169_));
  BUFFER     u1141(.A(men_men_n525_), .Y(men_men_n1170_));
  NA2        u1142(.A(men_men_n1170_), .B(men_men_n1169_), .Y(men_men_n1171_));
  AOI210     u1143(.A0(men_men_n189_), .A1(men_men_n79_), .B0(men_men_n198_), .Y(men_men_n1172_));
  OAI210     u1144(.A0(men_men_n768_), .A1(men_men_n403_), .B0(men_men_n1172_), .Y(men_men_n1173_));
  OAI210     u1145(.A0(men_men_n335_), .A1(men_men_n34_), .B0(l), .Y(men_men_n1174_));
  NA2        u1146(.A(men_men_n188_), .B(men_men_n34_), .Y(men_men_n1175_));
  AO210      u1147(.A0(men_men_n1175_), .A1(men_men_n1174_), .B0(men_men_n308_), .Y(men_men_n1176_));
  NA4        u1148(.A(men_men_n1176_), .B(men_men_n1173_), .C(men_men_n1171_), .D(men_men_n1168_), .Y(men_men_n1177_));
  AOI210     u1149(.A0(men_men_n559_), .A1(men_men_n109_), .B0(men_men_n565_), .Y(men_men_n1178_));
  OAI210     u1150(.A0(men_men_n1160_), .A1(men_men_n556_), .B0(men_men_n1178_), .Y(men_men_n1179_));
  NA2        u1151(.A(men_men_n262_), .B(men_men_n180_), .Y(men_men_n1180_));
  NA2        u1152(.A(men_men_n1180_), .B(men_men_n630_), .Y(men_men_n1181_));
  NO3        u1153(.A(men_men_n780_), .B(men_men_n189_), .C(men_men_n382_), .Y(men_men_n1182_));
  NO2        u1154(.A(men_men_n1182_), .B(men_men_n908_), .Y(men_men_n1183_));
  NA3        u1155(.A(men_men_n1183_), .B(men_men_n1181_), .C(men_men_n745_), .Y(men_men_n1184_));
  NO3        u1156(.A(men_men_n1184_), .B(men_men_n1179_), .C(men_men_n1177_), .Y(men_men_n1185_));
  NA3        u1157(.A(men_men_n568_), .B(men_men_n29_), .C(f), .Y(men_men_n1186_));
  NO2        u1158(.A(men_men_n1186_), .B(men_men_n189_), .Y(men_men_n1187_));
  INV        u1159(.A(men_men_n1187_), .Y(men_men_n1188_));
  OR3        u1160(.A(men_men_n1156_), .B(men_men_n569_), .C(i), .Y(men_men_n1189_));
  NO2        u1161(.A(men_men_n192_), .B(men_men_n102_), .Y(men_men_n1190_));
  NO2        u1162(.A(men_men_n1190_), .B(men_men_n1104_), .Y(men_men_n1191_));
  NA4        u1163(.A(men_men_n1191_), .B(men_men_n1189_), .C(men_men_n1188_), .D(men_men_n717_), .Y(men_men_n1192_));
  NA2        u1164(.A(men_men_n535_), .B(men_men_n533_), .Y(men_men_n1193_));
  NO3        u1165(.A(m), .B(men_men_n283_), .C(men_men_n45_), .Y(men_men_n1194_));
  NA2        u1166(.A(men_men_n1194_), .B(men_men_n516_), .Y(men_men_n1195_));
  NA3        u1167(.A(men_men_n1195_), .B(men_men_n1193_), .C(men_men_n634_), .Y(men_men_n1196_));
  INV        u1168(.A(men_men_n363_), .Y(men_men_n1197_));
  NO3        u1169(.A(men_men_n1197_), .B(men_men_n1196_), .C(men_men_n1192_), .Y(men_men_n1198_));
  AO220      u1170(.A0(i), .A1(men_men_n588_), .B0(i), .B1(men_men_n663_), .Y(men_men_n1199_));
  NO3        u1171(.A(men_men_n1032_), .B(men_men_n166_), .C(men_men_n77_), .Y(men_men_n1200_));
  NO2        u1172(.A(men_men_n579_), .B(men_men_n578_), .Y(men_men_n1201_));
  NO4        u1173(.A(men_men_n1032_), .B(men_men_n1201_), .C(men_men_n164_), .D(men_men_n77_), .Y(men_men_n1202_));
  NO3        u1174(.A(men_men_n1202_), .B(men_men_n1200_), .C(men_men_n606_), .Y(men_men_n1203_));
  NA4        u1175(.A(men_men_n1203_), .B(men_men_n1198_), .C(men_men_n1185_), .D(men_men_n1166_), .Y(men06));
  NO2        u1176(.A(men_men_n383_), .B(men_men_n522_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n249_), .B(men_men_n1205_), .Y(men_men_n1206_));
  NO2        u1178(.A(men_men_n210_), .B(men_men_n94_), .Y(men_men_n1207_));
  OAI210     u1179(.A0(men_men_n1207_), .A1(men_men_n1200_), .B0(men_men_n359_), .Y(men_men_n1208_));
  NO3        u1180(.A(men_men_n563_), .B(men_men_n766_), .C(men_men_n566_), .Y(men_men_n1209_));
  OR2        u1181(.A(men_men_n1209_), .B(men_men_n841_), .Y(men_men_n1210_));
  NA3        u1182(.A(men_men_n1210_), .B(men_men_n1208_), .C(men_men_n1206_), .Y(men_men_n1211_));
  NO3        u1183(.A(men_men_n1211_), .B(men_men_n1196_), .C(men_men_n240_), .Y(men_men_n1212_));
  NO2        u1184(.A(men_men_n283_), .B(men_men_n45_), .Y(men_men_n1213_));
  NA2        u1185(.A(men_men_n1213_), .B(men_men_n920_), .Y(men_men_n1214_));
  AOI210     u1186(.A0(men_men_n1213_), .A1(men_men_n519_), .B0(men_men_n1199_), .Y(men_men_n1215_));
  AOI210     u1187(.A0(men_men_n1215_), .A1(men_men_n1214_), .B0(men_men_n314_), .Y(men_men_n1216_));
  OAI210     u1188(.A0(men_men_n79_), .A1(men_men_n40_), .B0(men_men_n637_), .Y(men_men_n1217_));
  NA2        u1189(.A(men_men_n1217_), .B(men_men_n610_), .Y(men_men_n1218_));
  NO2        u1190(.A(men_men_n432_), .B(men_men_n231_), .Y(men_men_n1219_));
  NO2        u1191(.A(men_men_n1219_), .B(men_men_n125_), .Y(men_men_n1220_));
  OR2        u1192(.A(men_men_n564_), .B(men_men_n562_), .Y(men_men_n1221_));
  INV        u1193(.A(men_men_n1221_), .Y(men_men_n1222_));
  NA3        u1194(.A(men_men_n1222_), .B(men_men_n1220_), .C(men_men_n1218_), .Y(men_men_n1223_));
  NO2        u1195(.A(men_men_n708_), .B(men_men_n343_), .Y(men_men_n1224_));
  NO3        u1196(.A(men_men_n639_), .B(men_men_n719_), .C(men_men_n602_), .Y(men_men_n1225_));
  NOi21      u1197(.An(men_men_n1224_), .B(men_men_n1225_), .Y(men_men_n1226_));
  BUFFER     u1198(.A(men_men_n904_), .Y(men_men_n1227_));
  NO4        u1199(.A(men_men_n1227_), .B(men_men_n1226_), .C(men_men_n1223_), .D(men_men_n1216_), .Y(men_men_n1228_));
  NO2        u1200(.A(men_men_n760_), .B(men_men_n258_), .Y(men_men_n1229_));
  OAI220     u1201(.A0(men_men_n692_), .A1(men_men_n47_), .B0(men_men_n210_), .B1(men_men_n581_), .Y(men_men_n1230_));
  OAI210     u1202(.A0(men_men_n258_), .A1(c), .B0(men_men_n609_), .Y(men_men_n1231_));
  AOI220     u1203(.A0(men_men_n1231_), .A1(men_men_n1230_), .B0(men_men_n1229_), .B1(men_men_n249_), .Y(men_men_n1232_));
  NO2        u1204(.A(men_men_n94_), .B(men_men_n265_), .Y(men_men_n1233_));
  OAI220     u1205(.A0(men_men_n655_), .A1(men_men_n231_), .B0(men_men_n474_), .B1(men_men_n478_), .Y(men_men_n1234_));
  NO2        u1206(.A(men_men_n561_), .B(j), .Y(men_men_n1235_));
  NOi21      u1207(.An(men_men_n1235_), .B(men_men_n68_), .Y(men_men_n1236_));
  NO3        u1208(.A(men_men_n1236_), .B(men_men_n1234_), .C(men_men_n1233_), .Y(men_men_n1237_));
  NA4        u1209(.A(men_men_n752_), .B(men_men_n751_), .C(men_men_n411_), .D(men_men_n835_), .Y(men_men_n1238_));
  NAi31      u1210(.An(men_men_n708_), .B(men_men_n1238_), .C(men_men_n188_), .Y(men_men_n1239_));
  NA3        u1211(.A(men_men_n1239_), .B(men_men_n1237_), .C(men_men_n1232_), .Y(men_men_n1240_));
  OR2        u1212(.A(men_men_n741_), .B(men_men_n504_), .Y(men_men_n1241_));
  OR3        u1213(.A(men_men_n347_), .B(men_men_n210_), .C(men_men_n581_), .Y(men_men_n1242_));
  AOI210     u1214(.A0(men_men_n535_), .A1(men_men_n423_), .B0(men_men_n349_), .Y(men_men_n1243_));
  NA2        u1215(.A(men_men_n1235_), .B(men_men_n748_), .Y(men_men_n1244_));
  NA4        u1216(.A(men_men_n1244_), .B(men_men_n1243_), .C(men_men_n1242_), .D(men_men_n1241_), .Y(men_men_n1245_));
  NA2        u1217(.A(men_men_n1224_), .B(men_men_n718_), .Y(men_men_n1246_));
  INV        u1218(.A(men_men_n1246_), .Y(men_men_n1247_));
  NAi21      u1219(.An(j), .B(i), .Y(men_men_n1248_));
  NO4        u1220(.A(men_men_n1201_), .B(men_men_n1248_), .C(men_men_n417_), .D(men_men_n220_), .Y(men_men_n1249_));
  NO4        u1221(.A(men_men_n1249_), .B(men_men_n1247_), .C(men_men_n1245_), .D(men_men_n1240_), .Y(men_men_n1250_));
  NA4        u1222(.A(men_men_n1250_), .B(men_men_n1228_), .C(men_men_n1212_), .D(men_men_n1203_), .Y(men07));
  NOi21      u1223(.An(j), .B(k), .Y(men_men_n1252_));
  NAi32      u1224(.An(m), .Bn(b), .C(n), .Y(men_men_n1253_));
  NO3        u1225(.A(men_men_n1253_), .B(u), .C(f), .Y(men_men_n1254_));
  OAI210     u1226(.A0(i), .A1(men_men_n452_), .B0(men_men_n1254_), .Y(men_men_n1255_));
  NAi21      u1227(.An(f), .B(c), .Y(men_men_n1256_));
  OR2        u1228(.A(e), .B(d), .Y(men_men_n1257_));
  OAI220     u1229(.A0(men_men_n1257_), .A1(men_men_n1256_), .B0(men_men_n594_), .B1(men_men_n304_), .Y(men_men_n1258_));
  NA2        u1230(.A(men_men_n1258_), .B(men_men_n169_), .Y(men_men_n1259_));
  NOi31      u1231(.An(n), .B(m), .C(b), .Y(men_men_n1260_));
  NA2        u1232(.A(men_men_n1259_), .B(men_men_n1255_), .Y(men_men_n1261_));
  NOi41      u1233(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1262_));
  NA3        u1234(.A(men_men_n1262_), .B(men_men_n826_), .C(men_men_n385_), .Y(men_men_n1263_));
  NO2        u1235(.A(men_men_n1263_), .B(men_men_n54_), .Y(men_men_n1264_));
  NA2        u1236(.A(b), .B(men_men_n206_), .Y(men_men_n1265_));
  NO2        u1237(.A(men_men_n1265_), .B(men_men_n58_), .Y(men_men_n1266_));
  NO2        u1238(.A(k), .B(i), .Y(men_men_n1267_));
  NA2        u1239(.A(men_men_n1143_), .B(men_men_n273_), .Y(men_men_n1268_));
  INV        u1240(.A(men_men_n1268_), .Y(men_men_n1269_));
  NO4        u1241(.A(men_men_n1269_), .B(men_men_n1266_), .C(men_men_n1264_), .D(men_men_n1261_), .Y(men_men_n1270_));
  NO3        u1242(.A(e), .B(d), .C(c), .Y(men_men_n1271_));
  OAI210     u1243(.A0(men_men_n122_), .A1(men_men_n199_), .B0(men_men_n570_), .Y(men_men_n1272_));
  NA2        u1244(.A(men_men_n1272_), .B(men_men_n1271_), .Y(men_men_n1273_));
  INV        u1245(.A(men_men_n1273_), .Y(men_men_n1274_));
  NO3        u1246(.A(n), .B(m), .C(i), .Y(men_men_n1275_));
  OAI210     u1247(.A0(men_men_n1052_), .A1(men_men_n146_), .B0(men_men_n1275_), .Y(men_men_n1276_));
  NO2        u1248(.A(i), .B(u), .Y(men_men_n1277_));
  OR3        u1249(.A(men_men_n1277_), .B(men_men_n1253_), .C(e), .Y(men_men_n1278_));
  OAI220     u1250(.A0(men_men_n1278_), .A1(men_men_n452_), .B0(men_men_n1276_), .B1(f), .Y(men_men_n1279_));
  NA3        u1251(.A(men_men_n652_), .B(men_men_n1397_), .C(men_men_n103_), .Y(men_men_n1280_));
  NA3        u1252(.A(men_men_n1260_), .B(j), .C(h), .Y(men_men_n1281_));
  AOI210     u1253(.A0(men_men_n1281_), .A1(men_men_n1280_), .B0(men_men_n45_), .Y(men_men_n1282_));
  NA2        u1254(.A(men_men_n1275_), .B(men_men_n608_), .Y(men_men_n1283_));
  NO3        u1255(.A(men_men_n1282_), .B(men_men_n1279_), .C(men_men_n1274_), .Y(men_men_n1284_));
  NO2        u1256(.A(men_men_n136_), .B(h), .Y(men_men_n1285_));
  NO2        u1257(.A(men_men_n425_), .B(a), .Y(men_men_n1286_));
  NA3        u1258(.A(men_men_n1286_), .B(k), .C(men_men_n104_), .Y(men_men_n1287_));
  NO2        u1259(.A(i), .B(h), .Y(men_men_n1288_));
  NA2        u1260(.A(men_men_n1072_), .B(h), .Y(men_men_n1289_));
  NA2        u1261(.A(men_men_n127_), .B(men_men_n206_), .Y(men_men_n1290_));
  NO2        u1262(.A(men_men_n1290_), .B(men_men_n1289_), .Y(men_men_n1291_));
  NO2        u1263(.A(men_men_n715_), .B(men_men_n174_), .Y(men_men_n1292_));
  NOi31      u1264(.An(m), .B(n), .C(b), .Y(men_men_n1293_));
  NOi31      u1265(.An(f), .B(d), .C(c), .Y(men_men_n1294_));
  NA2        u1266(.A(men_men_n1294_), .B(men_men_n1293_), .Y(men_men_n1295_));
  INV        u1267(.A(men_men_n1295_), .Y(men_men_n1296_));
  NO3        u1268(.A(men_men_n1296_), .B(men_men_n1292_), .C(men_men_n1291_), .Y(men_men_n1297_));
  NA2        u1269(.A(men_men_n490_), .B(men_men_n1005_), .Y(men_men_n1298_));
  NO3        u1270(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1299_));
  AN3        u1271(.A(men_men_n1298_), .B(men_men_n1297_), .C(men_men_n1287_), .Y(men_men_n1300_));
  NA2        u1272(.A(men_men_n1260_), .B(men_men_n356_), .Y(men_men_n1301_));
  NO2        u1273(.A(men_men_n174_), .B(b), .Y(men_men_n1302_));
  NA2        u1274(.A(men_men_n1102_), .B(men_men_n1302_), .Y(men_men_n1303_));
  NO2        u1275(.A(i), .B(men_men_n198_), .Y(men_men_n1304_));
  NA4        u1276(.A(men_men_n1078_), .B(men_men_n1304_), .C(men_men_n95_), .D(m), .Y(men_men_n1305_));
  NA2        u1277(.A(men_men_n1305_), .B(men_men_n1303_), .Y(men_men_n1306_));
  NO4        u1278(.A(men_men_n122_), .B(u), .C(f), .D(e), .Y(men_men_n1307_));
  NA2        u1279(.A(men_men_n1267_), .B(h), .Y(men_men_n1308_));
  NA2        u1280(.A(men_men_n30_), .B(h), .Y(men_men_n1309_));
  NO2        u1281(.A(men_men_n1309_), .B(men_men_n1024_), .Y(men_men_n1310_));
  NOi41      u1282(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1311_));
  NA2        u1283(.A(men_men_n1311_), .B(men_men_n104_), .Y(men_men_n1312_));
  INV        u1284(.A(men_men_n1312_), .Y(men_men_n1313_));
  OR3        u1285(.A(men_men_n504_), .B(men_men_n503_), .C(men_men_n103_), .Y(men_men_n1314_));
  NA2        u1286(.A(men_men_n1051_), .B(men_men_n382_), .Y(men_men_n1315_));
  OAI220     u1287(.A0(men_men_n1315_), .A1(men_men_n410_), .B0(men_men_n1314_), .B1(men_men_n283_), .Y(men_men_n1316_));
  AO210      u1288(.A0(men_men_n1316_), .A1(men_men_n107_), .B0(men_men_n1313_), .Y(men_men_n1317_));
  NO3        u1289(.A(men_men_n1317_), .B(men_men_n1310_), .C(men_men_n1306_), .Y(men_men_n1318_));
  NA4        u1290(.A(men_men_n1318_), .B(men_men_n1300_), .C(men_men_n1284_), .D(men_men_n1270_), .Y(men_men_n1319_));
  NO2        u1291(.A(men_men_n1063_), .B(men_men_n101_), .Y(men_men_n1320_));
  AOI210     u1292(.A0(c), .A1(f), .B0(men_men_n1283_), .Y(men_men_n1321_));
  INV        u1293(.A(men_men_n1321_), .Y(men_men_n1322_));
  NA3        u1294(.A(men_men_n1299_), .B(men_men_n1257_), .C(men_men_n1051_), .Y(men_men_n1323_));
  NAi31      u1295(.An(men_men_n1288_), .B(men_men_n1017_), .C(men_men_n158_), .Y(men_men_n1324_));
  NA2        u1296(.A(men_men_n1324_), .B(men_men_n1323_), .Y(men_men_n1325_));
  NO3        u1297(.A(men_men_n708_), .B(men_men_n164_), .C(men_men_n385_), .Y(men_men_n1326_));
  NO2        u1298(.A(men_men_n1326_), .B(men_men_n1325_), .Y(men_men_n1327_));
  NO3        u1299(.A(men_men_n1024_), .B(men_men_n544_), .C(u), .Y(men_men_n1328_));
  INV        u1300(.A(men_men_n1328_), .Y(men_men_n1329_));
  NO2        u1301(.A(men_men_n1329_), .B(f), .Y(men_men_n1330_));
  INV        u1302(.A(men_men_n49_), .Y(men_men_n1331_));
  NA2        u1303(.A(men_men_n1331_), .B(men_men_n1108_), .Y(men_men_n1332_));
  INV        u1304(.A(men_men_n1332_), .Y(men_men_n1333_));
  NA2        u1305(.A(men_men_n1302_), .B(men_men_n41_), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n122_), .B(l), .Y(men_men_n1335_));
  NO2        u1307(.A(men_men_n210_), .B(k), .Y(men_men_n1336_));
  OAI210     u1308(.A0(men_men_n1336_), .A1(men_men_n1288_), .B0(men_men_n1335_), .Y(men_men_n1337_));
  OAI220     u1309(.A0(men_men_n1337_), .A1(men_men_n31_), .B0(men_men_n1334_), .B1(men_men_n166_), .Y(men_men_n1338_));
  NO3        u1310(.A(men_men_n1338_), .B(men_men_n1333_), .C(men_men_n1330_), .Y(men_men_n1339_));
  INV        u1311(.A(men_men_n49_), .Y(men_men_n1340_));
  NA2        u1312(.A(men_men_n1035_), .B(men_men_n1340_), .Y(men_men_n1341_));
  NO2        u1313(.A(men_men_n1024_), .B(h), .Y(men_men_n1342_));
  NA3        u1314(.A(men_men_n1342_), .B(d), .C(men_men_n990_), .Y(men_men_n1343_));
  OAI220     u1315(.A0(men_men_n1343_), .A1(c), .B0(men_men_n1341_), .B1(j), .Y(men_men_n1344_));
  NA3        u1316(.A(men_men_n1320_), .B(men_men_n438_), .C(f), .Y(men_men_n1345_));
  NA2        u1317(.A(men_men_n169_), .B(men_men_n103_), .Y(men_men_n1346_));
  NO2        u1318(.A(men_men_n1252_), .B(men_men_n42_), .Y(men_men_n1347_));
  AOI210     u1319(.A0(men_men_n104_), .A1(men_men_n40_), .B0(men_men_n1347_), .Y(men_men_n1348_));
  NO2        u1320(.A(men_men_n1348_), .B(men_men_n1345_), .Y(men_men_n1349_));
  AOI210     u1321(.A0(men_men_n490_), .A1(h), .B0(men_men_n66_), .Y(men_men_n1350_));
  NA2        u1322(.A(men_men_n1350_), .B(men_men_n1286_), .Y(men_men_n1351_));
  NA2        u1323(.A(men_men_n1286_), .B(men_men_n1347_), .Y(men_men_n1352_));
  NO2        u1324(.A(men_men_n283_), .B(c), .Y(men_men_n1353_));
  NA2        u1325(.A(men_men_n1353_), .B(men_men_n505_), .Y(men_men_n1354_));
  NA3        u1326(.A(men_men_n1354_), .B(men_men_n1352_), .C(men_men_n1351_), .Y(men_men_n1355_));
  NO3        u1327(.A(men_men_n1355_), .B(men_men_n1349_), .C(men_men_n1344_), .Y(men_men_n1356_));
  NA4        u1328(.A(men_men_n1356_), .B(men_men_n1339_), .C(men_men_n1327_), .D(men_men_n1322_), .Y(men_men_n1357_));
  NO2        u1329(.A(c), .B(men_men_n122_), .Y(men_men_n1358_));
  NA3        u1330(.A(b), .B(men_men_n99_), .C(men_men_n206_), .Y(men_men_n1359_));
  NO2        u1331(.A(men_men_n140_), .B(men_men_n171_), .Y(men_men_n1360_));
  OAI210     u1332(.A0(men_men_n1360_), .A1(men_men_n101_), .B0(men_men_n1293_), .Y(men_men_n1361_));
  NA2        u1333(.A(men_men_n1361_), .B(men_men_n1359_), .Y(men_men_n1362_));
  NO2        u1334(.A(men_men_n1362_), .B(men_men_n1358_), .Y(men_men_n1363_));
  NO2        u1335(.A(men_men_n1256_), .B(e), .Y(men_men_n1364_));
  NA2        u1336(.A(men_men_n1364_), .B(men_men_n380_), .Y(men_men_n1365_));
  NA2        u1337(.A(men_men_n1058_), .B(men_men_n598_), .Y(men_men_n1366_));
  OR3        u1338(.A(men_men_n1336_), .B(men_men_n1143_), .C(men_men_n122_), .Y(men_men_n1367_));
  OAI220     u1339(.A0(men_men_n1367_), .A1(men_men_n1365_), .B0(men_men_n1366_), .B1(men_men_n419_), .Y(men_men_n1368_));
  NO3        u1340(.A(men_men_n1314_), .B(men_men_n329_), .C(a), .Y(men_men_n1369_));
  NO2        u1341(.A(men_men_n1369_), .B(men_men_n1368_), .Y(men_men_n1370_));
  NO2        u1342(.A(men_men_n236_), .B(u), .Y(men_men_n1371_));
  NO2        u1343(.A(m), .B(i), .Y(men_men_n1372_));
  BUFFER     u1344(.A(men_men_n1372_), .Y(men_men_n1373_));
  AOI220     u1345(.A0(men_men_n1373_), .A1(men_men_n1285_), .B0(men_men_n1017_), .B1(men_men_n1371_), .Y(men_men_n1374_));
  NA3        u1346(.A(men_men_n1374_), .B(men_men_n1370_), .C(men_men_n1363_), .Y(men_men_n1375_));
  NA3        u1347(.A(men_men_n910_), .B(men_men_n127_), .C(men_men_n46_), .Y(men_men_n1376_));
  AOI210     u1348(.A0(men_men_n146_), .A1(men_men_n54_), .B0(men_men_n1364_), .Y(men_men_n1377_));
  NO2        u1349(.A(men_men_n1377_), .B(men_men_n1346_), .Y(men_men_n1378_));
  NO2        u1350(.A(men_men_n1376_), .B(men_men_n101_), .Y(men_men_n1379_));
  NO2        u1351(.A(men_men_n1379_), .B(men_men_n1378_), .Y(men_men_n1380_));
  NO2        u1352(.A(men_men_n1345_), .B(men_men_n66_), .Y(men_men_n1381_));
  NO2        u1353(.A(men_men_n1267_), .B(men_men_n109_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n1382_), .B(men_men_n1301_), .Y(men_men_n1383_));
  NO2        u1355(.A(men_men_n1383_), .B(men_men_n1381_), .Y(men_men_n1384_));
  NA2        u1356(.A(men_men_n1384_), .B(men_men_n1380_), .Y(men_men_n1385_));
  OR4        u1357(.A(men_men_n1385_), .B(men_men_n1375_), .C(men_men_n1357_), .D(men_men_n1319_), .Y(men04));
  NOi31      u1358(.An(men_men_n1307_), .B(men_men_n1308_), .C(men_men_n992_), .Y(men_men_n1387_));
  NO4        u1359(.A(men_men_n254_), .B(men_men_n984_), .C(men_men_n453_), .D(j), .Y(men_men_n1388_));
  OR3        u1360(.A(men_men_n1388_), .B(men_men_n1387_), .C(men_men_n1007_), .Y(men_men_n1389_));
  NO3        u1361(.A(i), .B(men_men_n81_), .C(k), .Y(men_men_n1390_));
  AOI210     u1362(.A0(men_men_n1390_), .A1(men_men_n1002_), .B0(men_men_n1119_), .Y(men_men_n1391_));
  NA2        u1363(.A(men_men_n1391_), .B(men_men_n1145_), .Y(men_men_n1392_));
  NO4        u1364(.A(men_men_n1392_), .B(men_men_n1389_), .C(men_men_n1015_), .D(men_men_n997_), .Y(men_men_n1393_));
  NA4        u1365(.A(men_men_n1393_), .B(men_men_n1060_), .C(men_men_n1049_), .D(men_men_n1037_), .Y(men05));
  INV        u1366(.A(n), .Y(men_men_n1397_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule