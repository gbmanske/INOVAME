library verilog;
use verilog.vl_types.all;
entity tb_data_driver is
end tb_data_driver;
