library verilog;
use verilog.vl_types.all;
entity freqdiv2_vlg_vec_tst is
end freqdiv2_vlg_vec_tst;
