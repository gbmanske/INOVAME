// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1040_, new_new_n1041_, new_new_n1042_, new_new_n1043_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g0028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g0029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g0032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(i_3_), .B(i_9_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_7_), .Y(new_new_n83_));
  NO3        g0061(.A(new_new_n83_), .B(new_new_n82_), .C(new_new_n63_), .Y(new_new_n84_));
  INV        g0062(.A(i_6_), .Y(new_new_n85_));
  NO2        g0063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  INV        g0064(.A(new_new_n86_), .Y(new_new_n87_));
  NA2        g0065(.A(new_new_n84_), .B(new_new_n87_), .Y(new_new_n88_));
  NAi21      g0066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g0067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g0068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n63_), .Y(new_new_n91_));
  NA2        g0069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g0070(.A(new_new_n92_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g0071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n88_), .B0(new_new_n80_), .Y(new_new_n95_));
  AN3        g0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g0074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g0075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g0076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g0077(.A0(new_new_n99_), .A1(new_new_n62_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g0078(.A(i_7_), .Y(new_new_n101_));
  NA2        g0079(.A(new_new_n46_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g0080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g0081(.A(new_new_n103_), .B(new_new_n85_), .Y(new_new_n104_));
  NA2        g0082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g0083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g0084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g0085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  AN2        g0086(.A(i_2_), .B(i_10_), .Y(new_new_n109_));
  NO2        g0087(.A(new_new_n109_), .B(i_7_), .Y(new_new_n110_));
  OR2        g0088(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n111_));
  NO2        g0089(.A(i_8_), .B(new_new_n101_), .Y(new_new_n112_));
  NO3        g0090(.A(new_new_n112_), .B(new_new_n111_), .C(new_new_n110_), .Y(new_new_n113_));
  NA2        g0091(.A(i_12_), .B(i_7_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n115_));
  NA2        g0093(.A(new_new_n115_), .B(i_0_), .Y(new_new_n116_));
  NA2        g0094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  OAI210     g0095(.A0(new_new_n116_), .A1(new_new_n114_), .B0(new_new_n117_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n118_), .B(new_new_n113_), .Y(new_new_n119_));
  NA3        g0097(.A(new_new_n119_), .B(new_new_n107_), .C(new_new_n100_), .Y(new_new_n120_));
  NOi21      g0098(.An(i_1_), .B(i_5_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n121_), .B(i_11_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g0101(.A(i_7_), .B(new_new_n25_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(new_new_n123_), .Y(new_new_n125_));
  NO2        g0103(.A(new_new_n125_), .B(new_new_n46_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n127_));
  NAi21      g0105(.An(i_3_), .B(i_8_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n62_), .Y(new_new_n129_));
  NOi31      g0107(.An(new_new_n129_), .B(new_new_n127_), .C(new_new_n126_), .Y(new_new_n130_));
  NO2        g0108(.A(i_1_), .B(new_new_n85_), .Y(new_new_n131_));
  NO2        g0109(.A(i_6_), .B(i_5_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(i_3_), .Y(new_new_n133_));
  AO210      g0111(.A0(new_new_n133_), .A1(new_new_n47_), .B0(new_new_n131_), .Y(new_new_n134_));
  OAI220     g0112(.A0(new_new_n134_), .A1(new_new_n108_), .B0(new_new_n130_), .B1(new_new_n122_), .Y(new_new_n135_));
  NO3        g0113(.A(new_new_n135_), .B(new_new_n120_), .C(new_new_n95_), .Y(new_new_n136_));
  NA3        g0114(.A(new_new_n136_), .B(new_new_n79_), .C(new_new_n56_), .Y(men2));
  NO2        g0115(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n138_));
  NA2        g0116(.A(i_6_), .B(new_new_n25_), .Y(new_new_n139_));
  NA2        g0117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g0118(.A(new_new_n140_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(men0));
  AN2        g0119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g0121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g0122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g0123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g0124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g0125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NO2        g0126(.A(new_new_n148_), .B(i_4_), .Y(new_new_n149_));
  NA3        g0127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  OR2        g0128(.A(new_new_n150_), .B(new_new_n25_), .Y(new_new_n151_));
  AN2        g0129(.A(new_new_n144_), .B(new_new_n82_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(new_new_n27_), .Y(new_new_n153_));
  NA2        g0131(.A(i_1_), .B(i_5_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n73_), .B(new_new_n46_), .Y(new_new_n155_));
  NA2        g0133(.A(new_new_n155_), .B(new_new_n36_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n156_), .B(new_new_n154_), .C(new_new_n153_), .Y(new_new_n157_));
  OR2        g0135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n159_));
  NAi32      g0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n160_));
  NAi21      g0138(.An(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NOi21      g0139(.An(i_4_), .B(i_10_), .Y(new_new_n162_));
  NA2        g0140(.A(new_new_n162_), .B(new_new_n40_), .Y(new_new_n163_));
  NO2        g0141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  NO3        g0142(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n165_));
  INV        g0143(.A(new_new_n165_), .Y(new_new_n166_));
  OAI210     g0144(.A0(new_new_n166_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n167_));
  NO2        g0145(.A(new_new_n167_), .B(new_new_n157_), .Y(new_new_n168_));
  AOI210     g0146(.A0(new_new_n168_), .A1(new_new_n151_), .B0(new_new_n143_), .Y(new_new_n169_));
  NA2        g0147(.A(new_new_n46_), .B(i_1_), .Y(new_new_n170_));
  NA2        g0148(.A(i_3_), .B(new_new_n48_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_4_), .B(i_9_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_11_), .B(i_13_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n173_), .B(new_new_n172_), .Y(new_new_n174_));
  OR2        g0152(.A(new_new_n174_), .B(new_new_n171_), .Y(new_new_n175_));
  NO2        g0153(.A(i_4_), .B(i_5_), .Y(new_new_n176_));
  NAi21      g0154(.An(i_12_), .B(i_11_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n177_), .B(i_13_), .Y(new_new_n178_));
  NA3        g0156(.A(new_new_n178_), .B(new_new_n176_), .C(new_new_n82_), .Y(new_new_n179_));
  AOI210     g0157(.A0(new_new_n179_), .A1(new_new_n175_), .B0(new_new_n170_), .Y(new_new_n180_));
  NO2        g0158(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n181_), .B(new_new_n46_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n36_), .B(i_5_), .Y(new_new_n183_));
  NAi31      g0161(.An(new_new_n183_), .B(new_new_n152_), .C(i_11_), .Y(new_new_n184_));
  NA2        g0162(.A(i_3_), .B(i_5_), .Y(new_new_n185_));
  OR2        g0163(.A(new_new_n185_), .B(new_new_n174_), .Y(new_new_n186_));
  AOI210     g0164(.A0(new_new_n186_), .A1(new_new_n184_), .B0(new_new_n182_), .Y(new_new_n187_));
  NO2        g0165(.A(new_new_n73_), .B(i_5_), .Y(new_new_n188_));
  NO2        g0166(.A(i_13_), .B(i_10_), .Y(new_new_n189_));
  NA3        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n44_), .Y(new_new_n190_));
  NO2        g0168(.A(i_2_), .B(i_1_), .Y(new_new_n191_));
  NA2        g0169(.A(new_new_n191_), .B(i_3_), .Y(new_new_n192_));
  NAi21      g0170(.An(i_4_), .B(i_12_), .Y(new_new_n193_));
  NO4        g0171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n190_), .D(new_new_n25_), .Y(new_new_n194_));
  NO3        g0172(.A(new_new_n194_), .B(new_new_n187_), .C(new_new_n180_), .Y(new_new_n195_));
  INV        g0173(.A(i_8_), .Y(new_new_n196_));
  NA2        g0174(.A(i_8_), .B(i_6_), .Y(new_new_n197_));
  NO3        g0175(.A(i_3_), .B(new_new_n85_), .C(new_new_n48_), .Y(new_new_n198_));
  NA2        g0176(.A(new_new_n198_), .B(new_new_n112_), .Y(new_new_n199_));
  NO3        g0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n200_));
  NA3        g0178(.A(new_new_n200_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n201_));
  NO3        g0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n202_));
  OAI210     g0180(.A0(new_new_n96_), .A1(i_12_), .B0(new_new_n202_), .Y(new_new_n203_));
  AOI210     g0181(.A0(new_new_n203_), .A1(new_new_n201_), .B0(new_new_n199_), .Y(new_new_n204_));
  NO2        g0182(.A(i_3_), .B(i_8_), .Y(new_new_n205_));
  NO3        g0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n206_));
  NA3        g0184(.A(new_new_n206_), .B(new_new_n205_), .C(new_new_n40_), .Y(new_new_n207_));
  NO2        g0185(.A(i_13_), .B(i_9_), .Y(new_new_n208_));
  NA3        g0186(.A(new_new_n208_), .B(i_6_), .C(new_new_n196_), .Y(new_new_n209_));
  NAi21      g0187(.An(i_12_), .B(i_3_), .Y(new_new_n210_));
  NO2        g0188(.A(new_new_n44_), .B(i_5_), .Y(new_new_n211_));
  NO3        g0189(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n212_));
  NA3        g0190(.A(new_new_n212_), .B(new_new_n211_), .C(i_10_), .Y(new_new_n213_));
  OAI220     g0191(.A0(new_new_n213_), .A1(new_new_n209_), .B0(new_new_n103_), .B1(new_new_n207_), .Y(new_new_n214_));
  AOI210     g0192(.A0(new_new_n214_), .A1(i_7_), .B0(new_new_n204_), .Y(new_new_n215_));
  OAI220     g0193(.A0(new_new_n215_), .A1(i_4_), .B0(new_new_n197_), .B1(new_new_n195_), .Y(new_new_n216_));
  NAi21      g0194(.An(i_12_), .B(i_7_), .Y(new_new_n217_));
  NA3        g0195(.A(i_13_), .B(new_new_n196_), .C(i_10_), .Y(new_new_n218_));
  NO2        g0196(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n219_));
  NA2        g0197(.A(i_0_), .B(i_5_), .Y(new_new_n220_));
  NA2        g0198(.A(new_new_n220_), .B(new_new_n104_), .Y(new_new_n221_));
  OAI220     g0199(.A0(new_new_n221_), .A1(new_new_n192_), .B0(new_new_n182_), .B1(new_new_n133_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n36_), .B(i_13_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n225_));
  NA3        g0203(.A(new_new_n225_), .B(new_new_n224_), .C(new_new_n223_), .Y(new_new_n226_));
  INV        g0204(.A(i_13_), .Y(new_new_n227_));
  NO2        g0205(.A(i_12_), .B(new_new_n227_), .Y(new_new_n228_));
  NA3        g0206(.A(new_new_n228_), .B(new_new_n200_), .C(new_new_n198_), .Y(new_new_n229_));
  OAI210     g0207(.A0(new_new_n226_), .A1(i_9_), .B0(new_new_n229_), .Y(new_new_n230_));
  AOI220     g0208(.A0(new_new_n230_), .A1(new_new_n142_), .B0(new_new_n222_), .B1(new_new_n219_), .Y(new_new_n231_));
  NO2        g0209(.A(i_12_), .B(new_new_n37_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n185_), .B(i_4_), .Y(new_new_n233_));
  NA2        g0211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  OR2        g0212(.A(i_8_), .B(i_7_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n235_), .B(new_new_n85_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n53_), .B(i_1_), .Y(new_new_n237_));
  NA2        g0215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  INV        g0216(.A(i_12_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n44_), .B(new_new_n239_), .Y(new_new_n240_));
  NO3        g0218(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n241_));
  NA2        g0219(.A(i_2_), .B(i_1_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n238_), .B(new_new_n234_), .Y(new_new_n243_));
  NO3        g0221(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n244_));
  NAi21      g0222(.An(i_4_), .B(i_3_), .Y(new_new_n245_));
  INV        g0223(.A(new_new_n75_), .Y(new_new_n246_));
  NO2        g0224(.A(i_0_), .B(i_6_), .Y(new_new_n247_));
  NOi41      g0225(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n248_));
  NA2        g0226(.A(new_new_n248_), .B(new_new_n247_), .Y(new_new_n249_));
  NO2        g0227(.A(new_new_n242_), .B(new_new_n185_), .Y(new_new_n250_));
  NAi21      g0228(.An(new_new_n249_), .B(new_new_n250_), .Y(new_new_n251_));
  INV        g0229(.A(new_new_n251_), .Y(new_new_n252_));
  AOI220     g0230(.A0(new_new_n252_), .A1(new_new_n40_), .B0(new_new_n243_), .B1(new_new_n208_), .Y(new_new_n253_));
  NO2        g0231(.A(i_11_), .B(new_new_n227_), .Y(new_new_n254_));
  NOi21      g0232(.An(i_1_), .B(i_6_), .Y(new_new_n255_));
  NAi21      g0233(.An(i_3_), .B(i_7_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n239_), .B(i_9_), .Y(new_new_n257_));
  OR4        g0235(.A(new_new_n257_), .B(new_new_n256_), .C(new_new_n255_), .D(new_new_n188_), .Y(new_new_n258_));
  NO2        g0236(.A(i_12_), .B(i_3_), .Y(new_new_n259_));
  NA2        g0237(.A(new_new_n73_), .B(i_5_), .Y(new_new_n260_));
  NA2        g0238(.A(i_3_), .B(i_9_), .Y(new_new_n261_));
  NAi21      g0239(.An(i_7_), .B(i_10_), .Y(new_new_n262_));
  NO2        g0240(.A(new_new_n262_), .B(new_new_n261_), .Y(new_new_n263_));
  NA3        g0241(.A(new_new_n263_), .B(new_new_n260_), .C(new_new_n64_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n264_), .B(new_new_n258_), .Y(new_new_n265_));
  NA3        g0243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n266_));
  INV        g0244(.A(new_new_n143_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n239_), .B(i_13_), .Y(new_new_n268_));
  NO2        g0246(.A(new_new_n268_), .B(new_new_n75_), .Y(new_new_n269_));
  AOI220     g0247(.A0(new_new_n269_), .A1(new_new_n267_), .B0(new_new_n265_), .B1(new_new_n254_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n235_), .B(new_new_n37_), .Y(new_new_n271_));
  NA2        g0249(.A(i_12_), .B(i_6_), .Y(new_new_n272_));
  OR2        g0250(.A(i_13_), .B(i_9_), .Y(new_new_n273_));
  NO3        g0251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n48_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n245_), .B(i_2_), .Y(new_new_n275_));
  NA3        g0253(.A(new_new_n275_), .B(new_new_n274_), .C(new_new_n44_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n254_), .B(i_9_), .Y(new_new_n277_));
  NA2        g0255(.A(new_new_n260_), .B(new_new_n64_), .Y(new_new_n278_));
  OAI210     g0256(.A0(new_new_n278_), .A1(new_new_n277_), .B0(new_new_n276_), .Y(new_new_n279_));
  NA2        g0257(.A(new_new_n155_), .B(new_new_n63_), .Y(new_new_n280_));
  NO3        g0258(.A(i_11_), .B(new_new_n227_), .C(new_new_n25_), .Y(new_new_n281_));
  NO2        g0259(.A(new_new_n256_), .B(i_8_), .Y(new_new_n282_));
  NO2        g0260(.A(i_6_), .B(new_new_n48_), .Y(new_new_n283_));
  NA3        g0261(.A(new_new_n283_), .B(new_new_n282_), .C(new_new_n281_), .Y(new_new_n284_));
  NO3        g0262(.A(new_new_n26_), .B(new_new_n85_), .C(i_5_), .Y(new_new_n285_));
  NA3        g0263(.A(new_new_n285_), .B(new_new_n271_), .C(new_new_n228_), .Y(new_new_n286_));
  AOI210     g0264(.A0(new_new_n286_), .A1(new_new_n284_), .B0(new_new_n280_), .Y(new_new_n287_));
  AOI210     g0265(.A0(new_new_n279_), .A1(new_new_n271_), .B0(new_new_n287_), .Y(new_new_n288_));
  NA4        g0266(.A(new_new_n288_), .B(new_new_n270_), .C(new_new_n253_), .D(new_new_n231_), .Y(new_new_n289_));
  NO3        g0267(.A(i_12_), .B(new_new_n227_), .C(new_new_n37_), .Y(new_new_n290_));
  INV        g0268(.A(new_new_n290_), .Y(new_new_n291_));
  NA2        g0269(.A(i_8_), .B(new_new_n101_), .Y(new_new_n292_));
  NO3        g0270(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n293_));
  AOI220     g0271(.A0(new_new_n293_), .A1(new_new_n198_), .B0(new_new_n164_), .B1(new_new_n237_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n294_), .B(new_new_n292_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n242_), .B(i_0_), .Y(new_new_n296_));
  AOI220     g0274(.A0(new_new_n296_), .A1(i_8_), .B0(i_1_), .B1(new_new_n142_), .Y(new_new_n297_));
  NA2        g0275(.A(new_new_n283_), .B(new_new_n26_), .Y(new_new_n298_));
  NO2        g0276(.A(new_new_n298_), .B(new_new_n297_), .Y(new_new_n299_));
  NA2        g0277(.A(i_0_), .B(i_1_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n300_), .B(i_2_), .Y(new_new_n301_));
  NO2        g0279(.A(new_new_n59_), .B(i_6_), .Y(new_new_n302_));
  NA3        g0280(.A(new_new_n302_), .B(new_new_n301_), .C(new_new_n164_), .Y(new_new_n303_));
  INV        g0281(.A(new_new_n303_), .Y(new_new_n304_));
  NO3        g0282(.A(new_new_n304_), .B(new_new_n299_), .C(new_new_n295_), .Y(new_new_n305_));
  NO2        g0283(.A(i_3_), .B(i_10_), .Y(new_new_n306_));
  NA3        g0284(.A(new_new_n306_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n307_));
  NO2        g0285(.A(i_2_), .B(new_new_n101_), .Y(new_new_n308_));
  NA2        g0286(.A(i_1_), .B(new_new_n36_), .Y(new_new_n309_));
  NOi21      g0287(.An(new_new_n220_), .B(new_new_n103_), .Y(new_new_n310_));
  NA3        g0288(.A(new_new_n310_), .B(new_new_n36_), .C(new_new_n308_), .Y(new_new_n311_));
  AN2        g0289(.A(i_3_), .B(i_10_), .Y(new_new_n312_));
  NA4        g0290(.A(new_new_n312_), .B(new_new_n200_), .C(new_new_n178_), .D(new_new_n176_), .Y(new_new_n313_));
  NO2        g0291(.A(i_5_), .B(new_new_n37_), .Y(new_new_n314_));
  NO2        g0292(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n315_));
  OR2        g0293(.A(new_new_n311_), .B(new_new_n307_), .Y(new_new_n316_));
  OAI220     g0294(.A0(new_new_n316_), .A1(i_6_), .B0(new_new_n305_), .B1(new_new_n291_), .Y(new_new_n317_));
  NO4        g0295(.A(new_new_n317_), .B(new_new_n289_), .C(new_new_n216_), .D(new_new_n169_), .Y(new_new_n318_));
  NO3        g0296(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n319_));
  NO2        g0297(.A(new_new_n59_), .B(new_new_n85_), .Y(new_new_n320_));
  NA2        g0298(.A(new_new_n296_), .B(new_new_n320_), .Y(new_new_n321_));
  NO3        g0299(.A(i_6_), .B(new_new_n196_), .C(i_7_), .Y(new_new_n322_));
  NA2        g0300(.A(new_new_n322_), .B(new_new_n200_), .Y(new_new_n323_));
  AOI210     g0301(.A0(new_new_n323_), .A1(new_new_n321_), .B0(new_new_n171_), .Y(new_new_n324_));
  NO2        g0302(.A(i_2_), .B(i_3_), .Y(new_new_n325_));
  OR2        g0303(.A(i_0_), .B(i_5_), .Y(new_new_n326_));
  NA2        g0304(.A(new_new_n220_), .B(new_new_n326_), .Y(new_new_n327_));
  NA4        g0305(.A(new_new_n327_), .B(new_new_n236_), .C(new_new_n325_), .D(i_1_), .Y(new_new_n328_));
  NA3        g0306(.A(new_new_n296_), .B(new_new_n164_), .C(new_new_n112_), .Y(new_new_n329_));
  NAi21      g0307(.An(i_8_), .B(i_7_), .Y(new_new_n330_));
  NO2        g0308(.A(new_new_n330_), .B(i_6_), .Y(new_new_n331_));
  NO2        g0309(.A(new_new_n158_), .B(new_new_n46_), .Y(new_new_n332_));
  NA3        g0310(.A(new_new_n332_), .B(new_new_n331_), .C(new_new_n164_), .Y(new_new_n333_));
  NA3        g0311(.A(new_new_n333_), .B(new_new_n329_), .C(new_new_n328_), .Y(new_new_n334_));
  OAI210     g0312(.A0(new_new_n334_), .A1(new_new_n324_), .B0(i_4_), .Y(new_new_n335_));
  NO2        g0313(.A(i_12_), .B(i_10_), .Y(new_new_n336_));
  NOi21      g0314(.An(i_5_), .B(i_0_), .Y(new_new_n337_));
  NO2        g0315(.A(new_new_n309_), .B(new_new_n128_), .Y(new_new_n338_));
  NA2        g0316(.A(new_new_n338_), .B(new_new_n336_), .Y(new_new_n339_));
  NO2        g0317(.A(i_6_), .B(i_8_), .Y(new_new_n340_));
  NOi21      g0318(.An(i_0_), .B(i_2_), .Y(new_new_n341_));
  AN2        g0319(.A(new_new_n341_), .B(new_new_n340_), .Y(new_new_n342_));
  NO2        g0320(.A(i_1_), .B(i_7_), .Y(new_new_n343_));
  AO220      g0321(.A0(new_new_n343_), .A1(new_new_n342_), .B0(new_new_n331_), .B1(new_new_n237_), .Y(new_new_n344_));
  NA2        g0322(.A(new_new_n344_), .B(i_4_), .Y(new_new_n345_));
  NA3        g0323(.A(new_new_n345_), .B(new_new_n339_), .C(new_new_n335_), .Y(new_new_n346_));
  NO3        g0324(.A(new_new_n235_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n347_));
  NO3        g0325(.A(new_new_n330_), .B(i_2_), .C(i_1_), .Y(new_new_n348_));
  OAI210     g0326(.A0(new_new_n348_), .A1(new_new_n347_), .B0(i_6_), .Y(new_new_n349_));
  NA2        g0327(.A(new_new_n255_), .B(new_new_n308_), .Y(new_new_n350_));
  AOI210     g0328(.A0(new_new_n350_), .A1(new_new_n349_), .B0(new_new_n327_), .Y(new_new_n351_));
  NOi21      g0329(.An(new_new_n154_), .B(new_new_n104_), .Y(new_new_n352_));
  NO2        g0330(.A(new_new_n352_), .B(new_new_n124_), .Y(new_new_n353_));
  OAI210     g0331(.A0(new_new_n353_), .A1(new_new_n351_), .B0(i_3_), .Y(new_new_n354_));
  INV        g0332(.A(new_new_n83_), .Y(new_new_n355_));
  NO2        g0333(.A(new_new_n300_), .B(new_new_n81_), .Y(new_new_n356_));
  NA2        g0334(.A(new_new_n356_), .B(new_new_n132_), .Y(new_new_n357_));
  NO2        g0335(.A(new_new_n92_), .B(new_new_n196_), .Y(new_new_n358_));
  NA3        g0336(.A(new_new_n310_), .B(new_new_n358_), .C(new_new_n63_), .Y(new_new_n359_));
  AOI210     g0337(.A0(new_new_n359_), .A1(new_new_n357_), .B0(new_new_n355_), .Y(new_new_n360_));
  NO2        g0338(.A(new_new_n196_), .B(i_9_), .Y(new_new_n361_));
  NO2        g0339(.A(new_new_n360_), .B(new_new_n299_), .Y(new_new_n362_));
  AOI210     g0340(.A0(new_new_n362_), .A1(new_new_n354_), .B0(new_new_n163_), .Y(new_new_n363_));
  AOI210     g0341(.A0(new_new_n346_), .A1(new_new_n319_), .B0(new_new_n363_), .Y(new_new_n364_));
  NOi32      g0342(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n365_));
  INV        g0343(.A(new_new_n365_), .Y(new_new_n366_));
  NAi21      g0344(.An(i_0_), .B(i_6_), .Y(new_new_n367_));
  NAi21      g0345(.An(i_1_), .B(i_5_), .Y(new_new_n368_));
  NA2        g0346(.A(new_new_n368_), .B(new_new_n367_), .Y(new_new_n369_));
  NA2        g0347(.A(new_new_n369_), .B(new_new_n25_), .Y(new_new_n370_));
  OAI210     g0348(.A0(new_new_n370_), .A1(new_new_n160_), .B0(new_new_n249_), .Y(new_new_n371_));
  NAi41      g0349(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n372_));
  AOI210     g0350(.A0(new_new_n372_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n373_));
  NOi32      g0351(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n374_));
  NO2        g0352(.A(i_1_), .B(new_new_n101_), .Y(new_new_n375_));
  NAi21      g0353(.An(i_3_), .B(i_4_), .Y(new_new_n376_));
  NO2        g0354(.A(new_new_n376_), .B(i_9_), .Y(new_new_n377_));
  AN2        g0355(.A(i_6_), .B(i_7_), .Y(new_new_n378_));
  OAI210     g0356(.A0(new_new_n378_), .A1(new_new_n375_), .B0(new_new_n377_), .Y(new_new_n379_));
  NA2        g0357(.A(i_2_), .B(i_7_), .Y(new_new_n380_));
  NO2        g0358(.A(new_new_n376_), .B(i_10_), .Y(new_new_n381_));
  NA3        g0359(.A(new_new_n381_), .B(new_new_n380_), .C(new_new_n247_), .Y(new_new_n382_));
  AOI210     g0360(.A0(new_new_n382_), .A1(new_new_n379_), .B0(new_new_n188_), .Y(new_new_n383_));
  AOI210     g0361(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n384_));
  AOI220     g0362(.A0(new_new_n381_), .A1(new_new_n343_), .B0(new_new_n241_), .B1(new_new_n191_), .Y(new_new_n385_));
  NO3        g0363(.A(new_new_n383_), .B(new_new_n373_), .C(new_new_n371_), .Y(new_new_n386_));
  NO2        g0364(.A(new_new_n386_), .B(new_new_n366_), .Y(new_new_n387_));
  NO2        g0365(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n388_));
  AN2        g0366(.A(i_12_), .B(i_5_), .Y(new_new_n389_));
  NO2        g0367(.A(i_4_), .B(new_new_n26_), .Y(new_new_n390_));
  NA2        g0368(.A(new_new_n390_), .B(new_new_n389_), .Y(new_new_n391_));
  NO2        g0369(.A(i_11_), .B(i_6_), .Y(new_new_n392_));
  NA3        g0370(.A(new_new_n392_), .B(new_new_n332_), .C(new_new_n227_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n393_), .B(new_new_n391_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n245_), .B(i_5_), .Y(new_new_n395_));
  NO2        g0373(.A(i_5_), .B(i_10_), .Y(new_new_n396_));
  NA2        g0374(.A(new_new_n395_), .B(new_new_n200_), .Y(new_new_n397_));
  NO2        g0375(.A(i_12_), .B(new_new_n397_), .Y(new_new_n398_));
  OAI210     g0376(.A0(new_new_n398_), .A1(new_new_n394_), .B0(new_new_n388_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n400_));
  INV        g0378(.A(new_new_n150_), .Y(new_new_n401_));
  OAI210     g0379(.A0(new_new_n401_), .A1(new_new_n394_), .B0(new_new_n400_), .Y(new_new_n402_));
  NO3        g0380(.A(new_new_n85_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n403_));
  NA2        g0381(.A(new_new_n306_), .B(new_new_n90_), .Y(new_new_n404_));
  NO2        g0382(.A(i_11_), .B(i_12_), .Y(new_new_n405_));
  NA2        g0383(.A(new_new_n405_), .B(new_new_n36_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n404_), .B(new_new_n406_), .Y(new_new_n407_));
  NA2        g0385(.A(new_new_n396_), .B(new_new_n239_), .Y(new_new_n408_));
  NA3        g0386(.A(new_new_n112_), .B(i_4_), .C(i_11_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n409_), .B(i_9_), .Y(new_new_n410_));
  NAi21      g0388(.An(i_13_), .B(i_0_), .Y(new_new_n411_));
  NO2        g0389(.A(new_new_n411_), .B(new_new_n242_), .Y(new_new_n412_));
  OAI210     g0390(.A0(new_new_n410_), .A1(new_new_n407_), .B0(new_new_n412_), .Y(new_new_n413_));
  NA3        g0391(.A(new_new_n413_), .B(new_new_n402_), .C(new_new_n399_), .Y(new_new_n414_));
  NO2        g0392(.A(i_0_), .B(i_11_), .Y(new_new_n415_));
  INV        g0393(.A(i_5_), .Y(new_new_n416_));
  AN2        g0394(.A(i_1_), .B(i_6_), .Y(new_new_n417_));
  NOi21      g0395(.An(i_2_), .B(i_12_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n418_), .B(new_new_n417_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n419_), .B(new_new_n416_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n142_), .B(i_9_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n421_), .B(i_4_), .Y(new_new_n422_));
  NA2        g0400(.A(new_new_n420_), .B(new_new_n422_), .Y(new_new_n423_));
  NAi21      g0401(.An(i_9_), .B(i_4_), .Y(new_new_n424_));
  OR2        g0402(.A(i_13_), .B(i_10_), .Y(new_new_n425_));
  NO3        g0403(.A(new_new_n425_), .B(new_new_n117_), .C(new_new_n424_), .Y(new_new_n426_));
  NO2        g0404(.A(new_new_n174_), .B(new_new_n123_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n290_), .B(new_new_n428_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n283_), .B(new_new_n212_), .Y(new_new_n430_));
  OAI220     g0408(.A0(new_new_n430_), .A1(new_new_n218_), .B0(new_new_n429_), .B1(new_new_n352_), .Y(new_new_n431_));
  INV        g0409(.A(new_new_n431_), .Y(new_new_n432_));
  AOI210     g0410(.A0(new_new_n432_), .A1(new_new_n423_), .B0(new_new_n26_), .Y(new_new_n433_));
  NA2        g0411(.A(new_new_n329_), .B(new_new_n328_), .Y(new_new_n434_));
  AOI220     g0412(.A0(new_new_n302_), .A1(new_new_n293_), .B0(new_new_n296_), .B1(new_new_n320_), .Y(new_new_n435_));
  NO2        g0413(.A(new_new_n435_), .B(new_new_n171_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n185_), .B(new_new_n85_), .Y(new_new_n437_));
  AOI220     g0415(.A0(new_new_n437_), .A1(new_new_n301_), .B0(new_new_n285_), .B1(new_new_n212_), .Y(new_new_n438_));
  NO2        g0416(.A(new_new_n438_), .B(new_new_n292_), .Y(new_new_n439_));
  NO3        g0417(.A(new_new_n439_), .B(new_new_n436_), .C(new_new_n434_), .Y(new_new_n440_));
  NA2        g0418(.A(new_new_n198_), .B(new_new_n96_), .Y(new_new_n441_));
  NA3        g0419(.A(new_new_n332_), .B(new_new_n164_), .C(new_new_n85_), .Y(new_new_n442_));
  AOI210     g0420(.A0(new_new_n442_), .A1(new_new_n441_), .B0(new_new_n330_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n302_), .B(new_new_n237_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n444_), .B(new_new_n185_), .Y(new_new_n445_));
  NO2        g0423(.A(i_3_), .B(new_new_n48_), .Y(new_new_n446_));
  NO2        g0424(.A(new_new_n445_), .B(new_new_n443_), .Y(new_new_n447_));
  AOI210     g0425(.A0(new_new_n447_), .A1(new_new_n440_), .B0(new_new_n277_), .Y(new_new_n448_));
  NO4        g0426(.A(new_new_n448_), .B(new_new_n433_), .C(new_new_n414_), .D(new_new_n387_), .Y(new_new_n449_));
  NO2        g0427(.A(new_new_n63_), .B(i_4_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n73_), .B(i_13_), .Y(new_new_n451_));
  NO2        g0429(.A(i_10_), .B(i_9_), .Y(new_new_n452_));
  NAi21      g0430(.An(i_12_), .B(i_8_), .Y(new_new_n453_));
  NO2        g0431(.A(new_new_n453_), .B(i_3_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n46_), .B(i_4_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n455_), .B(new_new_n104_), .Y(new_new_n456_));
  NO2        g0434(.A(new_new_n456_), .B(new_new_n207_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n315_), .B(i_0_), .Y(new_new_n458_));
  NO3        g0436(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n272_), .B(new_new_n97_), .Y(new_new_n460_));
  NA2        g0438(.A(new_new_n460_), .B(new_new_n459_), .Y(new_new_n461_));
  NA2        g0439(.A(i_8_), .B(i_9_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n461_), .B(new_new_n458_), .Y(new_new_n463_));
  NO3        g0441(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n464_));
  NA3        g0442(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n465_));
  NA4        g0443(.A(new_new_n145_), .B(new_new_n115_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n466_));
  NO2        g0444(.A(new_new_n466_), .B(new_new_n465_), .Y(new_new_n467_));
  NO3        g0445(.A(new_new_n467_), .B(new_new_n463_), .C(new_new_n457_), .Y(new_new_n468_));
  OR2        g0446(.A(new_new_n300_), .B(new_new_n209_), .Y(new_new_n469_));
  BUFFER     g0447(.A(new_new_n303_), .Y(new_new_n470_));
  OA220      g0448(.A0(new_new_n470_), .A1(new_new_n163_), .B0(new_new_n469_), .B1(new_new_n234_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n96_), .B(i_13_), .Y(new_new_n472_));
  NA2        g0450(.A(new_new_n437_), .B(new_new_n388_), .Y(new_new_n473_));
  NO2        g0451(.A(new_new_n473_), .B(new_new_n472_), .Y(new_new_n474_));
  NO3        g0452(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n475_));
  NO2        g0453(.A(i_6_), .B(i_7_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n476_), .B(new_new_n475_), .Y(new_new_n477_));
  NO2        g0455(.A(i_11_), .B(i_1_), .Y(new_new_n478_));
  NO2        g0456(.A(new_new_n73_), .B(i_3_), .Y(new_new_n479_));
  NOi21      g0457(.An(i_2_), .B(i_7_), .Y(new_new_n480_));
  NAi31      g0458(.An(i_11_), .B(new_new_n480_), .C(new_new_n479_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n425_), .B(i_6_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n482_), .B(new_new_n450_), .Y(new_new_n483_));
  NO2        g0461(.A(new_new_n483_), .B(new_new_n481_), .Y(new_new_n484_));
  NO2        g0462(.A(i_6_), .B(i_10_), .Y(new_new_n485_));
  NA4        g0463(.A(new_new_n485_), .B(new_new_n319_), .C(i_8_), .D(new_new_n239_), .Y(new_new_n486_));
  NO2        g0464(.A(new_new_n486_), .B(new_new_n156_), .Y(new_new_n487_));
  NA2        g0465(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n488_));
  NO2        g0466(.A(new_new_n158_), .B(i_3_), .Y(new_new_n489_));
  NAi31      g0467(.An(new_new_n488_), .B(new_new_n489_), .C(new_new_n228_), .Y(new_new_n490_));
  NA3        g0468(.A(new_new_n400_), .B(new_new_n181_), .C(new_new_n149_), .Y(new_new_n491_));
  NA2        g0469(.A(new_new_n491_), .B(new_new_n490_), .Y(new_new_n492_));
  NO4        g0470(.A(new_new_n492_), .B(new_new_n487_), .C(new_new_n484_), .D(new_new_n474_), .Y(new_new_n493_));
  NA2        g0471(.A(new_new_n464_), .B(new_new_n396_), .Y(new_new_n494_));
  NO2        g0472(.A(new_new_n494_), .B(new_new_n226_), .Y(new_new_n495_));
  NAi21      g0473(.An(new_new_n218_), .B(new_new_n405_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n343_), .B(new_new_n220_), .Y(new_new_n497_));
  NO2        g0475(.A(new_new_n26_), .B(i_5_), .Y(new_new_n498_));
  NO2        g0476(.A(i_0_), .B(new_new_n85_), .Y(new_new_n499_));
  NA3        g0477(.A(new_new_n499_), .B(new_new_n498_), .C(new_new_n142_), .Y(new_new_n500_));
  OR3        g0478(.A(new_new_n309_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n501_));
  OAI220     g0479(.A0(new_new_n501_), .A1(new_new_n500_), .B0(new_new_n497_), .B1(new_new_n496_), .Y(new_new_n502_));
  NA2        g0480(.A(new_new_n27_), .B(i_10_), .Y(new_new_n503_));
  NO2        g0481(.A(new_new_n503_), .B(new_new_n472_), .Y(new_new_n504_));
  NA3        g0482(.A(new_new_n312_), .B(new_new_n225_), .C(new_new_n73_), .Y(new_new_n505_));
  NO2        g0483(.A(new_new_n505_), .B(new_new_n477_), .Y(new_new_n506_));
  NO4        g0484(.A(new_new_n506_), .B(new_new_n504_), .C(new_new_n502_), .D(new_new_n495_), .Y(new_new_n507_));
  NA4        g0485(.A(new_new_n507_), .B(new_new_n493_), .C(new_new_n471_), .D(new_new_n468_), .Y(new_new_n508_));
  NA3        g0486(.A(new_new_n312_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n509_));
  INV        g0487(.A(new_new_n509_), .Y(new_new_n510_));
  AN2        g0488(.A(new_new_n293_), .B(new_new_n236_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n511_), .B(new_new_n510_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n122_), .B(new_new_n111_), .Y(new_new_n513_));
  AN2        g0491(.A(new_new_n513_), .B(new_new_n459_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n319_), .B(new_new_n165_), .Y(new_new_n515_));
  OAI210     g0493(.A0(new_new_n515_), .A1(new_new_n234_), .B0(new_new_n313_), .Y(new_new_n516_));
  AOI220     g0494(.A0(new_new_n516_), .A1(new_new_n331_), .B0(new_new_n514_), .B1(new_new_n315_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n389_), .B(new_new_n227_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n365_), .B(new_new_n73_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n378_), .B(new_new_n374_), .Y(new_new_n520_));
  AO210      g0498(.A0(new_new_n519_), .A1(new_new_n518_), .B0(new_new_n520_), .Y(new_new_n521_));
  NO2        g0499(.A(new_new_n36_), .B(i_8_), .Y(new_new_n522_));
  NAi41      g0500(.An(new_new_n519_), .B(new_new_n485_), .C(new_new_n522_), .D(new_new_n46_), .Y(new_new_n523_));
  AOI210     g0501(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n426_), .Y(new_new_n524_));
  NA3        g0502(.A(new_new_n524_), .B(new_new_n523_), .C(new_new_n521_), .Y(new_new_n525_));
  INV        g0503(.A(new_new_n525_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n260_), .B(new_new_n64_), .Y(new_new_n527_));
  OAI210     g0505(.A0(i_8_), .A1(new_new_n527_), .B0(new_new_n134_), .Y(new_new_n528_));
  NO2        g0506(.A(i_7_), .B(new_new_n201_), .Y(new_new_n529_));
  OR2        g0507(.A(new_new_n185_), .B(i_4_), .Y(new_new_n530_));
  NO2        g0508(.A(new_new_n530_), .B(new_new_n85_), .Y(new_new_n531_));
  AOI220     g0509(.A0(new_new_n531_), .A1(new_new_n529_), .B0(new_new_n528_), .B1(new_new_n427_), .Y(new_new_n532_));
  NA4        g0510(.A(new_new_n532_), .B(new_new_n526_), .C(new_new_n517_), .D(new_new_n512_), .Y(new_new_n533_));
  NA2        g0511(.A(new_new_n395_), .B(new_new_n301_), .Y(new_new_n534_));
  OAI210     g0512(.A0(new_new_n391_), .A1(new_new_n170_), .B0(new_new_n534_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n1041_), .B(new_new_n227_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n485_), .B(new_new_n27_), .Y(new_new_n537_));
  NO2        g0515(.A(new_new_n537_), .B(new_new_n536_), .Y(new_new_n538_));
  NOi31      g0516(.An(new_new_n322_), .B(new_new_n425_), .C(new_new_n38_), .Y(new_new_n539_));
  OAI210     g0517(.A0(new_new_n539_), .A1(new_new_n538_), .B0(new_new_n535_), .Y(new_new_n540_));
  NO2        g0518(.A(i_8_), .B(i_7_), .Y(new_new_n541_));
  OAI210     g0519(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n542_));
  NA2        g0520(.A(new_new_n542_), .B(new_new_n225_), .Y(new_new_n543_));
  OAI220     g0521(.A0(new_new_n46_), .A1(new_new_n530_), .B0(new_new_n543_), .B1(new_new_n245_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n44_), .B(i_10_), .Y(new_new_n545_));
  NO2        g0523(.A(new_new_n545_), .B(i_6_), .Y(new_new_n546_));
  NA3        g0524(.A(new_new_n546_), .B(new_new_n544_), .C(new_new_n541_), .Y(new_new_n547_));
  AOI220     g0525(.A0(new_new_n437_), .A1(new_new_n332_), .B0(new_new_n250_), .B1(new_new_n247_), .Y(new_new_n548_));
  NO2        g0526(.A(new_new_n548_), .B(new_new_n268_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n549_), .B(new_new_n271_), .Y(new_new_n550_));
  NO2        g0528(.A(new_new_n307_), .B(new_new_n183_), .Y(new_new_n551_));
  NA3        g0529(.A(new_new_n312_), .B(new_new_n176_), .C(new_new_n96_), .Y(new_new_n552_));
  NO2        g0530(.A(new_new_n223_), .B(new_new_n44_), .Y(new_new_n553_));
  NO2        g0531(.A(new_new_n158_), .B(i_5_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n554_), .B(new_new_n325_), .Y(new_new_n555_));
  OAI210     g0533(.A0(new_new_n555_), .A1(new_new_n553_), .B0(new_new_n552_), .Y(new_new_n556_));
  OAI210     g0534(.A0(new_new_n556_), .A1(new_new_n551_), .B0(new_new_n464_), .Y(new_new_n557_));
  NA4        g0535(.A(new_new_n557_), .B(new_new_n550_), .C(new_new_n547_), .D(new_new_n540_), .Y(new_new_n558_));
  NA3        g0536(.A(new_new_n220_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n559_));
  NA2        g0537(.A(new_new_n290_), .B(new_new_n83_), .Y(new_new_n560_));
  AOI210     g0538(.A0(new_new_n559_), .A1(new_new_n357_), .B0(new_new_n560_), .Y(new_new_n561_));
  NA2        g0539(.A(new_new_n302_), .B(new_new_n293_), .Y(new_new_n562_));
  NO2        g0540(.A(new_new_n562_), .B(new_new_n175_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n564_));
  NA2        g0542(.A(new_new_n452_), .B(new_new_n223_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n564_), .B(new_new_n565_), .Y(new_new_n566_));
  NA2        g0544(.A(i_0_), .B(new_new_n48_), .Y(new_new_n567_));
  NO3        g0545(.A(new_new_n566_), .B(new_new_n563_), .C(new_new_n561_), .Y(new_new_n568_));
  NO4        g0546(.A(new_new_n255_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n569_));
  NO3        g0547(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n570_));
  NO2        g0548(.A(new_new_n235_), .B(new_new_n36_), .Y(new_new_n571_));
  AN2        g0549(.A(new_new_n571_), .B(new_new_n570_), .Y(new_new_n572_));
  OA210      g0550(.A0(new_new_n572_), .A1(new_new_n569_), .B0(new_new_n365_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n425_), .B(i_1_), .Y(new_new_n574_));
  NOi31      g0552(.An(new_new_n574_), .B(new_new_n460_), .C(new_new_n73_), .Y(new_new_n575_));
  AN4        g0553(.A(new_new_n575_), .B(new_new_n422_), .C(new_new_n498_), .D(i_2_), .Y(new_new_n576_));
  NO2        g0554(.A(new_new_n435_), .B(new_new_n179_), .Y(new_new_n577_));
  NO3        g0555(.A(new_new_n577_), .B(new_new_n576_), .C(new_new_n573_), .Y(new_new_n578_));
  NOi21      g0556(.An(i_10_), .B(i_6_), .Y(new_new_n579_));
  NO2        g0557(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n580_));
  AOI220     g0558(.A0(new_new_n290_), .A1(new_new_n580_), .B0(new_new_n281_), .B1(new_new_n579_), .Y(new_new_n581_));
  NO2        g0559(.A(new_new_n581_), .B(new_new_n458_), .Y(new_new_n582_));
  NO2        g0560(.A(new_new_n114_), .B(new_new_n23_), .Y(new_new_n583_));
  NA2        g0561(.A(new_new_n322_), .B(new_new_n165_), .Y(new_new_n584_));
  AOI220     g0562(.A0(new_new_n584_), .A1(new_new_n444_), .B0(new_new_n186_), .B1(new_new_n184_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n585_), .B(new_new_n582_), .Y(new_new_n586_));
  NO2        g0564(.A(new_new_n519_), .B(new_new_n385_), .Y(new_new_n587_));
  INV        g0565(.A(new_new_n325_), .Y(new_new_n588_));
  NO2        g0566(.A(i_12_), .B(new_new_n85_), .Y(new_new_n589_));
  NO3        g0567(.A(i_4_), .B(new_new_n349_), .C(new_new_n307_), .Y(new_new_n590_));
  OR2        g0568(.A(i_2_), .B(i_5_), .Y(new_new_n591_));
  OR2        g0569(.A(new_new_n591_), .B(new_new_n417_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n592_), .B(new_new_n496_), .Y(new_new_n593_));
  NO3        g0571(.A(new_new_n593_), .B(new_new_n590_), .C(new_new_n587_), .Y(new_new_n594_));
  NA4        g0572(.A(new_new_n594_), .B(new_new_n586_), .C(new_new_n578_), .D(new_new_n568_), .Y(new_new_n595_));
  NO4        g0573(.A(new_new_n595_), .B(new_new_n558_), .C(new_new_n533_), .D(new_new_n508_), .Y(new_new_n596_));
  NA4        g0574(.A(new_new_n596_), .B(new_new_n449_), .C(new_new_n364_), .D(new_new_n318_), .Y(men7));
  NO2        g0575(.A(new_new_n92_), .B(new_new_n54_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n108_), .B(new_new_n89_), .Y(new_new_n599_));
  NA2        g0577(.A(i_11_), .B(new_new_n196_), .Y(new_new_n600_));
  NA3        g0578(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n601_));
  NO2        g0579(.A(new_new_n239_), .B(i_4_), .Y(new_new_n602_));
  NA2        g0580(.A(new_new_n602_), .B(i_8_), .Y(new_new_n603_));
  NO2        g0581(.A(new_new_n105_), .B(new_new_n601_), .Y(new_new_n604_));
  NA2        g0582(.A(i_2_), .B(new_new_n85_), .Y(new_new_n605_));
  OAI210     g0583(.A0(new_new_n86_), .A1(new_new_n205_), .B0(new_new_n206_), .Y(new_new_n606_));
  NO2        g0584(.A(i_7_), .B(new_new_n37_), .Y(new_new_n607_));
  NA2        g0585(.A(i_4_), .B(i_8_), .Y(new_new_n608_));
  AOI210     g0586(.A0(new_new_n608_), .A1(new_new_n312_), .B0(new_new_n607_), .Y(new_new_n609_));
  OAI220     g0587(.A0(new_new_n609_), .A1(new_new_n605_), .B0(new_new_n606_), .B1(i_13_), .Y(new_new_n610_));
  NO3        g0588(.A(new_new_n610_), .B(new_new_n604_), .C(new_new_n598_), .Y(new_new_n611_));
  OR2        g0589(.A(i_6_), .B(i_10_), .Y(new_new_n612_));
  NO2        g0590(.A(new_new_n612_), .B(new_new_n23_), .Y(new_new_n613_));
  OR3        g0591(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n614_));
  NO3        g0592(.A(new_new_n614_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n615_));
  INV        g0593(.A(new_new_n202_), .Y(new_new_n616_));
  NO2        g0594(.A(new_new_n615_), .B(new_new_n613_), .Y(new_new_n617_));
  OA220      g0595(.A0(new_new_n617_), .A1(new_new_n588_), .B0(new_new_n1043_), .B1(new_new_n273_), .Y(new_new_n618_));
  AOI210     g0596(.A0(new_new_n618_), .A1(new_new_n611_), .B0(new_new_n63_), .Y(new_new_n619_));
  NOi21      g0597(.An(i_11_), .B(i_7_), .Y(new_new_n620_));
  AO210      g0598(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n621_));
  NO2        g0599(.A(new_new_n621_), .B(new_new_n620_), .Y(new_new_n622_));
  NA2        g0600(.A(new_new_n622_), .B(new_new_n208_), .Y(new_new_n623_));
  NA3        g0601(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n624_));
  NAi31      g0602(.An(new_new_n624_), .B(new_new_n217_), .C(i_11_), .Y(new_new_n625_));
  AOI210     g0603(.A0(new_new_n625_), .A1(new_new_n623_), .B0(new_new_n63_), .Y(new_new_n626_));
  NO3        g0604(.A(new_new_n262_), .B(new_new_n210_), .C(new_new_n600_), .Y(new_new_n627_));
  OAI210     g0605(.A0(new_new_n627_), .A1(new_new_n228_), .B0(new_new_n63_), .Y(new_new_n628_));
  NA2        g0606(.A(new_new_n418_), .B(new_new_n31_), .Y(new_new_n629_));
  OR2        g0607(.A(new_new_n210_), .B(new_new_n108_), .Y(new_new_n630_));
  NA2        g0608(.A(new_new_n630_), .B(new_new_n629_), .Y(new_new_n631_));
  NO2        g0609(.A(new_new_n63_), .B(i_9_), .Y(new_new_n632_));
  NO2        g0610(.A(new_new_n632_), .B(i_4_), .Y(new_new_n633_));
  NA2        g0611(.A(new_new_n633_), .B(new_new_n631_), .Y(new_new_n634_));
  NO2        g0612(.A(i_1_), .B(i_12_), .Y(new_new_n635_));
  NA2        g0613(.A(new_new_n634_), .B(new_new_n628_), .Y(new_new_n636_));
  OAI210     g0614(.A0(new_new_n636_), .A1(new_new_n626_), .B0(i_6_), .Y(new_new_n637_));
  NO2        g0615(.A(new_new_n239_), .B(new_new_n85_), .Y(new_new_n638_));
  NO2        g0616(.A(new_new_n638_), .B(i_11_), .Y(new_new_n639_));
  INV        g0617(.A(new_new_n461_), .Y(new_new_n640_));
  NO4        g0618(.A(new_new_n217_), .B(new_new_n128_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n641_));
  NA2        g0619(.A(new_new_n641_), .B(new_new_n632_), .Y(new_new_n642_));
  NA2        g0620(.A(new_new_n239_), .B(i_6_), .Y(new_new_n643_));
  NO3        g0621(.A(new_new_n612_), .B(new_new_n235_), .C(new_new_n23_), .Y(new_new_n644_));
  AOI210     g0622(.A0(i_1_), .A1(new_new_n263_), .B0(new_new_n644_), .Y(new_new_n645_));
  OAI210     g0623(.A0(new_new_n645_), .A1(new_new_n44_), .B0(new_new_n642_), .Y(new_new_n646_));
  NA3        g0624(.A(new_new_n541_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n138_), .B(i_9_), .Y(new_new_n648_));
  NA3        g0626(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n649_));
  NO2        g0627(.A(new_new_n46_), .B(i_1_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n648_), .B(new_new_n1040_), .Y(new_new_n651_));
  AOI210     g0629(.A0(new_new_n478_), .A1(new_new_n428_), .B0(new_new_n244_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n652_), .B(new_new_n605_), .Y(new_new_n653_));
  NAi21      g0631(.An(new_new_n647_), .B(new_new_n91_), .Y(new_new_n654_));
  NA2        g0632(.A(new_new_n650_), .B(new_new_n272_), .Y(new_new_n655_));
  NO2        g0633(.A(i_11_), .B(new_new_n37_), .Y(new_new_n656_));
  NA2        g0634(.A(new_new_n656_), .B(new_new_n24_), .Y(new_new_n657_));
  OAI210     g0635(.A0(new_new_n657_), .A1(new_new_n655_), .B0(new_new_n654_), .Y(new_new_n658_));
  OR3        g0636(.A(new_new_n658_), .B(new_new_n653_), .C(new_new_n651_), .Y(new_new_n659_));
  NO3        g0637(.A(new_new_n659_), .B(new_new_n646_), .C(new_new_n640_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n239_), .B(new_new_n101_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n661_), .B(new_new_n620_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(i_1_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n663_), .B(new_new_n614_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n424_), .B(new_new_n85_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n664_), .B(new_new_n46_), .Y(new_new_n666_));
  NA2        g0644(.A(i_3_), .B(new_new_n196_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n667_), .B(new_new_n114_), .Y(new_new_n668_));
  AN2        g0646(.A(new_new_n668_), .B(new_new_n546_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n235_), .B(new_new_n44_), .Y(new_new_n670_));
  NO3        g0648(.A(new_new_n670_), .B(new_new_n315_), .C(new_new_n240_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n672_), .B(i_6_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n85_), .B(i_9_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n63_), .Y(new_new_n675_));
  NO2        g0653(.A(new_new_n675_), .B(new_new_n635_), .Y(new_new_n676_));
  NO4        g0654(.A(new_new_n676_), .B(new_new_n673_), .C(new_new_n671_), .D(i_4_), .Y(new_new_n677_));
  NA2        g0655(.A(i_1_), .B(i_3_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n462_), .B(new_new_n92_), .Y(new_new_n679_));
  AOI210     g0657(.A0(new_new_n670_), .A1(new_new_n579_), .B0(new_new_n679_), .Y(new_new_n680_));
  NO2        g0658(.A(new_new_n680_), .B(new_new_n678_), .Y(new_new_n681_));
  NO3        g0659(.A(new_new_n681_), .B(new_new_n677_), .C(new_new_n669_), .Y(new_new_n682_));
  NA4        g0660(.A(new_new_n682_), .B(new_new_n666_), .C(new_new_n660_), .D(new_new_n637_), .Y(new_new_n683_));
  NO3        g0661(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n684_));
  NOi21      g0662(.An(new_new_n684_), .B(i_10_), .Y(new_new_n685_));
  OA210      g0663(.A0(new_new_n685_), .A1(new_new_n248_), .B0(new_new_n85_), .Y(new_new_n686_));
  NA2        g0664(.A(new_new_n378_), .B(new_new_n377_), .Y(new_new_n687_));
  NA3        g0665(.A(new_new_n485_), .B(new_new_n522_), .C(new_new_n46_), .Y(new_new_n688_));
  NO3        g0666(.A(new_new_n480_), .B(new_new_n608_), .C(new_new_n85_), .Y(new_new_n689_));
  NA2        g0667(.A(new_new_n689_), .B(new_new_n25_), .Y(new_new_n690_));
  NA3        g0668(.A(new_new_n690_), .B(new_new_n688_), .C(new_new_n687_), .Y(new_new_n691_));
  OAI210     g0669(.A0(new_new_n691_), .A1(new_new_n686_), .B0(i_1_), .Y(new_new_n692_));
  AOI210     g0670(.A0(new_new_n272_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n376_), .B(i_2_), .Y(new_new_n694_));
  NA2        g0672(.A(new_new_n694_), .B(new_new_n693_), .Y(new_new_n695_));
  AOI210     g0673(.A0(new_new_n695_), .A1(new_new_n692_), .B0(i_13_), .Y(new_new_n696_));
  OR2        g0674(.A(i_11_), .B(i_7_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n54_), .B(i_12_), .Y(new_new_n698_));
  INV        g0676(.A(new_new_n698_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n480_), .B(new_new_n24_), .Y(new_new_n700_));
  AOI220     g0678(.A0(new_new_n700_), .A1(new_new_n665_), .B0(new_new_n248_), .B1(new_new_n131_), .Y(new_new_n701_));
  OAI220     g0679(.A0(new_new_n701_), .A1(new_new_n41_), .B0(new_new_n699_), .B1(new_new_n92_), .Y(new_new_n702_));
  INV        g0680(.A(new_new_n702_), .Y(new_new_n703_));
  NA2        g0681(.A(new_new_n392_), .B(new_new_n650_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n704_), .B(new_new_n245_), .Y(new_new_n705_));
  AOI210     g0683(.A0(new_new_n453_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n706_));
  NA2        g0684(.A(new_new_n127_), .B(i_13_), .Y(new_new_n707_));
  NO2        g0685(.A(new_new_n649_), .B(new_new_n114_), .Y(new_new_n708_));
  NO2        g0686(.A(new_new_n707_), .B(new_new_n693_), .Y(new_new_n709_));
  NA2        g0687(.A(new_new_n26_), .B(new_new_n196_), .Y(new_new_n710_));
  NA2        g0688(.A(new_new_n710_), .B(i_7_), .Y(new_new_n711_));
  NO3        g0689(.A(new_new_n480_), .B(new_new_n239_), .C(new_new_n85_), .Y(new_new_n712_));
  NA2        g0690(.A(new_new_n712_), .B(new_new_n711_), .Y(new_new_n713_));
  AOI220     g0691(.A0(new_new_n392_), .A1(new_new_n650_), .B0(new_new_n91_), .B1(new_new_n102_), .Y(new_new_n714_));
  OAI220     g0692(.A0(new_new_n714_), .A1(new_new_n603_), .B0(new_new_n713_), .B1(new_new_n616_), .Y(new_new_n715_));
  NO3        g0693(.A(new_new_n715_), .B(new_new_n709_), .C(new_new_n705_), .Y(new_new_n716_));
  OR2        g0694(.A(i_11_), .B(i_6_), .Y(new_new_n717_));
  NA3        g0695(.A(new_new_n418_), .B(new_new_n607_), .C(new_new_n97_), .Y(new_new_n718_));
  NA2        g0696(.A(new_new_n639_), .B(i_13_), .Y(new_new_n719_));
  NAi21      g0697(.An(i_11_), .B(i_12_), .Y(new_new_n720_));
  NA2        g0698(.A(new_new_n719_), .B(new_new_n718_), .Y(new_new_n721_));
  NA2        g0699(.A(new_new_n721_), .B(new_new_n63_), .Y(new_new_n722_));
  NO2        g0700(.A(i_2_), .B(i_12_), .Y(new_new_n723_));
  NA2        g0701(.A(new_new_n375_), .B(new_new_n723_), .Y(new_new_n724_));
  NA2        g0702(.A(i_8_), .B(new_new_n25_), .Y(new_new_n725_));
  NO3        g0703(.A(new_new_n725_), .B(new_new_n390_), .C(new_new_n602_), .Y(new_new_n726_));
  OAI210     g0704(.A0(new_new_n726_), .A1(new_new_n377_), .B0(new_new_n375_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n128_), .B(i_2_), .Y(new_new_n728_));
  NA2        g0706(.A(new_new_n728_), .B(new_new_n635_), .Y(new_new_n729_));
  NA3        g0707(.A(new_new_n729_), .B(new_new_n727_), .C(new_new_n724_), .Y(new_new_n730_));
  NA3        g0708(.A(new_new_n730_), .B(new_new_n45_), .C(new_new_n227_), .Y(new_new_n731_));
  NA4        g0709(.A(new_new_n731_), .B(new_new_n722_), .C(new_new_n716_), .D(new_new_n703_), .Y(new_new_n732_));
  OR4        g0710(.A(new_new_n732_), .B(new_new_n696_), .C(new_new_n683_), .D(new_new_n619_), .Y(men5));
  AOI210     g0711(.A0(new_new_n662_), .A1(new_new_n275_), .B0(new_new_n427_), .Y(new_new_n734_));
  AN2        g0712(.A(new_new_n24_), .B(i_10_), .Y(new_new_n735_));
  NA3        g0713(.A(new_new_n735_), .B(new_new_n723_), .C(new_new_n108_), .Y(new_new_n736_));
  NO2        g0714(.A(new_new_n603_), .B(i_11_), .Y(new_new_n737_));
  NA2        g0715(.A(new_new_n86_), .B(new_new_n737_), .Y(new_new_n738_));
  NA3        g0716(.A(new_new_n738_), .B(new_new_n736_), .C(new_new_n734_), .Y(new_new_n739_));
  NO3        g0717(.A(i_11_), .B(new_new_n239_), .C(i_13_), .Y(new_new_n740_));
  NO2        g0718(.A(new_new_n124_), .B(new_new_n23_), .Y(new_new_n741_));
  NA2        g0719(.A(i_12_), .B(i_8_), .Y(new_new_n742_));
  OAI210     g0720(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n742_), .Y(new_new_n743_));
  INV        g0721(.A(new_new_n452_), .Y(new_new_n744_));
  AOI220     g0722(.A0(new_new_n325_), .A1(new_new_n583_), .B0(new_new_n743_), .B1(new_new_n741_), .Y(new_new_n745_));
  INV        g0723(.A(new_new_n745_), .Y(new_new_n746_));
  NO2        g0724(.A(new_new_n746_), .B(new_new_n739_), .Y(new_new_n747_));
  INV        g0725(.A(new_new_n173_), .Y(new_new_n748_));
  INV        g0726(.A(new_new_n248_), .Y(new_new_n749_));
  OAI210     g0727(.A0(new_new_n694_), .A1(new_new_n454_), .B0(new_new_n110_), .Y(new_new_n750_));
  AOI210     g0728(.A0(new_new_n750_), .A1(new_new_n749_), .B0(new_new_n748_), .Y(new_new_n751_));
  NO2        g0729(.A(new_new_n462_), .B(new_new_n26_), .Y(new_new_n752_));
  NO2        g0730(.A(new_new_n752_), .B(new_new_n428_), .Y(new_new_n753_));
  NA2        g0731(.A(new_new_n753_), .B(i_2_), .Y(new_new_n754_));
  INV        g0732(.A(new_new_n754_), .Y(new_new_n755_));
  AOI210     g0733(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n425_), .Y(new_new_n756_));
  AOI210     g0734(.A0(new_new_n756_), .A1(new_new_n755_), .B0(new_new_n751_), .Y(new_new_n757_));
  NO2        g0735(.A(new_new_n193_), .B(new_new_n125_), .Y(new_new_n758_));
  OAI210     g0736(.A0(new_new_n758_), .A1(new_new_n741_), .B0(i_2_), .Y(new_new_n759_));
  NO2        g0737(.A(new_new_n759_), .B(new_new_n196_), .Y(new_new_n760_));
  OA210      g0738(.A0(new_new_n622_), .A1(new_new_n126_), .B0(i_13_), .Y(new_new_n761_));
  NA2        g0739(.A(new_new_n202_), .B(new_new_n205_), .Y(new_new_n762_));
  NA2        g0740(.A(new_new_n152_), .B(new_new_n600_), .Y(new_new_n763_));
  AOI210     g0741(.A0(new_new_n763_), .A1(new_new_n762_), .B0(new_new_n380_), .Y(new_new_n764_));
  AOI210     g0742(.A0(new_new_n210_), .A1(new_new_n148_), .B0(new_new_n522_), .Y(new_new_n765_));
  NA2        g0743(.A(new_new_n765_), .B(new_new_n428_), .Y(new_new_n766_));
  NO2        g0744(.A(new_new_n102_), .B(new_new_n44_), .Y(new_new_n767_));
  INV        g0745(.A(new_new_n308_), .Y(new_new_n768_));
  NA4        g0746(.A(new_new_n768_), .B(new_new_n312_), .C(new_new_n124_), .D(new_new_n42_), .Y(new_new_n769_));
  OAI210     g0747(.A0(new_new_n769_), .A1(new_new_n767_), .B0(new_new_n766_), .Y(new_new_n770_));
  NO4        g0748(.A(new_new_n770_), .B(new_new_n764_), .C(new_new_n761_), .D(new_new_n760_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n583_), .B(new_new_n28_), .Y(new_new_n772_));
  NA2        g0750(.A(new_new_n740_), .B(new_new_n282_), .Y(new_new_n773_));
  NA2        g0751(.A(new_new_n773_), .B(new_new_n772_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n62_), .B(i_12_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n775_), .B(new_new_n126_), .Y(new_new_n776_));
  NO2        g0754(.A(new_new_n776_), .B(new_new_n600_), .Y(new_new_n777_));
  AOI220     g0755(.A0(new_new_n777_), .A1(new_new_n36_), .B0(new_new_n774_), .B1(new_new_n46_), .Y(new_new_n778_));
  NA4        g0756(.A(new_new_n778_), .B(new_new_n771_), .C(new_new_n757_), .D(new_new_n747_), .Y(men6));
  NO3        g0757(.A(i_9_), .B(new_new_n314_), .C(i_1_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n188_), .B(new_new_n139_), .Y(new_new_n781_));
  OAI210     g0759(.A0(new_new_n781_), .A1(new_new_n780_), .B0(new_new_n728_), .Y(new_new_n782_));
  INV        g0760(.A(new_new_n337_), .Y(new_new_n783_));
  AO210      g0761(.A0(new_new_n783_), .A1(new_new_n782_), .B0(i_12_), .Y(new_new_n784_));
  NA2        g0762(.A(new_new_n589_), .B(new_new_n63_), .Y(new_new_n785_));
  NA2        g0763(.A(new_new_n685_), .B(new_new_n71_), .Y(new_new_n786_));
  NA2        g0764(.A(new_new_n786_), .B(new_new_n785_), .Y(new_new_n787_));
  NA2        g0765(.A(new_new_n787_), .B(new_new_n73_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n336_), .Y(new_new_n789_));
  NA2        g0767(.A(new_new_n75_), .B(new_new_n131_), .Y(new_new_n790_));
  NO2        g0768(.A(new_new_n790_), .B(new_new_n789_), .Y(new_new_n791_));
  NO2        g0769(.A(new_new_n255_), .B(i_9_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n792_), .B(new_new_n775_), .Y(new_new_n793_));
  AOI210     g0771(.A0(new_new_n793_), .A1(new_new_n520_), .B0(new_new_n188_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n32_), .B(i_11_), .Y(new_new_n795_));
  NA3        g0773(.A(new_new_n795_), .B(new_new_n476_), .C(new_new_n396_), .Y(new_new_n796_));
  NAi32      g0774(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n797_));
  NO2        g0775(.A(new_new_n717_), .B(new_new_n797_), .Y(new_new_n798_));
  OAI210     g0776(.A0(new_new_n684_), .A1(new_new_n571_), .B0(new_new_n570_), .Y(new_new_n799_));
  NAi31      g0777(.An(new_new_n798_), .B(new_new_n799_), .C(new_new_n796_), .Y(new_new_n800_));
  OR3        g0778(.A(new_new_n800_), .B(new_new_n794_), .C(new_new_n791_), .Y(new_new_n801_));
  NO2        g0779(.A(new_new_n697_), .B(i_2_), .Y(new_new_n802_));
  NA2        g0780(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n803_));
  OAI210     g0781(.A0(new_new_n803_), .A1(new_new_n417_), .B0(new_new_n370_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n804_), .B(new_new_n802_), .Y(new_new_n805_));
  AO210      g0783(.A0(new_new_n369_), .A1(new_new_n361_), .B0(new_new_n403_), .Y(new_new_n806_));
  NA3        g0784(.A(new_new_n806_), .B(new_new_n259_), .C(i_7_), .Y(new_new_n807_));
  NA3        g0785(.A(new_new_n454_), .B(new_new_n147_), .C(new_new_n69_), .Y(new_new_n808_));
  AO210      g0786(.A0(new_new_n494_), .A1(new_new_n744_), .B0(new_new_n36_), .Y(new_new_n809_));
  NA4        g0787(.A(new_new_n809_), .B(new_new_n808_), .C(new_new_n807_), .D(new_new_n805_), .Y(new_new_n810_));
  NO2        g0788(.A(new_new_n638_), .B(i_11_), .Y(new_new_n811_));
  NA2        g0789(.A(new_new_n811_), .B(new_new_n570_), .Y(new_new_n812_));
  NA3        g0790(.A(new_new_n380_), .B(new_new_n241_), .C(new_new_n147_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n403_), .B(new_new_n70_), .Y(new_new_n814_));
  NA4        g0792(.A(new_new_n814_), .B(new_new_n813_), .C(new_new_n812_), .D(new_new_n606_), .Y(new_new_n815_));
  AN2        g0793(.A(new_new_n522_), .B(new_new_n46_), .Y(new_new_n816_));
  NA3        g0794(.A(new_new_n816_), .B(new_new_n485_), .C(new_new_n220_), .Y(new_new_n817_));
  AOI210     g0795(.A0(new_new_n454_), .A1(new_new_n452_), .B0(new_new_n569_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n111_), .B(new_new_n415_), .Y(new_new_n819_));
  INV        g0797(.A(new_new_n592_), .Y(new_new_n820_));
  NA3        g0798(.A(new_new_n820_), .B(new_new_n336_), .C(i_7_), .Y(new_new_n821_));
  NA4        g0799(.A(new_new_n821_), .B(new_new_n819_), .C(new_new_n818_), .D(new_new_n817_), .Y(new_new_n822_));
  NO4        g0800(.A(new_new_n822_), .B(new_new_n815_), .C(new_new_n810_), .D(new_new_n801_), .Y(new_new_n823_));
  NA4        g0801(.A(new_new_n823_), .B(new_new_n788_), .C(new_new_n784_), .D(new_new_n386_), .Y(men3));
  NA2        g0802(.A(i_12_), .B(i_10_), .Y(new_new_n825_));
  NA2        g0803(.A(i_6_), .B(i_7_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n826_), .B(i_0_), .Y(new_new_n827_));
  NO2        g0805(.A(i_11_), .B(new_new_n239_), .Y(new_new_n828_));
  OAI210     g0806(.A0(new_new_n827_), .A1(new_new_n296_), .B0(new_new_n828_), .Y(new_new_n829_));
  NO2        g0807(.A(new_new_n829_), .B(new_new_n196_), .Y(new_new_n830_));
  NO3        g0808(.A(new_new_n458_), .B(new_new_n89_), .C(new_new_n44_), .Y(new_new_n831_));
  OA210      g0809(.A0(new_new_n831_), .A1(new_new_n830_), .B0(new_new_n176_), .Y(new_new_n832_));
  NA3        g0810(.A(new_new_n813_), .B(new_new_n606_), .C(new_new_n379_), .Y(new_new_n833_));
  NA2        g0811(.A(new_new_n833_), .B(new_new_n40_), .Y(new_new_n834_));
  NO3        g0812(.A(new_new_n630_), .B(new_new_n462_), .C(new_new_n131_), .Y(new_new_n835_));
  AN2        g0813(.A(new_new_n460_), .B(new_new_n55_), .Y(new_new_n836_));
  NO2        g0814(.A(new_new_n836_), .B(new_new_n835_), .Y(new_new_n837_));
  AOI210     g0815(.A0(new_new_n837_), .A1(new_new_n834_), .B0(new_new_n48_), .Y(new_new_n838_));
  NO4        g0816(.A(new_new_n384_), .B(new_new_n389_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n188_), .B(new_new_n579_), .Y(new_new_n840_));
  NOi21      g0818(.An(new_new_n840_), .B(new_new_n839_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n706_), .B(new_new_n674_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n341_), .B(new_new_n446_), .Y(new_new_n843_));
  OAI220     g0821(.A0(new_new_n843_), .A1(new_new_n842_), .B0(new_new_n841_), .B1(new_new_n63_), .Y(new_new_n844_));
  NOi21      g0822(.An(i_5_), .B(i_9_), .Y(new_new_n845_));
  NA2        g0823(.A(new_new_n845_), .B(new_new_n451_), .Y(new_new_n846_));
  AOI210     g0824(.A0(new_new_n272_), .A1(new_new_n478_), .B0(new_new_n689_), .Y(new_new_n847_));
  NO3        g0825(.A(new_new_n421_), .B(new_new_n272_), .C(new_new_n73_), .Y(new_new_n848_));
  NO2        g0826(.A(new_new_n177_), .B(new_new_n148_), .Y(new_new_n849_));
  AOI210     g0827(.A0(new_new_n849_), .A1(new_new_n247_), .B0(new_new_n848_), .Y(new_new_n850_));
  OAI220     g0828(.A0(new_new_n850_), .A1(new_new_n183_), .B0(new_new_n847_), .B1(new_new_n846_), .Y(new_new_n851_));
  NO4        g0829(.A(new_new_n851_), .B(new_new_n844_), .C(new_new_n838_), .D(new_new_n832_), .Y(new_new_n852_));
  NA2        g0830(.A(new_new_n188_), .B(new_new_n24_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n319_), .B(new_new_n129_), .Y(new_new_n854_));
  NAi21      g0832(.An(new_new_n163_), .B(new_new_n446_), .Y(new_new_n855_));
  NO2        g0833(.A(new_new_n854_), .B(new_new_n408_), .Y(new_new_n856_));
  INV        g0834(.A(new_new_n856_), .Y(new_new_n857_));
  NO2        g0835(.A(new_new_n396_), .B(new_new_n300_), .Y(new_new_n858_));
  NA2        g0836(.A(new_new_n858_), .B(new_new_n708_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n580_), .B(i_0_), .Y(new_new_n860_));
  NO2        g0838(.A(new_new_n860_), .B(new_new_n391_), .Y(new_new_n861_));
  NO4        g0839(.A(new_new_n591_), .B(new_new_n217_), .C(new_new_n425_), .D(new_new_n417_), .Y(new_new_n862_));
  AOI210     g0840(.A0(new_new_n862_), .A1(i_11_), .B0(new_new_n861_), .Y(new_new_n863_));
  AN2        g0841(.A(new_new_n96_), .B(new_new_n246_), .Y(new_new_n864_));
  NA2        g0842(.A(new_new_n740_), .B(new_new_n337_), .Y(new_new_n865_));
  INV        g0843(.A(new_new_n58_), .Y(new_new_n866_));
  OAI220     g0844(.A0(new_new_n866_), .A1(new_new_n865_), .B0(new_new_n657_), .B1(new_new_n543_), .Y(new_new_n867_));
  NO2        g0845(.A(new_new_n257_), .B(new_new_n154_), .Y(new_new_n868_));
  NA2        g0846(.A(i_0_), .B(i_10_), .Y(new_new_n869_));
  OAI210     g0847(.A0(new_new_n869_), .A1(new_new_n85_), .B0(new_new_n545_), .Y(new_new_n870_));
  NO4        g0848(.A(new_new_n114_), .B(new_new_n58_), .C(new_new_n667_), .D(i_5_), .Y(new_new_n871_));
  AO220      g0849(.A0(new_new_n871_), .A1(new_new_n870_), .B0(new_new_n868_), .B1(i_6_), .Y(new_new_n872_));
  AOI220     g0850(.A0(new_new_n341_), .A1(new_new_n98_), .B0(new_new_n188_), .B1(new_new_n83_), .Y(new_new_n873_));
  NA2        g0851(.A(new_new_n574_), .B(i_4_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n191_), .B(new_new_n205_), .Y(new_new_n875_));
  OAI220     g0853(.A0(new_new_n875_), .A1(new_new_n865_), .B0(new_new_n874_), .B1(new_new_n873_), .Y(new_new_n876_));
  NO4        g0854(.A(new_new_n876_), .B(new_new_n872_), .C(new_new_n867_), .D(new_new_n864_), .Y(new_new_n877_));
  NA4        g0855(.A(new_new_n877_), .B(new_new_n863_), .C(new_new_n859_), .D(new_new_n857_), .Y(new_new_n878_));
  NO2        g0856(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n879_));
  NA2        g0857(.A(i_11_), .B(i_9_), .Y(new_new_n880_));
  NO3        g0858(.A(i_12_), .B(new_new_n880_), .C(new_new_n605_), .Y(new_new_n881_));
  AN2        g0859(.A(new_new_n881_), .B(new_new_n879_), .Y(new_new_n882_));
  NO2        g0860(.A(new_new_n48_), .B(i_7_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n400_), .B(new_new_n181_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n884_), .B(new_new_n161_), .Y(new_new_n885_));
  NO2        g0863(.A(new_new_n880_), .B(new_new_n73_), .Y(new_new_n886_));
  NO2        g0864(.A(new_new_n177_), .B(i_0_), .Y(new_new_n887_));
  INV        g0865(.A(new_new_n887_), .Y(new_new_n888_));
  NA2        g0866(.A(new_new_n476_), .B(new_new_n233_), .Y(new_new_n889_));
  NO2        g0867(.A(new_new_n889_), .B(new_new_n888_), .Y(new_new_n890_));
  NO3        g0868(.A(new_new_n890_), .B(new_new_n885_), .C(new_new_n882_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n656_), .B(new_new_n121_), .Y(new_new_n892_));
  NO2        g0870(.A(i_6_), .B(new_new_n892_), .Y(new_new_n893_));
  AOI210     g0871(.A0(new_new_n453_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n894_));
  NA2        g0872(.A(new_new_n173_), .B(new_new_n103_), .Y(new_new_n895_));
  NOi32      g0873(.An(new_new_n894_), .Bn(new_new_n191_), .C(new_new_n895_), .Y(new_new_n896_));
  NO2        g0874(.A(new_new_n896_), .B(new_new_n893_), .Y(new_new_n897_));
  NOi21      g0875(.An(i_7_), .B(i_5_), .Y(new_new_n898_));
  NOi31      g0876(.An(new_new_n898_), .B(i_0_), .C(new_new_n720_), .Y(new_new_n899_));
  NA3        g0877(.A(new_new_n899_), .B(new_new_n390_), .C(i_6_), .Y(new_new_n900_));
  OA210      g0878(.A0(new_new_n895_), .A1(new_new_n520_), .B0(new_new_n900_), .Y(new_new_n901_));
  NO3        g0879(.A(new_new_n411_), .B(new_new_n372_), .C(new_new_n368_), .Y(new_new_n902_));
  NO2        g0880(.A(new_new_n266_), .B(new_new_n326_), .Y(new_new_n903_));
  NO2        g0881(.A(new_new_n720_), .B(new_new_n261_), .Y(new_new_n904_));
  AOI210     g0882(.A0(new_new_n904_), .A1(new_new_n903_), .B0(new_new_n902_), .Y(new_new_n905_));
  NA4        g0883(.A(new_new_n905_), .B(new_new_n901_), .C(new_new_n897_), .D(new_new_n891_), .Y(new_new_n906_));
  NO2        g0884(.A(new_new_n853_), .B(new_new_n242_), .Y(new_new_n907_));
  AN2        g0885(.A(new_new_n340_), .B(new_new_n337_), .Y(new_new_n908_));
  AN2        g0886(.A(new_new_n908_), .B(new_new_n849_), .Y(new_new_n909_));
  OAI210     g0887(.A0(new_new_n909_), .A1(new_new_n907_), .B0(i_10_), .Y(new_new_n910_));
  NO2        g0888(.A(new_new_n825_), .B(new_new_n325_), .Y(new_new_n911_));
  NA2        g0889(.A(new_new_n911_), .B(new_new_n886_), .Y(new_new_n912_));
  NA3        g0890(.A(new_new_n475_), .B(new_new_n418_), .C(new_new_n45_), .Y(new_new_n913_));
  OAI210     g0891(.A0(new_new_n855_), .A1(i_6_), .B0(new_new_n913_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n259_), .B(new_new_n46_), .Y(new_new_n915_));
  NO2        g0893(.A(new_new_n915_), .B(new_new_n190_), .Y(new_new_n916_));
  AOI220     g0894(.A0(new_new_n916_), .A1(new_new_n476_), .B0(new_new_n914_), .B1(new_new_n73_), .Y(new_new_n917_));
  NA3        g0895(.A(new_new_n803_), .B(new_new_n388_), .C(new_new_n638_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n92_), .B(new_new_n44_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n75_), .B(new_new_n742_), .Y(new_new_n920_));
  AOI220     g0898(.A0(new_new_n920_), .A1(new_new_n919_), .B0(new_new_n176_), .B1(new_new_n599_), .Y(new_new_n921_));
  AOI210     g0899(.A0(new_new_n921_), .A1(new_new_n918_), .B0(new_new_n47_), .Y(new_new_n922_));
  NO3        g0900(.A(new_new_n591_), .B(new_new_n367_), .C(new_new_n24_), .Y(new_new_n923_));
  AOI210     g0901(.A0(new_new_n700_), .A1(new_new_n554_), .B0(new_new_n923_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n601_), .B(new_new_n105_), .Y(new_new_n925_));
  NA2        g0903(.A(new_new_n925_), .B(i_0_), .Y(new_new_n926_));
  OAI220     g0904(.A0(new_new_n926_), .A1(new_new_n85_), .B0(new_new_n924_), .B1(new_new_n174_), .Y(new_new_n927_));
  NO3        g0905(.A(new_new_n927_), .B(new_new_n922_), .C(new_new_n525_), .Y(new_new_n928_));
  NA4        g0906(.A(new_new_n928_), .B(new_new_n917_), .C(new_new_n912_), .D(new_new_n910_), .Y(new_new_n929_));
  NO3        g0907(.A(new_new_n929_), .B(new_new_n906_), .C(new_new_n878_), .Y(new_new_n930_));
  NO2        g0908(.A(i_0_), .B(new_new_n720_), .Y(new_new_n931_));
  NA2        g0909(.A(new_new_n73_), .B(new_new_n44_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n869_), .B(new_new_n932_), .Y(new_new_n933_));
  NO3        g0911(.A(new_new_n105_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n934_));
  AO220      g0912(.A0(new_new_n934_), .A1(new_new_n933_), .B0(new_new_n931_), .B1(new_new_n176_), .Y(new_new_n935_));
  AOI210     g0913(.A0(new_new_n785_), .A1(new_new_n687_), .B0(new_new_n895_), .Y(new_new_n936_));
  AOI210     g0914(.A0(new_new_n935_), .A1(new_new_n358_), .B0(new_new_n936_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n728_), .B(new_new_n146_), .Y(new_new_n938_));
  INV        g0916(.A(new_new_n938_), .Y(new_new_n939_));
  NA3        g0917(.A(new_new_n939_), .B(new_new_n674_), .C(new_new_n73_), .Y(new_new_n940_));
  NO2        g0918(.A(new_new_n799_), .B(new_new_n411_), .Y(new_new_n941_));
  NA3        g0919(.A(new_new_n827_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n942_));
  NA2        g0920(.A(new_new_n828_), .B(i_9_), .Y(new_new_n943_));
  AOI210     g0921(.A0(new_new_n942_), .A1(new_new_n500_), .B0(new_new_n943_), .Y(new_new_n944_));
  NA2        g0922(.A(new_new_n247_), .B(new_new_n232_), .Y(new_new_n945_));
  AOI210     g0923(.A0(new_new_n945_), .A1(new_new_n860_), .B0(new_new_n154_), .Y(new_new_n946_));
  NO3        g0924(.A(new_new_n946_), .B(new_new_n944_), .C(new_new_n941_), .Y(new_new_n947_));
  NA3        g0925(.A(new_new_n947_), .B(new_new_n940_), .C(new_new_n937_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n908_), .B(new_new_n380_), .Y(new_new_n949_));
  AOI210     g0927(.A0(new_new_n307_), .A1(new_new_n163_), .B0(new_new_n949_), .Y(new_new_n950_));
  NA3        g0928(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n951_));
  NA2        g0929(.A(new_new_n883_), .B(new_new_n489_), .Y(new_new_n952_));
  AOI210     g0930(.A0(new_new_n951_), .A1(new_new_n163_), .B0(new_new_n952_), .Y(new_new_n953_));
  NO2        g0931(.A(new_new_n953_), .B(new_new_n950_), .Y(new_new_n954_));
  NO3        g0932(.A(new_new_n869_), .B(new_new_n845_), .C(new_new_n193_), .Y(new_new_n955_));
  AOI220     g0933(.A0(new_new_n955_), .A1(i_11_), .B0(new_new_n575_), .B1(new_new_n75_), .Y(new_new_n956_));
  NO3        g0934(.A(new_new_n211_), .B(new_new_n389_), .C(i_0_), .Y(new_new_n957_));
  OAI210     g0935(.A0(new_new_n957_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n958_));
  INV        g0936(.A(new_new_n220_), .Y(new_new_n959_));
  OAI220     g0937(.A0(new_new_n536_), .A1(new_new_n139_), .B0(new_new_n643_), .B1(new_new_n616_), .Y(new_new_n960_));
  NA3        g0938(.A(new_new_n960_), .B(i_7_), .C(new_new_n959_), .Y(new_new_n961_));
  NA4        g0939(.A(new_new_n961_), .B(new_new_n958_), .C(new_new_n956_), .D(new_new_n954_), .Y(new_new_n962_));
  NO2        g0940(.A(new_new_n245_), .B(new_new_n92_), .Y(new_new_n963_));
  NA2        g0941(.A(new_new_n963_), .B(new_new_n931_), .Y(new_new_n964_));
  AOI220     g0942(.A0(new_new_n898_), .A1(new_new_n489_), .B0(new_new_n827_), .B1(new_new_n164_), .Y(new_new_n965_));
  NA2        g0943(.A(new_new_n361_), .B(new_new_n178_), .Y(new_new_n966_));
  OA220      g0944(.A0(new_new_n966_), .A1(new_new_n965_), .B0(new_new_n964_), .B1(i_5_), .Y(new_new_n967_));
  AOI210     g0945(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n177_), .Y(new_new_n968_));
  NA3        g0946(.A(new_new_n613_), .B(new_new_n188_), .C(new_new_n83_), .Y(new_new_n969_));
  NA2        g0947(.A(new_new_n969_), .B(new_new_n552_), .Y(new_new_n970_));
  INV        g0948(.A(new_new_n970_), .Y(new_new_n971_));
  NA3        g0949(.A(new_new_n396_), .B(new_new_n342_), .C(new_new_n223_), .Y(new_new_n972_));
  INV        g0950(.A(new_new_n972_), .Y(new_new_n973_));
  NOi31      g0951(.An(new_new_n395_), .B(new_new_n932_), .C(new_new_n242_), .Y(new_new_n974_));
  NO2        g0952(.A(new_new_n974_), .B(new_new_n973_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n975_), .B(new_new_n971_), .C(new_new_n967_), .Y(new_new_n976_));
  INV        g0954(.A(new_new_n615_), .Y(new_new_n977_));
  NO3        g0955(.A(new_new_n977_), .B(new_new_n567_), .C(new_new_n355_), .Y(new_new_n978_));
  NO2        g0956(.A(new_new_n85_), .B(i_5_), .Y(new_new_n979_));
  NA3        g0957(.A(new_new_n828_), .B(new_new_n109_), .C(new_new_n124_), .Y(new_new_n980_));
  INV        g0958(.A(new_new_n980_), .Y(new_new_n981_));
  AOI210     g0959(.A0(new_new_n981_), .A1(new_new_n979_), .B0(new_new_n978_), .Y(new_new_n982_));
  NA3        g0960(.A(new_new_n312_), .B(i_5_), .C(new_new_n196_), .Y(new_new_n983_));
  NAi31      g0961(.An(new_new_n244_), .B(new_new_n983_), .C(new_new_n245_), .Y(new_new_n984_));
  NO4        g0962(.A(new_new_n242_), .B(new_new_n211_), .C(i_0_), .D(i_12_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n985_), .B(new_new_n984_), .Y(new_new_n986_));
  AN2        g0964(.A(new_new_n869_), .B(new_new_n154_), .Y(new_new_n987_));
  NO4        g0965(.A(new_new_n987_), .B(i_12_), .C(new_new_n647_), .D(new_new_n131_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n988_), .B(new_new_n220_), .Y(new_new_n989_));
  NA3        g0967(.A(new_new_n98_), .B(new_new_n579_), .C(i_11_), .Y(new_new_n990_));
  NO2        g0968(.A(new_new_n990_), .B(new_new_n156_), .Y(new_new_n991_));
  NO2        g0969(.A(i_7_), .B(new_new_n983_), .Y(new_new_n992_));
  AOI210     g0970(.A0(new_new_n992_), .A1(new_new_n887_), .B0(new_new_n991_), .Y(new_new_n993_));
  NA4        g0971(.A(new_new_n993_), .B(new_new_n989_), .C(new_new_n986_), .D(new_new_n982_), .Y(new_new_n994_));
  NO4        g0972(.A(new_new_n994_), .B(new_new_n976_), .C(new_new_n962_), .D(new_new_n948_), .Y(new_new_n995_));
  OAI210     g0973(.A0(new_new_n802_), .A1(new_new_n795_), .B0(new_new_n37_), .Y(new_new_n996_));
  NA3        g0974(.A(new_new_n894_), .B(new_new_n375_), .C(i_5_), .Y(new_new_n997_));
  NA3        g0975(.A(new_new_n997_), .B(new_new_n996_), .C(new_new_n1043_), .Y(new_new_n998_));
  NA2        g0976(.A(new_new_n998_), .B(new_new_n208_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n189_), .B(new_new_n191_), .Y(new_new_n1000_));
  AO210      g0978(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n1000_), .Y(new_new_n1001_));
  OAI210     g0979(.A0(new_new_n615_), .A1(new_new_n613_), .B0(new_new_n325_), .Y(new_new_n1002_));
  NAi31      g0980(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1003_));
  AOI210     g0981(.A0(new_new_n117_), .A1(new_new_n70_), .B0(new_new_n1003_), .Y(new_new_n1004_));
  NO2        g0982(.A(new_new_n1004_), .B(new_new_n644_), .Y(new_new_n1005_));
  NA3        g0983(.A(new_new_n1005_), .B(new_new_n1002_), .C(new_new_n1001_), .Y(new_new_n1006_));
  NO2        g0984(.A(new_new_n465_), .B(new_new_n272_), .Y(new_new_n1007_));
  NO4        g0985(.A(new_new_n235_), .B(new_new_n145_), .C(new_new_n678_), .D(new_new_n37_), .Y(new_new_n1008_));
  NO3        g0986(.A(new_new_n1008_), .B(new_new_n1007_), .C(new_new_n862_), .Y(new_new_n1009_));
  OAI210     g0987(.A0(new_new_n990_), .A1(new_new_n148_), .B0(new_new_n1009_), .Y(new_new_n1010_));
  AOI210     g0988(.A0(new_new_n1006_), .A1(new_new_n48_), .B0(new_new_n1010_), .Y(new_new_n1011_));
  AOI210     g0989(.A0(new_new_n1011_), .A1(new_new_n999_), .B0(new_new_n73_), .Y(new_new_n1012_));
  INV        g0990(.A(new_new_n572_), .Y(new_new_n1013_));
  NO2        g0991(.A(new_new_n1013_), .B(new_new_n748_), .Y(new_new_n1014_));
  OAI210     g0992(.A0(new_new_n80_), .A1(new_new_n54_), .B0(new_new_n108_), .Y(new_new_n1015_));
  NA2        g0993(.A(new_new_n1015_), .B(new_new_n76_), .Y(new_new_n1016_));
  AOI210     g0994(.A0(new_new_n968_), .A1(new_new_n883_), .B0(new_new_n899_), .Y(new_new_n1017_));
  AOI210     g0995(.A0(new_new_n1017_), .A1(new_new_n1016_), .B0(new_new_n678_), .Y(new_new_n1018_));
  NA2        g0996(.A(new_new_n266_), .B(new_new_n57_), .Y(new_new_n1019_));
  NA2        g0997(.A(new_new_n1019_), .B(new_new_n76_), .Y(new_new_n1020_));
  NO2        g0998(.A(new_new_n1020_), .B(new_new_n239_), .Y(new_new_n1021_));
  NA3        g0999(.A(new_new_n96_), .B(new_new_n314_), .C(new_new_n31_), .Y(new_new_n1022_));
  INV        g1000(.A(new_new_n1022_), .Y(new_new_n1023_));
  NO3        g1001(.A(new_new_n1023_), .B(new_new_n1021_), .C(new_new_n1018_), .Y(new_new_n1024_));
  OAI210     g1002(.A0(new_new_n274_), .A1(new_new_n159_), .B0(new_new_n86_), .Y(new_new_n1025_));
  NA3        g1003(.A(new_new_n752_), .B(new_new_n296_), .C(new_new_n80_), .Y(new_new_n1026_));
  AOI210     g1004(.A0(new_new_n1026_), .A1(new_new_n1025_), .B0(i_11_), .Y(new_new_n1027_));
  OAI210     g1005(.A0(new_new_n1042_), .A1(new_new_n894_), .B0(new_new_n208_), .Y(new_new_n1028_));
  NA2        g1006(.A(new_new_n165_), .B(i_5_), .Y(new_new_n1029_));
  NO2        g1007(.A(new_new_n1028_), .B(new_new_n1029_), .Y(new_new_n1030_));
  NO3        g1008(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1031_));
  OAI210     g1009(.A0(new_new_n903_), .A1(new_new_n314_), .B0(new_new_n1031_), .Y(new_new_n1032_));
  NO2        g1010(.A(new_new_n1032_), .B(new_new_n720_), .Y(new_new_n1033_));
  NO3        g1011(.A(new_new_n1033_), .B(new_new_n1030_), .C(new_new_n1027_), .Y(new_new_n1034_));
  OAI210     g1012(.A0(new_new_n1024_), .A1(i_4_), .B0(new_new_n1034_), .Y(new_new_n1035_));
  NO3        g1013(.A(new_new_n1035_), .B(new_new_n1014_), .C(new_new_n1012_), .Y(new_new_n1036_));
  NA4        g1014(.A(new_new_n1036_), .B(new_new_n995_), .C(new_new_n930_), .D(new_new_n852_), .Y(men4));
  INV        g1015(.A(i_2_), .Y(new_new_n1040_));
  INV        g1016(.A(i_12_), .Y(new_new_n1041_));
  INV        g1017(.A(i_12_), .Y(new_new_n1042_));
  INV        g1018(.A(new_new_n162_), .Y(new_new_n1043_));
endmodule


