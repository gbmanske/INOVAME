//Benchmark atmr_intb_466_0.125

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n286_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n323_, ori_ori_n324_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n310_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n363_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n436_, men_men_n437_, men_men_n438_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  INV        o035(.A(ori_ori_n55_), .Y(ori_ori_n58_));
  NO2        o036(.A(x02), .B(ori_ori_n58_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n60_));
  OAI210     o038(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n60_), .Y(ori_ori_n61_));
  AOI220     o039(.A0(ori_ori_n61_), .A1(ori_ori_n55_), .B0(ori_ori_n59_), .B1(ori_ori_n31_), .Y(ori_ori_n62_));
  NO2        o040(.A(ori_ori_n62_), .B(x05), .Y(ori_ori_n63_));
  NA2        o041(.A(x09), .B(x05), .Y(ori_ori_n64_));
  NA2        o042(.A(x10), .B(x06), .Y(ori_ori_n65_));
  NA3        o043(.A(ori_ori_n65_), .B(ori_ori_n64_), .C(ori_ori_n28_), .Y(ori_ori_n66_));
  OAI210     o044(.A0(ori_ori_n66_), .A1(x07), .B0(x03), .Y(ori_ori_n67_));
  NOi31      o045(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n68_));
  INV        o046(.A(x07), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n24_), .Y(ori_ori_n70_));
  NO2        o048(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n71_));
  OAI210     o049(.A0(ori_ori_n71_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n48_), .B(ori_ori_n72_), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n74_));
  NO2        o052(.A(x08), .B(x01), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n35_), .Y(ori_ori_n76_));
  NO3        o054(.A(ori_ori_n76_), .B(ori_ori_n73_), .C(ori_ori_n70_), .Y(ori_ori_n77_));
  AN2        o055(.A(ori_ori_n77_), .B(ori_ori_n67_), .Y(ori_ori_n78_));
  INV        o056(.A(ori_ori_n76_), .Y(ori_ori_n79_));
  NA2        o057(.A(x11), .B(x00), .Y(ori_ori_n80_));
  NO2        o058(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n81_));
  NOi21      o059(.An(ori_ori_n80_), .B(ori_ori_n81_), .Y(ori_ori_n82_));
  NOi21      o060(.An(x01), .B(x10), .Y(ori_ori_n83_));
  NO2        o061(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n84_));
  NO3        o062(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(x06), .Y(ori_ori_n85_));
  NA2        o063(.A(ori_ori_n85_), .B(ori_ori_n27_), .Y(ori_ori_n86_));
  OAI210     o064(.A0(ori_ori_n323_), .A1(x07), .B0(ori_ori_n86_), .Y(ori_ori_n87_));
  NO3        o065(.A(ori_ori_n87_), .B(ori_ori_n78_), .C(ori_ori_n63_), .Y(ori01));
  INV        o066(.A(x12), .Y(ori_ori_n89_));
  INV        o067(.A(x13), .Y(ori_ori_n90_));
  NO2        o068(.A(x10), .B(x01), .Y(ori_ori_n91_));
  NO2        o069(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  NA2        o071(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n95_));
  NOi21      o073(.An(ori_ori_n95_), .B(ori_ori_n54_), .Y(ori_ori_n96_));
  NA2        o074(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n97_));
  NA2        o075(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n98_), .B(x05), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n35_), .B(ori_ori_n53_), .Y(ori_ori_n100_));
  INV        o078(.A(ori_ori_n96_), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n101_), .B(ori_ori_n65_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n103_));
  NA2        o081(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n104_), .B(ori_ori_n103_), .Y(ori_ori_n105_));
  NA2        o083(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n107_));
  NA3        o085(.A(ori_ori_n107_), .B(ori_ori_n106_), .C(x13), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n109_));
  NOi21      o087(.An(ori_ori_n108_), .B(ori_ori_n105_), .Y(ori_ori_n110_));
  NO3        o088(.A(ori_ori_n110_), .B(x06), .C(x03), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(ori_ori_n102_), .Y(ori_ori_n112_));
  NA2        o090(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n113_));
  OAI210     o091(.A0(ori_ori_n75_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n114_), .B(ori_ori_n113_), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n117_));
  AOI210     o095(.A0(ori_ori_n117_), .A1(ori_ori_n49_), .B0(ori_ori_n116_), .Y(ori_ori_n118_));
  AN2        o096(.A(ori_ori_n118_), .B(ori_ori_n115_), .Y(ori_ori_n119_));
  NO2        o097(.A(x09), .B(x05), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(ori_ori_n47_), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n93_), .B(ori_ori_n49_), .Y(ori_ori_n122_));
  NA2        o100(.A(x09), .B(x00), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n95_), .B(ori_ori_n123_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n122_), .B(ori_ori_n119_), .Y(ori_ori_n125_));
  NO2        o103(.A(x03), .B(x02), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n76_), .B(ori_ori_n90_), .Y(ori_ori_n127_));
  OAI210     o105(.A0(ori_ori_n127_), .A1(ori_ori_n96_), .B0(ori_ori_n126_), .Y(ori_ori_n128_));
  OA210      o106(.A0(ori_ori_n125_), .A1(x11), .B0(ori_ori_n128_), .Y(ori_ori_n129_));
  OAI210     o107(.A0(ori_ori_n112_), .A1(ori_ori_n23_), .B0(ori_ori_n129_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n93_), .B(ori_ori_n40_), .Y(ori_ori_n131_));
  NO2        o109(.A(ori_ori_n131_), .B(ori_ori_n41_), .Y(ori_ori_n132_));
  NO2        o110(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n133_));
  NA2        o111(.A(ori_ori_n90_), .B(x01), .Y(ori_ori_n134_));
  NO2        o112(.A(ori_ori_n133_), .B(ori_ori_n48_), .Y(ori_ori_n135_));
  AOI210     o113(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n136_));
  OAI210     o114(.A0(ori_ori_n135_), .A1(ori_ori_n132_), .B0(ori_ori_n136_), .Y(ori_ori_n137_));
  NA2        o115(.A(x10), .B(x05), .Y(ori_ori_n138_));
  NO2        o116(.A(x09), .B(x01), .Y(ori_ori_n139_));
  NO2        o117(.A(ori_ori_n95_), .B(x08), .Y(ori_ori_n140_));
  NO2        o118(.A(ori_ori_n84_), .B(x06), .Y(ori_ori_n141_));
  NOi21      o119(.An(x09), .B(x00), .Y(ori_ori_n142_));
  NO3        o120(.A(ori_ori_n74_), .B(ori_ori_n142_), .C(ori_ori_n47_), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n143_), .B(ori_ori_n104_), .Y(ori_ori_n144_));
  NA2        o122(.A(x06), .B(x05), .Y(ori_ori_n145_));
  OAI210     o123(.A0(ori_ori_n145_), .A1(ori_ori_n35_), .B0(ori_ori_n89_), .Y(ori_ori_n146_));
  AOI210     o124(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n146_), .Y(ori_ori_n147_));
  NA2        o125(.A(ori_ori_n147_), .B(ori_ori_n144_), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n90_), .B(x12), .Y(ori_ori_n149_));
  AOI210     o127(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n149_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n151_));
  NA2        o129(.A(ori_ori_n151_), .B(x02), .Y(ori_ori_n152_));
  NA2        o130(.A(ori_ori_n150_), .B(ori_ori_n148_), .Y(ori_ori_n153_));
  NA2        o131(.A(ori_ori_n153_), .B(ori_ori_n137_), .Y(ori_ori_n154_));
  AOI210     o132(.A0(ori_ori_n130_), .A1(ori_ori_n89_), .B0(ori_ori_n154_), .Y(ori_ori_n155_));
  INV        o133(.A(ori_ori_n66_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n156_), .B(ori_ori_n115_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n103_), .B(x06), .Y(ori_ori_n158_));
  INV        o136(.A(ori_ori_n158_), .Y(ori_ori_n159_));
  AOI210     o137(.A0(ori_ori_n159_), .A1(ori_ori_n157_), .B0(x12), .Y(ori_ori_n160_));
  INV        o138(.A(ori_ori_n68_), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n83_), .B(x06), .Y(ori_ori_n162_));
  AOI210     o140(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n50_), .Y(ori_ori_n163_));
  NO3        o141(.A(ori_ori_n163_), .B(ori_ori_n162_), .C(ori_ori_n41_), .Y(ori_ori_n164_));
  INV        o142(.A(ori_ori_n117_), .Y(ori_ori_n165_));
  OAI210     o143(.A0(ori_ori_n165_), .A1(ori_ori_n164_), .B0(x02), .Y(ori_ori_n166_));
  AOI210     o144(.A0(ori_ori_n166_), .A1(ori_ori_n53_), .B0(ori_ori_n23_), .Y(ori_ori_n167_));
  OAI210     o145(.A0(ori_ori_n160_), .A1(ori_ori_n53_), .B0(ori_ori_n167_), .Y(ori_ori_n168_));
  INV        o146(.A(ori_ori_n117_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n170_));
  OAI210     o148(.A0(ori_ori_n71_), .A1(ori_ori_n36_), .B0(ori_ori_n97_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n90_), .B(x03), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n173_));
  NOi21      o151(.An(x13), .B(x04), .Y(ori_ori_n174_));
  NO3        o152(.A(ori_ori_n174_), .B(ori_ori_n68_), .C(ori_ori_n142_), .Y(ori_ori_n175_));
  NO2        o153(.A(ori_ori_n175_), .B(x05), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(ori_ori_n173_), .Y(ori_ori_n177_));
  INV        o155(.A(ori_ori_n177_), .Y(ori_ori_n178_));
  INV        o156(.A(ori_ori_n81_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n179_), .B(x12), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n181_));
  AOI210     o159(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n182_));
  NO2        o160(.A(x06), .B(x00), .Y(ori_ori_n183_));
  NO3        o161(.A(ori_ori_n183_), .B(ori_ori_n182_), .C(ori_ori_n41_), .Y(ori_ori_n184_));
  INV        o162(.A(ori_ori_n65_), .Y(ori_ori_n185_));
  NO2        o163(.A(ori_ori_n185_), .B(ori_ori_n184_), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n187_));
  INV        o165(.A(x03), .Y(ori_ori_n188_));
  OR2        o166(.A(ori_ori_n188_), .B(ori_ori_n186_), .Y(ori_ori_n189_));
  NA2        o167(.A(x13), .B(ori_ori_n89_), .Y(ori_ori_n190_));
  NA3        o168(.A(ori_ori_n190_), .B(ori_ori_n146_), .C(ori_ori_n82_), .Y(ori_ori_n191_));
  OAI210     o169(.A0(ori_ori_n189_), .A1(ori_ori_n181_), .B0(ori_ori_n191_), .Y(ori_ori_n192_));
  AOI210     o170(.A0(ori_ori_n180_), .A1(ori_ori_n178_), .B0(ori_ori_n192_), .Y(ori_ori_n193_));
  AOI210     o171(.A0(ori_ori_n193_), .A1(ori_ori_n168_), .B0(x07), .Y(ori_ori_n194_));
  NA2        o172(.A(ori_ori_n64_), .B(ori_ori_n29_), .Y(ori_ori_n195_));
  NOi31      o173(.An(ori_ori_n113_), .B(ori_ori_n174_), .C(ori_ori_n142_), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n196_), .B(ori_ori_n195_), .Y(ori_ori_n197_));
  OAI210     o175(.A0(ori_ori_n68_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n198_));
  INV        o176(.A(ori_ori_n198_), .Y(ori_ori_n199_));
  NO2        o177(.A(x12), .B(x02), .Y(ori_ori_n200_));
  INV        o178(.A(ori_ori_n200_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n201_), .B(ori_ori_n179_), .Y(ori_ori_n202_));
  OA210      o180(.A0(ori_ori_n199_), .A1(ori_ori_n197_), .B0(ori_ori_n202_), .Y(ori_ori_n203_));
  NA2        o181(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n204_), .B(x01), .Y(ori_ori_n205_));
  INV        o183(.A(ori_ori_n205_), .Y(ori_ori_n206_));
  AOI210     o184(.A0(ori_ori_n206_), .A1(ori_ori_n108_), .B0(ori_ori_n29_), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n90_), .B(x04), .Y(ori_ori_n208_));
  NO3        o186(.A(ori_ori_n80_), .B(x12), .C(x03), .Y(ori_ori_n209_));
  NA2        o187(.A(ori_ori_n207_), .B(ori_ori_n209_), .Y(ori_ori_n210_));
  NOi21      o188(.An(ori_ori_n195_), .B(ori_ori_n162_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n212_));
  NA2        o190(.A(ori_ori_n211_), .B(ori_ori_n212_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n214_));
  NO3        o192(.A(ori_ori_n214_), .B(ori_ori_n163_), .C(ori_ori_n141_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n181_), .B(ori_ori_n28_), .Y(ori_ori_n216_));
  OAI210     o194(.A0(ori_ori_n215_), .A1(ori_ori_n169_), .B0(ori_ori_n216_), .Y(ori_ori_n217_));
  NA3        o195(.A(ori_ori_n217_), .B(ori_ori_n213_), .C(ori_ori_n210_), .Y(ori_ori_n218_));
  NO3        o196(.A(ori_ori_n218_), .B(ori_ori_n203_), .C(ori_ori_n194_), .Y(ori_ori_n219_));
  OAI210     o197(.A0(ori_ori_n155_), .A1(ori_ori_n57_), .B0(ori_ori_n219_), .Y(ori02));
  AOI210     o198(.A0(ori_ori_n113_), .A1(ori_ori_n76_), .B0(ori_ori_n106_), .Y(ori_ori_n221_));
  NOi21      o199(.An(ori_ori_n175_), .B(ori_ori_n139_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n222_), .B(ori_ori_n32_), .Y(ori_ori_n223_));
  OAI210     o201(.A0(ori_ori_n223_), .A1(ori_ori_n221_), .B0(ori_ori_n138_), .Y(ori_ori_n224_));
  INV        o202(.A(ori_ori_n138_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n76_), .B(ori_ori_n50_), .Y(ori_ori_n226_));
  AOI220     o204(.A0(ori_ori_n226_), .A1(ori_ori_n225_), .B0(ori_ori_n127_), .B1(ori_ori_n126_), .Y(ori_ori_n227_));
  AOI210     o205(.A0(ori_ori_n227_), .A1(ori_ori_n224_), .B0(ori_ori_n48_), .Y(ori_ori_n228_));
  NO2        o206(.A(ori_ori_n187_), .B(ori_ori_n47_), .Y(ori_ori_n229_));
  NA2        o207(.A(ori_ori_n229_), .B(ori_ori_n176_), .Y(ori_ori_n230_));
  AN2        o208(.A(ori_ori_n172_), .B(ori_ori_n171_), .Y(ori_ori_n231_));
  OAI210     o209(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n232_));
  BUFFER     o210(.A(ori_ori_n121_), .Y(ori_ori_n233_));
  AOI210     o211(.A0(ori_ori_n233_), .A1(ori_ori_n114_), .B0(ori_ori_n232_), .Y(ori_ori_n234_));
  OAI210     o212(.A0(ori_ori_n234_), .A1(ori_ori_n231_), .B0(ori_ori_n84_), .Y(ori_ori_n235_));
  INV        o213(.A(ori_ori_n126_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(ori_ori_n105_), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n237_), .B(x13), .Y(ori_ori_n238_));
  NA3        o216(.A(ori_ori_n238_), .B(ori_ori_n235_), .C(ori_ori_n230_), .Y(ori_ori_n239_));
  NO2        o217(.A(ori_ori_n239_), .B(ori_ori_n228_), .Y(ori_ori_n240_));
  NA2        o218(.A(ori_ori_n116_), .B(x03), .Y(ori_ori_n241_));
  OAI210     o219(.A0(ori_ori_n324_), .A1(ori_ori_n214_), .B0(ori_ori_n241_), .Y(ori_ori_n242_));
  NA2        o220(.A(ori_ori_n242_), .B(ori_ori_n91_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n140_), .B(ori_ori_n92_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n208_), .B(ori_ori_n89_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n89_), .B(ori_ori_n41_), .Y(ori_ori_n246_));
  NA3        o224(.A(ori_ori_n246_), .B(ori_ori_n245_), .C(ori_ori_n105_), .Y(ori_ori_n247_));
  NA4        o225(.A(ori_ori_n247_), .B(ori_ori_n244_), .C(ori_ori_n243_), .D(ori_ori_n48_), .Y(ori_ori_n248_));
  INV        o226(.A(ori_ori_n151_), .Y(ori_ori_n249_));
  INV        o227(.A(ori_ori_n40_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n251_));
  OAI220     o229(.A0(ori_ori_n251_), .A1(ori_ori_n250_), .B0(ori_ori_n249_), .B1(ori_ori_n55_), .Y(ori_ori_n252_));
  NA2        o230(.A(ori_ori_n252_), .B(x02), .Y(ori_ori_n253_));
  NO3        o231(.A(ori_ori_n149_), .B(ori_ori_n133_), .C(ori_ori_n51_), .Y(ori_ori_n254_));
  OAI210     o232(.A0(ori_ori_n123_), .A1(ori_ori_n36_), .B0(ori_ori_n89_), .Y(ori_ori_n255_));
  OAI210     o233(.A0(ori_ori_n255_), .A1(ori_ori_n143_), .B0(ori_ori_n254_), .Y(ori_ori_n256_));
  NA3        o234(.A(ori_ori_n256_), .B(ori_ori_n253_), .C(x06), .Y(ori_ori_n257_));
  NO3        o235(.A(ori_ori_n214_), .B(ori_ori_n103_), .C(x08), .Y(ori_ori_n258_));
  INV        o236(.A(ori_ori_n258_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n260_));
  NO3        o238(.A(ori_ori_n95_), .B(ori_ori_n104_), .C(ori_ori_n38_), .Y(ori_ori_n261_));
  AOI210     o239(.A0(ori_ori_n254_), .A1(ori_ori_n260_), .B0(ori_ori_n261_), .Y(ori_ori_n262_));
  OAI210     o240(.A0(ori_ori_n259_), .A1(ori_ori_n28_), .B0(ori_ori_n262_), .Y(ori_ori_n263_));
  AN2        o241(.A(ori_ori_n263_), .B(x04), .Y(ori_ori_n264_));
  AOI210     o242(.A0(ori_ori_n257_), .A1(ori_ori_n248_), .B0(ori_ori_n264_), .Y(ori_ori_n265_));
  OAI210     o243(.A0(ori_ori_n240_), .A1(x12), .B0(ori_ori_n265_), .Y(ori03));
  OR2        o244(.A(ori_ori_n42_), .B(ori_ori_n170_), .Y(ori_ori_n267_));
  AOI210     o245(.A0(ori_ori_n127_), .A1(ori_ori_n89_), .B0(ori_ori_n267_), .Y(ori_ori_n268_));
  NA2        o246(.A(ori_ori_n149_), .B(ori_ori_n126_), .Y(ori_ori_n269_));
  NA2        o247(.A(ori_ori_n269_), .B(ori_ori_n152_), .Y(ori_ori_n270_));
  OAI210     o248(.A0(ori_ori_n270_), .A1(ori_ori_n268_), .B0(x05), .Y(ori_ori_n271_));
  NA2        o249(.A(ori_ori_n267_), .B(x05), .Y(ori_ori_n272_));
  AOI210     o250(.A0(ori_ori_n114_), .A1(ori_ori_n161_), .B0(ori_ori_n272_), .Y(ori_ori_n273_));
  AOI210     o251(.A0(ori_ori_n172_), .A1(ori_ori_n41_), .B0(ori_ori_n99_), .Y(ori_ori_n274_));
  NO2        o252(.A(ori_ori_n274_), .B(ori_ori_n55_), .Y(ori_ori_n275_));
  OAI210     o253(.A0(ori_ori_n275_), .A1(ori_ori_n273_), .B0(ori_ori_n89_), .Y(ori_ori_n276_));
  AOI210     o254(.A0(ori_ori_n121_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n277_));
  NO2        o255(.A(ori_ori_n139_), .B(ori_ori_n109_), .Y(ori_ori_n278_));
  OAI220     o256(.A0(ori_ori_n278_), .A1(ori_ori_n37_), .B0(ori_ori_n124_), .B1(x13), .Y(ori_ori_n279_));
  OAI210     o257(.A0(ori_ori_n279_), .A1(ori_ori_n277_), .B0(x04), .Y(ori_ori_n280_));
  NO3        o258(.A(ori_ori_n246_), .B(ori_ori_n76_), .C(ori_ori_n55_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n89_), .B(ori_ori_n121_), .Y(ori_ori_n282_));
  AN2        o260(.A(x12), .B(ori_ori_n109_), .Y(ori_ori_n283_));
  NO3        o261(.A(ori_ori_n283_), .B(ori_ori_n282_), .C(ori_ori_n281_), .Y(ori_ori_n284_));
  NA4        o262(.A(ori_ori_n284_), .B(ori_ori_n280_), .C(ori_ori_n276_), .D(ori_ori_n271_), .Y(ori04));
  NO2        o263(.A(ori_ori_n79_), .B(ori_ori_n39_), .Y(ori_ori_n286_));
  XO2        o264(.A(ori_ori_n286_), .B(ori_ori_n190_), .Y(ori05));
  NO2        o265(.A(x06), .B(ori_ori_n24_), .Y(ori_ori_n288_));
  OAI210     o266(.A0(ori_ori_n288_), .A1(x03), .B0(ori_ori_n89_), .Y(ori_ori_n289_));
  OAI210     o267(.A0(ori_ori_n26_), .A1(ori_ori_n89_), .B0(x07), .Y(ori_ori_n290_));
  INV        o268(.A(ori_ori_n290_), .Y(ori_ori_n291_));
  NA2        o269(.A(ori_ori_n183_), .B(ori_ori_n179_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n292_), .B(ori_ori_n181_), .Y(ori_ori_n293_));
  NA2        o271(.A(ori_ori_n293_), .B(ori_ori_n89_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n33_), .B(ori_ori_n89_), .Y(ori_ori_n295_));
  AOI210     o273(.A0(ori_ori_n295_), .A1(ori_ori_n81_), .B0(x07), .Y(ori_ori_n296_));
  AOI220     o274(.A0(ori_ori_n296_), .A1(ori_ori_n294_), .B0(ori_ori_n291_), .B1(ori_ori_n289_), .Y(ori_ori_n297_));
  NO2        o275(.A(ori_ori_n94_), .B(ori_ori_n200_), .Y(ori_ori_n298_));
  NOi21      o276(.An(ori_ori_n241_), .B(ori_ori_n109_), .Y(ori_ori_n299_));
  NO2        o277(.A(ori_ori_n299_), .B(ori_ori_n201_), .Y(ori_ori_n300_));
  AOI210     o278(.A0(ori_ori_n190_), .A1(ori_ori_n47_), .B0(x04), .Y(ori_ori_n301_));
  NO4        o279(.A(ori_ori_n301_), .B(ori_ori_n300_), .C(ori_ori_n298_), .D(x08), .Y(ori_ori_n302_));
  NO2        o280(.A(ori_ori_n106_), .B(ori_ori_n28_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n303_), .B(ori_ori_n205_), .Y(ori_ori_n304_));
  OR3        o282(.A(ori_ori_n304_), .B(x12), .C(x03), .Y(ori_ori_n305_));
  NA3        o283(.A(ori_ori_n249_), .B(ori_ori_n100_), .C(x12), .Y(ori_ori_n306_));
  AO210      o284(.A0(ori_ori_n249_), .A1(ori_ori_n100_), .B0(ori_ori_n190_), .Y(ori_ori_n307_));
  NA4        o285(.A(ori_ori_n307_), .B(ori_ori_n306_), .C(ori_ori_n305_), .D(x08), .Y(ori_ori_n308_));
  INV        o286(.A(ori_ori_n308_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n302_), .B(ori_ori_n309_), .Y(ori_ori_n310_));
  NA3        o288(.A(ori_ori_n304_), .B(ori_ori_n299_), .C(ori_ori_n245_), .Y(ori_ori_n311_));
  INV        o289(.A(x14), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n134_), .B(ori_ori_n53_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n313_), .B(ori_ori_n312_), .Y(ori_ori_n314_));
  NA2        o292(.A(ori_ori_n314_), .B(ori_ori_n311_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n295_), .B(ori_ori_n57_), .Y(ori_ori_n316_));
  INV        o294(.A(ori_ori_n124_), .Y(ori_ori_n317_));
  NA2        o295(.A(ori_ori_n317_), .B(ori_ori_n89_), .Y(ori_ori_n318_));
  OAI210     o296(.A0(ori_ori_n316_), .A1(ori_ori_n80_), .B0(ori_ori_n318_), .Y(ori_ori_n319_));
  NO4        o297(.A(ori_ori_n319_), .B(ori_ori_n315_), .C(ori_ori_n310_), .D(ori_ori_n297_), .Y(ori06));
  INV        o298(.A(ori_ori_n82_), .Y(ori_ori_n323_));
  INV        o299(.A(x08), .Y(ori_ori_n324_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO2        m027(.A(mai_mai_n49_), .B(x11), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NO2        m048(.A(mai_mai_n61_), .B(mai_mai_n23_), .Y(mai_mai_n71_));
  NA2        m049(.A(x09), .B(x05), .Y(mai_mai_n72_));
  NA2        m050(.A(x10), .B(x06), .Y(mai_mai_n73_));
  NA2        m051(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  NO2        m052(.A(mai_mai_n61_), .B(mai_mai_n41_), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n74_), .A1(mai_mai_n71_), .B0(x03), .Y(mai_mai_n76_));
  NOi31      m054(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n373_), .B(mai_mai_n24_), .Y(mai_mai_n78_));
  NO2        m056(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n79_));
  NO2        m057(.A(mai_mai_n79_), .B(mai_mai_n36_), .Y(mai_mai_n80_));
  OAI210     m058(.A0(mai_mai_n79_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n81_));
  AOI210     m059(.A0(mai_mai_n80_), .A1(mai_mai_n48_), .B0(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m060(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n83_));
  NO2        m061(.A(x08), .B(x01), .Y(mai_mai_n84_));
  OAI210     m062(.A0(mai_mai_n84_), .A1(mai_mai_n83_), .B0(mai_mai_n35_), .Y(mai_mai_n85_));
  NO3        m063(.A(mai_mai_n85_), .B(mai_mai_n82_), .C(mai_mai_n78_), .Y(mai_mai_n86_));
  AN2        m064(.A(mai_mai_n86_), .B(mai_mai_n76_), .Y(mai_mai_n87_));
  INV        m065(.A(mai_mai_n85_), .Y(mai_mai_n88_));
  NA2        m066(.A(x11), .B(x00), .Y(mai_mai_n89_));
  NO2        m067(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n90_));
  NOi21      m068(.An(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  NOi21      m069(.An(x01), .B(x10), .Y(mai_mai_n92_));
  NO2        m070(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n93_));
  NO3        m071(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(x06), .Y(mai_mai_n94_));
  NA2        m072(.A(mai_mai_n94_), .B(mai_mai_n27_), .Y(mai_mai_n95_));
  OAI210     m073(.A0(mai_mai_n374_), .A1(x07), .B0(mai_mai_n95_), .Y(mai_mai_n96_));
  NO3        m074(.A(mai_mai_n96_), .B(mai_mai_n87_), .C(mai_mai_n70_), .Y(mai01));
  INV        m075(.A(x12), .Y(mai_mai_n98_));
  INV        m076(.A(x13), .Y(mai_mai_n99_));
  NA2        m077(.A(x08), .B(x04), .Y(mai_mai_n100_));
  NA2        m078(.A(mai_mai_n92_), .B(mai_mai_n28_), .Y(mai_mai_n101_));
  NO2        m079(.A(x10), .B(x01), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NA2        m082(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n84_), .B(x13), .Y(mai_mai_n108_));
  NA2        m086(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(x05), .Y(mai_mai_n110_));
  NA2        m088(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n111_));
  NA2        m089(.A(mai_mai_n57_), .B(mai_mai_n80_), .Y(mai_mai_n112_));
  AOI210     m090(.A0(mai_mai_n112_), .A1(mai_mai_n108_), .B0(mai_mai_n73_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n114_));
  NA2        m092(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n115_));
  NA2        m093(.A(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n118_));
  NO3        m096(.A(x00), .B(x06), .C(x03), .Y(mai_mai_n119_));
  NO3        m097(.A(mai_mai_n119_), .B(mai_mai_n113_), .C(mai_mai_n106_), .Y(mai_mai_n120_));
  OAI210     m098(.A0(mai_mai_n84_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n121_));
  NO2        m099(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n123_));
  NO2        m101(.A(x09), .B(x05), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n124_), .B(mai_mai_n47_), .Y(mai_mai_n125_));
  AOI210     m103(.A0(mai_mai_n125_), .A1(mai_mai_n104_), .B0(mai_mai_n49_), .Y(mai_mai_n126_));
  NA2        m104(.A(x09), .B(x00), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n107_), .B(mai_mai_n127_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n77_), .B(mai_mai_n51_), .Y(mai_mai_n129_));
  AOI210     m107(.A0(mai_mai_n129_), .A1(mai_mai_n128_), .B0(mai_mai_n123_), .Y(mai_mai_n130_));
  NO2        m108(.A(mai_mai_n130_), .B(mai_mai_n126_), .Y(mai_mai_n131_));
  NO2        m109(.A(x03), .B(x02), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n85_), .B(mai_mai_n99_), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n134_));
  OA210      m112(.A0(mai_mai_n131_), .A1(x11), .B0(mai_mai_n134_), .Y(mai_mai_n135_));
  OAI210     m113(.A0(mai_mai_n120_), .A1(mai_mai_n23_), .B0(mai_mai_n135_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n104_), .B(mai_mai_n40_), .Y(mai_mai_n137_));
  NAi21      m115(.An(x06), .B(x10), .Y(mai_mai_n138_));
  NA2        m116(.A(x01), .B(mai_mai_n138_), .Y(mai_mai_n139_));
  BUFFER     m117(.A(mai_mai_n139_), .Y(mai_mai_n140_));
  AOI210     m118(.A0(mai_mai_n140_), .A1(mai_mai_n137_), .B0(mai_mai_n41_), .Y(mai_mai_n141_));
  NO2        m119(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n99_), .B(x01), .Y(mai_mai_n143_));
  NO2        m121(.A(mai_mai_n143_), .B(x08), .Y(mai_mai_n144_));
  AOI210     m122(.A0(x09), .A1(mai_mai_n142_), .B0(mai_mai_n48_), .Y(mai_mai_n145_));
  AOI210     m123(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n146_));
  OAI210     m124(.A0(mai_mai_n145_), .A1(mai_mai_n141_), .B0(mai_mai_n146_), .Y(mai_mai_n147_));
  NA2        m125(.A(x04), .B(x02), .Y(mai_mai_n148_));
  NA2        m126(.A(x10), .B(x05), .Y(mai_mai_n149_));
  INV        m127(.A(x03), .Y(mai_mai_n150_));
  NA2        m128(.A(x11), .B(mai_mai_n150_), .Y(mai_mai_n151_));
  NAi21      m129(.An(mai_mai_n148_), .B(mai_mai_n151_), .Y(mai_mai_n152_));
  INV        m130(.A(mai_mai_n25_), .Y(mai_mai_n153_));
  NAi21      m131(.An(x13), .B(x00), .Y(mai_mai_n154_));
  AOI210     m132(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n154_), .Y(mai_mai_n155_));
  AOI220     m133(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n156_));
  AN2        m134(.A(x04), .B(mai_mai_n155_), .Y(mai_mai_n157_));
  BUFFER     m135(.A(mai_mai_n72_), .Y(mai_mai_n158_));
  NO2        m136(.A(mai_mai_n154_), .B(mai_mai_n36_), .Y(mai_mai_n159_));
  INV        m137(.A(mai_mai_n159_), .Y(mai_mai_n160_));
  OAI210     m138(.A0(mai_mai_n57_), .A1(mai_mai_n158_), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  OAI210     m139(.A0(mai_mai_n161_), .A1(mai_mai_n157_), .B0(mai_mai_n153_), .Y(mai_mai_n162_));
  NOi21      m140(.An(x09), .B(x00), .Y(mai_mai_n163_));
  NO2        m141(.A(mai_mai_n163_), .B(mai_mai_n47_), .Y(mai_mai_n164_));
  NO2        m142(.A(mai_mai_n99_), .B(x12), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n167_));
  NA2        m145(.A(mai_mai_n166_), .B(x12), .Y(mai_mai_n168_));
  NA4        m146(.A(mai_mai_n168_), .B(mai_mai_n162_), .C(mai_mai_n152_), .D(mai_mai_n147_), .Y(mai_mai_n169_));
  AOI210     m147(.A0(mai_mai_n136_), .A1(mai_mai_n98_), .B0(mai_mai_n169_), .Y(mai_mai_n170_));
  NA2        m148(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n171_));
  NA2        m149(.A(mai_mai_n171_), .B(mai_mai_n121_), .Y(mai_mai_n172_));
  AOI210     m150(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n114_), .B(x06), .Y(mai_mai_n174_));
  AOI210     m152(.A0(mai_mai_n173_), .A1(mai_mai_n172_), .B0(mai_mai_n174_), .Y(mai_mai_n175_));
  NO2        m153(.A(mai_mai_n175_), .B(x12), .Y(mai_mai_n176_));
  INV        m154(.A(mai_mai_n77_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n139_), .B(mai_mai_n57_), .Y(mai_mai_n178_));
  INV        m156(.A(mai_mai_n178_), .Y(mai_mai_n179_));
  NA2        m157(.A(mai_mai_n56_), .B(x02), .Y(mai_mai_n180_));
  AOI210     m158(.A0(mai_mai_n180_), .A1(mai_mai_n179_), .B0(mai_mai_n23_), .Y(mai_mai_n181_));
  OAI210     m159(.A0(mai_mai_n176_), .A1(mai_mai_n57_), .B0(mai_mai_n181_), .Y(mai_mai_n182_));
  INV        m160(.A(mai_mai_n123_), .Y(mai_mai_n183_));
  NO2        m161(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n99_), .B(x03), .Y(mai_mai_n185_));
  AOI210     m163(.A0(mai_mai_n77_), .A1(mai_mai_n184_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  NA2        m164(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n187_));
  INV        m165(.A(mai_mai_n138_), .Y(mai_mai_n188_));
  NOi21      m166(.An(x13), .B(x04), .Y(mai_mai_n189_));
  NO3        m167(.A(mai_mai_n189_), .B(mai_mai_n77_), .C(mai_mai_n163_), .Y(mai_mai_n190_));
  NO2        m168(.A(mai_mai_n190_), .B(x05), .Y(mai_mai_n191_));
  AOI220     m169(.A0(mai_mai_n191_), .A1(mai_mai_n187_), .B0(mai_mai_n188_), .B1(mai_mai_n57_), .Y(mai_mai_n192_));
  OAI210     m170(.A0(mai_mai_n186_), .A1(mai_mai_n183_), .B0(mai_mai_n192_), .Y(mai_mai_n193_));
  INV        m171(.A(mai_mai_n90_), .Y(mai_mai_n194_));
  NO2        m172(.A(mai_mai_n194_), .B(x12), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n196_));
  OAI210     m174(.A0(x08), .A1(x04), .B0(mai_mai_n155_), .Y(mai_mai_n197_));
  AOI210     m175(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n127_), .B(mai_mai_n73_), .Y(mai_mai_n199_));
  INV        m177(.A(mai_mai_n199_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n201_));
  NA2        m179(.A(mai_mai_n201_), .B(x03), .Y(mai_mai_n202_));
  OA210      m180(.A0(mai_mai_n202_), .A1(mai_mai_n200_), .B0(mai_mai_n197_), .Y(mai_mai_n203_));
  NA2        m181(.A(x13), .B(mai_mai_n98_), .Y(mai_mai_n204_));
  NA3        m182(.A(mai_mai_n204_), .B(x12), .C(mai_mai_n91_), .Y(mai_mai_n205_));
  OAI210     m183(.A0(mai_mai_n203_), .A1(mai_mai_n196_), .B0(mai_mai_n205_), .Y(mai_mai_n206_));
  AOI210     m184(.A0(mai_mai_n195_), .A1(mai_mai_n193_), .B0(mai_mai_n206_), .Y(mai_mai_n207_));
  AOI210     m185(.A0(mai_mai_n207_), .A1(mai_mai_n182_), .B0(x07), .Y(mai_mai_n208_));
  NA2        m186(.A(mai_mai_n72_), .B(mai_mai_n29_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n189_), .B(mai_mai_n163_), .Y(mai_mai_n210_));
  AOI210     m188(.A0(mai_mai_n210_), .A1(mai_mai_n129_), .B0(mai_mai_n209_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n99_), .B(x06), .Y(mai_mai_n212_));
  INV        m190(.A(mai_mai_n212_), .Y(mai_mai_n213_));
  NO2        m191(.A(x08), .B(x05), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n214_), .B(mai_mai_n198_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n215_), .B(mai_mai_n213_), .Y(mai_mai_n216_));
  NO2        m194(.A(x12), .B(x02), .Y(mai_mai_n217_));
  INV        m195(.A(mai_mai_n217_), .Y(mai_mai_n218_));
  NO2        m196(.A(mai_mai_n218_), .B(mai_mai_n194_), .Y(mai_mai_n219_));
  OA210      m197(.A0(mai_mai_n216_), .A1(mai_mai_n211_), .B0(mai_mai_n219_), .Y(mai_mai_n220_));
  NA2        m198(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n221_), .B(x01), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n84_), .B(mai_mai_n222_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n223_), .B(mai_mai_n29_), .Y(mai_mai_n224_));
  INV        m202(.A(mai_mai_n212_), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n99_), .B(x04), .Y(mai_mai_n226_));
  OAI210     m204(.A0(x02), .A1(mai_mai_n108_), .B0(mai_mai_n225_), .Y(mai_mai_n227_));
  NO3        m205(.A(mai_mai_n89_), .B(x12), .C(x03), .Y(mai_mai_n228_));
  OAI210     m206(.A0(mai_mai_n227_), .A1(mai_mai_n224_), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  NO2        m207(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n230_));
  OAI210     m208(.A0(x06), .A1(mai_mai_n92_), .B0(mai_mai_n230_), .Y(mai_mai_n231_));
  NA2        m209(.A(mai_mai_n231_), .B(mai_mai_n229_), .Y(mai_mai_n232_));
  NO3        m210(.A(mai_mai_n232_), .B(mai_mai_n220_), .C(mai_mai_n208_), .Y(mai_mai_n233_));
  OAI210     m211(.A0(mai_mai_n170_), .A1(mai_mai_n61_), .B0(mai_mai_n233_), .Y(mai02));
  BUFFER     m212(.A(mai_mai_n190_), .Y(mai_mai_n235_));
  NO2        m213(.A(mai_mai_n99_), .B(mai_mai_n35_), .Y(mai_mai_n236_));
  NA3        m214(.A(mai_mai_n236_), .B(x10), .C(mai_mai_n56_), .Y(mai_mai_n237_));
  OAI210     m215(.A0(mai_mai_n235_), .A1(mai_mai_n32_), .B0(mai_mai_n237_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n238_), .B(mai_mai_n149_), .Y(mai_mai_n239_));
  INV        m217(.A(mai_mai_n149_), .Y(mai_mai_n240_));
  OAI220     m218(.A0(mai_mai_n376_), .A1(mai_mai_n99_), .B0(mai_mai_n85_), .B1(mai_mai_n51_), .Y(mai_mai_n241_));
  AOI220     m219(.A0(mai_mai_n241_), .A1(mai_mai_n240_), .B0(mai_mai_n133_), .B1(mai_mai_n132_), .Y(mai_mai_n242_));
  AOI210     m220(.A0(mai_mai_n242_), .A1(mai_mai_n239_), .B0(mai_mai_n48_), .Y(mai_mai_n243_));
  NO2        m221(.A(x05), .B(x02), .Y(mai_mai_n244_));
  OAI210     m222(.A0(mai_mai_n172_), .A1(mai_mai_n163_), .B0(mai_mai_n244_), .Y(mai_mai_n245_));
  AOI220     m223(.A0(mai_mai_n214_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n246_));
  NOi21      m224(.An(mai_mai_n236_), .B(mai_mai_n246_), .Y(mai_mai_n247_));
  AOI210     m225(.A0(mai_mai_n189_), .A1(mai_mai_n79_), .B0(mai_mai_n247_), .Y(mai_mai_n248_));
  AOI210     m226(.A0(mai_mai_n248_), .A1(mai_mai_n245_), .B0(mai_mai_n123_), .Y(mai_mai_n249_));
  NAi21      m227(.An(mai_mai_n191_), .B(mai_mai_n186_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n201_), .B(mai_mai_n47_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n251_), .B(mai_mai_n250_), .Y(mai_mai_n252_));
  OAI210     m230(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n253_));
  NA2        m231(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n254_));
  AOI210     m232(.A0(mai_mai_n254_), .A1(mai_mai_n121_), .B0(mai_mai_n253_), .Y(mai_mai_n255_));
  OAI210     m233(.A0(mai_mai_n255_), .A1(mai_mai_n185_), .B0(mai_mai_n93_), .Y(mai_mai_n256_));
  NA3        m234(.A(mai_mai_n93_), .B(mai_mai_n84_), .C(mai_mai_n184_), .Y(mai_mai_n257_));
  NA3        m235(.A(mai_mai_n92_), .B(mai_mai_n83_), .C(mai_mai_n42_), .Y(mai_mai_n258_));
  AOI210     m236(.A0(mai_mai_n258_), .A1(mai_mai_n257_), .B0(x04), .Y(mai_mai_n259_));
  NO2        m237(.A(mai_mai_n215_), .B(mai_mai_n101_), .Y(mai_mai_n260_));
  AOI210     m238(.A0(mai_mai_n260_), .A1(x13), .B0(mai_mai_n259_), .Y(mai_mai_n261_));
  NA3        m239(.A(mai_mai_n261_), .B(mai_mai_n256_), .C(mai_mai_n252_), .Y(mai_mai_n262_));
  NO3        m240(.A(mai_mai_n262_), .B(mai_mai_n249_), .C(mai_mai_n243_), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n122_), .B(x03), .Y(mai_mai_n264_));
  OAI210     m242(.A0(mai_mai_n154_), .A1(mai_mai_n51_), .B0(mai_mai_n264_), .Y(mai_mai_n265_));
  NA2        m243(.A(mai_mai_n265_), .B(mai_mai_n102_), .Y(mai_mai_n266_));
  OAI220     m244(.A0(mai_mai_n226_), .A1(x09), .B0(mai_mai_n117_), .B1(mai_mai_n28_), .Y(mai_mai_n267_));
  NA2        m245(.A(mai_mai_n267_), .B(mai_mai_n103_), .Y(mai_mai_n268_));
  NA2        m246(.A(mai_mai_n226_), .B(mai_mai_n98_), .Y(mai_mai_n269_));
  NA2        m247(.A(mai_mai_n98_), .B(mai_mai_n41_), .Y(mai_mai_n270_));
  NA3        m248(.A(mai_mai_n270_), .B(mai_mai_n269_), .C(mai_mai_n116_), .Y(mai_mai_n271_));
  NA4        m249(.A(mai_mai_n271_), .B(mai_mai_n268_), .C(mai_mai_n266_), .D(mai_mai_n48_), .Y(mai_mai_n272_));
  INV        m250(.A(mai_mai_n167_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n144_), .B(mai_mai_n40_), .Y(mai_mai_n274_));
  NA2        m252(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n275_));
  OAI220     m253(.A0(mai_mai_n275_), .A1(mai_mai_n274_), .B0(mai_mai_n273_), .B1(mai_mai_n59_), .Y(mai_mai_n276_));
  NA2        m254(.A(mai_mai_n276_), .B(x02), .Y(mai_mai_n277_));
  NA2        m255(.A(mai_mai_n165_), .B(x04), .Y(mai_mai_n278_));
  INV        m256(.A(mai_mai_n278_), .Y(mai_mai_n279_));
  NO3        m257(.A(mai_mai_n156_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n280_));
  OAI210     m258(.A0(mai_mai_n280_), .A1(mai_mai_n279_), .B0(mai_mai_n93_), .Y(mai_mai_n281_));
  NO3        m259(.A(mai_mai_n165_), .B(mai_mai_n142_), .C(mai_mai_n52_), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n127_), .A1(mai_mai_n36_), .B0(mai_mai_n98_), .Y(mai_mai_n283_));
  OAI210     m261(.A0(mai_mai_n283_), .A1(mai_mai_n164_), .B0(mai_mai_n282_), .Y(mai_mai_n284_));
  NA4        m262(.A(mai_mai_n284_), .B(mai_mai_n281_), .C(mai_mai_n277_), .D(x06), .Y(mai_mai_n285_));
  NA2        m263(.A(x09), .B(x03), .Y(mai_mai_n286_));
  OAI220     m264(.A0(mai_mai_n286_), .A1(mai_mai_n115_), .B0(mai_mai_n171_), .B1(mai_mai_n64_), .Y(mai_mai_n287_));
  OAI220     m265(.A0(mai_mai_n143_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n288_));
  NA2        m266(.A(mai_mai_n288_), .B(mai_mai_n183_), .Y(mai_mai_n289_));
  NO2        m267(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n290_));
  NA2        m268(.A(mai_mai_n282_), .B(mai_mai_n290_), .Y(mai_mai_n291_));
  OAI210     m269(.A0(mai_mai_n289_), .A1(mai_mai_n28_), .B0(mai_mai_n291_), .Y(mai_mai_n292_));
  AO220      m270(.A0(mai_mai_n292_), .A1(x04), .B0(mai_mai_n287_), .B1(x05), .Y(mai_mai_n293_));
  AOI210     m271(.A0(mai_mai_n285_), .A1(mai_mai_n272_), .B0(mai_mai_n293_), .Y(mai_mai_n294_));
  OAI210     m272(.A0(mai_mai_n263_), .A1(x12), .B0(mai_mai_n294_), .Y(mai03));
  OR2        m273(.A(mai_mai_n42_), .B(mai_mai_n184_), .Y(mai_mai_n296_));
  AOI210     m274(.A0(mai_mai_n133_), .A1(mai_mai_n98_), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  OAI210     m275(.A0(mai_mai_n375_), .A1(mai_mai_n297_), .B0(x05), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n296_), .B(x05), .Y(mai_mai_n299_));
  AOI210     m277(.A0(mai_mai_n121_), .A1(mai_mai_n177_), .B0(mai_mai_n299_), .Y(mai_mai_n300_));
  AOI210     m278(.A0(mai_mai_n185_), .A1(mai_mai_n80_), .B0(mai_mai_n110_), .Y(mai_mai_n301_));
  OAI220     m279(.A0(mai_mai_n301_), .A1(mai_mai_n59_), .B0(mai_mai_n254_), .B1(mai_mai_n246_), .Y(mai_mai_n302_));
  OAI210     m280(.A0(mai_mai_n302_), .A1(mai_mai_n300_), .B0(mai_mai_n98_), .Y(mai_mai_n303_));
  NO2        m281(.A(mai_mai_n128_), .B(x13), .Y(mai_mai_n304_));
  NA2        m282(.A(mai_mai_n304_), .B(x04), .Y(mai_mai_n305_));
  AOI210     m283(.A0(mai_mai_n160_), .A1(mai_mai_n98_), .B0(mai_mai_n125_), .Y(mai_mai_n306_));
  OA210      m284(.A0(mai_mai_n144_), .A1(x12), .B0(mai_mai_n118_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n307_), .B(mai_mai_n306_), .Y(mai_mai_n308_));
  NA4        m286(.A(mai_mai_n308_), .B(mai_mai_n305_), .C(mai_mai_n303_), .D(mai_mai_n298_), .Y(mai04));
  NO2        m287(.A(mai_mai_n88_), .B(mai_mai_n39_), .Y(mai_mai_n310_));
  XO2        m288(.A(mai_mai_n310_), .B(mai_mai_n204_), .Y(mai05));
  INV        m289(.A(mai_mai_n174_), .Y(mai_mai_n312_));
  AOI210     m290(.A0(mai_mai_n312_), .A1(mai_mai_n253_), .B0(mai_mai_n25_), .Y(mai_mai_n313_));
  NA3        m291(.A(mai_mai_n123_), .B(mai_mai_n117_), .C(mai_mai_n31_), .Y(mai_mai_n314_));
  NO2        m292(.A(mai_mai_n314_), .B(mai_mai_n24_), .Y(mai_mai_n315_));
  OAI210     m293(.A0(mai_mai_n315_), .A1(mai_mai_n313_), .B0(mai_mai_n98_), .Y(mai_mai_n316_));
  NA2        m294(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n317_));
  NA2        m295(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n318_));
  NA2        m296(.A(mai_mai_n209_), .B(x03), .Y(mai_mai_n319_));
  OAI220     m297(.A0(mai_mai_n319_), .A1(mai_mai_n318_), .B0(mai_mai_n317_), .B1(mai_mai_n81_), .Y(mai_mai_n320_));
  OAI210     m298(.A0(mai_mai_n26_), .A1(mai_mai_n98_), .B0(x07), .Y(mai_mai_n321_));
  AOI210     m299(.A0(mai_mai_n320_), .A1(x06), .B0(mai_mai_n321_), .Y(mai_mai_n322_));
  AOI220     m300(.A0(mai_mai_n81_), .A1(mai_mai_n31_), .B0(mai_mai_n52_), .B1(mai_mai_n51_), .Y(mai_mai_n323_));
  NO3        m301(.A(mai_mai_n323_), .B(mai_mai_n23_), .C(x00), .Y(mai_mai_n324_));
  INV        m302(.A(mai_mai_n212_), .Y(mai_mai_n325_));
  OR2        m303(.A(mai_mai_n325_), .B(mai_mai_n196_), .Y(mai_mai_n326_));
  NO2        m304(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n327_));
  OAI210     m305(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n328_));
  OR3        m306(.A(mai_mai_n328_), .B(mai_mai_n327_), .C(mai_mai_n44_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n329_), .B(mai_mai_n326_), .Y(mai_mai_n330_));
  OAI210     m308(.A0(mai_mai_n330_), .A1(mai_mai_n324_), .B0(mai_mai_n98_), .Y(mai_mai_n331_));
  NA2        m309(.A(mai_mai_n33_), .B(mai_mai_n98_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(mai_mai_n332_), .A1(mai_mai_n90_), .B0(x07), .Y(mai_mai_n333_));
  AOI220     m311(.A0(mai_mai_n333_), .A1(mai_mai_n331_), .B0(mai_mai_n322_), .B1(mai_mai_n316_), .Y(mai_mai_n334_));
  AOI210     m312(.A0(mai_mai_n327_), .A1(mai_mai_n75_), .B0(mai_mai_n122_), .Y(mai_mai_n335_));
  OR2        m313(.A(mai_mai_n335_), .B(x03), .Y(mai_mai_n336_));
  NA2        m314(.A(mai_mai_n290_), .B(mai_mai_n61_), .Y(mai_mai_n337_));
  NO2        m315(.A(mai_mai_n337_), .B(x11), .Y(mai_mai_n338_));
  NO3        m316(.A(mai_mai_n338_), .B(mai_mai_n124_), .C(mai_mai_n28_), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n339_), .A1(mai_mai_n336_), .B0(mai_mai_n47_), .Y(mai_mai_n340_));
  NA2        m318(.A(mai_mai_n340_), .B(mai_mai_n99_), .Y(mai_mai_n341_));
  AOI210     m319(.A0(mai_mai_n278_), .A1(mai_mai_n105_), .B0(mai_mai_n217_), .Y(mai_mai_n342_));
  NOi21      m320(.An(mai_mai_n264_), .B(mai_mai_n118_), .Y(mai_mai_n343_));
  NO2        m321(.A(mai_mai_n343_), .B(mai_mai_n218_), .Y(mai_mai_n344_));
  OAI210     m322(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n345_));
  AOI210     m323(.A0(mai_mai_n204_), .A1(mai_mai_n47_), .B0(mai_mai_n345_), .Y(mai_mai_n346_));
  NO4        m324(.A(mai_mai_n346_), .B(mai_mai_n344_), .C(mai_mai_n342_), .D(x08), .Y(mai_mai_n347_));
  NO2        m325(.A(mai_mai_n117_), .B(mai_mai_n28_), .Y(mai_mai_n348_));
  NO2        m326(.A(mai_mai_n348_), .B(mai_mai_n222_), .Y(mai_mai_n349_));
  NA3        m327(.A(mai_mai_n273_), .B(mai_mai_n111_), .C(x12), .Y(mai_mai_n350_));
  AO210      m328(.A0(mai_mai_n273_), .A1(mai_mai_n111_), .B0(mai_mai_n204_), .Y(mai_mai_n351_));
  NA3        m329(.A(mai_mai_n351_), .B(mai_mai_n350_), .C(x08), .Y(mai_mai_n352_));
  INV        m330(.A(mai_mai_n352_), .Y(mai_mai_n353_));
  AOI210     m331(.A0(mai_mai_n347_), .A1(mai_mai_n341_), .B0(mai_mai_n353_), .Y(mai_mai_n354_));
  OAI210     m332(.A0(mai_mai_n337_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n355_));
  NA2        m333(.A(mai_mai_n240_), .B(x07), .Y(mai_mai_n356_));
  OAI220     m334(.A0(mai_mai_n356_), .A1(mai_mai_n318_), .B0(mai_mai_n124_), .B1(mai_mai_n43_), .Y(mai_mai_n357_));
  OAI210     m335(.A0(mai_mai_n357_), .A1(mai_mai_n355_), .B0(mai_mai_n159_), .Y(mai_mai_n358_));
  NA3        m336(.A(mai_mai_n349_), .B(mai_mai_n343_), .C(mai_mai_n269_), .Y(mai_mai_n359_));
  INV        m337(.A(x14), .Y(mai_mai_n360_));
  NO3        m338(.A(mai_mai_n264_), .B(mai_mai_n101_), .C(x11), .Y(mai_mai_n361_));
  NO2        m339(.A(mai_mai_n361_), .B(mai_mai_n360_), .Y(mai_mai_n362_));
  NA3        m340(.A(mai_mai_n362_), .B(mai_mai_n359_), .C(mai_mai_n358_), .Y(mai_mai_n363_));
  AOI220     m341(.A0(mai_mai_n332_), .A1(mai_mai_n61_), .B0(mai_mai_n348_), .B1(mai_mai_n142_), .Y(mai_mai_n364_));
  NOi21      m342(.An(mai_mai_n226_), .B(mai_mai_n128_), .Y(mai_mai_n365_));
  NA2        m343(.A(mai_mai_n230_), .B(mai_mai_n188_), .Y(mai_mai_n366_));
  OAI210     m344(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n366_), .Y(mai_mai_n367_));
  OAI210     m345(.A0(mai_mai_n367_), .A1(mai_mai_n365_), .B0(mai_mai_n98_), .Y(mai_mai_n368_));
  OAI210     m346(.A0(mai_mai_n364_), .A1(mai_mai_n89_), .B0(mai_mai_n368_), .Y(mai_mai_n369_));
  NO4        m347(.A(mai_mai_n369_), .B(mai_mai_n363_), .C(mai_mai_n354_), .D(mai_mai_n334_), .Y(mai06));
  INV        m348(.A(x07), .Y(mai_mai_n373_));
  INV        m349(.A(mai_mai_n91_), .Y(mai_mai_n374_));
  INV        m350(.A(mai_mai_n278_), .Y(mai_mai_n375_));
  INV        m351(.A(x09), .Y(mai_mai_n376_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NO3        u026(.A(x02), .B(x11), .C(x09), .Y(men_men_n49_));
  INV        u027(.A(x09), .Y(men_men_n50_));
  NO2        u028(.A(x10), .B(x02), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x07), .Y(men_men_n52_));
  OAI210     u030(.A0(men_men_n52_), .A1(men_men_n49_), .B0(men_men_n47_), .Y(men_men_n53_));
  NOi21      u031(.An(x01), .B(x09), .Y(men_men_n54_));
  INV        u032(.A(x00), .Y(men_men_n55_));
  NO2        u033(.A(men_men_n50_), .B(men_men_n55_), .Y(men_men_n56_));
  NO2        u034(.A(men_men_n56_), .B(men_men_n54_), .Y(men_men_n57_));
  NA2        u035(.A(x09), .B(men_men_n55_), .Y(men_men_n58_));
  INV        u036(.A(x07), .Y(men_men_n59_));
  INV        u037(.A(men_men_n57_), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n29_), .B(x02), .Y(men_men_n61_));
  OAI210     u039(.A0(men_men_n23_), .A1(men_men_n60_), .B0(men_men_n58_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n62_), .B(men_men_n31_), .Y(men_men_n63_));
  AOI210     u041(.A0(men_men_n63_), .A1(men_men_n53_), .B0(x05), .Y(men_men_n64_));
  NA2        u042(.A(x10), .B(x09), .Y(men_men_n65_));
  NA2        u043(.A(x09), .B(x05), .Y(men_men_n66_));
  NA2        u044(.A(x10), .B(x06), .Y(men_men_n67_));
  NO2        u045(.A(men_men_n59_), .B(men_men_n41_), .Y(men_men_n68_));
  NA2        u046(.A(x11), .B(x03), .Y(men_men_n69_));
  NOi31      u047(.An(x08), .B(x04), .C(x00), .Y(men_men_n70_));
  NO2        u048(.A(x10), .B(x09), .Y(men_men_n71_));
  NO2        u049(.A(x09), .B(men_men_n41_), .Y(men_men_n72_));
  NO2        u050(.A(men_men_n72_), .B(men_men_n36_), .Y(men_men_n73_));
  OAI210     u051(.A0(men_men_n72_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n74_));
  NO2        u052(.A(men_men_n36_), .B(x00), .Y(men_men_n75_));
  NO2        u053(.A(x08), .B(x01), .Y(men_men_n76_));
  OAI210     u054(.A0(men_men_n76_), .A1(men_men_n75_), .B0(men_men_n35_), .Y(men_men_n77_));
  NA2        u055(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n77_), .B(x02), .Y(men_men_n79_));
  AN2        u057(.A(men_men_n79_), .B(men_men_n69_), .Y(men_men_n80_));
  INV        u058(.A(men_men_n77_), .Y(men_men_n81_));
  NO2        u059(.A(x06), .B(x05), .Y(men_men_n82_));
  NA2        u060(.A(x11), .B(x00), .Y(men_men_n83_));
  NO2        u061(.A(x11), .B(men_men_n47_), .Y(men_men_n84_));
  NOi21      u062(.An(men_men_n83_), .B(men_men_n84_), .Y(men_men_n85_));
  AOI210     u063(.A0(men_men_n82_), .A1(men_men_n81_), .B0(men_men_n85_), .Y(men_men_n86_));
  NOi21      u064(.An(x01), .B(x10), .Y(men_men_n87_));
  NO2        u065(.A(men_men_n29_), .B(men_men_n55_), .Y(men_men_n88_));
  NO3        u066(.A(men_men_n88_), .B(men_men_n87_), .C(x06), .Y(men_men_n89_));
  NA2        u067(.A(men_men_n89_), .B(men_men_n27_), .Y(men_men_n90_));
  OAI210     u068(.A0(men_men_n86_), .A1(x07), .B0(men_men_n90_), .Y(men_men_n91_));
  NO3        u069(.A(men_men_n91_), .B(men_men_n80_), .C(men_men_n64_), .Y(men01));
  INV        u070(.A(x12), .Y(men_men_n93_));
  INV        u071(.A(x13), .Y(men_men_n94_));
  NA2        u072(.A(men_men_n82_), .B(x01), .Y(men_men_n95_));
  NA2        u073(.A(men_men_n95_), .B(men_men_n65_), .Y(men_men_n96_));
  NA2        u074(.A(x08), .B(x04), .Y(men_men_n97_));
  NO2        u075(.A(men_men_n97_), .B(men_men_n55_), .Y(men_men_n98_));
  NA2        u076(.A(men_men_n98_), .B(men_men_n96_), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n87_), .B(men_men_n28_), .Y(men_men_n100_));
  NO2        u078(.A(men_men_n100_), .B(men_men_n66_), .Y(men_men_n101_));
  NO2        u079(.A(x10), .B(x01), .Y(men_men_n102_));
  NO2        u080(.A(men_men_n29_), .B(x00), .Y(men_men_n103_));
  NO2        u081(.A(men_men_n103_), .B(men_men_n102_), .Y(men_men_n104_));
  NA2        u082(.A(x04), .B(men_men_n28_), .Y(men_men_n105_));
  NO3        u083(.A(men_men_n105_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n106_));
  AOI210     u084(.A0(men_men_n106_), .A1(men_men_n104_), .B0(men_men_n101_), .Y(men_men_n107_));
  AOI210     u085(.A0(men_men_n107_), .A1(men_men_n99_), .B0(men_men_n94_), .Y(men_men_n108_));
  NO2        u086(.A(men_men_n54_), .B(x05), .Y(men_men_n109_));
  NOi21      u087(.An(men_men_n109_), .B(men_men_n56_), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n35_), .B(x02), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n94_), .B(men_men_n36_), .Y(men_men_n112_));
  NA3        u090(.A(men_men_n112_), .B(men_men_n111_), .C(x06), .Y(men_men_n113_));
  NO2        u091(.A(men_men_n113_), .B(men_men_n110_), .Y(men_men_n114_));
  NA2        u092(.A(x09), .B(men_men_n35_), .Y(men_men_n115_));
  INV        u093(.A(men_men_n115_), .Y(men_men_n116_));
  NA2        u094(.A(x13), .B(men_men_n35_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n117_), .B(x05), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n118_), .B(men_men_n116_), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n35_), .B(men_men_n55_), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n120_), .B(men_men_n94_), .Y(men_men_n121_));
  AOI210     u099(.A0(men_men_n121_), .A1(men_men_n73_), .B0(men_men_n110_), .Y(men_men_n122_));
  AOI210     u100(.A0(men_men_n122_), .A1(men_men_n119_), .B0(men_men_n67_), .Y(men_men_n123_));
  NA2        u101(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n124_));
  NA2        u102(.A(x10), .B(men_men_n55_), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n125_), .B(men_men_n124_), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n50_), .B(x05), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n36_), .B(x04), .Y(men_men_n128_));
  NA3        u106(.A(men_men_n128_), .B(men_men_n127_), .C(x13), .Y(men_men_n129_));
  NO3        u107(.A(men_men_n120_), .B(men_men_n72_), .C(men_men_n36_), .Y(men_men_n130_));
  NO2        u108(.A(men_men_n58_), .B(x05), .Y(men_men_n131_));
  NOi41      u109(.An(men_men_n129_), .B(men_men_n131_), .C(men_men_n130_), .D(men_men_n126_), .Y(men_men_n132_));
  NO3        u110(.A(men_men_n132_), .B(x06), .C(x03), .Y(men_men_n133_));
  NO4        u111(.A(men_men_n133_), .B(men_men_n123_), .C(men_men_n114_), .D(men_men_n108_), .Y(men_men_n134_));
  NA2        u112(.A(x13), .B(men_men_n36_), .Y(men_men_n135_));
  OAI210     u113(.A0(men_men_n76_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n136_));
  NA2        u114(.A(men_men_n136_), .B(men_men_n135_), .Y(men_men_n137_));
  NO2        u115(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n138_));
  OA210      u116(.A0(x00), .A1(men_men_n71_), .B0(men_men_n138_), .Y(men_men_n139_));
  NO2        u117(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n140_));
  NA2        u118(.A(men_men_n29_), .B(x06), .Y(men_men_n141_));
  OA210      u119(.A0(men_men_n28_), .A1(men_men_n139_), .B0(men_men_n137_), .Y(men_men_n142_));
  NO2        u120(.A(x09), .B(x05), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n143_), .B(men_men_n47_), .Y(men_men_n144_));
  AOI210     u122(.A0(men_men_n144_), .A1(men_men_n104_), .B0(x02), .Y(men_men_n145_));
  NA2        u123(.A(x09), .B(x00), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n109_), .B(men_men_n146_), .Y(men_men_n147_));
  NO2        u125(.A(men_men_n145_), .B(men_men_n142_), .Y(men_men_n148_));
  NO2        u126(.A(x03), .B(x02), .Y(men_men_n149_));
  NA2        u127(.A(men_men_n77_), .B(men_men_n94_), .Y(men_men_n150_));
  OAI210     u128(.A0(men_men_n150_), .A1(men_men_n110_), .B0(men_men_n149_), .Y(men_men_n151_));
  OA210      u129(.A0(men_men_n148_), .A1(x11), .B0(men_men_n151_), .Y(men_men_n152_));
  OAI210     u130(.A0(men_men_n134_), .A1(men_men_n23_), .B0(men_men_n152_), .Y(men_men_n153_));
  NAi21      u131(.An(x06), .B(x10), .Y(men_men_n154_));
  NOi21      u132(.An(x01), .B(x13), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  OR2        u134(.A(men_men_n156_), .B(x08), .Y(men_men_n157_));
  NO2        u135(.A(men_men_n157_), .B(men_men_n41_), .Y(men_men_n158_));
  NO2        u136(.A(men_men_n29_), .B(x03), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n94_), .B(x01), .Y(men_men_n160_));
  NO2        u138(.A(men_men_n160_), .B(x08), .Y(men_men_n161_));
  OAI210     u139(.A0(x05), .A1(men_men_n161_), .B0(men_men_n50_), .Y(men_men_n162_));
  AOI210     u140(.A0(men_men_n162_), .A1(men_men_n159_), .B0(men_men_n48_), .Y(men_men_n163_));
  AOI210     u141(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n164_));
  OAI210     u142(.A0(men_men_n163_), .A1(men_men_n158_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u143(.A(x04), .B(x02), .Y(men_men_n166_));
  NA2        u144(.A(x10), .B(x05), .Y(men_men_n167_));
  NA2        u145(.A(x09), .B(x06), .Y(men_men_n168_));
  NO2        u146(.A(x09), .B(x01), .Y(men_men_n169_));
  NO3        u147(.A(men_men_n169_), .B(men_men_n102_), .C(men_men_n31_), .Y(men_men_n170_));
  NA2        u148(.A(men_men_n170_), .B(x00), .Y(men_men_n171_));
  NO2        u149(.A(men_men_n109_), .B(x08), .Y(men_men_n172_));
  NA3        u150(.A(men_men_n155_), .B(men_men_n154_), .C(men_men_n50_), .Y(men_men_n173_));
  NA2        u151(.A(men_men_n87_), .B(x05), .Y(men_men_n174_));
  OAI210     u152(.A0(men_men_n174_), .A1(men_men_n112_), .B0(men_men_n173_), .Y(men_men_n175_));
  AOI210     u153(.A0(men_men_n172_), .A1(x06), .B0(men_men_n175_), .Y(men_men_n176_));
  OAI210     u154(.A0(men_men_n176_), .A1(x11), .B0(men_men_n171_), .Y(men_men_n177_));
  NAi21      u155(.An(men_men_n166_), .B(men_men_n177_), .Y(men_men_n178_));
  INV        u156(.A(men_men_n25_), .Y(men_men_n179_));
  NAi21      u157(.An(x13), .B(x00), .Y(men_men_n180_));
  AOI210     u158(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n180_), .Y(men_men_n181_));
  AOI220     u159(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n182_));
  OAI210     u160(.A0(men_men_n167_), .A1(men_men_n35_), .B0(men_men_n182_), .Y(men_men_n183_));
  AN2        u161(.A(men_men_n183_), .B(men_men_n181_), .Y(men_men_n184_));
  AN2        u162(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n185_));
  NO2        u163(.A(men_men_n88_), .B(x06), .Y(men_men_n186_));
  NO2        u164(.A(men_men_n180_), .B(men_men_n36_), .Y(men_men_n187_));
  INV        u165(.A(men_men_n187_), .Y(men_men_n188_));
  OAI220     u166(.A0(men_men_n188_), .A1(men_men_n168_), .B0(men_men_n186_), .B1(men_men_n185_), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n189_), .A1(men_men_n184_), .B0(men_men_n179_), .Y(men_men_n190_));
  NOi21      u168(.An(x09), .B(x00), .Y(men_men_n191_));
  NO3        u169(.A(men_men_n75_), .B(men_men_n191_), .C(men_men_n47_), .Y(men_men_n192_));
  NA2        u170(.A(men_men_n192_), .B(men_men_n125_), .Y(men_men_n193_));
  NA2        u171(.A(x10), .B(x08), .Y(men_men_n194_));
  INV        u172(.A(men_men_n194_), .Y(men_men_n195_));
  NA2        u173(.A(x06), .B(x05), .Y(men_men_n196_));
  OAI210     u174(.A0(men_men_n196_), .A1(men_men_n35_), .B0(men_men_n93_), .Y(men_men_n197_));
  AOI210     u175(.A0(men_men_n195_), .A1(men_men_n56_), .B0(men_men_n197_), .Y(men_men_n198_));
  NA2        u176(.A(men_men_n198_), .B(men_men_n193_), .Y(men_men_n199_));
  NO2        u177(.A(men_men_n94_), .B(x12), .Y(men_men_n200_));
  AOI210     u178(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n200_), .Y(men_men_n201_));
  NA2        u179(.A(men_men_n87_), .B(men_men_n50_), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n203_));
  NA2        u181(.A(men_men_n203_), .B(x02), .Y(men_men_n204_));
  NO2        u182(.A(men_men_n204_), .B(men_men_n202_), .Y(men_men_n205_));
  AOI210     u183(.A0(men_men_n201_), .A1(men_men_n199_), .B0(men_men_n205_), .Y(men_men_n206_));
  NA4        u184(.A(men_men_n206_), .B(men_men_n190_), .C(men_men_n178_), .D(men_men_n165_), .Y(men_men_n207_));
  AOI210     u185(.A0(men_men_n153_), .A1(men_men_n93_), .B0(men_men_n207_), .Y(men_men_n208_));
  NA2        u186(.A(men_men_n28_), .B(men_men_n137_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n50_), .B(men_men_n47_), .Y(men_men_n210_));
  NA2        u188(.A(men_men_n210_), .B(men_men_n136_), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n124_), .B(x06), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n438_), .A1(men_men_n211_), .B0(men_men_n212_), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n213_), .A1(men_men_n209_), .B0(x12), .Y(men_men_n214_));
  INV        u192(.A(men_men_n70_), .Y(men_men_n215_));
  AOI210     u193(.A0(men_men_n194_), .A1(x05), .B0(men_men_n50_), .Y(men_men_n216_));
  OAI210     u194(.A0(men_men_n216_), .A1(men_men_n156_), .B0(men_men_n55_), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n217_), .B(men_men_n215_), .Y(men_men_n218_));
  NO2        u196(.A(men_men_n87_), .B(x06), .Y(men_men_n219_));
  AOI210     u197(.A0(men_men_n36_), .A1(x04), .B0(men_men_n50_), .Y(men_men_n220_));
  NO3        u198(.A(men_men_n220_), .B(men_men_n219_), .C(men_men_n41_), .Y(men_men_n221_));
  NA4        u199(.A(men_men_n154_), .B(men_men_n54_), .C(men_men_n36_), .D(x04), .Y(men_men_n222_));
  NA2        u200(.A(men_men_n222_), .B(men_men_n141_), .Y(men_men_n223_));
  OAI210     u201(.A0(men_men_n223_), .A1(men_men_n221_), .B0(x02), .Y(men_men_n224_));
  AOI210     u202(.A0(men_men_n224_), .A1(men_men_n218_), .B0(men_men_n23_), .Y(men_men_n225_));
  OAI210     u203(.A0(men_men_n214_), .A1(men_men_n55_), .B0(men_men_n225_), .Y(men_men_n226_));
  INV        u204(.A(men_men_n141_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n50_), .B(x03), .Y(men_men_n228_));
  OAI210     u206(.A0(men_men_n72_), .A1(men_men_n36_), .B0(men_men_n115_), .Y(men_men_n229_));
  NO2        u207(.A(men_men_n94_), .B(x03), .Y(men_men_n230_));
  AOI220     u208(.A0(men_men_n230_), .A1(men_men_n229_), .B0(men_men_n70_), .B1(men_men_n228_), .Y(men_men_n231_));
  INV        u209(.A(men_men_n154_), .Y(men_men_n232_));
  NA2        u210(.A(men_men_n232_), .B(men_men_n55_), .Y(men_men_n233_));
  NA2        u211(.A(men_men_n231_), .B(men_men_n233_), .Y(men_men_n234_));
  INV        u212(.A(men_men_n84_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n235_), .B(x12), .Y(men_men_n236_));
  NA2        u214(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n238_));
  OAI210     u216(.A0(men_men_n238_), .A1(men_men_n183_), .B0(men_men_n181_), .Y(men_men_n239_));
  NO2        u217(.A(x06), .B(x00), .Y(men_men_n240_));
  OAI210     u218(.A0(men_men_n97_), .A1(men_men_n146_), .B0(men_men_n67_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n241_), .B(x05), .Y(men_men_n242_));
  NA2        u220(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n243_));
  NA2        u221(.A(men_men_n243_), .B(x03), .Y(men_men_n244_));
  OA210      u222(.A0(men_men_n244_), .A1(men_men_n242_), .B0(men_men_n239_), .Y(men_men_n245_));
  NA2        u223(.A(x13), .B(men_men_n93_), .Y(men_men_n246_));
  NA3        u224(.A(men_men_n246_), .B(men_men_n197_), .C(men_men_n85_), .Y(men_men_n247_));
  OAI210     u225(.A0(men_men_n245_), .A1(men_men_n237_), .B0(men_men_n247_), .Y(men_men_n248_));
  AOI210     u226(.A0(men_men_n236_), .A1(men_men_n234_), .B0(men_men_n248_), .Y(men_men_n249_));
  AOI210     u227(.A0(men_men_n249_), .A1(men_men_n226_), .B0(x07), .Y(men_men_n250_));
  NA2        u228(.A(men_men_n66_), .B(men_men_n29_), .Y(men_men_n251_));
  NO2        u229(.A(men_men_n94_), .B(x06), .Y(men_men_n252_));
  NO2        u230(.A(x08), .B(x05), .Y(men_men_n253_));
  NO2        u231(.A(x12), .B(x02), .Y(men_men_n254_));
  INV        u232(.A(men_men_n254_), .Y(men_men_n255_));
  NO2        u233(.A(men_men_n255_), .B(men_men_n235_), .Y(men_men_n256_));
  OA210      u234(.A0(x13), .A1(men_men_n70_), .B0(men_men_n256_), .Y(men_men_n257_));
  NA2        u235(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n258_));
  NO2        u236(.A(men_men_n258_), .B(x01), .Y(men_men_n259_));
  AOI210     u237(.A0(men_men_n115_), .A1(men_men_n129_), .B0(men_men_n29_), .Y(men_men_n260_));
  NA2        u238(.A(men_men_n252_), .B(men_men_n229_), .Y(men_men_n261_));
  NA2        u239(.A(men_men_n94_), .B(x04), .Y(men_men_n262_));
  NA2        u240(.A(men_men_n262_), .B(men_men_n28_), .Y(men_men_n263_));
  NA2        u241(.A(men_men_n263_), .B(men_men_n261_), .Y(men_men_n264_));
  NO3        u242(.A(men_men_n83_), .B(x12), .C(x03), .Y(men_men_n265_));
  OAI210     u243(.A0(men_men_n264_), .A1(men_men_n260_), .B0(men_men_n265_), .Y(men_men_n266_));
  AOI210     u244(.A0(men_men_n202_), .A1(men_men_n196_), .B0(men_men_n97_), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n25_), .B(x00), .Y(men_men_n268_));
  NA2        u246(.A(men_men_n267_), .B(men_men_n268_), .Y(men_men_n269_));
  NO2        u247(.A(men_men_n56_), .B(x05), .Y(men_men_n270_));
  NO3        u248(.A(men_men_n270_), .B(men_men_n220_), .C(men_men_n186_), .Y(men_men_n271_));
  NO2        u249(.A(men_men_n237_), .B(men_men_n28_), .Y(men_men_n272_));
  OAI210     u250(.A0(men_men_n271_), .A1(men_men_n227_), .B0(men_men_n272_), .Y(men_men_n273_));
  NA3        u251(.A(men_men_n273_), .B(men_men_n269_), .C(men_men_n266_), .Y(men_men_n274_));
  NO3        u252(.A(men_men_n274_), .B(men_men_n257_), .C(men_men_n250_), .Y(men_men_n275_));
  OAI210     u253(.A0(men_men_n208_), .A1(men_men_n59_), .B0(men_men_n275_), .Y(men02));
  NO2        u254(.A(men_men_n77_), .B(men_men_n127_), .Y(men_men_n277_));
  NA3        u255(.A(x13), .B(men_men_n195_), .C(men_men_n54_), .Y(men_men_n278_));
  OAI210     u256(.A0(men_men_n437_), .A1(men_men_n32_), .B0(men_men_n278_), .Y(men_men_n279_));
  OAI210     u257(.A0(men_men_n279_), .A1(men_men_n277_), .B0(men_men_n167_), .Y(men_men_n280_));
  INV        u258(.A(men_men_n167_), .Y(men_men_n281_));
  AOI210     u259(.A0(men_men_n111_), .A1(men_men_n78_), .B0(men_men_n220_), .Y(men_men_n282_));
  NO2        u260(.A(men_men_n282_), .B(men_men_n94_), .Y(men_men_n283_));
  AOI220     u261(.A0(men_men_n283_), .A1(men_men_n281_), .B0(men_men_n150_), .B1(men_men_n149_), .Y(men_men_n284_));
  AOI210     u262(.A0(men_men_n284_), .A1(men_men_n280_), .B0(men_men_n48_), .Y(men_men_n285_));
  NO2        u263(.A(x05), .B(x02), .Y(men_men_n286_));
  OAI210     u264(.A0(men_men_n211_), .A1(men_men_n191_), .B0(men_men_n286_), .Y(men_men_n287_));
  AOI220     u265(.A0(men_men_n253_), .A1(men_men_n56_), .B0(men_men_n54_), .B1(men_men_n36_), .Y(men_men_n288_));
  NOi21      u266(.An(x13), .B(men_men_n288_), .Y(men_men_n289_));
  AOI210     u267(.A0(x13), .A1(men_men_n72_), .B0(men_men_n289_), .Y(men_men_n290_));
  AOI210     u268(.A0(men_men_n290_), .A1(men_men_n287_), .B0(men_men_n141_), .Y(men_men_n291_));
  INV        u269(.A(men_men_n231_), .Y(men_men_n292_));
  NO2        u270(.A(men_men_n243_), .B(men_men_n47_), .Y(men_men_n293_));
  NA2        u271(.A(men_men_n293_), .B(men_men_n292_), .Y(men_men_n294_));
  OAI210     u272(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n295_));
  NA2        u273(.A(x13), .B(men_men_n28_), .Y(men_men_n296_));
  OA210      u274(.A0(men_men_n296_), .A1(x08), .B0(men_men_n144_), .Y(men_men_n297_));
  AOI210     u275(.A0(men_men_n297_), .A1(men_men_n136_), .B0(men_men_n295_), .Y(men_men_n298_));
  NA2        u276(.A(men_men_n298_), .B(men_men_n88_), .Y(men_men_n299_));
  NA2        u277(.A(men_men_n88_), .B(men_men_n228_), .Y(men_men_n300_));
  NA3        u278(.A(men_men_n87_), .B(men_men_n75_), .C(men_men_n42_), .Y(men_men_n301_));
  AOI210     u279(.A0(men_men_n301_), .A1(men_men_n300_), .B0(x04), .Y(men_men_n302_));
  INV        u280(.A(men_men_n100_), .Y(men_men_n303_));
  AOI210     u281(.A0(men_men_n303_), .A1(x13), .B0(men_men_n302_), .Y(men_men_n304_));
  NA3        u282(.A(men_men_n304_), .B(men_men_n299_), .C(men_men_n294_), .Y(men_men_n305_));
  NO3        u283(.A(men_men_n305_), .B(men_men_n291_), .C(men_men_n285_), .Y(men_men_n306_));
  NA2        u284(.A(men_men_n140_), .B(x03), .Y(men_men_n307_));
  INV        u285(.A(men_men_n180_), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n50_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n309_));
  AOI220     u287(.A0(men_men_n309_), .A1(men_men_n308_), .B0(men_men_n203_), .B1(x08), .Y(men_men_n310_));
  OAI210     u288(.A0(men_men_n310_), .A1(men_men_n270_), .B0(men_men_n307_), .Y(men_men_n311_));
  NA2        u289(.A(men_men_n311_), .B(men_men_n102_), .Y(men_men_n312_));
  NA2        u290(.A(men_men_n166_), .B(men_men_n160_), .Y(men_men_n313_));
  AN2        u291(.A(men_men_n313_), .B(men_men_n172_), .Y(men_men_n314_));
  INV        u292(.A(men_men_n54_), .Y(men_men_n315_));
  OAI220     u293(.A0(men_men_n262_), .A1(men_men_n315_), .B0(men_men_n127_), .B1(men_men_n28_), .Y(men_men_n316_));
  OAI210     u294(.A0(men_men_n316_), .A1(men_men_n314_), .B0(men_men_n103_), .Y(men_men_n317_));
  NA2        u295(.A(men_men_n262_), .B(men_men_n93_), .Y(men_men_n318_));
  NA2        u296(.A(men_men_n93_), .B(men_men_n41_), .Y(men_men_n319_));
  NA3        u297(.A(men_men_n319_), .B(men_men_n318_), .C(men_men_n126_), .Y(men_men_n320_));
  NA4        u298(.A(men_men_n320_), .B(men_men_n317_), .C(men_men_n312_), .D(men_men_n48_), .Y(men_men_n321_));
  INV        u299(.A(men_men_n203_), .Y(men_men_n322_));
  NA2        u300(.A(men_men_n32_), .B(x05), .Y(men_men_n323_));
  NA2        u301(.A(men_men_n436_), .B(x02), .Y(men_men_n324_));
  INV        u302(.A(men_men_n238_), .Y(men_men_n325_));
  NA2        u303(.A(men_men_n200_), .B(x04), .Y(men_men_n326_));
  NO2        u304(.A(men_men_n326_), .B(men_men_n325_), .Y(men_men_n327_));
  NO2        u305(.A(x13), .B(men_men_n31_), .Y(men_men_n328_));
  OAI210     u306(.A0(men_men_n328_), .A1(men_men_n327_), .B0(men_men_n88_), .Y(men_men_n329_));
  NO3        u307(.A(men_men_n200_), .B(men_men_n159_), .C(men_men_n51_), .Y(men_men_n330_));
  OAI210     u308(.A0(x12), .A1(men_men_n192_), .B0(men_men_n330_), .Y(men_men_n331_));
  NA4        u309(.A(men_men_n331_), .B(men_men_n329_), .C(men_men_n324_), .D(x06), .Y(men_men_n332_));
  NA2        u310(.A(x09), .B(x03), .Y(men_men_n333_));
  OAI220     u311(.A0(men_men_n333_), .A1(men_men_n125_), .B0(men_men_n210_), .B1(men_men_n61_), .Y(men_men_n334_));
  NO3        u312(.A(men_men_n270_), .B(men_men_n124_), .C(x08), .Y(men_men_n335_));
  AOI210     u313(.A0(x01), .A1(men_men_n227_), .B0(men_men_n335_), .Y(men_men_n336_));
  NO3        u314(.A(men_men_n109_), .B(men_men_n125_), .C(men_men_n38_), .Y(men_men_n337_));
  INV        u315(.A(men_men_n337_), .Y(men_men_n338_));
  OAI210     u316(.A0(men_men_n336_), .A1(men_men_n28_), .B0(men_men_n338_), .Y(men_men_n339_));
  AO220      u317(.A0(men_men_n339_), .A1(x04), .B0(men_men_n334_), .B1(x05), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n332_), .A1(men_men_n321_), .B0(men_men_n340_), .Y(men_men_n341_));
  OAI210     u319(.A0(men_men_n306_), .A1(x12), .B0(men_men_n341_), .Y(men03));
  OR2        u320(.A(men_men_n42_), .B(men_men_n228_), .Y(men_men_n343_));
  AOI210     u321(.A0(men_men_n150_), .A1(men_men_n93_), .B0(men_men_n343_), .Y(men_men_n344_));
  AO210      u322(.A0(men_men_n325_), .A1(men_men_n78_), .B0(men_men_n326_), .Y(men_men_n345_));
  NA2        u323(.A(men_men_n200_), .B(men_men_n149_), .Y(men_men_n346_));
  NA3        u324(.A(men_men_n346_), .B(men_men_n345_), .C(men_men_n204_), .Y(men_men_n347_));
  OAI210     u325(.A0(men_men_n347_), .A1(men_men_n344_), .B0(x05), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n343_), .B(x05), .Y(men_men_n349_));
  AOI210     u327(.A0(men_men_n136_), .A1(men_men_n215_), .B0(men_men_n349_), .Y(men_men_n350_));
  AOI210     u328(.A0(men_men_n230_), .A1(men_men_n73_), .B0(men_men_n118_), .Y(men_men_n351_));
  OAI220     u329(.A0(men_men_n351_), .A1(men_men_n57_), .B0(men_men_n296_), .B1(men_men_n288_), .Y(men_men_n352_));
  OAI210     u330(.A0(men_men_n352_), .A1(men_men_n350_), .B0(men_men_n93_), .Y(men_men_n353_));
  AOI210     u331(.A0(men_men_n144_), .A1(men_men_n58_), .B0(men_men_n38_), .Y(men_men_n354_));
  NO2        u332(.A(men_men_n169_), .B(men_men_n131_), .Y(men_men_n355_));
  OAI220     u333(.A0(men_men_n355_), .A1(men_men_n37_), .B0(men_men_n147_), .B1(x13), .Y(men_men_n356_));
  OAI210     u334(.A0(men_men_n356_), .A1(men_men_n354_), .B0(x04), .Y(men_men_n357_));
  NO3        u335(.A(men_men_n319_), .B(men_men_n77_), .C(men_men_n57_), .Y(men_men_n358_));
  AOI210     u336(.A0(men_men_n188_), .A1(men_men_n93_), .B0(men_men_n144_), .Y(men_men_n359_));
  OA210      u337(.A0(men_men_n161_), .A1(x12), .B0(men_men_n131_), .Y(men_men_n360_));
  NO3        u338(.A(men_men_n360_), .B(men_men_n359_), .C(men_men_n358_), .Y(men_men_n361_));
  NA4        u339(.A(men_men_n361_), .B(men_men_n357_), .C(men_men_n353_), .D(men_men_n348_), .Y(men04));
  NO2        u340(.A(men_men_n81_), .B(men_men_n39_), .Y(men_men_n363_));
  XO2        u341(.A(men_men_n363_), .B(men_men_n246_), .Y(men05));
  AOI210     u342(.A0(men_men_n66_), .A1(men_men_n51_), .B0(men_men_n212_), .Y(men_men_n365_));
  NO2        u343(.A(men_men_n365_), .B(men_men_n25_), .Y(men_men_n366_));
  NA3        u344(.A(men_men_n141_), .B(men_men_n127_), .C(men_men_n31_), .Y(men_men_n367_));
  AOI210     u345(.A0(men_men_n232_), .A1(men_men_n55_), .B0(men_men_n82_), .Y(men_men_n368_));
  AOI210     u346(.A0(men_men_n368_), .A1(men_men_n367_), .B0(men_men_n24_), .Y(men_men_n369_));
  OAI210     u347(.A0(men_men_n369_), .A1(men_men_n366_), .B0(men_men_n93_), .Y(men_men_n370_));
  NA2        u348(.A(x11), .B(men_men_n31_), .Y(men_men_n371_));
  NA2        u349(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n372_));
  NA2        u350(.A(men_men_n251_), .B(x03), .Y(men_men_n373_));
  OAI220     u351(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n371_), .B1(men_men_n74_), .Y(men_men_n374_));
  OAI210     u352(.A0(men_men_n26_), .A1(men_men_n93_), .B0(x07), .Y(men_men_n375_));
  AOI210     u353(.A0(men_men_n374_), .A1(x06), .B0(men_men_n375_), .Y(men_men_n376_));
  AOI220     u354(.A0(men_men_n74_), .A1(men_men_n31_), .B0(men_men_n51_), .B1(men_men_n50_), .Y(men_men_n377_));
  NO3        u355(.A(men_men_n377_), .B(men_men_n23_), .C(x00), .Y(men_men_n378_));
  NA2        u356(.A(men_men_n65_), .B(x02), .Y(men_men_n379_));
  NA2        u357(.A(men_men_n379_), .B(men_men_n373_), .Y(men_men_n380_));
  OR2        u358(.A(men_men_n380_), .B(men_men_n237_), .Y(men_men_n381_));
  NA2        u359(.A(men_men_n155_), .B(x05), .Y(men_men_n382_));
  NA3        u360(.A(men_men_n382_), .B(men_men_n240_), .C(men_men_n235_), .Y(men_men_n383_));
  NO2        u361(.A(men_men_n23_), .B(x10), .Y(men_men_n384_));
  OAI210     u362(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n385_));
  OR3        u363(.A(men_men_n385_), .B(men_men_n384_), .C(men_men_n44_), .Y(men_men_n386_));
  NA3        u364(.A(men_men_n386_), .B(men_men_n383_), .C(men_men_n381_), .Y(men_men_n387_));
  OAI210     u365(.A0(men_men_n387_), .A1(men_men_n378_), .B0(men_men_n93_), .Y(men_men_n388_));
  AOI210     u366(.A0(x12), .A1(men_men_n84_), .B0(x07), .Y(men_men_n389_));
  AOI220     u367(.A0(men_men_n389_), .A1(men_men_n388_), .B0(men_men_n376_), .B1(men_men_n370_), .Y(men_men_n390_));
  NA3        u368(.A(men_men_n23_), .B(men_men_n59_), .C(men_men_n48_), .Y(men_men_n391_));
  AO210      u369(.A0(men_men_n391_), .A1(men_men_n258_), .B0(men_men_n255_), .Y(men_men_n392_));
  AOI210     u370(.A0(men_men_n384_), .A1(men_men_n68_), .B0(men_men_n140_), .Y(men_men_n393_));
  OR2        u371(.A(men_men_n393_), .B(x03), .Y(men_men_n394_));
  NA2        u372(.A(x05), .B(men_men_n59_), .Y(men_men_n395_));
  NO2        u373(.A(men_men_n395_), .B(x11), .Y(men_men_n396_));
  NO3        u374(.A(men_men_n396_), .B(men_men_n143_), .C(men_men_n28_), .Y(men_men_n397_));
  AOI220     u375(.A0(men_men_n397_), .A1(men_men_n394_), .B0(men_men_n392_), .B1(men_men_n47_), .Y(men_men_n398_));
  NO4        u376(.A(men_men_n319_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n399_));
  OAI210     u377(.A0(men_men_n399_), .A1(men_men_n398_), .B0(men_men_n94_), .Y(men_men_n400_));
  AOI210     u378(.A0(men_men_n326_), .A1(men_men_n105_), .B0(men_men_n254_), .Y(men_men_n401_));
  NOi21      u379(.An(men_men_n307_), .B(men_men_n131_), .Y(men_men_n402_));
  NO2        u380(.A(men_men_n401_), .B(x08), .Y(men_men_n403_));
  AOI210     u381(.A0(men_men_n384_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n404_));
  NA2        u382(.A(x09), .B(men_men_n41_), .Y(men_men_n405_));
  OAI210     u383(.A0(men_men_n405_), .A1(men_men_n404_), .B0(men_men_n371_), .Y(men_men_n406_));
  NO2        u384(.A(x13), .B(x12), .Y(men_men_n407_));
  NO2        u385(.A(men_men_n127_), .B(men_men_n28_), .Y(men_men_n408_));
  NO2        u386(.A(men_men_n408_), .B(men_men_n259_), .Y(men_men_n409_));
  OR3        u387(.A(men_men_n409_), .B(x12), .C(x03), .Y(men_men_n410_));
  NA3        u388(.A(men_men_n322_), .B(men_men_n120_), .C(x12), .Y(men_men_n411_));
  NA3        u389(.A(men_men_n411_), .B(men_men_n410_), .C(x08), .Y(men_men_n412_));
  AOI210     u390(.A0(men_men_n407_), .A1(men_men_n406_), .B0(men_men_n412_), .Y(men_men_n413_));
  AOI210     u391(.A0(men_men_n403_), .A1(men_men_n400_), .B0(men_men_n413_), .Y(men_men_n414_));
  OAI210     u392(.A0(men_men_n395_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n415_));
  NA2        u393(.A(men_men_n281_), .B(x07), .Y(men_men_n416_));
  OAI220     u394(.A0(men_men_n416_), .A1(men_men_n372_), .B0(men_men_n143_), .B1(men_men_n43_), .Y(men_men_n417_));
  OAI210     u395(.A0(men_men_n417_), .A1(men_men_n415_), .B0(men_men_n187_), .Y(men_men_n418_));
  NA3        u396(.A(men_men_n409_), .B(men_men_n402_), .C(men_men_n318_), .Y(men_men_n419_));
  INV        u397(.A(x14), .Y(men_men_n420_));
  NO3        u398(.A(men_men_n307_), .B(men_men_n100_), .C(x11), .Y(men_men_n421_));
  NO3        u399(.A(men_men_n160_), .B(men_men_n68_), .C(men_men_n55_), .Y(men_men_n422_));
  NO3        u400(.A(men_men_n391_), .B(men_men_n319_), .C(men_men_n180_), .Y(men_men_n423_));
  NO4        u401(.A(men_men_n423_), .B(men_men_n422_), .C(men_men_n421_), .D(men_men_n420_), .Y(men_men_n424_));
  NA3        u402(.A(men_men_n424_), .B(men_men_n419_), .C(men_men_n418_), .Y(men_men_n425_));
  AOI220     u403(.A0(x12), .A1(men_men_n59_), .B0(men_men_n408_), .B1(men_men_n159_), .Y(men_men_n426_));
  NOi21      u404(.An(men_men_n262_), .B(men_men_n147_), .Y(men_men_n427_));
  NO3        u405(.A(men_men_n124_), .B(men_men_n24_), .C(x06), .Y(men_men_n428_));
  AOI210     u406(.A0(men_men_n268_), .A1(men_men_n232_), .B0(men_men_n428_), .Y(men_men_n429_));
  OAI210     u407(.A0(men_men_n44_), .A1(x04), .B0(men_men_n429_), .Y(men_men_n430_));
  OAI210     u408(.A0(men_men_n430_), .A1(men_men_n427_), .B0(men_men_n93_), .Y(men_men_n431_));
  OAI210     u409(.A0(men_men_n426_), .A1(men_men_n83_), .B0(men_men_n431_), .Y(men_men_n432_));
  NO4        u410(.A(men_men_n432_), .B(men_men_n425_), .C(men_men_n414_), .D(men_men_n390_), .Y(men06));
  INV        u411(.A(men_men_n323_), .Y(men_men_n436_));
  INV        u412(.A(men_men_n169_), .Y(men_men_n437_));
  INV        u413(.A(x05), .Y(men_men_n438_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule