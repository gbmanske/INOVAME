// Benchmark "top" written by ABC on Thu Jun 20 14:59:19 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n135_,
    new_new_n136_, new_new_n137_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n617_, new_new_n618_,
    new_new_n619_, new_new_n620_, new_new_n621_, new_new_n622_,
    new_new_n623_, new_new_n624_, new_new_n625_, new_new_n626_,
    new_new_n627_, new_new_n628_, new_new_n629_, new_new_n630_,
    new_new_n631_, new_new_n632_, new_new_n633_, new_new_n634_,
    new_new_n635_, new_new_n636_, new_new_n637_, new_new_n638_,
    new_new_n639_, new_new_n640_, new_new_n641_, new_new_n642_,
    new_new_n643_, new_new_n644_, new_new_n645_, new_new_n646_,
    new_new_n647_, new_new_n648_, new_new_n649_, new_new_n650_,
    new_new_n651_, new_new_n652_, new_new_n653_, new_new_n654_,
    new_new_n655_, new_new_n656_, new_new_n657_, new_new_n658_,
    new_new_n659_, new_new_n660_, new_new_n661_, new_new_n662_,
    new_new_n663_, new_new_n665_, new_new_n666_, new_new_n667_,
    new_new_n668_, new_new_n669_, new_new_n670_, new_new_n671_,
    new_new_n672_, new_new_n673_, new_new_n674_, new_new_n675_,
    new_new_n676_, new_new_n677_, new_new_n678_, new_new_n679_,
    new_new_n680_, new_new_n681_, new_new_n682_, new_new_n683_,
    new_new_n684_, new_new_n685_, new_new_n686_, new_new_n687_,
    new_new_n688_, new_new_n689_, new_new_n690_, new_new_n691_,
    new_new_n692_, new_new_n693_, new_new_n694_, new_new_n695_,
    new_new_n696_, new_new_n697_, new_new_n698_, new_new_n699_,
    new_new_n700_, new_new_n701_, new_new_n702_, new_new_n703_,
    new_new_n704_, new_new_n705_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n873_, new_new_n874_, new_new_n875_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n55_));
  NO2        g033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  NAi21      g035(.An(i_2_), .B(i_7_), .Y(new_new_n58_));
  INV        g036(.A(i_1_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_6_), .Y(new_new_n60_));
  NA3        g038(.A(new_new_n60_), .B(new_new_n58_), .C(new_new_n31_), .Y(new_new_n61_));
  NA2        g039(.A(i_1_), .B(i_10_), .Y(new_new_n62_));
  NO2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NAi21      g041(.An(new_new_n63_), .B(new_new_n61_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n50_), .B(i_2_), .Y(new_new_n65_));
  AOI210     g043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_6_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(new_new_n25_), .Y(new_new_n68_));
  INV        g046(.A(i_0_), .Y(new_new_n69_));
  NAi21      g047(.An(i_5_), .B(i_10_), .Y(new_new_n70_));
  NA2        g048(.A(i_5_), .B(i_9_), .Y(new_new_n71_));
  AOI210     g049(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n69_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n72_), .B(new_new_n68_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n66_), .A1(new_new_n65_), .B0(new_new_n73_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n74_), .A1(new_new_n64_), .B0(i_0_), .Y(new_new_n75_));
  NA2        g053(.A(i_12_), .B(i_5_), .Y(new_new_n76_));
  NA2        g054(.A(i_2_), .B(i_8_), .Y(new_new_n77_));
  NO2        g055(.A(new_new_n77_), .B(new_new_n56_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_9_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_7_), .Y(new_new_n80_));
  INV        g058(.A(i_6_), .Y(new_new_n81_));
  OR4        g059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n82_));
  INV        g060(.A(new_new_n82_), .Y(new_new_n83_));
  NO2        g061(.A(i_2_), .B(i_7_), .Y(new_new_n84_));
  NAi21      g062(.An(i_6_), .B(i_10_), .Y(new_new_n85_));
  NA2        g063(.A(i_6_), .B(i_9_), .Y(new_new_n86_));
  AOI210     g064(.A0(new_new_n86_), .A1(new_new_n85_), .B0(new_new_n59_), .Y(new_new_n87_));
  NA2        g065(.A(i_2_), .B(i_6_), .Y(new_new_n88_));
  NO3        g066(.A(new_new_n88_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n89_));
  NO2        g067(.A(new_new_n89_), .B(new_new_n87_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n874_), .B0(new_new_n76_), .Y(new_new_n91_));
  AN3        g069(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n92_));
  NAi21      g070(.An(i_6_), .B(i_11_), .Y(new_new_n93_));
  NO2        g071(.A(i_5_), .B(i_8_), .Y(new_new_n94_));
  NOi21      g072(.An(new_new_n94_), .B(new_new_n93_), .Y(new_new_n95_));
  AOI220     g073(.A0(new_new_n95_), .A1(new_new_n58_), .B0(new_new_n92_), .B1(new_new_n32_), .Y(new_new_n96_));
  INV        g074(.A(i_7_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n46_), .B(new_new_n97_), .Y(new_new_n98_));
  NO2        g076(.A(i_0_), .B(i_5_), .Y(new_new_n99_));
  NO2        g077(.A(new_new_n99_), .B(new_new_n81_), .Y(new_new_n100_));
  NA2        g078(.A(i_12_), .B(i_3_), .Y(new_new_n101_));
  INV        g079(.A(new_new_n101_), .Y(new_new_n102_));
  NA3        g080(.A(new_new_n102_), .B(new_new_n100_), .C(new_new_n98_), .Y(new_new_n103_));
  NAi21      g081(.An(i_7_), .B(i_11_), .Y(new_new_n104_));
  NO3        g082(.A(new_new_n104_), .B(new_new_n85_), .C(new_new_n53_), .Y(new_new_n105_));
  AN2        g083(.A(i_2_), .B(i_10_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(i_7_), .Y(new_new_n107_));
  OR2        g085(.A(new_new_n76_), .B(new_new_n56_), .Y(new_new_n108_));
  NO2        g086(.A(i_8_), .B(new_new_n97_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n108_), .C(new_new_n107_), .Y(new_new_n110_));
  NA2        g088(.A(i_12_), .B(i_7_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n59_), .B(new_new_n26_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n112_), .B(i_0_), .Y(new_new_n113_));
  NA2        g091(.A(i_11_), .B(i_12_), .Y(new_new_n114_));
  OAI210     g092(.A0(new_new_n113_), .A1(new_new_n111_), .B0(new_new_n114_), .Y(new_new_n115_));
  NO2        g093(.A(new_new_n115_), .B(new_new_n110_), .Y(new_new_n116_));
  NAi41      g094(.An(new_new_n105_), .B(new_new_n116_), .C(new_new_n103_), .D(new_new_n96_), .Y(new_new_n117_));
  NOi21      g095(.An(i_1_), .B(i_5_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n118_), .B(i_11_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n120_));
  NA2        g098(.A(i_7_), .B(new_new_n25_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n121_), .B(new_new_n120_), .Y(new_new_n122_));
  NO2        g100(.A(new_new_n122_), .B(new_new_n46_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n86_), .B(new_new_n85_), .Y(new_new_n124_));
  NAi21      g102(.An(i_3_), .B(i_8_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n125_), .B(new_new_n58_), .Y(new_new_n126_));
  NOi31      g104(.An(new_new_n126_), .B(new_new_n124_), .C(new_new_n123_), .Y(new_new_n127_));
  NO2        g105(.A(i_1_), .B(new_new_n81_), .Y(new_new_n128_));
  NO2        g106(.A(i_6_), .B(i_5_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n129_), .B(i_3_), .Y(new_new_n130_));
  AO210      g108(.A0(new_new_n130_), .A1(new_new_n47_), .B0(new_new_n128_), .Y(new_new_n131_));
  OAI220     g109(.A0(new_new_n131_), .A1(new_new_n104_), .B0(new_new_n127_), .B1(new_new_n119_), .Y(new_new_n132_));
  NO3        g110(.A(new_new_n132_), .B(new_new_n117_), .C(new_new_n91_), .Y(new_new_n133_));
  NA3        g111(.A(new_new_n133_), .B(new_new_n75_), .C(new_new_n55_), .Y(ori2));
  NO2        g112(.A(new_new_n59_), .B(new_new_n37_), .Y(new_new_n135_));
  NA2        g113(.A(i_6_), .B(new_new_n25_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(new_new_n135_), .Y(new_new_n137_));
  NA4        g115(.A(new_new_n137_), .B(new_new_n73_), .C(new_new_n65_), .D(new_new_n30_), .Y(ori0));
  AN2        g116(.A(i_8_), .B(i_7_), .Y(new_new_n139_));
  NA2        g117(.A(new_new_n139_), .B(i_6_), .Y(new_new_n140_));
  NO2        g118(.A(i_12_), .B(i_13_), .Y(new_new_n141_));
  NAi21      g119(.An(i_5_), .B(i_11_), .Y(new_new_n142_));
  NOi21      g120(.An(new_new_n141_), .B(new_new_n142_), .Y(new_new_n143_));
  NO2        g121(.A(i_0_), .B(i_1_), .Y(new_new_n144_));
  NA2        g122(.A(i_2_), .B(i_3_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(i_4_), .Y(new_new_n146_));
  NA3        g124(.A(new_new_n146_), .B(new_new_n144_), .C(new_new_n143_), .Y(new_new_n147_));
  AN2        g125(.A(new_new_n141_), .B(new_new_n79_), .Y(new_new_n148_));
  NA2        g126(.A(i_1_), .B(i_5_), .Y(new_new_n149_));
  OR2        g127(.A(i_0_), .B(i_1_), .Y(new_new_n150_));
  NO3        g128(.A(new_new_n150_), .B(new_new_n76_), .C(i_13_), .Y(new_new_n151_));
  NAi32      g129(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n152_));
  NAi21      g130(.An(new_new_n152_), .B(new_new_n151_), .Y(new_new_n153_));
  NOi21      g131(.An(i_4_), .B(i_10_), .Y(new_new_n154_));
  NA2        g132(.A(new_new_n154_), .B(new_new_n40_), .Y(new_new_n155_));
  NO2        g133(.A(i_3_), .B(i_5_), .Y(new_new_n156_));
  NO3        g134(.A(new_new_n69_), .B(i_2_), .C(i_1_), .Y(new_new_n157_));
  NA2        g135(.A(new_new_n157_), .B(new_new_n156_), .Y(new_new_n158_));
  OAI210     g136(.A0(new_new_n158_), .A1(new_new_n155_), .B0(new_new_n153_), .Y(new_new_n159_));
  INV        g137(.A(new_new_n159_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n160_), .B(new_new_n140_), .Y(new_new_n161_));
  NOi21      g139(.An(i_4_), .B(i_9_), .Y(new_new_n162_));
  NOi21      g140(.An(i_11_), .B(i_13_), .Y(new_new_n163_));
  NA2        g141(.A(new_new_n163_), .B(new_new_n162_), .Y(new_new_n164_));
  NO2        g142(.A(i_4_), .B(i_5_), .Y(new_new_n165_));
  NAi21      g143(.An(i_12_), .B(i_11_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n69_), .B(new_new_n59_), .Y(new_new_n167_));
  NA2        g145(.A(new_new_n167_), .B(new_new_n46_), .Y(new_new_n168_));
  NA2        g146(.A(new_new_n36_), .B(i_5_), .Y(new_new_n169_));
  NAi31      g147(.An(new_new_n169_), .B(new_new_n148_), .C(i_11_), .Y(new_new_n170_));
  NA2        g148(.A(i_3_), .B(i_5_), .Y(new_new_n171_));
  OR2        g149(.A(new_new_n171_), .B(new_new_n164_), .Y(new_new_n172_));
  AOI210     g150(.A0(new_new_n172_), .A1(new_new_n170_), .B0(new_new_n168_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n69_), .B(i_5_), .Y(new_new_n174_));
  NO2        g152(.A(i_13_), .B(i_10_), .Y(new_new_n175_));
  NA3        g153(.A(new_new_n175_), .B(new_new_n174_), .C(new_new_n44_), .Y(new_new_n176_));
  NO2        g154(.A(i_2_), .B(i_1_), .Y(new_new_n177_));
  NA2        g155(.A(new_new_n177_), .B(i_3_), .Y(new_new_n178_));
  NAi21      g156(.An(i_4_), .B(i_12_), .Y(new_new_n179_));
  INV        g157(.A(new_new_n173_), .Y(new_new_n180_));
  INV        g158(.A(i_8_), .Y(new_new_n181_));
  NO2        g159(.A(new_new_n181_), .B(i_7_), .Y(new_new_n182_));
  NO3        g160(.A(i_3_), .B(new_new_n81_), .C(new_new_n48_), .Y(new_new_n183_));
  NA2        g161(.A(new_new_n183_), .B(new_new_n109_), .Y(new_new_n184_));
  NO3        g162(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n185_));
  NA3        g163(.A(new_new_n185_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n186_));
  NO3        g164(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n186_), .B(new_new_n184_), .Y(new_new_n188_));
  NO2        g166(.A(i_3_), .B(i_8_), .Y(new_new_n189_));
  NO3        g167(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n190_));
  NA3        g168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n40_), .Y(new_new_n191_));
  NO2        g169(.A(new_new_n99_), .B(new_new_n56_), .Y(new_new_n192_));
  INV        g170(.A(new_new_n192_), .Y(new_new_n193_));
  NO2        g171(.A(i_13_), .B(i_9_), .Y(new_new_n194_));
  NAi21      g172(.An(i_12_), .B(i_3_), .Y(new_new_n195_));
  NO2        g173(.A(new_new_n44_), .B(i_5_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n193_), .B(new_new_n191_), .Y(new_new_n197_));
  AOI210     g175(.A0(new_new_n197_), .A1(i_7_), .B0(new_new_n188_), .Y(new_new_n198_));
  OAI220     g176(.A0(new_new_n198_), .A1(i_4_), .B0(i_7_), .B1(new_new_n180_), .Y(new_new_n199_));
  NAi21      g177(.An(i_12_), .B(i_7_), .Y(new_new_n200_));
  NA3        g178(.A(i_13_), .B(new_new_n181_), .C(i_10_), .Y(new_new_n201_));
  NO2        g179(.A(new_new_n201_), .B(new_new_n200_), .Y(new_new_n202_));
  NA2        g180(.A(i_0_), .B(i_5_), .Y(new_new_n203_));
  OAI220     g181(.A0(new_new_n81_), .A1(new_new_n178_), .B0(new_new_n168_), .B1(new_new_n130_), .Y(new_new_n204_));
  NAi31      g182(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n36_), .B(i_13_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n46_), .B(new_new_n59_), .Y(new_new_n207_));
  NA3        g185(.A(new_new_n207_), .B(i_0_), .C(new_new_n206_), .Y(new_new_n208_));
  INV        g186(.A(i_13_), .Y(new_new_n209_));
  NO2        g187(.A(i_12_), .B(new_new_n209_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n208_), .B(new_new_n205_), .Y(new_new_n211_));
  AOI220     g189(.A0(new_new_n211_), .A1(new_new_n139_), .B0(new_new_n204_), .B1(new_new_n202_), .Y(new_new_n212_));
  NO2        g190(.A(i_12_), .B(new_new_n37_), .Y(new_new_n213_));
  OR2        g191(.A(i_8_), .B(i_7_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n53_), .B(i_1_), .Y(new_new_n215_));
  INV        g193(.A(i_12_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n44_), .B(new_new_n216_), .Y(new_new_n217_));
  NO3        g195(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n218_));
  NA2        g196(.A(i_2_), .B(i_1_), .Y(new_new_n219_));
  NO3        g197(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n220_));
  NAi21      g198(.An(i_4_), .B(i_3_), .Y(new_new_n221_));
  NO2        g199(.A(i_0_), .B(i_6_), .Y(new_new_n222_));
  NOi41      g200(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n219_), .B(new_new_n171_), .Y(new_new_n224_));
  NO2        g202(.A(i_11_), .B(new_new_n209_), .Y(new_new_n225_));
  NOi21      g203(.An(i_1_), .B(i_6_), .Y(new_new_n226_));
  NAi21      g204(.An(i_3_), .B(i_7_), .Y(new_new_n227_));
  NA2        g205(.A(new_new_n216_), .B(i_9_), .Y(new_new_n228_));
  OR4        g206(.A(new_new_n228_), .B(new_new_n227_), .C(new_new_n226_), .D(new_new_n174_), .Y(new_new_n229_));
  NO2        g207(.A(i_12_), .B(i_3_), .Y(new_new_n230_));
  NA2        g208(.A(new_new_n69_), .B(i_5_), .Y(new_new_n231_));
  NA2        g209(.A(i_3_), .B(i_9_), .Y(new_new_n232_));
  NAi21      g210(.An(i_7_), .B(i_10_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  NA3        g212(.A(new_new_n234_), .B(new_new_n231_), .C(new_new_n60_), .Y(new_new_n235_));
  NA2        g213(.A(new_new_n235_), .B(new_new_n229_), .Y(new_new_n236_));
  INV        g214(.A(new_new_n140_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n216_), .B(i_13_), .Y(new_new_n238_));
  NO2        g216(.A(new_new_n238_), .B(new_new_n71_), .Y(new_new_n239_));
  AOI220     g217(.A0(new_new_n239_), .A1(new_new_n237_), .B0(new_new_n236_), .B1(new_new_n225_), .Y(new_new_n240_));
  NO2        g218(.A(new_new_n214_), .B(new_new_n37_), .Y(new_new_n241_));
  NA2        g219(.A(i_12_), .B(i_6_), .Y(new_new_n242_));
  OR2        g220(.A(i_13_), .B(i_9_), .Y(new_new_n243_));
  NO3        g221(.A(new_new_n243_), .B(new_new_n242_), .C(new_new_n48_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n221_), .B(i_2_), .Y(new_new_n245_));
  NA3        g223(.A(new_new_n245_), .B(new_new_n244_), .C(new_new_n44_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n225_), .B(i_9_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n231_), .B(new_new_n60_), .Y(new_new_n248_));
  OAI210     g226(.A0(new_new_n248_), .A1(new_new_n247_), .B0(new_new_n246_), .Y(new_new_n249_));
  NO3        g227(.A(i_11_), .B(new_new_n209_), .C(new_new_n25_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n227_), .B(i_8_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n249_), .B(new_new_n241_), .Y(new_new_n252_));
  NA3        g230(.A(new_new_n252_), .B(new_new_n240_), .C(new_new_n212_), .Y(new_new_n253_));
  NO3        g231(.A(i_12_), .B(new_new_n209_), .C(new_new_n37_), .Y(new_new_n254_));
  INV        g232(.A(new_new_n254_), .Y(new_new_n255_));
  NA2        g233(.A(i_8_), .B(new_new_n97_), .Y(new_new_n256_));
  AOI220     g234(.A0(i_2_), .A1(new_new_n183_), .B0(new_new_n156_), .B1(new_new_n215_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n257_), .B(new_new_n256_), .Y(new_new_n258_));
  NO3        g236(.A(i_0_), .B(i_2_), .C(new_new_n59_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n219_), .B(i_0_), .Y(new_new_n260_));
  AOI220     g238(.A0(new_new_n260_), .A1(new_new_n182_), .B0(new_new_n259_), .B1(new_new_n139_), .Y(new_new_n261_));
  NA2        g239(.A(i_5_), .B(new_new_n26_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n262_), .B(new_new_n261_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n57_), .B(i_6_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n158_), .B(new_new_n140_), .Y(new_new_n265_));
  NO3        g243(.A(new_new_n265_), .B(new_new_n263_), .C(new_new_n258_), .Y(new_new_n266_));
  NO2        g244(.A(i_3_), .B(i_10_), .Y(new_new_n267_));
  NO2        g245(.A(i_2_), .B(new_new_n97_), .Y(new_new_n268_));
  AN2        g246(.A(i_3_), .B(i_10_), .Y(new_new_n269_));
  NO2        g247(.A(i_5_), .B(new_new_n37_), .Y(new_new_n270_));
  NO2        g248(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n266_), .B(new_new_n255_), .Y(new_new_n272_));
  NO4        g250(.A(new_new_n272_), .B(new_new_n253_), .C(new_new_n199_), .D(new_new_n161_), .Y(new_new_n273_));
  NO3        g251(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n274_));
  NA2        g252(.A(new_new_n260_), .B(i_7_), .Y(new_new_n275_));
  NO3        g253(.A(i_6_), .B(new_new_n181_), .C(i_7_), .Y(new_new_n276_));
  NA2        g254(.A(new_new_n276_), .B(new_new_n185_), .Y(new_new_n277_));
  AOI210     g255(.A0(new_new_n277_), .A1(new_new_n275_), .B0(i_5_), .Y(new_new_n278_));
  NO2        g256(.A(i_2_), .B(i_3_), .Y(new_new_n279_));
  OR2        g257(.A(i_0_), .B(i_5_), .Y(new_new_n280_));
  NA3        g258(.A(new_new_n260_), .B(new_new_n156_), .C(new_new_n109_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n150_), .B(new_new_n46_), .Y(new_new_n282_));
  INV        g260(.A(new_new_n281_), .Y(new_new_n283_));
  OAI210     g261(.A0(new_new_n283_), .A1(new_new_n278_), .B0(i_4_), .Y(new_new_n284_));
  NO2        g262(.A(i_12_), .B(i_10_), .Y(new_new_n285_));
  NOi21      g263(.An(i_5_), .B(i_0_), .Y(new_new_n286_));
  NO2        g264(.A(i_2_), .B(new_new_n97_), .Y(new_new_n287_));
  NO4        g265(.A(new_new_n287_), .B(i_4_), .C(new_new_n286_), .D(new_new_n125_), .Y(new_new_n288_));
  NA4        g266(.A(new_new_n80_), .B(new_new_n36_), .C(new_new_n81_), .D(i_8_), .Y(new_new_n289_));
  NA2        g267(.A(new_new_n288_), .B(new_new_n285_), .Y(new_new_n290_));
  NO2        g268(.A(i_6_), .B(i_8_), .Y(new_new_n291_));
  NOi21      g269(.An(i_0_), .B(i_2_), .Y(new_new_n292_));
  AN2        g270(.A(new_new_n292_), .B(new_new_n291_), .Y(new_new_n293_));
  NO2        g271(.A(i_1_), .B(i_7_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n290_), .B(new_new_n284_), .Y(new_new_n295_));
  NA3        g273(.A(new_new_n226_), .B(new_new_n268_), .C(new_new_n181_), .Y(new_new_n296_));
  INV        g274(.A(new_new_n88_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n181_), .B(i_9_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n298_), .B(new_new_n192_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n299_), .B(new_new_n46_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n300_), .B(new_new_n263_), .Y(new_new_n301_));
  AOI210     g279(.A0(new_new_n301_), .A1(new_new_n296_), .B0(new_new_n155_), .Y(new_new_n302_));
  AOI210     g280(.A0(new_new_n295_), .A1(new_new_n274_), .B0(new_new_n302_), .Y(new_new_n303_));
  NOi32      g281(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n304_));
  INV        g282(.A(new_new_n304_), .Y(new_new_n305_));
  NAi21      g283(.An(i_0_), .B(i_6_), .Y(new_new_n306_));
  NAi21      g284(.An(i_1_), .B(i_5_), .Y(new_new_n307_));
  NA2        g285(.A(new_new_n307_), .B(new_new_n306_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n308_), .B(new_new_n25_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n309_), .B(new_new_n152_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n152_), .B(new_new_n150_), .Y(new_new_n311_));
  NOi32      g289(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n312_));
  NAi21      g290(.An(i_6_), .B(i_1_), .Y(new_new_n313_));
  NA3        g291(.A(new_new_n313_), .B(new_new_n312_), .C(new_new_n46_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n314_), .B(i_0_), .Y(new_new_n315_));
  OR2        g293(.A(new_new_n315_), .B(new_new_n311_), .Y(new_new_n316_));
  NO2        g294(.A(i_1_), .B(new_new_n97_), .Y(new_new_n317_));
  NAi21      g295(.An(i_3_), .B(i_4_), .Y(new_new_n318_));
  NO2        g296(.A(new_new_n318_), .B(i_9_), .Y(new_new_n319_));
  AN2        g297(.A(i_6_), .B(i_7_), .Y(new_new_n320_));
  OAI210     g298(.A0(new_new_n320_), .A1(new_new_n317_), .B0(new_new_n319_), .Y(new_new_n321_));
  NA2        g299(.A(i_2_), .B(i_7_), .Y(new_new_n322_));
  NO2        g300(.A(new_new_n318_), .B(i_10_), .Y(new_new_n323_));
  NA3        g301(.A(new_new_n323_), .B(new_new_n322_), .C(new_new_n222_), .Y(new_new_n324_));
  AOI210     g302(.A0(new_new_n324_), .A1(new_new_n321_), .B0(new_new_n174_), .Y(new_new_n325_));
  AOI210     g303(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n326_));
  AOI220     g304(.A0(new_new_n323_), .A1(new_new_n294_), .B0(new_new_n218_), .B1(new_new_n177_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n327_), .B(i_5_), .Y(new_new_n328_));
  NO4        g306(.A(new_new_n328_), .B(new_new_n325_), .C(new_new_n316_), .D(new_new_n310_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n329_), .B(new_new_n305_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n331_));
  AN2        g309(.A(i_12_), .B(i_5_), .Y(new_new_n332_));
  NO2        g310(.A(i_4_), .B(new_new_n26_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n333_), .B(new_new_n332_), .Y(new_new_n334_));
  NO2        g312(.A(i_11_), .B(i_6_), .Y(new_new_n335_));
  NA3        g313(.A(new_new_n335_), .B(new_new_n282_), .C(new_new_n209_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n336_), .B(new_new_n334_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n221_), .B(i_5_), .Y(new_new_n338_));
  NO2        g316(.A(i_5_), .B(i_10_), .Y(new_new_n339_));
  AOI220     g317(.A0(new_new_n339_), .A1(new_new_n245_), .B0(new_new_n338_), .B1(new_new_n185_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n141_), .B(new_new_n45_), .Y(new_new_n341_));
  NO2        g319(.A(new_new_n341_), .B(new_new_n340_), .Y(new_new_n342_));
  OAI210     g320(.A0(new_new_n342_), .A1(new_new_n337_), .B0(new_new_n331_), .Y(new_new_n343_));
  NO2        g321(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n147_), .B(new_new_n81_), .Y(new_new_n345_));
  OAI210     g323(.A0(new_new_n345_), .A1(new_new_n337_), .B0(new_new_n344_), .Y(new_new_n346_));
  NO3        g324(.A(new_new_n81_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n347_));
  NA3        g325(.A(new_new_n267_), .B(new_new_n86_), .C(new_new_n71_), .Y(new_new_n348_));
  NO2        g326(.A(i_11_), .B(i_12_), .Y(new_new_n349_));
  NA2        g327(.A(new_new_n349_), .B(new_new_n36_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n348_), .B(new_new_n350_), .Y(new_new_n351_));
  NA2        g329(.A(new_new_n339_), .B(new_new_n216_), .Y(new_new_n352_));
  NAi21      g330(.An(i_13_), .B(i_0_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n353_), .B(new_new_n219_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n351_), .B(new_new_n354_), .Y(new_new_n355_));
  NA3        g333(.A(new_new_n355_), .B(new_new_n346_), .C(new_new_n343_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n44_), .B(new_new_n209_), .Y(new_new_n357_));
  NO2        g335(.A(i_0_), .B(i_11_), .Y(new_new_n358_));
  AN2        g336(.A(i_1_), .B(i_6_), .Y(new_new_n359_));
  NOi21      g337(.An(i_2_), .B(i_12_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n139_), .B(i_9_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n361_), .B(i_4_), .Y(new_new_n362_));
  OR2        g340(.A(i_13_), .B(i_10_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n164_), .B(new_new_n120_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n97_), .B(new_new_n25_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n171_), .B(new_new_n81_), .Y(new_new_n366_));
  NA2        g344(.A(new_new_n181_), .B(i_10_), .Y(new_new_n367_));
  NA3        g345(.A(new_new_n231_), .B(new_new_n60_), .C(i_2_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n264_), .B(new_new_n215_), .Y(new_new_n369_));
  OAI220     g347(.A0(new_new_n369_), .A1(new_new_n171_), .B0(new_new_n368_), .B1(new_new_n367_), .Y(new_new_n370_));
  INV        g348(.A(new_new_n370_), .Y(new_new_n371_));
  AOI210     g349(.A0(new_new_n371_), .A1(new_new_n281_), .B0(new_new_n247_), .Y(new_new_n372_));
  NO3        g350(.A(new_new_n372_), .B(new_new_n356_), .C(new_new_n330_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n69_), .B(i_13_), .Y(new_new_n374_));
  NO2        g352(.A(i_10_), .B(i_9_), .Y(new_new_n375_));
  NAi21      g353(.An(i_12_), .B(i_8_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n376_), .B(i_3_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n46_), .B(i_4_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n378_), .B(new_new_n100_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n191_), .Y(new_new_n380_));
  NA2        g358(.A(new_new_n271_), .B(i_0_), .Y(new_new_n381_));
  NO3        g359(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n242_), .B(new_new_n93_), .Y(new_new_n383_));
  NA2        g361(.A(new_new_n383_), .B(new_new_n382_), .Y(new_new_n384_));
  NA2        g362(.A(i_8_), .B(i_9_), .Y(new_new_n385_));
  AOI210     g363(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n386_));
  OR2        g364(.A(new_new_n386_), .B(new_new_n385_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n254_), .B(new_new_n192_), .Y(new_new_n388_));
  OAI220     g366(.A0(new_new_n388_), .A1(new_new_n387_), .B0(new_new_n384_), .B1(new_new_n381_), .Y(new_new_n389_));
  NO3        g367(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n389_), .B(new_new_n380_), .Y(new_new_n391_));
  OR2        g369(.A(new_new_n299_), .B(new_new_n97_), .Y(new_new_n392_));
  OR2        g370(.A(new_new_n392_), .B(new_new_n155_), .Y(new_new_n393_));
  NA2        g371(.A(new_new_n92_), .B(i_13_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n366_), .B(new_new_n331_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n395_), .B(new_new_n394_), .Y(new_new_n396_));
  NO3        g374(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n397_));
  NO2        g375(.A(i_6_), .B(i_7_), .Y(new_new_n398_));
  NO2        g376(.A(i_11_), .B(i_1_), .Y(new_new_n399_));
  OR2        g377(.A(i_11_), .B(i_8_), .Y(new_new_n400_));
  NOi21      g378(.An(i_2_), .B(i_7_), .Y(new_new_n401_));
  NO2        g379(.A(i_6_), .B(i_10_), .Y(new_new_n402_));
  NA3        g380(.A(new_new_n223_), .B(new_new_n163_), .C(new_new_n129_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n404_));
  NA3        g382(.A(new_new_n344_), .B(new_new_n167_), .C(new_new_n146_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n405_), .B(new_new_n403_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n406_), .B(new_new_n396_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n382_), .B(new_new_n332_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n390_), .B(new_new_n339_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n409_), .B(new_new_n208_), .Y(new_new_n410_));
  NAi21      g388(.An(new_new_n201_), .B(new_new_n349_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n294_), .B(new_new_n203_), .Y(new_new_n412_));
  NO2        g390(.A(new_new_n412_), .B(new_new_n411_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n27_), .B(i_10_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n274_), .B(new_new_n218_), .Y(new_new_n415_));
  OAI220     g393(.A0(new_new_n415_), .A1(new_new_n368_), .B0(new_new_n414_), .B1(new_new_n394_), .Y(new_new_n416_));
  NO3        g394(.A(new_new_n416_), .B(new_new_n413_), .C(new_new_n410_), .Y(new_new_n417_));
  NA4        g395(.A(new_new_n417_), .B(new_new_n407_), .C(new_new_n393_), .D(new_new_n391_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n119_), .B(new_new_n108_), .Y(new_new_n419_));
  AN2        g397(.A(new_new_n419_), .B(new_new_n382_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n420_), .B(new_new_n271_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n304_), .B(new_new_n69_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n320_), .B(new_new_n312_), .Y(new_new_n423_));
  NO2        g401(.A(new_new_n36_), .B(i_8_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n39_), .B(i_13_), .Y(new_new_n425_));
  OAI210     g403(.A0(i_8_), .A1(new_new_n59_), .B0(new_new_n131_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n426_), .B(new_new_n364_), .Y(new_new_n427_));
  NA3        g405(.A(new_new_n427_), .B(new_new_n425_), .C(new_new_n421_), .Y(new_new_n428_));
  NO2        g406(.A(i_12_), .B(new_new_n181_), .Y(new_new_n429_));
  NO2        g407(.A(i_8_), .B(i_7_), .Y(new_new_n430_));
  OAI210     g408(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n431_), .B(new_new_n207_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n432_), .B(new_new_n221_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n44_), .B(i_10_), .Y(new_new_n434_));
  NO2        g412(.A(new_new_n434_), .B(i_6_), .Y(new_new_n435_));
  NA3        g413(.A(new_new_n435_), .B(new_new_n433_), .C(new_new_n430_), .Y(new_new_n436_));
  AOI220     g414(.A0(new_new_n366_), .A1(new_new_n282_), .B0(new_new_n224_), .B1(new_new_n222_), .Y(new_new_n437_));
  OAI220     g415(.A0(new_new_n437_), .A1(new_new_n238_), .B0(new_new_n394_), .B1(new_new_n130_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n438_), .B(new_new_n241_), .Y(new_new_n439_));
  NA3        g417(.A(new_new_n269_), .B(new_new_n165_), .C(new_new_n92_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n206_), .B(new_new_n44_), .Y(new_new_n441_));
  NO2        g419(.A(new_new_n150_), .B(i_5_), .Y(new_new_n442_));
  NA3        g420(.A(new_new_n442_), .B(new_new_n357_), .C(new_new_n279_), .Y(new_new_n443_));
  OAI210     g421(.A0(new_new_n443_), .A1(new_new_n441_), .B0(new_new_n440_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n444_), .B(new_new_n390_), .Y(new_new_n445_));
  NA3        g423(.A(new_new_n445_), .B(new_new_n439_), .C(new_new_n436_), .Y(new_new_n446_));
  AOI210     g424(.A0(new_new_n313_), .A1(new_new_n46_), .B0(new_new_n317_), .Y(new_new_n447_));
  NA2        g425(.A(i_0_), .B(new_new_n48_), .Y(new_new_n448_));
  NA3        g426(.A(new_new_n429_), .B(new_new_n250_), .C(new_new_n448_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n447_), .B(new_new_n449_), .Y(new_new_n450_));
  INV        g428(.A(new_new_n450_), .Y(new_new_n451_));
  NO4        g429(.A(new_new_n226_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n452_));
  NO3        g430(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n453_));
  NO2        g431(.A(new_new_n214_), .B(new_new_n36_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n363_), .B(i_1_), .Y(new_new_n455_));
  NOi31      g433(.An(new_new_n455_), .B(new_new_n383_), .C(new_new_n69_), .Y(new_new_n456_));
  AN4        g434(.A(new_new_n456_), .B(new_new_n362_), .C(i_3_), .D(i_2_), .Y(new_new_n457_));
  INV        g435(.A(new_new_n457_), .Y(new_new_n458_));
  NOi21      g436(.An(i_10_), .B(i_6_), .Y(new_new_n459_));
  NO2        g437(.A(new_new_n81_), .B(new_new_n25_), .Y(new_new_n460_));
  AOI220     g438(.A0(new_new_n254_), .A1(new_new_n460_), .B0(new_new_n250_), .B1(new_new_n459_), .Y(new_new_n461_));
  NO2        g439(.A(new_new_n461_), .B(new_new_n381_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n111_), .B(new_new_n23_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n276_), .B(new_new_n157_), .Y(new_new_n464_));
  AOI220     g442(.A0(new_new_n464_), .A1(new_new_n369_), .B0(new_new_n172_), .B1(new_new_n170_), .Y(new_new_n465_));
  NO2        g443(.A(new_new_n185_), .B(new_new_n37_), .Y(new_new_n466_));
  NOi31      g444(.An(new_new_n143_), .B(new_new_n466_), .C(new_new_n289_), .Y(new_new_n467_));
  NO3        g445(.A(new_new_n467_), .B(new_new_n465_), .C(new_new_n462_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n422_), .B(new_new_n327_), .Y(new_new_n469_));
  INV        g447(.A(new_new_n279_), .Y(new_new_n470_));
  NO2        g448(.A(i_12_), .B(new_new_n81_), .Y(new_new_n471_));
  NA3        g449(.A(new_new_n471_), .B(new_new_n250_), .C(new_new_n448_), .Y(new_new_n472_));
  NA3        g450(.A(new_new_n335_), .B(new_new_n254_), .C(new_new_n203_), .Y(new_new_n473_));
  AOI210     g451(.A0(new_new_n473_), .A1(new_new_n472_), .B0(new_new_n470_), .Y(new_new_n474_));
  OR2        g452(.A(i_2_), .B(i_5_), .Y(new_new_n475_));
  OR2        g453(.A(new_new_n475_), .B(new_new_n359_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n322_), .B(new_new_n222_), .Y(new_new_n477_));
  AOI210     g455(.A0(new_new_n477_), .A1(new_new_n476_), .B0(new_new_n411_), .Y(new_new_n478_));
  NO3        g456(.A(new_new_n478_), .B(new_new_n474_), .C(new_new_n469_), .Y(new_new_n479_));
  NA4        g457(.A(new_new_n479_), .B(new_new_n468_), .C(new_new_n458_), .D(new_new_n451_), .Y(new_new_n480_));
  NO4        g458(.A(new_new_n480_), .B(new_new_n446_), .C(new_new_n428_), .D(new_new_n418_), .Y(new_new_n481_));
  NA4        g459(.A(new_new_n481_), .B(new_new_n373_), .C(new_new_n303_), .D(new_new_n273_), .Y(ori7));
  NO2        g460(.A(new_new_n88_), .B(new_new_n54_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n104_), .B(new_new_n85_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n333_), .B(new_new_n484_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n402_), .B(new_new_n80_), .Y(new_new_n486_));
  NA2        g464(.A(i_11_), .B(new_new_n181_), .Y(new_new_n487_));
  NA2        g465(.A(new_new_n141_), .B(new_new_n487_), .Y(new_new_n488_));
  OAI210     g466(.A0(new_new_n488_), .A1(new_new_n486_), .B0(new_new_n485_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n216_), .B(i_4_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n490_), .B(i_8_), .Y(new_new_n491_));
  NA2        g469(.A(i_2_), .B(new_new_n81_), .Y(new_new_n492_));
  OAI210     g470(.A0(new_new_n84_), .A1(new_new_n189_), .B0(new_new_n190_), .Y(new_new_n493_));
  NO2        g471(.A(i_7_), .B(new_new_n37_), .Y(new_new_n494_));
  NA2        g472(.A(i_4_), .B(i_8_), .Y(new_new_n495_));
  AOI210     g473(.A0(new_new_n495_), .A1(new_new_n269_), .B0(new_new_n494_), .Y(new_new_n496_));
  OAI220     g474(.A0(new_new_n496_), .A1(new_new_n492_), .B0(new_new_n493_), .B1(i_13_), .Y(new_new_n497_));
  NO3        g475(.A(new_new_n497_), .B(new_new_n489_), .C(new_new_n483_), .Y(new_new_n498_));
  AOI210     g476(.A0(new_new_n125_), .A1(new_new_n58_), .B0(i_10_), .Y(new_new_n499_));
  AOI210     g477(.A0(new_new_n499_), .A1(new_new_n216_), .B0(new_new_n154_), .Y(new_new_n500_));
  OR2        g478(.A(i_6_), .B(i_10_), .Y(new_new_n501_));
  OR3        g479(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n502_));
  INV        g480(.A(new_new_n187_), .Y(new_new_n503_));
  OR2        g481(.A(new_new_n500_), .B(new_new_n243_), .Y(new_new_n504_));
  AOI210     g482(.A0(new_new_n504_), .A1(new_new_n498_), .B0(new_new_n59_), .Y(new_new_n505_));
  NOi21      g483(.An(i_11_), .B(i_7_), .Y(new_new_n506_));
  AO210      g484(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(new_new_n506_), .Y(new_new_n508_));
  NA2        g486(.A(new_new_n508_), .B(new_new_n194_), .Y(new_new_n509_));
  NA3        g487(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n510_));
  NAi31      g488(.An(new_new_n510_), .B(new_new_n200_), .C(i_11_), .Y(new_new_n511_));
  AOI210     g489(.A0(new_new_n511_), .A1(new_new_n509_), .B0(new_new_n59_), .Y(new_new_n512_));
  NA2        g490(.A(new_new_n83_), .B(new_new_n59_), .Y(new_new_n513_));
  AO210      g491(.A0(new_new_n513_), .A1(new_new_n327_), .B0(new_new_n41_), .Y(new_new_n514_));
  NO3        g492(.A(new_new_n233_), .B(new_new_n195_), .C(new_new_n487_), .Y(new_new_n515_));
  OAI210     g493(.A0(new_new_n515_), .A1(new_new_n210_), .B0(new_new_n59_), .Y(new_new_n516_));
  NA2        g494(.A(new_new_n360_), .B(new_new_n31_), .Y(new_new_n517_));
  OR2        g495(.A(new_new_n195_), .B(new_new_n104_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n518_), .B(new_new_n517_), .Y(new_new_n519_));
  NO2        g497(.A(i_1_), .B(i_4_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n520_), .B(new_new_n519_), .Y(new_new_n521_));
  NO2        g499(.A(i_1_), .B(i_12_), .Y(new_new_n522_));
  NA3        g500(.A(new_new_n521_), .B(new_new_n516_), .C(new_new_n514_), .Y(new_new_n523_));
  OAI210     g501(.A0(new_new_n523_), .A1(new_new_n512_), .B0(i_6_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n510_), .B(new_new_n104_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n525_), .B(new_new_n471_), .Y(new_new_n526_));
  NO2        g504(.A(i_6_), .B(i_11_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n526_), .B(new_new_n384_), .Y(new_new_n528_));
  NO3        g506(.A(new_new_n501_), .B(new_new_n214_), .C(new_new_n23_), .Y(new_new_n529_));
  AOI210     g507(.A0(i_1_), .A1(new_new_n234_), .B0(new_new_n529_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n530_), .B(new_new_n44_), .Y(new_new_n531_));
  NA3        g509(.A(new_new_n430_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n532_));
  INV        g510(.A(i_2_), .Y(new_new_n533_));
  NA2        g511(.A(new_new_n135_), .B(i_9_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n46_), .B(i_1_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n534_), .B(new_new_n533_), .Y(new_new_n536_));
  AOI210     g514(.A0(new_new_n399_), .A1(new_new_n365_), .B0(new_new_n220_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n537_), .B(new_new_n492_), .Y(new_new_n538_));
  NAi21      g516(.An(new_new_n532_), .B(new_new_n87_), .Y(new_new_n539_));
  NA2        g517(.A(new_new_n535_), .B(new_new_n242_), .Y(new_new_n540_));
  NO2        g518(.A(i_11_), .B(new_new_n37_), .Y(new_new_n541_));
  NA2        g519(.A(new_new_n541_), .B(new_new_n24_), .Y(new_new_n542_));
  OAI210     g520(.A0(new_new_n542_), .A1(new_new_n540_), .B0(new_new_n539_), .Y(new_new_n543_));
  OR3        g521(.A(new_new_n543_), .B(new_new_n538_), .C(new_new_n536_), .Y(new_new_n544_));
  NO3        g522(.A(new_new_n544_), .B(new_new_n531_), .C(new_new_n528_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n216_), .B(new_new_n97_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n546_), .B(new_new_n506_), .Y(new_new_n547_));
  NA2        g525(.A(new_new_n547_), .B(i_1_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n548_), .B(new_new_n502_), .Y(new_new_n549_));
  NA2        g527(.A(new_new_n549_), .B(new_new_n46_), .Y(new_new_n550_));
  NA2        g528(.A(i_3_), .B(new_new_n181_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n551_), .B(new_new_n111_), .Y(new_new_n552_));
  AN2        g530(.A(new_new_n552_), .B(new_new_n435_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n214_), .B(new_new_n44_), .Y(new_new_n554_));
  NO3        g532(.A(new_new_n554_), .B(new_new_n271_), .C(new_new_n217_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n114_), .B(new_new_n37_), .Y(new_new_n556_));
  NO2        g534(.A(new_new_n556_), .B(i_6_), .Y(new_new_n557_));
  NO2        g535(.A(new_new_n81_), .B(i_9_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n558_), .B(new_new_n59_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n559_), .B(new_new_n522_), .Y(new_new_n560_));
  NO4        g538(.A(new_new_n560_), .B(new_new_n557_), .C(new_new_n555_), .D(i_4_), .Y(new_new_n561_));
  NA2        g539(.A(i_1_), .B(i_3_), .Y(new_new_n562_));
  NO2        g540(.A(new_new_n385_), .B(new_new_n88_), .Y(new_new_n563_));
  AOI210     g541(.A0(new_new_n554_), .A1(new_new_n459_), .B0(new_new_n563_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n564_), .B(new_new_n562_), .Y(new_new_n565_));
  NO3        g543(.A(new_new_n565_), .B(new_new_n561_), .C(new_new_n553_), .Y(new_new_n566_));
  NA4        g544(.A(new_new_n566_), .B(new_new_n550_), .C(new_new_n545_), .D(new_new_n524_), .Y(new_new_n567_));
  NO3        g545(.A(new_new_n400_), .B(i_3_), .C(i_7_), .Y(new_new_n568_));
  NOi21      g546(.An(new_new_n568_), .B(i_10_), .Y(new_new_n569_));
  OA210      g547(.A0(new_new_n569_), .A1(new_new_n223_), .B0(new_new_n81_), .Y(new_new_n570_));
  NA3        g548(.A(new_new_n402_), .B(new_new_n424_), .C(new_new_n46_), .Y(new_new_n571_));
  NO3        g549(.A(new_new_n401_), .B(new_new_n495_), .C(new_new_n81_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n572_), .B(new_new_n25_), .Y(new_new_n573_));
  NA2        g551(.A(new_new_n573_), .B(new_new_n571_), .Y(new_new_n574_));
  OAI210     g552(.A0(new_new_n574_), .A1(new_new_n570_), .B0(i_1_), .Y(new_new_n575_));
  AOI210     g553(.A0(new_new_n242_), .A1(new_new_n93_), .B0(i_1_), .Y(new_new_n576_));
  NO2        g554(.A(new_new_n318_), .B(i_2_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n577_), .B(new_new_n576_), .Y(new_new_n578_));
  AOI210     g556(.A0(new_new_n578_), .A1(new_new_n575_), .B0(i_13_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n54_), .B(i_12_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n401_), .B(new_new_n24_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n873_), .B(new_new_n88_), .Y(new_new_n582_));
  INV        g560(.A(new_new_n582_), .Y(new_new_n583_));
  INV        g561(.A(new_new_n111_), .Y(new_new_n584_));
  AOI220     g562(.A0(new_new_n584_), .A1(new_new_n68_), .B0(new_new_n335_), .B1(new_new_n535_), .Y(new_new_n585_));
  NO2        g563(.A(new_new_n585_), .B(new_new_n221_), .Y(new_new_n586_));
  AOI210     g564(.A0(new_new_n376_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n587_));
  NOi31      g565(.An(new_new_n587_), .B(new_new_n486_), .C(new_new_n44_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n124_), .B(i_13_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n589_), .B(new_new_n576_), .Y(new_new_n590_));
  NO3        g568(.A(new_new_n67_), .B(new_new_n32_), .C(new_new_n97_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n26_), .B(new_new_n181_), .Y(new_new_n592_));
  NA2        g570(.A(new_new_n592_), .B(i_7_), .Y(new_new_n593_));
  NO3        g571(.A(new_new_n401_), .B(new_new_n216_), .C(new_new_n81_), .Y(new_new_n594_));
  AOI210     g572(.A0(new_new_n594_), .A1(new_new_n593_), .B0(new_new_n591_), .Y(new_new_n595_));
  AOI220     g573(.A0(new_new_n335_), .A1(new_new_n535_), .B0(new_new_n87_), .B1(new_new_n98_), .Y(new_new_n596_));
  OAI220     g574(.A0(new_new_n596_), .A1(new_new_n491_), .B0(new_new_n595_), .B1(new_new_n503_), .Y(new_new_n597_));
  NO4        g575(.A(new_new_n597_), .B(new_new_n590_), .C(new_new_n588_), .D(new_new_n586_), .Y(new_new_n598_));
  OR2        g576(.A(i_11_), .B(i_6_), .Y(new_new_n599_));
  NA3        g577(.A(new_new_n490_), .B(new_new_n592_), .C(i_7_), .Y(new_new_n600_));
  NO2        g578(.A(new_new_n600_), .B(new_new_n599_), .Y(new_new_n601_));
  NA3        g579(.A(new_new_n360_), .B(new_new_n494_), .C(new_new_n93_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n527_), .B(i_13_), .Y(new_new_n603_));
  NAi21      g581(.An(i_11_), .B(i_12_), .Y(new_new_n604_));
  NO3        g582(.A(new_new_n401_), .B(new_new_n471_), .C(new_new_n495_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n605_), .B(new_new_n274_), .Y(new_new_n606_));
  NA3        g584(.A(new_new_n606_), .B(new_new_n603_), .C(new_new_n602_), .Y(new_new_n607_));
  OAI210     g585(.A0(new_new_n607_), .A1(new_new_n601_), .B0(new_new_n59_), .Y(new_new_n608_));
  NO2        g586(.A(i_2_), .B(i_12_), .Y(new_new_n609_));
  NA2        g587(.A(new_new_n317_), .B(new_new_n609_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n125_), .B(i_2_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n611_), .B(new_new_n522_), .Y(new_new_n612_));
  NA2        g590(.A(new_new_n612_), .B(new_new_n610_), .Y(new_new_n613_));
  NA3        g591(.A(new_new_n613_), .B(new_new_n45_), .C(new_new_n209_), .Y(new_new_n614_));
  NA4        g592(.A(new_new_n614_), .B(new_new_n608_), .C(new_new_n598_), .D(new_new_n583_), .Y(new_new_n615_));
  OR4        g593(.A(new_new_n615_), .B(new_new_n579_), .C(new_new_n567_), .D(new_new_n505_), .Y(ori5));
  NA2        g594(.A(new_new_n547_), .B(new_new_n245_), .Y(new_new_n617_));
  AN2        g595(.A(new_new_n24_), .B(i_10_), .Y(new_new_n618_));
  NA3        g596(.A(new_new_n618_), .B(new_new_n609_), .C(new_new_n104_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n491_), .B(i_11_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n84_), .B(new_new_n620_), .Y(new_new_n621_));
  NA3        g599(.A(new_new_n621_), .B(new_new_n619_), .C(new_new_n617_), .Y(new_new_n622_));
  NO3        g600(.A(i_11_), .B(new_new_n216_), .C(i_13_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n121_), .B(new_new_n23_), .Y(new_new_n624_));
  NA2        g602(.A(i_12_), .B(i_8_), .Y(new_new_n625_));
  OAI210     g603(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n625_), .Y(new_new_n626_));
  INV        g604(.A(new_new_n375_), .Y(new_new_n627_));
  AOI220     g605(.A0(new_new_n279_), .A1(new_new_n463_), .B0(new_new_n626_), .B1(new_new_n624_), .Y(new_new_n628_));
  INV        g606(.A(new_new_n628_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n629_), .B(new_new_n622_), .Y(new_new_n630_));
  INV        g608(.A(new_new_n163_), .Y(new_new_n631_));
  INV        g609(.A(new_new_n223_), .Y(new_new_n632_));
  OAI210     g610(.A0(new_new_n577_), .A1(new_new_n377_), .B0(new_new_n107_), .Y(new_new_n633_));
  AOI210     g611(.A0(new_new_n633_), .A1(new_new_n632_), .B0(new_new_n631_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n385_), .B(new_new_n26_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n635_), .B(new_new_n365_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n636_), .B(i_2_), .Y(new_new_n637_));
  INV        g615(.A(new_new_n637_), .Y(new_new_n638_));
  AOI210     g616(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n363_), .Y(new_new_n639_));
  AOI210     g617(.A0(new_new_n639_), .A1(new_new_n638_), .B0(new_new_n634_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n179_), .B(new_new_n122_), .Y(new_new_n641_));
  OAI210     g619(.A0(new_new_n641_), .A1(new_new_n624_), .B0(i_2_), .Y(new_new_n642_));
  INV        g620(.A(new_new_n164_), .Y(new_new_n643_));
  NA2        g621(.A(new_new_n643_), .B(new_new_n84_), .Y(new_new_n644_));
  AOI210     g622(.A0(new_new_n644_), .A1(new_new_n642_), .B0(new_new_n181_), .Y(new_new_n645_));
  OA210      g623(.A0(new_new_n508_), .A1(new_new_n123_), .B0(i_13_), .Y(new_new_n646_));
  NA2        g624(.A(new_new_n187_), .B(new_new_n189_), .Y(new_new_n647_));
  NA2        g625(.A(new_new_n148_), .B(new_new_n487_), .Y(new_new_n648_));
  AOI210     g626(.A0(new_new_n648_), .A1(new_new_n647_), .B0(new_new_n322_), .Y(new_new_n649_));
  AOI210     g627(.A0(new_new_n195_), .A1(new_new_n145_), .B0(new_new_n424_), .Y(new_new_n650_));
  NA2        g628(.A(new_new_n650_), .B(new_new_n365_), .Y(new_new_n651_));
  NO2        g629(.A(new_new_n98_), .B(new_new_n44_), .Y(new_new_n652_));
  INV        g630(.A(new_new_n268_), .Y(new_new_n653_));
  NA4        g631(.A(new_new_n653_), .B(new_new_n269_), .C(new_new_n121_), .D(new_new_n42_), .Y(new_new_n654_));
  OAI210     g632(.A0(new_new_n654_), .A1(new_new_n652_), .B0(new_new_n651_), .Y(new_new_n655_));
  NO4        g633(.A(new_new_n655_), .B(new_new_n649_), .C(new_new_n646_), .D(new_new_n645_), .Y(new_new_n656_));
  NA2        g634(.A(new_new_n463_), .B(new_new_n28_), .Y(new_new_n657_));
  NA2        g635(.A(new_new_n623_), .B(new_new_n251_), .Y(new_new_n658_));
  NA2        g636(.A(new_new_n658_), .B(new_new_n657_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n58_), .B(i_12_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n660_), .B(new_new_n123_), .Y(new_new_n661_));
  NO2        g639(.A(new_new_n661_), .B(new_new_n487_), .Y(new_new_n662_));
  AOI220     g640(.A0(new_new_n662_), .A1(new_new_n36_), .B0(new_new_n659_), .B1(new_new_n46_), .Y(new_new_n663_));
  NA4        g641(.A(new_new_n663_), .B(new_new_n656_), .C(new_new_n640_), .D(new_new_n630_), .Y(ori6));
  NO3        g642(.A(i_9_), .B(new_new_n270_), .C(i_1_), .Y(new_new_n665_));
  NO2        g643(.A(new_new_n174_), .B(new_new_n136_), .Y(new_new_n666_));
  OAI210     g644(.A0(new_new_n666_), .A1(new_new_n665_), .B0(new_new_n611_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n205_), .B(new_new_n404_), .Y(new_new_n668_));
  INV        g646(.A(new_new_n286_), .Y(new_new_n669_));
  AO210      g647(.A0(new_new_n669_), .A1(new_new_n667_), .B0(i_12_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n471_), .B(new_new_n59_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n569_), .B(new_new_n67_), .Y(new_new_n672_));
  BUFFER     g650(.A(new_new_n513_), .Y(new_new_n673_));
  NA3        g651(.A(new_new_n673_), .B(new_new_n672_), .C(new_new_n671_), .Y(new_new_n674_));
  NA2        g652(.A(new_new_n674_), .B(new_new_n69_), .Y(new_new_n675_));
  INV        g653(.A(new_new_n285_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n71_), .B(new_new_n128_), .Y(new_new_n677_));
  NO2        g655(.A(new_new_n677_), .B(new_new_n676_), .Y(new_new_n678_));
  NO2        g656(.A(new_new_n226_), .B(i_9_), .Y(new_new_n679_));
  NA2        g657(.A(new_new_n679_), .B(new_new_n660_), .Y(new_new_n680_));
  AOI210     g658(.A0(new_new_n680_), .A1(new_new_n423_), .B0(new_new_n174_), .Y(new_new_n681_));
  NO2        g659(.A(new_new_n32_), .B(i_11_), .Y(new_new_n682_));
  NA3        g660(.A(new_new_n682_), .B(new_new_n398_), .C(new_new_n339_), .Y(new_new_n683_));
  NAi32      g661(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n684_));
  NO2        g662(.A(new_new_n599_), .B(new_new_n684_), .Y(new_new_n685_));
  OAI210     g663(.A0(new_new_n568_), .A1(new_new_n454_), .B0(new_new_n453_), .Y(new_new_n686_));
  NAi31      g664(.An(new_new_n685_), .B(new_new_n686_), .C(new_new_n683_), .Y(new_new_n687_));
  OR3        g665(.A(new_new_n687_), .B(new_new_n681_), .C(new_new_n678_), .Y(new_new_n688_));
  AO220      g666(.A0(new_new_n308_), .A1(new_new_n298_), .B0(new_new_n347_), .B1(new_new_n487_), .Y(new_new_n689_));
  NA3        g667(.A(new_new_n689_), .B(new_new_n230_), .C(i_7_), .Y(new_new_n690_));
  NA3        g668(.A(new_new_n377_), .B(new_new_n144_), .C(new_new_n65_), .Y(new_new_n691_));
  AO210      g669(.A0(new_new_n409_), .A1(new_new_n627_), .B0(new_new_n36_), .Y(new_new_n692_));
  NA3        g670(.A(new_new_n692_), .B(new_new_n691_), .C(new_new_n690_), .Y(new_new_n693_));
  OAI210     g671(.A0(i_6_), .A1(i_11_), .B0(new_new_n82_), .Y(new_new_n694_));
  AOI220     g672(.A0(new_new_n694_), .A1(new_new_n453_), .B0(new_new_n668_), .B1(new_new_n593_), .Y(new_new_n695_));
  NA3        g673(.A(new_new_n322_), .B(new_new_n218_), .C(new_new_n144_), .Y(new_new_n696_));
  NA2        g674(.A(new_new_n347_), .B(new_new_n66_), .Y(new_new_n697_));
  NA4        g675(.A(new_new_n697_), .B(new_new_n696_), .C(new_new_n695_), .D(new_new_n493_), .Y(new_new_n698_));
  AO210      g676(.A0(new_new_n424_), .A1(new_new_n46_), .B0(new_new_n83_), .Y(new_new_n699_));
  NA3        g677(.A(new_new_n699_), .B(new_new_n402_), .C(new_new_n203_), .Y(new_new_n700_));
  AOI210     g678(.A0(new_new_n377_), .A1(new_new_n375_), .B0(new_new_n452_), .Y(new_new_n701_));
  NO2        g679(.A(new_new_n501_), .B(new_new_n98_), .Y(new_new_n702_));
  OAI210     g680(.A0(new_new_n702_), .A1(new_new_n108_), .B0(new_new_n358_), .Y(new_new_n703_));
  NA2        g681(.A(new_new_n222_), .B(new_new_n46_), .Y(new_new_n704_));
  INV        g682(.A(new_new_n476_), .Y(new_new_n705_));
  NA3        g683(.A(new_new_n705_), .B(new_new_n285_), .C(i_7_), .Y(new_new_n706_));
  NA4        g684(.A(new_new_n706_), .B(new_new_n703_), .C(new_new_n701_), .D(new_new_n700_), .Y(new_new_n707_));
  NO4        g685(.A(new_new_n707_), .B(new_new_n698_), .C(new_new_n693_), .D(new_new_n688_), .Y(new_new_n708_));
  NA4        g686(.A(new_new_n708_), .B(new_new_n675_), .C(new_new_n670_), .D(new_new_n329_), .Y(ori3));
  NA2        g687(.A(i_12_), .B(i_10_), .Y(new_new_n710_));
  NO2        g688(.A(i_11_), .B(new_new_n216_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n696_), .B(new_new_n493_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n712_), .B(new_new_n40_), .Y(new_new_n713_));
  NO3        g691(.A(new_new_n518_), .B(new_new_n385_), .C(new_new_n128_), .Y(new_new_n714_));
  NA2        g692(.A(new_new_n360_), .B(new_new_n45_), .Y(new_new_n715_));
  INV        g693(.A(new_new_n714_), .Y(new_new_n716_));
  AOI210     g694(.A0(new_new_n716_), .A1(new_new_n713_), .B0(new_new_n48_), .Y(new_new_n717_));
  NO4        g695(.A(new_new_n326_), .B(new_new_n332_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n718_));
  NA2        g696(.A(new_new_n587_), .B(new_new_n558_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n292_), .B(i_5_), .Y(new_new_n720_));
  OAI220     g698(.A0(new_new_n720_), .A1(new_new_n719_), .B0(new_new_n875_), .B1(new_new_n59_), .Y(new_new_n721_));
  NOi21      g699(.An(i_5_), .B(i_9_), .Y(new_new_n722_));
  NA2        g700(.A(new_new_n722_), .B(new_new_n374_), .Y(new_new_n723_));
  BUFFER     g701(.A(new_new_n242_), .Y(new_new_n724_));
  AOI210     g702(.A0(new_new_n724_), .A1(new_new_n399_), .B0(new_new_n572_), .Y(new_new_n725_));
  NO3        g703(.A(new_new_n361_), .B(new_new_n242_), .C(new_new_n69_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n166_), .B(new_new_n145_), .Y(new_new_n727_));
  AOI210     g705(.A0(new_new_n727_), .A1(new_new_n222_), .B0(new_new_n726_), .Y(new_new_n728_));
  OAI220     g706(.A0(new_new_n728_), .A1(new_new_n169_), .B0(new_new_n725_), .B1(new_new_n723_), .Y(new_new_n729_));
  NO3        g707(.A(new_new_n729_), .B(new_new_n721_), .C(new_new_n717_), .Y(new_new_n730_));
  NA2        g708(.A(new_new_n174_), .B(new_new_n24_), .Y(new_new_n731_));
  NO2        g709(.A(new_new_n556_), .B(new_new_n484_), .Y(new_new_n732_));
  NO2        g710(.A(new_new_n732_), .B(new_new_n731_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n274_), .B(new_new_n126_), .Y(new_new_n734_));
  NAi21      g712(.An(new_new_n155_), .B(i_5_), .Y(new_new_n735_));
  OAI220     g713(.A0(new_new_n735_), .A1(new_new_n704_), .B0(new_new_n734_), .B1(new_new_n352_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n736_), .B(new_new_n733_), .Y(new_new_n737_));
  NA2        g715(.A(new_new_n460_), .B(i_0_), .Y(new_new_n738_));
  NO3        g716(.A(new_new_n738_), .B(new_new_n334_), .C(new_new_n84_), .Y(new_new_n739_));
  NO4        g717(.A(new_new_n475_), .B(new_new_n200_), .C(new_new_n363_), .D(new_new_n359_), .Y(new_new_n740_));
  AOI210     g718(.A0(new_new_n740_), .A1(i_11_), .B0(new_new_n739_), .Y(new_new_n741_));
  INV        g719(.A(new_new_n398_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n623_), .B(new_new_n286_), .Y(new_new_n743_));
  AOI210     g721(.A0(new_new_n402_), .A1(new_new_n84_), .B0(new_new_n56_), .Y(new_new_n744_));
  OAI220     g722(.A0(new_new_n744_), .A1(new_new_n743_), .B0(new_new_n542_), .B1(new_new_n432_), .Y(new_new_n745_));
  NO2        g723(.A(new_new_n228_), .B(new_new_n149_), .Y(new_new_n746_));
  NA2        g724(.A(i_0_), .B(i_10_), .Y(new_new_n747_));
  INV        g725(.A(new_new_n434_), .Y(new_new_n748_));
  NO4        g726(.A(new_new_n111_), .B(new_new_n56_), .C(new_new_n551_), .D(i_5_), .Y(new_new_n749_));
  AO220      g727(.A0(new_new_n749_), .A1(new_new_n748_), .B0(new_new_n746_), .B1(i_6_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n177_), .B(new_new_n189_), .Y(new_new_n751_));
  NO2        g729(.A(new_new_n751_), .B(new_new_n743_), .Y(new_new_n752_));
  NO3        g730(.A(new_new_n752_), .B(new_new_n750_), .C(new_new_n745_), .Y(new_new_n753_));
  NA3        g731(.A(new_new_n753_), .B(new_new_n741_), .C(new_new_n737_), .Y(new_new_n754_));
  NA2        g732(.A(i_11_), .B(i_9_), .Y(new_new_n755_));
  NA2        g733(.A(new_new_n344_), .B(new_new_n167_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n756_), .B(new_new_n153_), .Y(new_new_n757_));
  NO2        g735(.A(new_new_n755_), .B(new_new_n69_), .Y(new_new_n758_));
  NO2        g736(.A(new_new_n166_), .B(i_0_), .Y(new_new_n759_));
  INV        g737(.A(new_new_n757_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n541_), .B(new_new_n118_), .Y(new_new_n761_));
  NO2        g739(.A(i_6_), .B(new_new_n761_), .Y(new_new_n762_));
  AOI210     g740(.A0(new_new_n376_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n763_));
  NA2        g741(.A(new_new_n163_), .B(new_new_n99_), .Y(new_new_n764_));
  NOi32      g742(.An(new_new_n763_), .Bn(new_new_n177_), .C(new_new_n764_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n494_), .B(new_new_n286_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n766_), .B(new_new_n715_), .Y(new_new_n767_));
  NO3        g745(.A(new_new_n767_), .B(new_new_n765_), .C(new_new_n762_), .Y(new_new_n768_));
  NOi21      g746(.An(i_7_), .B(i_5_), .Y(new_new_n769_));
  NOi31      g747(.An(new_new_n769_), .B(i_0_), .C(new_new_n604_), .Y(new_new_n770_));
  NA3        g748(.A(new_new_n770_), .B(new_new_n333_), .C(i_6_), .Y(new_new_n771_));
  OA210      g749(.A0(new_new_n764_), .A1(new_new_n423_), .B0(new_new_n771_), .Y(new_new_n772_));
  INV        g750(.A(new_new_n280_), .Y(new_new_n773_));
  NA3        g751(.A(new_new_n772_), .B(new_new_n768_), .C(new_new_n760_), .Y(new_new_n774_));
  NO2        g752(.A(new_new_n710_), .B(new_new_n279_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n775_), .B(new_new_n758_), .Y(new_new_n776_));
  NA3        g754(.A(new_new_n397_), .B(new_new_n360_), .C(new_new_n45_), .Y(new_new_n777_));
  OAI210     g755(.A0(new_new_n735_), .A1(new_new_n742_), .B0(new_new_n777_), .Y(new_new_n778_));
  NO2        g756(.A(new_new_n230_), .B(new_new_n46_), .Y(new_new_n779_));
  NA2        g757(.A(new_new_n758_), .B(new_new_n269_), .Y(new_new_n780_));
  OAI210     g758(.A0(new_new_n779_), .A1(new_new_n176_), .B0(new_new_n780_), .Y(new_new_n781_));
  AOI220     g759(.A0(new_new_n781_), .A1(new_new_n398_), .B0(new_new_n778_), .B1(new_new_n69_), .Y(new_new_n782_));
  NO2        g760(.A(new_new_n71_), .B(new_new_n625_), .Y(new_new_n783_));
  AOI210     g761(.A0(new_new_n165_), .A1(new_new_n484_), .B0(new_new_n783_), .Y(new_new_n784_));
  NO2        g762(.A(new_new_n784_), .B(new_new_n47_), .Y(new_new_n785_));
  NO3        g763(.A(new_new_n475_), .B(new_new_n306_), .C(new_new_n24_), .Y(new_new_n786_));
  AOI210     g764(.A0(new_new_n581_), .A1(new_new_n442_), .B0(new_new_n786_), .Y(new_new_n787_));
  NAi21      g765(.An(i_9_), .B(i_5_), .Y(new_new_n788_));
  NO2        g766(.A(new_new_n787_), .B(new_new_n164_), .Y(new_new_n789_));
  NO2        g767(.A(new_new_n789_), .B(new_new_n785_), .Y(new_new_n790_));
  NA3        g768(.A(new_new_n790_), .B(new_new_n782_), .C(new_new_n776_), .Y(new_new_n791_));
  NO3        g769(.A(new_new_n791_), .B(new_new_n774_), .C(new_new_n754_), .Y(new_new_n792_));
  NO2        g770(.A(i_0_), .B(new_new_n604_), .Y(new_new_n793_));
  NA2        g771(.A(new_new_n69_), .B(new_new_n44_), .Y(new_new_n794_));
  AN2        g772(.A(new_new_n793_), .B(new_new_n165_), .Y(new_new_n795_));
  NO2        g773(.A(new_new_n671_), .B(new_new_n764_), .Y(new_new_n796_));
  AOI210     g774(.A0(new_new_n795_), .A1(new_new_n297_), .B0(new_new_n796_), .Y(new_new_n797_));
  NO2        g775(.A(new_new_n686_), .B(new_new_n353_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n222_), .B(new_new_n213_), .Y(new_new_n799_));
  AOI210     g777(.A0(new_new_n799_), .A1(new_new_n738_), .B0(new_new_n149_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n800_), .B(new_new_n798_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n801_), .B(new_new_n797_), .Y(new_new_n802_));
  NO3        g780(.A(new_new_n747_), .B(new_new_n722_), .C(new_new_n179_), .Y(new_new_n803_));
  AOI220     g781(.A0(new_new_n803_), .A1(i_11_), .B0(new_new_n456_), .B1(new_new_n71_), .Y(new_new_n804_));
  NO3        g782(.A(new_new_n196_), .B(new_new_n332_), .C(i_0_), .Y(new_new_n805_));
  OAI210     g783(.A0(new_new_n805_), .A1(new_new_n72_), .B0(i_13_), .Y(new_new_n806_));
  NA2        g784(.A(new_new_n806_), .B(new_new_n804_), .Y(new_new_n807_));
  INV        g785(.A(new_new_n105_), .Y(new_new_n808_));
  OR2        g786(.A(new_new_n808_), .B(i_5_), .Y(new_new_n809_));
  NO3        g787(.A(new_new_n715_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n408_), .B(new_new_n403_), .Y(new_new_n811_));
  NO2        g789(.A(new_new_n811_), .B(new_new_n810_), .Y(new_new_n812_));
  NA3        g790(.A(new_new_n339_), .B(new_new_n163_), .C(new_new_n162_), .Y(new_new_n813_));
  INV        g791(.A(new_new_n813_), .Y(new_new_n814_));
  NA3        g792(.A(new_new_n339_), .B(new_new_n293_), .C(new_new_n206_), .Y(new_new_n815_));
  INV        g793(.A(new_new_n815_), .Y(new_new_n816_));
  NOi31      g794(.An(new_new_n338_), .B(new_new_n794_), .C(new_new_n219_), .Y(new_new_n817_));
  NO3        g795(.A(new_new_n755_), .B(new_new_n203_), .C(new_new_n179_), .Y(new_new_n818_));
  NO4        g796(.A(new_new_n818_), .B(new_new_n817_), .C(new_new_n816_), .D(new_new_n814_), .Y(new_new_n819_));
  NA3        g797(.A(new_new_n819_), .B(new_new_n812_), .C(new_new_n809_), .Y(new_new_n820_));
  NO2        g798(.A(new_new_n81_), .B(i_5_), .Y(new_new_n821_));
  NA3        g799(.A(new_new_n711_), .B(new_new_n106_), .C(new_new_n121_), .Y(new_new_n822_));
  INV        g800(.A(new_new_n822_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n823_), .B(new_new_n821_), .Y(new_new_n824_));
  NA3        g802(.A(new_new_n269_), .B(i_5_), .C(new_new_n181_), .Y(new_new_n825_));
  NAi31      g803(.An(new_new_n220_), .B(new_new_n825_), .C(new_new_n221_), .Y(new_new_n826_));
  NO4        g804(.A(new_new_n219_), .B(new_new_n196_), .C(i_0_), .D(i_12_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n827_), .B(new_new_n826_), .Y(new_new_n828_));
  AN2        g806(.A(new_new_n747_), .B(new_new_n149_), .Y(new_new_n829_));
  NO4        g807(.A(new_new_n829_), .B(i_12_), .C(new_new_n532_), .D(new_new_n128_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n830_), .B(new_new_n203_), .Y(new_new_n831_));
  NA3        g809(.A(new_new_n94_), .B(new_new_n459_), .C(i_11_), .Y(new_new_n832_));
  NO2        g810(.A(new_new_n832_), .B(new_new_n69_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n60_), .B(new_new_n97_), .Y(new_new_n834_));
  NO2        g812(.A(new_new_n834_), .B(new_new_n825_), .Y(new_new_n835_));
  AOI210     g813(.A0(new_new_n835_), .A1(new_new_n759_), .B0(new_new_n833_), .Y(new_new_n836_));
  NA4        g814(.A(new_new_n836_), .B(new_new_n831_), .C(new_new_n828_), .D(new_new_n824_), .Y(new_new_n837_));
  NO4        g815(.A(new_new_n837_), .B(new_new_n820_), .C(new_new_n807_), .D(new_new_n802_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n682_), .B(new_new_n37_), .Y(new_new_n839_));
  NA3        g817(.A(new_new_n763_), .B(new_new_n317_), .C(i_5_), .Y(new_new_n840_));
  NA3        g818(.A(new_new_n840_), .B(new_new_n839_), .C(new_new_n500_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n841_), .B(new_new_n194_), .Y(new_new_n842_));
  BUFFER     g820(.A(new_new_n318_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n175_), .B(new_new_n177_), .Y(new_new_n844_));
  AO210      g822(.A0(new_new_n843_), .A1(new_new_n33_), .B0(new_new_n844_), .Y(new_new_n845_));
  INV        g823(.A(new_new_n529_), .Y(new_new_n846_));
  NA2        g824(.A(new_new_n846_), .B(new_new_n845_), .Y(new_new_n847_));
  AOI210     g825(.A0(new_new_n847_), .A1(new_new_n48_), .B0(new_new_n740_), .Y(new_new_n848_));
  AOI210     g826(.A0(new_new_n848_), .A1(new_new_n842_), .B0(new_new_n69_), .Y(new_new_n849_));
  INV        g827(.A(new_new_n72_), .Y(new_new_n850_));
  INV        g828(.A(new_new_n770_), .Y(new_new_n851_));
  AOI210     g829(.A0(new_new_n851_), .A1(new_new_n850_), .B0(new_new_n562_), .Y(new_new_n852_));
  INV        g830(.A(new_new_n852_), .Y(new_new_n853_));
  OAI210     g831(.A0(new_new_n244_), .A1(new_new_n151_), .B0(new_new_n84_), .Y(new_new_n854_));
  NA3        g832(.A(new_new_n635_), .B(new_new_n260_), .C(new_new_n76_), .Y(new_new_n855_));
  AOI210     g833(.A0(new_new_n855_), .A1(new_new_n854_), .B0(i_11_), .Y(new_new_n856_));
  NA2        g834(.A(new_new_n495_), .B(new_new_n200_), .Y(new_new_n857_));
  OAI210     g835(.A0(new_new_n857_), .A1(new_new_n763_), .B0(new_new_n194_), .Y(new_new_n858_));
  NA2        g836(.A(new_new_n157_), .B(i_5_), .Y(new_new_n859_));
  NO2        g837(.A(new_new_n858_), .B(new_new_n859_), .Y(new_new_n860_));
  NO3        g838(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n861_));
  OAI210     g839(.A0(new_new_n773_), .A1(new_new_n270_), .B0(new_new_n861_), .Y(new_new_n862_));
  NO2        g840(.A(new_new_n862_), .B(new_new_n604_), .Y(new_new_n863_));
  NO4        g841(.A(new_new_n788_), .B(new_new_n400_), .C(new_new_n227_), .D(new_new_n226_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n864_), .B(new_new_n452_), .Y(new_new_n865_));
  NO2        g843(.A(new_new_n865_), .B(new_new_n41_), .Y(new_new_n866_));
  NO4        g844(.A(new_new_n866_), .B(new_new_n863_), .C(new_new_n860_), .D(new_new_n856_), .Y(new_new_n867_));
  OAI210     g845(.A0(new_new_n853_), .A1(i_4_), .B0(new_new_n867_), .Y(new_new_n868_));
  NO2        g846(.A(new_new_n868_), .B(new_new_n849_), .Y(new_new_n869_));
  NA4        g847(.A(new_new_n869_), .B(new_new_n838_), .C(new_new_n792_), .D(new_new_n730_), .Y(ori4));
  INV        g848(.A(new_new_n580_), .Y(new_new_n873_));
  INV        g849(.A(new_new_n78_), .Y(new_new_n874_));
  INV        g850(.A(new_new_n718_), .Y(new_new_n875_));
endmodule


