//Benchmark atmr_alu4_1266_0.0625

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n137_, ori_ori_n138_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n56_));
  NO2        o034(.A(i_1_), .B(i_6_), .Y(ori_ori_n57_));
  NA2        o035(.A(i_8_), .B(i_7_), .Y(ori_ori_n58_));
  NAi21      o036(.An(i_2_), .B(i_7_), .Y(ori_ori_n59_));
  INV        o037(.A(i_1_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(i_6_), .Y(ori_ori_n61_));
  NA3        o039(.A(ori_ori_n61_), .B(ori_ori_n59_), .C(ori_ori_n31_), .Y(ori_ori_n62_));
  NA2        o040(.A(i_1_), .B(i_10_), .Y(ori_ori_n63_));
  NO2        o041(.A(ori_ori_n63_), .B(i_6_), .Y(ori_ori_n64_));
  NAi21      o042(.An(ori_ori_n64_), .B(ori_ori_n62_), .Y(ori_ori_n65_));
  NA2        o043(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n66_));
  AOI210     o044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n67_));
  NA2        o045(.A(i_1_), .B(i_6_), .Y(ori_ori_n68_));
  NO2        o046(.A(ori_ori_n68_), .B(ori_ori_n25_), .Y(ori_ori_n69_));
  INV        o047(.A(i_0_), .Y(ori_ori_n70_));
  NAi21      o048(.An(i_5_), .B(i_10_), .Y(ori_ori_n71_));
  NA2        o049(.A(i_5_), .B(i_9_), .Y(ori_ori_n72_));
  AOI210     o050(.A0(ori_ori_n72_), .A1(ori_ori_n71_), .B0(ori_ori_n70_), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n73_), .B(ori_ori_n69_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n67_), .A1(ori_ori_n66_), .B0(ori_ori_n74_), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n65_), .B0(i_0_), .Y(ori_ori_n76_));
  NA2        o054(.A(i_12_), .B(i_5_), .Y(ori_ori_n77_));
  NA2        o055(.A(i_2_), .B(i_8_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n78_), .B(ori_ori_n57_), .Y(ori_ori_n79_));
  NO2        o057(.A(i_3_), .B(i_9_), .Y(ori_ori_n80_));
  NO2        o058(.A(i_3_), .B(i_7_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n80_), .B(ori_ori_n60_), .Y(ori_ori_n82_));
  INV        o060(.A(i_6_), .Y(ori_ori_n83_));
  OR4        o061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n84_), .Y(ori_ori_n85_));
  NO2        o063(.A(i_2_), .B(i_7_), .Y(ori_ori_n86_));
  NO2        o064(.A(ori_ori_n85_), .B(ori_ori_n86_), .Y(ori_ori_n87_));
  OAI210     o065(.A0(ori_ori_n82_), .A1(ori_ori_n79_), .B0(ori_ori_n87_), .Y(ori_ori_n88_));
  NAi21      o066(.An(i_6_), .B(i_10_), .Y(ori_ori_n89_));
  NA2        o067(.A(i_6_), .B(i_9_), .Y(ori_ori_n90_));
  AOI210     o068(.A0(ori_ori_n90_), .A1(ori_ori_n89_), .B0(ori_ori_n60_), .Y(ori_ori_n91_));
  NA2        o069(.A(i_2_), .B(i_6_), .Y(ori_ori_n92_));
  NO3        o070(.A(ori_ori_n92_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n93_), .B(ori_ori_n91_), .Y(ori_ori_n94_));
  AOI210     o072(.A0(ori_ori_n94_), .A1(ori_ori_n88_), .B0(ori_ori_n77_), .Y(ori_ori_n95_));
  AN3        o073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n96_));
  NAi21      o074(.An(i_6_), .B(i_11_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n96_), .B(ori_ori_n32_), .Y(ori_ori_n98_));
  INV        o076(.A(i_7_), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n46_), .B(ori_ori_n99_), .Y(ori_ori_n100_));
  NO2        o078(.A(i_0_), .B(i_5_), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n101_), .B(ori_ori_n83_), .Y(ori_ori_n102_));
  NA2        o080(.A(i_12_), .B(i_3_), .Y(ori_ori_n103_));
  INV        o081(.A(ori_ori_n103_), .Y(ori_ori_n104_));
  NA3        o082(.A(ori_ori_n104_), .B(ori_ori_n102_), .C(ori_ori_n100_), .Y(ori_ori_n105_));
  NAi21      o083(.An(i_7_), .B(i_11_), .Y(ori_ori_n106_));
  NO3        o084(.A(ori_ori_n106_), .B(ori_ori_n89_), .C(ori_ori_n53_), .Y(ori_ori_n107_));
  AN2        o085(.A(i_2_), .B(i_10_), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n108_), .B(i_7_), .Y(ori_ori_n109_));
  OR2        o087(.A(ori_ori_n77_), .B(ori_ori_n57_), .Y(ori_ori_n110_));
  NO2        o088(.A(i_8_), .B(ori_ori_n99_), .Y(ori_ori_n111_));
  NO3        o089(.A(ori_ori_n111_), .B(ori_ori_n110_), .C(ori_ori_n109_), .Y(ori_ori_n112_));
  NA2        o090(.A(i_12_), .B(i_7_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n60_), .B(ori_ori_n26_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n114_), .B(i_0_), .Y(ori_ori_n115_));
  NA2        o093(.A(i_11_), .B(i_12_), .Y(ori_ori_n116_));
  OAI210     o094(.A0(ori_ori_n115_), .A1(ori_ori_n113_), .B0(ori_ori_n116_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n117_), .B(ori_ori_n112_), .Y(ori_ori_n118_));
  NAi41      o096(.An(ori_ori_n107_), .B(ori_ori_n118_), .C(ori_ori_n105_), .D(ori_ori_n98_), .Y(ori_ori_n119_));
  NOi21      o097(.An(i_1_), .B(i_5_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(i_11_), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n99_), .B(ori_ori_n37_), .Y(ori_ori_n122_));
  NA2        o100(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(ori_ori_n122_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n124_), .B(ori_ori_n46_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n90_), .B(ori_ori_n89_), .Y(ori_ori_n126_));
  NAi21      o104(.An(i_3_), .B(i_8_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n127_), .B(ori_ori_n59_), .Y(ori_ori_n128_));
  NOi31      o106(.An(ori_ori_n128_), .B(ori_ori_n126_), .C(ori_ori_n125_), .Y(ori_ori_n129_));
  NO2        o107(.A(i_1_), .B(ori_ori_n83_), .Y(ori_ori_n130_));
  NO2        o108(.A(i_6_), .B(i_5_), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n131_), .B(i_3_), .Y(ori_ori_n132_));
  AO210      o110(.A0(ori_ori_n132_), .A1(ori_ori_n47_), .B0(ori_ori_n130_), .Y(ori_ori_n133_));
  OAI220     o111(.A0(ori_ori_n133_), .A1(ori_ori_n106_), .B0(ori_ori_n129_), .B1(ori_ori_n121_), .Y(ori_ori_n134_));
  NO3        o112(.A(ori_ori_n134_), .B(ori_ori_n119_), .C(ori_ori_n95_), .Y(ori_ori_n135_));
  NA3        o113(.A(ori_ori_n135_), .B(ori_ori_n76_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o114(.A(ori_ori_n60_), .B(ori_ori_n37_), .Y(ori_ori_n137_));
  NA2        o115(.A(ori_ori_n754_), .B(ori_ori_n137_), .Y(ori_ori_n138_));
  NA4        o116(.A(ori_ori_n138_), .B(ori_ori_n74_), .C(ori_ori_n66_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o117(.A(i_12_), .B(i_13_), .Y(ori_ori_n140_));
  NAi21      o118(.An(i_5_), .B(i_11_), .Y(ori_ori_n141_));
  NO2        o119(.A(i_0_), .B(i_1_), .Y(ori_ori_n142_));
  NA2        o120(.A(i_2_), .B(i_3_), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n143_), .B(i_4_), .Y(ori_ori_n144_));
  NA2        o122(.A(i_1_), .B(i_5_), .Y(ori_ori_n145_));
  OR2        o123(.A(i_0_), .B(i_1_), .Y(ori_ori_n146_));
  NAi32      o124(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n147_));
  NOi21      o125(.An(i_4_), .B(i_10_), .Y(ori_ori_n148_));
  NA2        o126(.A(ori_ori_n148_), .B(ori_ori_n40_), .Y(ori_ori_n149_));
  NOi21      o127(.An(i_4_), .B(i_9_), .Y(ori_ori_n150_));
  NOi21      o128(.An(i_11_), .B(i_13_), .Y(ori_ori_n151_));
  NA2        o129(.A(ori_ori_n151_), .B(ori_ori_n150_), .Y(ori_ori_n152_));
  NO2        o130(.A(i_4_), .B(i_5_), .Y(ori_ori_n153_));
  NAi21      o131(.An(i_12_), .B(i_11_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n154_), .B(i_13_), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n70_), .B(ori_ori_n60_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n70_), .B(i_5_), .Y(ori_ori_n157_));
  NO2        o135(.A(i_13_), .B(i_10_), .Y(ori_ori_n158_));
  NO2        o136(.A(i_2_), .B(i_1_), .Y(ori_ori_n159_));
  NAi21      o137(.An(i_4_), .B(i_12_), .Y(ori_ori_n160_));
  INV        o138(.A(i_8_), .Y(ori_ori_n161_));
  NO3        o139(.A(i_3_), .B(ori_ori_n83_), .C(ori_ori_n48_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n162_), .B(ori_ori_n111_), .Y(ori_ori_n163_));
  NO3        o141(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n164_));
  NO2        o142(.A(i_3_), .B(i_8_), .Y(ori_ori_n165_));
  NO3        o143(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n166_));
  NA3        o144(.A(ori_ori_n166_), .B(ori_ori_n165_), .C(ori_ori_n40_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n101_), .B(ori_ori_n57_), .Y(ori_ori_n168_));
  INV        o146(.A(ori_ori_n168_), .Y(ori_ori_n169_));
  NO2        o147(.A(i_13_), .B(i_9_), .Y(ori_ori_n170_));
  NAi21      o148(.An(i_12_), .B(i_3_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n169_), .B(ori_ori_n167_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n173_), .B(i_7_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n174_), .B(i_4_), .Y(ori_ori_n175_));
  NAi21      o153(.An(i_12_), .B(i_7_), .Y(ori_ori_n176_));
  NA3        o154(.A(i_13_), .B(ori_ori_n161_), .C(i_10_), .Y(ori_ori_n177_));
  NA2        o155(.A(i_0_), .B(i_5_), .Y(ori_ori_n178_));
  NAi31      o156(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n70_), .B(ori_ori_n26_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n46_), .B(ori_ori_n60_), .Y(ori_ori_n182_));
  INV        o160(.A(i_13_), .Y(ori_ori_n183_));
  NO2        o161(.A(i_12_), .B(ori_ori_n183_), .Y(ori_ori_n184_));
  NO2        o162(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n185_));
  OR2        o163(.A(i_8_), .B(i_7_), .Y(ori_ori_n186_));
  INV        o164(.A(i_12_), .Y(ori_ori_n187_));
  NO3        o165(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n188_));
  NA2        o166(.A(i_2_), .B(i_1_), .Y(ori_ori_n189_));
  NO3        o167(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n190_));
  NAi21      o168(.An(i_4_), .B(i_3_), .Y(ori_ori_n191_));
  NO2        o169(.A(i_0_), .B(i_6_), .Y(ori_ori_n192_));
  NOi41      o170(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n193_));
  NA2        o171(.A(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n194_));
  NO2        o172(.A(i_11_), .B(ori_ori_n183_), .Y(ori_ori_n195_));
  NOi21      o173(.An(i_1_), .B(i_6_), .Y(ori_ori_n196_));
  NAi21      o174(.An(i_3_), .B(i_7_), .Y(ori_ori_n197_));
  NA2        o175(.A(ori_ori_n187_), .B(i_9_), .Y(ori_ori_n198_));
  OR4        o176(.A(ori_ori_n198_), .B(ori_ori_n197_), .C(ori_ori_n196_), .D(ori_ori_n157_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n70_), .B(i_5_), .Y(ori_ori_n200_));
  NA2        o178(.A(i_3_), .B(i_9_), .Y(ori_ori_n201_));
  NAi21      o179(.An(i_7_), .B(i_10_), .Y(ori_ori_n202_));
  NO2        o180(.A(ori_ori_n202_), .B(ori_ori_n201_), .Y(ori_ori_n203_));
  NA3        o181(.A(ori_ori_n203_), .B(ori_ori_n200_), .C(ori_ori_n61_), .Y(ori_ori_n204_));
  NA2        o182(.A(ori_ori_n204_), .B(ori_ori_n199_), .Y(ori_ori_n205_));
  NA2        o183(.A(ori_ori_n205_), .B(ori_ori_n195_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n186_), .B(ori_ori_n37_), .Y(ori_ori_n207_));
  NA2        o185(.A(i_12_), .B(i_6_), .Y(ori_ori_n208_));
  OR2        o186(.A(i_13_), .B(i_9_), .Y(ori_ori_n209_));
  NO3        o187(.A(ori_ori_n209_), .B(ori_ori_n208_), .C(ori_ori_n48_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n191_), .B(i_2_), .Y(ori_ori_n211_));
  NA3        o189(.A(ori_ori_n211_), .B(ori_ori_n210_), .C(ori_ori_n44_), .Y(ori_ori_n212_));
  NA2        o190(.A(ori_ori_n195_), .B(i_9_), .Y(ori_ori_n213_));
  NA2        o191(.A(ori_ori_n200_), .B(ori_ori_n61_), .Y(ori_ori_n214_));
  OAI210     o192(.A0(ori_ori_n214_), .A1(ori_ori_n213_), .B0(ori_ori_n212_), .Y(ori_ori_n215_));
  NO3        o193(.A(i_11_), .B(ori_ori_n183_), .C(ori_ori_n25_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n197_), .B(i_8_), .Y(ori_ori_n217_));
  NA2        o195(.A(ori_ori_n215_), .B(ori_ori_n207_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n218_), .B(ori_ori_n206_), .Y(ori_ori_n219_));
  NO3        o197(.A(i_12_), .B(ori_ori_n183_), .C(ori_ori_n37_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n189_), .B(i_0_), .Y(ori_ori_n221_));
  NO2        o199(.A(i_3_), .B(i_10_), .Y(ori_ori_n222_));
  NO2        o200(.A(i_2_), .B(ori_ori_n99_), .Y(ori_ori_n223_));
  AN2        o201(.A(i_3_), .B(i_10_), .Y(ori_ori_n224_));
  NO2        o202(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n219_), .B(ori_ori_n175_), .Y(ori_ori_n227_));
  NO3        o205(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n228_));
  NO2        o206(.A(i_2_), .B(i_3_), .Y(ori_ori_n229_));
  OR2        o207(.A(i_0_), .B(i_5_), .Y(ori_ori_n230_));
  NO2        o208(.A(i_12_), .B(i_10_), .Y(ori_ori_n231_));
  NOi21      o209(.An(i_5_), .B(i_0_), .Y(ori_ori_n232_));
  NO2        o210(.A(i_2_), .B(ori_ori_n99_), .Y(ori_ori_n233_));
  NO4        o211(.A(ori_ori_n233_), .B(i_4_), .C(ori_ori_n232_), .D(ori_ori_n127_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n234_), .B(ori_ori_n231_), .Y(ori_ori_n235_));
  NO2        o213(.A(i_6_), .B(i_8_), .Y(ori_ori_n236_));
  NO2        o214(.A(i_1_), .B(i_7_), .Y(ori_ori_n237_));
  INV        o215(.A(ori_ori_n235_), .Y(ori_ori_n238_));
  NOi21      o216(.An(ori_ori_n145_), .B(ori_ori_n102_), .Y(ori_ori_n239_));
  NO2        o217(.A(ori_ori_n239_), .B(ori_ori_n123_), .Y(ori_ori_n240_));
  NA2        o218(.A(ori_ori_n240_), .B(i_3_), .Y(ori_ori_n241_));
  NO2        o219(.A(ori_ori_n161_), .B(i_9_), .Y(ori_ori_n242_));
  NA2        o220(.A(ori_ori_n242_), .B(ori_ori_n168_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n243_), .B(ori_ori_n46_), .Y(ori_ori_n244_));
  INV        o222(.A(ori_ori_n244_), .Y(ori_ori_n245_));
  AOI210     o223(.A0(ori_ori_n245_), .A1(ori_ori_n241_), .B0(ori_ori_n149_), .Y(ori_ori_n246_));
  AOI210     o224(.A0(ori_ori_n238_), .A1(ori_ori_n228_), .B0(ori_ori_n246_), .Y(ori_ori_n247_));
  NOi32      o225(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n248_));
  INV        o226(.A(ori_ori_n248_), .Y(ori_ori_n249_));
  NAi21      o227(.An(i_0_), .B(i_6_), .Y(ori_ori_n250_));
  NAi21      o228(.An(i_1_), .B(i_5_), .Y(ori_ori_n251_));
  NA2        o229(.A(ori_ori_n251_), .B(ori_ori_n250_), .Y(ori_ori_n252_));
  NA2        o230(.A(ori_ori_n252_), .B(ori_ori_n25_), .Y(ori_ori_n253_));
  OAI210     o231(.A0(ori_ori_n253_), .A1(ori_ori_n147_), .B0(ori_ori_n194_), .Y(ori_ori_n254_));
  NAi41      o232(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n255_));
  OAI220     o233(.A0(ori_ori_n255_), .A1(ori_ori_n251_), .B0(ori_ori_n179_), .B1(ori_ori_n147_), .Y(ori_ori_n256_));
  AOI210     o234(.A0(ori_ori_n255_), .A1(ori_ori_n147_), .B0(ori_ori_n146_), .Y(ori_ori_n257_));
  NOi32      o235(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n258_));
  NAi21      o236(.An(i_6_), .B(i_1_), .Y(ori_ori_n259_));
  NA3        o237(.A(ori_ori_n259_), .B(ori_ori_n258_), .C(ori_ori_n46_), .Y(ori_ori_n260_));
  NO2        o238(.A(ori_ori_n260_), .B(i_0_), .Y(ori_ori_n261_));
  OR3        o239(.A(ori_ori_n261_), .B(ori_ori_n257_), .C(ori_ori_n256_), .Y(ori_ori_n262_));
  NO2        o240(.A(i_1_), .B(ori_ori_n99_), .Y(ori_ori_n263_));
  NAi21      o241(.An(i_3_), .B(i_4_), .Y(ori_ori_n264_));
  NO2        o242(.A(ori_ori_n264_), .B(i_9_), .Y(ori_ori_n265_));
  AN2        o243(.A(i_6_), .B(i_7_), .Y(ori_ori_n266_));
  NA2        o244(.A(i_2_), .B(i_7_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n264_), .B(i_10_), .Y(ori_ori_n268_));
  AOI210     o246(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n269_));
  OAI210     o247(.A0(ori_ori_n269_), .A1(ori_ori_n159_), .B0(ori_ori_n268_), .Y(ori_ori_n270_));
  AOI220     o248(.A0(ori_ori_n268_), .A1(ori_ori_n237_), .B0(ori_ori_n188_), .B1(ori_ori_n159_), .Y(ori_ori_n271_));
  AOI210     o249(.A0(ori_ori_n271_), .A1(ori_ori_n270_), .B0(i_5_), .Y(ori_ori_n272_));
  NO3        o250(.A(ori_ori_n272_), .B(ori_ori_n262_), .C(ori_ori_n254_), .Y(ori_ori_n273_));
  NO2        o251(.A(ori_ori_n273_), .B(ori_ori_n249_), .Y(ori_ori_n274_));
  AN2        o252(.A(i_12_), .B(i_5_), .Y(ori_ori_n275_));
  NA2        o253(.A(i_3_), .B(ori_ori_n275_), .Y(ori_ori_n276_));
  NO2        o254(.A(i_11_), .B(i_6_), .Y(ori_ori_n277_));
  NO2        o255(.A(i_5_), .B(i_10_), .Y(ori_ori_n278_));
  NO2        o256(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n279_));
  NO3        o257(.A(ori_ori_n83_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n280_));
  NA3        o258(.A(ori_ori_n222_), .B(ori_ori_n90_), .C(ori_ori_n72_), .Y(ori_ori_n281_));
  NO2        o259(.A(i_11_), .B(i_12_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n282_), .B(ori_ori_n36_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n281_), .B(ori_ori_n283_), .Y(ori_ori_n284_));
  NAi21      o262(.An(i_13_), .B(i_0_), .Y(ori_ori_n285_));
  NO2        o263(.A(ori_ori_n285_), .B(ori_ori_n189_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n284_), .B(ori_ori_n286_), .Y(ori_ori_n287_));
  INV        o265(.A(ori_ori_n287_), .Y(ori_ori_n288_));
  NO2        o266(.A(i_0_), .B(i_11_), .Y(ori_ori_n289_));
  NOi21      o267(.An(i_2_), .B(i_12_), .Y(ori_ori_n290_));
  NAi21      o268(.An(i_9_), .B(i_4_), .Y(ori_ori_n291_));
  OR2        o269(.A(i_13_), .B(i_10_), .Y(ori_ori_n292_));
  NO3        o270(.A(ori_ori_n292_), .B(ori_ori_n116_), .C(ori_ori_n291_), .Y(ori_ori_n293_));
  NO2        o271(.A(ori_ori_n152_), .B(ori_ori_n122_), .Y(ori_ori_n294_));
  NO2        o272(.A(ori_ori_n99_), .B(ori_ori_n25_), .Y(ori_ori_n295_));
  NA2        o273(.A(ori_ori_n220_), .B(ori_ori_n295_), .Y(ori_ori_n296_));
  NO2        o274(.A(ori_ori_n296_), .B(ori_ori_n239_), .Y(ori_ori_n297_));
  INV        o275(.A(ori_ori_n297_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n298_), .B(ori_ori_n26_), .Y(ori_ori_n299_));
  NA2        o277(.A(ori_ori_n161_), .B(i_10_), .Y(ori_ori_n300_));
  NA3        o278(.A(ori_ori_n200_), .B(ori_ori_n61_), .C(i_2_), .Y(ori_ori_n301_));
  NO2        o279(.A(ori_ori_n301_), .B(ori_ori_n300_), .Y(ori_ori_n302_));
  INV        o280(.A(ori_ori_n302_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n303_), .B(ori_ori_n213_), .Y(ori_ori_n304_));
  NO4        o282(.A(ori_ori_n304_), .B(ori_ori_n299_), .C(ori_ori_n288_), .D(ori_ori_n274_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n70_), .B(i_13_), .Y(ori_ori_n306_));
  NO2        o284(.A(i_10_), .B(i_9_), .Y(ori_ori_n307_));
  NAi21      o285(.An(i_12_), .B(i_8_), .Y(ori_ori_n308_));
  NO2        o286(.A(ori_ori_n308_), .B(i_3_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n310_));
  NA2        o288(.A(ori_ori_n310_), .B(ori_ori_n102_), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n311_), .B(ori_ori_n167_), .Y(ori_ori_n312_));
  NA2        o290(.A(ori_ori_n226_), .B(i_0_), .Y(ori_ori_n313_));
  NO3        o291(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n314_));
  NA2        o292(.A(ori_ori_n208_), .B(ori_ori_n97_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n315_), .B(ori_ori_n314_), .Y(ori_ori_n316_));
  NA2        o294(.A(i_8_), .B(i_9_), .Y(ori_ori_n317_));
  NA2        o295(.A(ori_ori_n220_), .B(ori_ori_n168_), .Y(ori_ori_n318_));
  OAI220     o296(.A0(ori_ori_n318_), .A1(ori_ori_n317_), .B0(ori_ori_n316_), .B1(ori_ori_n313_), .Y(ori_ori_n319_));
  NA2        o297(.A(ori_ori_n195_), .B(ori_ori_n225_), .Y(ori_ori_n320_));
  NO3        o298(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n321_));
  INV        o299(.A(ori_ori_n321_), .Y(ori_ori_n322_));
  NA3        o300(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n323_));
  NA4        o301(.A(ori_ori_n141_), .B(ori_ori_n114_), .C(ori_ori_n77_), .D(ori_ori_n23_), .Y(ori_ori_n324_));
  OAI220     o302(.A0(ori_ori_n324_), .A1(ori_ori_n323_), .B0(ori_ori_n322_), .B1(ori_ori_n320_), .Y(ori_ori_n325_));
  NO3        o303(.A(ori_ori_n325_), .B(ori_ori_n319_), .C(ori_ori_n312_), .Y(ori_ori_n326_));
  OR2        o304(.A(ori_ori_n243_), .B(ori_ori_n99_), .Y(ori_ori_n327_));
  OR2        o305(.A(ori_ori_n327_), .B(ori_ori_n149_), .Y(ori_ori_n328_));
  NO2        o306(.A(i_2_), .B(i_13_), .Y(ori_ori_n329_));
  NO3        o307(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n330_));
  NO2        o308(.A(i_6_), .B(i_7_), .Y(ori_ori_n331_));
  NO2        o309(.A(i_11_), .B(i_1_), .Y(ori_ori_n332_));
  OR2        o310(.A(i_11_), .B(i_8_), .Y(ori_ori_n333_));
  NOi21      o311(.An(i_2_), .B(i_7_), .Y(ori_ori_n334_));
  NO2        o312(.A(i_3_), .B(ori_ori_n161_), .Y(ori_ori_n335_));
  NO2        o313(.A(i_6_), .B(i_10_), .Y(ori_ori_n336_));
  NA3        o314(.A(ori_ori_n193_), .B(ori_ori_n151_), .C(ori_ori_n131_), .Y(ori_ori_n337_));
  NA2        o315(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n338_));
  NO2        o316(.A(ori_ori_n146_), .B(i_3_), .Y(ori_ori_n339_));
  NAi31      o317(.An(ori_ori_n338_), .B(ori_ori_n339_), .C(ori_ori_n184_), .Y(ori_ori_n340_));
  NA3        o318(.A(ori_ori_n279_), .B(ori_ori_n156_), .C(ori_ori_n144_), .Y(ori_ori_n341_));
  NA3        o319(.A(ori_ori_n341_), .B(ori_ori_n340_), .C(ori_ori_n337_), .Y(ori_ori_n342_));
  INV        o320(.A(ori_ori_n342_), .Y(ori_ori_n343_));
  NA2        o321(.A(ori_ori_n314_), .B(ori_ori_n275_), .Y(ori_ori_n344_));
  NAi21      o322(.An(ori_ori_n177_), .B(ori_ori_n282_), .Y(ori_ori_n345_));
  NA2        o323(.A(ori_ori_n237_), .B(ori_ori_n178_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n346_), .B(ori_ori_n345_), .Y(ori_ori_n347_));
  NA2        o325(.A(ori_ori_n228_), .B(ori_ori_n188_), .Y(ori_ori_n348_));
  NO2        o326(.A(ori_ori_n348_), .B(ori_ori_n301_), .Y(ori_ori_n349_));
  NO2        o327(.A(ori_ori_n349_), .B(ori_ori_n347_), .Y(ori_ori_n350_));
  NA4        o328(.A(ori_ori_n350_), .B(ori_ori_n343_), .C(ori_ori_n328_), .D(ori_ori_n326_), .Y(ori_ori_n351_));
  NA2        o329(.A(ori_ori_n121_), .B(ori_ori_n110_), .Y(ori_ori_n352_));
  AN2        o330(.A(ori_ori_n352_), .B(ori_ori_n314_), .Y(ori_ori_n353_));
  NA2        o331(.A(ori_ori_n353_), .B(ori_ori_n226_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n275_), .B(ori_ori_n183_), .Y(ori_ori_n355_));
  NA2        o333(.A(ori_ori_n248_), .B(ori_ori_n70_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n266_), .B(ori_ori_n258_), .Y(ori_ori_n357_));
  OR2        o335(.A(ori_ori_n355_), .B(ori_ori_n357_), .Y(ori_ori_n358_));
  NO2        o336(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n359_));
  AOI210     o337(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n293_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n360_), .B(ori_ori_n358_), .Y(ori_ori_n361_));
  INV        o339(.A(ori_ori_n361_), .Y(ori_ori_n362_));
  NA2        o340(.A(ori_ori_n200_), .B(ori_ori_n61_), .Y(ori_ori_n363_));
  OAI210     o341(.A0(i_8_), .A1(ori_ori_n363_), .B0(ori_ori_n133_), .Y(ori_ori_n364_));
  NA2        o342(.A(ori_ori_n364_), .B(ori_ori_n294_), .Y(ori_ori_n365_));
  NA3        o343(.A(ori_ori_n365_), .B(ori_ori_n362_), .C(ori_ori_n354_), .Y(ori_ori_n366_));
  NO2        o344(.A(i_12_), .B(ori_ori_n161_), .Y(ori_ori_n367_));
  NO2        o345(.A(i_8_), .B(i_7_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n369_));
  NO2        o347(.A(ori_ori_n369_), .B(i_6_), .Y(ori_ori_n370_));
  NA3        o348(.A(ori_ori_n224_), .B(ori_ori_n153_), .C(ori_ori_n96_), .Y(ori_ori_n371_));
  NO2        o349(.A(ori_ori_n146_), .B(i_5_), .Y(ori_ori_n372_));
  INV        o350(.A(ori_ori_n371_), .Y(ori_ori_n373_));
  NA2        o351(.A(ori_ori_n373_), .B(ori_ori_n321_), .Y(ori_ori_n374_));
  INV        o352(.A(ori_ori_n374_), .Y(ori_ori_n375_));
  NA2        o353(.A(ori_ori_n182_), .B(ori_ori_n181_), .Y(ori_ori_n376_));
  NA2        o354(.A(ori_ori_n307_), .B(ori_ori_n180_), .Y(ori_ori_n377_));
  NO2        o355(.A(ori_ori_n376_), .B(ori_ori_n377_), .Y(ori_ori_n378_));
  AOI210     o356(.A0(ori_ori_n259_), .A1(ori_ori_n46_), .B0(ori_ori_n263_), .Y(ori_ori_n379_));
  NA2        o357(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n380_));
  NA3        o358(.A(ori_ori_n367_), .B(ori_ori_n216_), .C(ori_ori_n380_), .Y(ori_ori_n381_));
  NO2        o359(.A(ori_ori_n379_), .B(ori_ori_n381_), .Y(ori_ori_n382_));
  NO2        o360(.A(ori_ori_n382_), .B(ori_ori_n378_), .Y(ori_ori_n383_));
  NO4        o361(.A(ori_ori_n196_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n384_));
  NO3        o362(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n292_), .B(i_1_), .Y(ori_ori_n386_));
  NOi31      o364(.An(ori_ori_n386_), .B(ori_ori_n315_), .C(ori_ori_n70_), .Y(ori_ori_n387_));
  NOi21      o365(.An(i_10_), .B(i_6_), .Y(ori_ori_n388_));
  NO2        o366(.A(ori_ori_n83_), .B(ori_ori_n25_), .Y(ori_ori_n389_));
  AOI220     o367(.A0(ori_ori_n220_), .A1(ori_ori_n389_), .B0(ori_ori_n216_), .B1(ori_ori_n388_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n390_), .B(ori_ori_n313_), .Y(ori_ori_n391_));
  NO2        o369(.A(ori_ori_n113_), .B(ori_ori_n23_), .Y(ori_ori_n392_));
  INV        o370(.A(ori_ori_n391_), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n356_), .B(ori_ori_n271_), .Y(ori_ori_n394_));
  INV        o372(.A(ori_ori_n229_), .Y(ori_ori_n395_));
  NO2        o373(.A(i_12_), .B(ori_ori_n83_), .Y(ori_ori_n396_));
  NA3        o374(.A(ori_ori_n396_), .B(ori_ori_n216_), .C(ori_ori_n380_), .Y(ori_ori_n397_));
  NA3        o375(.A(ori_ori_n277_), .B(ori_ori_n220_), .C(ori_ori_n178_), .Y(ori_ori_n398_));
  AOI210     o376(.A0(ori_ori_n398_), .A1(ori_ori_n397_), .B0(ori_ori_n395_), .Y(ori_ori_n399_));
  OR2        o377(.A(i_2_), .B(i_5_), .Y(ori_ori_n400_));
  NA2        o378(.A(ori_ori_n267_), .B(ori_ori_n192_), .Y(ori_ori_n401_));
  NO2        o379(.A(ori_ori_n401_), .B(ori_ori_n345_), .Y(ori_ori_n402_));
  NO3        o380(.A(ori_ori_n402_), .B(ori_ori_n399_), .C(ori_ori_n394_), .Y(ori_ori_n403_));
  NA3        o381(.A(ori_ori_n403_), .B(ori_ori_n393_), .C(ori_ori_n383_), .Y(ori_ori_n404_));
  NO4        o382(.A(ori_ori_n404_), .B(ori_ori_n375_), .C(ori_ori_n366_), .D(ori_ori_n351_), .Y(ori_ori_n405_));
  NA4        o383(.A(ori_ori_n405_), .B(ori_ori_n305_), .C(ori_ori_n247_), .D(ori_ori_n227_), .Y(ori7));
  NO2        o384(.A(ori_ori_n92_), .B(ori_ori_n54_), .Y(ori_ori_n407_));
  NO2        o385(.A(ori_ori_n106_), .B(ori_ori_n89_), .Y(ori_ori_n408_));
  NA2        o386(.A(i_3_), .B(ori_ori_n408_), .Y(ori_ori_n409_));
  NA2        o387(.A(ori_ori_n336_), .B(ori_ori_n81_), .Y(ori_ori_n410_));
  NA2        o388(.A(i_11_), .B(ori_ori_n161_), .Y(ori_ori_n411_));
  NA2        o389(.A(ori_ori_n140_), .B(ori_ori_n411_), .Y(ori_ori_n412_));
  OAI210     o390(.A0(ori_ori_n412_), .A1(ori_ori_n410_), .B0(ori_ori_n409_), .Y(ori_ori_n413_));
  NO2        o391(.A(ori_ori_n187_), .B(i_4_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n414_), .B(i_8_), .Y(ori_ori_n415_));
  NA2        o393(.A(i_2_), .B(ori_ori_n83_), .Y(ori_ori_n416_));
  OAI210     o394(.A0(ori_ori_n86_), .A1(ori_ori_n165_), .B0(ori_ori_n166_), .Y(ori_ori_n417_));
  NO2        o395(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n418_));
  NA2        o396(.A(i_4_), .B(i_8_), .Y(ori_ori_n419_));
  AOI210     o397(.A0(ori_ori_n419_), .A1(ori_ori_n224_), .B0(ori_ori_n418_), .Y(ori_ori_n420_));
  OAI220     o398(.A0(ori_ori_n420_), .A1(ori_ori_n416_), .B0(ori_ori_n417_), .B1(i_13_), .Y(ori_ori_n421_));
  NO3        o399(.A(ori_ori_n421_), .B(ori_ori_n413_), .C(ori_ori_n407_), .Y(ori_ori_n422_));
  AOI210     o400(.A0(ori_ori_n127_), .A1(ori_ori_n59_), .B0(i_10_), .Y(ori_ori_n423_));
  AOI210     o401(.A0(ori_ori_n423_), .A1(ori_ori_n187_), .B0(ori_ori_n148_), .Y(ori_ori_n424_));
  OR2        o402(.A(i_6_), .B(i_10_), .Y(ori_ori_n425_));
  OR3        o403(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n426_));
  INV        o404(.A(ori_ori_n164_), .Y(ori_ori_n427_));
  OR2        o405(.A(ori_ori_n424_), .B(ori_ori_n209_), .Y(ori_ori_n428_));
  AOI210     o406(.A0(ori_ori_n428_), .A1(ori_ori_n422_), .B0(ori_ori_n60_), .Y(ori_ori_n429_));
  NOi21      o407(.An(i_11_), .B(i_7_), .Y(ori_ori_n430_));
  AO210      o408(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n431_));
  NO2        o409(.A(ori_ori_n431_), .B(ori_ori_n430_), .Y(ori_ori_n432_));
  NA2        o410(.A(ori_ori_n432_), .B(ori_ori_n170_), .Y(ori_ori_n433_));
  NA3        o411(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n434_));
  NAi31      o412(.An(ori_ori_n434_), .B(ori_ori_n176_), .C(i_11_), .Y(ori_ori_n435_));
  AOI210     o413(.A0(ori_ori_n435_), .A1(ori_ori_n433_), .B0(ori_ori_n60_), .Y(ori_ori_n436_));
  NA2        o414(.A(ori_ori_n85_), .B(ori_ori_n60_), .Y(ori_ori_n437_));
  AO210      o415(.A0(ori_ori_n437_), .A1(ori_ori_n271_), .B0(ori_ori_n41_), .Y(ori_ori_n438_));
  NO3        o416(.A(ori_ori_n202_), .B(ori_ori_n171_), .C(ori_ori_n411_), .Y(ori_ori_n439_));
  OAI210     o417(.A0(ori_ori_n439_), .A1(ori_ori_n184_), .B0(ori_ori_n60_), .Y(ori_ori_n440_));
  NA2        o418(.A(ori_ori_n290_), .B(ori_ori_n31_), .Y(ori_ori_n441_));
  OR2        o419(.A(ori_ori_n171_), .B(ori_ori_n106_), .Y(ori_ori_n442_));
  NA2        o420(.A(ori_ori_n442_), .B(ori_ori_n441_), .Y(ori_ori_n443_));
  NO2        o421(.A(i_1_), .B(i_4_), .Y(ori_ori_n444_));
  NA2        o422(.A(ori_ori_n444_), .B(ori_ori_n443_), .Y(ori_ori_n445_));
  NO2        o423(.A(i_1_), .B(i_12_), .Y(ori_ori_n446_));
  NA3        o424(.A(ori_ori_n446_), .B(ori_ori_n108_), .C(ori_ori_n24_), .Y(ori_ori_n447_));
  BUFFER     o425(.A(ori_ori_n447_), .Y(ori_ori_n448_));
  NA4        o426(.A(ori_ori_n448_), .B(ori_ori_n445_), .C(ori_ori_n440_), .D(ori_ori_n438_), .Y(ori_ori_n449_));
  OAI210     o427(.A0(ori_ori_n449_), .A1(ori_ori_n436_), .B0(i_6_), .Y(ori_ori_n450_));
  NO2        o428(.A(ori_ori_n434_), .B(ori_ori_n106_), .Y(ori_ori_n451_));
  NA2        o429(.A(ori_ori_n451_), .B(ori_ori_n396_), .Y(ori_ori_n452_));
  NO2        o430(.A(i_6_), .B(i_11_), .Y(ori_ori_n453_));
  NA2        o431(.A(ori_ori_n452_), .B(ori_ori_n316_), .Y(ori_ori_n454_));
  NO3        o432(.A(ori_ori_n425_), .B(ori_ori_n186_), .C(ori_ori_n23_), .Y(ori_ori_n455_));
  AOI210     o433(.A0(i_1_), .A1(ori_ori_n203_), .B0(ori_ori_n455_), .Y(ori_ori_n456_));
  NO2        o434(.A(ori_ori_n456_), .B(ori_ori_n44_), .Y(ori_ori_n457_));
  NA3        o435(.A(ori_ori_n368_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n458_));
  INV        o436(.A(i_2_), .Y(ori_ori_n459_));
  NA2        o437(.A(ori_ori_n137_), .B(i_9_), .Y(ori_ori_n460_));
  NA3        o438(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n461_));
  NO2        o439(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n462_));
  NA3        o440(.A(ori_ori_n462_), .B(ori_ori_n208_), .C(ori_ori_n44_), .Y(ori_ori_n463_));
  OAI220     o441(.A0(ori_ori_n463_), .A1(ori_ori_n461_), .B0(ori_ori_n460_), .B1(ori_ori_n459_), .Y(ori_ori_n464_));
  AOI210     o442(.A0(ori_ori_n332_), .A1(ori_ori_n295_), .B0(ori_ori_n190_), .Y(ori_ori_n465_));
  NO2        o443(.A(ori_ori_n465_), .B(ori_ori_n416_), .Y(ori_ori_n466_));
  NAi21      o444(.An(ori_ori_n458_), .B(ori_ori_n91_), .Y(ori_ori_n467_));
  NO2        o445(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n468_));
  INV        o446(.A(ori_ori_n467_), .Y(ori_ori_n469_));
  OR3        o447(.A(ori_ori_n469_), .B(ori_ori_n466_), .C(ori_ori_n464_), .Y(ori_ori_n470_));
  NO3        o448(.A(ori_ori_n470_), .B(ori_ori_n457_), .C(ori_ori_n454_), .Y(ori_ori_n471_));
  NO2        o449(.A(ori_ori_n187_), .B(ori_ori_n99_), .Y(ori_ori_n472_));
  NO2        o450(.A(ori_ori_n472_), .B(ori_ori_n430_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n473_), .B(i_1_), .Y(ori_ori_n474_));
  NO2        o452(.A(ori_ori_n474_), .B(ori_ori_n426_), .Y(ori_ori_n475_));
  NA2        o453(.A(ori_ori_n475_), .B(ori_ori_n46_), .Y(ori_ori_n476_));
  NA2        o454(.A(i_3_), .B(ori_ori_n161_), .Y(ori_ori_n477_));
  NO2        o455(.A(ori_ori_n477_), .B(ori_ori_n113_), .Y(ori_ori_n478_));
  AN2        o456(.A(ori_ori_n478_), .B(ori_ori_n370_), .Y(ori_ori_n479_));
  NO2        o457(.A(ori_ori_n116_), .B(ori_ori_n37_), .Y(ori_ori_n480_));
  NA2        o458(.A(i_1_), .B(i_3_), .Y(ori_ori_n481_));
  NO2        o459(.A(ori_ori_n317_), .B(ori_ori_n92_), .Y(ori_ori_n482_));
  INV        o460(.A(ori_ori_n482_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n483_), .B(ori_ori_n481_), .Y(ori_ori_n484_));
  NO2        o462(.A(ori_ori_n484_), .B(ori_ori_n479_), .Y(ori_ori_n485_));
  NA4        o463(.A(ori_ori_n485_), .B(ori_ori_n476_), .C(ori_ori_n471_), .D(ori_ori_n450_), .Y(ori_ori_n486_));
  NA2        o464(.A(ori_ori_n266_), .B(ori_ori_n265_), .Y(ori_ori_n487_));
  NO3        o465(.A(ori_ori_n334_), .B(ori_ori_n419_), .C(ori_ori_n83_), .Y(ori_ori_n488_));
  NA2        o466(.A(ori_ori_n488_), .B(ori_ori_n25_), .Y(ori_ori_n489_));
  NA2        o467(.A(ori_ori_n489_), .B(ori_ori_n487_), .Y(ori_ori_n490_));
  NA2        o468(.A(ori_ori_n490_), .B(i_1_), .Y(ori_ori_n491_));
  AOI210     o469(.A0(ori_ori_n208_), .A1(ori_ori_n97_), .B0(i_1_), .Y(ori_ori_n492_));
  NO2        o470(.A(ori_ori_n264_), .B(i_2_), .Y(ori_ori_n493_));
  NA2        o471(.A(ori_ori_n493_), .B(ori_ori_n492_), .Y(ori_ori_n494_));
  AOI210     o472(.A0(ori_ori_n494_), .A1(ori_ori_n491_), .B0(i_13_), .Y(ori_ori_n495_));
  OR2        o473(.A(i_11_), .B(i_7_), .Y(ori_ori_n496_));
  NA3        o474(.A(ori_ori_n496_), .B(ori_ori_n104_), .C(ori_ori_n137_), .Y(ori_ori_n497_));
  AOI220     o475(.A0(ori_ori_n329_), .A1(ori_ori_n148_), .B0(ori_ori_n310_), .B1(ori_ori_n137_), .Y(ori_ori_n498_));
  OAI210     o476(.A0(ori_ori_n498_), .A1(ori_ori_n44_), .B0(ori_ori_n497_), .Y(ori_ori_n499_));
  NO2        o477(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n500_));
  NO2        o478(.A(ori_ori_n334_), .B(ori_ori_n24_), .Y(ori_ori_n501_));
  NO2        o479(.A(ori_ori_n752_), .B(ori_ori_n92_), .Y(ori_ori_n502_));
  AOI210     o480(.A0(ori_ori_n499_), .A1(ori_ori_n236_), .B0(ori_ori_n502_), .Y(ori_ori_n503_));
  INV        o481(.A(ori_ori_n113_), .Y(ori_ori_n504_));
  AOI220     o482(.A0(ori_ori_n504_), .A1(ori_ori_n69_), .B0(ori_ori_n277_), .B1(ori_ori_n462_), .Y(ori_ori_n505_));
  NO2        o483(.A(ori_ori_n505_), .B(ori_ori_n191_), .Y(ori_ori_n506_));
  NA2        o484(.A(ori_ori_n126_), .B(i_13_), .Y(ori_ori_n507_));
  NO2        o485(.A(ori_ori_n461_), .B(ori_ori_n113_), .Y(ori_ori_n508_));
  INV        o486(.A(ori_ori_n508_), .Y(ori_ori_n509_));
  OAI220     o487(.A0(ori_ori_n509_), .A1(ori_ori_n68_), .B0(ori_ori_n507_), .B1(ori_ori_n492_), .Y(ori_ori_n510_));
  NO3        o488(.A(ori_ori_n68_), .B(ori_ori_n32_), .C(ori_ori_n99_), .Y(ori_ori_n511_));
  NA2        o489(.A(ori_ori_n26_), .B(ori_ori_n161_), .Y(ori_ori_n512_));
  NA2        o490(.A(ori_ori_n512_), .B(i_7_), .Y(ori_ori_n513_));
  NO3        o491(.A(ori_ori_n334_), .B(ori_ori_n187_), .C(ori_ori_n83_), .Y(ori_ori_n514_));
  AOI210     o492(.A0(ori_ori_n514_), .A1(ori_ori_n513_), .B0(ori_ori_n511_), .Y(ori_ori_n515_));
  AOI220     o493(.A0(ori_ori_n277_), .A1(ori_ori_n462_), .B0(ori_ori_n91_), .B1(ori_ori_n100_), .Y(ori_ori_n516_));
  OAI220     o494(.A0(ori_ori_n516_), .A1(ori_ori_n415_), .B0(ori_ori_n515_), .B1(ori_ori_n427_), .Y(ori_ori_n517_));
  NO3        o495(.A(ori_ori_n517_), .B(ori_ori_n510_), .C(ori_ori_n506_), .Y(ori_ori_n518_));
  OR2        o496(.A(i_11_), .B(i_6_), .Y(ori_ori_n519_));
  NA3        o497(.A(ori_ori_n414_), .B(ori_ori_n512_), .C(i_7_), .Y(ori_ori_n520_));
  AOI210     o498(.A0(ori_ori_n520_), .A1(ori_ori_n509_), .B0(ori_ori_n519_), .Y(ori_ori_n521_));
  NA3        o499(.A(ori_ori_n290_), .B(ori_ori_n418_), .C(ori_ori_n97_), .Y(ori_ori_n522_));
  NA2        o500(.A(ori_ori_n453_), .B(i_13_), .Y(ori_ori_n523_));
  NAi21      o501(.An(i_11_), .B(i_12_), .Y(ori_ori_n524_));
  NO3        o502(.A(ori_ori_n334_), .B(ori_ori_n396_), .C(ori_ori_n419_), .Y(ori_ori_n525_));
  NA2        o503(.A(ori_ori_n525_), .B(ori_ori_n228_), .Y(ori_ori_n526_));
  NA3        o504(.A(ori_ori_n526_), .B(ori_ori_n523_), .C(ori_ori_n522_), .Y(ori_ori_n527_));
  OAI210     o505(.A0(ori_ori_n527_), .A1(ori_ori_n521_), .B0(ori_ori_n60_), .Y(ori_ori_n528_));
  NO2        o506(.A(i_2_), .B(i_12_), .Y(ori_ori_n529_));
  NA2        o507(.A(ori_ori_n263_), .B(ori_ori_n529_), .Y(ori_ori_n530_));
  NO2        o508(.A(ori_ori_n127_), .B(i_2_), .Y(ori_ori_n531_));
  NA2        o509(.A(ori_ori_n531_), .B(ori_ori_n446_), .Y(ori_ori_n532_));
  NA2        o510(.A(ori_ori_n532_), .B(ori_ori_n530_), .Y(ori_ori_n533_));
  NA3        o511(.A(ori_ori_n533_), .B(ori_ori_n45_), .C(ori_ori_n183_), .Y(ori_ori_n534_));
  NA4        o512(.A(ori_ori_n534_), .B(ori_ori_n528_), .C(ori_ori_n518_), .D(ori_ori_n503_), .Y(ori_ori_n535_));
  OR4        o513(.A(ori_ori_n535_), .B(ori_ori_n495_), .C(ori_ori_n486_), .D(ori_ori_n429_), .Y(ori5));
  NA2        o514(.A(ori_ori_n473_), .B(ori_ori_n211_), .Y(ori_ori_n537_));
  AN2        o515(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n538_));
  NA3        o516(.A(ori_ori_n538_), .B(ori_ori_n529_), .C(ori_ori_n106_), .Y(ori_ori_n539_));
  NO2        o517(.A(ori_ori_n415_), .B(i_11_), .Y(ori_ori_n540_));
  NA2        o518(.A(ori_ori_n86_), .B(ori_ori_n540_), .Y(ori_ori_n541_));
  NA3        o519(.A(ori_ori_n541_), .B(ori_ori_n539_), .C(ori_ori_n537_), .Y(ori_ori_n542_));
  NO3        o520(.A(i_11_), .B(ori_ori_n187_), .C(i_13_), .Y(ori_ori_n543_));
  NO2        o521(.A(ori_ori_n123_), .B(ori_ori_n23_), .Y(ori_ori_n544_));
  NA2        o522(.A(i_12_), .B(i_8_), .Y(ori_ori_n545_));
  OAI210     o523(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n545_), .Y(ori_ori_n546_));
  INV        o524(.A(ori_ori_n307_), .Y(ori_ori_n547_));
  AOI220     o525(.A0(ori_ori_n229_), .A1(ori_ori_n392_), .B0(ori_ori_n546_), .B1(ori_ori_n544_), .Y(ori_ori_n548_));
  INV        o526(.A(ori_ori_n548_), .Y(ori_ori_n549_));
  NO2        o527(.A(ori_ori_n549_), .B(ori_ori_n542_), .Y(ori_ori_n550_));
  INV        o528(.A(ori_ori_n151_), .Y(ori_ori_n551_));
  INV        o529(.A(ori_ori_n193_), .Y(ori_ori_n552_));
  OAI210     o530(.A0(ori_ori_n493_), .A1(ori_ori_n309_), .B0(ori_ori_n109_), .Y(ori_ori_n553_));
  AOI210     o531(.A0(ori_ori_n553_), .A1(ori_ori_n552_), .B0(ori_ori_n551_), .Y(ori_ori_n554_));
  NO2        o532(.A(ori_ori_n317_), .B(ori_ori_n26_), .Y(ori_ori_n555_));
  NO2        o533(.A(ori_ori_n555_), .B(ori_ori_n295_), .Y(ori_ori_n556_));
  NA2        o534(.A(ori_ori_n556_), .B(i_2_), .Y(ori_ori_n557_));
  INV        o535(.A(ori_ori_n557_), .Y(ori_ori_n558_));
  AOI210     o536(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n292_), .Y(ori_ori_n559_));
  AOI210     o537(.A0(ori_ori_n559_), .A1(ori_ori_n558_), .B0(ori_ori_n554_), .Y(ori_ori_n560_));
  NO2        o538(.A(ori_ori_n160_), .B(ori_ori_n124_), .Y(ori_ori_n561_));
  OAI210     o539(.A0(ori_ori_n561_), .A1(ori_ori_n544_), .B0(i_2_), .Y(ori_ori_n562_));
  INV        o540(.A(ori_ori_n152_), .Y(ori_ori_n563_));
  NO3        o541(.A(ori_ori_n431_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n564_));
  AOI210     o542(.A0(ori_ori_n563_), .A1(ori_ori_n86_), .B0(ori_ori_n564_), .Y(ori_ori_n565_));
  AOI210     o543(.A0(ori_ori_n565_), .A1(ori_ori_n562_), .B0(ori_ori_n161_), .Y(ori_ori_n566_));
  OA210      o544(.A0(ori_ori_n432_), .A1(ori_ori_n125_), .B0(i_13_), .Y(ori_ori_n567_));
  NA2        o545(.A(ori_ori_n164_), .B(ori_ori_n165_), .Y(ori_ori_n568_));
  NO2        o546(.A(ori_ori_n568_), .B(ori_ori_n267_), .Y(ori_ori_n569_));
  AOI210     o547(.A0(ori_ori_n171_), .A1(ori_ori_n143_), .B0(ori_ori_n359_), .Y(ori_ori_n570_));
  NA2        o548(.A(ori_ori_n570_), .B(ori_ori_n295_), .Y(ori_ori_n571_));
  NO2        o549(.A(ori_ori_n100_), .B(ori_ori_n44_), .Y(ori_ori_n572_));
  INV        o550(.A(ori_ori_n223_), .Y(ori_ori_n573_));
  NA4        o551(.A(ori_ori_n573_), .B(ori_ori_n224_), .C(ori_ori_n123_), .D(ori_ori_n42_), .Y(ori_ori_n574_));
  OAI210     o552(.A0(ori_ori_n574_), .A1(ori_ori_n572_), .B0(ori_ori_n571_), .Y(ori_ori_n575_));
  NO4        o553(.A(ori_ori_n575_), .B(ori_ori_n569_), .C(ori_ori_n567_), .D(ori_ori_n566_), .Y(ori_ori_n576_));
  NA2        o554(.A(ori_ori_n392_), .B(ori_ori_n28_), .Y(ori_ori_n577_));
  NA2        o555(.A(ori_ori_n543_), .B(ori_ori_n217_), .Y(ori_ori_n578_));
  NA2        o556(.A(ori_ori_n578_), .B(ori_ori_n577_), .Y(ori_ori_n579_));
  NO2        o557(.A(ori_ori_n59_), .B(i_12_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n580_), .B(ori_ori_n125_), .Y(ori_ori_n581_));
  NO2        o559(.A(ori_ori_n581_), .B(ori_ori_n411_), .Y(ori_ori_n582_));
  AOI220     o560(.A0(ori_ori_n582_), .A1(ori_ori_n36_), .B0(ori_ori_n579_), .B1(ori_ori_n46_), .Y(ori_ori_n583_));
  NA4        o561(.A(ori_ori_n583_), .B(ori_ori_n576_), .C(ori_ori_n560_), .D(ori_ori_n550_), .Y(ori6));
  NA4        o562(.A(ori_ori_n278_), .B(ori_ori_n335_), .C(ori_ori_n68_), .D(ori_ori_n99_), .Y(ori_ori_n585_));
  INV        o563(.A(ori_ori_n585_), .Y(ori_ori_n586_));
  NO2        o564(.A(ori_ori_n179_), .B(ori_ori_n338_), .Y(ori_ori_n587_));
  NO2        o565(.A(i_11_), .B(i_9_), .Y(ori_ori_n588_));
  NO2        o566(.A(ori_ori_n586_), .B(ori_ori_n232_), .Y(ori_ori_n589_));
  OR2        o567(.A(ori_ori_n589_), .B(i_12_), .Y(ori_ori_n590_));
  NA2        o568(.A(ori_ori_n396_), .B(ori_ori_n60_), .Y(ori_ori_n591_));
  BUFFER     o569(.A(ori_ori_n437_), .Y(ori_ori_n592_));
  NA2        o570(.A(ori_ori_n592_), .B(ori_ori_n591_), .Y(ori_ori_n593_));
  INV        o571(.A(ori_ori_n163_), .Y(ori_ori_n594_));
  AOI220     o572(.A0(ori_ori_n594_), .A1(ori_ori_n588_), .B0(ori_ori_n593_), .B1(ori_ori_n70_), .Y(ori_ori_n595_));
  INV        o573(.A(ori_ori_n231_), .Y(ori_ori_n596_));
  NA2        o574(.A(ori_ori_n72_), .B(ori_ori_n130_), .Y(ori_ori_n597_));
  INV        o575(.A(ori_ori_n123_), .Y(ori_ori_n598_));
  NA2        o576(.A(ori_ori_n598_), .B(ori_ori_n46_), .Y(ori_ori_n599_));
  AOI210     o577(.A0(ori_ori_n599_), .A1(ori_ori_n597_), .B0(ori_ori_n596_), .Y(ori_ori_n600_));
  NO2        o578(.A(ori_ori_n196_), .B(i_9_), .Y(ori_ori_n601_));
  NA2        o579(.A(ori_ori_n601_), .B(ori_ori_n580_), .Y(ori_ori_n602_));
  AOI210     o580(.A0(ori_ori_n602_), .A1(ori_ori_n357_), .B0(ori_ori_n157_), .Y(ori_ori_n603_));
  NO2        o581(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n604_));
  NAi32      o582(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n605_));
  NO2        o583(.A(ori_ori_n519_), .B(ori_ori_n605_), .Y(ori_ori_n606_));
  OR3        o584(.A(ori_ori_n606_), .B(ori_ori_n603_), .C(ori_ori_n600_), .Y(ori_ori_n607_));
  NO2        o585(.A(ori_ori_n496_), .B(i_2_), .Y(ori_ori_n608_));
  OR2        o586(.A(ori_ori_n432_), .B(ori_ori_n309_), .Y(ori_ori_n609_));
  NA3        o587(.A(ori_ori_n609_), .B(ori_ori_n142_), .C(ori_ori_n66_), .Y(ori_ori_n610_));
  OR2        o588(.A(ori_ori_n547_), .B(ori_ori_n36_), .Y(ori_ori_n611_));
  NA2        o589(.A(ori_ori_n611_), .B(ori_ori_n610_), .Y(ori_ori_n612_));
  OAI210     o590(.A0(i_6_), .A1(i_11_), .B0(ori_ori_n84_), .Y(ori_ori_n613_));
  AOI220     o591(.A0(ori_ori_n613_), .A1(ori_ori_n385_), .B0(ori_ori_n587_), .B1(ori_ori_n513_), .Y(ori_ori_n614_));
  NA3        o592(.A(ori_ori_n267_), .B(ori_ori_n188_), .C(ori_ori_n142_), .Y(ori_ori_n615_));
  NA2        o593(.A(ori_ori_n280_), .B(ori_ori_n67_), .Y(ori_ori_n616_));
  NA4        o594(.A(ori_ori_n616_), .B(ori_ori_n615_), .C(ori_ori_n614_), .D(ori_ori_n417_), .Y(ori_ori_n617_));
  AO210      o595(.A0(ori_ori_n359_), .A1(ori_ori_n46_), .B0(ori_ori_n85_), .Y(ori_ori_n618_));
  NA3        o596(.A(ori_ori_n618_), .B(ori_ori_n336_), .C(ori_ori_n178_), .Y(ori_ori_n619_));
  AOI210     o597(.A0(ori_ori_n309_), .A1(ori_ori_n307_), .B0(ori_ori_n384_), .Y(ori_ori_n620_));
  NO2        o598(.A(ori_ori_n425_), .B(ori_ori_n100_), .Y(ori_ori_n621_));
  OAI210     o599(.A0(ori_ori_n621_), .A1(ori_ori_n110_), .B0(ori_ori_n289_), .Y(ori_ori_n622_));
  NA3        o600(.A(ori_ori_n622_), .B(ori_ori_n620_), .C(ori_ori_n619_), .Y(ori_ori_n623_));
  NO4        o601(.A(ori_ori_n623_), .B(ori_ori_n617_), .C(ori_ori_n612_), .D(ori_ori_n607_), .Y(ori_ori_n624_));
  NA4        o602(.A(ori_ori_n624_), .B(ori_ori_n595_), .C(ori_ori_n590_), .D(ori_ori_n273_), .Y(ori3));
  NA2        o603(.A(i_12_), .B(i_10_), .Y(ori_ori_n626_));
  NA2        o604(.A(ori_ori_n615_), .B(ori_ori_n417_), .Y(ori_ori_n627_));
  NA2        o605(.A(ori_ori_n627_), .B(ori_ori_n40_), .Y(ori_ori_n628_));
  NOi21      o606(.An(ori_ori_n96_), .B(ori_ori_n556_), .Y(ori_ori_n629_));
  NO3        o607(.A(ori_ori_n442_), .B(ori_ori_n317_), .C(ori_ori_n130_), .Y(ori_ori_n630_));
  NA2        o608(.A(ori_ori_n290_), .B(ori_ori_n45_), .Y(ori_ori_n631_));
  AN2        o609(.A(ori_ori_n315_), .B(ori_ori_n55_), .Y(ori_ori_n632_));
  NO3        o610(.A(ori_ori_n632_), .B(ori_ori_n630_), .C(ori_ori_n629_), .Y(ori_ori_n633_));
  AOI210     o611(.A0(ori_ori_n633_), .A1(ori_ori_n628_), .B0(ori_ori_n48_), .Y(ori_ori_n634_));
  NO4        o612(.A(ori_ori_n269_), .B(ori_ori_n275_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n635_));
  NA2        o613(.A(ori_ori_n157_), .B(ori_ori_n388_), .Y(ori_ori_n636_));
  NOi21      o614(.An(ori_ori_n636_), .B(ori_ori_n635_), .Y(ori_ori_n637_));
  NO2        o615(.A(ori_ori_n637_), .B(ori_ori_n60_), .Y(ori_ori_n638_));
  NOi21      o616(.An(i_5_), .B(i_9_), .Y(ori_ori_n639_));
  NA2        o617(.A(ori_ori_n639_), .B(ori_ori_n306_), .Y(ori_ori_n640_));
  BUFFER     o618(.A(ori_ori_n208_), .Y(ori_ori_n641_));
  AOI210     o619(.A0(ori_ori_n641_), .A1(ori_ori_n332_), .B0(ori_ori_n488_), .Y(ori_ori_n642_));
  NO2        o620(.A(ori_ori_n642_), .B(ori_ori_n640_), .Y(ori_ori_n643_));
  NO3        o621(.A(ori_ori_n643_), .B(ori_ori_n638_), .C(ori_ori_n634_), .Y(ori_ori_n644_));
  NA2        o622(.A(ori_ori_n157_), .B(ori_ori_n24_), .Y(ori_ori_n645_));
  NO2        o623(.A(ori_ori_n480_), .B(ori_ori_n408_), .Y(ori_ori_n646_));
  NO2        o624(.A(ori_ori_n646_), .B(ori_ori_n645_), .Y(ori_ori_n647_));
  INV        o625(.A(ori_ori_n647_), .Y(ori_ori_n648_));
  NA2        o626(.A(ori_ori_n389_), .B(i_0_), .Y(ori_ori_n649_));
  NO3        o627(.A(ori_ori_n649_), .B(ori_ori_n276_), .C(ori_ori_n86_), .Y(ori_ori_n650_));
  NO4        o628(.A(ori_ori_n400_), .B(ori_ori_n176_), .C(ori_ori_n292_), .D(i_6_), .Y(ori_ori_n651_));
  AOI210     o629(.A0(ori_ori_n651_), .A1(i_11_), .B0(ori_ori_n650_), .Y(ori_ori_n652_));
  NA2        o630(.A(ori_ori_n543_), .B(ori_ori_n232_), .Y(ori_ori_n653_));
  AOI210     o631(.A0(ori_ori_n336_), .A1(ori_ori_n86_), .B0(ori_ori_n57_), .Y(ori_ori_n654_));
  NO2        o632(.A(ori_ori_n654_), .B(ori_ori_n653_), .Y(ori_ori_n655_));
  NO2        o633(.A(ori_ori_n198_), .B(ori_ori_n145_), .Y(ori_ori_n656_));
  NA2        o634(.A(i_0_), .B(i_10_), .Y(ori_ori_n657_));
  INV        o635(.A(ori_ori_n369_), .Y(ori_ori_n658_));
  NO4        o636(.A(ori_ori_n113_), .B(ori_ori_n57_), .C(ori_ori_n477_), .D(i_5_), .Y(ori_ori_n659_));
  AO220      o637(.A0(ori_ori_n659_), .A1(ori_ori_n658_), .B0(ori_ori_n656_), .B1(i_6_), .Y(ori_ori_n660_));
  NO2        o638(.A(ori_ori_n660_), .B(ori_ori_n655_), .Y(ori_ori_n661_));
  NA3        o639(.A(ori_ori_n661_), .B(ori_ori_n652_), .C(ori_ori_n648_), .Y(ori_ori_n662_));
  NO2        o640(.A(ori_ori_n101_), .B(ori_ori_n37_), .Y(ori_ori_n663_));
  NA2        o641(.A(i_11_), .B(i_9_), .Y(ori_ori_n664_));
  NO3        o642(.A(i_12_), .B(ori_ori_n664_), .C(ori_ori_n416_), .Y(ori_ori_n665_));
  AN2        o643(.A(ori_ori_n665_), .B(ori_ori_n663_), .Y(ori_ori_n666_));
  NA2        o644(.A(ori_ori_n279_), .B(ori_ori_n156_), .Y(ori_ori_n667_));
  INV        o645(.A(ori_ori_n667_), .Y(ori_ori_n668_));
  NO2        o646(.A(ori_ori_n664_), .B(ori_ori_n70_), .Y(ori_ori_n669_));
  NO2        o647(.A(ori_ori_n668_), .B(ori_ori_n666_), .Y(ori_ori_n670_));
  NA2        o648(.A(ori_ori_n468_), .B(ori_ori_n120_), .Y(ori_ori_n671_));
  NO2        o649(.A(i_6_), .B(ori_ori_n671_), .Y(ori_ori_n672_));
  NA2        o650(.A(ori_ori_n151_), .B(ori_ori_n101_), .Y(ori_ori_n673_));
  NA2        o651(.A(ori_ori_n418_), .B(ori_ori_n232_), .Y(ori_ori_n674_));
  NO2        o652(.A(ori_ori_n674_), .B(ori_ori_n631_), .Y(ori_ori_n675_));
  NO2        o653(.A(ori_ori_n675_), .B(ori_ori_n672_), .Y(ori_ori_n676_));
  INV        o654(.A(ori_ori_n230_), .Y(ori_ori_n677_));
  NA2        o655(.A(ori_ori_n676_), .B(ori_ori_n670_), .Y(ori_ori_n678_));
  NO2        o656(.A(ori_ori_n626_), .B(ori_ori_n229_), .Y(ori_ori_n679_));
  OA210      o657(.A0(ori_ori_n331_), .A1(ori_ori_n182_), .B0(ori_ori_n330_), .Y(ori_ori_n680_));
  NA2        o658(.A(ori_ori_n679_), .B(ori_ori_n669_), .Y(ori_ori_n681_));
  NA2        o659(.A(ori_ori_n669_), .B(ori_ori_n224_), .Y(ori_ori_n682_));
  INV        o660(.A(ori_ori_n682_), .Y(ori_ori_n683_));
  NA2        o661(.A(ori_ori_n683_), .B(ori_ori_n331_), .Y(ori_ori_n684_));
  NO3        o662(.A(ori_ori_n400_), .B(ori_ori_n250_), .C(ori_ori_n24_), .Y(ori_ori_n685_));
  AOI210     o663(.A0(ori_ori_n501_), .A1(ori_ori_n372_), .B0(ori_ori_n685_), .Y(ori_ori_n686_));
  NAi21      o664(.An(i_9_), .B(i_5_), .Y(ori_ori_n687_));
  NO2        o665(.A(ori_ori_n687_), .B(ori_ori_n285_), .Y(ori_ori_n688_));
  NA2        o666(.A(ori_ori_n688_), .B(ori_ori_n432_), .Y(ori_ori_n689_));
  OAI220     o667(.A0(ori_ori_n689_), .A1(ori_ori_n83_), .B0(ori_ori_n686_), .B1(ori_ori_n152_), .Y(ori_ori_n690_));
  NO2        o668(.A(ori_ori_n690_), .B(ori_ori_n361_), .Y(ori_ori_n691_));
  NA3        o669(.A(ori_ori_n691_), .B(ori_ori_n684_), .C(ori_ori_n681_), .Y(ori_ori_n692_));
  NO3        o670(.A(ori_ori_n692_), .B(ori_ori_n678_), .C(ori_ori_n662_), .Y(ori_ori_n693_));
  NO2        o671(.A(i_0_), .B(ori_ori_n524_), .Y(ori_ori_n694_));
  AOI210     o672(.A0(ori_ori_n591_), .A1(ori_ori_n487_), .B0(ori_ori_n673_), .Y(ori_ori_n695_));
  INV        o673(.A(ori_ori_n695_), .Y(ori_ori_n696_));
  NA2        o674(.A(ori_ori_n192_), .B(ori_ori_n185_), .Y(ori_ori_n697_));
  AOI210     o675(.A0(ori_ori_n697_), .A1(ori_ori_n649_), .B0(ori_ori_n145_), .Y(ori_ori_n698_));
  INV        o676(.A(ori_ori_n698_), .Y(ori_ori_n699_));
  NA2        o677(.A(ori_ori_n699_), .B(ori_ori_n696_), .Y(ori_ori_n700_));
  NO3        o678(.A(ori_ori_n657_), .B(ori_ori_n639_), .C(ori_ori_n160_), .Y(ori_ori_n701_));
  AOI220     o679(.A0(ori_ori_n701_), .A1(i_11_), .B0(ori_ori_n387_), .B1(ori_ori_n72_), .Y(ori_ori_n702_));
  NO3        o680(.A(ori_ori_n172_), .B(ori_ori_n275_), .C(i_0_), .Y(ori_ori_n703_));
  OAI210     o681(.A0(ori_ori_n703_), .A1(ori_ori_n73_), .B0(i_13_), .Y(ori_ori_n704_));
  NA2        o682(.A(ori_ori_n704_), .B(ori_ori_n702_), .Y(ori_ori_n705_));
  INV        o683(.A(ori_ori_n92_), .Y(ori_ori_n706_));
  AOI210     o684(.A0(ori_ori_n706_), .A1(ori_ori_n694_), .B0(ori_ori_n107_), .Y(ori_ori_n707_));
  OR2        o685(.A(ori_ori_n707_), .B(i_5_), .Y(ori_ori_n708_));
  AOI210     o686(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n154_), .Y(ori_ori_n709_));
  NA2        o687(.A(ori_ori_n709_), .B(ori_ori_n680_), .Y(ori_ori_n710_));
  NO3        o688(.A(ori_ori_n631_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n711_));
  NA2        o689(.A(ori_ori_n344_), .B(ori_ori_n337_), .Y(ori_ori_n712_));
  NO3        o690(.A(ori_ori_n712_), .B(ori_ori_n711_), .C(ori_ori_n753_), .Y(ori_ori_n713_));
  NA3        o691(.A(ori_ori_n278_), .B(ori_ori_n151_), .C(ori_ori_n150_), .Y(ori_ori_n714_));
  NA3        o692(.A(i_5_), .B(ori_ori_n221_), .C(ori_ori_n185_), .Y(ori_ori_n715_));
  NA2        o693(.A(ori_ori_n715_), .B(ori_ori_n714_), .Y(ori_ori_n716_));
  NO3        o694(.A(ori_ori_n664_), .B(ori_ori_n178_), .C(ori_ori_n160_), .Y(ori_ori_n717_));
  NO2        o695(.A(ori_ori_n717_), .B(ori_ori_n716_), .Y(ori_ori_n718_));
  NA4        o696(.A(ori_ori_n718_), .B(ori_ori_n713_), .C(ori_ori_n710_), .D(ori_ori_n708_), .Y(ori_ori_n719_));
  NA2        o697(.A(ori_ori_n586_), .B(ori_ori_n155_), .Y(ori_ori_n720_));
  INV        o698(.A(ori_ori_n720_), .Y(ori_ori_n721_));
  NO4        o699(.A(ori_ori_n721_), .B(ori_ori_n719_), .C(ori_ori_n705_), .D(ori_ori_n700_), .Y(ori_ori_n722_));
  OAI210     o700(.A0(ori_ori_n608_), .A1(ori_ori_n604_), .B0(ori_ori_n37_), .Y(ori_ori_n723_));
  NA2        o701(.A(ori_ori_n723_), .B(ori_ori_n424_), .Y(ori_ori_n724_));
  NA2        o702(.A(ori_ori_n724_), .B(ori_ori_n170_), .Y(ori_ori_n725_));
  NA2        o703(.A(ori_ori_n158_), .B(ori_ori_n159_), .Y(ori_ori_n726_));
  AO210      o704(.A0(ori_ori_n496_), .A1(ori_ori_n33_), .B0(ori_ori_n726_), .Y(ori_ori_n727_));
  NAi31      o705(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n728_));
  AOI210     o706(.A0(ori_ori_n116_), .A1(ori_ori_n67_), .B0(ori_ori_n728_), .Y(ori_ori_n729_));
  NO2        o707(.A(ori_ori_n729_), .B(ori_ori_n455_), .Y(ori_ori_n730_));
  NA2        o708(.A(ori_ori_n730_), .B(ori_ori_n727_), .Y(ori_ori_n731_));
  NO2        o709(.A(ori_ori_n323_), .B(ori_ori_n208_), .Y(ori_ori_n732_));
  AOI210     o710(.A0(ori_ori_n731_), .A1(ori_ori_n48_), .B0(ori_ori_n732_), .Y(ori_ori_n733_));
  AOI210     o711(.A0(ori_ori_n733_), .A1(ori_ori_n725_), .B0(ori_ori_n70_), .Y(ori_ori_n734_));
  INV        o712(.A(ori_ori_n272_), .Y(ori_ori_n735_));
  NO2        o713(.A(ori_ori_n735_), .B(ori_ori_n551_), .Y(ori_ori_n736_));
  NA3        o714(.A(ori_ori_n555_), .B(ori_ori_n221_), .C(ori_ori_n77_), .Y(ori_ori_n737_));
  NO2        o715(.A(ori_ori_n737_), .B(i_11_), .Y(ori_ori_n738_));
  NO3        o716(.A(ori_ori_n58_), .B(ori_ori_n57_), .C(i_4_), .Y(ori_ori_n739_));
  OAI210     o717(.A0(ori_ori_n677_), .A1(ori_ori_n225_), .B0(ori_ori_n739_), .Y(ori_ori_n740_));
  NO2        o718(.A(ori_ori_n740_), .B(ori_ori_n524_), .Y(ori_ori_n741_));
  NO4        o719(.A(ori_ori_n687_), .B(ori_ori_n333_), .C(ori_ori_n197_), .D(ori_ori_n196_), .Y(ori_ori_n742_));
  NO2        o720(.A(ori_ori_n742_), .B(ori_ori_n384_), .Y(ori_ori_n743_));
  INV        o721(.A(ori_ori_n256_), .Y(ori_ori_n744_));
  AOI210     o722(.A0(ori_ori_n744_), .A1(ori_ori_n743_), .B0(ori_ori_n41_), .Y(ori_ori_n745_));
  NO3        o723(.A(ori_ori_n745_), .B(ori_ori_n741_), .C(ori_ori_n738_), .Y(ori_ori_n746_));
  INV        o724(.A(ori_ori_n746_), .Y(ori_ori_n747_));
  NO3        o725(.A(ori_ori_n747_), .B(ori_ori_n736_), .C(ori_ori_n734_), .Y(ori_ori_n748_));
  NA4        o726(.A(ori_ori_n748_), .B(ori_ori_n722_), .C(ori_ori_n693_), .D(ori_ori_n644_), .Y(ori4));
  INV        o727(.A(ori_ori_n500_), .Y(ori_ori_n752_));
  INV        o728(.A(ori_ori_n371_), .Y(ori_ori_n753_));
  INV        o729(.A(i_6_), .Y(ori_ori_n754_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NA2        m028(.A(i_0_), .B(i_2_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_7_), .B(i_9_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NA3        m031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n54_));
  NO2        m032(.A(i_1_), .B(i_6_), .Y(mai_mai_n55_));
  NA2        m033(.A(i_8_), .B(i_7_), .Y(mai_mai_n56_));
  OAI210     m034(.A0(mai_mai_n56_), .A1(mai_mai_n55_), .B0(mai_mai_n54_), .Y(mai_mai_n57_));
  NA2        m035(.A(mai_mai_n57_), .B(i_12_), .Y(mai_mai_n58_));
  NAi21      m036(.An(i_2_), .B(i_7_), .Y(mai_mai_n59_));
  INV        m037(.A(i_1_), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n61_));
  NA3        m039(.A(mai_mai_n61_), .B(mai_mai_n59_), .C(mai_mai_n31_), .Y(mai_mai_n62_));
  NA2        m040(.A(i_1_), .B(i_10_), .Y(mai_mai_n63_));
  NO2        m041(.A(mai_mai_n63_), .B(i_6_), .Y(mai_mai_n64_));
  NAi31      m042(.An(mai_mai_n64_), .B(mai_mai_n62_), .C(mai_mai_n58_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n66_));
  AOI210     m044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n67_));
  NA2        m045(.A(i_1_), .B(i_6_), .Y(mai_mai_n68_));
  NO2        m046(.A(mai_mai_n68_), .B(mai_mai_n25_), .Y(mai_mai_n69_));
  INV        m047(.A(i_0_), .Y(mai_mai_n70_));
  NAi21      m048(.An(i_5_), .B(i_10_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_5_), .B(i_9_), .Y(mai_mai_n72_));
  AOI210     m050(.A0(mai_mai_n72_), .A1(mai_mai_n71_), .B0(mai_mai_n70_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n69_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n74_), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n75_), .A1(mai_mai_n65_), .B0(i_0_), .Y(mai_mai_n76_));
  NA2        m054(.A(i_12_), .B(i_5_), .Y(mai_mai_n77_));
  NA2        m055(.A(i_2_), .B(i_8_), .Y(mai_mai_n78_));
  NO2        m056(.A(i_3_), .B(i_9_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_3_), .B(i_7_), .Y(mai_mai_n80_));
  NO3        m058(.A(mai_mai_n80_), .B(mai_mai_n79_), .C(mai_mai_n60_), .Y(mai_mai_n81_));
  INV        m059(.A(i_6_), .Y(mai_mai_n82_));
  NO2        m060(.A(i_2_), .B(i_7_), .Y(mai_mai_n83_));
  INV        m061(.A(mai_mai_n83_), .Y(mai_mai_n84_));
  NA2        m062(.A(mai_mai_n81_), .B(mai_mai_n84_), .Y(mai_mai_n85_));
  NAi21      m063(.An(i_6_), .B(i_10_), .Y(mai_mai_n86_));
  NA2        m064(.A(i_6_), .B(i_9_), .Y(mai_mai_n87_));
  AOI210     m065(.A0(mai_mai_n87_), .A1(mai_mai_n86_), .B0(mai_mai_n60_), .Y(mai_mai_n88_));
  NA2        m066(.A(i_2_), .B(i_6_), .Y(mai_mai_n89_));
  NO3        m067(.A(mai_mai_n89_), .B(mai_mai_n49_), .C(mai_mai_n25_), .Y(mai_mai_n90_));
  NO2        m068(.A(mai_mai_n90_), .B(mai_mai_n88_), .Y(mai_mai_n91_));
  AOI210     m069(.A0(mai_mai_n91_), .A1(mai_mai_n85_), .B0(mai_mai_n77_), .Y(mai_mai_n92_));
  AN3        m070(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n93_));
  NAi21      m071(.An(i_6_), .B(i_11_), .Y(mai_mai_n94_));
  NO2        m072(.A(i_5_), .B(i_8_), .Y(mai_mai_n95_));
  NOi21      m073(.An(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  AOI220     m074(.A0(mai_mai_n96_), .A1(mai_mai_n59_), .B0(mai_mai_n93_), .B1(mai_mai_n32_), .Y(mai_mai_n97_));
  INV        m075(.A(i_7_), .Y(mai_mai_n98_));
  NA2        m076(.A(mai_mai_n46_), .B(mai_mai_n98_), .Y(mai_mai_n99_));
  NO2        m077(.A(i_0_), .B(i_5_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n82_), .Y(mai_mai_n101_));
  NA2        m079(.A(i_12_), .B(i_3_), .Y(mai_mai_n102_));
  INV        m080(.A(mai_mai_n102_), .Y(mai_mai_n103_));
  NA3        m081(.A(mai_mai_n103_), .B(mai_mai_n101_), .C(mai_mai_n99_), .Y(mai_mai_n104_));
  NAi21      m082(.An(i_7_), .B(i_11_), .Y(mai_mai_n105_));
  AN2        m083(.A(i_2_), .B(i_10_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(i_7_), .Y(mai_mai_n107_));
  OR2        m085(.A(mai_mai_n77_), .B(mai_mai_n55_), .Y(mai_mai_n108_));
  NO2        m086(.A(i_8_), .B(mai_mai_n98_), .Y(mai_mai_n109_));
  NO3        m087(.A(mai_mai_n109_), .B(mai_mai_n108_), .C(mai_mai_n107_), .Y(mai_mai_n110_));
  NA2        m088(.A(i_12_), .B(i_7_), .Y(mai_mai_n111_));
  NA2        m089(.A(i_11_), .B(i_12_), .Y(mai_mai_n112_));
  INV        m090(.A(mai_mai_n112_), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n113_), .B(mai_mai_n110_), .Y(mai_mai_n114_));
  NA3        m092(.A(mai_mai_n114_), .B(mai_mai_n104_), .C(mai_mai_n97_), .Y(mai_mai_n115_));
  NOi21      m093(.An(i_1_), .B(i_5_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n116_), .B(i_11_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n98_), .B(mai_mai_n37_), .Y(mai_mai_n118_));
  NA2        m096(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n120_), .B(mai_mai_n46_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n87_), .B(mai_mai_n86_), .Y(mai_mai_n122_));
  NAi21      m100(.An(i_3_), .B(i_8_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n123_), .B(mai_mai_n59_), .Y(mai_mai_n124_));
  NOi31      m102(.An(mai_mai_n124_), .B(mai_mai_n122_), .C(mai_mai_n121_), .Y(mai_mai_n125_));
  NO2        m103(.A(i_1_), .B(mai_mai_n82_), .Y(mai_mai_n126_));
  NO2        m104(.A(i_6_), .B(i_5_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(i_3_), .Y(mai_mai_n128_));
  OAI220     m106(.A0(mai_mai_n128_), .A1(mai_mai_n105_), .B0(mai_mai_n125_), .B1(mai_mai_n117_), .Y(mai_mai_n129_));
  NO3        m107(.A(mai_mai_n129_), .B(mai_mai_n115_), .C(mai_mai_n92_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(mai_mai_n76_), .Y(mai2));
  NO2        m109(.A(mai_mai_n60_), .B(mai_mai_n37_), .Y(mai_mai_n132_));
  NA2        m110(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n134_));
  NA4        m112(.A(mai_mai_n134_), .B(mai_mai_n74_), .C(mai_mai_n66_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m113(.A(i_8_), .B(i_7_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n136_), .B(i_6_), .Y(mai_mai_n137_));
  NO2        m115(.A(i_12_), .B(i_13_), .Y(mai_mai_n138_));
  NAi21      m116(.An(i_5_), .B(i_11_), .Y(mai_mai_n139_));
  NOi21      m117(.An(mai_mai_n138_), .B(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m118(.A(i_0_), .B(i_1_), .Y(mai_mai_n141_));
  NA2        m119(.A(i_2_), .B(i_3_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n142_), .B(i_4_), .Y(mai_mai_n143_));
  NA3        m121(.A(mai_mai_n143_), .B(mai_mai_n141_), .C(mai_mai_n140_), .Y(mai_mai_n144_));
  AN2        m122(.A(mai_mai_n138_), .B(mai_mai_n79_), .Y(mai_mai_n145_));
  NO2        m123(.A(mai_mai_n145_), .B(mai_mai_n27_), .Y(mai_mai_n146_));
  NA2        m124(.A(i_1_), .B(i_5_), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n70_), .B(mai_mai_n46_), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n36_), .Y(mai_mai_n149_));
  NO3        m127(.A(mai_mai_n149_), .B(mai_mai_n147_), .C(mai_mai_n146_), .Y(mai_mai_n150_));
  OR2        m128(.A(i_0_), .B(i_1_), .Y(mai_mai_n151_));
  NO3        m129(.A(mai_mai_n151_), .B(mai_mai_n77_), .C(i_13_), .Y(mai_mai_n152_));
  NAi32      m130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n153_));
  NAi21      m131(.An(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NOi21      m132(.An(i_4_), .B(i_10_), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n155_), .B(mai_mai_n40_), .Y(mai_mai_n156_));
  NO2        m134(.A(i_3_), .B(i_5_), .Y(mai_mai_n157_));
  NO3        m135(.A(mai_mai_n70_), .B(i_2_), .C(i_1_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  OAI210     m137(.A0(mai_mai_n159_), .A1(mai_mai_n156_), .B0(mai_mai_n154_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n160_), .B(mai_mai_n150_), .Y(mai_mai_n161_));
  AOI210     m139(.A0(mai_mai_n161_), .A1(mai_mai_n144_), .B0(mai_mai_n137_), .Y(mai_mai_n162_));
  NA2        m140(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n163_));
  NOi21      m141(.An(i_4_), .B(i_9_), .Y(mai_mai_n164_));
  NOi21      m142(.An(i_11_), .B(i_13_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  OR2        m144(.A(mai_mai_n166_), .B(mai_mai_n163_), .Y(mai_mai_n167_));
  NO2        m145(.A(i_4_), .B(i_5_), .Y(mai_mai_n168_));
  NAi21      m146(.An(i_12_), .B(i_11_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n169_), .B(i_13_), .Y(mai_mai_n170_));
  NA3        m148(.A(mai_mai_n170_), .B(mai_mai_n168_), .C(mai_mai_n79_), .Y(mai_mai_n171_));
  AOI210     m149(.A0(mai_mai_n171_), .A1(mai_mai_n167_), .B0(mai_mai_n1001_), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n70_), .B(mai_mai_n60_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n173_), .B(mai_mai_n46_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n175_));
  NAi31      m153(.An(mai_mai_n175_), .B(mai_mai_n145_), .C(i_11_), .Y(mai_mai_n176_));
  NA2        m154(.A(i_3_), .B(i_5_), .Y(mai_mai_n177_));
  AOI210     m155(.A0(mai_mai_n166_), .A1(mai_mai_n176_), .B0(mai_mai_n174_), .Y(mai_mai_n178_));
  NO2        m156(.A(mai_mai_n70_), .B(i_5_), .Y(mai_mai_n179_));
  NO2        m157(.A(i_13_), .B(i_10_), .Y(mai_mai_n180_));
  NA3        m158(.A(mai_mai_n180_), .B(mai_mai_n179_), .C(mai_mai_n44_), .Y(mai_mai_n181_));
  NO2        m159(.A(i_2_), .B(i_1_), .Y(mai_mai_n182_));
  NA2        m160(.A(mai_mai_n182_), .B(i_3_), .Y(mai_mai_n183_));
  NAi21      m161(.An(i_4_), .B(i_12_), .Y(mai_mai_n184_));
  NO4        m162(.A(mai_mai_n184_), .B(mai_mai_n183_), .C(mai_mai_n181_), .D(mai_mai_n25_), .Y(mai_mai_n185_));
  NO3        m163(.A(mai_mai_n185_), .B(mai_mai_n178_), .C(mai_mai_n172_), .Y(mai_mai_n186_));
  INV        m164(.A(i_8_), .Y(mai_mai_n187_));
  NO2        m165(.A(mai_mai_n187_), .B(i_7_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n188_), .B(i_6_), .Y(mai_mai_n189_));
  NO3        m167(.A(i_3_), .B(mai_mai_n82_), .C(mai_mai_n48_), .Y(mai_mai_n190_));
  NA2        m168(.A(mai_mai_n190_), .B(mai_mai_n109_), .Y(mai_mai_n191_));
  NO3        m169(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n192_));
  NA3        m170(.A(mai_mai_n192_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n193_));
  NO3        m171(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n194_));
  OAI210     m172(.A0(mai_mai_n93_), .A1(i_12_), .B0(mai_mai_n194_), .Y(mai_mai_n195_));
  AOI210     m173(.A0(mai_mai_n195_), .A1(mai_mai_n193_), .B0(mai_mai_n191_), .Y(mai_mai_n196_));
  NO2        m174(.A(i_3_), .B(i_8_), .Y(mai_mai_n197_));
  NO3        m175(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n198_));
  NO2        m176(.A(i_13_), .B(i_9_), .Y(mai_mai_n199_));
  NA3        m177(.A(mai_mai_n199_), .B(i_6_), .C(mai_mai_n187_), .Y(mai_mai_n200_));
  NAi21      m178(.An(i_12_), .B(i_3_), .Y(mai_mai_n201_));
  NO2        m179(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n202_));
  NO3        m180(.A(i_0_), .B(i_2_), .C(mai_mai_n60_), .Y(mai_mai_n203_));
  NA3        m181(.A(mai_mai_n203_), .B(mai_mai_n202_), .C(i_10_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n204_), .B(mai_mai_n200_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n205_), .B(mai_mai_n196_), .Y(mai_mai_n206_));
  OAI220     m184(.A0(mai_mai_n206_), .A1(i_4_), .B0(mai_mai_n189_), .B1(mai_mai_n186_), .Y(mai_mai_n207_));
  NAi21      m185(.An(i_12_), .B(i_7_), .Y(mai_mai_n208_));
  NA3        m186(.A(i_13_), .B(mai_mai_n187_), .C(i_10_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n210_));
  NA2        m188(.A(i_0_), .B(i_5_), .Y(mai_mai_n211_));
  NA2        m189(.A(mai_mai_n211_), .B(mai_mai_n101_), .Y(mai_mai_n212_));
  OAI220     m190(.A0(mai_mai_n212_), .A1(mai_mai_n183_), .B0(mai_mai_n174_), .B1(mai_mai_n128_), .Y(mai_mai_n213_));
  NAi31      m191(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n70_), .B(mai_mai_n26_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n46_), .B(mai_mai_n60_), .Y(mai_mai_n217_));
  NA3        m195(.A(mai_mai_n217_), .B(mai_mai_n216_), .C(mai_mai_n215_), .Y(mai_mai_n218_));
  INV        m196(.A(i_13_), .Y(mai_mai_n219_));
  NO2        m197(.A(i_12_), .B(mai_mai_n219_), .Y(mai_mai_n220_));
  NA3        m198(.A(mai_mai_n220_), .B(mai_mai_n192_), .C(mai_mai_n190_), .Y(mai_mai_n221_));
  OAI210     m199(.A0(mai_mai_n218_), .A1(mai_mai_n214_), .B0(mai_mai_n221_), .Y(mai_mai_n222_));
  AOI220     m200(.A0(mai_mai_n222_), .A1(mai_mai_n136_), .B0(mai_mai_n213_), .B1(mai_mai_n210_), .Y(mai_mai_n223_));
  NO2        m201(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n177_), .B(i_4_), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n226_));
  OR2        m204(.A(i_8_), .B(i_7_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n227_), .B(mai_mai_n82_), .Y(mai_mai_n228_));
  NO2        m206(.A(mai_mai_n51_), .B(i_1_), .Y(mai_mai_n229_));
  NA2        m207(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n230_));
  INV        m208(.A(i_12_), .Y(mai_mai_n231_));
  NO2        m209(.A(mai_mai_n44_), .B(mai_mai_n231_), .Y(mai_mai_n232_));
  NO3        m210(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n233_));
  NA2        m211(.A(i_2_), .B(i_1_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n230_), .B(mai_mai_n226_), .Y(mai_mai_n235_));
  NO3        m213(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n236_));
  NAi21      m214(.An(i_4_), .B(i_3_), .Y(mai_mai_n237_));
  NO2        m215(.A(i_0_), .B(i_6_), .Y(mai_mai_n238_));
  NOi41      m216(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n239_));
  NA2        m217(.A(mai_mai_n239_), .B(mai_mai_n238_), .Y(mai_mai_n240_));
  NO2        m218(.A(mai_mai_n234_), .B(mai_mai_n177_), .Y(mai_mai_n241_));
  NAi21      m219(.An(mai_mai_n240_), .B(mai_mai_n241_), .Y(mai_mai_n242_));
  INV        m220(.A(mai_mai_n242_), .Y(mai_mai_n243_));
  AOI210     m221(.A0(mai_mai_n243_), .A1(mai_mai_n40_), .B0(mai_mai_n235_), .Y(mai_mai_n244_));
  NO2        m222(.A(i_11_), .B(mai_mai_n219_), .Y(mai_mai_n245_));
  NOi21      m223(.An(i_1_), .B(i_6_), .Y(mai_mai_n246_));
  NAi21      m224(.An(i_3_), .B(i_7_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n231_), .B(i_9_), .Y(mai_mai_n248_));
  OR4        m226(.A(mai_mai_n248_), .B(mai_mai_n247_), .C(mai_mai_n246_), .D(mai_mai_n179_), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n48_), .B(mai_mai_n25_), .Y(mai_mai_n250_));
  NO2        m228(.A(i_12_), .B(i_3_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n70_), .B(i_5_), .Y(mai_mai_n252_));
  NA2        m230(.A(i_3_), .B(i_9_), .Y(mai_mai_n253_));
  NAi21      m231(.An(i_7_), .B(i_10_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n254_), .B(mai_mai_n253_), .Y(mai_mai_n255_));
  NA3        m233(.A(mai_mai_n255_), .B(mai_mai_n252_), .C(mai_mai_n61_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n256_), .B(mai_mai_n249_), .Y(mai_mai_n257_));
  NA3        m235(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n258_));
  INV        m236(.A(mai_mai_n137_), .Y(mai_mai_n259_));
  NA2        m237(.A(mai_mai_n231_), .B(i_13_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n260_), .B(mai_mai_n72_), .Y(mai_mai_n261_));
  AOI220     m239(.A0(mai_mai_n261_), .A1(mai_mai_n259_), .B0(mai_mai_n257_), .B1(mai_mai_n245_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n227_), .B(mai_mai_n37_), .Y(mai_mai_n263_));
  NA2        m241(.A(i_12_), .B(i_6_), .Y(mai_mai_n264_));
  OR2        m242(.A(i_13_), .B(i_9_), .Y(mai_mai_n265_));
  NO3        m243(.A(mai_mai_n265_), .B(mai_mai_n264_), .C(mai_mai_n48_), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n237_), .B(i_2_), .Y(mai_mai_n267_));
  NA2        m245(.A(mai_mai_n245_), .B(i_9_), .Y(mai_mai_n268_));
  NA2        m246(.A(mai_mai_n148_), .B(mai_mai_n60_), .Y(mai_mai_n269_));
  NO3        m247(.A(i_11_), .B(mai_mai_n219_), .C(mai_mai_n25_), .Y(mai_mai_n270_));
  NO2        m248(.A(mai_mai_n247_), .B(i_8_), .Y(mai_mai_n271_));
  NO2        m249(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n272_));
  NA3        m250(.A(mai_mai_n272_), .B(mai_mai_n271_), .C(mai_mai_n270_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n26_), .B(mai_mai_n82_), .Y(mai_mai_n274_));
  NA3        m252(.A(mai_mai_n274_), .B(mai_mai_n263_), .C(mai_mai_n220_), .Y(mai_mai_n275_));
  AOI210     m253(.A0(mai_mai_n275_), .A1(mai_mai_n273_), .B0(mai_mai_n269_), .Y(mai_mai_n276_));
  INV        m254(.A(mai_mai_n276_), .Y(mai_mai_n277_));
  NA4        m255(.A(mai_mai_n277_), .B(mai_mai_n262_), .C(mai_mai_n244_), .D(mai_mai_n223_), .Y(mai_mai_n278_));
  NO3        m256(.A(i_12_), .B(mai_mai_n219_), .C(mai_mai_n37_), .Y(mai_mai_n279_));
  INV        m257(.A(mai_mai_n279_), .Y(mai_mai_n280_));
  NA2        m258(.A(i_8_), .B(mai_mai_n98_), .Y(mai_mai_n281_));
  NOi21      m259(.An(mai_mai_n157_), .B(mai_mai_n82_), .Y(mai_mai_n282_));
  NO3        m260(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n283_));
  AOI220     m261(.A0(mai_mai_n283_), .A1(mai_mai_n190_), .B0(mai_mai_n282_), .B1(mai_mai_n229_), .Y(mai_mai_n284_));
  NO2        m262(.A(mai_mai_n284_), .B(mai_mai_n281_), .Y(mai_mai_n285_));
  NO2        m263(.A(mai_mai_n234_), .B(i_0_), .Y(mai_mai_n286_));
  AOI220     m264(.A0(mai_mai_n286_), .A1(mai_mai_n188_), .B0(i_1_), .B1(mai_mai_n136_), .Y(mai_mai_n287_));
  NA2        m265(.A(mai_mai_n272_), .B(mai_mai_n26_), .Y(mai_mai_n288_));
  NO2        m266(.A(mai_mai_n288_), .B(mai_mai_n287_), .Y(mai_mai_n289_));
  NA2        m267(.A(i_0_), .B(i_1_), .Y(mai_mai_n290_));
  NO2        m268(.A(mai_mai_n290_), .B(i_2_), .Y(mai_mai_n291_));
  NO2        m269(.A(mai_mai_n56_), .B(i_6_), .Y(mai_mai_n292_));
  NA3        m270(.A(mai_mai_n292_), .B(mai_mai_n291_), .C(mai_mai_n157_), .Y(mai_mai_n293_));
  OAI210     m271(.A0(mai_mai_n159_), .A1(mai_mai_n137_), .B0(mai_mai_n293_), .Y(mai_mai_n294_));
  NO3        m272(.A(mai_mai_n294_), .B(mai_mai_n289_), .C(mai_mai_n285_), .Y(mai_mai_n295_));
  NO2        m273(.A(i_3_), .B(i_10_), .Y(mai_mai_n296_));
  NA3        m274(.A(mai_mai_n296_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n297_));
  NO2        m275(.A(i_2_), .B(mai_mai_n98_), .Y(mai_mai_n298_));
  NA2        m276(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n299_));
  NO2        m277(.A(mai_mai_n299_), .B(i_8_), .Y(mai_mai_n300_));
  NA2        m278(.A(mai_mai_n300_), .B(mai_mai_n298_), .Y(mai_mai_n301_));
  AN2        m279(.A(i_3_), .B(i_10_), .Y(mai_mai_n302_));
  NA4        m280(.A(mai_mai_n302_), .B(mai_mai_n192_), .C(mai_mai_n170_), .D(mai_mai_n168_), .Y(mai_mai_n303_));
  NO2        m281(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n304_));
  NO2        m282(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n305_));
  OR2        m283(.A(mai_mai_n301_), .B(mai_mai_n297_), .Y(mai_mai_n306_));
  OAI220     m284(.A0(mai_mai_n306_), .A1(i_6_), .B0(mai_mai_n295_), .B1(mai_mai_n280_), .Y(mai_mai_n307_));
  NO4        m285(.A(mai_mai_n307_), .B(mai_mai_n278_), .C(mai_mai_n207_), .D(mai_mai_n162_), .Y(mai_mai_n308_));
  NO3        m286(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n309_));
  NO2        m287(.A(mai_mai_n56_), .B(mai_mai_n82_), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n286_), .B(mai_mai_n310_), .Y(mai_mai_n311_));
  NO3        m289(.A(i_6_), .B(mai_mai_n187_), .C(i_7_), .Y(mai_mai_n312_));
  NA2        m290(.A(mai_mai_n312_), .B(mai_mai_n192_), .Y(mai_mai_n313_));
  AOI210     m291(.A0(mai_mai_n313_), .A1(mai_mai_n311_), .B0(mai_mai_n163_), .Y(mai_mai_n314_));
  NO2        m292(.A(i_2_), .B(i_3_), .Y(mai_mai_n315_));
  OR2        m293(.A(i_0_), .B(i_5_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n211_), .B(mai_mai_n316_), .Y(mai_mai_n317_));
  NA4        m295(.A(mai_mai_n317_), .B(mai_mai_n228_), .C(mai_mai_n315_), .D(i_1_), .Y(mai_mai_n318_));
  NA3        m296(.A(mai_mai_n286_), .B(mai_mai_n282_), .C(mai_mai_n109_), .Y(mai_mai_n319_));
  NAi21      m297(.An(i_8_), .B(i_7_), .Y(mai_mai_n320_));
  NO2        m298(.A(mai_mai_n320_), .B(i_6_), .Y(mai_mai_n321_));
  NO2        m299(.A(mai_mai_n151_), .B(mai_mai_n46_), .Y(mai_mai_n322_));
  NA3        m300(.A(mai_mai_n322_), .B(mai_mai_n321_), .C(mai_mai_n157_), .Y(mai_mai_n323_));
  NA3        m301(.A(mai_mai_n323_), .B(mai_mai_n319_), .C(mai_mai_n318_), .Y(mai_mai_n324_));
  OAI210     m302(.A0(mai_mai_n324_), .A1(mai_mai_n314_), .B0(i_4_), .Y(mai_mai_n325_));
  NO2        m303(.A(i_12_), .B(i_10_), .Y(mai_mai_n326_));
  NOi21      m304(.An(i_5_), .B(i_0_), .Y(mai_mai_n327_));
  NA4        m305(.A(mai_mai_n80_), .B(mai_mai_n36_), .C(mai_mai_n82_), .D(i_8_), .Y(mai_mai_n328_));
  NO2        m306(.A(i_6_), .B(i_8_), .Y(mai_mai_n329_));
  NOi21      m307(.An(i_0_), .B(i_2_), .Y(mai_mai_n330_));
  AN2        m308(.A(mai_mai_n330_), .B(mai_mai_n329_), .Y(mai_mai_n331_));
  NO2        m309(.A(i_1_), .B(i_7_), .Y(mai_mai_n332_));
  AO220      m310(.A0(mai_mai_n332_), .A1(mai_mai_n331_), .B0(mai_mai_n321_), .B1(mai_mai_n229_), .Y(mai_mai_n333_));
  NA3        m311(.A(mai_mai_n333_), .B(i_4_), .C(i_5_), .Y(mai_mai_n334_));
  NA2        m312(.A(mai_mai_n334_), .B(mai_mai_n325_), .Y(mai_mai_n335_));
  NO3        m313(.A(mai_mai_n227_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n336_));
  NO3        m314(.A(mai_mai_n320_), .B(i_2_), .C(i_1_), .Y(mai_mai_n337_));
  OAI210     m315(.A0(mai_mai_n337_), .A1(mai_mai_n336_), .B0(i_6_), .Y(mai_mai_n338_));
  NA3        m316(.A(mai_mai_n246_), .B(mai_mai_n298_), .C(mai_mai_n187_), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(mai_mai_n317_), .Y(mai_mai_n340_));
  NOi21      m318(.An(mai_mai_n147_), .B(mai_mai_n101_), .Y(mai_mai_n341_));
  NO2        m319(.A(mai_mai_n341_), .B(mai_mai_n119_), .Y(mai_mai_n342_));
  OAI210     m320(.A0(mai_mai_n342_), .A1(mai_mai_n340_), .B0(i_3_), .Y(mai_mai_n343_));
  INV        m321(.A(mai_mai_n80_), .Y(mai_mai_n344_));
  NO2        m322(.A(mai_mai_n290_), .B(mai_mai_n78_), .Y(mai_mai_n345_));
  NA2        m323(.A(mai_mai_n345_), .B(mai_mai_n127_), .Y(mai_mai_n346_));
  NO2        m324(.A(mai_mai_n89_), .B(mai_mai_n187_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n347_), .B(mai_mai_n60_), .Y(mai_mai_n348_));
  AOI210     m326(.A0(mai_mai_n348_), .A1(mai_mai_n346_), .B0(mai_mai_n344_), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n187_), .B(i_9_), .Y(mai_mai_n350_));
  NA2        m328(.A(mai_mai_n350_), .B(i_1_), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n351_), .B(mai_mai_n46_), .Y(mai_mai_n352_));
  NO3        m330(.A(mai_mai_n352_), .B(mai_mai_n349_), .C(mai_mai_n289_), .Y(mai_mai_n353_));
  AOI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n343_), .B0(mai_mai_n156_), .Y(mai_mai_n354_));
  AOI210     m332(.A0(mai_mai_n335_), .A1(mai_mai_n309_), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  NOi32      m333(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n356_));
  INV        m334(.A(mai_mai_n356_), .Y(mai_mai_n357_));
  NAi21      m335(.An(i_0_), .B(i_6_), .Y(mai_mai_n358_));
  NAi21      m336(.An(i_1_), .B(i_5_), .Y(mai_mai_n359_));
  NA2        m337(.A(mai_mai_n359_), .B(mai_mai_n358_), .Y(mai_mai_n360_));
  NA2        m338(.A(mai_mai_n360_), .B(mai_mai_n25_), .Y(mai_mai_n361_));
  OAI210     m339(.A0(mai_mai_n361_), .A1(mai_mai_n153_), .B0(mai_mai_n240_), .Y(mai_mai_n362_));
  NAi41      m340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n363_));
  NO2        m341(.A(mai_mai_n153_), .B(mai_mai_n151_), .Y(mai_mai_n364_));
  NOi32      m342(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n365_));
  NO2        m343(.A(i_1_), .B(mai_mai_n98_), .Y(mai_mai_n366_));
  NAi21      m344(.An(i_3_), .B(i_4_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n367_), .B(i_9_), .Y(mai_mai_n368_));
  AN2        m346(.A(i_6_), .B(i_7_), .Y(mai_mai_n369_));
  OAI210     m347(.A0(mai_mai_n369_), .A1(mai_mai_n366_), .B0(mai_mai_n368_), .Y(mai_mai_n370_));
  NA2        m348(.A(i_2_), .B(i_7_), .Y(mai_mai_n371_));
  NO2        m349(.A(mai_mai_n367_), .B(i_10_), .Y(mai_mai_n372_));
  NA3        m350(.A(mai_mai_n372_), .B(mai_mai_n371_), .C(mai_mai_n238_), .Y(mai_mai_n373_));
  AOI210     m351(.A0(mai_mai_n373_), .A1(mai_mai_n370_), .B0(mai_mai_n179_), .Y(mai_mai_n374_));
  AOI210     m352(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n375_));
  OAI210     m353(.A0(mai_mai_n375_), .A1(mai_mai_n182_), .B0(mai_mai_n372_), .Y(mai_mai_n376_));
  NO2        m354(.A(mai_mai_n376_), .B(i_5_), .Y(mai_mai_n377_));
  NO4        m355(.A(mai_mai_n377_), .B(mai_mai_n374_), .C(mai_mai_n364_), .D(mai_mai_n362_), .Y(mai_mai_n378_));
  NO2        m356(.A(mai_mai_n378_), .B(mai_mai_n357_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n56_), .B(mai_mai_n25_), .Y(mai_mai_n380_));
  AN2        m358(.A(i_12_), .B(i_5_), .Y(mai_mai_n381_));
  NO2        m359(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n382_));
  NA2        m360(.A(mai_mai_n382_), .B(mai_mai_n381_), .Y(mai_mai_n383_));
  NO2        m361(.A(i_11_), .B(i_6_), .Y(mai_mai_n384_));
  NA3        m362(.A(mai_mai_n384_), .B(mai_mai_n322_), .C(mai_mai_n219_), .Y(mai_mai_n385_));
  NO2        m363(.A(mai_mai_n385_), .B(mai_mai_n383_), .Y(mai_mai_n386_));
  NO2        m364(.A(mai_mai_n237_), .B(i_5_), .Y(mai_mai_n387_));
  NO2        m365(.A(i_5_), .B(i_10_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n138_), .B(mai_mai_n45_), .Y(mai_mai_n389_));
  NO2        m367(.A(mai_mai_n389_), .B(mai_mai_n237_), .Y(mai_mai_n390_));
  OAI210     m368(.A0(mai_mai_n390_), .A1(mai_mai_n386_), .B0(mai_mai_n380_), .Y(mai_mai_n391_));
  NO2        m369(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n392_));
  NA2        m370(.A(mai_mai_n386_), .B(mai_mai_n392_), .Y(mai_mai_n393_));
  NO3        m371(.A(mai_mai_n82_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n394_));
  NO2        m372(.A(i_11_), .B(i_12_), .Y(mai_mai_n395_));
  NA2        m373(.A(mai_mai_n388_), .B(mai_mai_n231_), .Y(mai_mai_n396_));
  NA3        m374(.A(mai_mai_n109_), .B(i_4_), .C(i_11_), .Y(mai_mai_n397_));
  NO2        m375(.A(mai_mai_n397_), .B(mai_mai_n214_), .Y(mai_mai_n398_));
  NAi21      m376(.An(i_13_), .B(i_0_), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n399_), .B(mai_mai_n234_), .Y(mai_mai_n400_));
  NA2        m378(.A(mai_mai_n398_), .B(mai_mai_n400_), .Y(mai_mai_n401_));
  NA3        m379(.A(mai_mai_n401_), .B(mai_mai_n393_), .C(mai_mai_n391_), .Y(mai_mai_n402_));
  NA2        m380(.A(mai_mai_n44_), .B(mai_mai_n219_), .Y(mai_mai_n403_));
  NO3        m381(.A(i_1_), .B(i_12_), .C(mai_mai_n82_), .Y(mai_mai_n404_));
  NO2        m382(.A(i_0_), .B(i_11_), .Y(mai_mai_n405_));
  INV        m383(.A(i_5_), .Y(mai_mai_n406_));
  AN2        m384(.A(i_1_), .B(i_6_), .Y(mai_mai_n407_));
  NOi21      m385(.An(i_2_), .B(i_12_), .Y(mai_mai_n408_));
  NA2        m386(.A(mai_mai_n408_), .B(mai_mai_n407_), .Y(mai_mai_n409_));
  NO2        m387(.A(mai_mai_n409_), .B(mai_mai_n406_), .Y(mai_mai_n410_));
  NA2        m388(.A(mai_mai_n136_), .B(i_9_), .Y(mai_mai_n411_));
  NO2        m389(.A(mai_mai_n411_), .B(i_4_), .Y(mai_mai_n412_));
  NA2        m390(.A(mai_mai_n410_), .B(mai_mai_n412_), .Y(mai_mai_n413_));
  NAi21      m391(.An(i_9_), .B(i_4_), .Y(mai_mai_n414_));
  OR2        m392(.A(i_13_), .B(i_10_), .Y(mai_mai_n415_));
  NO3        m393(.A(mai_mai_n415_), .B(mai_mai_n112_), .C(mai_mai_n414_), .Y(mai_mai_n416_));
  OR2        m394(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n417_));
  NO2        m395(.A(mai_mai_n98_), .B(mai_mai_n25_), .Y(mai_mai_n418_));
  NA2        m396(.A(mai_mai_n279_), .B(mai_mai_n418_), .Y(mai_mai_n419_));
  NA2        m397(.A(mai_mai_n272_), .B(mai_mai_n203_), .Y(mai_mai_n420_));
  OAI220     m398(.A0(mai_mai_n420_), .A1(mai_mai_n417_), .B0(mai_mai_n419_), .B1(mai_mai_n341_), .Y(mai_mai_n421_));
  INV        m399(.A(mai_mai_n421_), .Y(mai_mai_n422_));
  AOI210     m400(.A0(mai_mai_n422_), .A1(mai_mai_n413_), .B0(mai_mai_n26_), .Y(mai_mai_n423_));
  NA2        m401(.A(mai_mai_n319_), .B(mai_mai_n318_), .Y(mai_mai_n424_));
  AOI220     m402(.A0(mai_mai_n292_), .A1(mai_mai_n283_), .B0(mai_mai_n286_), .B1(mai_mai_n310_), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n425_), .B(mai_mai_n163_), .Y(mai_mai_n426_));
  NO2        m404(.A(mai_mai_n177_), .B(mai_mai_n82_), .Y(mai_mai_n427_));
  AOI220     m405(.A0(mai_mai_n427_), .A1(mai_mai_n291_), .B0(mai_mai_n274_), .B1(mai_mai_n203_), .Y(mai_mai_n428_));
  NO2        m406(.A(mai_mai_n428_), .B(mai_mai_n281_), .Y(mai_mai_n429_));
  NO3        m407(.A(mai_mai_n429_), .B(mai_mai_n426_), .C(mai_mai_n424_), .Y(mai_mai_n430_));
  NA2        m408(.A(mai_mai_n190_), .B(mai_mai_n93_), .Y(mai_mai_n431_));
  NA3        m409(.A(mai_mai_n322_), .B(mai_mai_n157_), .C(mai_mai_n82_), .Y(mai_mai_n432_));
  AOI210     m410(.A0(mai_mai_n432_), .A1(mai_mai_n431_), .B0(mai_mai_n320_), .Y(mai_mai_n433_));
  NA2        m411(.A(mai_mai_n187_), .B(i_10_), .Y(mai_mai_n434_));
  NA3        m412(.A(mai_mai_n252_), .B(mai_mai_n61_), .C(i_2_), .Y(mai_mai_n435_));
  NA2        m413(.A(mai_mai_n292_), .B(mai_mai_n229_), .Y(mai_mai_n436_));
  OAI220     m414(.A0(mai_mai_n436_), .A1(mai_mai_n177_), .B0(mai_mai_n435_), .B1(mai_mai_n434_), .Y(mai_mai_n437_));
  NO2        m415(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n438_));
  NA3        m416(.A(mai_mai_n332_), .B(mai_mai_n331_), .C(mai_mai_n438_), .Y(mai_mai_n439_));
  NA2        m417(.A(mai_mai_n312_), .B(mai_mai_n317_), .Y(mai_mai_n440_));
  OAI210     m418(.A0(mai_mai_n440_), .A1(mai_mai_n183_), .B0(mai_mai_n439_), .Y(mai_mai_n441_));
  NO3        m419(.A(mai_mai_n441_), .B(mai_mai_n437_), .C(mai_mai_n433_), .Y(mai_mai_n442_));
  AOI210     m420(.A0(mai_mai_n442_), .A1(mai_mai_n430_), .B0(mai_mai_n268_), .Y(mai_mai_n443_));
  NO4        m421(.A(mai_mai_n443_), .B(mai_mai_n423_), .C(mai_mai_n402_), .D(mai_mai_n379_), .Y(mai_mai_n444_));
  NO2        m422(.A(mai_mai_n60_), .B(i_4_), .Y(mai_mai_n445_));
  NO2        m423(.A(mai_mai_n70_), .B(i_13_), .Y(mai_mai_n446_));
  NO2        m424(.A(i_10_), .B(i_9_), .Y(mai_mai_n447_));
  NAi21      m425(.An(i_12_), .B(i_8_), .Y(mai_mai_n448_));
  NO2        m426(.A(mai_mai_n448_), .B(i_3_), .Y(mai_mai_n449_));
  INV        m427(.A(i_0_), .Y(mai_mai_n450_));
  NO3        m428(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n451_));
  NA2        m429(.A(mai_mai_n264_), .B(mai_mai_n94_), .Y(mai_mai_n452_));
  NA2        m430(.A(mai_mai_n452_), .B(mai_mai_n451_), .Y(mai_mai_n453_));
  NA2        m431(.A(i_8_), .B(i_9_), .Y(mai_mai_n454_));
  NO3        m432(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n455_));
  NA3        m433(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n456_));
  OR2        m434(.A(mai_mai_n290_), .B(mai_mai_n200_), .Y(mai_mai_n457_));
  BUFFER     m435(.A(mai_mai_n293_), .Y(mai_mai_n458_));
  OA220      m436(.A0(mai_mai_n458_), .A1(mai_mai_n156_), .B0(mai_mai_n457_), .B1(mai_mai_n226_), .Y(mai_mai_n459_));
  NA2        m437(.A(mai_mai_n93_), .B(i_13_), .Y(mai_mai_n460_));
  NA2        m438(.A(mai_mai_n427_), .B(mai_mai_n380_), .Y(mai_mai_n461_));
  NO2        m439(.A(i_2_), .B(i_13_), .Y(mai_mai_n462_));
  NO2        m440(.A(mai_mai_n461_), .B(mai_mai_n460_), .Y(mai_mai_n463_));
  NO3        m441(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n464_));
  NO2        m442(.A(i_6_), .B(i_7_), .Y(mai_mai_n465_));
  NA2        m443(.A(mai_mai_n465_), .B(mai_mai_n464_), .Y(mai_mai_n466_));
  NO2        m444(.A(i_11_), .B(i_1_), .Y(mai_mai_n467_));
  NO2        m445(.A(mai_mai_n70_), .B(i_3_), .Y(mai_mai_n468_));
  NOi21      m446(.An(i_2_), .B(i_7_), .Y(mai_mai_n469_));
  NAi31      m447(.An(i_11_), .B(mai_mai_n469_), .C(mai_mai_n468_), .Y(mai_mai_n470_));
  INV        m448(.A(mai_mai_n415_), .Y(mai_mai_n471_));
  NA3        m449(.A(mai_mai_n471_), .B(mai_mai_n445_), .C(mai_mai_n72_), .Y(mai_mai_n472_));
  NO2        m450(.A(mai_mai_n472_), .B(mai_mai_n470_), .Y(mai_mai_n473_));
  NO2        m451(.A(i_6_), .B(i_10_), .Y(mai_mai_n474_));
  NA4        m452(.A(mai_mai_n474_), .B(mai_mai_n309_), .C(i_8_), .D(mai_mai_n231_), .Y(mai_mai_n475_));
  NO2        m453(.A(mai_mai_n475_), .B(mai_mai_n149_), .Y(mai_mai_n476_));
  NA2        m454(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n477_));
  NO2        m455(.A(mai_mai_n151_), .B(i_3_), .Y(mai_mai_n478_));
  NAi31      m456(.An(mai_mai_n477_), .B(mai_mai_n478_), .C(mai_mai_n220_), .Y(mai_mai_n479_));
  NA3        m457(.A(mai_mai_n392_), .B(mai_mai_n173_), .C(mai_mai_n143_), .Y(mai_mai_n480_));
  NA2        m458(.A(mai_mai_n480_), .B(mai_mai_n479_), .Y(mai_mai_n481_));
  NO4        m459(.A(mai_mai_n481_), .B(mai_mai_n476_), .C(mai_mai_n473_), .D(mai_mai_n463_), .Y(mai_mai_n482_));
  NA2        m460(.A(mai_mai_n455_), .B(mai_mai_n388_), .Y(mai_mai_n483_));
  NO2        m461(.A(mai_mai_n483_), .B(mai_mai_n218_), .Y(mai_mai_n484_));
  NAi21      m462(.An(mai_mai_n209_), .B(mai_mai_n395_), .Y(mai_mai_n485_));
  NO2        m463(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n486_));
  NO2        m464(.A(i_0_), .B(mai_mai_n82_), .Y(mai_mai_n487_));
  NA3        m465(.A(mai_mai_n487_), .B(mai_mai_n486_), .C(mai_mai_n136_), .Y(mai_mai_n488_));
  OR3        m466(.A(mai_mai_n299_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n489_));
  NO2        m467(.A(mai_mai_n489_), .B(mai_mai_n488_), .Y(mai_mai_n490_));
  NA2        m468(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n491_));
  NA2        m469(.A(mai_mai_n309_), .B(mai_mai_n233_), .Y(mai_mai_n492_));
  OAI220     m470(.A0(mai_mai_n492_), .A1(mai_mai_n435_), .B0(mai_mai_n491_), .B1(mai_mai_n460_), .Y(mai_mai_n493_));
  NA3        m471(.A(mai_mai_n302_), .B(mai_mai_n217_), .C(mai_mai_n70_), .Y(mai_mai_n494_));
  NO2        m472(.A(mai_mai_n494_), .B(mai_mai_n466_), .Y(mai_mai_n495_));
  NO4        m473(.A(mai_mai_n495_), .B(mai_mai_n493_), .C(mai_mai_n490_), .D(mai_mai_n484_), .Y(mai_mai_n496_));
  NA3        m474(.A(mai_mai_n496_), .B(mai_mai_n482_), .C(mai_mai_n459_), .Y(mai_mai_n497_));
  NA3        m475(.A(mai_mai_n302_), .B(mai_mai_n170_), .C(mai_mai_n168_), .Y(mai_mai_n498_));
  INV        m476(.A(mai_mai_n498_), .Y(mai_mai_n499_));
  BUFFER     m477(.A(mai_mai_n283_), .Y(mai_mai_n500_));
  NA2        m478(.A(mai_mai_n500_), .B(mai_mai_n499_), .Y(mai_mai_n501_));
  NA2        m479(.A(mai_mai_n309_), .B(mai_mai_n158_), .Y(mai_mai_n502_));
  OAI210     m480(.A0(mai_mai_n502_), .A1(mai_mai_n226_), .B0(mai_mai_n303_), .Y(mai_mai_n503_));
  NA2        m481(.A(mai_mai_n503_), .B(mai_mai_n321_), .Y(mai_mai_n504_));
  NA2        m482(.A(mai_mai_n381_), .B(mai_mai_n219_), .Y(mai_mai_n505_));
  NA2        m483(.A(mai_mai_n356_), .B(mai_mai_n70_), .Y(mai_mai_n506_));
  NA2        m484(.A(mai_mai_n369_), .B(mai_mai_n365_), .Y(mai_mai_n507_));
  OR2        m485(.A(mai_mai_n505_), .B(mai_mai_n507_), .Y(mai_mai_n508_));
  NO2        m486(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n509_));
  NAi41      m487(.An(mai_mai_n506_), .B(mai_mai_n474_), .C(mai_mai_n509_), .D(mai_mai_n46_), .Y(mai_mai_n510_));
  AOI210     m488(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n416_), .Y(mai_mai_n511_));
  NA3        m489(.A(mai_mai_n511_), .B(mai_mai_n510_), .C(mai_mai_n508_), .Y(mai_mai_n512_));
  INV        m490(.A(mai_mai_n512_), .Y(mai_mai_n513_));
  NO2        m491(.A(i_7_), .B(mai_mai_n193_), .Y(mai_mai_n514_));
  OR2        m492(.A(mai_mai_n177_), .B(i_4_), .Y(mai_mai_n515_));
  NO2        m493(.A(mai_mai_n515_), .B(mai_mai_n82_), .Y(mai_mai_n516_));
  NA2        m494(.A(mai_mai_n516_), .B(mai_mai_n514_), .Y(mai_mai_n517_));
  NA4        m495(.A(mai_mai_n517_), .B(mai_mai_n513_), .C(mai_mai_n504_), .D(mai_mai_n501_), .Y(mai_mai_n518_));
  NA2        m496(.A(mai_mai_n387_), .B(mai_mai_n291_), .Y(mai_mai_n519_));
  NA2        m497(.A(mai_mai_n383_), .B(mai_mai_n519_), .Y(mai_mai_n520_));
  NA2        m498(.A(mai_mai_n997_), .B(mai_mai_n219_), .Y(mai_mai_n521_));
  NA2        m499(.A(mai_mai_n474_), .B(mai_mai_n27_), .Y(mai_mai_n522_));
  NO2        m500(.A(mai_mai_n522_), .B(mai_mai_n521_), .Y(mai_mai_n523_));
  NOi31      m501(.An(mai_mai_n312_), .B(mai_mai_n415_), .C(mai_mai_n38_), .Y(mai_mai_n524_));
  OAI210     m502(.A0(mai_mai_n524_), .A1(mai_mai_n523_), .B0(mai_mai_n520_), .Y(mai_mai_n525_));
  NO2        m503(.A(i_8_), .B(i_7_), .Y(mai_mai_n526_));
  OAI210     m504(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n527_));
  NA2        m505(.A(mai_mai_n527_), .B(mai_mai_n217_), .Y(mai_mai_n528_));
  OAI220     m506(.A0(mai_mai_n46_), .A1(mai_mai_n515_), .B0(mai_mai_n528_), .B1(mai_mai_n237_), .Y(mai_mai_n529_));
  NA2        m507(.A(mai_mai_n44_), .B(i_10_), .Y(mai_mai_n530_));
  NO2        m508(.A(mai_mai_n530_), .B(i_6_), .Y(mai_mai_n531_));
  NA3        m509(.A(mai_mai_n531_), .B(mai_mai_n529_), .C(mai_mai_n526_), .Y(mai_mai_n532_));
  AOI220     m510(.A0(mai_mai_n427_), .A1(mai_mai_n322_), .B0(mai_mai_n241_), .B1(mai_mai_n238_), .Y(mai_mai_n533_));
  OAI220     m511(.A0(mai_mai_n533_), .A1(mai_mai_n260_), .B0(mai_mai_n460_), .B1(mai_mai_n128_), .Y(mai_mai_n534_));
  NA2        m512(.A(mai_mai_n534_), .B(mai_mai_n263_), .Y(mai_mai_n535_));
  NOi31      m513(.An(mai_mai_n286_), .B(mai_mai_n297_), .C(mai_mai_n175_), .Y(mai_mai_n536_));
  NO2        m514(.A(mai_mai_n215_), .B(mai_mai_n44_), .Y(mai_mai_n537_));
  NO2        m515(.A(mai_mai_n151_), .B(i_5_), .Y(mai_mai_n538_));
  NA3        m516(.A(mai_mai_n538_), .B(mai_mai_n403_), .C(mai_mai_n315_), .Y(mai_mai_n539_));
  NO2        m517(.A(mai_mai_n539_), .B(mai_mai_n537_), .Y(mai_mai_n540_));
  OAI210     m518(.A0(mai_mai_n540_), .A1(mai_mai_n536_), .B0(mai_mai_n455_), .Y(mai_mai_n541_));
  NA4        m519(.A(mai_mai_n541_), .B(mai_mai_n535_), .C(mai_mai_n532_), .D(mai_mai_n525_), .Y(mai_mai_n542_));
  NA3        m520(.A(mai_mai_n211_), .B(mai_mai_n68_), .C(mai_mai_n44_), .Y(mai_mai_n543_));
  NA2        m521(.A(mai_mai_n279_), .B(mai_mai_n80_), .Y(mai_mai_n544_));
  AOI210     m522(.A0(mai_mai_n543_), .A1(mai_mai_n346_), .B0(mai_mai_n544_), .Y(mai_mai_n545_));
  NA2        m523(.A(mai_mai_n292_), .B(mai_mai_n283_), .Y(mai_mai_n546_));
  NO2        m524(.A(mai_mai_n546_), .B(mai_mai_n167_), .Y(mai_mai_n547_));
  NA2        m525(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n548_));
  NA2        m526(.A(mai_mai_n447_), .B(mai_mai_n215_), .Y(mai_mai_n549_));
  NO2        m527(.A(mai_mai_n548_), .B(mai_mai_n549_), .Y(mai_mai_n550_));
  NO3        m528(.A(mai_mai_n550_), .B(mai_mai_n547_), .C(mai_mai_n545_), .Y(mai_mai_n551_));
  NO4        m529(.A(mai_mai_n246_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n552_));
  NO3        m530(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n553_));
  NO2        m531(.A(mai_mai_n227_), .B(mai_mai_n36_), .Y(mai_mai_n554_));
  AN2        m532(.A(mai_mai_n554_), .B(mai_mai_n553_), .Y(mai_mai_n555_));
  OA210      m533(.A0(mai_mai_n555_), .A1(mai_mai_n552_), .B0(mai_mai_n356_), .Y(mai_mai_n556_));
  NO2        m534(.A(mai_mai_n415_), .B(i_1_), .Y(mai_mai_n557_));
  NOi31      m535(.An(mai_mai_n557_), .B(mai_mai_n452_), .C(mai_mai_n70_), .Y(mai_mai_n558_));
  AN4        m536(.A(mai_mai_n558_), .B(mai_mai_n412_), .C(mai_mai_n486_), .D(i_2_), .Y(mai_mai_n559_));
  NO2        m537(.A(mai_mai_n425_), .B(mai_mai_n171_), .Y(mai_mai_n560_));
  NO3        m538(.A(mai_mai_n560_), .B(mai_mai_n559_), .C(mai_mai_n556_), .Y(mai_mai_n561_));
  NOi21      m539(.An(i_10_), .B(i_6_), .Y(mai_mai_n562_));
  NO2        m540(.A(mai_mai_n111_), .B(mai_mai_n23_), .Y(mai_mai_n563_));
  NA2        m541(.A(mai_mai_n312_), .B(mai_mai_n158_), .Y(mai_mai_n564_));
  AOI220     m542(.A0(mai_mai_n564_), .A1(mai_mai_n436_), .B0(mai_mai_n166_), .B1(mai_mai_n176_), .Y(mai_mai_n565_));
  NOi21      m543(.An(mai_mai_n140_), .B(mai_mai_n328_), .Y(mai_mai_n566_));
  NO2        m544(.A(mai_mai_n566_), .B(mai_mai_n565_), .Y(mai_mai_n567_));
  INV        m545(.A(mai_mai_n315_), .Y(mai_mai_n568_));
  NO2        m546(.A(i_12_), .B(mai_mai_n82_), .Y(mai_mai_n569_));
  NO3        m547(.A(i_4_), .B(mai_mai_n338_), .C(mai_mai_n297_), .Y(mai_mai_n570_));
  OR2        m548(.A(i_2_), .B(i_5_), .Y(mai_mai_n571_));
  OR2        m549(.A(mai_mai_n571_), .B(mai_mai_n407_), .Y(mai_mai_n572_));
  NA2        m550(.A(mai_mai_n371_), .B(mai_mai_n238_), .Y(mai_mai_n573_));
  AOI210     m551(.A0(mai_mai_n573_), .A1(mai_mai_n572_), .B0(mai_mai_n485_), .Y(mai_mai_n574_));
  NO2        m552(.A(mai_mai_n574_), .B(mai_mai_n570_), .Y(mai_mai_n575_));
  NA4        m553(.A(mai_mai_n575_), .B(mai_mai_n567_), .C(mai_mai_n561_), .D(mai_mai_n551_), .Y(mai_mai_n576_));
  NO4        m554(.A(mai_mai_n576_), .B(mai_mai_n542_), .C(mai_mai_n518_), .D(mai_mai_n497_), .Y(mai_mai_n577_));
  NA4        m555(.A(mai_mai_n577_), .B(mai_mai_n444_), .C(mai_mai_n355_), .D(mai_mai_n308_), .Y(mai7));
  NO2        m556(.A(mai_mai_n89_), .B(mai_mai_n52_), .Y(mai_mai_n579_));
  NA2        m557(.A(mai_mai_n474_), .B(mai_mai_n80_), .Y(mai_mai_n580_));
  NA2        m558(.A(i_11_), .B(mai_mai_n187_), .Y(mai_mai_n581_));
  NA3        m559(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n582_));
  NO2        m560(.A(mai_mai_n231_), .B(i_4_), .Y(mai_mai_n583_));
  NA2        m561(.A(mai_mai_n583_), .B(i_8_), .Y(mai_mai_n584_));
  NO2        m562(.A(mai_mai_n102_), .B(mai_mai_n582_), .Y(mai_mai_n585_));
  NA2        m563(.A(i_2_), .B(mai_mai_n82_), .Y(mai_mai_n586_));
  OAI210     m564(.A0(mai_mai_n83_), .A1(mai_mai_n197_), .B0(mai_mai_n198_), .Y(mai_mai_n587_));
  NO2        m565(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n588_));
  NA2        m566(.A(i_4_), .B(i_8_), .Y(mai_mai_n589_));
  AOI210     m567(.A0(mai_mai_n589_), .A1(mai_mai_n302_), .B0(mai_mai_n588_), .Y(mai_mai_n590_));
  OAI220     m568(.A0(mai_mai_n590_), .A1(mai_mai_n586_), .B0(mai_mai_n587_), .B1(i_13_), .Y(mai_mai_n591_));
  NO3        m569(.A(mai_mai_n591_), .B(mai_mai_n585_), .C(mai_mai_n579_), .Y(mai_mai_n592_));
  AOI210     m570(.A0(mai_mai_n123_), .A1(mai_mai_n59_), .B0(i_10_), .Y(mai_mai_n593_));
  AOI210     m571(.A0(mai_mai_n593_), .A1(mai_mai_n231_), .B0(mai_mai_n155_), .Y(mai_mai_n594_));
  OR2        m572(.A(i_6_), .B(i_10_), .Y(mai_mai_n595_));
  NO2        m573(.A(mai_mai_n595_), .B(mai_mai_n23_), .Y(mai_mai_n596_));
  OR3        m574(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n597_));
  NO3        m575(.A(mai_mai_n597_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n598_));
  INV        m576(.A(mai_mai_n194_), .Y(mai_mai_n599_));
  NO2        m577(.A(mai_mai_n598_), .B(mai_mai_n596_), .Y(mai_mai_n600_));
  OA220      m578(.A0(mai_mai_n600_), .A1(mai_mai_n568_), .B0(mai_mai_n594_), .B1(mai_mai_n265_), .Y(mai_mai_n601_));
  AOI210     m579(.A0(mai_mai_n601_), .A1(mai_mai_n592_), .B0(mai_mai_n60_), .Y(mai_mai_n602_));
  NOi21      m580(.An(i_11_), .B(i_7_), .Y(mai_mai_n603_));
  AO210      m581(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n604_));
  NO2        m582(.A(mai_mai_n604_), .B(mai_mai_n603_), .Y(mai_mai_n605_));
  NA2        m583(.A(mai_mai_n605_), .B(mai_mai_n199_), .Y(mai_mai_n606_));
  NA3        m584(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n607_));
  NO2        m585(.A(mai_mai_n606_), .B(mai_mai_n60_), .Y(mai_mai_n608_));
  NO3        m586(.A(mai_mai_n254_), .B(mai_mai_n201_), .C(mai_mai_n581_), .Y(mai_mai_n609_));
  OAI210     m587(.A0(mai_mai_n609_), .A1(mai_mai_n220_), .B0(mai_mai_n60_), .Y(mai_mai_n610_));
  OR2        m588(.A(mai_mai_n201_), .B(mai_mai_n105_), .Y(mai_mai_n611_));
  NO2        m589(.A(mai_mai_n60_), .B(i_9_), .Y(mai_mai_n612_));
  NO2        m590(.A(i_1_), .B(i_12_), .Y(mai_mai_n613_));
  INV        m591(.A(mai_mai_n610_), .Y(mai_mai_n614_));
  OAI210     m592(.A0(mai_mai_n614_), .A1(mai_mai_n608_), .B0(i_6_), .Y(mai_mai_n615_));
  NO2        m593(.A(mai_mai_n607_), .B(mai_mai_n105_), .Y(mai_mai_n616_));
  NA2        m594(.A(mai_mai_n616_), .B(mai_mai_n569_), .Y(mai_mai_n617_));
  NO2        m595(.A(i_6_), .B(i_11_), .Y(mai_mai_n618_));
  NA2        m596(.A(mai_mai_n617_), .B(mai_mai_n453_), .Y(mai_mai_n619_));
  NO4        m597(.A(mai_mai_n208_), .B(mai_mai_n123_), .C(i_13_), .D(mai_mai_n82_), .Y(mai_mai_n620_));
  NA2        m598(.A(mai_mai_n620_), .B(mai_mai_n612_), .Y(mai_mai_n621_));
  NA2        m599(.A(mai_mai_n231_), .B(i_6_), .Y(mai_mai_n622_));
  NO3        m600(.A(mai_mai_n595_), .B(mai_mai_n227_), .C(mai_mai_n23_), .Y(mai_mai_n623_));
  AOI210     m601(.A0(i_1_), .A1(mai_mai_n255_), .B0(mai_mai_n623_), .Y(mai_mai_n624_));
  OAI210     m602(.A0(mai_mai_n624_), .A1(mai_mai_n44_), .B0(mai_mai_n621_), .Y(mai_mai_n625_));
  NA3        m603(.A(mai_mai_n526_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n626_));
  NA2        m604(.A(mai_mai_n132_), .B(i_9_), .Y(mai_mai_n627_));
  NA3        m605(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n629_));
  NA3        m607(.A(mai_mai_n629_), .B(mai_mai_n264_), .C(mai_mai_n44_), .Y(mai_mai_n630_));
  OAI220     m608(.A0(mai_mai_n630_), .A1(mai_mai_n628_), .B0(mai_mai_n627_), .B1(mai_mai_n996_), .Y(mai_mai_n631_));
  NA3        m609(.A(mai_mai_n612_), .B(mai_mai_n315_), .C(i_6_), .Y(mai_mai_n632_));
  NO2        m610(.A(mai_mai_n632_), .B(mai_mai_n23_), .Y(mai_mai_n633_));
  AOI210     m611(.A0(mai_mai_n467_), .A1(mai_mai_n418_), .B0(mai_mai_n236_), .Y(mai_mai_n634_));
  NO2        m612(.A(mai_mai_n634_), .B(mai_mai_n586_), .Y(mai_mai_n635_));
  NAi21      m613(.An(mai_mai_n626_), .B(mai_mai_n88_), .Y(mai_mai_n636_));
  NA2        m614(.A(mai_mai_n629_), .B(mai_mai_n264_), .Y(mai_mai_n637_));
  NO2        m615(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n638_));
  NA2        m616(.A(mai_mai_n638_), .B(mai_mai_n24_), .Y(mai_mai_n639_));
  OAI210     m617(.A0(mai_mai_n639_), .A1(mai_mai_n637_), .B0(mai_mai_n636_), .Y(mai_mai_n640_));
  OR4        m618(.A(mai_mai_n640_), .B(mai_mai_n635_), .C(mai_mai_n633_), .D(mai_mai_n631_), .Y(mai_mai_n641_));
  NO3        m619(.A(mai_mai_n641_), .B(mai_mai_n625_), .C(mai_mai_n619_), .Y(mai_mai_n642_));
  NO2        m620(.A(mai_mai_n231_), .B(mai_mai_n98_), .Y(mai_mai_n643_));
  NO2        m621(.A(mai_mai_n643_), .B(mai_mai_n603_), .Y(mai_mai_n644_));
  NA2        m622(.A(mai_mai_n644_), .B(i_1_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n645_), .B(mai_mai_n597_), .Y(mai_mai_n646_));
  NO2        m624(.A(mai_mai_n414_), .B(mai_mai_n82_), .Y(mai_mai_n647_));
  NA2        m625(.A(mai_mai_n646_), .B(mai_mai_n46_), .Y(mai_mai_n648_));
  NA2        m626(.A(i_3_), .B(mai_mai_n187_), .Y(mai_mai_n649_));
  NO2        m627(.A(mai_mai_n649_), .B(mai_mai_n111_), .Y(mai_mai_n650_));
  AN2        m628(.A(mai_mai_n650_), .B(mai_mai_n531_), .Y(mai_mai_n651_));
  NO2        m629(.A(mai_mai_n227_), .B(mai_mai_n44_), .Y(mai_mai_n652_));
  NO3        m630(.A(mai_mai_n652_), .B(mai_mai_n305_), .C(mai_mai_n232_), .Y(mai_mai_n653_));
  NO2        m631(.A(mai_mai_n112_), .B(mai_mai_n37_), .Y(mai_mai_n654_));
  NO2        m632(.A(mai_mai_n654_), .B(i_6_), .Y(mai_mai_n655_));
  NO2        m633(.A(mai_mai_n82_), .B(i_9_), .Y(mai_mai_n656_));
  NO2        m634(.A(mai_mai_n656_), .B(mai_mai_n60_), .Y(mai_mai_n657_));
  NO2        m635(.A(mai_mai_n657_), .B(mai_mai_n613_), .Y(mai_mai_n658_));
  NO4        m636(.A(mai_mai_n658_), .B(mai_mai_n655_), .C(mai_mai_n653_), .D(i_4_), .Y(mai_mai_n659_));
  NA2        m637(.A(i_1_), .B(i_3_), .Y(mai_mai_n660_));
  NO2        m638(.A(mai_mai_n454_), .B(mai_mai_n89_), .Y(mai_mai_n661_));
  AOI210     m639(.A0(mai_mai_n652_), .A1(mai_mai_n562_), .B0(mai_mai_n661_), .Y(mai_mai_n662_));
  NO2        m640(.A(mai_mai_n662_), .B(mai_mai_n660_), .Y(mai_mai_n663_));
  NO3        m641(.A(mai_mai_n663_), .B(mai_mai_n659_), .C(mai_mai_n651_), .Y(mai_mai_n664_));
  NA4        m642(.A(mai_mai_n664_), .B(mai_mai_n648_), .C(mai_mai_n642_), .D(mai_mai_n615_), .Y(mai_mai_n665_));
  NO3        m643(.A(i_11_), .B(i_3_), .C(i_7_), .Y(mai_mai_n666_));
  NOi21      m644(.An(mai_mai_n666_), .B(i_10_), .Y(mai_mai_n667_));
  OA210      m645(.A0(mai_mai_n667_), .A1(mai_mai_n239_), .B0(mai_mai_n82_), .Y(mai_mai_n668_));
  NA2        m646(.A(mai_mai_n369_), .B(mai_mai_n368_), .Y(mai_mai_n669_));
  NA3        m647(.A(mai_mai_n474_), .B(mai_mai_n509_), .C(mai_mai_n46_), .Y(mai_mai_n670_));
  NA2        m648(.A(mai_mai_n670_), .B(mai_mai_n669_), .Y(mai_mai_n671_));
  OAI210     m649(.A0(mai_mai_n671_), .A1(mai_mai_n668_), .B0(i_1_), .Y(mai_mai_n672_));
  AOI210     m650(.A0(mai_mai_n264_), .A1(mai_mai_n94_), .B0(i_1_), .Y(mai_mai_n673_));
  NO2        m651(.A(mai_mai_n367_), .B(i_2_), .Y(mai_mai_n674_));
  NA2        m652(.A(mai_mai_n674_), .B(mai_mai_n673_), .Y(mai_mai_n675_));
  OAI210     m653(.A0(mai_mai_n632_), .A1(mai_mai_n448_), .B0(mai_mai_n675_), .Y(mai_mai_n676_));
  INV        m654(.A(mai_mai_n676_), .Y(mai_mai_n677_));
  AOI210     m655(.A0(mai_mai_n677_), .A1(mai_mai_n672_), .B0(i_13_), .Y(mai_mai_n678_));
  OR2        m656(.A(i_11_), .B(i_7_), .Y(mai_mai_n679_));
  NO2        m657(.A(mai_mai_n52_), .B(i_12_), .Y(mai_mai_n680_));
  INV        m658(.A(mai_mai_n680_), .Y(mai_mai_n681_));
  NO2        m659(.A(mai_mai_n469_), .B(mai_mai_n24_), .Y(mai_mai_n682_));
  AOI220     m660(.A0(mai_mai_n682_), .A1(mai_mai_n647_), .B0(mai_mai_n239_), .B1(mai_mai_n126_), .Y(mai_mai_n683_));
  OAI220     m661(.A0(mai_mai_n683_), .A1(mai_mai_n41_), .B0(mai_mai_n681_), .B1(mai_mai_n89_), .Y(mai_mai_n684_));
  INV        m662(.A(mai_mai_n684_), .Y(mai_mai_n685_));
  NA2        m663(.A(mai_mai_n384_), .B(mai_mai_n629_), .Y(mai_mai_n686_));
  NO2        m664(.A(mai_mai_n686_), .B(mai_mai_n237_), .Y(mai_mai_n687_));
  AOI210     m665(.A0(mai_mai_n448_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n688_));
  NOi31      m666(.An(mai_mai_n688_), .B(mai_mai_n580_), .C(mai_mai_n44_), .Y(mai_mai_n689_));
  NA2        m667(.A(mai_mai_n122_), .B(i_13_), .Y(mai_mai_n690_));
  NO2        m668(.A(mai_mai_n628_), .B(mai_mai_n111_), .Y(mai_mai_n691_));
  INV        m669(.A(mai_mai_n691_), .Y(mai_mai_n692_));
  OAI220     m670(.A0(mai_mai_n692_), .A1(mai_mai_n68_), .B0(mai_mai_n690_), .B1(mai_mai_n673_), .Y(mai_mai_n693_));
  NA2        m671(.A(mai_mai_n26_), .B(mai_mai_n187_), .Y(mai_mai_n694_));
  NA2        m672(.A(mai_mai_n694_), .B(i_7_), .Y(mai_mai_n695_));
  NO3        m673(.A(mai_mai_n469_), .B(mai_mai_n231_), .C(mai_mai_n82_), .Y(mai_mai_n696_));
  NA2        m674(.A(mai_mai_n696_), .B(mai_mai_n695_), .Y(mai_mai_n697_));
  AOI220     m675(.A0(mai_mai_n384_), .A1(mai_mai_n629_), .B0(mai_mai_n88_), .B1(mai_mai_n99_), .Y(mai_mai_n698_));
  OAI220     m676(.A0(mai_mai_n698_), .A1(mai_mai_n584_), .B0(mai_mai_n697_), .B1(mai_mai_n599_), .Y(mai_mai_n699_));
  NO4        m677(.A(mai_mai_n699_), .B(mai_mai_n693_), .C(mai_mai_n689_), .D(mai_mai_n687_), .Y(mai_mai_n700_));
  OR2        m678(.A(i_11_), .B(i_6_), .Y(mai_mai_n701_));
  NA3        m679(.A(mai_mai_n583_), .B(mai_mai_n694_), .C(i_7_), .Y(mai_mai_n702_));
  AOI210     m680(.A0(mai_mai_n702_), .A1(mai_mai_n692_), .B0(mai_mai_n701_), .Y(mai_mai_n703_));
  NA3        m681(.A(mai_mai_n408_), .B(mai_mai_n588_), .C(mai_mai_n94_), .Y(mai_mai_n704_));
  NA2        m682(.A(mai_mai_n618_), .B(i_13_), .Y(mai_mai_n705_));
  NA2        m683(.A(mai_mai_n99_), .B(mai_mai_n694_), .Y(mai_mai_n706_));
  NAi21      m684(.An(i_11_), .B(i_12_), .Y(mai_mai_n707_));
  NOi41      m685(.An(mai_mai_n107_), .B(mai_mai_n707_), .C(i_13_), .D(mai_mai_n82_), .Y(mai_mai_n708_));
  NA2        m686(.A(mai_mai_n708_), .B(mai_mai_n706_), .Y(mai_mai_n709_));
  NA3        m687(.A(mai_mai_n709_), .B(mai_mai_n705_), .C(mai_mai_n704_), .Y(mai_mai_n710_));
  OAI210     m688(.A0(mai_mai_n710_), .A1(mai_mai_n703_), .B0(mai_mai_n60_), .Y(mai_mai_n711_));
  NO2        m689(.A(i_2_), .B(i_12_), .Y(mai_mai_n712_));
  NA2        m690(.A(mai_mai_n366_), .B(mai_mai_n712_), .Y(mai_mai_n713_));
  NA2        m691(.A(i_8_), .B(mai_mai_n25_), .Y(mai_mai_n714_));
  NO3        m692(.A(mai_mai_n714_), .B(mai_mai_n382_), .C(mai_mai_n583_), .Y(mai_mai_n715_));
  OAI210     m693(.A0(mai_mai_n715_), .A1(mai_mai_n368_), .B0(mai_mai_n366_), .Y(mai_mai_n716_));
  NO2        m694(.A(mai_mai_n123_), .B(i_2_), .Y(mai_mai_n717_));
  NA2        m695(.A(mai_mai_n717_), .B(mai_mai_n613_), .Y(mai_mai_n718_));
  NA3        m696(.A(mai_mai_n718_), .B(mai_mai_n716_), .C(mai_mai_n713_), .Y(mai_mai_n719_));
  NA3        m697(.A(mai_mai_n719_), .B(mai_mai_n45_), .C(mai_mai_n219_), .Y(mai_mai_n720_));
  NA4        m698(.A(mai_mai_n720_), .B(mai_mai_n711_), .C(mai_mai_n700_), .D(mai_mai_n685_), .Y(mai_mai_n721_));
  OR4        m699(.A(mai_mai_n721_), .B(mai_mai_n678_), .C(mai_mai_n665_), .D(mai_mai_n602_), .Y(mai5));
  NA2        m700(.A(mai_mai_n644_), .B(mai_mai_n267_), .Y(mai_mai_n723_));
  AN2        m701(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n724_));
  NA3        m702(.A(mai_mai_n724_), .B(mai_mai_n712_), .C(mai_mai_n105_), .Y(mai_mai_n725_));
  NO2        m703(.A(mai_mai_n584_), .B(i_11_), .Y(mai_mai_n726_));
  NA2        m704(.A(mai_mai_n83_), .B(mai_mai_n726_), .Y(mai_mai_n727_));
  NA3        m705(.A(mai_mai_n727_), .B(mai_mai_n725_), .C(mai_mai_n723_), .Y(mai_mai_n728_));
  NO3        m706(.A(i_11_), .B(mai_mai_n231_), .C(i_13_), .Y(mai_mai_n729_));
  NO2        m707(.A(mai_mai_n119_), .B(mai_mai_n23_), .Y(mai_mai_n730_));
  NA2        m708(.A(i_12_), .B(i_8_), .Y(mai_mai_n731_));
  OAI210     m709(.A0(mai_mai_n46_), .A1(i_3_), .B0(mai_mai_n731_), .Y(mai_mai_n732_));
  INV        m710(.A(mai_mai_n447_), .Y(mai_mai_n733_));
  AOI220     m711(.A0(mai_mai_n315_), .A1(mai_mai_n563_), .B0(mai_mai_n732_), .B1(mai_mai_n730_), .Y(mai_mai_n734_));
  INV        m712(.A(mai_mai_n734_), .Y(mai_mai_n735_));
  NO2        m713(.A(mai_mai_n735_), .B(mai_mai_n728_), .Y(mai_mai_n736_));
  INV        m714(.A(mai_mai_n165_), .Y(mai_mai_n737_));
  INV        m715(.A(mai_mai_n239_), .Y(mai_mai_n738_));
  OAI210     m716(.A0(mai_mai_n674_), .A1(mai_mai_n449_), .B0(mai_mai_n107_), .Y(mai_mai_n739_));
  AOI210     m717(.A0(mai_mai_n739_), .A1(mai_mai_n738_), .B0(mai_mai_n737_), .Y(mai_mai_n740_));
  NO2        m718(.A(mai_mai_n454_), .B(mai_mai_n26_), .Y(mai_mai_n741_));
  NO2        m719(.A(mai_mai_n741_), .B(mai_mai_n418_), .Y(mai_mai_n742_));
  NA2        m720(.A(mai_mai_n742_), .B(i_2_), .Y(mai_mai_n743_));
  INV        m721(.A(mai_mai_n743_), .Y(mai_mai_n744_));
  AOI210     m722(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n415_), .Y(mai_mai_n745_));
  AOI210     m723(.A0(mai_mai_n745_), .A1(mai_mai_n744_), .B0(mai_mai_n740_), .Y(mai_mai_n746_));
  NO2        m724(.A(mai_mai_n184_), .B(mai_mai_n120_), .Y(mai_mai_n747_));
  OAI210     m725(.A0(mai_mai_n747_), .A1(mai_mai_n730_), .B0(i_2_), .Y(mai_mai_n748_));
  INV        m726(.A(mai_mai_n166_), .Y(mai_mai_n749_));
  NO3        m727(.A(mai_mai_n604_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n750_));
  AOI210     m728(.A0(mai_mai_n749_), .A1(mai_mai_n83_), .B0(mai_mai_n750_), .Y(mai_mai_n751_));
  AOI210     m729(.A0(mai_mai_n751_), .A1(mai_mai_n748_), .B0(mai_mai_n187_), .Y(mai_mai_n752_));
  OA210      m730(.A0(mai_mai_n605_), .A1(mai_mai_n121_), .B0(i_13_), .Y(mai_mai_n753_));
  NA2        m731(.A(mai_mai_n145_), .B(mai_mai_n581_), .Y(mai_mai_n754_));
  NO2        m732(.A(mai_mai_n754_), .B(mai_mai_n371_), .Y(mai_mai_n755_));
  AOI210     m733(.A0(mai_mai_n201_), .A1(mai_mai_n142_), .B0(mai_mai_n509_), .Y(mai_mai_n756_));
  NA2        m734(.A(mai_mai_n756_), .B(mai_mai_n418_), .Y(mai_mai_n757_));
  NO2        m735(.A(mai_mai_n99_), .B(mai_mai_n44_), .Y(mai_mai_n758_));
  INV        m736(.A(mai_mai_n298_), .Y(mai_mai_n759_));
  NA4        m737(.A(mai_mai_n759_), .B(mai_mai_n302_), .C(mai_mai_n119_), .D(mai_mai_n42_), .Y(mai_mai_n760_));
  OAI210     m738(.A0(mai_mai_n760_), .A1(mai_mai_n758_), .B0(mai_mai_n757_), .Y(mai_mai_n761_));
  NO4        m739(.A(mai_mai_n761_), .B(mai_mai_n755_), .C(mai_mai_n753_), .D(mai_mai_n752_), .Y(mai_mai_n762_));
  NA2        m740(.A(mai_mai_n563_), .B(mai_mai_n28_), .Y(mai_mai_n763_));
  NA2        m741(.A(mai_mai_n729_), .B(mai_mai_n271_), .Y(mai_mai_n764_));
  NA2        m742(.A(mai_mai_n764_), .B(mai_mai_n763_), .Y(mai_mai_n765_));
  NO2        m743(.A(mai_mai_n59_), .B(i_12_), .Y(mai_mai_n766_));
  NO2        m744(.A(mai_mai_n766_), .B(mai_mai_n121_), .Y(mai_mai_n767_));
  NO2        m745(.A(mai_mai_n767_), .B(mai_mai_n581_), .Y(mai_mai_n768_));
  AOI220     m746(.A0(mai_mai_n768_), .A1(mai_mai_n36_), .B0(mai_mai_n765_), .B1(mai_mai_n46_), .Y(mai_mai_n769_));
  NA4        m747(.A(mai_mai_n769_), .B(mai_mai_n762_), .C(mai_mai_n746_), .D(mai_mai_n736_), .Y(mai6));
  NO3        m748(.A(mai_mai_n250_), .B(mai_mai_n304_), .C(i_1_), .Y(mai_mai_n771_));
  NO2        m749(.A(mai_mai_n179_), .B(mai_mai_n133_), .Y(mai_mai_n772_));
  OAI210     m750(.A0(mai_mai_n772_), .A1(mai_mai_n771_), .B0(mai_mai_n717_), .Y(mai_mai_n773_));
  NO2        m751(.A(mai_mai_n214_), .B(mai_mai_n477_), .Y(mai_mai_n774_));
  INV        m752(.A(mai_mai_n327_), .Y(mai_mai_n775_));
  AO210      m753(.A0(mai_mai_n775_), .A1(mai_mai_n773_), .B0(i_12_), .Y(mai_mai_n776_));
  NA2        m754(.A(mai_mai_n372_), .B(mai_mai_n332_), .Y(mai_mai_n777_));
  NA2        m755(.A(mai_mai_n569_), .B(mai_mai_n60_), .Y(mai_mai_n778_));
  NA2        m756(.A(mai_mai_n667_), .B(mai_mai_n68_), .Y(mai_mai_n779_));
  NA3        m757(.A(mai_mai_n779_), .B(mai_mai_n778_), .C(mai_mai_n777_), .Y(mai_mai_n780_));
  NA2        m758(.A(mai_mai_n780_), .B(mai_mai_n70_), .Y(mai_mai_n781_));
  INV        m759(.A(mai_mai_n326_), .Y(mai_mai_n782_));
  NA2        m760(.A(mai_mai_n72_), .B(mai_mai_n126_), .Y(mai_mai_n783_));
  INV        m761(.A(mai_mai_n119_), .Y(mai_mai_n784_));
  NA2        m762(.A(mai_mai_n784_), .B(mai_mai_n46_), .Y(mai_mai_n785_));
  AOI210     m763(.A0(mai_mai_n785_), .A1(mai_mai_n783_), .B0(mai_mai_n782_), .Y(mai_mai_n786_));
  NO2        m764(.A(mai_mai_n507_), .B(mai_mai_n179_), .Y(mai_mai_n787_));
  NO2        m765(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n788_));
  NA3        m766(.A(mai_mai_n788_), .B(mai_mai_n465_), .C(mai_mai_n388_), .Y(mai_mai_n789_));
  NAi32      m767(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n790_));
  NO2        m768(.A(mai_mai_n701_), .B(mai_mai_n790_), .Y(mai_mai_n791_));
  OAI210     m769(.A0(mai_mai_n666_), .A1(mai_mai_n554_), .B0(mai_mai_n553_), .Y(mai_mai_n792_));
  NAi31      m770(.An(mai_mai_n791_), .B(mai_mai_n792_), .C(mai_mai_n789_), .Y(mai_mai_n793_));
  OR3        m771(.A(mai_mai_n793_), .B(mai_mai_n787_), .C(mai_mai_n786_), .Y(mai_mai_n794_));
  NO2        m772(.A(mai_mai_n679_), .B(i_2_), .Y(mai_mai_n795_));
  NA2        m773(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n796_));
  NO2        m774(.A(mai_mai_n796_), .B(mai_mai_n407_), .Y(mai_mai_n797_));
  NA2        m775(.A(mai_mai_n797_), .B(mai_mai_n795_), .Y(mai_mai_n798_));
  AO210      m776(.A0(mai_mai_n360_), .A1(mai_mai_n350_), .B0(mai_mai_n394_), .Y(mai_mai_n799_));
  NA3        m777(.A(mai_mai_n799_), .B(mai_mai_n251_), .C(i_7_), .Y(mai_mai_n800_));
  OR2        m778(.A(mai_mai_n605_), .B(mai_mai_n449_), .Y(mai_mai_n801_));
  NA3        m779(.A(mai_mai_n801_), .B(mai_mai_n141_), .C(mai_mai_n66_), .Y(mai_mai_n802_));
  AO210      m780(.A0(mai_mai_n483_), .A1(mai_mai_n733_), .B0(mai_mai_n36_), .Y(mai_mai_n803_));
  NA4        m781(.A(mai_mai_n803_), .B(mai_mai_n802_), .C(mai_mai_n800_), .D(mai_mai_n798_), .Y(mai_mai_n804_));
  NO2        m782(.A(i_6_), .B(i_11_), .Y(mai_mai_n805_));
  AOI220     m783(.A0(mai_mai_n805_), .A1(mai_mai_n553_), .B0(mai_mai_n774_), .B1(mai_mai_n695_), .Y(mai_mai_n806_));
  NA3        m784(.A(mai_mai_n371_), .B(mai_mai_n233_), .C(mai_mai_n141_), .Y(mai_mai_n807_));
  NA2        m785(.A(mai_mai_n394_), .B(mai_mai_n67_), .Y(mai_mai_n808_));
  NA4        m786(.A(mai_mai_n808_), .B(mai_mai_n807_), .C(mai_mai_n806_), .D(mai_mai_n587_), .Y(mai_mai_n809_));
  AOI210     m787(.A0(mai_mai_n449_), .A1(mai_mai_n447_), .B0(mai_mai_n552_), .Y(mai_mai_n810_));
  NO2        m788(.A(mai_mai_n595_), .B(mai_mai_n99_), .Y(mai_mai_n811_));
  OAI210     m789(.A0(mai_mai_n811_), .A1(mai_mai_n108_), .B0(mai_mai_n405_), .Y(mai_mai_n812_));
  INV        m790(.A(mai_mai_n238_), .Y(mai_mai_n813_));
  INV        m791(.A(mai_mai_n572_), .Y(mai_mai_n814_));
  NA3        m792(.A(mai_mai_n814_), .B(mai_mai_n326_), .C(i_7_), .Y(mai_mai_n815_));
  NA3        m793(.A(mai_mai_n815_), .B(mai_mai_n812_), .C(mai_mai_n810_), .Y(mai_mai_n816_));
  NO4        m794(.A(mai_mai_n816_), .B(mai_mai_n809_), .C(mai_mai_n804_), .D(mai_mai_n794_), .Y(mai_mai_n817_));
  NA4        m795(.A(mai_mai_n817_), .B(mai_mai_n781_), .C(mai_mai_n776_), .D(mai_mai_n378_), .Y(mai3));
  NA2        m796(.A(i_6_), .B(i_7_), .Y(mai_mai_n819_));
  NO2        m797(.A(mai_mai_n819_), .B(i_0_), .Y(mai_mai_n820_));
  NO2        m798(.A(i_11_), .B(mai_mai_n231_), .Y(mai_mai_n821_));
  OAI210     m799(.A0(mai_mai_n820_), .A1(mai_mai_n286_), .B0(mai_mai_n821_), .Y(mai_mai_n822_));
  NO2        m800(.A(mai_mai_n822_), .B(mai_mai_n187_), .Y(mai_mai_n823_));
  NO3        m801(.A(mai_mai_n450_), .B(mai_mai_n86_), .C(mai_mai_n44_), .Y(mai_mai_n824_));
  OA210      m802(.A0(mai_mai_n824_), .A1(mai_mai_n823_), .B0(mai_mai_n168_), .Y(mai_mai_n825_));
  NA2        m803(.A(mai_mai_n807_), .B(mai_mai_n370_), .Y(mai_mai_n826_));
  NA2        m804(.A(mai_mai_n826_), .B(mai_mai_n40_), .Y(mai_mai_n827_));
  NO3        m805(.A(mai_mai_n611_), .B(mai_mai_n454_), .C(mai_mai_n126_), .Y(mai_mai_n828_));
  AN2        m806(.A(mai_mai_n452_), .B(mai_mai_n53_), .Y(mai_mai_n829_));
  NO2        m807(.A(mai_mai_n829_), .B(mai_mai_n828_), .Y(mai_mai_n830_));
  AOI210     m808(.A0(mai_mai_n830_), .A1(mai_mai_n827_), .B0(mai_mai_n48_), .Y(mai_mai_n831_));
  NO4        m809(.A(mai_mai_n375_), .B(mai_mai_n381_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n832_));
  NA2        m810(.A(mai_mai_n688_), .B(mai_mai_n656_), .Y(mai_mai_n833_));
  NA2        m811(.A(mai_mai_n330_), .B(mai_mai_n438_), .Y(mai_mai_n834_));
  OAI220     m812(.A0(mai_mai_n834_), .A1(mai_mai_n833_), .B0(mai_mai_n999_), .B1(mai_mai_n60_), .Y(mai_mai_n835_));
  NOi21      m813(.An(i_5_), .B(i_9_), .Y(mai_mai_n836_));
  NA2        m814(.A(mai_mai_n836_), .B(mai_mai_n446_), .Y(mai_mai_n837_));
  BUFFER     m815(.A(mai_mai_n264_), .Y(mai_mai_n838_));
  NA2        m816(.A(mai_mai_n838_), .B(mai_mai_n467_), .Y(mai_mai_n839_));
  NO3        m817(.A(mai_mai_n411_), .B(mai_mai_n264_), .C(mai_mai_n70_), .Y(mai_mai_n840_));
  NO2        m818(.A(mai_mai_n169_), .B(mai_mai_n142_), .Y(mai_mai_n841_));
  AOI210     m819(.A0(mai_mai_n841_), .A1(mai_mai_n238_), .B0(mai_mai_n840_), .Y(mai_mai_n842_));
  OAI220     m820(.A0(mai_mai_n842_), .A1(mai_mai_n175_), .B0(mai_mai_n839_), .B1(mai_mai_n837_), .Y(mai_mai_n843_));
  NO4        m821(.A(mai_mai_n843_), .B(mai_mai_n835_), .C(mai_mai_n831_), .D(mai_mai_n825_), .Y(mai_mai_n844_));
  NA2        m822(.A(mai_mai_n179_), .B(mai_mai_n24_), .Y(mai_mai_n845_));
  NA2        m823(.A(mai_mai_n309_), .B(mai_mai_n124_), .Y(mai_mai_n846_));
  NAi21      m824(.An(mai_mai_n156_), .B(mai_mai_n438_), .Y(mai_mai_n847_));
  OAI220     m825(.A0(mai_mai_n847_), .A1(mai_mai_n813_), .B0(mai_mai_n846_), .B1(mai_mai_n396_), .Y(mai_mai_n848_));
  INV        m826(.A(mai_mai_n848_), .Y(mai_mai_n849_));
  NO4        m827(.A(mai_mai_n571_), .B(mai_mai_n208_), .C(mai_mai_n415_), .D(mai_mai_n407_), .Y(mai_mai_n850_));
  NA2        m828(.A(mai_mai_n729_), .B(mai_mai_n327_), .Y(mai_mai_n851_));
  AOI210     m829(.A0(mai_mai_n474_), .A1(mai_mai_n83_), .B0(mai_mai_n55_), .Y(mai_mai_n852_));
  OAI220     m830(.A0(mai_mai_n852_), .A1(mai_mai_n851_), .B0(mai_mai_n639_), .B1(mai_mai_n528_), .Y(mai_mai_n853_));
  NO2        m831(.A(mai_mai_n248_), .B(mai_mai_n147_), .Y(mai_mai_n854_));
  NA2        m832(.A(i_0_), .B(i_10_), .Y(mai_mai_n855_));
  AN2        m833(.A(mai_mai_n854_), .B(i_6_), .Y(mai_mai_n856_));
  AOI220     m834(.A0(mai_mai_n330_), .A1(mai_mai_n95_), .B0(mai_mai_n179_), .B1(mai_mai_n80_), .Y(mai_mai_n857_));
  NA2        m835(.A(mai_mai_n557_), .B(i_4_), .Y(mai_mai_n858_));
  NA2        m836(.A(mai_mai_n182_), .B(mai_mai_n197_), .Y(mai_mai_n859_));
  OAI220     m837(.A0(mai_mai_n859_), .A1(mai_mai_n851_), .B0(mai_mai_n858_), .B1(mai_mai_n857_), .Y(mai_mai_n860_));
  NO3        m838(.A(mai_mai_n860_), .B(mai_mai_n856_), .C(mai_mai_n853_), .Y(mai_mai_n861_));
  NA2        m839(.A(mai_mai_n861_), .B(mai_mai_n849_), .Y(mai_mai_n862_));
  NA2        m840(.A(mai_mai_n392_), .B(mai_mai_n173_), .Y(mai_mai_n863_));
  NA2        m841(.A(mai_mai_n863_), .B(mai_mai_n154_), .Y(mai_mai_n864_));
  NO2        m842(.A(mai_mai_n169_), .B(i_0_), .Y(mai_mai_n865_));
  INV        m843(.A(mai_mai_n865_), .Y(mai_mai_n866_));
  NA2        m844(.A(mai_mai_n465_), .B(mai_mai_n225_), .Y(mai_mai_n867_));
  INV        m845(.A(mai_mai_n404_), .Y(mai_mai_n868_));
  OAI220     m846(.A0(mai_mai_n868_), .A1(mai_mai_n837_), .B0(mai_mai_n867_), .B1(mai_mai_n866_), .Y(mai_mai_n869_));
  NO2        m847(.A(mai_mai_n869_), .B(mai_mai_n864_), .Y(mai_mai_n870_));
  NA2        m848(.A(mai_mai_n638_), .B(mai_mai_n116_), .Y(mai_mai_n871_));
  NO2        m849(.A(i_6_), .B(mai_mai_n871_), .Y(mai_mai_n872_));
  AOI210     m850(.A0(mai_mai_n448_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n873_));
  NA2        m851(.A(mai_mai_n165_), .B(mai_mai_n100_), .Y(mai_mai_n874_));
  NOi32      m852(.An(mai_mai_n873_), .Bn(mai_mai_n182_), .C(mai_mai_n874_), .Y(mai_mai_n875_));
  NO2        m853(.A(mai_mai_n875_), .B(mai_mai_n872_), .Y(mai_mai_n876_));
  NOi21      m854(.An(i_7_), .B(i_5_), .Y(mai_mai_n877_));
  NOi31      m855(.An(mai_mai_n877_), .B(i_0_), .C(mai_mai_n707_), .Y(mai_mai_n878_));
  NA3        m856(.A(mai_mai_n878_), .B(mai_mai_n382_), .C(i_6_), .Y(mai_mai_n879_));
  OA210      m857(.A0(mai_mai_n874_), .A1(mai_mai_n507_), .B0(mai_mai_n879_), .Y(mai_mai_n880_));
  NO3        m858(.A(mai_mai_n399_), .B(mai_mai_n363_), .C(mai_mai_n359_), .Y(mai_mai_n881_));
  NO2        m859(.A(mai_mai_n258_), .B(mai_mai_n316_), .Y(mai_mai_n882_));
  NO2        m860(.A(mai_mai_n707_), .B(mai_mai_n253_), .Y(mai_mai_n883_));
  AOI210     m861(.A0(mai_mai_n883_), .A1(mai_mai_n882_), .B0(mai_mai_n881_), .Y(mai_mai_n884_));
  NA4        m862(.A(mai_mai_n884_), .B(mai_mai_n880_), .C(mai_mai_n876_), .D(mai_mai_n870_), .Y(mai_mai_n885_));
  NO2        m863(.A(mai_mai_n845_), .B(mai_mai_n234_), .Y(mai_mai_n886_));
  AN2        m864(.A(mai_mai_n329_), .B(mai_mai_n327_), .Y(mai_mai_n887_));
  AN2        m865(.A(mai_mai_n887_), .B(mai_mai_n841_), .Y(mai_mai_n888_));
  OAI210     m866(.A0(mai_mai_n888_), .A1(mai_mai_n886_), .B0(i_10_), .Y(mai_mai_n889_));
  OA210      m867(.A0(mai_mai_n465_), .A1(mai_mai_n217_), .B0(mai_mai_n464_), .Y(mai_mai_n890_));
  NA3        m868(.A(mai_mai_n464_), .B(mai_mai_n408_), .C(mai_mai_n45_), .Y(mai_mai_n891_));
  INV        m869(.A(mai_mai_n891_), .Y(mai_mai_n892_));
  INV        m870(.A(mai_mai_n181_), .Y(mai_mai_n893_));
  AOI220     m871(.A0(mai_mai_n893_), .A1(mai_mai_n465_), .B0(mai_mai_n892_), .B1(mai_mai_n70_), .Y(mai_mai_n894_));
  NO2        m872(.A(mai_mai_n72_), .B(mai_mai_n731_), .Y(mai_mai_n895_));
  INV        m873(.A(mai_mai_n895_), .Y(mai_mai_n896_));
  NO2        m874(.A(mai_mai_n896_), .B(mai_mai_n47_), .Y(mai_mai_n897_));
  NO2        m875(.A(mai_mai_n582_), .B(mai_mai_n102_), .Y(mai_mai_n898_));
  NA2        m876(.A(mai_mai_n898_), .B(i_0_), .Y(mai_mai_n899_));
  NO2        m877(.A(mai_mai_n899_), .B(mai_mai_n82_), .Y(mai_mai_n900_));
  NO3        m878(.A(mai_mai_n900_), .B(mai_mai_n897_), .C(mai_mai_n512_), .Y(mai_mai_n901_));
  NA3        m879(.A(mai_mai_n901_), .B(mai_mai_n894_), .C(mai_mai_n889_), .Y(mai_mai_n902_));
  NO3        m880(.A(mai_mai_n902_), .B(mai_mai_n885_), .C(mai_mai_n862_), .Y(mai_mai_n903_));
  NO2        m881(.A(i_0_), .B(mai_mai_n707_), .Y(mai_mai_n904_));
  NA2        m882(.A(mai_mai_n70_), .B(mai_mai_n44_), .Y(mai_mai_n905_));
  NA2        m883(.A(mai_mai_n855_), .B(mai_mai_n905_), .Y(mai_mai_n906_));
  NO3        m884(.A(mai_mai_n102_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n907_));
  AO220      m885(.A0(mai_mai_n907_), .A1(mai_mai_n906_), .B0(mai_mai_n904_), .B1(mai_mai_n168_), .Y(mai_mai_n908_));
  AOI210     m886(.A0(mai_mai_n778_), .A1(mai_mai_n669_), .B0(mai_mai_n874_), .Y(mai_mai_n909_));
  AOI210     m887(.A0(mai_mai_n908_), .A1(mai_mai_n347_), .B0(mai_mai_n909_), .Y(mai_mai_n910_));
  NO2        m888(.A(mai_mai_n792_), .B(mai_mai_n399_), .Y(mai_mai_n911_));
  NA3        m889(.A(mai_mai_n820_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n912_));
  NA2        m890(.A(mai_mai_n821_), .B(i_9_), .Y(mai_mai_n913_));
  AOI210     m891(.A0(mai_mai_n912_), .A1(mai_mai_n488_), .B0(mai_mai_n913_), .Y(mai_mai_n914_));
  NA2        m892(.A(mai_mai_n238_), .B(mai_mai_n224_), .Y(mai_mai_n915_));
  NO2        m893(.A(mai_mai_n915_), .B(mai_mai_n147_), .Y(mai_mai_n916_));
  NO3        m894(.A(mai_mai_n916_), .B(mai_mai_n914_), .C(mai_mai_n911_), .Y(mai_mai_n917_));
  NA2        m895(.A(mai_mai_n917_), .B(mai_mai_n910_), .Y(mai_mai_n918_));
  NA2        m896(.A(mai_mai_n887_), .B(mai_mai_n371_), .Y(mai_mai_n919_));
  AOI210     m897(.A0(mai_mai_n297_), .A1(mai_mai_n156_), .B0(mai_mai_n919_), .Y(mai_mai_n920_));
  NA3        m898(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n44_), .Y(mai_mai_n921_));
  NA2        m899(.A(i_5_), .B(mai_mai_n478_), .Y(mai_mai_n922_));
  AOI210     m900(.A0(mai_mai_n921_), .A1(mai_mai_n156_), .B0(mai_mai_n922_), .Y(mai_mai_n923_));
  NO2        m901(.A(mai_mai_n923_), .B(mai_mai_n920_), .Y(mai_mai_n924_));
  NO3        m902(.A(mai_mai_n855_), .B(mai_mai_n836_), .C(mai_mai_n184_), .Y(mai_mai_n925_));
  AOI220     m903(.A0(mai_mai_n925_), .A1(i_11_), .B0(mai_mai_n558_), .B1(mai_mai_n72_), .Y(mai_mai_n926_));
  NO3        m904(.A(mai_mai_n202_), .B(mai_mai_n381_), .C(i_0_), .Y(mai_mai_n927_));
  OAI210     m905(.A0(mai_mai_n927_), .A1(mai_mai_n73_), .B0(i_13_), .Y(mai_mai_n928_));
  INV        m906(.A(mai_mai_n211_), .Y(mai_mai_n929_));
  OAI220     m907(.A0(mai_mai_n521_), .A1(mai_mai_n133_), .B0(mai_mai_n622_), .B1(mai_mai_n599_), .Y(mai_mai_n930_));
  NA3        m908(.A(mai_mai_n930_), .B(i_7_), .C(mai_mai_n929_), .Y(mai_mai_n931_));
  NA4        m909(.A(mai_mai_n931_), .B(mai_mai_n928_), .C(mai_mai_n926_), .D(mai_mai_n924_), .Y(mai_mai_n932_));
  NA2        m910(.A(mai_mai_n350_), .B(mai_mai_n170_), .Y(mai_mai_n933_));
  OR2        m911(.A(mai_mai_n933_), .B(mai_mai_n1000_), .Y(mai_mai_n934_));
  AOI210     m912(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n169_), .Y(mai_mai_n935_));
  NA2        m913(.A(mai_mai_n935_), .B(mai_mai_n890_), .Y(mai_mai_n936_));
  NA3        m914(.A(mai_mai_n388_), .B(mai_mai_n331_), .C(mai_mai_n215_), .Y(mai_mai_n937_));
  INV        m915(.A(mai_mai_n937_), .Y(mai_mai_n938_));
  NOi31      m916(.An(mai_mai_n387_), .B(mai_mai_n905_), .C(mai_mai_n234_), .Y(mai_mai_n939_));
  NO2        m917(.A(mai_mai_n939_), .B(mai_mai_n938_), .Y(mai_mai_n940_));
  NA3        m918(.A(mai_mai_n940_), .B(mai_mai_n936_), .C(mai_mai_n934_), .Y(mai_mai_n941_));
  NA3        m919(.A(mai_mai_n302_), .B(i_5_), .C(mai_mai_n187_), .Y(mai_mai_n942_));
  NAi31      m920(.An(mai_mai_n236_), .B(mai_mai_n942_), .C(mai_mai_n237_), .Y(mai_mai_n943_));
  NO4        m921(.A(mai_mai_n234_), .B(mai_mai_n202_), .C(i_0_), .D(i_12_), .Y(mai_mai_n944_));
  NA2        m922(.A(mai_mai_n944_), .B(mai_mai_n943_), .Y(mai_mai_n945_));
  AN2        m923(.A(mai_mai_n855_), .B(mai_mai_n147_), .Y(mai_mai_n946_));
  NO4        m924(.A(mai_mai_n946_), .B(i_12_), .C(mai_mai_n626_), .D(mai_mai_n126_), .Y(mai_mai_n947_));
  NA2        m925(.A(mai_mai_n947_), .B(mai_mai_n211_), .Y(mai_mai_n948_));
  NA3        m926(.A(mai_mai_n95_), .B(mai_mai_n562_), .C(i_11_), .Y(mai_mai_n949_));
  NA2        m927(.A(mai_mai_n877_), .B(mai_mai_n462_), .Y(mai_mai_n950_));
  NA2        m928(.A(mai_mai_n61_), .B(mai_mai_n98_), .Y(mai_mai_n951_));
  OAI220     m929(.A0(mai_mai_n951_), .A1(mai_mai_n942_), .B0(mai_mai_n950_), .B1(mai_mai_n657_), .Y(mai_mai_n952_));
  NA2        m930(.A(mai_mai_n952_), .B(mai_mai_n865_), .Y(mai_mai_n953_));
  NA3        m931(.A(mai_mai_n953_), .B(mai_mai_n948_), .C(mai_mai_n945_), .Y(mai_mai_n954_));
  NO4        m932(.A(mai_mai_n954_), .B(mai_mai_n941_), .C(mai_mai_n932_), .D(mai_mai_n918_), .Y(mai_mai_n955_));
  OAI210     m933(.A0(mai_mai_n795_), .A1(mai_mai_n788_), .B0(mai_mai_n37_), .Y(mai_mai_n956_));
  NA3        m934(.A(mai_mai_n873_), .B(mai_mai_n366_), .C(i_5_), .Y(mai_mai_n957_));
  NA3        m935(.A(mai_mai_n957_), .B(mai_mai_n956_), .C(mai_mai_n594_), .Y(mai_mai_n958_));
  NA2        m936(.A(mai_mai_n958_), .B(mai_mai_n199_), .Y(mai_mai_n959_));
  BUFFER     m937(.A(mai_mai_n367_), .Y(mai_mai_n960_));
  NA2        m938(.A(mai_mai_n180_), .B(mai_mai_n182_), .Y(mai_mai_n961_));
  AO210      m939(.A0(mai_mai_n960_), .A1(mai_mai_n33_), .B0(mai_mai_n961_), .Y(mai_mai_n962_));
  OAI210     m940(.A0(mai_mai_n598_), .A1(mai_mai_n596_), .B0(mai_mai_n315_), .Y(mai_mai_n963_));
  NAi31      m941(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n964_));
  AOI210     m942(.A0(mai_mai_n112_), .A1(mai_mai_n67_), .B0(mai_mai_n964_), .Y(mai_mai_n965_));
  NO2        m943(.A(mai_mai_n965_), .B(mai_mai_n623_), .Y(mai_mai_n966_));
  NA3        m944(.A(mai_mai_n966_), .B(mai_mai_n963_), .C(mai_mai_n962_), .Y(mai_mai_n967_));
  NO2        m945(.A(mai_mai_n456_), .B(mai_mai_n264_), .Y(mai_mai_n968_));
  NO4        m946(.A(mai_mai_n227_), .B(mai_mai_n139_), .C(mai_mai_n660_), .D(mai_mai_n37_), .Y(mai_mai_n969_));
  NO3        m947(.A(mai_mai_n969_), .B(mai_mai_n968_), .C(mai_mai_n850_), .Y(mai_mai_n970_));
  OAI210     m948(.A0(mai_mai_n949_), .A1(mai_mai_n142_), .B0(mai_mai_n970_), .Y(mai_mai_n971_));
  AOI210     m949(.A0(mai_mai_n967_), .A1(mai_mai_n48_), .B0(mai_mai_n971_), .Y(mai_mai_n972_));
  AOI210     m950(.A0(mai_mai_n972_), .A1(mai_mai_n959_), .B0(mai_mai_n70_), .Y(mai_mai_n973_));
  NO2        m951(.A(mai_mai_n555_), .B(mai_mai_n377_), .Y(mai_mai_n974_));
  NO2        m952(.A(mai_mai_n974_), .B(mai_mai_n737_), .Y(mai_mai_n975_));
  INV        m953(.A(mai_mai_n73_), .Y(mai_mai_n976_));
  AOI210     m954(.A0(mai_mai_n935_), .A1(i_5_), .B0(mai_mai_n878_), .Y(mai_mai_n977_));
  AOI210     m955(.A0(mai_mai_n977_), .A1(mai_mai_n976_), .B0(mai_mai_n660_), .Y(mai_mai_n978_));
  NA2        m956(.A(mai_mai_n258_), .B(mai_mai_n54_), .Y(mai_mai_n979_));
  AOI220     m957(.A0(mai_mai_n979_), .A1(mai_mai_n73_), .B0(mai_mai_n345_), .B1(mai_mai_n250_), .Y(mai_mai_n980_));
  NO2        m958(.A(mai_mai_n980_), .B(mai_mai_n231_), .Y(mai_mai_n981_));
  NA3        m959(.A(mai_mai_n93_), .B(mai_mai_n304_), .C(mai_mai_n31_), .Y(mai_mai_n982_));
  INV        m960(.A(mai_mai_n982_), .Y(mai_mai_n983_));
  NO3        m961(.A(mai_mai_n983_), .B(mai_mai_n981_), .C(mai_mai_n978_), .Y(mai_mai_n984_));
  OAI210     m962(.A0(mai_mai_n266_), .A1(mai_mai_n152_), .B0(mai_mai_n83_), .Y(mai_mai_n985_));
  NO2        m963(.A(mai_mai_n985_), .B(i_11_), .Y(mai_mai_n986_));
  OAI210     m964(.A0(mai_mai_n998_), .A1(mai_mai_n873_), .B0(mai_mai_n199_), .Y(mai_mai_n987_));
  NA2        m965(.A(mai_mai_n158_), .B(i_5_), .Y(mai_mai_n988_));
  NO2        m966(.A(mai_mai_n987_), .B(mai_mai_n988_), .Y(mai_mai_n989_));
  NO2        m967(.A(mai_mai_n989_), .B(mai_mai_n986_), .Y(mai_mai_n990_));
  OAI210     m968(.A0(mai_mai_n984_), .A1(i_4_), .B0(mai_mai_n990_), .Y(mai_mai_n991_));
  NO3        m969(.A(mai_mai_n991_), .B(mai_mai_n975_), .C(mai_mai_n973_), .Y(mai_mai_n992_));
  NA4        m970(.A(mai_mai_n992_), .B(mai_mai_n955_), .C(mai_mai_n903_), .D(mai_mai_n844_), .Y(mai4));
  INV        m971(.A(i_2_), .Y(mai_mai_n996_));
  INV        m972(.A(i_12_), .Y(mai_mai_n997_));
  INV        m973(.A(i_12_), .Y(mai_mai_n998_));
  INV        m974(.A(mai_mai_n832_), .Y(mai_mai_n999_));
  INV        m975(.A(mai_mai_n157_), .Y(mai_mai_n1000_));
  INV        m976(.A(i_1_), .Y(mai_mai_n1001_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n51_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(men_men_n81_), .B(men_men_n58_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_9_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_7_), .Y(men_men_n84_));
  INV        u0062(.A(i_6_), .Y(men_men_n85_));
  OR4        u0063(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n86_));
  INV        u0064(.A(men_men_n86_), .Y(men_men_n87_));
  NO2        u0065(.A(i_2_), .B(i_7_), .Y(men_men_n88_));
  NAi21      u0066(.An(i_6_), .B(i_10_), .Y(men_men_n89_));
  NA2        u0067(.A(i_6_), .B(i_9_), .Y(men_men_n90_));
  AOI210     u0068(.A0(men_men_n90_), .A1(men_men_n89_), .B0(men_men_n63_), .Y(men_men_n91_));
  NA2        u0069(.A(i_2_), .B(i_6_), .Y(men_men_n92_));
  INV        u0070(.A(men_men_n91_), .Y(men_men_n93_));
  AOI210     u0071(.A0(men_men_n93_), .A1(men_men_n1078_), .B0(men_men_n80_), .Y(men_men_n94_));
  AN3        u0072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n95_));
  NAi21      u0073(.An(i_6_), .B(i_11_), .Y(men_men_n96_));
  NO2        u0074(.A(i_5_), .B(i_8_), .Y(men_men_n97_));
  NOi21      u0075(.An(men_men_n97_), .B(men_men_n96_), .Y(men_men_n98_));
  AOI220     u0076(.A0(men_men_n98_), .A1(men_men_n62_), .B0(men_men_n95_), .B1(men_men_n32_), .Y(men_men_n99_));
  INV        u0077(.A(i_7_), .Y(men_men_n100_));
  NA2        u0078(.A(men_men_n47_), .B(men_men_n100_), .Y(men_men_n101_));
  NO2        u0079(.A(i_0_), .B(i_5_), .Y(men_men_n102_));
  NO2        u0080(.A(men_men_n102_), .B(men_men_n85_), .Y(men_men_n103_));
  NA2        u0081(.A(i_12_), .B(i_3_), .Y(men_men_n104_));
  INV        u0082(.A(men_men_n104_), .Y(men_men_n105_));
  NA3        u0083(.A(men_men_n105_), .B(men_men_n103_), .C(men_men_n101_), .Y(men_men_n106_));
  NAi21      u0084(.An(i_7_), .B(i_11_), .Y(men_men_n107_));
  NO3        u0085(.A(men_men_n107_), .B(men_men_n89_), .C(men_men_n54_), .Y(men_men_n108_));
  AN2        u0086(.A(i_2_), .B(i_10_), .Y(men_men_n109_));
  NO2        u0087(.A(men_men_n109_), .B(i_7_), .Y(men_men_n110_));
  OR2        u0088(.A(men_men_n80_), .B(men_men_n58_), .Y(men_men_n111_));
  NO2        u0089(.A(i_8_), .B(men_men_n100_), .Y(men_men_n112_));
  NO3        u0090(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n110_), .Y(men_men_n113_));
  NA2        u0091(.A(i_12_), .B(i_7_), .Y(men_men_n114_));
  NO2        u0092(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n115_));
  NA2        u0093(.A(men_men_n115_), .B(i_0_), .Y(men_men_n116_));
  NA2        u0094(.A(i_11_), .B(i_12_), .Y(men_men_n117_));
  OAI210     u0095(.A0(men_men_n116_), .A1(men_men_n114_), .B0(men_men_n117_), .Y(men_men_n118_));
  NO2        u0096(.A(men_men_n118_), .B(men_men_n113_), .Y(men_men_n119_));
  NAi41      u0097(.An(men_men_n108_), .B(men_men_n119_), .C(men_men_n106_), .D(men_men_n99_), .Y(men_men_n120_));
  NOi21      u0098(.An(i_1_), .B(i_5_), .Y(men_men_n121_));
  NA2        u0099(.A(men_men_n121_), .B(i_11_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n100_), .B(men_men_n37_), .Y(men_men_n123_));
  NA2        u0101(.A(i_7_), .B(men_men_n25_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NO2        u0103(.A(men_men_n125_), .B(men_men_n47_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n127_));
  NAi21      u0105(.An(i_3_), .B(i_8_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n128_), .B(men_men_n62_), .Y(men_men_n129_));
  NOi31      u0107(.An(men_men_n129_), .B(men_men_n127_), .C(men_men_n126_), .Y(men_men_n130_));
  NO2        u0108(.A(i_1_), .B(men_men_n85_), .Y(men_men_n131_));
  NO2        u0109(.A(i_6_), .B(i_5_), .Y(men_men_n132_));
  NA2        u0110(.A(men_men_n132_), .B(i_3_), .Y(men_men_n133_));
  AO210      u0111(.A0(men_men_n133_), .A1(men_men_n48_), .B0(men_men_n131_), .Y(men_men_n134_));
  OAI220     u0112(.A0(men_men_n134_), .A1(men_men_n107_), .B0(men_men_n130_), .B1(men_men_n122_), .Y(men_men_n135_));
  NO3        u0113(.A(men_men_n135_), .B(men_men_n120_), .C(men_men_n94_), .Y(men_men_n136_));
  NA3        u0114(.A(men_men_n136_), .B(men_men_n79_), .C(men_men_n56_), .Y(men2));
  NO2        u0115(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n138_));
  NA2        u0116(.A(i_6_), .B(men_men_n25_), .Y(men_men_n139_));
  NA2        u0117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NA4        u0118(.A(men_men_n140_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n30_), .Y(men0));
  AN2        u0119(.A(i_8_), .B(i_7_), .Y(men_men_n142_));
  NA2        u0120(.A(men_men_n142_), .B(i_6_), .Y(men_men_n143_));
  NO2        u0121(.A(i_12_), .B(i_13_), .Y(men_men_n144_));
  NAi21      u0122(.An(i_5_), .B(i_11_), .Y(men_men_n145_));
  NOi21      u0123(.An(men_men_n144_), .B(men_men_n145_), .Y(men_men_n146_));
  NO2        u0124(.A(i_0_), .B(i_1_), .Y(men_men_n147_));
  NA2        u0125(.A(i_2_), .B(i_3_), .Y(men_men_n148_));
  NA3        u0126(.A(i_3_), .B(men_men_n147_), .C(men_men_n146_), .Y(men_men_n149_));
  OR2        u0127(.A(men_men_n149_), .B(men_men_n25_), .Y(men_men_n150_));
  AN2        u0128(.A(men_men_n144_), .B(men_men_n83_), .Y(men_men_n151_));
  NO2        u0129(.A(men_men_n151_), .B(men_men_n27_), .Y(men_men_n152_));
  NA2        u0130(.A(i_1_), .B(i_5_), .Y(men_men_n153_));
  NO2        u0131(.A(men_men_n73_), .B(men_men_n47_), .Y(men_men_n154_));
  NA2        u0132(.A(men_men_n154_), .B(men_men_n36_), .Y(men_men_n155_));
  NO3        u0133(.A(men_men_n155_), .B(men_men_n153_), .C(men_men_n152_), .Y(men_men_n156_));
  OR2        u0134(.A(i_0_), .B(i_1_), .Y(men_men_n157_));
  NO3        u0135(.A(men_men_n157_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n158_));
  NAi32      u0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n159_));
  NAi21      u0137(.An(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  NOi21      u0138(.An(i_4_), .B(i_10_), .Y(men_men_n161_));
  NA2        u0139(.A(men_men_n161_), .B(men_men_n40_), .Y(men_men_n162_));
  NO2        u0140(.A(i_3_), .B(i_5_), .Y(men_men_n163_));
  NO3        u0141(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n164_));
  NA2        u0142(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  OAI210     u0143(.A0(men_men_n165_), .A1(men_men_n162_), .B0(men_men_n160_), .Y(men_men_n166_));
  NO2        u0144(.A(men_men_n166_), .B(men_men_n156_), .Y(men_men_n167_));
  AOI210     u0145(.A0(men_men_n167_), .A1(men_men_n150_), .B0(men_men_n143_), .Y(men_men_n168_));
  NA3        u0146(.A(men_men_n73_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n169_));
  NOi21      u0147(.An(i_4_), .B(i_9_), .Y(men_men_n170_));
  NOi21      u0148(.An(i_11_), .B(i_13_), .Y(men_men_n171_));
  NA2        u0149(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  NO2        u0150(.A(i_4_), .B(i_5_), .Y(men_men_n173_));
  NAi21      u0151(.An(i_12_), .B(i_11_), .Y(men_men_n174_));
  NO2        u0152(.A(men_men_n174_), .B(i_13_), .Y(men_men_n175_));
  NA3        u0153(.A(men_men_n175_), .B(men_men_n173_), .C(men_men_n83_), .Y(men_men_n176_));
  AOI210     u0154(.A0(men_men_n176_), .A1(men_men_n172_), .B0(men_men_n169_), .Y(men_men_n177_));
  NO2        u0155(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n178_));
  NA2        u0156(.A(men_men_n178_), .B(men_men_n47_), .Y(men_men_n179_));
  NA2        u0157(.A(men_men_n36_), .B(i_5_), .Y(men_men_n180_));
  NAi31      u0158(.An(men_men_n180_), .B(men_men_n151_), .C(i_11_), .Y(men_men_n181_));
  NA2        u0159(.A(i_3_), .B(i_5_), .Y(men_men_n182_));
  OR2        u0160(.A(men_men_n182_), .B(men_men_n172_), .Y(men_men_n183_));
  AOI210     u0161(.A0(men_men_n183_), .A1(men_men_n181_), .B0(men_men_n179_), .Y(men_men_n184_));
  NO2        u0162(.A(men_men_n73_), .B(i_5_), .Y(men_men_n185_));
  NO2        u0163(.A(i_13_), .B(i_10_), .Y(men_men_n186_));
  NA3        u0164(.A(men_men_n186_), .B(men_men_n185_), .C(men_men_n45_), .Y(men_men_n187_));
  NO2        u0165(.A(i_2_), .B(i_1_), .Y(men_men_n188_));
  NA2        u0166(.A(men_men_n188_), .B(i_3_), .Y(men_men_n189_));
  NAi21      u0167(.An(i_4_), .B(i_12_), .Y(men_men_n190_));
  NO4        u0168(.A(men_men_n190_), .B(men_men_n189_), .C(men_men_n187_), .D(men_men_n25_), .Y(men_men_n191_));
  NO3        u0169(.A(men_men_n191_), .B(men_men_n184_), .C(men_men_n177_), .Y(men_men_n192_));
  INV        u0170(.A(i_8_), .Y(men_men_n193_));
  NO2        u0171(.A(men_men_n193_), .B(i_7_), .Y(men_men_n194_));
  NA2        u0172(.A(men_men_n194_), .B(i_6_), .Y(men_men_n195_));
  NO3        u0173(.A(i_3_), .B(men_men_n85_), .C(men_men_n49_), .Y(men_men_n196_));
  NA2        u0174(.A(men_men_n196_), .B(men_men_n112_), .Y(men_men_n197_));
  NO3        u0175(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n198_));
  NA3        u0176(.A(men_men_n198_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n199_));
  NO3        u0177(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n200_));
  OAI210     u0178(.A0(men_men_n95_), .A1(i_12_), .B0(men_men_n200_), .Y(men_men_n201_));
  AOI210     u0179(.A0(men_men_n201_), .A1(men_men_n199_), .B0(men_men_n197_), .Y(men_men_n202_));
  NO2        u0180(.A(i_3_), .B(i_8_), .Y(men_men_n203_));
  NO3        u0181(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n204_));
  NA3        u0182(.A(men_men_n204_), .B(men_men_n203_), .C(men_men_n40_), .Y(men_men_n205_));
  NO2        u0183(.A(men_men_n102_), .B(men_men_n58_), .Y(men_men_n206_));
  NO2        u0184(.A(i_13_), .B(i_9_), .Y(men_men_n207_));
  NA3        u0185(.A(men_men_n207_), .B(i_6_), .C(men_men_n193_), .Y(men_men_n208_));
  NAi21      u0186(.An(i_12_), .B(i_3_), .Y(men_men_n209_));
  OR2        u0187(.A(men_men_n209_), .B(men_men_n208_), .Y(men_men_n210_));
  NO2        u0188(.A(men_men_n45_), .B(i_5_), .Y(men_men_n211_));
  NO3        u0189(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n212_));
  INV        u0190(.A(men_men_n212_), .Y(men_men_n213_));
  OAI220     u0191(.A0(men_men_n213_), .A1(men_men_n210_), .B0(men_men_n102_), .B1(men_men_n205_), .Y(men_men_n214_));
  AOI210     u0192(.A0(men_men_n214_), .A1(i_7_), .B0(men_men_n202_), .Y(men_men_n215_));
  OAI220     u0193(.A0(men_men_n215_), .A1(i_4_), .B0(men_men_n195_), .B1(men_men_n192_), .Y(men_men_n216_));
  NAi21      u0194(.An(i_12_), .B(i_7_), .Y(men_men_n217_));
  NA3        u0195(.A(i_13_), .B(men_men_n193_), .C(i_10_), .Y(men_men_n218_));
  NO2        u0196(.A(men_men_n218_), .B(men_men_n217_), .Y(men_men_n219_));
  NA2        u0197(.A(i_0_), .B(i_5_), .Y(men_men_n220_));
  OAI220     u0198(.A0(men_men_n85_), .A1(men_men_n189_), .B0(men_men_n179_), .B1(men_men_n133_), .Y(men_men_n221_));
  NAi31      u0199(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n36_), .B(i_13_), .Y(men_men_n223_));
  NO2        u0201(.A(men_men_n47_), .B(men_men_n63_), .Y(men_men_n224_));
  NA3        u0202(.A(men_men_n224_), .B(i_0_), .C(men_men_n223_), .Y(men_men_n225_));
  INV        u0203(.A(i_13_), .Y(men_men_n226_));
  NO2        u0204(.A(i_12_), .B(men_men_n226_), .Y(men_men_n227_));
  NA3        u0205(.A(men_men_n227_), .B(men_men_n198_), .C(men_men_n196_), .Y(men_men_n228_));
  OAI210     u0206(.A0(men_men_n225_), .A1(men_men_n222_), .B0(men_men_n228_), .Y(men_men_n229_));
  AOI220     u0207(.A0(men_men_n229_), .A1(men_men_n142_), .B0(men_men_n221_), .B1(men_men_n219_), .Y(men_men_n230_));
  NO2        u0208(.A(i_12_), .B(men_men_n37_), .Y(men_men_n231_));
  NO2        u0209(.A(men_men_n182_), .B(i_4_), .Y(men_men_n232_));
  NA2        u0210(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n233_));
  OR2        u0211(.A(i_8_), .B(i_7_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n234_), .B(men_men_n85_), .Y(men_men_n235_));
  NO2        u0213(.A(men_men_n54_), .B(i_1_), .Y(men_men_n236_));
  NA2        u0214(.A(men_men_n236_), .B(men_men_n235_), .Y(men_men_n237_));
  INV        u0215(.A(i_12_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n45_), .B(men_men_n238_), .Y(men_men_n239_));
  NO3        u0217(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n240_));
  NA2        u0218(.A(i_2_), .B(i_1_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n237_), .B(men_men_n233_), .Y(men_men_n242_));
  NO3        u0220(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n243_));
  NAi21      u0221(.An(i_4_), .B(i_3_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n244_), .B(men_men_n75_), .Y(men_men_n245_));
  NO2        u0223(.A(i_0_), .B(i_6_), .Y(men_men_n246_));
  NOi41      u0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n247_));
  NA2        u0225(.A(men_men_n247_), .B(men_men_n246_), .Y(men_men_n248_));
  NO2        u0226(.A(men_men_n241_), .B(men_men_n182_), .Y(men_men_n249_));
  NAi21      u0227(.An(men_men_n248_), .B(men_men_n249_), .Y(men_men_n250_));
  INV        u0228(.A(men_men_n250_), .Y(men_men_n251_));
  AOI220     u0229(.A0(men_men_n251_), .A1(men_men_n40_), .B0(men_men_n242_), .B1(men_men_n207_), .Y(men_men_n252_));
  NO2        u0230(.A(i_11_), .B(men_men_n226_), .Y(men_men_n253_));
  NOi21      u0231(.An(i_1_), .B(i_6_), .Y(men_men_n254_));
  NAi21      u0232(.An(i_3_), .B(i_7_), .Y(men_men_n255_));
  NO2        u0233(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n256_));
  NO2        u0234(.A(i_12_), .B(i_3_), .Y(men_men_n257_));
  NA2        u0235(.A(i_3_), .B(i_9_), .Y(men_men_n258_));
  NA3        u0236(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n259_));
  INV        u0237(.A(men_men_n143_), .Y(men_men_n260_));
  NA2        u0238(.A(men_men_n238_), .B(i_13_), .Y(men_men_n261_));
  NO2        u0239(.A(men_men_n261_), .B(men_men_n75_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n262_), .B(men_men_n260_), .Y(men_men_n263_));
  NO2        u0241(.A(men_men_n234_), .B(men_men_n37_), .Y(men_men_n264_));
  NA2        u0242(.A(i_12_), .B(i_6_), .Y(men_men_n265_));
  OR2        u0243(.A(i_13_), .B(i_9_), .Y(men_men_n266_));
  NO3        u0244(.A(men_men_n266_), .B(men_men_n265_), .C(men_men_n49_), .Y(men_men_n267_));
  NO2        u0245(.A(men_men_n244_), .B(i_2_), .Y(men_men_n268_));
  NA3        u0246(.A(men_men_n268_), .B(men_men_n267_), .C(men_men_n45_), .Y(men_men_n269_));
  NA2        u0247(.A(men_men_n253_), .B(i_9_), .Y(men_men_n270_));
  NA2        u0248(.A(i_0_), .B(men_men_n64_), .Y(men_men_n271_));
  OAI210     u0249(.A0(men_men_n271_), .A1(men_men_n270_), .B0(men_men_n269_), .Y(men_men_n272_));
  NA2        u0250(.A(men_men_n154_), .B(men_men_n63_), .Y(men_men_n273_));
  NO3        u0251(.A(i_11_), .B(men_men_n226_), .C(men_men_n25_), .Y(men_men_n274_));
  NO2        u0252(.A(men_men_n255_), .B(i_8_), .Y(men_men_n275_));
  NO2        u0253(.A(i_6_), .B(men_men_n49_), .Y(men_men_n276_));
  NA3        u0254(.A(men_men_n276_), .B(men_men_n275_), .C(men_men_n274_), .Y(men_men_n277_));
  NO3        u0255(.A(men_men_n26_), .B(men_men_n85_), .C(i_5_), .Y(men_men_n278_));
  NA3        u0256(.A(men_men_n278_), .B(men_men_n264_), .C(men_men_n227_), .Y(men_men_n279_));
  AOI210     u0257(.A0(men_men_n279_), .A1(men_men_n277_), .B0(men_men_n273_), .Y(men_men_n280_));
  AOI210     u0258(.A0(men_men_n272_), .A1(men_men_n264_), .B0(men_men_n280_), .Y(men_men_n281_));
  NA4        u0259(.A(men_men_n281_), .B(men_men_n263_), .C(men_men_n252_), .D(men_men_n230_), .Y(men_men_n282_));
  NO3        u0260(.A(i_12_), .B(men_men_n226_), .C(men_men_n37_), .Y(men_men_n283_));
  INV        u0261(.A(men_men_n283_), .Y(men_men_n284_));
  NA2        u0262(.A(i_8_), .B(men_men_n100_), .Y(men_men_n285_));
  NO3        u0263(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n286_));
  AOI220     u0264(.A0(men_men_n286_), .A1(men_men_n196_), .B0(men_men_n163_), .B1(men_men_n236_), .Y(men_men_n287_));
  NO2        u0265(.A(men_men_n287_), .B(men_men_n285_), .Y(men_men_n288_));
  NO3        u0266(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n289_));
  NO2        u0267(.A(men_men_n241_), .B(i_0_), .Y(men_men_n290_));
  AOI220     u0268(.A0(men_men_n290_), .A1(men_men_n194_), .B0(men_men_n289_), .B1(men_men_n142_), .Y(men_men_n291_));
  NA2        u0269(.A(men_men_n276_), .B(men_men_n26_), .Y(men_men_n292_));
  NO2        u0270(.A(men_men_n292_), .B(men_men_n291_), .Y(men_men_n293_));
  NA2        u0271(.A(i_0_), .B(i_1_), .Y(men_men_n294_));
  NO2        u0272(.A(men_men_n294_), .B(i_2_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n59_), .B(i_6_), .Y(men_men_n296_));
  NA3        u0274(.A(men_men_n296_), .B(men_men_n295_), .C(men_men_n163_), .Y(men_men_n297_));
  OAI210     u0275(.A0(men_men_n165_), .A1(men_men_n143_), .B0(men_men_n297_), .Y(men_men_n298_));
  NO3        u0276(.A(men_men_n298_), .B(men_men_n293_), .C(men_men_n288_), .Y(men_men_n299_));
  NO2        u0277(.A(i_3_), .B(i_10_), .Y(men_men_n300_));
  NA3        u0278(.A(men_men_n300_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n301_));
  NO2        u0279(.A(i_2_), .B(men_men_n100_), .Y(men_men_n302_));
  NA2        u0280(.A(i_1_), .B(men_men_n36_), .Y(men_men_n303_));
  NOi21      u0281(.An(men_men_n220_), .B(men_men_n102_), .Y(men_men_n304_));
  NA3        u0282(.A(men_men_n304_), .B(i_1_), .C(men_men_n302_), .Y(men_men_n305_));
  AN2        u0283(.A(i_3_), .B(i_10_), .Y(men_men_n306_));
  NA4        u0284(.A(men_men_n306_), .B(men_men_n198_), .C(men_men_n175_), .D(men_men_n173_), .Y(men_men_n307_));
  NO2        u0285(.A(i_5_), .B(men_men_n37_), .Y(men_men_n308_));
  NO2        u0286(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n309_));
  OR2        u0287(.A(men_men_n305_), .B(men_men_n301_), .Y(men_men_n310_));
  OAI220     u0288(.A0(men_men_n310_), .A1(i_6_), .B0(men_men_n299_), .B1(men_men_n284_), .Y(men_men_n311_));
  NO4        u0289(.A(men_men_n311_), .B(men_men_n282_), .C(men_men_n216_), .D(men_men_n168_), .Y(men_men_n312_));
  NO3        u0290(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n313_));
  NO2        u0291(.A(men_men_n59_), .B(men_men_n85_), .Y(men_men_n314_));
  NA2        u0292(.A(men_men_n290_), .B(men_men_n314_), .Y(men_men_n315_));
  NO3        u0293(.A(i_6_), .B(men_men_n193_), .C(i_7_), .Y(men_men_n316_));
  NA2        u0294(.A(men_men_n316_), .B(men_men_n198_), .Y(men_men_n317_));
  AOI210     u0295(.A0(men_men_n317_), .A1(men_men_n315_), .B0(i_5_), .Y(men_men_n318_));
  NO2        u0296(.A(i_2_), .B(i_3_), .Y(men_men_n319_));
  OR2        u0297(.A(i_0_), .B(i_5_), .Y(men_men_n320_));
  NA2        u0298(.A(men_men_n220_), .B(men_men_n320_), .Y(men_men_n321_));
  NA4        u0299(.A(men_men_n321_), .B(men_men_n235_), .C(men_men_n319_), .D(i_1_), .Y(men_men_n322_));
  NA3        u0300(.A(men_men_n290_), .B(men_men_n163_), .C(men_men_n112_), .Y(men_men_n323_));
  NO2        u0301(.A(i_8_), .B(i_6_), .Y(men_men_n324_));
  NO2        u0302(.A(men_men_n157_), .B(men_men_n47_), .Y(men_men_n325_));
  NA3        u0303(.A(men_men_n325_), .B(men_men_n324_), .C(men_men_n163_), .Y(men_men_n326_));
  NA3        u0304(.A(men_men_n326_), .B(men_men_n323_), .C(men_men_n322_), .Y(men_men_n327_));
  OAI210     u0305(.A0(men_men_n327_), .A1(men_men_n318_), .B0(i_4_), .Y(men_men_n328_));
  NO2        u0306(.A(i_12_), .B(i_10_), .Y(men_men_n329_));
  NOi21      u0307(.An(i_5_), .B(i_0_), .Y(men_men_n330_));
  NO3        u0308(.A(men_men_n303_), .B(men_men_n330_), .C(men_men_n128_), .Y(men_men_n331_));
  NA4        u0309(.A(men_men_n84_), .B(men_men_n36_), .C(men_men_n85_), .D(i_8_), .Y(men_men_n332_));
  NA2        u0310(.A(men_men_n331_), .B(men_men_n329_), .Y(men_men_n333_));
  NO2        u0311(.A(i_6_), .B(i_8_), .Y(men_men_n334_));
  NOi21      u0312(.An(i_0_), .B(i_2_), .Y(men_men_n335_));
  AN2        u0313(.A(men_men_n335_), .B(men_men_n334_), .Y(men_men_n336_));
  NO2        u0314(.A(i_1_), .B(i_7_), .Y(men_men_n337_));
  AO220      u0315(.A0(men_men_n337_), .A1(men_men_n336_), .B0(men_men_n324_), .B1(men_men_n236_), .Y(men_men_n338_));
  NA2        u0316(.A(men_men_n338_), .B(men_men_n42_), .Y(men_men_n339_));
  NA3        u0317(.A(men_men_n339_), .B(men_men_n333_), .C(men_men_n328_), .Y(men_men_n340_));
  NO3        u0318(.A(men_men_n234_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n341_));
  NO3        u0319(.A(i_8_), .B(i_2_), .C(i_1_), .Y(men_men_n342_));
  OAI210     u0320(.A0(men_men_n342_), .A1(men_men_n341_), .B0(i_6_), .Y(men_men_n343_));
  NA3        u0321(.A(men_men_n254_), .B(men_men_n302_), .C(men_men_n193_), .Y(men_men_n344_));
  AOI210     u0322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n321_), .Y(men_men_n345_));
  NA2        u0323(.A(men_men_n345_), .B(i_3_), .Y(men_men_n346_));
  INV        u0324(.A(men_men_n84_), .Y(men_men_n347_));
  NO2        u0325(.A(men_men_n294_), .B(men_men_n81_), .Y(men_men_n348_));
  NA2        u0326(.A(men_men_n348_), .B(men_men_n132_), .Y(men_men_n349_));
  NO2        u0327(.A(men_men_n92_), .B(men_men_n193_), .Y(men_men_n350_));
  NA3        u0328(.A(men_men_n304_), .B(men_men_n350_), .C(men_men_n63_), .Y(men_men_n351_));
  AOI210     u0329(.A0(men_men_n351_), .A1(men_men_n349_), .B0(men_men_n347_), .Y(men_men_n352_));
  NO2        u0330(.A(men_men_n193_), .B(i_9_), .Y(men_men_n353_));
  NA2        u0331(.A(men_men_n353_), .B(men_men_n206_), .Y(men_men_n354_));
  NO2        u0332(.A(men_men_n352_), .B(men_men_n293_), .Y(men_men_n355_));
  AOI210     u0333(.A0(men_men_n355_), .A1(men_men_n346_), .B0(men_men_n162_), .Y(men_men_n356_));
  AOI210     u0334(.A0(men_men_n340_), .A1(men_men_n313_), .B0(men_men_n356_), .Y(men_men_n357_));
  NOi32      u0335(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n358_));
  INV        u0336(.A(men_men_n358_), .Y(men_men_n359_));
  NAi21      u0337(.An(i_0_), .B(i_6_), .Y(men_men_n360_));
  NAi21      u0338(.An(i_1_), .B(i_5_), .Y(men_men_n361_));
  NA2        u0339(.A(men_men_n361_), .B(men_men_n360_), .Y(men_men_n362_));
  NAi41      u0340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n363_));
  OAI220     u0341(.A0(men_men_n363_), .A1(men_men_n361_), .B0(men_men_n222_), .B1(men_men_n159_), .Y(men_men_n364_));
  AOI210     u0342(.A0(men_men_n363_), .A1(men_men_n159_), .B0(men_men_n157_), .Y(men_men_n365_));
  NOi32      u0343(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n366_));
  NAi21      u0344(.An(i_6_), .B(i_1_), .Y(men_men_n367_));
  NA3        u0345(.A(men_men_n367_), .B(men_men_n366_), .C(men_men_n47_), .Y(men_men_n368_));
  NO2        u0346(.A(men_men_n368_), .B(i_0_), .Y(men_men_n369_));
  OR3        u0347(.A(men_men_n369_), .B(men_men_n365_), .C(men_men_n364_), .Y(men_men_n370_));
  NO2        u0348(.A(i_1_), .B(men_men_n100_), .Y(men_men_n371_));
  NAi21      u0349(.An(i_3_), .B(i_4_), .Y(men_men_n372_));
  NO2        u0350(.A(men_men_n372_), .B(i_9_), .Y(men_men_n373_));
  AN2        u0351(.A(i_6_), .B(i_7_), .Y(men_men_n374_));
  OAI210     u0352(.A0(men_men_n374_), .A1(men_men_n371_), .B0(men_men_n373_), .Y(men_men_n375_));
  NA2        u0353(.A(i_2_), .B(i_7_), .Y(men_men_n376_));
  NO2        u0354(.A(men_men_n372_), .B(i_10_), .Y(men_men_n377_));
  NA3        u0355(.A(men_men_n377_), .B(men_men_n376_), .C(men_men_n246_), .Y(men_men_n378_));
  AOI210     u0356(.A0(men_men_n378_), .A1(men_men_n375_), .B0(men_men_n185_), .Y(men_men_n379_));
  AOI210     u0357(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n380_));
  AOI220     u0358(.A0(men_men_n377_), .A1(men_men_n337_), .B0(men_men_n240_), .B1(men_men_n188_), .Y(men_men_n381_));
  NO2        u0359(.A(men_men_n381_), .B(i_5_), .Y(men_men_n382_));
  NO3        u0360(.A(men_men_n382_), .B(men_men_n379_), .C(men_men_n370_), .Y(men_men_n383_));
  NO2        u0361(.A(men_men_n383_), .B(men_men_n359_), .Y(men_men_n384_));
  NO2        u0362(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n385_));
  AN2        u0363(.A(i_12_), .B(i_5_), .Y(men_men_n386_));
  NO2        u0364(.A(i_4_), .B(men_men_n26_), .Y(men_men_n387_));
  NA2        u0365(.A(men_men_n387_), .B(men_men_n386_), .Y(men_men_n388_));
  NO2        u0366(.A(i_11_), .B(i_6_), .Y(men_men_n389_));
  NA3        u0367(.A(men_men_n389_), .B(men_men_n325_), .C(men_men_n226_), .Y(men_men_n390_));
  NO2        u0368(.A(men_men_n390_), .B(men_men_n388_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n244_), .B(i_5_), .Y(men_men_n392_));
  NO2        u0370(.A(i_5_), .B(i_10_), .Y(men_men_n393_));
  AOI220     u0371(.A0(men_men_n393_), .A1(men_men_n268_), .B0(men_men_n392_), .B1(men_men_n198_), .Y(men_men_n394_));
  NA2        u0372(.A(men_men_n144_), .B(men_men_n46_), .Y(men_men_n395_));
  NO2        u0373(.A(men_men_n395_), .B(men_men_n394_), .Y(men_men_n396_));
  OAI210     u0374(.A0(men_men_n396_), .A1(men_men_n391_), .B0(men_men_n385_), .Y(men_men_n397_));
  NO2        u0375(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n398_));
  NO2        u0376(.A(men_men_n149_), .B(men_men_n85_), .Y(men_men_n399_));
  OAI210     u0377(.A0(men_men_n399_), .A1(men_men_n391_), .B0(men_men_n398_), .Y(men_men_n400_));
  NO3        u0378(.A(men_men_n85_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n401_));
  NO2        u0379(.A(i_3_), .B(men_men_n100_), .Y(men_men_n402_));
  NO2        u0380(.A(i_11_), .B(i_12_), .Y(men_men_n403_));
  NA2        u0381(.A(men_men_n393_), .B(men_men_n238_), .Y(men_men_n404_));
  NA2        u0382(.A(men_men_n42_), .B(i_11_), .Y(men_men_n405_));
  OAI220     u0383(.A0(men_men_n405_), .A1(men_men_n222_), .B0(men_men_n404_), .B1(men_men_n332_), .Y(men_men_n406_));
  NAi21      u0384(.An(i_13_), .B(i_0_), .Y(men_men_n407_));
  NO2        u0385(.A(men_men_n407_), .B(men_men_n241_), .Y(men_men_n408_));
  NA2        u0386(.A(men_men_n406_), .B(men_men_n408_), .Y(men_men_n409_));
  NA3        u0387(.A(men_men_n409_), .B(men_men_n400_), .C(men_men_n397_), .Y(men_men_n410_));
  NO3        u0388(.A(i_1_), .B(i_12_), .C(men_men_n85_), .Y(men_men_n411_));
  NO2        u0389(.A(i_0_), .B(i_11_), .Y(men_men_n412_));
  AN2        u0390(.A(i_1_), .B(i_6_), .Y(men_men_n413_));
  NOi21      u0391(.An(i_2_), .B(i_12_), .Y(men_men_n414_));
  NA2        u0392(.A(men_men_n414_), .B(men_men_n413_), .Y(men_men_n415_));
  INV        u0393(.A(men_men_n415_), .Y(men_men_n416_));
  NA2        u0394(.A(men_men_n142_), .B(i_9_), .Y(men_men_n417_));
  NO2        u0395(.A(men_men_n417_), .B(i_4_), .Y(men_men_n418_));
  NA2        u0396(.A(men_men_n416_), .B(men_men_n418_), .Y(men_men_n419_));
  NAi21      u0397(.An(i_9_), .B(i_4_), .Y(men_men_n420_));
  OR2        u0398(.A(i_13_), .B(i_10_), .Y(men_men_n421_));
  NO2        u0399(.A(men_men_n172_), .B(men_men_n123_), .Y(men_men_n422_));
  BUFFER     u0400(.A(men_men_n218_), .Y(men_men_n423_));
  NO2        u0401(.A(men_men_n100_), .B(men_men_n25_), .Y(men_men_n424_));
  NA2        u0402(.A(men_men_n276_), .B(men_men_n212_), .Y(men_men_n425_));
  NO2        u0403(.A(men_men_n425_), .B(men_men_n423_), .Y(men_men_n426_));
  INV        u0404(.A(men_men_n426_), .Y(men_men_n427_));
  AOI210     u0405(.A0(men_men_n427_), .A1(men_men_n419_), .B0(men_men_n26_), .Y(men_men_n428_));
  NA2        u0406(.A(men_men_n323_), .B(men_men_n322_), .Y(men_men_n429_));
  AOI220     u0407(.A0(men_men_n296_), .A1(men_men_n286_), .B0(men_men_n290_), .B1(men_men_n314_), .Y(men_men_n430_));
  NO2        u0408(.A(men_men_n430_), .B(i_5_), .Y(men_men_n431_));
  NO2        u0409(.A(men_men_n182_), .B(men_men_n85_), .Y(men_men_n432_));
  AOI220     u0410(.A0(men_men_n432_), .A1(men_men_n295_), .B0(men_men_n278_), .B1(men_men_n212_), .Y(men_men_n433_));
  NO2        u0411(.A(men_men_n433_), .B(men_men_n285_), .Y(men_men_n434_));
  NO3        u0412(.A(men_men_n434_), .B(men_men_n431_), .C(men_men_n429_), .Y(men_men_n435_));
  NA2        u0413(.A(men_men_n196_), .B(men_men_n95_), .Y(men_men_n436_));
  NA3        u0414(.A(men_men_n325_), .B(men_men_n163_), .C(men_men_n85_), .Y(men_men_n437_));
  AOI210     u0415(.A0(men_men_n437_), .A1(men_men_n436_), .B0(i_8_), .Y(men_men_n438_));
  NA2        u0416(.A(men_men_n296_), .B(men_men_n236_), .Y(men_men_n439_));
  NO2        u0417(.A(men_men_n439_), .B(men_men_n182_), .Y(men_men_n440_));
  NO2        u0418(.A(i_3_), .B(men_men_n49_), .Y(men_men_n441_));
  NA3        u0419(.A(men_men_n337_), .B(men_men_n336_), .C(men_men_n441_), .Y(men_men_n442_));
  INV        u0420(.A(men_men_n316_), .Y(men_men_n443_));
  OAI210     u0421(.A0(men_men_n443_), .A1(men_men_n189_), .B0(men_men_n442_), .Y(men_men_n444_));
  NO3        u0422(.A(men_men_n444_), .B(men_men_n440_), .C(men_men_n438_), .Y(men_men_n445_));
  AOI210     u0423(.A0(men_men_n445_), .A1(men_men_n435_), .B0(men_men_n270_), .Y(men_men_n446_));
  NO4        u0424(.A(men_men_n446_), .B(men_men_n428_), .C(men_men_n410_), .D(men_men_n384_), .Y(men_men_n447_));
  NO2        u0425(.A(men_men_n63_), .B(i_4_), .Y(men_men_n448_));
  NO2        u0426(.A(men_men_n73_), .B(i_13_), .Y(men_men_n449_));
  NA3        u0427(.A(men_men_n449_), .B(men_men_n448_), .C(i_2_), .Y(men_men_n450_));
  NO2        u0428(.A(i_10_), .B(i_9_), .Y(men_men_n451_));
  NAi21      u0429(.An(i_12_), .B(i_8_), .Y(men_men_n452_));
  NO2        u0430(.A(men_men_n452_), .B(i_3_), .Y(men_men_n453_));
  NA2        u0431(.A(men_men_n453_), .B(men_men_n451_), .Y(men_men_n454_));
  NO2        u0432(.A(men_men_n47_), .B(i_4_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n455_), .B(men_men_n103_), .Y(men_men_n456_));
  OAI220     u0434(.A0(men_men_n456_), .A1(men_men_n205_), .B0(men_men_n454_), .B1(men_men_n450_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n309_), .B(i_0_), .Y(men_men_n458_));
  NO3        u0436(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n459_));
  NA2        u0437(.A(men_men_n265_), .B(men_men_n96_), .Y(men_men_n460_));
  NA2        u0438(.A(men_men_n460_), .B(men_men_n459_), .Y(men_men_n461_));
  NA2        u0439(.A(i_8_), .B(i_9_), .Y(men_men_n462_));
  AOI210     u0440(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n463_));
  OR2        u0441(.A(men_men_n463_), .B(men_men_n462_), .Y(men_men_n464_));
  NA2        u0442(.A(men_men_n283_), .B(men_men_n206_), .Y(men_men_n465_));
  OAI220     u0443(.A0(men_men_n465_), .A1(men_men_n464_), .B0(men_men_n461_), .B1(men_men_n458_), .Y(men_men_n466_));
  NA2        u0444(.A(men_men_n253_), .B(men_men_n308_), .Y(men_men_n467_));
  NO3        u0445(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n468_));
  INV        u0446(.A(men_men_n468_), .Y(men_men_n469_));
  NA3        u0447(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n470_));
  NA4        u0448(.A(men_men_n145_), .B(men_men_n115_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n471_));
  OAI220     u0449(.A0(men_men_n471_), .A1(men_men_n470_), .B0(men_men_n469_), .B1(men_men_n467_), .Y(men_men_n472_));
  NO3        u0450(.A(men_men_n472_), .B(men_men_n466_), .C(men_men_n457_), .Y(men_men_n473_));
  NA2        u0451(.A(men_men_n295_), .B(men_men_n107_), .Y(men_men_n474_));
  OR2        u0452(.A(men_men_n474_), .B(men_men_n208_), .Y(men_men_n475_));
  BUFFER     u0453(.A(men_men_n354_), .Y(men_men_n476_));
  OA220      u0454(.A0(men_men_n476_), .A1(men_men_n162_), .B0(men_men_n475_), .B1(men_men_n233_), .Y(men_men_n477_));
  NA2        u0455(.A(men_men_n95_), .B(i_13_), .Y(men_men_n478_));
  NA2        u0456(.A(men_men_n432_), .B(men_men_n385_), .Y(men_men_n479_));
  NO2        u0457(.A(i_2_), .B(i_13_), .Y(men_men_n480_));
  NO2        u0458(.A(men_men_n479_), .B(men_men_n478_), .Y(men_men_n481_));
  NO3        u0459(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n482_));
  NO2        u0460(.A(i_6_), .B(i_7_), .Y(men_men_n483_));
  NA2        u0461(.A(men_men_n483_), .B(men_men_n482_), .Y(men_men_n484_));
  NO2        u0462(.A(i_11_), .B(i_1_), .Y(men_men_n485_));
  OR2        u0463(.A(i_11_), .B(i_8_), .Y(men_men_n486_));
  NOi21      u0464(.An(i_2_), .B(i_7_), .Y(men_men_n487_));
  NAi31      u0465(.An(men_men_n486_), .B(men_men_n487_), .C(i_0_), .Y(men_men_n488_));
  NO2        u0466(.A(men_men_n421_), .B(i_6_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n489_), .B(men_men_n448_), .Y(men_men_n490_));
  NO2        u0468(.A(men_men_n490_), .B(men_men_n488_), .Y(men_men_n491_));
  NO2        u0469(.A(i_3_), .B(men_men_n193_), .Y(men_men_n492_));
  NO2        u0470(.A(i_6_), .B(i_10_), .Y(men_men_n493_));
  NA4        u0471(.A(men_men_n493_), .B(men_men_n313_), .C(men_men_n492_), .D(men_men_n238_), .Y(men_men_n494_));
  NO2        u0472(.A(men_men_n494_), .B(men_men_n155_), .Y(men_men_n495_));
  NA3        u0473(.A(men_men_n247_), .B(men_men_n171_), .C(men_men_n132_), .Y(men_men_n496_));
  NO2        u0474(.A(men_men_n157_), .B(i_3_), .Y(men_men_n497_));
  NO4        u0475(.A(men_men_n1080_), .B(men_men_n495_), .C(men_men_n491_), .D(men_men_n481_), .Y(men_men_n498_));
  NA2        u0476(.A(men_men_n459_), .B(men_men_n386_), .Y(men_men_n499_));
  NA2        u0477(.A(men_men_n468_), .B(men_men_n393_), .Y(men_men_n500_));
  NO2        u0478(.A(men_men_n500_), .B(men_men_n225_), .Y(men_men_n501_));
  NAi21      u0479(.An(men_men_n218_), .B(men_men_n403_), .Y(men_men_n502_));
  NA2        u0480(.A(men_men_n337_), .B(men_men_n220_), .Y(men_men_n503_));
  NO2        u0481(.A(men_men_n26_), .B(i_5_), .Y(men_men_n504_));
  NA3        u0482(.A(i_6_), .B(men_men_n504_), .C(men_men_n142_), .Y(men_men_n505_));
  OR3        u0483(.A(men_men_n303_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n506_));
  OAI220     u0484(.A0(men_men_n506_), .A1(men_men_n505_), .B0(men_men_n503_), .B1(men_men_n502_), .Y(men_men_n507_));
  NA2        u0485(.A(men_men_n27_), .B(i_10_), .Y(men_men_n508_));
  NO2        u0486(.A(men_men_n508_), .B(men_men_n478_), .Y(men_men_n509_));
  NA4        u0487(.A(men_men_n306_), .B(men_men_n224_), .C(men_men_n73_), .D(men_men_n238_), .Y(men_men_n510_));
  NO2        u0488(.A(men_men_n510_), .B(men_men_n484_), .Y(men_men_n511_));
  NO4        u0489(.A(men_men_n511_), .B(men_men_n509_), .C(men_men_n507_), .D(men_men_n501_), .Y(men_men_n512_));
  NA4        u0490(.A(men_men_n512_), .B(men_men_n498_), .C(men_men_n477_), .D(men_men_n473_), .Y(men_men_n513_));
  NA3        u0491(.A(men_men_n306_), .B(men_men_n175_), .C(men_men_n173_), .Y(men_men_n514_));
  OAI210     u0492(.A0(men_men_n301_), .A1(men_men_n180_), .B0(men_men_n514_), .Y(men_men_n515_));
  AN2        u0493(.A(men_men_n286_), .B(men_men_n235_), .Y(men_men_n516_));
  NA2        u0494(.A(men_men_n516_), .B(men_men_n515_), .Y(men_men_n517_));
  NA2        u0495(.A(men_men_n122_), .B(men_men_n111_), .Y(men_men_n518_));
  AN2        u0496(.A(men_men_n518_), .B(men_men_n459_), .Y(men_men_n519_));
  NA2        u0497(.A(men_men_n313_), .B(men_men_n164_), .Y(men_men_n520_));
  OAI210     u0498(.A0(men_men_n520_), .A1(men_men_n233_), .B0(men_men_n307_), .Y(men_men_n521_));
  AOI220     u0499(.A0(men_men_n521_), .A1(men_men_n324_), .B0(men_men_n519_), .B1(men_men_n309_), .Y(men_men_n522_));
  NA4        u0500(.A(men_men_n449_), .B(men_men_n448_), .C(men_men_n203_), .D(i_2_), .Y(men_men_n523_));
  INV        u0501(.A(men_men_n523_), .Y(men_men_n524_));
  NA2        u0502(.A(men_men_n358_), .B(men_men_n73_), .Y(men_men_n525_));
  NA2        u0503(.A(men_men_n374_), .B(men_men_n366_), .Y(men_men_n526_));
  NO2        u0504(.A(men_men_n36_), .B(i_8_), .Y(men_men_n527_));
  NAi41      u0505(.An(men_men_n525_), .B(men_men_n493_), .C(men_men_n527_), .D(men_men_n47_), .Y(men_men_n528_));
  NA2        u0506(.A(men_men_n39_), .B(i_13_), .Y(men_men_n529_));
  NA2        u0507(.A(men_men_n529_), .B(men_men_n528_), .Y(men_men_n530_));
  AOI210     u0508(.A0(men_men_n524_), .A1(men_men_n204_), .B0(men_men_n530_), .Y(men_men_n531_));
  OAI210     u0509(.A0(i_8_), .A1(men_men_n63_), .B0(men_men_n134_), .Y(men_men_n532_));
  AOI210     u0510(.A0(men_men_n194_), .A1(i_9_), .B0(men_men_n264_), .Y(men_men_n533_));
  NO2        u0511(.A(men_men_n533_), .B(men_men_n199_), .Y(men_men_n534_));
  NO2        u0512(.A(men_men_n182_), .B(men_men_n85_), .Y(men_men_n535_));
  AOI220     u0513(.A0(men_men_n535_), .A1(men_men_n534_), .B0(men_men_n532_), .B1(men_men_n422_), .Y(men_men_n536_));
  NA4        u0514(.A(men_men_n536_), .B(men_men_n531_), .C(men_men_n522_), .D(men_men_n517_), .Y(men_men_n537_));
  NA2        u0515(.A(men_men_n392_), .B(men_men_n295_), .Y(men_men_n538_));
  OAI210     u0516(.A0(men_men_n388_), .A1(men_men_n169_), .B0(men_men_n538_), .Y(men_men_n539_));
  NO2        u0517(.A(i_12_), .B(men_men_n193_), .Y(men_men_n540_));
  NA2        u0518(.A(men_men_n540_), .B(men_men_n226_), .Y(men_men_n541_));
  NO3        u0519(.A(i_10_), .B(men_men_n541_), .C(men_men_n474_), .Y(men_men_n542_));
  NOi31      u0520(.An(men_men_n316_), .B(men_men_n421_), .C(men_men_n38_), .Y(men_men_n543_));
  OAI210     u0521(.A0(men_men_n543_), .A1(men_men_n542_), .B0(men_men_n539_), .Y(men_men_n544_));
  NO2        u0522(.A(i_8_), .B(i_7_), .Y(men_men_n545_));
  OAI210     u0523(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n546_));
  NA2        u0524(.A(men_men_n546_), .B(men_men_n224_), .Y(men_men_n547_));
  AOI220     u0525(.A0(men_men_n325_), .A1(men_men_n40_), .B0(men_men_n236_), .B1(men_men_n207_), .Y(men_men_n548_));
  OAI220     u0526(.A0(men_men_n548_), .A1(men_men_n182_), .B0(men_men_n547_), .B1(men_men_n244_), .Y(men_men_n549_));
  NA2        u0527(.A(men_men_n45_), .B(i_10_), .Y(men_men_n550_));
  NO2        u0528(.A(men_men_n550_), .B(i_6_), .Y(men_men_n551_));
  NA3        u0529(.A(men_men_n551_), .B(men_men_n549_), .C(men_men_n545_), .Y(men_men_n552_));
  AOI220     u0530(.A0(men_men_n432_), .A1(men_men_n325_), .B0(men_men_n249_), .B1(men_men_n246_), .Y(men_men_n553_));
  OAI220     u0531(.A0(men_men_n553_), .A1(men_men_n261_), .B0(men_men_n478_), .B1(men_men_n133_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n554_), .B(men_men_n264_), .Y(men_men_n555_));
  NO2        u0533(.A(men_men_n301_), .B(men_men_n180_), .Y(men_men_n556_));
  NA3        u0534(.A(men_men_n306_), .B(men_men_n173_), .C(men_men_n95_), .Y(men_men_n557_));
  NO2        u0535(.A(men_men_n223_), .B(men_men_n45_), .Y(men_men_n558_));
  NO2        u0536(.A(men_men_n157_), .B(i_5_), .Y(men_men_n559_));
  NA2        u0537(.A(men_men_n559_), .B(men_men_n319_), .Y(men_men_n560_));
  OAI210     u0538(.A0(men_men_n560_), .A1(men_men_n558_), .B0(men_men_n557_), .Y(men_men_n561_));
  OAI210     u0539(.A0(men_men_n561_), .A1(men_men_n556_), .B0(men_men_n468_), .Y(men_men_n562_));
  NA4        u0540(.A(men_men_n562_), .B(men_men_n555_), .C(men_men_n552_), .D(men_men_n544_), .Y(men_men_n563_));
  NA3        u0541(.A(men_men_n220_), .B(men_men_n71_), .C(men_men_n45_), .Y(men_men_n564_));
  NA2        u0542(.A(men_men_n283_), .B(men_men_n84_), .Y(men_men_n565_));
  AOI210     u0543(.A0(men_men_n564_), .A1(men_men_n349_), .B0(men_men_n565_), .Y(men_men_n566_));
  NA2        u0544(.A(men_men_n296_), .B(men_men_n286_), .Y(men_men_n567_));
  NO2        u0545(.A(men_men_n567_), .B(men_men_n172_), .Y(men_men_n568_));
  AOI210     u0546(.A0(men_men_n367_), .A1(men_men_n47_), .B0(men_men_n371_), .Y(men_men_n569_));
  NA2        u0547(.A(i_0_), .B(men_men_n49_), .Y(men_men_n570_));
  NA3        u0548(.A(men_men_n540_), .B(men_men_n274_), .C(men_men_n570_), .Y(men_men_n571_));
  NO2        u0549(.A(men_men_n569_), .B(men_men_n571_), .Y(men_men_n572_));
  NO3        u0550(.A(men_men_n572_), .B(men_men_n568_), .C(men_men_n566_), .Y(men_men_n573_));
  NO4        u0551(.A(men_men_n254_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n574_));
  NO3        u0552(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n575_));
  NO2        u0553(.A(men_men_n234_), .B(men_men_n36_), .Y(men_men_n576_));
  AN2        u0554(.A(men_men_n576_), .B(men_men_n575_), .Y(men_men_n577_));
  OA210      u0555(.A0(men_men_n577_), .A1(men_men_n574_), .B0(men_men_n358_), .Y(men_men_n578_));
  NO2        u0556(.A(men_men_n421_), .B(i_1_), .Y(men_men_n579_));
  NOi31      u0557(.An(men_men_n579_), .B(men_men_n460_), .C(men_men_n73_), .Y(men_men_n580_));
  AN4        u0558(.A(men_men_n580_), .B(men_men_n418_), .C(men_men_n504_), .D(i_2_), .Y(men_men_n581_));
  NO2        u0559(.A(men_men_n430_), .B(men_men_n176_), .Y(men_men_n582_));
  NO3        u0560(.A(men_men_n582_), .B(men_men_n581_), .C(men_men_n578_), .Y(men_men_n583_));
  NOi21      u0561(.An(i_10_), .B(i_6_), .Y(men_men_n584_));
  NO2        u0562(.A(men_men_n85_), .B(men_men_n25_), .Y(men_men_n585_));
  AOI220     u0563(.A0(men_men_n283_), .A1(men_men_n585_), .B0(men_men_n274_), .B1(men_men_n584_), .Y(men_men_n586_));
  NO2        u0564(.A(men_men_n586_), .B(men_men_n458_), .Y(men_men_n587_));
  NO2        u0565(.A(men_men_n114_), .B(men_men_n23_), .Y(men_men_n588_));
  NA2        u0566(.A(men_men_n316_), .B(men_men_n164_), .Y(men_men_n589_));
  AOI220     u0567(.A0(men_men_n589_), .A1(men_men_n439_), .B0(men_men_n183_), .B1(men_men_n181_), .Y(men_men_n590_));
  NO2        u0568(.A(men_men_n198_), .B(men_men_n37_), .Y(men_men_n591_));
  NOi31      u0569(.An(men_men_n146_), .B(men_men_n591_), .C(men_men_n332_), .Y(men_men_n592_));
  NO3        u0570(.A(men_men_n592_), .B(men_men_n590_), .C(men_men_n587_), .Y(men_men_n593_));
  NO2        u0571(.A(men_men_n525_), .B(men_men_n381_), .Y(men_men_n594_));
  INV        u0572(.A(men_men_n319_), .Y(men_men_n595_));
  NO2        u0573(.A(i_12_), .B(men_men_n85_), .Y(men_men_n596_));
  NA3        u0574(.A(men_men_n596_), .B(men_men_n274_), .C(men_men_n570_), .Y(men_men_n597_));
  NA3        u0575(.A(men_men_n389_), .B(men_men_n283_), .C(men_men_n220_), .Y(men_men_n598_));
  AOI210     u0576(.A0(men_men_n598_), .A1(men_men_n597_), .B0(men_men_n595_), .Y(men_men_n599_));
  NA2        u0577(.A(men_men_n173_), .B(i_0_), .Y(men_men_n600_));
  NO3        u0578(.A(men_men_n600_), .B(men_men_n343_), .C(men_men_n301_), .Y(men_men_n601_));
  OR2        u0579(.A(i_2_), .B(i_5_), .Y(men_men_n602_));
  OR2        u0580(.A(men_men_n602_), .B(men_men_n413_), .Y(men_men_n603_));
  NO2        u0581(.A(men_men_n603_), .B(men_men_n502_), .Y(men_men_n604_));
  NO4        u0582(.A(men_men_n604_), .B(men_men_n601_), .C(men_men_n599_), .D(men_men_n594_), .Y(men_men_n605_));
  NA4        u0583(.A(men_men_n605_), .B(men_men_n593_), .C(men_men_n583_), .D(men_men_n573_), .Y(men_men_n606_));
  NO4        u0584(.A(men_men_n606_), .B(men_men_n563_), .C(men_men_n537_), .D(men_men_n513_), .Y(men_men_n607_));
  NA4        u0585(.A(men_men_n607_), .B(men_men_n447_), .C(men_men_n357_), .D(men_men_n312_), .Y(men7));
  NO2        u0586(.A(men_men_n92_), .B(men_men_n55_), .Y(men_men_n609_));
  NO2        u0587(.A(men_men_n107_), .B(men_men_n89_), .Y(men_men_n610_));
  NA2        u0588(.A(men_men_n387_), .B(men_men_n610_), .Y(men_men_n611_));
  NA2        u0589(.A(men_men_n493_), .B(men_men_n84_), .Y(men_men_n612_));
  NA2        u0590(.A(i_11_), .B(men_men_n193_), .Y(men_men_n613_));
  NA2        u0591(.A(men_men_n144_), .B(men_men_n613_), .Y(men_men_n614_));
  OAI210     u0592(.A0(men_men_n614_), .A1(men_men_n612_), .B0(men_men_n611_), .Y(men_men_n615_));
  NA3        u0593(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n616_));
  NO2        u0594(.A(men_men_n238_), .B(i_4_), .Y(men_men_n617_));
  NA2        u0595(.A(men_men_n617_), .B(i_8_), .Y(men_men_n618_));
  NO2        u0596(.A(men_men_n104_), .B(men_men_n616_), .Y(men_men_n619_));
  NA2        u0597(.A(i_2_), .B(men_men_n85_), .Y(men_men_n620_));
  OAI210     u0598(.A0(men_men_n88_), .A1(men_men_n203_), .B0(men_men_n204_), .Y(men_men_n621_));
  NO2        u0599(.A(i_7_), .B(men_men_n37_), .Y(men_men_n622_));
  NA2        u0600(.A(i_4_), .B(i_8_), .Y(men_men_n623_));
  AOI210     u0601(.A0(men_men_n623_), .A1(men_men_n306_), .B0(men_men_n622_), .Y(men_men_n624_));
  NO2        u0602(.A(men_men_n624_), .B(men_men_n620_), .Y(men_men_n625_));
  NO4        u0603(.A(men_men_n625_), .B(men_men_n619_), .C(men_men_n615_), .D(men_men_n609_), .Y(men_men_n626_));
  OR2        u0604(.A(i_6_), .B(i_10_), .Y(men_men_n627_));
  NO2        u0605(.A(men_men_n627_), .B(men_men_n23_), .Y(men_men_n628_));
  OR3        u0606(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n629_));
  NO3        u0607(.A(men_men_n629_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n630_));
  INV        u0608(.A(men_men_n200_), .Y(men_men_n631_));
  NO2        u0609(.A(men_men_n630_), .B(men_men_n628_), .Y(men_men_n632_));
  OA220      u0610(.A0(men_men_n632_), .A1(men_men_n595_), .B0(men_men_n1079_), .B1(men_men_n266_), .Y(men_men_n633_));
  AOI210     u0611(.A0(men_men_n633_), .A1(men_men_n626_), .B0(men_men_n63_), .Y(men_men_n634_));
  NOi21      u0612(.An(i_11_), .B(i_7_), .Y(men_men_n635_));
  AO210      u0613(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n636_));
  NO2        u0614(.A(men_men_n636_), .B(men_men_n635_), .Y(men_men_n637_));
  NA2        u0615(.A(men_men_n637_), .B(men_men_n207_), .Y(men_men_n638_));
  NA3        u0616(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n639_));
  NAi31      u0617(.An(men_men_n639_), .B(men_men_n217_), .C(i_11_), .Y(men_men_n640_));
  AOI210     u0618(.A0(men_men_n640_), .A1(men_men_n638_), .B0(men_men_n63_), .Y(men_men_n641_));
  NA2        u0619(.A(men_men_n87_), .B(men_men_n63_), .Y(men_men_n642_));
  AO210      u0620(.A0(men_men_n642_), .A1(men_men_n381_), .B0(men_men_n41_), .Y(men_men_n643_));
  NA2        u0621(.A(men_men_n227_), .B(men_men_n63_), .Y(men_men_n644_));
  NA2        u0622(.A(men_men_n414_), .B(men_men_n31_), .Y(men_men_n645_));
  OR2        u0623(.A(men_men_n209_), .B(men_men_n107_), .Y(men_men_n646_));
  NA2        u0624(.A(men_men_n646_), .B(men_men_n645_), .Y(men_men_n647_));
  NO2        u0625(.A(men_men_n63_), .B(i_9_), .Y(men_men_n648_));
  NO2        u0626(.A(men_men_n648_), .B(i_4_), .Y(men_men_n649_));
  NA2        u0627(.A(men_men_n649_), .B(men_men_n647_), .Y(men_men_n650_));
  NO2        u0628(.A(i_1_), .B(i_12_), .Y(men_men_n651_));
  NA3        u0629(.A(men_men_n651_), .B(men_men_n109_), .C(men_men_n24_), .Y(men_men_n652_));
  NA4        u0630(.A(men_men_n652_), .B(men_men_n650_), .C(men_men_n644_), .D(men_men_n643_), .Y(men_men_n653_));
  OAI210     u0631(.A0(men_men_n653_), .A1(men_men_n641_), .B0(i_6_), .Y(men_men_n654_));
  NO2        u0632(.A(men_men_n238_), .B(men_men_n85_), .Y(men_men_n655_));
  NO2        u0633(.A(men_men_n655_), .B(i_11_), .Y(men_men_n656_));
  INV        u0634(.A(men_men_n461_), .Y(men_men_n657_));
  NO4        u0635(.A(men_men_n217_), .B(men_men_n128_), .C(i_13_), .D(men_men_n85_), .Y(men_men_n658_));
  NA2        u0636(.A(men_men_n658_), .B(men_men_n648_), .Y(men_men_n659_));
  INV        u0637(.A(men_men_n659_), .Y(men_men_n660_));
  NA3        u0638(.A(men_men_n545_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n661_));
  NA2        u0639(.A(men_men_n138_), .B(i_9_), .Y(men_men_n662_));
  NA3        u0640(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n663_));
  NO2        u0641(.A(men_men_n47_), .B(i_1_), .Y(men_men_n664_));
  NO2        u0642(.A(men_men_n662_), .B(men_men_n1077_), .Y(men_men_n665_));
  NA3        u0643(.A(men_men_n648_), .B(men_men_n319_), .C(i_6_), .Y(men_men_n666_));
  NO2        u0644(.A(men_men_n666_), .B(men_men_n23_), .Y(men_men_n667_));
  AOI210     u0645(.A0(men_men_n485_), .A1(men_men_n424_), .B0(men_men_n243_), .Y(men_men_n668_));
  NO2        u0646(.A(men_men_n668_), .B(men_men_n620_), .Y(men_men_n669_));
  NA2        u0647(.A(men_men_n664_), .B(men_men_n265_), .Y(men_men_n670_));
  NO2        u0648(.A(i_11_), .B(men_men_n37_), .Y(men_men_n671_));
  NA2        u0649(.A(men_men_n671_), .B(men_men_n24_), .Y(men_men_n672_));
  NO2        u0650(.A(men_men_n672_), .B(men_men_n670_), .Y(men_men_n673_));
  OR4        u0651(.A(men_men_n673_), .B(men_men_n669_), .C(men_men_n667_), .D(men_men_n665_), .Y(men_men_n674_));
  NO3        u0652(.A(men_men_n674_), .B(men_men_n660_), .C(men_men_n657_), .Y(men_men_n675_));
  NO2        u0653(.A(men_men_n238_), .B(men_men_n100_), .Y(men_men_n676_));
  NO2        u0654(.A(men_men_n676_), .B(men_men_n635_), .Y(men_men_n677_));
  NA2        u0655(.A(men_men_n677_), .B(i_1_), .Y(men_men_n678_));
  NO2        u0656(.A(men_men_n678_), .B(men_men_n629_), .Y(men_men_n679_));
  NO2        u0657(.A(men_men_n420_), .B(men_men_n85_), .Y(men_men_n680_));
  NA2        u0658(.A(men_men_n679_), .B(men_men_n47_), .Y(men_men_n681_));
  NA2        u0659(.A(i_3_), .B(men_men_n193_), .Y(men_men_n682_));
  NO2        u0660(.A(men_men_n234_), .B(men_men_n45_), .Y(men_men_n683_));
  NO3        u0661(.A(men_men_n683_), .B(men_men_n309_), .C(men_men_n239_), .Y(men_men_n684_));
  NO2        u0662(.A(men_men_n117_), .B(men_men_n37_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n685_), .B(i_6_), .Y(men_men_n686_));
  NO2        u0664(.A(men_men_n85_), .B(i_9_), .Y(men_men_n687_));
  NO2        u0665(.A(men_men_n687_), .B(men_men_n63_), .Y(men_men_n688_));
  NO2        u0666(.A(men_men_n688_), .B(men_men_n651_), .Y(men_men_n689_));
  NO4        u0667(.A(men_men_n689_), .B(men_men_n686_), .C(men_men_n684_), .D(i_4_), .Y(men_men_n690_));
  NA2        u0668(.A(i_1_), .B(i_3_), .Y(men_men_n691_));
  INV        u0669(.A(men_men_n690_), .Y(men_men_n692_));
  NA4        u0670(.A(men_men_n692_), .B(men_men_n681_), .C(men_men_n675_), .D(men_men_n654_), .Y(men_men_n693_));
  NO3        u0671(.A(men_men_n486_), .B(i_3_), .C(i_7_), .Y(men_men_n694_));
  NOi21      u0672(.An(men_men_n694_), .B(i_10_), .Y(men_men_n695_));
  OA210      u0673(.A0(men_men_n695_), .A1(men_men_n247_), .B0(men_men_n85_), .Y(men_men_n696_));
  NA3        u0674(.A(men_men_n493_), .B(men_men_n527_), .C(men_men_n47_), .Y(men_men_n697_));
  NO3        u0675(.A(men_men_n487_), .B(men_men_n623_), .C(men_men_n85_), .Y(men_men_n698_));
  NA2        u0676(.A(men_men_n698_), .B(men_men_n25_), .Y(men_men_n699_));
  NA3        u0677(.A(men_men_n161_), .B(men_men_n84_), .C(men_men_n85_), .Y(men_men_n700_));
  NA3        u0678(.A(men_men_n700_), .B(men_men_n699_), .C(men_men_n697_), .Y(men_men_n701_));
  OAI210     u0679(.A0(men_men_n701_), .A1(men_men_n696_), .B0(i_1_), .Y(men_men_n702_));
  AOI210     u0680(.A0(men_men_n265_), .A1(men_men_n96_), .B0(i_1_), .Y(men_men_n703_));
  NO2        u0681(.A(men_men_n372_), .B(i_2_), .Y(men_men_n704_));
  NA2        u0682(.A(men_men_n704_), .B(men_men_n703_), .Y(men_men_n705_));
  OAI210     u0683(.A0(men_men_n666_), .A1(men_men_n452_), .B0(men_men_n705_), .Y(men_men_n706_));
  INV        u0684(.A(men_men_n706_), .Y(men_men_n707_));
  AOI210     u0685(.A0(men_men_n707_), .A1(men_men_n702_), .B0(i_13_), .Y(men_men_n708_));
  NA3        u0686(.A(i_11_), .B(men_men_n105_), .C(men_men_n138_), .Y(men_men_n709_));
  AOI220     u0687(.A0(men_men_n480_), .A1(men_men_n161_), .B0(men_men_n455_), .B1(men_men_n138_), .Y(men_men_n710_));
  OAI210     u0688(.A0(men_men_n710_), .A1(men_men_n45_), .B0(men_men_n709_), .Y(men_men_n711_));
  NO2        u0689(.A(men_men_n55_), .B(i_12_), .Y(men_men_n712_));
  INV        u0690(.A(men_men_n712_), .Y(men_men_n713_));
  NO2        u0691(.A(men_men_n487_), .B(men_men_n24_), .Y(men_men_n714_));
  AOI220     u0692(.A0(men_men_n714_), .A1(men_men_n680_), .B0(men_men_n247_), .B1(men_men_n131_), .Y(men_men_n715_));
  OAI220     u0693(.A0(men_men_n715_), .A1(men_men_n41_), .B0(men_men_n713_), .B1(men_men_n92_), .Y(men_men_n716_));
  AOI210     u0694(.A0(men_men_n711_), .A1(men_men_n334_), .B0(men_men_n716_), .Y(men_men_n717_));
  AOI220     u0695(.A0(i_12_), .A1(men_men_n72_), .B0(men_men_n389_), .B1(men_men_n664_), .Y(men_men_n718_));
  NO2        u0696(.A(men_men_n718_), .B(men_men_n244_), .Y(men_men_n719_));
  AOI210     u0697(.A0(men_men_n452_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n720_));
  NOi31      u0698(.An(men_men_n720_), .B(men_men_n612_), .C(men_men_n45_), .Y(men_men_n721_));
  NA2        u0699(.A(men_men_n127_), .B(i_13_), .Y(men_men_n722_));
  NO2        u0700(.A(men_men_n663_), .B(men_men_n114_), .Y(men_men_n723_));
  NO2        u0701(.A(men_men_n722_), .B(men_men_n703_), .Y(men_men_n724_));
  NO3        u0702(.A(men_men_n71_), .B(men_men_n32_), .C(men_men_n100_), .Y(men_men_n725_));
  NA2        u0703(.A(men_men_n26_), .B(men_men_n193_), .Y(men_men_n726_));
  INV        u0704(.A(men_men_n725_), .Y(men_men_n727_));
  NO2        u0705(.A(men_men_n727_), .B(men_men_n631_), .Y(men_men_n728_));
  NO4        u0706(.A(men_men_n728_), .B(men_men_n724_), .C(men_men_n721_), .D(men_men_n719_), .Y(men_men_n729_));
  OR2        u0707(.A(i_11_), .B(i_6_), .Y(men_men_n730_));
  NA3        u0708(.A(men_men_n617_), .B(men_men_n726_), .C(i_7_), .Y(men_men_n731_));
  NO2        u0709(.A(men_men_n731_), .B(men_men_n730_), .Y(men_men_n732_));
  NA3        u0710(.A(men_men_n414_), .B(men_men_n622_), .C(men_men_n96_), .Y(men_men_n733_));
  NA2        u0711(.A(men_men_n656_), .B(i_13_), .Y(men_men_n734_));
  NA2        u0712(.A(men_men_n101_), .B(men_men_n726_), .Y(men_men_n735_));
  NAi21      u0713(.An(i_11_), .B(i_12_), .Y(men_men_n736_));
  NOi41      u0714(.An(men_men_n110_), .B(men_men_n736_), .C(i_13_), .D(men_men_n85_), .Y(men_men_n737_));
  NO3        u0715(.A(men_men_n487_), .B(men_men_n596_), .C(men_men_n623_), .Y(men_men_n738_));
  AOI220     u0716(.A0(men_men_n738_), .A1(men_men_n313_), .B0(men_men_n737_), .B1(men_men_n735_), .Y(men_men_n739_));
  NA3        u0717(.A(men_men_n739_), .B(men_men_n734_), .C(men_men_n733_), .Y(men_men_n740_));
  OAI210     u0718(.A0(men_men_n740_), .A1(men_men_n732_), .B0(men_men_n63_), .Y(men_men_n741_));
  NO2        u0719(.A(i_2_), .B(i_12_), .Y(men_men_n742_));
  NA2        u0720(.A(men_men_n371_), .B(men_men_n742_), .Y(men_men_n743_));
  NA2        u0721(.A(i_8_), .B(men_men_n25_), .Y(men_men_n744_));
  NO3        u0722(.A(men_men_n744_), .B(men_men_n387_), .C(men_men_n617_), .Y(men_men_n745_));
  OAI210     u0723(.A0(men_men_n745_), .A1(men_men_n373_), .B0(men_men_n371_), .Y(men_men_n746_));
  NO2        u0724(.A(men_men_n128_), .B(i_2_), .Y(men_men_n747_));
  NA2        u0725(.A(men_men_n746_), .B(men_men_n743_), .Y(men_men_n748_));
  NA3        u0726(.A(men_men_n748_), .B(men_men_n46_), .C(men_men_n226_), .Y(men_men_n749_));
  NA4        u0727(.A(men_men_n749_), .B(men_men_n741_), .C(men_men_n729_), .D(men_men_n717_), .Y(men_men_n750_));
  OR4        u0728(.A(men_men_n750_), .B(men_men_n708_), .C(men_men_n693_), .D(men_men_n634_), .Y(men5));
  AOI210     u0729(.A0(men_men_n677_), .A1(men_men_n268_), .B0(men_men_n422_), .Y(men_men_n752_));
  AN2        u0730(.A(men_men_n24_), .B(i_10_), .Y(men_men_n753_));
  NA3        u0731(.A(men_men_n753_), .B(men_men_n742_), .C(men_men_n107_), .Y(men_men_n754_));
  NO2        u0732(.A(men_men_n618_), .B(i_11_), .Y(men_men_n755_));
  NA2        u0733(.A(men_men_n88_), .B(men_men_n755_), .Y(men_men_n756_));
  NA3        u0734(.A(men_men_n756_), .B(men_men_n754_), .C(men_men_n752_), .Y(men_men_n757_));
  NO3        u0735(.A(i_11_), .B(men_men_n238_), .C(i_13_), .Y(men_men_n758_));
  NO2        u0736(.A(men_men_n124_), .B(men_men_n23_), .Y(men_men_n759_));
  NA2        u0737(.A(i_12_), .B(i_8_), .Y(men_men_n760_));
  OAI210     u0738(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n760_), .Y(men_men_n761_));
  INV        u0739(.A(men_men_n451_), .Y(men_men_n762_));
  AOI220     u0740(.A0(men_men_n319_), .A1(men_men_n588_), .B0(men_men_n761_), .B1(men_men_n759_), .Y(men_men_n763_));
  INV        u0741(.A(men_men_n763_), .Y(men_men_n764_));
  NO2        u0742(.A(men_men_n764_), .B(men_men_n757_), .Y(men_men_n765_));
  INV        u0743(.A(men_men_n171_), .Y(men_men_n766_));
  INV        u0744(.A(men_men_n247_), .Y(men_men_n767_));
  OAI210     u0745(.A0(men_men_n704_), .A1(men_men_n453_), .B0(men_men_n110_), .Y(men_men_n768_));
  AOI210     u0746(.A0(men_men_n768_), .A1(men_men_n767_), .B0(men_men_n766_), .Y(men_men_n769_));
  NO2        u0747(.A(men_men_n462_), .B(men_men_n26_), .Y(men_men_n770_));
  NO2        u0748(.A(men_men_n770_), .B(men_men_n424_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n771_), .B(i_2_), .Y(men_men_n772_));
  INV        u0750(.A(men_men_n772_), .Y(men_men_n773_));
  AOI210     u0751(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n421_), .Y(men_men_n774_));
  AOI210     u0752(.A0(men_men_n774_), .A1(men_men_n773_), .B0(men_men_n769_), .Y(men_men_n775_));
  NO2        u0753(.A(men_men_n190_), .B(men_men_n125_), .Y(men_men_n776_));
  OAI210     u0754(.A0(men_men_n776_), .A1(men_men_n759_), .B0(i_2_), .Y(men_men_n777_));
  NO2        u0755(.A(men_men_n777_), .B(men_men_n193_), .Y(men_men_n778_));
  OA210      u0756(.A0(men_men_n637_), .A1(men_men_n126_), .B0(i_13_), .Y(men_men_n779_));
  NA2        u0757(.A(men_men_n200_), .B(men_men_n203_), .Y(men_men_n780_));
  NA2        u0758(.A(men_men_n151_), .B(men_men_n613_), .Y(men_men_n781_));
  AOI210     u0759(.A0(men_men_n781_), .A1(men_men_n780_), .B0(men_men_n376_), .Y(men_men_n782_));
  AOI210     u0760(.A0(men_men_n209_), .A1(men_men_n148_), .B0(men_men_n527_), .Y(men_men_n783_));
  NA2        u0761(.A(men_men_n783_), .B(men_men_n424_), .Y(men_men_n784_));
  NO2        u0762(.A(men_men_n101_), .B(men_men_n45_), .Y(men_men_n785_));
  INV        u0763(.A(men_men_n302_), .Y(men_men_n786_));
  NA4        u0764(.A(men_men_n786_), .B(men_men_n306_), .C(men_men_n124_), .D(men_men_n43_), .Y(men_men_n787_));
  OAI210     u0765(.A0(men_men_n787_), .A1(men_men_n785_), .B0(men_men_n784_), .Y(men_men_n788_));
  NO4        u0766(.A(men_men_n788_), .B(men_men_n782_), .C(men_men_n779_), .D(men_men_n778_), .Y(men_men_n789_));
  NA2        u0767(.A(men_men_n588_), .B(men_men_n28_), .Y(men_men_n790_));
  NA2        u0768(.A(men_men_n758_), .B(men_men_n275_), .Y(men_men_n791_));
  NA2        u0769(.A(men_men_n791_), .B(men_men_n790_), .Y(men_men_n792_));
  NO2        u0770(.A(men_men_n62_), .B(i_12_), .Y(men_men_n793_));
  NO2        u0771(.A(men_men_n793_), .B(men_men_n126_), .Y(men_men_n794_));
  NO2        u0772(.A(men_men_n794_), .B(men_men_n613_), .Y(men_men_n795_));
  AOI220     u0773(.A0(men_men_n795_), .A1(men_men_n36_), .B0(men_men_n792_), .B1(men_men_n47_), .Y(men_men_n796_));
  NA4        u0774(.A(men_men_n796_), .B(men_men_n789_), .C(men_men_n775_), .D(men_men_n765_), .Y(men6));
  NO3        u0775(.A(men_men_n256_), .B(men_men_n308_), .C(i_1_), .Y(men_men_n798_));
  NO2        u0776(.A(men_men_n185_), .B(men_men_n139_), .Y(men_men_n799_));
  OAI210     u0777(.A0(men_men_n799_), .A1(men_men_n798_), .B0(men_men_n747_), .Y(men_men_n800_));
  NA4        u0778(.A(men_men_n393_), .B(men_men_n492_), .C(men_men_n71_), .D(men_men_n100_), .Y(men_men_n801_));
  INV        u0779(.A(men_men_n801_), .Y(men_men_n802_));
  NO2        u0780(.A(i_11_), .B(i_9_), .Y(men_men_n803_));
  NO2        u0781(.A(men_men_n802_), .B(men_men_n330_), .Y(men_men_n804_));
  AO210      u0782(.A0(men_men_n804_), .A1(men_men_n800_), .B0(i_12_), .Y(men_men_n805_));
  NA2        u0783(.A(men_men_n377_), .B(men_men_n337_), .Y(men_men_n806_));
  NA2        u0784(.A(men_men_n596_), .B(men_men_n63_), .Y(men_men_n807_));
  NA2        u0785(.A(men_men_n695_), .B(men_men_n71_), .Y(men_men_n808_));
  NA4        u0786(.A(men_men_n642_), .B(men_men_n808_), .C(men_men_n807_), .D(men_men_n806_), .Y(men_men_n809_));
  INV        u0787(.A(men_men_n197_), .Y(men_men_n810_));
  AOI220     u0788(.A0(men_men_n810_), .A1(men_men_n803_), .B0(men_men_n809_), .B1(men_men_n73_), .Y(men_men_n811_));
  INV        u0789(.A(men_men_n329_), .Y(men_men_n812_));
  NA2        u0790(.A(men_men_n75_), .B(men_men_n131_), .Y(men_men_n813_));
  NO2        u0791(.A(men_men_n813_), .B(men_men_n812_), .Y(men_men_n814_));
  NO2        u0792(.A(men_men_n254_), .B(i_9_), .Y(men_men_n815_));
  NA2        u0793(.A(men_men_n815_), .B(men_men_n793_), .Y(men_men_n816_));
  AOI210     u0794(.A0(men_men_n816_), .A1(men_men_n526_), .B0(men_men_n185_), .Y(men_men_n817_));
  NO2        u0795(.A(men_men_n32_), .B(i_11_), .Y(men_men_n818_));
  NA3        u0796(.A(men_men_n818_), .B(men_men_n483_), .C(men_men_n393_), .Y(men_men_n819_));
  NAi32      u0797(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n820_));
  AOI210     u0798(.A0(men_men_n730_), .A1(men_men_n86_), .B0(men_men_n820_), .Y(men_men_n821_));
  OAI210     u0799(.A0(men_men_n694_), .A1(men_men_n576_), .B0(men_men_n575_), .Y(men_men_n822_));
  NAi31      u0800(.An(men_men_n821_), .B(men_men_n822_), .C(men_men_n819_), .Y(men_men_n823_));
  OR3        u0801(.A(men_men_n823_), .B(men_men_n817_), .C(men_men_n814_), .Y(men_men_n824_));
  NO2        u0802(.A(i_11_), .B(i_2_), .Y(men_men_n825_));
  NA2        u0803(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n826_), .B(men_men_n413_), .Y(men_men_n827_));
  NA2        u0805(.A(men_men_n827_), .B(men_men_n825_), .Y(men_men_n828_));
  AO220      u0806(.A0(men_men_n362_), .A1(men_men_n353_), .B0(men_men_n401_), .B1(men_men_n613_), .Y(men_men_n829_));
  NA3        u0807(.A(men_men_n829_), .B(men_men_n257_), .C(i_7_), .Y(men_men_n830_));
  BUFFER     u0808(.A(men_men_n637_), .Y(men_men_n831_));
  NA3        u0809(.A(men_men_n831_), .B(men_men_n147_), .C(men_men_n69_), .Y(men_men_n832_));
  AO210      u0810(.A0(men_men_n500_), .A1(men_men_n762_), .B0(men_men_n36_), .Y(men_men_n833_));
  NA4        u0811(.A(men_men_n833_), .B(men_men_n832_), .C(men_men_n830_), .D(men_men_n828_), .Y(men_men_n834_));
  OAI210     u0812(.A0(men_men_n655_), .A1(i_11_), .B0(men_men_n86_), .Y(men_men_n835_));
  NA2        u0813(.A(men_men_n835_), .B(men_men_n575_), .Y(men_men_n836_));
  NA2        u0814(.A(men_men_n401_), .B(men_men_n70_), .Y(men_men_n837_));
  NA3        u0815(.A(men_men_n837_), .B(men_men_n836_), .C(men_men_n621_), .Y(men_men_n838_));
  AO210      u0816(.A0(men_men_n527_), .A1(men_men_n47_), .B0(men_men_n87_), .Y(men_men_n839_));
  NA3        u0817(.A(men_men_n839_), .B(men_men_n493_), .C(men_men_n220_), .Y(men_men_n840_));
  AOI210     u0818(.A0(men_men_n453_), .A1(men_men_n451_), .B0(men_men_n574_), .Y(men_men_n841_));
  NA2        u0819(.A(men_men_n111_), .B(men_men_n412_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n246_), .B(men_men_n47_), .Y(men_men_n843_));
  INV        u0821(.A(men_men_n603_), .Y(men_men_n844_));
  NA3        u0822(.A(men_men_n844_), .B(men_men_n329_), .C(i_7_), .Y(men_men_n845_));
  NA4        u0823(.A(men_men_n845_), .B(men_men_n842_), .C(men_men_n841_), .D(men_men_n840_), .Y(men_men_n846_));
  NO4        u0824(.A(men_men_n846_), .B(men_men_n838_), .C(men_men_n834_), .D(men_men_n824_), .Y(men_men_n847_));
  NA4        u0825(.A(men_men_n847_), .B(men_men_n811_), .C(men_men_n805_), .D(men_men_n383_), .Y(men3));
  NA2        u0826(.A(i_12_), .B(i_10_), .Y(men_men_n849_));
  NA2        u0827(.A(i_6_), .B(i_7_), .Y(men_men_n850_));
  NO2        u0828(.A(men_men_n850_), .B(i_0_), .Y(men_men_n851_));
  NO2        u0829(.A(i_11_), .B(men_men_n238_), .Y(men_men_n852_));
  OAI210     u0830(.A0(men_men_n851_), .A1(men_men_n290_), .B0(men_men_n852_), .Y(men_men_n853_));
  NO2        u0831(.A(men_men_n853_), .B(men_men_n193_), .Y(men_men_n854_));
  NO3        u0832(.A(men_men_n458_), .B(men_men_n89_), .C(men_men_n45_), .Y(men_men_n855_));
  OA210      u0833(.A0(men_men_n855_), .A1(men_men_n854_), .B0(men_men_n173_), .Y(men_men_n856_));
  NA2        u0834(.A(men_men_n621_), .B(men_men_n375_), .Y(men_men_n857_));
  NA2        u0835(.A(men_men_n857_), .B(men_men_n40_), .Y(men_men_n858_));
  NOi21      u0836(.An(men_men_n95_), .B(men_men_n771_), .Y(men_men_n859_));
  NA2        u0837(.A(men_men_n414_), .B(men_men_n46_), .Y(men_men_n860_));
  INV        u0838(.A(men_men_n859_), .Y(men_men_n861_));
  AOI210     u0839(.A0(men_men_n861_), .A1(men_men_n858_), .B0(men_men_n49_), .Y(men_men_n862_));
  NO4        u0840(.A(men_men_n380_), .B(men_men_n386_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n863_));
  NA2        u0841(.A(men_men_n185_), .B(men_men_n584_), .Y(men_men_n864_));
  NOi21      u0842(.An(men_men_n864_), .B(men_men_n863_), .Y(men_men_n865_));
  NA2        u0843(.A(men_men_n720_), .B(men_men_n687_), .Y(men_men_n866_));
  NA2        u0844(.A(men_men_n335_), .B(men_men_n441_), .Y(men_men_n867_));
  OAI220     u0845(.A0(men_men_n867_), .A1(men_men_n866_), .B0(men_men_n865_), .B1(men_men_n63_), .Y(men_men_n868_));
  NOi21      u0846(.An(i_5_), .B(i_9_), .Y(men_men_n869_));
  NA2        u0847(.A(men_men_n869_), .B(men_men_n449_), .Y(men_men_n870_));
  AOI210     u0848(.A0(men_men_n265_), .A1(men_men_n485_), .B0(men_men_n698_), .Y(men_men_n871_));
  NO3        u0849(.A(men_men_n417_), .B(men_men_n265_), .C(men_men_n73_), .Y(men_men_n872_));
  NO2        u0850(.A(men_men_n174_), .B(men_men_n148_), .Y(men_men_n873_));
  AOI210     u0851(.A0(men_men_n873_), .A1(men_men_n246_), .B0(men_men_n872_), .Y(men_men_n874_));
  OAI220     u0852(.A0(men_men_n874_), .A1(men_men_n180_), .B0(men_men_n871_), .B1(men_men_n870_), .Y(men_men_n875_));
  NO4        u0853(.A(men_men_n875_), .B(men_men_n868_), .C(men_men_n862_), .D(men_men_n856_), .Y(men_men_n876_));
  NA2        u0854(.A(men_men_n185_), .B(men_men_n24_), .Y(men_men_n877_));
  NO2        u0855(.A(men_men_n685_), .B(men_men_n610_), .Y(men_men_n878_));
  NO2        u0856(.A(men_men_n878_), .B(men_men_n877_), .Y(men_men_n879_));
  NA2        u0857(.A(men_men_n313_), .B(men_men_n129_), .Y(men_men_n880_));
  NAi21      u0858(.An(men_men_n162_), .B(men_men_n441_), .Y(men_men_n881_));
  OAI220     u0859(.A0(men_men_n881_), .A1(men_men_n843_), .B0(men_men_n880_), .B1(men_men_n404_), .Y(men_men_n882_));
  NO2        u0860(.A(men_men_n882_), .B(men_men_n879_), .Y(men_men_n883_));
  NO2        u0861(.A(men_men_n393_), .B(men_men_n294_), .Y(men_men_n884_));
  NA2        u0862(.A(men_men_n884_), .B(men_men_n723_), .Y(men_men_n885_));
  NA2        u0863(.A(men_men_n585_), .B(i_0_), .Y(men_men_n886_));
  NO3        u0864(.A(men_men_n886_), .B(men_men_n388_), .C(men_men_n88_), .Y(men_men_n887_));
  NO4        u0865(.A(men_men_n602_), .B(men_men_n217_), .C(men_men_n421_), .D(men_men_n413_), .Y(men_men_n888_));
  AOI210     u0866(.A0(men_men_n888_), .A1(i_11_), .B0(men_men_n887_), .Y(men_men_n889_));
  INV        u0867(.A(men_men_n483_), .Y(men_men_n890_));
  AN2        u0868(.A(men_men_n95_), .B(men_men_n245_), .Y(men_men_n891_));
  NA2        u0869(.A(men_men_n758_), .B(men_men_n330_), .Y(men_men_n892_));
  INV        u0870(.A(men_men_n58_), .Y(men_men_n893_));
  OAI220     u0871(.A0(men_men_n893_), .A1(men_men_n892_), .B0(men_men_n672_), .B1(men_men_n547_), .Y(men_men_n894_));
  NA2        u0872(.A(i_0_), .B(i_10_), .Y(men_men_n895_));
  OAI210     u0873(.A0(men_men_n895_), .A1(men_men_n85_), .B0(men_men_n550_), .Y(men_men_n896_));
  NO4        u0874(.A(men_men_n114_), .B(men_men_n58_), .C(men_men_n682_), .D(i_5_), .Y(men_men_n897_));
  AN2        u0875(.A(men_men_n897_), .B(men_men_n896_), .Y(men_men_n898_));
  AOI220     u0876(.A0(men_men_n335_), .A1(men_men_n97_), .B0(men_men_n185_), .B1(men_men_n84_), .Y(men_men_n899_));
  NA2        u0877(.A(men_men_n579_), .B(i_4_), .Y(men_men_n900_));
  NA2        u0878(.A(men_men_n188_), .B(men_men_n203_), .Y(men_men_n901_));
  OAI220     u0879(.A0(men_men_n901_), .A1(men_men_n892_), .B0(men_men_n900_), .B1(men_men_n899_), .Y(men_men_n902_));
  NO4        u0880(.A(men_men_n902_), .B(men_men_n898_), .C(men_men_n894_), .D(men_men_n891_), .Y(men_men_n903_));
  NA4        u0881(.A(men_men_n903_), .B(men_men_n889_), .C(men_men_n885_), .D(men_men_n883_), .Y(men_men_n904_));
  NO2        u0882(.A(men_men_n102_), .B(men_men_n37_), .Y(men_men_n905_));
  NA2        u0883(.A(i_11_), .B(i_9_), .Y(men_men_n906_));
  NO3        u0884(.A(i_12_), .B(men_men_n906_), .C(men_men_n620_), .Y(men_men_n907_));
  AO220      u0885(.A0(men_men_n907_), .A1(men_men_n905_), .B0(men_men_n267_), .B1(men_men_n87_), .Y(men_men_n908_));
  NO2        u0886(.A(men_men_n49_), .B(i_7_), .Y(men_men_n909_));
  NA2        u0887(.A(men_men_n398_), .B(men_men_n178_), .Y(men_men_n910_));
  NA2        u0888(.A(men_men_n910_), .B(men_men_n160_), .Y(men_men_n911_));
  NO2        u0889(.A(men_men_n906_), .B(men_men_n73_), .Y(men_men_n912_));
  NO2        u0890(.A(men_men_n174_), .B(i_0_), .Y(men_men_n913_));
  INV        u0891(.A(men_men_n913_), .Y(men_men_n914_));
  NA2        u0892(.A(men_men_n483_), .B(men_men_n232_), .Y(men_men_n915_));
  AOI210     u0893(.A0(men_men_n374_), .A1(men_men_n42_), .B0(men_men_n411_), .Y(men_men_n916_));
  OAI220     u0894(.A0(men_men_n916_), .A1(men_men_n870_), .B0(men_men_n915_), .B1(men_men_n914_), .Y(men_men_n917_));
  NO3        u0895(.A(men_men_n917_), .B(men_men_n911_), .C(men_men_n908_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n671_), .B(men_men_n121_), .Y(men_men_n919_));
  NO2        u0897(.A(i_6_), .B(men_men_n919_), .Y(men_men_n920_));
  AOI210     u0898(.A0(men_men_n452_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n921_));
  NA2        u0899(.A(men_men_n171_), .B(men_men_n102_), .Y(men_men_n922_));
  NOi32      u0900(.An(men_men_n921_), .Bn(men_men_n188_), .C(men_men_n922_), .Y(men_men_n923_));
  NA2        u0901(.A(men_men_n622_), .B(men_men_n330_), .Y(men_men_n924_));
  NO2        u0902(.A(men_men_n924_), .B(men_men_n860_), .Y(men_men_n925_));
  NO3        u0903(.A(men_men_n925_), .B(men_men_n923_), .C(men_men_n920_), .Y(men_men_n926_));
  NOi21      u0904(.An(i_7_), .B(i_5_), .Y(men_men_n927_));
  NOi31      u0905(.An(men_men_n927_), .B(i_0_), .C(men_men_n736_), .Y(men_men_n928_));
  NA3        u0906(.A(men_men_n928_), .B(men_men_n387_), .C(i_6_), .Y(men_men_n929_));
  OA210      u0907(.A0(men_men_n922_), .A1(men_men_n526_), .B0(men_men_n929_), .Y(men_men_n930_));
  NO3        u0908(.A(men_men_n407_), .B(men_men_n363_), .C(men_men_n361_), .Y(men_men_n931_));
  NO2        u0909(.A(men_men_n259_), .B(men_men_n320_), .Y(men_men_n932_));
  NO2        u0910(.A(men_men_n736_), .B(men_men_n258_), .Y(men_men_n933_));
  AOI210     u0911(.A0(men_men_n933_), .A1(men_men_n932_), .B0(men_men_n931_), .Y(men_men_n934_));
  NA4        u0912(.A(men_men_n934_), .B(men_men_n930_), .C(men_men_n926_), .D(men_men_n918_), .Y(men_men_n935_));
  NO2        u0913(.A(men_men_n877_), .B(men_men_n241_), .Y(men_men_n936_));
  AN2        u0914(.A(men_men_n334_), .B(men_men_n330_), .Y(men_men_n937_));
  AN2        u0915(.A(men_men_n937_), .B(men_men_n873_), .Y(men_men_n938_));
  OAI210     u0916(.A0(men_men_n938_), .A1(men_men_n936_), .B0(i_10_), .Y(men_men_n939_));
  NO2        u0917(.A(men_men_n849_), .B(men_men_n319_), .Y(men_men_n940_));
  NA2        u0918(.A(men_men_n940_), .B(men_men_n912_), .Y(men_men_n941_));
  NA3        u0919(.A(men_men_n482_), .B(men_men_n414_), .C(men_men_n46_), .Y(men_men_n942_));
  OAI210     u0920(.A0(men_men_n881_), .A1(men_men_n890_), .B0(men_men_n942_), .Y(men_men_n943_));
  NO2        u0921(.A(men_men_n257_), .B(men_men_n47_), .Y(men_men_n944_));
  NA2        u0922(.A(men_men_n912_), .B(men_men_n306_), .Y(men_men_n945_));
  OAI210     u0923(.A0(men_men_n944_), .A1(men_men_n187_), .B0(men_men_n945_), .Y(men_men_n946_));
  AOI220     u0924(.A0(men_men_n946_), .A1(men_men_n483_), .B0(men_men_n943_), .B1(men_men_n73_), .Y(men_men_n947_));
  NA3        u0925(.A(men_men_n826_), .B(men_men_n385_), .C(men_men_n655_), .Y(men_men_n948_));
  NA2        u0926(.A(men_men_n92_), .B(men_men_n45_), .Y(men_men_n949_));
  NO2        u0927(.A(men_men_n75_), .B(men_men_n760_), .Y(men_men_n950_));
  AOI220     u0928(.A0(men_men_n950_), .A1(men_men_n949_), .B0(men_men_n173_), .B1(men_men_n610_), .Y(men_men_n951_));
  AOI210     u0929(.A0(men_men_n951_), .A1(men_men_n948_), .B0(men_men_n48_), .Y(men_men_n952_));
  NO3        u0930(.A(men_men_n602_), .B(men_men_n360_), .C(men_men_n24_), .Y(men_men_n953_));
  AOI210     u0931(.A0(men_men_n714_), .A1(men_men_n559_), .B0(men_men_n953_), .Y(men_men_n954_));
  NAi21      u0932(.An(i_9_), .B(i_5_), .Y(men_men_n955_));
  NO2        u0933(.A(men_men_n955_), .B(men_men_n407_), .Y(men_men_n956_));
  NO2        u0934(.A(men_men_n616_), .B(men_men_n104_), .Y(men_men_n957_));
  AOI220     u0935(.A0(men_men_n957_), .A1(i_0_), .B0(men_men_n956_), .B1(men_men_n637_), .Y(men_men_n958_));
  OAI220     u0936(.A0(men_men_n958_), .A1(men_men_n85_), .B0(men_men_n954_), .B1(men_men_n172_), .Y(men_men_n959_));
  NO3        u0937(.A(men_men_n959_), .B(men_men_n952_), .C(men_men_n530_), .Y(men_men_n960_));
  NA4        u0938(.A(men_men_n960_), .B(men_men_n947_), .C(men_men_n941_), .D(men_men_n939_), .Y(men_men_n961_));
  NO3        u0939(.A(men_men_n961_), .B(men_men_n935_), .C(men_men_n904_), .Y(men_men_n962_));
  NO2        u0940(.A(i_0_), .B(men_men_n736_), .Y(men_men_n963_));
  NA2        u0941(.A(men_men_n73_), .B(men_men_n45_), .Y(men_men_n964_));
  NO3        u0942(.A(men_men_n104_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n965_));
  AO220      u0943(.A0(men_men_n965_), .A1(men_men_n45_), .B0(men_men_n963_), .B1(men_men_n173_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n807_), .B(men_men_n922_), .Y(men_men_n967_));
  AOI210     u0945(.A0(men_men_n966_), .A1(men_men_n350_), .B0(men_men_n967_), .Y(men_men_n968_));
  NA2        u0946(.A(men_men_n747_), .B(men_men_n146_), .Y(men_men_n969_));
  INV        u0947(.A(men_men_n969_), .Y(men_men_n970_));
  NA3        u0948(.A(men_men_n970_), .B(men_men_n687_), .C(men_men_n73_), .Y(men_men_n971_));
  NO2        u0949(.A(men_men_n822_), .B(men_men_n407_), .Y(men_men_n972_));
  NA3        u0950(.A(men_men_n851_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n973_));
  NA2        u0951(.A(men_men_n852_), .B(i_9_), .Y(men_men_n974_));
  AOI210     u0952(.A0(men_men_n973_), .A1(men_men_n505_), .B0(men_men_n974_), .Y(men_men_n975_));
  OAI210     u0953(.A0(men_men_n246_), .A1(i_9_), .B0(men_men_n231_), .Y(men_men_n976_));
  AOI210     u0954(.A0(men_men_n976_), .A1(men_men_n886_), .B0(men_men_n153_), .Y(men_men_n977_));
  NO3        u0955(.A(men_men_n977_), .B(men_men_n975_), .C(men_men_n972_), .Y(men_men_n978_));
  NA3        u0956(.A(men_men_n978_), .B(men_men_n971_), .C(men_men_n968_), .Y(men_men_n979_));
  NA2        u0957(.A(men_men_n937_), .B(men_men_n376_), .Y(men_men_n980_));
  AOI210     u0958(.A0(men_men_n301_), .A1(men_men_n162_), .B0(men_men_n980_), .Y(men_men_n981_));
  NA3        u0959(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n982_));
  NA2        u0960(.A(men_men_n909_), .B(men_men_n497_), .Y(men_men_n983_));
  AOI210     u0961(.A0(men_men_n982_), .A1(men_men_n162_), .B0(men_men_n983_), .Y(men_men_n984_));
  NO2        u0962(.A(men_men_n984_), .B(men_men_n981_), .Y(men_men_n985_));
  NA2        u0963(.A(men_men_n580_), .B(men_men_n75_), .Y(men_men_n986_));
  NO3        u0964(.A(men_men_n211_), .B(men_men_n386_), .C(i_0_), .Y(men_men_n987_));
  OAI210     u0965(.A0(men_men_n987_), .A1(men_men_n76_), .B0(i_13_), .Y(men_men_n988_));
  INV        u0966(.A(men_men_n220_), .Y(men_men_n989_));
  OAI220     u0967(.A0(men_men_n541_), .A1(men_men_n139_), .B0(i_12_), .B1(men_men_n631_), .Y(men_men_n990_));
  NA3        u0968(.A(men_men_n990_), .B(men_men_n402_), .C(men_men_n989_), .Y(men_men_n991_));
  NA4        u0969(.A(men_men_n991_), .B(men_men_n988_), .C(men_men_n986_), .D(men_men_n985_), .Y(men_men_n992_));
  NO2        u0970(.A(men_men_n244_), .B(men_men_n92_), .Y(men_men_n993_));
  AOI210     u0971(.A0(men_men_n993_), .A1(men_men_n963_), .B0(men_men_n108_), .Y(men_men_n994_));
  AOI220     u0972(.A0(men_men_n927_), .A1(men_men_n497_), .B0(men_men_n851_), .B1(men_men_n163_), .Y(men_men_n995_));
  NA2        u0973(.A(men_men_n353_), .B(men_men_n175_), .Y(men_men_n996_));
  OA220      u0974(.A0(men_men_n996_), .A1(men_men_n995_), .B0(men_men_n994_), .B1(i_5_), .Y(men_men_n997_));
  AOI210     u0975(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n174_), .Y(men_men_n998_));
  NA3        u0976(.A(men_men_n628_), .B(men_men_n185_), .C(men_men_n84_), .Y(men_men_n999_));
  NA2        u0977(.A(men_men_n999_), .B(men_men_n557_), .Y(men_men_n1000_));
  NO3        u0978(.A(men_men_n860_), .B(men_men_n55_), .C(men_men_n49_), .Y(men_men_n1001_));
  NA2        u0979(.A(men_men_n499_), .B(men_men_n496_), .Y(men_men_n1002_));
  NO3        u0980(.A(men_men_n1002_), .B(men_men_n1001_), .C(men_men_n1000_), .Y(men_men_n1003_));
  NA3        u0981(.A(men_men_n393_), .B(men_men_n171_), .C(men_men_n170_), .Y(men_men_n1004_));
  NA3        u0982(.A(men_men_n909_), .B(men_men_n290_), .C(men_men_n231_), .Y(men_men_n1005_));
  NA2        u0983(.A(men_men_n1005_), .B(men_men_n1004_), .Y(men_men_n1006_));
  NA3        u0984(.A(men_men_n393_), .B(men_men_n336_), .C(men_men_n223_), .Y(men_men_n1007_));
  INV        u0985(.A(men_men_n1007_), .Y(men_men_n1008_));
  NOi31      u0986(.An(men_men_n392_), .B(men_men_n964_), .C(men_men_n241_), .Y(men_men_n1009_));
  NO3        u0987(.A(men_men_n906_), .B(men_men_n220_), .C(men_men_n190_), .Y(men_men_n1010_));
  NO4        u0988(.A(men_men_n1010_), .B(men_men_n1009_), .C(men_men_n1008_), .D(men_men_n1006_), .Y(men_men_n1011_));
  NA3        u0989(.A(men_men_n1011_), .B(men_men_n1003_), .C(men_men_n997_), .Y(men_men_n1012_));
  INV        u0990(.A(men_men_n630_), .Y(men_men_n1013_));
  NO3        u0991(.A(men_men_n1013_), .B(men_men_n570_), .C(men_men_n347_), .Y(men_men_n1014_));
  NO2        u0992(.A(men_men_n85_), .B(i_5_), .Y(men_men_n1015_));
  NA3        u0993(.A(men_men_n852_), .B(men_men_n109_), .C(men_men_n124_), .Y(men_men_n1016_));
  INV        u0994(.A(men_men_n1016_), .Y(men_men_n1017_));
  AOI210     u0995(.A0(men_men_n1017_), .A1(men_men_n1015_), .B0(men_men_n1014_), .Y(men_men_n1018_));
  NA3        u0996(.A(men_men_n306_), .B(i_5_), .C(men_men_n193_), .Y(men_men_n1019_));
  NAi31      u0997(.An(men_men_n243_), .B(men_men_n1019_), .C(men_men_n244_), .Y(men_men_n1020_));
  NO4        u0998(.A(men_men_n241_), .B(men_men_n211_), .C(i_0_), .D(i_12_), .Y(men_men_n1021_));
  AOI220     u0999(.A0(men_men_n1021_), .A1(men_men_n1020_), .B0(men_men_n802_), .B1(men_men_n175_), .Y(men_men_n1022_));
  AN2        u1000(.A(men_men_n895_), .B(men_men_n153_), .Y(men_men_n1023_));
  NO4        u1001(.A(men_men_n1023_), .B(i_12_), .C(men_men_n661_), .D(men_men_n131_), .Y(men_men_n1024_));
  NA2        u1002(.A(men_men_n1024_), .B(men_men_n220_), .Y(men_men_n1025_));
  NA3        u1003(.A(men_men_n97_), .B(men_men_n584_), .C(i_11_), .Y(men_men_n1026_));
  NO2        u1004(.A(men_men_n1026_), .B(men_men_n155_), .Y(men_men_n1027_));
  NA2        u1005(.A(men_men_n927_), .B(men_men_n480_), .Y(men_men_n1028_));
  OAI220     u1006(.A0(i_7_), .A1(men_men_n1019_), .B0(men_men_n1028_), .B1(men_men_n688_), .Y(men_men_n1029_));
  AOI210     u1007(.A0(men_men_n1029_), .A1(men_men_n913_), .B0(men_men_n1027_), .Y(men_men_n1030_));
  NA4        u1008(.A(men_men_n1030_), .B(men_men_n1025_), .C(men_men_n1022_), .D(men_men_n1018_), .Y(men_men_n1031_));
  NO4        u1009(.A(men_men_n1031_), .B(men_men_n1012_), .C(men_men_n992_), .D(men_men_n979_), .Y(men_men_n1032_));
  NA3        u1010(.A(men_men_n921_), .B(men_men_n371_), .C(i_5_), .Y(men_men_n1033_));
  NA2        u1011(.A(men_men_n1033_), .B(men_men_n1079_), .Y(men_men_n1034_));
  NA2        u1012(.A(men_men_n1034_), .B(men_men_n207_), .Y(men_men_n1035_));
  NA2        u1013(.A(men_men_n186_), .B(men_men_n188_), .Y(men_men_n1036_));
  AO210      u1014(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n1036_), .Y(men_men_n1037_));
  OAI210     u1015(.A0(men_men_n630_), .A1(men_men_n628_), .B0(men_men_n319_), .Y(men_men_n1038_));
  NA2        u1016(.A(men_men_n1038_), .B(men_men_n1037_), .Y(men_men_n1039_));
  NO4        u1017(.A(men_men_n234_), .B(men_men_n145_), .C(men_men_n691_), .D(men_men_n37_), .Y(men_men_n1040_));
  NO2        u1018(.A(men_men_n1040_), .B(men_men_n888_), .Y(men_men_n1041_));
  OAI210     u1019(.A0(men_men_n1026_), .A1(men_men_n148_), .B0(men_men_n1041_), .Y(men_men_n1042_));
  AOI210     u1020(.A0(men_men_n1039_), .A1(men_men_n49_), .B0(men_men_n1042_), .Y(men_men_n1043_));
  AOI210     u1021(.A0(men_men_n1043_), .A1(men_men_n1035_), .B0(men_men_n73_), .Y(men_men_n1044_));
  NO2        u1022(.A(men_men_n577_), .B(men_men_n382_), .Y(men_men_n1045_));
  NO2        u1023(.A(men_men_n1045_), .B(men_men_n766_), .Y(men_men_n1046_));
  OAI210     u1024(.A0(men_men_n80_), .A1(men_men_n55_), .B0(men_men_n107_), .Y(men_men_n1047_));
  NA2        u1025(.A(men_men_n1047_), .B(men_men_n76_), .Y(men_men_n1048_));
  AOI210     u1026(.A0(men_men_n998_), .A1(men_men_n909_), .B0(men_men_n928_), .Y(men_men_n1049_));
  AOI210     u1027(.A0(men_men_n1049_), .A1(men_men_n1048_), .B0(men_men_n691_), .Y(men_men_n1050_));
  NA2        u1028(.A(men_men_n259_), .B(men_men_n57_), .Y(men_men_n1051_));
  AOI220     u1029(.A0(men_men_n1051_), .A1(men_men_n76_), .B0(men_men_n348_), .B1(men_men_n256_), .Y(men_men_n1052_));
  NO2        u1030(.A(men_men_n1052_), .B(men_men_n238_), .Y(men_men_n1053_));
  NA3        u1031(.A(men_men_n95_), .B(men_men_n308_), .C(men_men_n31_), .Y(men_men_n1054_));
  INV        u1032(.A(men_men_n1054_), .Y(men_men_n1055_));
  NO3        u1033(.A(men_men_n1055_), .B(men_men_n1053_), .C(men_men_n1050_), .Y(men_men_n1056_));
  OAI210     u1034(.A0(men_men_n267_), .A1(men_men_n158_), .B0(men_men_n88_), .Y(men_men_n1057_));
  NA3        u1035(.A(men_men_n770_), .B(men_men_n290_), .C(men_men_n80_), .Y(men_men_n1058_));
  AOI210     u1036(.A0(men_men_n1058_), .A1(men_men_n1057_), .B0(i_11_), .Y(men_men_n1059_));
  NA2        u1037(.A(men_men_n623_), .B(men_men_n217_), .Y(men_men_n1060_));
  OAI210     u1038(.A0(men_men_n1060_), .A1(men_men_n921_), .B0(men_men_n207_), .Y(men_men_n1061_));
  NA2        u1039(.A(men_men_n164_), .B(i_5_), .Y(men_men_n1062_));
  NO2        u1040(.A(men_men_n1061_), .B(men_men_n1062_), .Y(men_men_n1063_));
  NO3        u1041(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1064_));
  OAI210     u1042(.A0(men_men_n932_), .A1(men_men_n308_), .B0(men_men_n1064_), .Y(men_men_n1065_));
  NO2        u1043(.A(men_men_n1065_), .B(men_men_n736_), .Y(men_men_n1066_));
  NO4        u1044(.A(men_men_n955_), .B(men_men_n486_), .C(men_men_n255_), .D(men_men_n254_), .Y(men_men_n1067_));
  NO2        u1045(.A(men_men_n1067_), .B(men_men_n574_), .Y(men_men_n1068_));
  INV        u1046(.A(men_men_n364_), .Y(men_men_n1069_));
  AOI210     u1047(.A0(men_men_n1069_), .A1(men_men_n1068_), .B0(men_men_n41_), .Y(men_men_n1070_));
  NO4        u1048(.A(men_men_n1070_), .B(men_men_n1066_), .C(men_men_n1063_), .D(men_men_n1059_), .Y(men_men_n1071_));
  OAI210     u1049(.A0(men_men_n1056_), .A1(i_4_), .B0(men_men_n1071_), .Y(men_men_n1072_));
  NO3        u1050(.A(men_men_n1072_), .B(men_men_n1046_), .C(men_men_n1044_), .Y(men_men_n1073_));
  NA4        u1051(.A(men_men_n1073_), .B(men_men_n1032_), .C(men_men_n962_), .D(men_men_n876_), .Y(men4));
  INV        u1052(.A(i_2_), .Y(men_men_n1077_));
  INV        u1053(.A(men_men_n82_), .Y(men_men_n1078_));
  INV        u1054(.A(men_men_n161_), .Y(men_men_n1079_));
  INV        u1055(.A(men_men_n496_), .Y(men_men_n1080_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule