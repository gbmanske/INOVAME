//Benchmark atmr_intb_466_0.0313

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n331_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n381_, ori_ori_n382_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n370_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n380_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n456_, men_men_n457_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  INV        o035(.A(ori_ori_n55_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(ori_ori_n24_), .Y(ori_ori_n60_));
  NO2        o038(.A(ori_ori_n60_), .B(ori_ori_n58_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n62_));
  OAI210     o040(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n62_), .Y(ori_ori_n63_));
  AOI220     o041(.A0(ori_ori_n63_), .A1(ori_ori_n55_), .B0(ori_ori_n61_), .B1(ori_ori_n31_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(x05), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n57_), .B(ori_ori_n23_), .Y(ori_ori_n66_));
  NA2        o044(.A(x09), .B(x05), .Y(ori_ori_n67_));
  NA2        o045(.A(x10), .B(x06), .Y(ori_ori_n68_));
  NA3        o046(.A(ori_ori_n68_), .B(ori_ori_n67_), .C(ori_ori_n28_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n57_), .B(ori_ori_n41_), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n69_), .A1(ori_ori_n66_), .B0(x03), .Y(ori_ori_n71_));
  NOi31      o049(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n72_));
  INV        o050(.A(x07), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n73_), .B(ori_ori_n24_), .Y(ori_ori_n74_));
  NO2        o052(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n75_), .B(ori_ori_n36_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n75_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n77_));
  AOI210     o055(.A0(ori_ori_n76_), .A1(ori_ori_n48_), .B0(ori_ori_n77_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n79_));
  NO2        o057(.A(x08), .B(x01), .Y(ori_ori_n80_));
  OAI210     o058(.A0(ori_ori_n80_), .A1(ori_ori_n79_), .B0(ori_ori_n35_), .Y(ori_ori_n81_));
  NA2        o059(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n82_));
  NO3        o060(.A(ori_ori_n81_), .B(ori_ori_n78_), .C(ori_ori_n74_), .Y(ori_ori_n83_));
  AN2        o061(.A(ori_ori_n83_), .B(ori_ori_n71_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n81_), .Y(ori_ori_n85_));
  NA2        o063(.A(x11), .B(x00), .Y(ori_ori_n86_));
  NO2        o064(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n87_));
  NOi21      o065(.An(ori_ori_n86_), .B(ori_ori_n87_), .Y(ori_ori_n88_));
  NOi21      o066(.An(x01), .B(x10), .Y(ori_ori_n89_));
  NO2        o067(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n90_));
  NO3        o068(.A(ori_ori_n90_), .B(ori_ori_n89_), .C(x06), .Y(ori_ori_n91_));
  NA2        o069(.A(ori_ori_n91_), .B(ori_ori_n27_), .Y(ori_ori_n92_));
  OAI210     o070(.A0(ori_ori_n381_), .A1(x07), .B0(ori_ori_n92_), .Y(ori_ori_n93_));
  NO3        o071(.A(ori_ori_n93_), .B(ori_ori_n84_), .C(ori_ori_n65_), .Y(ori01));
  INV        o072(.A(x12), .Y(ori_ori_n95_));
  INV        o073(.A(x13), .Y(ori_ori_n96_));
  NA2        o074(.A(ori_ori_n89_), .B(ori_ori_n28_), .Y(ori_ori_n97_));
  NO2        o075(.A(x10), .B(x01), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n100_));
  NA2        o078(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n102_));
  NOi21      o080(.An(ori_ori_n102_), .B(ori_ori_n54_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n35_), .B(x02), .Y(ori_ori_n104_));
  INV        o082(.A(x13), .Y(ori_ori_n105_));
  NA2        o083(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n106_));
  NA2        o084(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n107_));
  NO2        o085(.A(ori_ori_n107_), .B(x05), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n35_), .B(ori_ori_n53_), .Y(ori_ori_n109_));
  INV        o087(.A(ori_ori_n103_), .Y(ori_ori_n110_));
  NO2        o088(.A(ori_ori_n110_), .B(ori_ori_n68_), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n112_));
  NA2        o090(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n113_), .B(ori_ori_n112_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n115_));
  NA2        o093(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n116_));
  NA3        o094(.A(ori_ori_n116_), .B(ori_ori_n115_), .C(x13), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n118_));
  NOi31      o096(.An(ori_ori_n117_), .B(ori_ori_n118_), .C(ori_ori_n114_), .Y(ori_ori_n119_));
  NO3        o097(.A(ori_ori_n119_), .B(x06), .C(x03), .Y(ori_ori_n120_));
  NO2        o098(.A(ori_ori_n120_), .B(ori_ori_n111_), .Y(ori_ori_n121_));
  NA2        o099(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n122_));
  OAI210     o100(.A0(ori_ori_n80_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(ori_ori_n122_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n126_));
  AOI210     o104(.A0(ori_ori_n126_), .A1(ori_ori_n49_), .B0(ori_ori_n125_), .Y(ori_ori_n127_));
  AN2        o105(.A(ori_ori_n127_), .B(ori_ori_n124_), .Y(ori_ori_n128_));
  NO2        o106(.A(x09), .B(x05), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n129_), .B(ori_ori_n47_), .Y(ori_ori_n130_));
  NO2        o108(.A(ori_ori_n100_), .B(ori_ori_n49_), .Y(ori_ori_n131_));
  NA2        o109(.A(x09), .B(x00), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n102_), .B(ori_ori_n132_), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n133_), .B(ori_ori_n126_), .Y(ori_ori_n134_));
  NO3        o112(.A(ori_ori_n134_), .B(ori_ori_n131_), .C(ori_ori_n128_), .Y(ori_ori_n135_));
  NO2        o113(.A(x03), .B(x02), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n81_), .B(ori_ori_n96_), .Y(ori_ori_n137_));
  OAI210     o115(.A0(ori_ori_n137_), .A1(ori_ori_n103_), .B0(ori_ori_n136_), .Y(ori_ori_n138_));
  OA210      o116(.A0(ori_ori_n135_), .A1(x11), .B0(ori_ori_n138_), .Y(ori_ori_n139_));
  OAI210     o117(.A0(ori_ori_n121_), .A1(ori_ori_n23_), .B0(ori_ori_n139_), .Y(ori_ori_n140_));
  NA2        o118(.A(ori_ori_n100_), .B(ori_ori_n40_), .Y(ori_ori_n141_));
  NAi21      o119(.An(x06), .B(x10), .Y(ori_ori_n142_));
  NO2        o120(.A(ori_ori_n141_), .B(ori_ori_n41_), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n144_));
  NA2        o122(.A(ori_ori_n96_), .B(x01), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n145_), .B(x08), .Y(ori_ori_n146_));
  NO2        o124(.A(ori_ori_n144_), .B(ori_ori_n48_), .Y(ori_ori_n147_));
  AOI210     o125(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n148_));
  OAI210     o126(.A0(ori_ori_n147_), .A1(ori_ori_n143_), .B0(ori_ori_n148_), .Y(ori_ori_n149_));
  NA2        o127(.A(x04), .B(x02), .Y(ori_ori_n150_));
  NA2        o128(.A(x10), .B(x05), .Y(ori_ori_n151_));
  NO2        o129(.A(x09), .B(x01), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n102_), .B(x08), .Y(ori_ori_n153_));
  INV        o131(.A(ori_ori_n25_), .Y(ori_ori_n154_));
  NAi21      o132(.An(x13), .B(x00), .Y(ori_ori_n155_));
  AN2        o133(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n90_), .B(x06), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n155_), .B(ori_ori_n36_), .Y(ori_ori_n158_));
  INV        o136(.A(ori_ori_n158_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n157_), .B(ori_ori_n156_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(ori_ori_n154_), .Y(ori_ori_n161_));
  NOi21      o139(.An(x09), .B(x00), .Y(ori_ori_n162_));
  NO3        o140(.A(ori_ori_n79_), .B(ori_ori_n162_), .C(ori_ori_n47_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n163_), .B(ori_ori_n113_), .Y(ori_ori_n164_));
  NA2        o142(.A(x06), .B(x05), .Y(ori_ori_n165_));
  OAI210     o143(.A0(ori_ori_n165_), .A1(ori_ori_n35_), .B0(ori_ori_n95_), .Y(ori_ori_n166_));
  AOI210     o144(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  NA2        o145(.A(ori_ori_n167_), .B(ori_ori_n164_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n96_), .B(x12), .Y(ori_ori_n169_));
  AOI210     o147(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n169_), .Y(ori_ori_n170_));
  NO2        o148(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n171_), .B(x02), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n170_), .B(ori_ori_n168_), .Y(ori_ori_n173_));
  NA3        o151(.A(ori_ori_n173_), .B(ori_ori_n161_), .C(ori_ori_n149_), .Y(ori_ori_n174_));
  AOI210     o152(.A0(ori_ori_n140_), .A1(ori_ori_n95_), .B0(ori_ori_n174_), .Y(ori_ori_n175_));
  INV        o153(.A(ori_ori_n69_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(ori_ori_n124_), .Y(ori_ori_n177_));
  NA2        o155(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n178_));
  NA2        o156(.A(ori_ori_n178_), .B(ori_ori_n123_), .Y(ori_ori_n179_));
  AOI210     o157(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n112_), .B(x06), .Y(ori_ori_n181_));
  AOI210     o159(.A0(ori_ori_n180_), .A1(ori_ori_n179_), .B0(ori_ori_n181_), .Y(ori_ori_n182_));
  AOI210     o160(.A0(ori_ori_n182_), .A1(ori_ori_n177_), .B0(x12), .Y(ori_ori_n183_));
  INV        o161(.A(ori_ori_n72_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n89_), .B(x06), .Y(ori_ori_n185_));
  AOI210     o163(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n50_), .Y(ori_ori_n186_));
  NO3        o164(.A(ori_ori_n186_), .B(ori_ori_n185_), .C(ori_ori_n41_), .Y(ori_ori_n187_));
  INV        o165(.A(ori_ori_n126_), .Y(ori_ori_n188_));
  OAI210     o166(.A0(ori_ori_n188_), .A1(ori_ori_n187_), .B0(x02), .Y(ori_ori_n189_));
  AOI210     o167(.A0(ori_ori_n189_), .A1(ori_ori_n53_), .B0(ori_ori_n23_), .Y(ori_ori_n190_));
  OAI210     o168(.A0(ori_ori_n183_), .A1(ori_ori_n53_), .B0(ori_ori_n190_), .Y(ori_ori_n191_));
  INV        o169(.A(ori_ori_n126_), .Y(ori_ori_n192_));
  NO2        o170(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n193_));
  OAI210     o171(.A0(ori_ori_n75_), .A1(ori_ori_n36_), .B0(ori_ori_n106_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n96_), .B(x03), .Y(ori_ori_n195_));
  AOI220     o173(.A0(ori_ori_n195_), .A1(ori_ori_n194_), .B0(ori_ori_n72_), .B1(ori_ori_n193_), .Y(ori_ori_n196_));
  NA2        o174(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n197_));
  INV        o175(.A(ori_ori_n142_), .Y(ori_ori_n198_));
  NOi21      o176(.An(x13), .B(x04), .Y(ori_ori_n199_));
  NO3        o177(.A(ori_ori_n199_), .B(ori_ori_n72_), .C(ori_ori_n162_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n200_), .B(x05), .Y(ori_ori_n201_));
  AOI220     o179(.A0(ori_ori_n201_), .A1(ori_ori_n197_), .B0(ori_ori_n198_), .B1(ori_ori_n53_), .Y(ori_ori_n202_));
  OAI210     o180(.A0(ori_ori_n196_), .A1(ori_ori_n192_), .B0(ori_ori_n202_), .Y(ori_ori_n203_));
  INV        o181(.A(ori_ori_n87_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n204_), .B(x12), .Y(ori_ori_n205_));
  NA2        o183(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n207_));
  AOI210     o185(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n208_));
  NO2        o186(.A(x06), .B(x00), .Y(ori_ori_n209_));
  NO3        o187(.A(ori_ori_n209_), .B(ori_ori_n208_), .C(ori_ori_n41_), .Y(ori_ori_n210_));
  INV        o188(.A(ori_ori_n68_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n211_), .B(ori_ori_n210_), .Y(ori_ori_n212_));
  NA2        o190(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n213_));
  NA2        o191(.A(ori_ori_n213_), .B(x03), .Y(ori_ori_n214_));
  OR2        o192(.A(ori_ori_n214_), .B(ori_ori_n212_), .Y(ori_ori_n215_));
  NA2        o193(.A(x13), .B(ori_ori_n95_), .Y(ori_ori_n216_));
  NA3        o194(.A(ori_ori_n216_), .B(ori_ori_n166_), .C(ori_ori_n88_), .Y(ori_ori_n217_));
  OAI210     o195(.A0(ori_ori_n215_), .A1(ori_ori_n206_), .B0(ori_ori_n217_), .Y(ori_ori_n218_));
  AOI210     o196(.A0(ori_ori_n205_), .A1(ori_ori_n203_), .B0(ori_ori_n218_), .Y(ori_ori_n219_));
  AOI210     o197(.A0(ori_ori_n219_), .A1(ori_ori_n191_), .B0(x07), .Y(ori_ori_n220_));
  NA2        o198(.A(ori_ori_n67_), .B(ori_ori_n29_), .Y(ori_ori_n221_));
  NOi31      o199(.An(ori_ori_n122_), .B(ori_ori_n199_), .C(ori_ori_n162_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n222_), .B(ori_ori_n221_), .Y(ori_ori_n223_));
  NO2        o201(.A(x08), .B(x05), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n224_), .B(ori_ori_n208_), .Y(ori_ori_n225_));
  OAI210     o203(.A0(ori_ori_n72_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n226_));
  INV        o204(.A(ori_ori_n226_), .Y(ori_ori_n227_));
  NO2        o205(.A(x12), .B(x02), .Y(ori_ori_n228_));
  INV        o206(.A(ori_ori_n228_), .Y(ori_ori_n229_));
  NO2        o207(.A(ori_ori_n229_), .B(ori_ori_n204_), .Y(ori_ori_n230_));
  OA210      o208(.A0(ori_ori_n227_), .A1(ori_ori_n223_), .B0(ori_ori_n230_), .Y(ori_ori_n231_));
  NA2        o209(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n232_), .B(x01), .Y(ori_ori_n233_));
  INV        o211(.A(ori_ori_n233_), .Y(ori_ori_n234_));
  AOI210     o212(.A0(ori_ori_n234_), .A1(ori_ori_n117_), .B0(ori_ori_n29_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n96_), .B(x04), .Y(ori_ori_n236_));
  NO2        o214(.A(x02), .B(ori_ori_n105_), .Y(ori_ori_n237_));
  NO3        o215(.A(ori_ori_n86_), .B(x12), .C(x03), .Y(ori_ori_n238_));
  OAI210     o216(.A0(ori_ori_n237_), .A1(ori_ori_n235_), .B0(ori_ori_n238_), .Y(ori_ori_n239_));
  NOi21      o217(.An(ori_ori_n221_), .B(ori_ori_n185_), .Y(ori_ori_n240_));
  NO2        o218(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n241_));
  NA2        o219(.A(ori_ori_n240_), .B(ori_ori_n241_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n243_));
  NO3        o221(.A(ori_ori_n243_), .B(ori_ori_n186_), .C(ori_ori_n157_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n206_), .B(ori_ori_n28_), .Y(ori_ori_n245_));
  OAI210     o223(.A0(ori_ori_n244_), .A1(ori_ori_n192_), .B0(ori_ori_n245_), .Y(ori_ori_n246_));
  NA3        o224(.A(ori_ori_n246_), .B(ori_ori_n242_), .C(ori_ori_n239_), .Y(ori_ori_n247_));
  NO3        o225(.A(ori_ori_n247_), .B(ori_ori_n231_), .C(ori_ori_n220_), .Y(ori_ori_n248_));
  OAI210     o226(.A0(ori_ori_n175_), .A1(ori_ori_n57_), .B0(ori_ori_n248_), .Y(ori02));
  AOI210     o227(.A0(ori_ori_n122_), .A1(ori_ori_n81_), .B0(ori_ori_n115_), .Y(ori_ori_n250_));
  NOi21      o228(.An(ori_ori_n200_), .B(ori_ori_n152_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n251_), .B(ori_ori_n32_), .Y(ori_ori_n252_));
  OAI210     o230(.A0(ori_ori_n252_), .A1(ori_ori_n250_), .B0(ori_ori_n151_), .Y(ori_ori_n253_));
  INV        o231(.A(ori_ori_n151_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n104_), .A1(ori_ori_n82_), .B0(ori_ori_n186_), .Y(ori_ori_n255_));
  OAI220     o233(.A0(ori_ori_n255_), .A1(ori_ori_n96_), .B0(ori_ori_n81_), .B1(ori_ori_n50_), .Y(ori_ori_n256_));
  AOI220     o234(.A0(ori_ori_n256_), .A1(ori_ori_n254_), .B0(ori_ori_n137_), .B1(ori_ori_n136_), .Y(ori_ori_n257_));
  AOI210     o235(.A0(ori_ori_n257_), .A1(ori_ori_n253_), .B0(ori_ori_n48_), .Y(ori_ori_n258_));
  NO2        o236(.A(x05), .B(x02), .Y(ori_ori_n259_));
  OAI210     o237(.A0(ori_ori_n179_), .A1(ori_ori_n162_), .B0(ori_ori_n259_), .Y(ori_ori_n260_));
  AOI220     o238(.A0(ori_ori_n224_), .A1(ori_ori_n54_), .B0(ori_ori_n52_), .B1(ori_ori_n36_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n260_), .B(ori_ori_n126_), .Y(ori_ori_n262_));
  NAi21      o240(.An(ori_ori_n201_), .B(ori_ori_n196_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n213_), .B(ori_ori_n47_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n264_), .B(ori_ori_n263_), .Y(ori_ori_n265_));
  AN2        o243(.A(ori_ori_n195_), .B(ori_ori_n194_), .Y(ori_ori_n266_));
  OAI210     o244(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n267_));
  NA2        o245(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n268_));
  OA210      o246(.A0(ori_ori_n268_), .A1(x08), .B0(ori_ori_n130_), .Y(ori_ori_n269_));
  AOI210     o247(.A0(ori_ori_n269_), .A1(ori_ori_n123_), .B0(ori_ori_n267_), .Y(ori_ori_n270_));
  OAI210     o248(.A0(ori_ori_n270_), .A1(ori_ori_n266_), .B0(ori_ori_n90_), .Y(ori_ori_n271_));
  INV        o249(.A(ori_ori_n136_), .Y(ori_ori_n272_));
  OAI220     o250(.A0(ori_ori_n225_), .A1(ori_ori_n97_), .B0(ori_ori_n272_), .B1(ori_ori_n114_), .Y(ori_ori_n273_));
  NA2        o251(.A(ori_ori_n273_), .B(x13), .Y(ori_ori_n274_));
  NA3        o252(.A(ori_ori_n274_), .B(ori_ori_n271_), .C(ori_ori_n265_), .Y(ori_ori_n275_));
  NO3        o253(.A(ori_ori_n275_), .B(ori_ori_n262_), .C(ori_ori_n258_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n125_), .B(x03), .Y(ori_ori_n277_));
  INV        o255(.A(ori_ori_n155_), .Y(ori_ori_n278_));
  AOI220     o256(.A0(x08), .A1(ori_ori_n278_), .B0(ori_ori_n171_), .B1(x08), .Y(ori_ori_n279_));
  OAI210     o257(.A0(ori_ori_n279_), .A1(ori_ori_n243_), .B0(ori_ori_n277_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n280_), .B(ori_ori_n98_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n150_), .B(ori_ori_n145_), .Y(ori_ori_n282_));
  AN2        o260(.A(ori_ori_n282_), .B(ori_ori_n153_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n115_), .B(ori_ori_n28_), .Y(ori_ori_n284_));
  OAI210     o262(.A0(ori_ori_n284_), .A1(ori_ori_n283_), .B0(ori_ori_n99_), .Y(ori_ori_n285_));
  NA2        o263(.A(ori_ori_n236_), .B(ori_ori_n95_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n95_), .B(ori_ori_n41_), .Y(ori_ori_n287_));
  NA3        o265(.A(ori_ori_n287_), .B(ori_ori_n286_), .C(ori_ori_n114_), .Y(ori_ori_n288_));
  NA4        o266(.A(ori_ori_n288_), .B(ori_ori_n285_), .C(ori_ori_n281_), .D(ori_ori_n48_), .Y(ori_ori_n289_));
  INV        o267(.A(ori_ori_n171_), .Y(ori_ori_n290_));
  NA2        o268(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n291_));
  OAI220     o269(.A0(ori_ori_n291_), .A1(ori_ori_n382_), .B0(ori_ori_n290_), .B1(ori_ori_n55_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n292_), .B(x02), .Y(ori_ori_n293_));
  INV        o271(.A(ori_ori_n207_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n169_), .B(x04), .Y(ori_ori_n295_));
  NO3        o273(.A(ori_ori_n169_), .B(ori_ori_n144_), .C(ori_ori_n51_), .Y(ori_ori_n296_));
  OAI210     o274(.A0(ori_ori_n132_), .A1(ori_ori_n36_), .B0(ori_ori_n95_), .Y(ori_ori_n297_));
  OAI210     o275(.A0(ori_ori_n297_), .A1(ori_ori_n163_), .B0(ori_ori_n296_), .Y(ori_ori_n298_));
  NA3        o276(.A(ori_ori_n298_), .B(ori_ori_n293_), .C(x06), .Y(ori_ori_n299_));
  NA2        o277(.A(x09), .B(x03), .Y(ori_ori_n300_));
  OAI220     o278(.A0(ori_ori_n300_), .A1(ori_ori_n113_), .B0(ori_ori_n178_), .B1(ori_ori_n59_), .Y(ori_ori_n301_));
  NO3        o279(.A(ori_ori_n243_), .B(ori_ori_n112_), .C(x08), .Y(ori_ori_n302_));
  INV        o280(.A(ori_ori_n302_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n304_));
  NO3        o282(.A(ori_ori_n102_), .B(ori_ori_n113_), .C(ori_ori_n38_), .Y(ori_ori_n305_));
  AOI210     o283(.A0(ori_ori_n296_), .A1(ori_ori_n304_), .B0(ori_ori_n305_), .Y(ori_ori_n306_));
  OAI210     o284(.A0(ori_ori_n303_), .A1(ori_ori_n28_), .B0(ori_ori_n306_), .Y(ori_ori_n307_));
  AO220      o285(.A0(ori_ori_n307_), .A1(x04), .B0(ori_ori_n301_), .B1(x05), .Y(ori_ori_n308_));
  AOI210     o286(.A0(ori_ori_n299_), .A1(ori_ori_n289_), .B0(ori_ori_n308_), .Y(ori_ori_n309_));
  OAI210     o287(.A0(ori_ori_n276_), .A1(x12), .B0(ori_ori_n309_), .Y(ori03));
  OR2        o288(.A(ori_ori_n42_), .B(ori_ori_n193_), .Y(ori_ori_n311_));
  AOI210     o289(.A0(ori_ori_n137_), .A1(ori_ori_n95_), .B0(ori_ori_n311_), .Y(ori_ori_n312_));
  AO210      o290(.A0(ori_ori_n294_), .A1(ori_ori_n82_), .B0(ori_ori_n295_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n169_), .B(ori_ori_n136_), .Y(ori_ori_n314_));
  NA3        o292(.A(ori_ori_n314_), .B(ori_ori_n313_), .C(ori_ori_n172_), .Y(ori_ori_n315_));
  OAI210     o293(.A0(ori_ori_n315_), .A1(ori_ori_n312_), .B0(x05), .Y(ori_ori_n316_));
  NA2        o294(.A(ori_ori_n311_), .B(x05), .Y(ori_ori_n317_));
  AOI210     o295(.A0(ori_ori_n123_), .A1(ori_ori_n184_), .B0(ori_ori_n317_), .Y(ori_ori_n318_));
  AOI210     o296(.A0(ori_ori_n195_), .A1(ori_ori_n76_), .B0(ori_ori_n108_), .Y(ori_ori_n319_));
  OAI220     o297(.A0(ori_ori_n319_), .A1(ori_ori_n55_), .B0(ori_ori_n268_), .B1(ori_ori_n261_), .Y(ori_ori_n320_));
  OAI210     o298(.A0(ori_ori_n320_), .A1(ori_ori_n318_), .B0(ori_ori_n95_), .Y(ori_ori_n321_));
  AOI210     o299(.A0(ori_ori_n130_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n152_), .B(ori_ori_n118_), .Y(ori_ori_n323_));
  OAI220     o301(.A0(ori_ori_n323_), .A1(ori_ori_n37_), .B0(ori_ori_n133_), .B1(x13), .Y(ori_ori_n324_));
  OAI210     o302(.A0(ori_ori_n324_), .A1(ori_ori_n322_), .B0(x04), .Y(ori_ori_n325_));
  NO3        o303(.A(ori_ori_n287_), .B(ori_ori_n81_), .C(ori_ori_n55_), .Y(ori_ori_n326_));
  AOI210     o304(.A0(ori_ori_n159_), .A1(ori_ori_n95_), .B0(ori_ori_n130_), .Y(ori_ori_n327_));
  OA210      o305(.A0(ori_ori_n146_), .A1(x12), .B0(ori_ori_n118_), .Y(ori_ori_n328_));
  NO3        o306(.A(ori_ori_n328_), .B(ori_ori_n327_), .C(ori_ori_n326_), .Y(ori_ori_n329_));
  NA4        o307(.A(ori_ori_n329_), .B(ori_ori_n325_), .C(ori_ori_n321_), .D(ori_ori_n316_), .Y(ori04));
  NO2        o308(.A(ori_ori_n85_), .B(ori_ori_n39_), .Y(ori_ori_n331_));
  XO2        o309(.A(ori_ori_n331_), .B(ori_ori_n216_), .Y(ori05));
  NO2        o310(.A(ori_ori_n51_), .B(ori_ori_n181_), .Y(ori_ori_n333_));
  AOI210     o311(.A0(ori_ori_n333_), .A1(ori_ori_n267_), .B0(ori_ori_n25_), .Y(ori_ori_n334_));
  NO2        o312(.A(x06), .B(ori_ori_n24_), .Y(ori_ori_n335_));
  OAI210     o313(.A0(ori_ori_n335_), .A1(ori_ori_n334_), .B0(ori_ori_n95_), .Y(ori_ori_n336_));
  OAI210     o314(.A0(ori_ori_n26_), .A1(ori_ori_n95_), .B0(x07), .Y(ori_ori_n337_));
  INV        o315(.A(ori_ori_n337_), .Y(ori_ori_n338_));
  AOI210     o316(.A0(ori_ori_n77_), .A1(ori_ori_n31_), .B0(ori_ori_n51_), .Y(ori_ori_n339_));
  NO3        o317(.A(ori_ori_n339_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n209_), .B(ori_ori_n204_), .Y(ori_ori_n341_));
  NA2        o319(.A(ori_ori_n341_), .B(ori_ori_n206_), .Y(ori_ori_n342_));
  OAI210     o320(.A0(ori_ori_n342_), .A1(ori_ori_n340_), .B0(ori_ori_n95_), .Y(ori_ori_n343_));
  NA2        o321(.A(ori_ori_n33_), .B(ori_ori_n95_), .Y(ori_ori_n344_));
  AOI210     o322(.A0(ori_ori_n344_), .A1(ori_ori_n87_), .B0(x07), .Y(ori_ori_n345_));
  AOI220     o323(.A0(ori_ori_n345_), .A1(ori_ori_n343_), .B0(ori_ori_n338_), .B1(ori_ori_n336_), .Y(ori_ori_n346_));
  OR2        o324(.A(ori_ori_n232_), .B(ori_ori_n229_), .Y(ori_ori_n347_));
  NO2        o325(.A(ori_ori_n129_), .B(ori_ori_n28_), .Y(ori_ori_n348_));
  AOI210     o326(.A0(ori_ori_n347_), .A1(ori_ori_n47_), .B0(ori_ori_n348_), .Y(ori_ori_n349_));
  NA2        o327(.A(ori_ori_n349_), .B(ori_ori_n96_), .Y(ori_ori_n350_));
  AOI210     o328(.A0(ori_ori_n295_), .A1(ori_ori_n101_), .B0(ori_ori_n228_), .Y(ori_ori_n351_));
  NOi21      o329(.An(ori_ori_n277_), .B(ori_ori_n118_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n352_), .B(ori_ori_n229_), .Y(ori_ori_n353_));
  OAI210     o331(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n354_));
  AOI210     o332(.A0(ori_ori_n216_), .A1(ori_ori_n47_), .B0(ori_ori_n354_), .Y(ori_ori_n355_));
  NO4        o333(.A(ori_ori_n355_), .B(ori_ori_n353_), .C(ori_ori_n351_), .D(x08), .Y(ori_ori_n356_));
  NO2        o334(.A(ori_ori_n115_), .B(ori_ori_n28_), .Y(ori_ori_n357_));
  NO2        o335(.A(ori_ori_n357_), .B(ori_ori_n233_), .Y(ori_ori_n358_));
  OR3        o336(.A(ori_ori_n358_), .B(x12), .C(x03), .Y(ori_ori_n359_));
  NA3        o337(.A(ori_ori_n290_), .B(ori_ori_n109_), .C(x12), .Y(ori_ori_n360_));
  AO210      o338(.A0(ori_ori_n290_), .A1(ori_ori_n109_), .B0(ori_ori_n216_), .Y(ori_ori_n361_));
  NA4        o339(.A(ori_ori_n361_), .B(ori_ori_n360_), .C(ori_ori_n359_), .D(x08), .Y(ori_ori_n362_));
  INV        o340(.A(ori_ori_n362_), .Y(ori_ori_n363_));
  AOI210     o341(.A0(ori_ori_n356_), .A1(ori_ori_n350_), .B0(ori_ori_n363_), .Y(ori_ori_n364_));
  INV        o342(.A(x03), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n129_), .B(ori_ori_n43_), .Y(ori_ori_n366_));
  OAI210     o344(.A0(ori_ori_n366_), .A1(ori_ori_n365_), .B0(ori_ori_n158_), .Y(ori_ori_n367_));
  NA3        o345(.A(ori_ori_n358_), .B(ori_ori_n352_), .C(ori_ori_n286_), .Y(ori_ori_n368_));
  INV        o346(.A(x14), .Y(ori_ori_n369_));
  NO3        o347(.A(ori_ori_n145_), .B(ori_ori_n70_), .C(ori_ori_n53_), .Y(ori_ori_n370_));
  NO2        o348(.A(ori_ori_n370_), .B(ori_ori_n369_), .Y(ori_ori_n371_));
  NA3        o349(.A(ori_ori_n371_), .B(ori_ori_n368_), .C(ori_ori_n367_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n344_), .B(ori_ori_n57_), .Y(ori_ori_n373_));
  NOi21      o351(.An(ori_ori_n236_), .B(ori_ori_n133_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n44_), .B(x04), .Y(ori_ori_n375_));
  OAI210     o353(.A0(ori_ori_n375_), .A1(ori_ori_n374_), .B0(ori_ori_n95_), .Y(ori_ori_n376_));
  OAI210     o354(.A0(ori_ori_n373_), .A1(ori_ori_n86_), .B0(ori_ori_n376_), .Y(ori_ori_n377_));
  NO4        o355(.A(ori_ori_n377_), .B(ori_ori_n372_), .C(ori_ori_n364_), .D(ori_ori_n346_), .Y(ori06));
  INV        o356(.A(ori_ori_n88_), .Y(ori_ori_n381_));
  INV        o357(.A(ori_ori_n40_), .Y(ori_ori_n382_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x09), .B(x05), .Y(mai_mai_n71_));
  NA2        m049(.A(x10), .B(x06), .Y(mai_mai_n72_));
  NA2        m050(.A(mai_mai_n72_), .B(mai_mai_n71_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n73_), .A1(x11), .B0(x03), .Y(mai_mai_n74_));
  NOi31      m052(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n75_));
  INV        m053(.A(mai_mai_n24_), .Y(mai_mai_n76_));
  NO2        m054(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n77_), .B(mai_mai_n36_), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n77_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n79_));
  INV        m057(.A(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m058(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n81_));
  NO2        m059(.A(x08), .B(x01), .Y(mai_mai_n82_));
  OAI210     m060(.A0(mai_mai_n82_), .A1(mai_mai_n81_), .B0(mai_mai_n35_), .Y(mai_mai_n83_));
  NA2        m061(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n84_));
  NO3        m062(.A(mai_mai_n83_), .B(mai_mai_n80_), .C(mai_mai_n76_), .Y(mai_mai_n85_));
  AN2        m063(.A(mai_mai_n85_), .B(mai_mai_n74_), .Y(mai_mai_n86_));
  INV        m064(.A(mai_mai_n83_), .Y(mai_mai_n87_));
  NO2        m065(.A(x06), .B(x05), .Y(mai_mai_n88_));
  NA2        m066(.A(x11), .B(x00), .Y(mai_mai_n89_));
  NO2        m067(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n90_));
  NOi21      m068(.An(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  AOI210     m069(.A0(mai_mai_n88_), .A1(mai_mai_n87_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NOi21      m070(.An(x01), .B(x10), .Y(mai_mai_n93_));
  NO2        m071(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n94_));
  NO3        m072(.A(mai_mai_n94_), .B(mai_mai_n93_), .C(x06), .Y(mai_mai_n95_));
  NA2        m073(.A(mai_mai_n95_), .B(mai_mai_n27_), .Y(mai_mai_n96_));
  OAI210     m074(.A0(mai_mai_n92_), .A1(x07), .B0(mai_mai_n96_), .Y(mai_mai_n97_));
  NO3        m075(.A(mai_mai_n97_), .B(mai_mai_n86_), .C(mai_mai_n70_), .Y(mai01));
  INV        m076(.A(x12), .Y(mai_mai_n99_));
  INV        m077(.A(x13), .Y(mai_mai_n100_));
  NA2        m078(.A(x08), .B(x04), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n101_), .B(mai_mai_n57_), .Y(mai_mai_n102_));
  NA2        m080(.A(mai_mai_n102_), .B(mai_mai_n88_), .Y(mai_mai_n103_));
  NA2        m081(.A(mai_mai_n93_), .B(mai_mai_n28_), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n104_), .B(mai_mai_n71_), .Y(mai_mai_n105_));
  NO2        m083(.A(x10), .B(x01), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n107_), .B(mai_mai_n106_), .Y(mai_mai_n108_));
  NA2        m086(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n109_));
  NO3        m087(.A(mai_mai_n109_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n110_));
  AOI210     m088(.A0(mai_mai_n110_), .A1(mai_mai_n108_), .B0(mai_mai_n105_), .Y(mai_mai_n111_));
  AOI210     m089(.A0(mai_mai_n111_), .A1(mai_mai_n103_), .B0(mai_mai_n100_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n113_));
  NOi21      m091(.An(mai_mai_n113_), .B(mai_mai_n58_), .Y(mai_mai_n114_));
  NA3        m092(.A(x13), .B(mai_mai_n436_), .C(x06), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n82_), .B(x13), .Y(mai_mai_n117_));
  NA2        m095(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n118_), .B(mai_mai_n117_), .Y(mai_mai_n119_));
  NA2        m097(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n120_), .B(x05), .Y(mai_mai_n121_));
  NO2        m099(.A(mai_mai_n121_), .B(mai_mai_n119_), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n123_));
  AOI210     m101(.A0(mai_mai_n57_), .A1(mai_mai_n78_), .B0(mai_mai_n114_), .Y(mai_mai_n124_));
  AOI210     m102(.A0(mai_mai_n124_), .A1(mai_mai_n122_), .B0(mai_mai_n72_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n126_));
  NA2        m104(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n129_));
  NO3        m107(.A(mai_mai_n123_), .B(mai_mai_n77_), .C(mai_mai_n36_), .Y(mai_mai_n130_));
  NO2        m108(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n131_));
  NO3        m109(.A(mai_mai_n131_), .B(mai_mai_n130_), .C(mai_mai_n128_), .Y(mai_mai_n132_));
  NO3        m110(.A(mai_mai_n132_), .B(x06), .C(x03), .Y(mai_mai_n133_));
  NO4        m111(.A(mai_mai_n133_), .B(mai_mai_n125_), .C(mai_mai_n116_), .D(mai_mai_n112_), .Y(mai_mai_n134_));
  OAI210     m112(.A0(mai_mai_n82_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n135_));
  NO2        m113(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n137_));
  NO2        m115(.A(x09), .B(x05), .Y(mai_mai_n138_));
  NA2        m116(.A(mai_mai_n138_), .B(mai_mai_n47_), .Y(mai_mai_n139_));
  AOI210     m117(.A0(mai_mai_n139_), .A1(mai_mai_n108_), .B0(mai_mai_n49_), .Y(mai_mai_n140_));
  NA2        m118(.A(x09), .B(x00), .Y(mai_mai_n141_));
  NA2        m119(.A(mai_mai_n113_), .B(mai_mai_n141_), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n75_), .B(mai_mai_n51_), .Y(mai_mai_n143_));
  AOI210     m121(.A0(mai_mai_n143_), .A1(mai_mai_n142_), .B0(mai_mai_n137_), .Y(mai_mai_n144_));
  NO2        m122(.A(mai_mai_n144_), .B(mai_mai_n140_), .Y(mai_mai_n145_));
  NO2        m123(.A(x03), .B(x02), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n83_), .B(mai_mai_n100_), .Y(mai_mai_n147_));
  OAI210     m125(.A0(mai_mai_n147_), .A1(mai_mai_n114_), .B0(mai_mai_n146_), .Y(mai_mai_n148_));
  OA210      m126(.A0(mai_mai_n145_), .A1(x11), .B0(mai_mai_n148_), .Y(mai_mai_n149_));
  OAI210     m127(.A0(mai_mai_n134_), .A1(mai_mai_n23_), .B0(mai_mai_n149_), .Y(mai_mai_n150_));
  NA2        m128(.A(mai_mai_n108_), .B(mai_mai_n40_), .Y(mai_mai_n151_));
  NAi21      m129(.An(x06), .B(x10), .Y(mai_mai_n152_));
  NOi21      m130(.An(x01), .B(x13), .Y(mai_mai_n153_));
  NA2        m131(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  BUFFER     m132(.A(mai_mai_n154_), .Y(mai_mai_n155_));
  AOI210     m133(.A0(mai_mai_n155_), .A1(mai_mai_n151_), .B0(mai_mai_n41_), .Y(mai_mai_n156_));
  NO2        m134(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n157_));
  NA2        m135(.A(mai_mai_n100_), .B(x01), .Y(mai_mai_n158_));
  NO2        m136(.A(mai_mai_n158_), .B(x08), .Y(mai_mai_n159_));
  OAI210     m137(.A0(x05), .A1(mai_mai_n159_), .B0(mai_mai_n51_), .Y(mai_mai_n160_));
  AOI210     m138(.A0(mai_mai_n160_), .A1(mai_mai_n157_), .B0(mai_mai_n48_), .Y(mai_mai_n161_));
  AOI210     m139(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n162_));
  OAI210     m140(.A0(mai_mai_n161_), .A1(mai_mai_n156_), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  NA2        m141(.A(x04), .B(x02), .Y(mai_mai_n164_));
  NA2        m142(.A(x10), .B(x05), .Y(mai_mai_n165_));
  INV        m143(.A(x06), .Y(mai_mai_n166_));
  NO2        m144(.A(x09), .B(x01), .Y(mai_mai_n167_));
  NO3        m145(.A(mai_mai_n167_), .B(mai_mai_n106_), .C(mai_mai_n31_), .Y(mai_mai_n168_));
  NA2        m146(.A(mai_mai_n168_), .B(x00), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n113_), .B(x08), .Y(mai_mai_n170_));
  OAI210     m148(.A0(mai_mai_n435_), .A1(x11), .B0(mai_mai_n169_), .Y(mai_mai_n171_));
  NAi21      m149(.An(mai_mai_n164_), .B(mai_mai_n171_), .Y(mai_mai_n172_));
  INV        m150(.A(mai_mai_n25_), .Y(mai_mai_n173_));
  NAi21      m151(.An(x13), .B(x00), .Y(mai_mai_n174_));
  AOI210     m152(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n174_), .Y(mai_mai_n175_));
  AOI220     m153(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n176_));
  OAI210     m154(.A0(mai_mai_n165_), .A1(mai_mai_n35_), .B0(mai_mai_n176_), .Y(mai_mai_n177_));
  AN2        m155(.A(mai_mai_n177_), .B(mai_mai_n175_), .Y(mai_mai_n178_));
  NO2        m156(.A(mai_mai_n174_), .B(mai_mai_n36_), .Y(mai_mai_n179_));
  INV        m157(.A(mai_mai_n179_), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n180_), .B(mai_mai_n166_), .Y(mai_mai_n181_));
  OAI210     m159(.A0(mai_mai_n181_), .A1(mai_mai_n178_), .B0(mai_mai_n173_), .Y(mai_mai_n182_));
  NOi21      m160(.An(x09), .B(x00), .Y(mai_mai_n183_));
  NO3        m161(.A(mai_mai_n81_), .B(mai_mai_n183_), .C(mai_mai_n47_), .Y(mai_mai_n184_));
  NA2        m162(.A(mai_mai_n184_), .B(mai_mai_n127_), .Y(mai_mai_n185_));
  NA2        m163(.A(x10), .B(x08), .Y(mai_mai_n186_));
  INV        m164(.A(mai_mai_n186_), .Y(mai_mai_n187_));
  NA2        m165(.A(x06), .B(x05), .Y(mai_mai_n188_));
  OAI210     m166(.A0(mai_mai_n188_), .A1(mai_mai_n35_), .B0(mai_mai_n99_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n99_), .B(mai_mai_n185_), .Y(mai_mai_n190_));
  NO2        m168(.A(mai_mai_n100_), .B(x12), .Y(mai_mai_n191_));
  AOI210     m169(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n191_), .Y(mai_mai_n192_));
  NA2        m170(.A(mai_mai_n93_), .B(mai_mai_n51_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n194_), .B(x02), .Y(mai_mai_n195_));
  NO2        m173(.A(mai_mai_n195_), .B(mai_mai_n193_), .Y(mai_mai_n196_));
  AOI210     m174(.A0(mai_mai_n192_), .A1(mai_mai_n190_), .B0(mai_mai_n196_), .Y(mai_mai_n197_));
  NA4        m175(.A(mai_mai_n197_), .B(mai_mai_n182_), .C(mai_mai_n172_), .D(mai_mai_n163_), .Y(mai_mai_n198_));
  AOI210     m176(.A0(mai_mai_n150_), .A1(mai_mai_n99_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  NA2        m177(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n200_), .B(mai_mai_n135_), .Y(mai_mai_n201_));
  AOI210     m179(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n126_), .B(x06), .Y(mai_mai_n203_));
  AOI210     m181(.A0(mai_mai_n202_), .A1(mai_mai_n201_), .B0(mai_mai_n203_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n204_), .B(x12), .Y(mai_mai_n205_));
  INV        m183(.A(mai_mai_n75_), .Y(mai_mai_n206_));
  NO2        m184(.A(x05), .B(mai_mai_n51_), .Y(mai_mai_n207_));
  OAI210     m185(.A0(mai_mai_n207_), .A1(mai_mai_n154_), .B0(mai_mai_n57_), .Y(mai_mai_n208_));
  NA2        m186(.A(mai_mai_n208_), .B(mai_mai_n206_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n93_), .B(x06), .Y(mai_mai_n210_));
  NA4        m188(.A(mai_mai_n152_), .B(mai_mai_n56_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n211_));
  NA2        m189(.A(mai_mai_n211_), .B(mai_mai_n137_), .Y(mai_mai_n212_));
  NA2        m190(.A(mai_mai_n212_), .B(x02), .Y(mai_mai_n213_));
  AOI210     m191(.A0(mai_mai_n213_), .A1(mai_mai_n209_), .B0(mai_mai_n23_), .Y(mai_mai_n214_));
  OAI210     m192(.A0(mai_mai_n205_), .A1(mai_mai_n57_), .B0(mai_mai_n214_), .Y(mai_mai_n215_));
  INV        m193(.A(mai_mai_n137_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n217_));
  OAI210     m195(.A0(mai_mai_n77_), .A1(mai_mai_n36_), .B0(mai_mai_n118_), .Y(mai_mai_n218_));
  NO2        m196(.A(mai_mai_n100_), .B(x03), .Y(mai_mai_n219_));
  NA2        m197(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n220_));
  NA2        m198(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n221_));
  INV        m199(.A(mai_mai_n152_), .Y(mai_mai_n222_));
  NOi21      m200(.An(x13), .B(x04), .Y(mai_mai_n223_));
  NO3        m201(.A(mai_mai_n223_), .B(mai_mai_n75_), .C(mai_mai_n183_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n224_), .B(x05), .Y(mai_mai_n225_));
  AOI220     m203(.A0(mai_mai_n225_), .A1(mai_mai_n221_), .B0(mai_mai_n222_), .B1(mai_mai_n57_), .Y(mai_mai_n226_));
  OAI210     m204(.A0(mai_mai_n220_), .A1(mai_mai_n216_), .B0(mai_mai_n226_), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n90_), .Y(mai_mai_n228_));
  NO2        m206(.A(mai_mai_n228_), .B(x12), .Y(mai_mai_n229_));
  NA2        m207(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n231_));
  OAI210     m209(.A0(mai_mai_n231_), .A1(mai_mai_n177_), .B0(mai_mai_n175_), .Y(mai_mai_n232_));
  AOI210     m210(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n233_));
  NO2        m211(.A(x06), .B(x00), .Y(mai_mai_n234_));
  NO3        m212(.A(mai_mai_n234_), .B(mai_mai_n233_), .C(mai_mai_n41_), .Y(mai_mai_n235_));
  OAI210     m213(.A0(mai_mai_n101_), .A1(mai_mai_n141_), .B0(mai_mai_n72_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n236_), .B(mai_mai_n235_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n238_), .B(x03), .Y(mai_mai_n239_));
  OA210      m217(.A0(mai_mai_n239_), .A1(mai_mai_n237_), .B0(mai_mai_n232_), .Y(mai_mai_n240_));
  NA2        m218(.A(x13), .B(mai_mai_n99_), .Y(mai_mai_n241_));
  NA3        m219(.A(mai_mai_n241_), .B(mai_mai_n189_), .C(mai_mai_n91_), .Y(mai_mai_n242_));
  OAI210     m220(.A0(mai_mai_n240_), .A1(mai_mai_n230_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  AOI210     m221(.A0(mai_mai_n229_), .A1(mai_mai_n227_), .B0(mai_mai_n243_), .Y(mai_mai_n244_));
  AOI210     m222(.A0(mai_mai_n244_), .A1(mai_mai_n215_), .B0(x07), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n71_), .B(mai_mai_n29_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n223_), .B(mai_mai_n183_), .Y(mai_mai_n247_));
  AOI210     m225(.A0(mai_mai_n247_), .A1(mai_mai_n143_), .B0(mai_mai_n246_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n100_), .B(x06), .Y(mai_mai_n249_));
  INV        m227(.A(mai_mai_n249_), .Y(mai_mai_n250_));
  NO2        m228(.A(x08), .B(x05), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n251_), .B(mai_mai_n233_), .Y(mai_mai_n252_));
  NA2        m230(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n253_));
  OAI210     m231(.A0(mai_mai_n252_), .A1(mai_mai_n250_), .B0(mai_mai_n253_), .Y(mai_mai_n254_));
  NO2        m232(.A(x12), .B(x02), .Y(mai_mai_n255_));
  INV        m233(.A(mai_mai_n255_), .Y(mai_mai_n256_));
  NO2        m234(.A(mai_mai_n256_), .B(mai_mai_n228_), .Y(mai_mai_n257_));
  OA210      m235(.A0(mai_mai_n254_), .A1(mai_mai_n248_), .B0(mai_mai_n257_), .Y(mai_mai_n258_));
  NA2        m236(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n259_));
  NO2        m237(.A(mai_mai_n259_), .B(x01), .Y(mai_mai_n260_));
  NOi21      m238(.An(mai_mai_n82_), .B(mai_mai_n118_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n261_), .B(mai_mai_n260_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n262_), .B(mai_mai_n29_), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n249_), .B(mai_mai_n218_), .Y(mai_mai_n264_));
  NA2        m242(.A(mai_mai_n100_), .B(x04), .Y(mai_mai_n265_));
  NA2        m243(.A(mai_mai_n265_), .B(mai_mai_n28_), .Y(mai_mai_n266_));
  OAI210     m244(.A0(mai_mai_n266_), .A1(mai_mai_n117_), .B0(mai_mai_n264_), .Y(mai_mai_n267_));
  NO3        m245(.A(mai_mai_n89_), .B(x12), .C(x03), .Y(mai_mai_n268_));
  OAI210     m246(.A0(mai_mai_n267_), .A1(mai_mai_n263_), .B0(mai_mai_n268_), .Y(mai_mai_n269_));
  AOI210     m247(.A0(mai_mai_n193_), .A1(mai_mai_n188_), .B0(mai_mai_n101_), .Y(mai_mai_n270_));
  NOi21      m248(.An(mai_mai_n246_), .B(mai_mai_n210_), .Y(mai_mai_n271_));
  NO2        m249(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n272_));
  OAI210     m250(.A0(mai_mai_n271_), .A1(mai_mai_n270_), .B0(mai_mai_n272_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n230_), .B(mai_mai_n28_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n216_), .B(mai_mai_n275_), .Y(mai_mai_n276_));
  NA3        m254(.A(mai_mai_n276_), .B(mai_mai_n273_), .C(mai_mai_n269_), .Y(mai_mai_n277_));
  NO3        m255(.A(mai_mai_n277_), .B(mai_mai_n258_), .C(mai_mai_n245_), .Y(mai_mai_n278_));
  OAI210     m256(.A0(mai_mai_n199_), .A1(mai_mai_n61_), .B0(mai_mai_n278_), .Y(mai02));
  NOi21      m257(.An(mai_mai_n224_), .B(mai_mai_n167_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n100_), .B(mai_mai_n35_), .Y(mai_mai_n281_));
  NA3        m259(.A(mai_mai_n281_), .B(mai_mai_n187_), .C(mai_mai_n56_), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n280_), .A1(mai_mai_n32_), .B0(mai_mai_n282_), .Y(mai_mai_n283_));
  NA2        m261(.A(mai_mai_n283_), .B(mai_mai_n165_), .Y(mai_mai_n284_));
  INV        m262(.A(mai_mai_n165_), .Y(mai_mai_n285_));
  OAI220     m263(.A0(mai_mai_n51_), .A1(mai_mai_n100_), .B0(mai_mai_n83_), .B1(mai_mai_n51_), .Y(mai_mai_n286_));
  AOI220     m264(.A0(mai_mai_n286_), .A1(mai_mai_n285_), .B0(mai_mai_n147_), .B1(mai_mai_n146_), .Y(mai_mai_n287_));
  AOI210     m265(.A0(mai_mai_n287_), .A1(mai_mai_n284_), .B0(mai_mai_n48_), .Y(mai_mai_n288_));
  NO2        m266(.A(x05), .B(x02), .Y(mai_mai_n289_));
  OAI210     m267(.A0(mai_mai_n201_), .A1(mai_mai_n183_), .B0(mai_mai_n289_), .Y(mai_mai_n290_));
  AOI220     m268(.A0(mai_mai_n251_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n291_));
  NOi21      m269(.An(mai_mai_n281_), .B(mai_mai_n291_), .Y(mai_mai_n292_));
  AOI210     m270(.A0(mai_mai_n223_), .A1(mai_mai_n77_), .B0(mai_mai_n292_), .Y(mai_mai_n293_));
  AOI210     m271(.A0(mai_mai_n293_), .A1(mai_mai_n290_), .B0(mai_mai_n137_), .Y(mai_mai_n294_));
  NAi21      m272(.An(mai_mai_n225_), .B(mai_mai_n220_), .Y(mai_mai_n295_));
  NO2        m273(.A(mai_mai_n238_), .B(mai_mai_n47_), .Y(mai_mai_n296_));
  NA2        m274(.A(mai_mai_n296_), .B(mai_mai_n295_), .Y(mai_mai_n297_));
  AN2        m275(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n298_));
  OAI210     m276(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n299_));
  NA2        m277(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n300_));
  AOI210     m278(.A0(mai_mai_n139_), .A1(mai_mai_n135_), .B0(mai_mai_n299_), .Y(mai_mai_n301_));
  OAI210     m279(.A0(mai_mai_n301_), .A1(mai_mai_n298_), .B0(mai_mai_n94_), .Y(mai_mai_n302_));
  NA3        m280(.A(mai_mai_n94_), .B(mai_mai_n82_), .C(mai_mai_n217_), .Y(mai_mai_n303_));
  NA3        m281(.A(mai_mai_n93_), .B(mai_mai_n81_), .C(mai_mai_n42_), .Y(mai_mai_n304_));
  AOI210     m282(.A0(mai_mai_n304_), .A1(mai_mai_n303_), .B0(x04), .Y(mai_mai_n305_));
  INV        m283(.A(mai_mai_n146_), .Y(mai_mai_n306_));
  OAI220     m284(.A0(mai_mai_n252_), .A1(mai_mai_n104_), .B0(mai_mai_n306_), .B1(mai_mai_n128_), .Y(mai_mai_n307_));
  AOI210     m285(.A0(mai_mai_n307_), .A1(x13), .B0(mai_mai_n305_), .Y(mai_mai_n308_));
  NA3        m286(.A(mai_mai_n308_), .B(mai_mai_n302_), .C(mai_mai_n297_), .Y(mai_mai_n309_));
  NO3        m287(.A(mai_mai_n309_), .B(mai_mai_n294_), .C(mai_mai_n288_), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n136_), .B(x03), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n174_), .Y(mai_mai_n312_));
  OAI210     m290(.A0(mai_mai_n51_), .A1(mai_mai_n35_), .B0(mai_mai_n36_), .Y(mai_mai_n313_));
  AOI220     m291(.A0(mai_mai_n313_), .A1(mai_mai_n312_), .B0(mai_mai_n194_), .B1(x08), .Y(mai_mai_n314_));
  OAI210     m292(.A0(mai_mai_n314_), .A1(mai_mai_n274_), .B0(mai_mai_n311_), .Y(mai_mai_n315_));
  NA2        m293(.A(mai_mai_n315_), .B(mai_mai_n106_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n164_), .B(mai_mai_n158_), .Y(mai_mai_n317_));
  AN2        m295(.A(mai_mai_n317_), .B(mai_mai_n170_), .Y(mai_mai_n318_));
  INV        m296(.A(mai_mai_n56_), .Y(mai_mai_n319_));
  OAI220     m297(.A0(mai_mai_n265_), .A1(mai_mai_n319_), .B0(mai_mai_n129_), .B1(mai_mai_n28_), .Y(mai_mai_n320_));
  OAI210     m298(.A0(mai_mai_n320_), .A1(mai_mai_n318_), .B0(mai_mai_n107_), .Y(mai_mai_n321_));
  NA2        m299(.A(mai_mai_n265_), .B(mai_mai_n99_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n99_), .B(mai_mai_n41_), .Y(mai_mai_n323_));
  NA3        m301(.A(mai_mai_n323_), .B(mai_mai_n322_), .C(mai_mai_n128_), .Y(mai_mai_n324_));
  NA4        m302(.A(mai_mai_n324_), .B(mai_mai_n321_), .C(mai_mai_n316_), .D(mai_mai_n48_), .Y(mai_mai_n325_));
  INV        m303(.A(mai_mai_n194_), .Y(mai_mai_n326_));
  NO2        m304(.A(mai_mai_n159_), .B(mai_mai_n40_), .Y(mai_mai_n327_));
  NA2        m305(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n328_));
  OAI220     m306(.A0(mai_mai_n328_), .A1(mai_mai_n327_), .B0(mai_mai_n326_), .B1(mai_mai_n59_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n329_), .B(x02), .Y(mai_mai_n330_));
  INV        m308(.A(mai_mai_n231_), .Y(mai_mai_n331_));
  NA2        m309(.A(mai_mai_n191_), .B(x04), .Y(mai_mai_n332_));
  NO2        m310(.A(mai_mai_n332_), .B(mai_mai_n331_), .Y(mai_mai_n333_));
  NO3        m311(.A(mai_mai_n176_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n334_));
  OAI210     m312(.A0(mai_mai_n334_), .A1(mai_mai_n333_), .B0(mai_mai_n94_), .Y(mai_mai_n335_));
  NO3        m313(.A(mai_mai_n191_), .B(mai_mai_n157_), .C(mai_mai_n52_), .Y(mai_mai_n336_));
  OAI210     m314(.A0(mai_mai_n141_), .A1(mai_mai_n36_), .B0(mai_mai_n99_), .Y(mai_mai_n337_));
  OAI210     m315(.A0(mai_mai_n337_), .A1(mai_mai_n184_), .B0(mai_mai_n336_), .Y(mai_mai_n338_));
  NA4        m316(.A(mai_mai_n338_), .B(mai_mai_n335_), .C(mai_mai_n330_), .D(x06), .Y(mai_mai_n339_));
  NA2        m317(.A(x09), .B(x03), .Y(mai_mai_n340_));
  OAI220     m318(.A0(mai_mai_n340_), .A1(mai_mai_n127_), .B0(mai_mai_n200_), .B1(mai_mai_n64_), .Y(mai_mai_n341_));
  OAI220     m319(.A0(mai_mai_n158_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n342_));
  NA2        m320(.A(mai_mai_n342_), .B(mai_mai_n216_), .Y(mai_mai_n343_));
  NO3        m321(.A(mai_mai_n113_), .B(mai_mai_n127_), .C(mai_mai_n38_), .Y(mai_mai_n344_));
  INV        m322(.A(mai_mai_n344_), .Y(mai_mai_n345_));
  OAI210     m323(.A0(mai_mai_n343_), .A1(mai_mai_n28_), .B0(mai_mai_n345_), .Y(mai_mai_n346_));
  AO220      m324(.A0(mai_mai_n346_), .A1(x04), .B0(mai_mai_n341_), .B1(x05), .Y(mai_mai_n347_));
  AOI210     m325(.A0(mai_mai_n339_), .A1(mai_mai_n325_), .B0(mai_mai_n347_), .Y(mai_mai_n348_));
  OAI210     m326(.A0(mai_mai_n310_), .A1(x12), .B0(mai_mai_n348_), .Y(mai03));
  OR2        m327(.A(mai_mai_n42_), .B(mai_mai_n217_), .Y(mai_mai_n350_));
  AOI210     m328(.A0(mai_mai_n147_), .A1(mai_mai_n99_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  AO210      m329(.A0(mai_mai_n331_), .A1(mai_mai_n84_), .B0(mai_mai_n332_), .Y(mai_mai_n352_));
  NA2        m330(.A(mai_mai_n191_), .B(mai_mai_n146_), .Y(mai_mai_n353_));
  NA3        m331(.A(mai_mai_n353_), .B(mai_mai_n352_), .C(mai_mai_n195_), .Y(mai_mai_n354_));
  OAI210     m332(.A0(mai_mai_n354_), .A1(mai_mai_n351_), .B0(x05), .Y(mai_mai_n355_));
  NA2        m333(.A(mai_mai_n350_), .B(x05), .Y(mai_mai_n356_));
  AOI210     m334(.A0(mai_mai_n135_), .A1(mai_mai_n206_), .B0(mai_mai_n356_), .Y(mai_mai_n357_));
  AOI210     m335(.A0(mai_mai_n219_), .A1(mai_mai_n78_), .B0(mai_mai_n121_), .Y(mai_mai_n358_));
  OAI220     m336(.A0(mai_mai_n358_), .A1(mai_mai_n59_), .B0(mai_mai_n300_), .B1(mai_mai_n291_), .Y(mai_mai_n359_));
  OAI210     m337(.A0(mai_mai_n359_), .A1(mai_mai_n357_), .B0(mai_mai_n99_), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n139_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n361_));
  NO2        m339(.A(mai_mai_n167_), .B(mai_mai_n131_), .Y(mai_mai_n362_));
  OAI220     m340(.A0(mai_mai_n362_), .A1(mai_mai_n37_), .B0(mai_mai_n142_), .B1(x13), .Y(mai_mai_n363_));
  OAI210     m341(.A0(mai_mai_n363_), .A1(mai_mai_n361_), .B0(x04), .Y(mai_mai_n364_));
  NO3        m342(.A(mai_mai_n323_), .B(mai_mai_n83_), .C(mai_mai_n59_), .Y(mai_mai_n365_));
  AOI210     m343(.A0(mai_mai_n180_), .A1(mai_mai_n99_), .B0(mai_mai_n139_), .Y(mai_mai_n366_));
  OA210      m344(.A0(mai_mai_n159_), .A1(x12), .B0(mai_mai_n131_), .Y(mai_mai_n367_));
  NO3        m345(.A(mai_mai_n367_), .B(mai_mai_n366_), .C(mai_mai_n365_), .Y(mai_mai_n368_));
  NA4        m346(.A(mai_mai_n368_), .B(mai_mai_n364_), .C(mai_mai_n360_), .D(mai_mai_n355_), .Y(mai04));
  NO2        m347(.A(mai_mai_n87_), .B(mai_mai_n39_), .Y(mai_mai_n370_));
  XO2        m348(.A(mai_mai_n370_), .B(mai_mai_n241_), .Y(mai05));
  NO2        m349(.A(mai_mai_n299_), .B(mai_mai_n25_), .Y(mai_mai_n372_));
  NA3        m350(.A(mai_mai_n137_), .B(mai_mai_n129_), .C(mai_mai_n31_), .Y(mai_mai_n373_));
  INV        m351(.A(mai_mai_n88_), .Y(mai_mai_n374_));
  AOI210     m352(.A0(mai_mai_n374_), .A1(mai_mai_n373_), .B0(mai_mai_n24_), .Y(mai_mai_n375_));
  OAI210     m353(.A0(mai_mai_n375_), .A1(mai_mai_n372_), .B0(mai_mai_n99_), .Y(mai_mai_n376_));
  NA2        m354(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n377_));
  NA2        m355(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n378_));
  NA2        m356(.A(mai_mai_n246_), .B(x03), .Y(mai_mai_n379_));
  OAI220     m357(.A0(mai_mai_n379_), .A1(mai_mai_n378_), .B0(mai_mai_n377_), .B1(mai_mai_n79_), .Y(mai_mai_n380_));
  OAI210     m358(.A0(mai_mai_n26_), .A1(mai_mai_n99_), .B0(x07), .Y(mai_mai_n381_));
  AOI210     m359(.A0(mai_mai_n380_), .A1(x06), .B0(mai_mai_n381_), .Y(mai_mai_n382_));
  AOI210     m360(.A0(mai_mai_n433_), .A1(mai_mai_n379_), .B0(mai_mai_n249_), .Y(mai_mai_n383_));
  OR2        m361(.A(mai_mai_n383_), .B(mai_mai_n230_), .Y(mai_mai_n384_));
  NA2        m362(.A(mai_mai_n153_), .B(x05), .Y(mai_mai_n385_));
  NA3        m363(.A(mai_mai_n385_), .B(mai_mai_n234_), .C(mai_mai_n228_), .Y(mai_mai_n386_));
  NO2        m364(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n387_));
  OAI210     m365(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n388_));
  OR3        m366(.A(mai_mai_n388_), .B(mai_mai_n387_), .C(mai_mai_n44_), .Y(mai_mai_n389_));
  NA3        m367(.A(mai_mai_n389_), .B(mai_mai_n386_), .C(mai_mai_n384_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n390_), .B(mai_mai_n99_), .Y(mai_mai_n391_));
  NA2        m369(.A(mai_mai_n33_), .B(mai_mai_n99_), .Y(mai_mai_n392_));
  AOI210     m370(.A0(mai_mai_n392_), .A1(mai_mai_n90_), .B0(x07), .Y(mai_mai_n393_));
  AOI220     m371(.A0(mai_mai_n393_), .A1(mai_mai_n391_), .B0(mai_mai_n382_), .B1(mai_mai_n376_), .Y(mai_mai_n394_));
  AOI210     m372(.A0(mai_mai_n387_), .A1(x07), .B0(mai_mai_n136_), .Y(mai_mai_n395_));
  OR2        m373(.A(mai_mai_n395_), .B(x03), .Y(mai_mai_n396_));
  NO2        m374(.A(x07), .B(x11), .Y(mai_mai_n397_));
  NO3        m375(.A(mai_mai_n397_), .B(mai_mai_n138_), .C(mai_mai_n28_), .Y(mai_mai_n398_));
  AOI210     m376(.A0(mai_mai_n398_), .A1(mai_mai_n396_), .B0(mai_mai_n47_), .Y(mai_mai_n399_));
  NA2        m377(.A(mai_mai_n399_), .B(mai_mai_n100_), .Y(mai_mai_n400_));
  AOI210     m378(.A0(mai_mai_n332_), .A1(mai_mai_n109_), .B0(mai_mai_n255_), .Y(mai_mai_n401_));
  NOi21      m379(.An(mai_mai_n311_), .B(mai_mai_n131_), .Y(mai_mai_n402_));
  NO2        m380(.A(mai_mai_n402_), .B(mai_mai_n256_), .Y(mai_mai_n403_));
  OAI210     m381(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n404_));
  AOI210     m382(.A0(mai_mai_n241_), .A1(mai_mai_n47_), .B0(mai_mai_n404_), .Y(mai_mai_n405_));
  NO4        m383(.A(mai_mai_n405_), .B(mai_mai_n403_), .C(mai_mai_n401_), .D(x08), .Y(mai_mai_n406_));
  NO2        m384(.A(x05), .B(x03), .Y(mai_mai_n407_));
  NO2        m385(.A(x13), .B(x12), .Y(mai_mai_n408_));
  NO2        m386(.A(mai_mai_n129_), .B(mai_mai_n28_), .Y(mai_mai_n409_));
  NO2        m387(.A(mai_mai_n409_), .B(mai_mai_n260_), .Y(mai_mai_n410_));
  NA3        m388(.A(mai_mai_n326_), .B(mai_mai_n123_), .C(x12), .Y(mai_mai_n411_));
  AO210      m389(.A0(mai_mai_n326_), .A1(mai_mai_n123_), .B0(mai_mai_n241_), .Y(mai_mai_n412_));
  NA3        m390(.A(mai_mai_n412_), .B(mai_mai_n411_), .C(x08), .Y(mai_mai_n413_));
  AOI210     m391(.A0(mai_mai_n408_), .A1(mai_mai_n407_), .B0(mai_mai_n413_), .Y(mai_mai_n414_));
  AOI210     m392(.A0(mai_mai_n406_), .A1(mai_mai_n400_), .B0(mai_mai_n414_), .Y(mai_mai_n415_));
  OAI210     m393(.A0(x07), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n416_));
  OAI220     m394(.A0(mai_mai_n434_), .A1(mai_mai_n378_), .B0(mai_mai_n138_), .B1(mai_mai_n43_), .Y(mai_mai_n417_));
  OAI210     m395(.A0(mai_mai_n417_), .A1(mai_mai_n416_), .B0(mai_mai_n179_), .Y(mai_mai_n418_));
  NA3        m396(.A(mai_mai_n410_), .B(mai_mai_n402_), .C(mai_mai_n322_), .Y(mai_mai_n419_));
  INV        m397(.A(x14), .Y(mai_mai_n420_));
  NO3        m398(.A(mai_mai_n311_), .B(mai_mai_n104_), .C(x11), .Y(mai_mai_n421_));
  NO2        m399(.A(mai_mai_n421_), .B(mai_mai_n420_), .Y(mai_mai_n422_));
  NA3        m400(.A(mai_mai_n422_), .B(mai_mai_n419_), .C(mai_mai_n418_), .Y(mai_mai_n423_));
  AOI220     m401(.A0(mai_mai_n392_), .A1(mai_mai_n61_), .B0(mai_mai_n409_), .B1(mai_mai_n157_), .Y(mai_mai_n424_));
  NOi21      m402(.An(mai_mai_n265_), .B(mai_mai_n142_), .Y(mai_mai_n425_));
  NA2        m403(.A(mai_mai_n272_), .B(mai_mai_n222_), .Y(mai_mai_n426_));
  OAI210     m404(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n426_), .Y(mai_mai_n427_));
  OAI210     m405(.A0(mai_mai_n427_), .A1(mai_mai_n425_), .B0(mai_mai_n99_), .Y(mai_mai_n428_));
  OAI210     m406(.A0(mai_mai_n424_), .A1(mai_mai_n89_), .B0(mai_mai_n428_), .Y(mai_mai_n429_));
  NO4        m407(.A(mai_mai_n429_), .B(mai_mai_n423_), .C(mai_mai_n415_), .D(mai_mai_n394_), .Y(mai06));
  INV        m408(.A(x02), .Y(mai_mai_n433_));
  INV        m409(.A(x07), .Y(mai_mai_n434_));
  INV        m410(.A(x01), .Y(mai_mai_n435_));
  INV        m411(.A(x02), .Y(mai_mai_n436_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  AOI220     u039(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n61_), .Y(men_men_n62_));
  INV        u040(.A(men_men_n59_), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n29_), .B(x02), .Y(men_men_n64_));
  NA2        u042(.A(men_men_n64_), .B(men_men_n24_), .Y(men_men_n65_));
  OAI220     u043(.A0(men_men_n65_), .A1(men_men_n63_), .B0(men_men_n62_), .B1(men_men_n60_), .Y(men_men_n66_));
  NA2        u044(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n67_));
  OAI210     u045(.A0(men_men_n30_), .A1(x11), .B0(men_men_n67_), .Y(men_men_n68_));
  AOI220     u046(.A0(men_men_n68_), .A1(men_men_n59_), .B0(men_men_n66_), .B1(men_men_n31_), .Y(men_men_n69_));
  AOI210     u047(.A0(men_men_n69_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n70_));
  NA2        u048(.A(x10), .B(x09), .Y(men_men_n71_));
  NO2        u049(.A(men_men_n61_), .B(men_men_n23_), .Y(men_men_n72_));
  NA2        u050(.A(x09), .B(x05), .Y(men_men_n73_));
  NA2        u051(.A(x10), .B(x06), .Y(men_men_n74_));
  NA3        u052(.A(men_men_n74_), .B(men_men_n73_), .C(men_men_n28_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n76_));
  OAI210     u054(.A0(men_men_n75_), .A1(men_men_n72_), .B0(x03), .Y(men_men_n77_));
  NOi31      u055(.An(x08), .B(x04), .C(x00), .Y(men_men_n78_));
  NO2        u056(.A(x10), .B(x09), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n456_), .B(men_men_n24_), .Y(men_men_n80_));
  NO2        u058(.A(x09), .B(men_men_n41_), .Y(men_men_n81_));
  NO2        u059(.A(men_men_n81_), .B(men_men_n36_), .Y(men_men_n82_));
  OAI210     u060(.A0(men_men_n81_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n83_));
  NO2        u061(.A(men_men_n48_), .B(men_men_n83_), .Y(men_men_n84_));
  NO2        u062(.A(men_men_n36_), .B(x00), .Y(men_men_n85_));
  NO2        u063(.A(x08), .B(x01), .Y(men_men_n86_));
  OAI210     u064(.A0(men_men_n86_), .A1(men_men_n85_), .B0(men_men_n35_), .Y(men_men_n87_));
  NA2        u065(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n88_));
  NO3        u066(.A(men_men_n87_), .B(men_men_n84_), .C(men_men_n80_), .Y(men_men_n89_));
  AN2        u067(.A(men_men_n89_), .B(men_men_n77_), .Y(men_men_n90_));
  INV        u068(.A(men_men_n87_), .Y(men_men_n91_));
  NO2        u069(.A(x06), .B(x05), .Y(men_men_n92_));
  NA2        u070(.A(x11), .B(x00), .Y(men_men_n93_));
  NO2        u071(.A(x11), .B(men_men_n47_), .Y(men_men_n94_));
  NOi21      u072(.An(men_men_n93_), .B(men_men_n94_), .Y(men_men_n95_));
  AOI210     u073(.A0(men_men_n92_), .A1(men_men_n91_), .B0(men_men_n95_), .Y(men_men_n96_));
  NOi21      u074(.An(x01), .B(x10), .Y(men_men_n97_));
  NO2        u075(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n98_));
  NO3        u076(.A(men_men_n98_), .B(men_men_n97_), .C(x06), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n99_), .B(men_men_n27_), .Y(men_men_n100_));
  OAI210     u078(.A0(men_men_n96_), .A1(x07), .B0(men_men_n100_), .Y(men_men_n101_));
  NO3        u079(.A(men_men_n101_), .B(men_men_n90_), .C(men_men_n70_), .Y(men01));
  INV        u080(.A(x12), .Y(men_men_n103_));
  INV        u081(.A(x13), .Y(men_men_n104_));
  NA2        u082(.A(men_men_n457_), .B(men_men_n71_), .Y(men_men_n105_));
  NA2        u083(.A(x08), .B(x04), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n57_), .Y(men_men_n107_));
  NA2        u085(.A(men_men_n107_), .B(men_men_n105_), .Y(men_men_n108_));
  NA2        u086(.A(men_men_n97_), .B(men_men_n28_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(men_men_n73_), .Y(men_men_n110_));
  NO2        u088(.A(x10), .B(x01), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n29_), .B(x00), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n112_), .B(men_men_n111_), .Y(men_men_n113_));
  NA2        u091(.A(x04), .B(men_men_n28_), .Y(men_men_n114_));
  NO3        u092(.A(men_men_n114_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n115_));
  AOI210     u093(.A0(men_men_n115_), .A1(men_men_n113_), .B0(men_men_n110_), .Y(men_men_n116_));
  AOI210     u094(.A0(men_men_n116_), .A1(men_men_n108_), .B0(men_men_n104_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n56_), .B(x05), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n35_), .B(x02), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n104_), .B(men_men_n36_), .Y(men_men_n120_));
  NA3        u098(.A(men_men_n120_), .B(men_men_n119_), .C(x06), .Y(men_men_n121_));
  INV        u099(.A(men_men_n121_), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n86_), .B(x13), .Y(men_men_n123_));
  NA2        u101(.A(x09), .B(men_men_n35_), .Y(men_men_n124_));
  NA2        u102(.A(x13), .B(men_men_n35_), .Y(men_men_n125_));
  NO2        u103(.A(men_men_n125_), .B(x05), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n127_));
  AOI210     u105(.A0(men_men_n127_), .A1(men_men_n123_), .B0(men_men_n74_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n129_));
  NA2        u107(.A(x10), .B(men_men_n57_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n130_), .B(men_men_n129_), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n51_), .B(x05), .Y(men_men_n132_));
  NA2        u110(.A(men_men_n132_), .B(x13), .Y(men_men_n133_));
  NO2        u111(.A(men_men_n60_), .B(x05), .Y(men_men_n134_));
  NOi41      u112(.An(men_men_n133_), .B(men_men_n134_), .C(men_men_n57_), .D(men_men_n131_), .Y(men_men_n135_));
  NO3        u113(.A(men_men_n135_), .B(x06), .C(x03), .Y(men_men_n136_));
  NO4        u114(.A(men_men_n136_), .B(men_men_n128_), .C(men_men_n122_), .D(men_men_n117_), .Y(men_men_n137_));
  NA2        u115(.A(x13), .B(men_men_n36_), .Y(men_men_n138_));
  OAI210     u116(.A0(men_men_n86_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NO2        u118(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n141_));
  OA210      u119(.A0(x00), .A1(men_men_n79_), .B0(men_men_n141_), .Y(men_men_n142_));
  NO2        u120(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n29_), .B(x06), .Y(men_men_n144_));
  AOI210     u122(.A0(men_men_n144_), .A1(men_men_n49_), .B0(men_men_n143_), .Y(men_men_n145_));
  OA210      u123(.A0(men_men_n145_), .A1(men_men_n142_), .B0(men_men_n140_), .Y(men_men_n146_));
  NO2        u124(.A(x09), .B(x05), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n147_), .B(men_men_n47_), .Y(men_men_n148_));
  AOI210     u126(.A0(men_men_n148_), .A1(men_men_n113_), .B0(men_men_n49_), .Y(men_men_n149_));
  NA2        u127(.A(x09), .B(x00), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n118_), .B(men_men_n150_), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n78_), .B(men_men_n51_), .Y(men_men_n152_));
  AOI210     u130(.A0(men_men_n152_), .A1(men_men_n151_), .B0(men_men_n144_), .Y(men_men_n153_));
  NO3        u131(.A(men_men_n153_), .B(men_men_n149_), .C(men_men_n146_), .Y(men_men_n154_));
  NO2        u132(.A(x03), .B(x02), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n87_), .B(men_men_n104_), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n156_), .B(men_men_n155_), .Y(men_men_n157_));
  OA210      u135(.A0(men_men_n154_), .A1(x11), .B0(men_men_n157_), .Y(men_men_n158_));
  OAI210     u136(.A0(men_men_n137_), .A1(men_men_n23_), .B0(men_men_n158_), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n113_), .B(men_men_n40_), .Y(men_men_n160_));
  NAi21      u138(.An(x06), .B(x10), .Y(men_men_n161_));
  NOi21      u139(.An(x01), .B(x13), .Y(men_men_n162_));
  NA2        u140(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  OR2        u141(.A(men_men_n163_), .B(x08), .Y(men_men_n164_));
  AOI210     u142(.A0(men_men_n164_), .A1(men_men_n160_), .B0(men_men_n41_), .Y(men_men_n165_));
  NO2        u143(.A(men_men_n29_), .B(x03), .Y(men_men_n166_));
  NA2        u144(.A(men_men_n104_), .B(x01), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n167_), .B(x08), .Y(men_men_n168_));
  OAI210     u146(.A0(x05), .A1(men_men_n168_), .B0(men_men_n51_), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n169_), .A1(men_men_n166_), .B0(men_men_n48_), .Y(men_men_n170_));
  AOI210     u148(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n170_), .A1(men_men_n165_), .B0(men_men_n171_), .Y(men_men_n172_));
  NA2        u150(.A(x04), .B(x02), .Y(men_men_n173_));
  NA2        u151(.A(x10), .B(x05), .Y(men_men_n174_));
  NA2        u152(.A(x09), .B(x06), .Y(men_men_n175_));
  NO2        u153(.A(x09), .B(x01), .Y(men_men_n176_));
  NO3        u154(.A(men_men_n176_), .B(men_men_n111_), .C(men_men_n31_), .Y(men_men_n177_));
  NA2        u155(.A(men_men_n177_), .B(x00), .Y(men_men_n178_));
  NO2        u156(.A(men_men_n118_), .B(x08), .Y(men_men_n179_));
  NA3        u157(.A(men_men_n162_), .B(men_men_n161_), .C(men_men_n51_), .Y(men_men_n180_));
  NA2        u158(.A(men_men_n97_), .B(x05), .Y(men_men_n181_));
  OAI210     u159(.A0(men_men_n181_), .A1(men_men_n120_), .B0(men_men_n180_), .Y(men_men_n182_));
  AOI210     u160(.A0(men_men_n179_), .A1(x06), .B0(men_men_n182_), .Y(men_men_n183_));
  OAI210     u161(.A0(men_men_n183_), .A1(x11), .B0(men_men_n178_), .Y(men_men_n184_));
  NAi21      u162(.An(men_men_n173_), .B(men_men_n184_), .Y(men_men_n185_));
  INV        u163(.A(men_men_n25_), .Y(men_men_n186_));
  NAi21      u164(.An(x13), .B(x00), .Y(men_men_n187_));
  AOI210     u165(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n187_), .Y(men_men_n188_));
  AOI220     u166(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n174_), .A1(men_men_n35_), .B0(men_men_n189_), .Y(men_men_n190_));
  AN2        u168(.A(men_men_n190_), .B(men_men_n188_), .Y(men_men_n191_));
  NO2        u169(.A(men_men_n98_), .B(x06), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n187_), .B(men_men_n36_), .Y(men_men_n193_));
  INV        u171(.A(men_men_n193_), .Y(men_men_n194_));
  OAI220     u172(.A0(men_men_n194_), .A1(men_men_n175_), .B0(men_men_n192_), .B1(men_men_n73_), .Y(men_men_n195_));
  OAI210     u173(.A0(men_men_n195_), .A1(men_men_n191_), .B0(men_men_n186_), .Y(men_men_n196_));
  NOi21      u174(.An(x09), .B(x00), .Y(men_men_n197_));
  NO3        u175(.A(men_men_n85_), .B(men_men_n197_), .C(men_men_n47_), .Y(men_men_n198_));
  NA2        u176(.A(men_men_n198_), .B(men_men_n130_), .Y(men_men_n199_));
  NA2        u177(.A(x10), .B(x08), .Y(men_men_n200_));
  INV        u178(.A(men_men_n200_), .Y(men_men_n201_));
  NA2        u179(.A(x06), .B(x05), .Y(men_men_n202_));
  OAI210     u180(.A0(men_men_n202_), .A1(men_men_n35_), .B0(men_men_n103_), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n201_), .A1(men_men_n58_), .B0(men_men_n203_), .Y(men_men_n204_));
  NA2        u182(.A(men_men_n204_), .B(men_men_n199_), .Y(men_men_n205_));
  NO2        u183(.A(men_men_n104_), .B(x12), .Y(men_men_n206_));
  AOI210     u184(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n206_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n97_), .B(men_men_n51_), .Y(men_men_n208_));
  NO2        u186(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n209_), .B(x02), .Y(men_men_n210_));
  NO2        u188(.A(men_men_n210_), .B(men_men_n208_), .Y(men_men_n211_));
  AOI210     u189(.A0(men_men_n207_), .A1(men_men_n205_), .B0(men_men_n211_), .Y(men_men_n212_));
  NA4        u190(.A(men_men_n212_), .B(men_men_n196_), .C(men_men_n185_), .D(men_men_n172_), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n159_), .A1(men_men_n103_), .B0(men_men_n213_), .Y(men_men_n214_));
  INV        u192(.A(men_men_n75_), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n215_), .B(men_men_n140_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n217_), .B(men_men_n139_), .Y(men_men_n218_));
  NO2        u196(.A(men_men_n129_), .B(x06), .Y(men_men_n219_));
  INV        u197(.A(men_men_n219_), .Y(men_men_n220_));
  AOI210     u198(.A0(men_men_n220_), .A1(men_men_n216_), .B0(x12), .Y(men_men_n221_));
  INV        u199(.A(men_men_n78_), .Y(men_men_n222_));
  NA2        u200(.A(men_men_n163_), .B(men_men_n57_), .Y(men_men_n223_));
  NA2        u201(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n97_), .B(x06), .Y(men_men_n225_));
  AOI210     u203(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n226_));
  NO3        u204(.A(men_men_n226_), .B(men_men_n225_), .C(men_men_n41_), .Y(men_men_n227_));
  NA4        u205(.A(men_men_n161_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n228_));
  NA2        u206(.A(men_men_n228_), .B(men_men_n144_), .Y(men_men_n229_));
  OAI210     u207(.A0(men_men_n229_), .A1(men_men_n227_), .B0(x02), .Y(men_men_n230_));
  AOI210     u208(.A0(men_men_n230_), .A1(men_men_n224_), .B0(men_men_n23_), .Y(men_men_n231_));
  OAI210     u209(.A0(men_men_n221_), .A1(men_men_n57_), .B0(men_men_n231_), .Y(men_men_n232_));
  INV        u210(.A(men_men_n144_), .Y(men_men_n233_));
  NO2        u211(.A(men_men_n51_), .B(x03), .Y(men_men_n234_));
  OAI210     u212(.A0(men_men_n81_), .A1(men_men_n36_), .B0(men_men_n124_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n104_), .B(x03), .Y(men_men_n236_));
  AOI220     u214(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n78_), .B1(men_men_n234_), .Y(men_men_n237_));
  NA2        u215(.A(men_men_n32_), .B(x06), .Y(men_men_n238_));
  INV        u216(.A(men_men_n161_), .Y(men_men_n239_));
  NOi21      u217(.An(x13), .B(x04), .Y(men_men_n240_));
  NO3        u218(.A(men_men_n240_), .B(men_men_n78_), .C(men_men_n197_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n241_), .B(x05), .Y(men_men_n242_));
  AOI220     u220(.A0(men_men_n242_), .A1(men_men_n238_), .B0(men_men_n239_), .B1(men_men_n57_), .Y(men_men_n243_));
  OAI210     u221(.A0(men_men_n237_), .A1(men_men_n233_), .B0(men_men_n243_), .Y(men_men_n244_));
  INV        u222(.A(men_men_n94_), .Y(men_men_n245_));
  NO2        u223(.A(men_men_n245_), .B(x12), .Y(men_men_n246_));
  NA2        u224(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n248_));
  OAI210     u226(.A0(men_men_n248_), .A1(men_men_n190_), .B0(men_men_n188_), .Y(men_men_n249_));
  AOI210     u227(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n250_));
  OAI210     u228(.A0(men_men_n106_), .A1(men_men_n150_), .B0(men_men_n74_), .Y(men_men_n251_));
  INV        u229(.A(men_men_n251_), .Y(men_men_n252_));
  NA2        u230(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n253_));
  INV        u231(.A(x03), .Y(men_men_n254_));
  OA210      u232(.A0(men_men_n254_), .A1(men_men_n252_), .B0(men_men_n249_), .Y(men_men_n255_));
  NA2        u233(.A(x13), .B(men_men_n103_), .Y(men_men_n256_));
  NA3        u234(.A(men_men_n256_), .B(men_men_n203_), .C(men_men_n95_), .Y(men_men_n257_));
  OAI210     u235(.A0(men_men_n255_), .A1(men_men_n247_), .B0(men_men_n257_), .Y(men_men_n258_));
  AOI210     u236(.A0(men_men_n246_), .A1(men_men_n244_), .B0(men_men_n258_), .Y(men_men_n259_));
  AOI210     u237(.A0(men_men_n259_), .A1(men_men_n232_), .B0(x07), .Y(men_men_n260_));
  NA2        u238(.A(men_men_n73_), .B(men_men_n29_), .Y(men_men_n261_));
  AOI210     u239(.A0(men_men_n138_), .A1(men_men_n152_), .B0(men_men_n261_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n104_), .B(x06), .Y(men_men_n263_));
  INV        u241(.A(men_men_n263_), .Y(men_men_n264_));
  NO2        u242(.A(x08), .B(x05), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n265_), .B(men_men_n250_), .Y(men_men_n266_));
  OAI210     u244(.A0(men_men_n78_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n267_));
  OAI210     u245(.A0(men_men_n266_), .A1(men_men_n264_), .B0(men_men_n267_), .Y(men_men_n268_));
  NO2        u246(.A(x12), .B(x02), .Y(men_men_n269_));
  INV        u247(.A(men_men_n269_), .Y(men_men_n270_));
  NO2        u248(.A(men_men_n270_), .B(men_men_n245_), .Y(men_men_n271_));
  OA210      u249(.A0(men_men_n268_), .A1(men_men_n262_), .B0(men_men_n271_), .Y(men_men_n272_));
  NA2        u250(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n273_), .B(x01), .Y(men_men_n274_));
  NO2        u252(.A(men_men_n86_), .B(men_men_n274_), .Y(men_men_n275_));
  AOI210     u253(.A0(men_men_n275_), .A1(men_men_n133_), .B0(men_men_n29_), .Y(men_men_n276_));
  NA2        u254(.A(men_men_n263_), .B(men_men_n235_), .Y(men_men_n277_));
  NA2        u255(.A(men_men_n104_), .B(x04), .Y(men_men_n278_));
  OAI210     u256(.A0(x02), .A1(men_men_n123_), .B0(men_men_n277_), .Y(men_men_n279_));
  NO3        u257(.A(men_men_n93_), .B(x12), .C(x03), .Y(men_men_n280_));
  OAI210     u258(.A0(men_men_n279_), .A1(men_men_n276_), .B0(men_men_n280_), .Y(men_men_n281_));
  AOI210     u259(.A0(men_men_n208_), .A1(men_men_n202_), .B0(men_men_n106_), .Y(men_men_n282_));
  NOi21      u260(.An(men_men_n261_), .B(men_men_n225_), .Y(men_men_n283_));
  NO2        u261(.A(men_men_n25_), .B(x00), .Y(men_men_n284_));
  OAI210     u262(.A0(men_men_n283_), .A1(men_men_n282_), .B0(men_men_n284_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n58_), .B(x05), .Y(men_men_n286_));
  NO3        u264(.A(men_men_n286_), .B(men_men_n226_), .C(men_men_n192_), .Y(men_men_n287_));
  NO2        u265(.A(men_men_n247_), .B(men_men_n28_), .Y(men_men_n288_));
  OAI210     u266(.A0(men_men_n287_), .A1(men_men_n233_), .B0(men_men_n288_), .Y(men_men_n289_));
  NA3        u267(.A(men_men_n289_), .B(men_men_n285_), .C(men_men_n281_), .Y(men_men_n290_));
  NO3        u268(.A(men_men_n290_), .B(men_men_n272_), .C(men_men_n260_), .Y(men_men_n291_));
  OAI210     u269(.A0(men_men_n214_), .A1(men_men_n61_), .B0(men_men_n291_), .Y(men02));
  AOI210     u270(.A0(men_men_n138_), .A1(men_men_n87_), .B0(men_men_n132_), .Y(men_men_n293_));
  NOi21      u271(.An(men_men_n241_), .B(men_men_n176_), .Y(men_men_n294_));
  NO2        u272(.A(men_men_n104_), .B(men_men_n35_), .Y(men_men_n295_));
  NA3        u273(.A(men_men_n295_), .B(men_men_n201_), .C(men_men_n56_), .Y(men_men_n296_));
  OAI210     u274(.A0(men_men_n294_), .A1(men_men_n32_), .B0(men_men_n296_), .Y(men_men_n297_));
  OAI210     u275(.A0(men_men_n297_), .A1(men_men_n293_), .B0(men_men_n174_), .Y(men_men_n298_));
  INV        u276(.A(men_men_n174_), .Y(men_men_n299_));
  AOI210     u277(.A0(men_men_n119_), .A1(men_men_n88_), .B0(men_men_n226_), .Y(men_men_n300_));
  NO2        u278(.A(men_men_n300_), .B(men_men_n104_), .Y(men_men_n301_));
  AOI220     u279(.A0(men_men_n301_), .A1(men_men_n299_), .B0(men_men_n156_), .B1(men_men_n155_), .Y(men_men_n302_));
  AOI210     u280(.A0(men_men_n302_), .A1(men_men_n298_), .B0(men_men_n48_), .Y(men_men_n303_));
  NO2        u281(.A(x05), .B(x02), .Y(men_men_n304_));
  OAI210     u282(.A0(men_men_n218_), .A1(men_men_n197_), .B0(men_men_n304_), .Y(men_men_n305_));
  AOI220     u283(.A0(men_men_n265_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n306_));
  NOi21      u284(.An(men_men_n295_), .B(men_men_n306_), .Y(men_men_n307_));
  AOI210     u285(.A0(men_men_n240_), .A1(men_men_n81_), .B0(men_men_n307_), .Y(men_men_n308_));
  AOI210     u286(.A0(men_men_n308_), .A1(men_men_n305_), .B0(men_men_n144_), .Y(men_men_n309_));
  NAi21      u287(.An(men_men_n242_), .B(men_men_n237_), .Y(men_men_n310_));
  NO2        u288(.A(men_men_n253_), .B(men_men_n47_), .Y(men_men_n311_));
  NA2        u289(.A(men_men_n311_), .B(men_men_n310_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n313_));
  NA2        u291(.A(x13), .B(men_men_n28_), .Y(men_men_n314_));
  OA210      u292(.A0(men_men_n314_), .A1(x08), .B0(men_men_n148_), .Y(men_men_n315_));
  AOI210     u293(.A0(men_men_n315_), .A1(men_men_n139_), .B0(men_men_n313_), .Y(men_men_n316_));
  NA2        u294(.A(men_men_n316_), .B(men_men_n98_), .Y(men_men_n317_));
  NA3        u295(.A(men_men_n98_), .B(men_men_n86_), .C(men_men_n234_), .Y(men_men_n318_));
  NA3        u296(.A(men_men_n97_), .B(men_men_n85_), .C(men_men_n42_), .Y(men_men_n319_));
  AOI210     u297(.A0(men_men_n319_), .A1(men_men_n318_), .B0(x04), .Y(men_men_n320_));
  INV        u298(.A(men_men_n155_), .Y(men_men_n321_));
  OAI220     u299(.A0(men_men_n266_), .A1(men_men_n109_), .B0(men_men_n321_), .B1(men_men_n131_), .Y(men_men_n322_));
  AOI210     u300(.A0(men_men_n322_), .A1(x13), .B0(men_men_n320_), .Y(men_men_n323_));
  NA3        u301(.A(men_men_n323_), .B(men_men_n317_), .C(men_men_n312_), .Y(men_men_n324_));
  NO3        u302(.A(men_men_n324_), .B(men_men_n309_), .C(men_men_n303_), .Y(men_men_n325_));
  NA2        u303(.A(men_men_n143_), .B(x03), .Y(men_men_n326_));
  OAI210     u304(.A0(men_men_n187_), .A1(men_men_n286_), .B0(men_men_n326_), .Y(men_men_n327_));
  NA2        u305(.A(men_men_n327_), .B(men_men_n111_), .Y(men_men_n328_));
  INV        u306(.A(men_men_n56_), .Y(men_men_n329_));
  OAI220     u307(.A0(men_men_n278_), .A1(men_men_n329_), .B0(men_men_n132_), .B1(men_men_n28_), .Y(men_men_n330_));
  NA2        u308(.A(men_men_n330_), .B(men_men_n112_), .Y(men_men_n331_));
  NA2        u309(.A(men_men_n278_), .B(men_men_n103_), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n103_), .B(men_men_n41_), .Y(men_men_n333_));
  NA3        u311(.A(men_men_n333_), .B(men_men_n332_), .C(men_men_n131_), .Y(men_men_n334_));
  NA4        u312(.A(men_men_n334_), .B(men_men_n331_), .C(men_men_n328_), .D(men_men_n48_), .Y(men_men_n335_));
  INV        u313(.A(men_men_n209_), .Y(men_men_n336_));
  NO2        u314(.A(men_men_n168_), .B(men_men_n40_), .Y(men_men_n337_));
  NA2        u315(.A(men_men_n32_), .B(x05), .Y(men_men_n338_));
  OAI220     u316(.A0(men_men_n338_), .A1(men_men_n337_), .B0(men_men_n336_), .B1(men_men_n59_), .Y(men_men_n339_));
  NA2        u317(.A(men_men_n339_), .B(x02), .Y(men_men_n340_));
  INV        u318(.A(men_men_n248_), .Y(men_men_n341_));
  NA2        u319(.A(men_men_n206_), .B(x04), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n342_), .B(men_men_n341_), .Y(men_men_n343_));
  NO3        u321(.A(men_men_n189_), .B(x13), .C(men_men_n31_), .Y(men_men_n344_));
  OAI210     u322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n98_), .Y(men_men_n345_));
  NO3        u323(.A(men_men_n206_), .B(men_men_n166_), .C(men_men_n52_), .Y(men_men_n346_));
  OAI210     u324(.A0(x12), .A1(men_men_n198_), .B0(men_men_n346_), .Y(men_men_n347_));
  NA4        u325(.A(men_men_n347_), .B(men_men_n345_), .C(men_men_n340_), .D(x06), .Y(men_men_n348_));
  NA2        u326(.A(x09), .B(x03), .Y(men_men_n349_));
  OAI220     u327(.A0(men_men_n349_), .A1(men_men_n130_), .B0(men_men_n217_), .B1(men_men_n64_), .Y(men_men_n350_));
  OAI220     u328(.A0(men_men_n167_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n351_));
  NO3        u329(.A(men_men_n286_), .B(men_men_n129_), .C(x08), .Y(men_men_n352_));
  AOI210     u330(.A0(men_men_n351_), .A1(men_men_n233_), .B0(men_men_n352_), .Y(men_men_n353_));
  NO2        u331(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n354_));
  NA2        u332(.A(men_men_n346_), .B(men_men_n354_), .Y(men_men_n355_));
  OAI210     u333(.A0(men_men_n353_), .A1(men_men_n28_), .B0(men_men_n355_), .Y(men_men_n356_));
  AO220      u334(.A0(men_men_n356_), .A1(x04), .B0(men_men_n350_), .B1(x05), .Y(men_men_n357_));
  AOI210     u335(.A0(men_men_n348_), .A1(men_men_n335_), .B0(men_men_n357_), .Y(men_men_n358_));
  OAI210     u336(.A0(men_men_n325_), .A1(x12), .B0(men_men_n358_), .Y(men03));
  OR2        u337(.A(men_men_n42_), .B(men_men_n234_), .Y(men_men_n360_));
  AOI210     u338(.A0(men_men_n156_), .A1(men_men_n103_), .B0(men_men_n360_), .Y(men_men_n361_));
  AO210      u339(.A0(men_men_n341_), .A1(men_men_n88_), .B0(men_men_n342_), .Y(men_men_n362_));
  NA2        u340(.A(men_men_n206_), .B(men_men_n155_), .Y(men_men_n363_));
  NA3        u341(.A(men_men_n363_), .B(men_men_n362_), .C(men_men_n210_), .Y(men_men_n364_));
  OAI210     u342(.A0(men_men_n364_), .A1(men_men_n361_), .B0(x05), .Y(men_men_n365_));
  NA2        u343(.A(men_men_n360_), .B(x05), .Y(men_men_n366_));
  AOI210     u344(.A0(men_men_n139_), .A1(men_men_n222_), .B0(men_men_n366_), .Y(men_men_n367_));
  AOI210     u345(.A0(men_men_n236_), .A1(men_men_n82_), .B0(men_men_n126_), .Y(men_men_n368_));
  OAI220     u346(.A0(men_men_n368_), .A1(men_men_n59_), .B0(men_men_n314_), .B1(men_men_n306_), .Y(men_men_n369_));
  OAI210     u347(.A0(men_men_n369_), .A1(men_men_n367_), .B0(men_men_n103_), .Y(men_men_n370_));
  AOI210     u348(.A0(men_men_n148_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n371_));
  NO2        u349(.A(men_men_n176_), .B(men_men_n134_), .Y(men_men_n372_));
  OAI220     u350(.A0(men_men_n372_), .A1(men_men_n37_), .B0(men_men_n151_), .B1(x13), .Y(men_men_n373_));
  OAI210     u351(.A0(men_men_n373_), .A1(men_men_n371_), .B0(x04), .Y(men_men_n374_));
  NO3        u352(.A(men_men_n333_), .B(men_men_n87_), .C(men_men_n59_), .Y(men_men_n375_));
  AOI210     u353(.A0(men_men_n194_), .A1(men_men_n103_), .B0(men_men_n148_), .Y(men_men_n376_));
  OA210      u354(.A0(men_men_n168_), .A1(x12), .B0(men_men_n134_), .Y(men_men_n377_));
  NO3        u355(.A(men_men_n377_), .B(men_men_n376_), .C(men_men_n375_), .Y(men_men_n378_));
  NA4        u356(.A(men_men_n378_), .B(men_men_n374_), .C(men_men_n370_), .D(men_men_n365_), .Y(men04));
  NO2        u357(.A(men_men_n91_), .B(men_men_n39_), .Y(men_men_n380_));
  XO2        u358(.A(men_men_n380_), .B(men_men_n256_), .Y(men05));
  AOI210     u359(.A0(men_men_n73_), .A1(men_men_n52_), .B0(men_men_n219_), .Y(men_men_n382_));
  AOI210     u360(.A0(men_men_n382_), .A1(men_men_n313_), .B0(men_men_n25_), .Y(men_men_n383_));
  NAi31      u361(.An(men_men_n79_), .B(men_men_n132_), .C(men_men_n31_), .Y(men_men_n384_));
  AOI210     u362(.A0(men_men_n239_), .A1(men_men_n57_), .B0(men_men_n92_), .Y(men_men_n385_));
  AOI210     u363(.A0(men_men_n385_), .A1(men_men_n384_), .B0(men_men_n24_), .Y(men_men_n386_));
  OAI210     u364(.A0(men_men_n386_), .A1(men_men_n383_), .B0(men_men_n103_), .Y(men_men_n387_));
  NA2        u365(.A(x11), .B(men_men_n31_), .Y(men_men_n388_));
  NA2        u366(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n389_));
  NA2        u367(.A(men_men_n261_), .B(x03), .Y(men_men_n390_));
  OAI220     u368(.A0(men_men_n390_), .A1(men_men_n389_), .B0(men_men_n388_), .B1(men_men_n83_), .Y(men_men_n391_));
  OAI210     u369(.A0(men_men_n26_), .A1(men_men_n103_), .B0(x07), .Y(men_men_n392_));
  AOI210     u370(.A0(men_men_n391_), .A1(x06), .B0(men_men_n392_), .Y(men_men_n393_));
  AOI220     u371(.A0(men_men_n83_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n394_));
  NO3        u372(.A(men_men_n394_), .B(men_men_n23_), .C(x00), .Y(men_men_n395_));
  NA2        u373(.A(men_men_n71_), .B(x02), .Y(men_men_n396_));
  NA2        u374(.A(men_men_n396_), .B(men_men_n390_), .Y(men_men_n397_));
  OR2        u375(.A(men_men_n397_), .B(men_men_n247_), .Y(men_men_n398_));
  NO2        u376(.A(men_men_n23_), .B(x10), .Y(men_men_n399_));
  OAI210     u377(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n400_));
  OR3        u378(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n44_), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n401_), .B(men_men_n398_), .Y(men_men_n402_));
  OAI210     u380(.A0(men_men_n402_), .A1(men_men_n395_), .B0(men_men_n103_), .Y(men_men_n403_));
  NA2        u381(.A(men_men_n33_), .B(men_men_n103_), .Y(men_men_n404_));
  AOI210     u382(.A0(men_men_n404_), .A1(men_men_n94_), .B0(x07), .Y(men_men_n405_));
  AOI220     u383(.A0(men_men_n405_), .A1(men_men_n403_), .B0(men_men_n393_), .B1(men_men_n387_), .Y(men_men_n406_));
  NA3        u384(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n407_));
  AO210      u385(.A0(men_men_n407_), .A1(men_men_n273_), .B0(men_men_n270_), .Y(men_men_n408_));
  AOI210     u386(.A0(men_men_n399_), .A1(men_men_n76_), .B0(men_men_n143_), .Y(men_men_n409_));
  OR2        u387(.A(men_men_n409_), .B(x03), .Y(men_men_n410_));
  NA2        u388(.A(men_men_n354_), .B(men_men_n61_), .Y(men_men_n411_));
  NO2        u389(.A(men_men_n411_), .B(x11), .Y(men_men_n412_));
  NO2        u390(.A(men_men_n412_), .B(men_men_n28_), .Y(men_men_n413_));
  AOI220     u391(.A0(men_men_n413_), .A1(men_men_n410_), .B0(men_men_n408_), .B1(men_men_n47_), .Y(men_men_n414_));
  NO4        u392(.A(men_men_n333_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n415_));
  OAI210     u393(.A0(men_men_n415_), .A1(men_men_n414_), .B0(men_men_n104_), .Y(men_men_n416_));
  AOI210     u394(.A0(men_men_n342_), .A1(men_men_n114_), .B0(men_men_n269_), .Y(men_men_n417_));
  NOi21      u395(.An(men_men_n326_), .B(men_men_n134_), .Y(men_men_n418_));
  NO2        u396(.A(men_men_n418_), .B(men_men_n270_), .Y(men_men_n419_));
  OAI210     u397(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n420_));
  AOI210     u398(.A0(men_men_n256_), .A1(men_men_n47_), .B0(men_men_n420_), .Y(men_men_n421_));
  NO4        u399(.A(men_men_n421_), .B(men_men_n419_), .C(men_men_n417_), .D(x08), .Y(men_men_n422_));
  AOI210     u400(.A0(men_men_n399_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n423_));
  NA2        u401(.A(x09), .B(men_men_n41_), .Y(men_men_n424_));
  OAI220     u402(.A0(men_men_n424_), .A1(men_men_n423_), .B0(men_men_n388_), .B1(men_men_n67_), .Y(men_men_n425_));
  NO2        u403(.A(x13), .B(x12), .Y(men_men_n426_));
  NO2        u404(.A(men_men_n132_), .B(men_men_n28_), .Y(men_men_n427_));
  NO2        u405(.A(men_men_n427_), .B(men_men_n274_), .Y(men_men_n428_));
  OR3        u406(.A(men_men_n428_), .B(x12), .C(x03), .Y(men_men_n429_));
  NA3        u407(.A(men_men_n336_), .B(men_men_n127_), .C(x12), .Y(men_men_n430_));
  AO210      u408(.A0(men_men_n336_), .A1(men_men_n127_), .B0(men_men_n256_), .Y(men_men_n431_));
  NA4        u409(.A(men_men_n431_), .B(men_men_n430_), .C(men_men_n429_), .D(x08), .Y(men_men_n432_));
  AOI210     u410(.A0(men_men_n426_), .A1(men_men_n425_), .B0(men_men_n432_), .Y(men_men_n433_));
  AOI210     u411(.A0(men_men_n422_), .A1(men_men_n416_), .B0(men_men_n433_), .Y(men_men_n434_));
  OAI210     u412(.A0(men_men_n411_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n435_));
  NA2        u413(.A(men_men_n299_), .B(x07), .Y(men_men_n436_));
  NO2        u414(.A(men_men_n436_), .B(men_men_n389_), .Y(men_men_n437_));
  OAI210     u415(.A0(men_men_n437_), .A1(men_men_n435_), .B0(men_men_n193_), .Y(men_men_n438_));
  NA3        u416(.A(men_men_n428_), .B(men_men_n418_), .C(men_men_n332_), .Y(men_men_n439_));
  INV        u417(.A(x14), .Y(men_men_n440_));
  NO3        u418(.A(men_men_n326_), .B(men_men_n109_), .C(x11), .Y(men_men_n441_));
  NO3        u419(.A(men_men_n167_), .B(men_men_n76_), .C(men_men_n57_), .Y(men_men_n442_));
  NO3        u420(.A(men_men_n407_), .B(men_men_n333_), .C(men_men_n187_), .Y(men_men_n443_));
  NO4        u421(.A(men_men_n443_), .B(men_men_n442_), .C(men_men_n441_), .D(men_men_n440_), .Y(men_men_n444_));
  NA3        u422(.A(men_men_n444_), .B(men_men_n439_), .C(men_men_n438_), .Y(men_men_n445_));
  AOI220     u423(.A0(men_men_n404_), .A1(men_men_n61_), .B0(men_men_n427_), .B1(men_men_n166_), .Y(men_men_n446_));
  NOi21      u424(.An(men_men_n278_), .B(men_men_n151_), .Y(men_men_n447_));
  NO3        u425(.A(men_men_n129_), .B(men_men_n24_), .C(x06), .Y(men_men_n448_));
  AOI210     u426(.A0(men_men_n284_), .A1(men_men_n239_), .B0(men_men_n448_), .Y(men_men_n449_));
  OAI210     u427(.A0(men_men_n44_), .A1(x04), .B0(men_men_n449_), .Y(men_men_n450_));
  OAI210     u428(.A0(men_men_n450_), .A1(men_men_n447_), .B0(men_men_n103_), .Y(men_men_n451_));
  OAI210     u429(.A0(men_men_n446_), .A1(men_men_n93_), .B0(men_men_n451_), .Y(men_men_n452_));
  NO4        u430(.A(men_men_n452_), .B(men_men_n445_), .C(men_men_n434_), .D(men_men_n406_), .Y(men06));
  INV        u431(.A(x07), .Y(men_men_n456_));
  INV        u432(.A(x01), .Y(men_men_n457_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule