module cla_32bits #(
    parameter int WIDTH = 32   
)(
    input  logic [WIDTH-1:0] A, B,
    input  logic Cin,
    output logic [WIDTH-1:0] S,
    output logic Cout
);
    logic [WIDTH-1:0] G, P, C;
    logic G0300, G0200, G0100, G0704, G0604, G0504, G1108, G1008, G0908, G1512, G1412, G1312, G1500, G1100, G0700, G1400, G1300, G1200, G1000, G0900, G0800, G0600, G0500, G0400;  
    logic P0300, P0200, P0100, P0704, P0604, P0504, P1108, P1008, P0908, P1512, P1412, P1312, P1500, P1100, P0700, P1400, P1300, P1200, P1000, P0900, P0800, P0600, P0500, P0400;


    genvar i;

    generate    
        for (i = 0; i < WIDTH; i = i + 1) begin : GENERATE_PROPAGATE
            generate_i  GENERATE  (.Ai(A[i]),.Bi(B[i]),.Gi(G[i]));
            propagate_i PROPAGATE (.Ai(A[i]),.Bi(B[i]),.Pi(P[i]));
        end
    endgenerate

    cla4x3 CLA1 (.G3(G[3]), .G2(G[2]), .G1(G[1]), .G0(G[0]), 
                 .P3(P[3]), .P2(P[2]), .P1(P[1]), .P0(P[0]), 
                 .G30(G0300), .G20(G0200), .G10(G0100), 
                 .P30(P0300), .P20(P0200), .P10(P0100)
    );

    cla4x3 CLA2 (.G3(G[7]), .G2(G[6]), .G1(G[5]), .G0(G[4]), 
                 .P3(P[7]), .P2(P[6]), .P1(P[5]), .P0(P[4]), 
                 .G30(G0704), .G20(G0604), .G10(G0504), 
                 .P30(P0704), .P20(P0604), .P10(P0504)
    );

    cla4x3 CLA3 (.G3(G[11]), .G2(G[10]), .G1(G[9]), .G0(G[8]), 
                 .P3(P[11]), .P2(P[10]), .P1(P[9]), .P0(P[8]), 
                 .G30(G1108), .G20(G1008), .G10(G0908), 
                 .P30(P1108), .P20(P1008), .P10(P0908)
    );

    cla4x3 CLA4 (.G3(G[15]), .G2(G[14]), .G1(G[13]), .G0(G[12]), 
                 .P3(P[15]), .P2(P[14]), .P1(P[13]), .P0(P[12]), 
                 .G30(G1512), .G20(G1412), .G10(G1312), 
                 .P30(P1512), .P20(P1412), .P10(P1312)
    );

    cla4x3 CLA5 (.G3(G[19]), .G2(G[18]), .G1(G[17]), .G0(G[16]), 
                 .P3(P[19]), .P2(P[18]), .P1(P[17]), .P0(P[16]), 
                 .G30(G1916), .G20(G1816), .G10(G1716), 
                 .P30(P1916), .P20(P1816), .P10(P1716)
    );

    cla4x3 CLA6 (.G3(G[23]), .G2(G[22]), .G1(G[21]), .G0(G[20]), 
                 .P3(P[23]), .P2(P[22]), .P1(P[21]), .P0(P[20]), 
                 .G30(G2320), .G20(G2220), .G10(G2120), 
                 .P30(P2320), .P20(P2220), .P10(P2120)
    );

    cla4x3 CLA7 (.G3(G[27]), .G2(G[26]), .G1(G[25]), .G0(G[24]), 
                 .P3(P[27]), .P2(P[26]), .P1(P[25]), .P0(P[24]), 
                 .G30(G2724), .G20(G2624), .G10(G2524), 
                 .P30(P2724), .P20(P2624), .P10(P2524)
    );

    cla4x3 CLA8 (.G3(G[31]), .G2(G[30]), .G1(G[29]), .G0(G[28]), 
                 .P3(P[31]), .P2(P[30]), .P1(P[29]), .P0(P[28]), 
                 .G30(G3128), .G20(G3028), .G10(G2928), 
                 .P30(P3128), .P20(P3028), .P10(P2928)
    );

    cla4x3 CLA9 (.G3(G1512), .G2(G1108), .G1(G0704), .G0(G0300), 
                 .P3(P1512), .P2(P1108), .P1(P0704), .P0(P0300), 
                 .G30(G1500), .G20(G1100), .G10(G0700), 
                 .P30(P1500), .P20(P1100), .P10(P0700)
    );

    cla4x3 CLA10 (.G3(G1412), .G2(G1312), .G1(G[12]), .G0(G1100), 
                 .P3(P1412), .P2(P1312), .P1(P[12]), .P0(P1100), 
                 .G30(G1400), .G20(G1300), .G10(G1200), 
                 .P30(P1400), .P20(P1300), .P10(P1200)
    );

    cla4x3 CLA11 (.G3(G1008), .G2(G0908), .G1(G[8]), .G0(G0700), 
                  .P3(P1008), .P2(P0908), .P1(P[8]), .P0(P0700), 
                  .G30(G1000), .G20(G0900), .G10(G0800), 
                  .P30(P1000), .P20(P0900), .P10(P0800)
    );

    cla4x3 CLA12 (.G3(G0604), .G2(G0504), .G1(G[4]), .G0(G0300), 
                  .P3(P0604), .P2(P0504), .P1(P[4]), .P0(P0300), 
                  .G30(G0600), .G20(G0500), .G10(G0400), 
                  .P30(P0600), .P20(P0500), .P10(P0400)
    );  

    cla4x3 CLA13 (.G3(G2724), .G2(G2320), .G1(G1916), .G0(G1500), 
                  .P3(P2724), .P2(P2320), .P1(P1916), .P0(P1500), 
                  .G30(G2700), .G20(G2300), .G10(G1900), 
                  .P30(P2700), .P20(P2300), .P10(P1900)
    );

    cla4x3 CLA14 (.G3(G2624), .G2(G2524), .G1(G[24]), .G0(G2300), 
                  .P3(P2624), .P2(P2524), .P1(P[24]), .P0(P2300), 
                  .G30(G2600), .G20(G2500), .G10(G2400), 
                  .P30(P2600), .P20(P2500), .P10(P2400)
    );

    cla4x3 CLA15 (.G3(G2220), .G2(G2120), .G1(G[20]), .G0(G1900), 
                  .P3(P2220), .P2(P2120), .P1(P[20]), .P0(P1900), 
                  .G30(G2200), .G20(G2100), .G10(G2000), 
                  .P30(P2200), .P20(P2100), .P10(P2000)
    );

    cla4x3 CLA16 (.G3(G1816), .G2(G1716), .G1(G[16]), .G0(G1500), 
                  .P3(P1816), .P2(P1716), .P1(P[16]), .P0(P1500), 
                  .G30(G1800), .G20(G1700), .G10(G1600), 
                  .P30(P1800), .P20(P1700), .P10(P1600)
    );

    cla4x3 CLA17 (.G3(G3028), .G2(G2928), .G1(G[28]), .G0(G2700), 
                  .P3(P3028), .P2(P2928), .P1(P[28]), .P0(P2700), 
                  .G30(G3000), .G20(G2900), .G10(G2800), 
                  .P30(P3000), .P20(P2900), .P10(P2800)
    );

    bolinha B10 (.Gi(G[31]),.Gj(G3000),.Pi(P[31]),.Pj(P3000),.Gij(G3100),.Pij(P3100));

    
    carry_output #(.N(32)) cs32 (
    .Cin(Cin),
    .G(G),
    .P(P),

    .Go_00({G3100, G3000, G2900, G2800, G2700, G2600, G2500, G2400,
            G2300, G2200, G2100, G2000, G1900, G1800, G1700, G1600,
            G1500, G1400, G1300, G1200, G1100, G1000, G0900, G0800,
            G0700, G0600, G0500, G0400, G0300, G0200, G0100, G0000}),

    .Po_00({P3100, P3000, P2900, P2800, P2700, P2600, P2500, P2400,
            P2300, P2200, P2100, P2000, P1900, P1800, P1700, P1600,
            P1500, P1400, P1300, P1200, P1100, P1000, P0900, P0800,
            P0700, P0600, P0500, P0400, P0300, P0200, P0100, P0000}),

    .C(C),
    .S(S)
);

    assign Cout = C[WIDTH-1];

endmodule