library verilog;
use verilog.vl_types.all;
entity memory_tb is
end memory_tb;
