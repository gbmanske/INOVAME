library verilog;
use verilog.vl_types.all;
entity tb_compare_concat is
end tb_compare_concat;
