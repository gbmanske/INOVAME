// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n132_, new_new_n133_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n974_, new_new_n975_,
    new_new_n976_, new_new_n977_, new_new_n978_, new_new_n979_,
    new_new_n980_, new_new_n981_, new_new_n982_, new_new_n983_,
    new_new_n984_, new_new_n985_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  BUFFER     g015(.A(i_11_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(men1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA3        g031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  OAI210     g034(.A0(new_new_n56_), .A1(new_new_n55_), .B0(new_new_n54_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_12_), .Y(new_new_n58_));
  NAi21      g036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g037(.A(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA3        g039(.A(new_new_n61_), .B(new_new_n59_), .C(new_new_n31_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(new_new_n58_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n50_), .B(i_2_), .Y(new_new_n64_));
  AOI210     g042(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_6_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(new_new_n25_), .Y(new_new_n67_));
  INV        g045(.A(i_0_), .Y(new_new_n68_));
  NAi21      g046(.An(i_5_), .B(i_10_), .Y(new_new_n69_));
  NA2        g047(.A(i_5_), .B(i_9_), .Y(new_new_n70_));
  AOI210     g048(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n68_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n67_), .Y(new_new_n72_));
  OAI210     g050(.A0(new_new_n65_), .A1(new_new_n64_), .B0(new_new_n72_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n73_), .A1(new_new_n63_), .B0(i_0_), .Y(new_new_n74_));
  NA2        g052(.A(i_12_), .B(i_5_), .Y(new_new_n75_));
  NA2        g053(.A(i_2_), .B(i_8_), .Y(new_new_n76_));
  NO2        g054(.A(i_3_), .B(i_9_), .Y(new_new_n77_));
  NO2        g055(.A(i_3_), .B(i_7_), .Y(new_new_n78_));
  INV        g056(.A(i_6_), .Y(new_new_n79_));
  OR4        g057(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n80_));
  INV        g058(.A(new_new_n80_), .Y(new_new_n81_));
  NO2        g059(.A(i_2_), .B(i_7_), .Y(new_new_n82_));
  NAi21      g060(.An(i_6_), .B(i_10_), .Y(new_new_n83_));
  NA2        g061(.A(i_6_), .B(i_9_), .Y(new_new_n84_));
  AOI210     g062(.A0(new_new_n84_), .A1(new_new_n83_), .B0(new_new_n60_), .Y(new_new_n85_));
  NA2        g063(.A(i_2_), .B(i_6_), .Y(new_new_n86_));
  NO3        g064(.A(new_new_n86_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n87_));
  NO2        g065(.A(new_new_n87_), .B(new_new_n85_), .Y(new_new_n88_));
  AOI210     g066(.A0(new_new_n88_), .A1(new_new_n76_), .B0(new_new_n75_), .Y(new_new_n89_));
  AN3        g067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n90_));
  NAi21      g068(.An(i_6_), .B(i_11_), .Y(new_new_n91_));
  NO2        g069(.A(i_5_), .B(i_8_), .Y(new_new_n92_));
  NOi21      g070(.An(new_new_n92_), .B(new_new_n91_), .Y(new_new_n93_));
  AOI220     g071(.A0(new_new_n93_), .A1(new_new_n59_), .B0(new_new_n90_), .B1(new_new_n32_), .Y(new_new_n94_));
  INV        g072(.A(i_7_), .Y(new_new_n95_));
  NA2        g073(.A(new_new_n46_), .B(new_new_n95_), .Y(new_new_n96_));
  NO2        g074(.A(i_0_), .B(i_5_), .Y(new_new_n97_));
  NO2        g075(.A(new_new_n97_), .B(new_new_n79_), .Y(new_new_n98_));
  NA2        g076(.A(i_12_), .B(i_3_), .Y(new_new_n99_));
  INV        g077(.A(new_new_n99_), .Y(new_new_n100_));
  NA3        g078(.A(new_new_n100_), .B(new_new_n98_), .C(new_new_n96_), .Y(new_new_n101_));
  NAi21      g079(.An(i_7_), .B(i_11_), .Y(new_new_n102_));
  NO3        g080(.A(new_new_n102_), .B(new_new_n83_), .C(new_new_n51_), .Y(new_new_n103_));
  AN2        g081(.A(i_2_), .B(i_10_), .Y(new_new_n104_));
  NO2        g082(.A(new_new_n104_), .B(i_7_), .Y(new_new_n105_));
  OR2        g083(.A(new_new_n75_), .B(new_new_n55_), .Y(new_new_n106_));
  NO2        g084(.A(i_8_), .B(new_new_n95_), .Y(new_new_n107_));
  NO3        g085(.A(new_new_n107_), .B(new_new_n106_), .C(new_new_n105_), .Y(new_new_n108_));
  NA2        g086(.A(i_12_), .B(i_7_), .Y(new_new_n109_));
  NA2        g087(.A(i_3_), .B(i_0_), .Y(new_new_n110_));
  NA2        g088(.A(i_11_), .B(i_12_), .Y(new_new_n111_));
  OAI210     g089(.A0(new_new_n110_), .A1(new_new_n109_), .B0(new_new_n111_), .Y(new_new_n112_));
  NO2        g090(.A(new_new_n112_), .B(new_new_n108_), .Y(new_new_n113_));
  NAi41      g091(.An(new_new_n103_), .B(new_new_n113_), .C(new_new_n101_), .D(new_new_n94_), .Y(new_new_n114_));
  NOi21      g092(.An(i_1_), .B(i_5_), .Y(new_new_n115_));
  NA2        g093(.A(new_new_n115_), .B(i_11_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n95_), .B(new_new_n37_), .Y(new_new_n117_));
  NA2        g095(.A(i_7_), .B(new_new_n25_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n118_), .B(new_new_n117_), .Y(new_new_n119_));
  NO2        g097(.A(new_new_n119_), .B(new_new_n46_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n84_), .B(new_new_n83_), .Y(new_new_n121_));
  NAi21      g099(.An(i_3_), .B(i_8_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n122_), .B(new_new_n59_), .Y(new_new_n123_));
  NOi31      g101(.An(new_new_n123_), .B(new_new_n121_), .C(new_new_n120_), .Y(new_new_n124_));
  NO2        g102(.A(i_1_), .B(new_new_n79_), .Y(new_new_n125_));
  NO2        g103(.A(i_6_), .B(i_5_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(i_3_), .Y(new_new_n127_));
  AO210      g105(.A0(new_new_n127_), .A1(new_new_n47_), .B0(new_new_n125_), .Y(new_new_n128_));
  OAI220     g106(.A0(new_new_n128_), .A1(new_new_n102_), .B0(new_new_n124_), .B1(new_new_n116_), .Y(new_new_n129_));
  NO3        g107(.A(new_new_n129_), .B(new_new_n114_), .C(new_new_n89_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n74_), .Y(men2));
  NO2        g109(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n132_));
  NA2        g110(.A(new_new_n982_), .B(new_new_n132_), .Y(new_new_n133_));
  NA4        g111(.A(new_new_n133_), .B(new_new_n72_), .C(new_new_n64_), .D(new_new_n30_), .Y(men0));
  AN2        g112(.A(i_8_), .B(i_7_), .Y(new_new_n135_));
  NA2        g113(.A(new_new_n135_), .B(i_6_), .Y(new_new_n136_));
  NO2        g114(.A(i_12_), .B(i_13_), .Y(new_new_n137_));
  NAi21      g115(.An(i_5_), .B(i_11_), .Y(new_new_n138_));
  NOi21      g116(.An(new_new_n137_), .B(new_new_n138_), .Y(new_new_n139_));
  NO2        g117(.A(i_0_), .B(i_1_), .Y(new_new_n140_));
  NA2        g118(.A(i_2_), .B(i_3_), .Y(new_new_n141_));
  NO2        g119(.A(new_new_n141_), .B(i_4_), .Y(new_new_n142_));
  NA3        g120(.A(new_new_n142_), .B(new_new_n140_), .C(new_new_n139_), .Y(new_new_n143_));
  OR2        g121(.A(new_new_n143_), .B(new_new_n25_), .Y(new_new_n144_));
  AN2        g122(.A(new_new_n137_), .B(new_new_n77_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(new_new_n27_), .Y(new_new_n146_));
  NA2        g124(.A(i_1_), .B(i_5_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n68_), .B(new_new_n46_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n36_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  OR2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NO3        g129(.A(new_new_n151_), .B(new_new_n75_), .C(i_13_), .Y(new_new_n152_));
  NAi32      g130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n153_));
  NAi21      g131(.An(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  NOi21      g132(.An(i_4_), .B(i_10_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n39_), .Y(new_new_n156_));
  NO2        g134(.A(i_3_), .B(i_5_), .Y(new_new_n157_));
  NO3        g135(.A(new_new_n68_), .B(i_2_), .C(i_1_), .Y(new_new_n158_));
  OAI210     g136(.A0(i_2_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n159_));
  NO2        g137(.A(new_new_n159_), .B(new_new_n150_), .Y(new_new_n160_));
  AOI210     g138(.A0(new_new_n160_), .A1(new_new_n144_), .B0(new_new_n136_), .Y(new_new_n161_));
  NA3        g139(.A(new_new_n68_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n162_));
  NOi21      g140(.An(i_4_), .B(i_9_), .Y(new_new_n163_));
  NOi21      g141(.An(i_11_), .B(i_13_), .Y(new_new_n164_));
  NA2        g142(.A(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  NO2        g143(.A(i_4_), .B(i_5_), .Y(new_new_n166_));
  NAi21      g144(.An(i_12_), .B(i_11_), .Y(new_new_n167_));
  NO2        g145(.A(new_new_n167_), .B(i_13_), .Y(new_new_n168_));
  NA2        g146(.A(new_new_n168_), .B(new_new_n166_), .Y(new_new_n169_));
  AOI210     g147(.A0(new_new_n169_), .A1(new_new_n165_), .B0(new_new_n162_), .Y(new_new_n170_));
  NO2        g148(.A(new_new_n68_), .B(new_new_n60_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n36_), .B(i_5_), .Y(new_new_n172_));
  NAi31      g150(.An(new_new_n172_), .B(new_new_n145_), .C(i_11_), .Y(new_new_n173_));
  NA2        g151(.A(i_3_), .B(i_5_), .Y(new_new_n174_));
  OR2        g152(.A(new_new_n174_), .B(new_new_n165_), .Y(new_new_n175_));
  AOI210     g153(.A0(new_new_n175_), .A1(new_new_n173_), .B0(i_2_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n68_), .B(i_5_), .Y(new_new_n177_));
  NO2        g155(.A(i_13_), .B(i_10_), .Y(new_new_n178_));
  NA3        g156(.A(new_new_n178_), .B(new_new_n177_), .C(new_new_n44_), .Y(new_new_n179_));
  NO2        g157(.A(i_2_), .B(i_1_), .Y(new_new_n180_));
  NA2        g158(.A(new_new_n180_), .B(i_3_), .Y(new_new_n181_));
  NAi21      g159(.An(i_4_), .B(i_12_), .Y(new_new_n182_));
  NO3        g160(.A(new_new_n182_), .B(new_new_n181_), .C(new_new_n25_), .Y(new_new_n183_));
  NO3        g161(.A(new_new_n183_), .B(new_new_n176_), .C(new_new_n170_), .Y(new_new_n184_));
  INV        g162(.A(i_8_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n185_), .B(i_7_), .Y(new_new_n186_));
  NA2        g164(.A(new_new_n186_), .B(i_6_), .Y(new_new_n187_));
  NO3        g165(.A(i_3_), .B(new_new_n79_), .C(new_new_n48_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n188_), .B(new_new_n107_), .Y(new_new_n189_));
  NO3        g167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n190_));
  NA3        g168(.A(new_new_n190_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n191_));
  NO3        g169(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n192_));
  OAI210     g170(.A0(new_new_n90_), .A1(i_12_), .B0(new_new_n192_), .Y(new_new_n193_));
  AOI210     g171(.A0(new_new_n193_), .A1(new_new_n191_), .B0(new_new_n189_), .Y(new_new_n194_));
  NO2        g172(.A(i_3_), .B(i_8_), .Y(new_new_n195_));
  NO3        g173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n196_));
  NA3        g174(.A(new_new_n196_), .B(new_new_n195_), .C(new_new_n39_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n97_), .B(new_new_n55_), .Y(new_new_n198_));
  INV        g176(.A(new_new_n198_), .Y(new_new_n199_));
  NO2        g177(.A(i_13_), .B(i_9_), .Y(new_new_n200_));
  NAi21      g178(.An(i_12_), .B(i_3_), .Y(new_new_n201_));
  NO2        g179(.A(new_new_n44_), .B(i_5_), .Y(new_new_n202_));
  NO3        g180(.A(i_0_), .B(i_2_), .C(new_new_n60_), .Y(new_new_n203_));
  NA2        g181(.A(new_new_n203_), .B(i_10_), .Y(new_new_n204_));
  OAI220     g182(.A0(new_new_n204_), .A1(new_new_n201_), .B0(new_new_n199_), .B1(new_new_n197_), .Y(new_new_n205_));
  AOI210     g183(.A0(new_new_n205_), .A1(i_7_), .B0(new_new_n194_), .Y(new_new_n206_));
  OAI220     g184(.A0(new_new_n206_), .A1(i_4_), .B0(new_new_n187_), .B1(new_new_n184_), .Y(new_new_n207_));
  NAi21      g185(.An(i_12_), .B(i_7_), .Y(new_new_n208_));
  NA3        g186(.A(i_13_), .B(new_new_n185_), .C(i_10_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n209_), .B(new_new_n208_), .Y(new_new_n210_));
  NA2        g188(.A(i_0_), .B(i_5_), .Y(new_new_n211_));
  NA2        g189(.A(new_new_n211_), .B(new_new_n98_), .Y(new_new_n212_));
  OAI220     g190(.A0(new_new_n212_), .A1(new_new_n181_), .B0(i_2_), .B1(new_new_n127_), .Y(new_new_n213_));
  NAi31      g191(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n36_), .B(i_13_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n68_), .B(new_new_n26_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n46_), .B(new_new_n60_), .Y(new_new_n217_));
  NA3        g195(.A(new_new_n217_), .B(new_new_n216_), .C(new_new_n215_), .Y(new_new_n218_));
  INV        g196(.A(i_13_), .Y(new_new_n219_));
  NO2        g197(.A(i_12_), .B(new_new_n219_), .Y(new_new_n220_));
  NA3        g198(.A(new_new_n220_), .B(new_new_n190_), .C(new_new_n188_), .Y(new_new_n221_));
  OAI210     g199(.A0(new_new_n218_), .A1(new_new_n214_), .B0(new_new_n221_), .Y(new_new_n222_));
  AOI220     g200(.A0(new_new_n222_), .A1(new_new_n135_), .B0(new_new_n213_), .B1(new_new_n210_), .Y(new_new_n223_));
  NO2        g201(.A(i_12_), .B(new_new_n37_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n174_), .B(i_4_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  OR2        g204(.A(i_8_), .B(i_7_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n79_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n51_), .B(i_1_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n230_));
  INV        g208(.A(i_12_), .Y(new_new_n231_));
  NO3        g209(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n232_));
  NA2        g210(.A(i_2_), .B(i_1_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n230_), .B(new_new_n226_), .Y(new_new_n234_));
  NO3        g212(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n235_));
  NAi21      g213(.An(i_4_), .B(i_3_), .Y(new_new_n236_));
  NO2        g214(.A(i_0_), .B(i_6_), .Y(new_new_n237_));
  NOi41      g215(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n238_), .B(new_new_n237_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n233_), .B(new_new_n174_), .Y(new_new_n240_));
  NAi21      g218(.An(new_new_n239_), .B(new_new_n240_), .Y(new_new_n241_));
  INV        g219(.A(new_new_n241_), .Y(new_new_n242_));
  AOI220     g220(.A0(new_new_n242_), .A1(new_new_n39_), .B0(new_new_n234_), .B1(new_new_n200_), .Y(new_new_n243_));
  NO2        g221(.A(i_11_), .B(new_new_n219_), .Y(new_new_n244_));
  NOi21      g222(.An(i_1_), .B(i_6_), .Y(new_new_n245_));
  NAi21      g223(.An(i_3_), .B(i_7_), .Y(new_new_n246_));
  OR4        g224(.A(i_12_), .B(new_new_n246_), .C(new_new_n245_), .D(new_new_n177_), .Y(new_new_n247_));
  NO2        g225(.A(i_12_), .B(i_3_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n68_), .B(i_5_), .Y(new_new_n249_));
  NA2        g227(.A(i_3_), .B(i_9_), .Y(new_new_n250_));
  NAi21      g228(.An(i_7_), .B(i_10_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n251_), .B(new_new_n250_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n252_), .B(new_new_n249_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n253_), .B(new_new_n247_), .Y(new_new_n254_));
  INV        g232(.A(new_new_n136_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n231_), .B(i_13_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n256_), .B(new_new_n70_), .Y(new_new_n257_));
  AOI220     g235(.A0(new_new_n257_), .A1(new_new_n255_), .B0(new_new_n254_), .B1(new_new_n244_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n227_), .B(new_new_n37_), .Y(new_new_n259_));
  NA2        g237(.A(i_12_), .B(i_6_), .Y(new_new_n260_));
  OR2        g238(.A(i_13_), .B(i_9_), .Y(new_new_n261_));
  NO3        g239(.A(new_new_n261_), .B(new_new_n260_), .C(new_new_n48_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n236_), .B(i_2_), .Y(new_new_n263_));
  NA3        g241(.A(new_new_n263_), .B(new_new_n262_), .C(new_new_n44_), .Y(new_new_n264_));
  NA2        g242(.A(new_new_n244_), .B(i_9_), .Y(new_new_n265_));
  OAI210     g243(.A0(new_new_n68_), .A1(new_new_n265_), .B0(new_new_n264_), .Y(new_new_n266_));
  NO3        g244(.A(i_11_), .B(new_new_n219_), .C(new_new_n25_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n246_), .B(i_8_), .Y(new_new_n268_));
  NO2        g246(.A(i_6_), .B(new_new_n48_), .Y(new_new_n269_));
  NA3        g247(.A(new_new_n269_), .B(new_new_n268_), .C(new_new_n267_), .Y(new_new_n270_));
  NO3        g248(.A(new_new_n26_), .B(new_new_n79_), .C(i_5_), .Y(new_new_n271_));
  NA3        g249(.A(new_new_n271_), .B(new_new_n259_), .C(new_new_n220_), .Y(new_new_n272_));
  AOI210     g250(.A0(new_new_n272_), .A1(new_new_n270_), .B0(new_new_n46_), .Y(new_new_n273_));
  AOI210     g251(.A0(new_new_n266_), .A1(new_new_n259_), .B0(new_new_n273_), .Y(new_new_n274_));
  NA4        g252(.A(new_new_n274_), .B(new_new_n258_), .C(new_new_n243_), .D(new_new_n223_), .Y(new_new_n275_));
  NO3        g253(.A(i_12_), .B(new_new_n219_), .C(new_new_n37_), .Y(new_new_n276_));
  INV        g254(.A(new_new_n276_), .Y(new_new_n277_));
  NOi21      g255(.An(new_new_n157_), .B(new_new_n79_), .Y(new_new_n278_));
  NO3        g256(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n279_));
  AOI220     g257(.A0(new_new_n279_), .A1(new_new_n188_), .B0(new_new_n278_), .B1(new_new_n229_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(i_7_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n233_), .B(i_0_), .Y(new_new_n282_));
  AOI220     g260(.A0(new_new_n282_), .A1(new_new_n186_), .B0(i_1_), .B1(new_new_n135_), .Y(new_new_n283_));
  NA2        g261(.A(new_new_n269_), .B(new_new_n26_), .Y(new_new_n284_));
  NO2        g262(.A(new_new_n284_), .B(new_new_n283_), .Y(new_new_n285_));
  NA2        g263(.A(i_0_), .B(i_1_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n286_), .B(i_2_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n56_), .B(i_6_), .Y(new_new_n288_));
  NO3        g266(.A(new_new_n135_), .B(new_new_n285_), .C(new_new_n281_), .Y(new_new_n289_));
  NO2        g267(.A(i_3_), .B(i_10_), .Y(new_new_n290_));
  NA3        g268(.A(new_new_n290_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n291_));
  NO2        g269(.A(i_2_), .B(new_new_n95_), .Y(new_new_n292_));
  NA2        g270(.A(i_1_), .B(new_new_n36_), .Y(new_new_n293_));
  NOi21      g271(.An(new_new_n211_), .B(new_new_n97_), .Y(new_new_n294_));
  NA3        g272(.A(new_new_n294_), .B(i_1_), .C(new_new_n292_), .Y(new_new_n295_));
  AN2        g273(.A(i_3_), .B(i_10_), .Y(new_new_n296_));
  NA3        g274(.A(new_new_n296_), .B(new_new_n168_), .C(new_new_n166_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n298_));
  OR2        g276(.A(new_new_n295_), .B(new_new_n291_), .Y(new_new_n299_));
  OAI220     g277(.A0(new_new_n299_), .A1(i_6_), .B0(new_new_n289_), .B1(new_new_n277_), .Y(new_new_n300_));
  NO4        g278(.A(new_new_n300_), .B(new_new_n275_), .C(new_new_n207_), .D(new_new_n161_), .Y(new_new_n301_));
  NO3        g279(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n302_));
  NO2        g280(.A(new_new_n56_), .B(new_new_n79_), .Y(new_new_n303_));
  NA2        g281(.A(new_new_n282_), .B(new_new_n303_), .Y(new_new_n304_));
  NO3        g282(.A(i_6_), .B(new_new_n185_), .C(i_7_), .Y(new_new_n305_));
  NA2        g283(.A(new_new_n305_), .B(new_new_n190_), .Y(new_new_n306_));
  AOI210     g284(.A0(new_new_n306_), .A1(new_new_n304_), .B0(i_5_), .Y(new_new_n307_));
  NO2        g285(.A(i_2_), .B(i_3_), .Y(new_new_n308_));
  OR2        g286(.A(i_0_), .B(i_5_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n211_), .B(new_new_n309_), .Y(new_new_n310_));
  NA4        g288(.A(new_new_n310_), .B(new_new_n228_), .C(new_new_n308_), .D(i_1_), .Y(new_new_n311_));
  NA3        g289(.A(new_new_n282_), .B(new_new_n278_), .C(new_new_n107_), .Y(new_new_n312_));
  NAi21      g290(.An(i_8_), .B(i_7_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n313_), .B(i_6_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n151_), .B(new_new_n46_), .Y(new_new_n315_));
  NA3        g293(.A(new_new_n315_), .B(new_new_n314_), .C(new_new_n157_), .Y(new_new_n316_));
  NA3        g294(.A(new_new_n316_), .B(new_new_n312_), .C(new_new_n311_), .Y(new_new_n317_));
  OAI210     g295(.A0(new_new_n317_), .A1(new_new_n307_), .B0(i_4_), .Y(new_new_n318_));
  NO2        g296(.A(i_12_), .B(i_10_), .Y(new_new_n319_));
  NOi21      g297(.An(i_5_), .B(i_0_), .Y(new_new_n320_));
  AOI210     g298(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n95_), .Y(new_new_n321_));
  NO3        g299(.A(new_new_n321_), .B(new_new_n293_), .C(new_new_n122_), .Y(new_new_n322_));
  NA4        g300(.A(new_new_n78_), .B(new_new_n36_), .C(new_new_n79_), .D(i_8_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n322_), .B(new_new_n319_), .Y(new_new_n324_));
  NO2        g302(.A(i_6_), .B(i_8_), .Y(new_new_n325_));
  NOi21      g303(.An(i_0_), .B(i_2_), .Y(new_new_n326_));
  AN2        g304(.A(new_new_n326_), .B(new_new_n325_), .Y(new_new_n327_));
  NO2        g305(.A(i_1_), .B(i_7_), .Y(new_new_n328_));
  NA3        g306(.A(new_new_n325_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n329_));
  NA3        g307(.A(new_new_n329_), .B(new_new_n324_), .C(new_new_n318_), .Y(new_new_n330_));
  NO2        g308(.A(i_8_), .B(new_new_n310_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n97_), .B(new_new_n118_), .Y(new_new_n332_));
  OAI210     g310(.A0(new_new_n332_), .A1(new_new_n331_), .B0(i_3_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n286_), .B(new_new_n76_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(new_new_n126_), .Y(new_new_n335_));
  NA3        g313(.A(new_new_n294_), .B(i_8_), .C(new_new_n60_), .Y(new_new_n336_));
  AOI210     g314(.A0(new_new_n336_), .A1(new_new_n335_), .B0(i_7_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n185_), .B(i_9_), .Y(new_new_n338_));
  NA2        g316(.A(new_new_n338_), .B(new_new_n198_), .Y(new_new_n339_));
  NO2        g317(.A(new_new_n337_), .B(new_new_n285_), .Y(new_new_n340_));
  AOI210     g318(.A0(new_new_n340_), .A1(new_new_n333_), .B0(new_new_n156_), .Y(new_new_n341_));
  AOI210     g319(.A0(new_new_n330_), .A1(new_new_n302_), .B0(new_new_n341_), .Y(new_new_n342_));
  NOi32      g320(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n343_));
  INV        g321(.A(new_new_n343_), .Y(new_new_n344_));
  NAi21      g322(.An(i_0_), .B(i_6_), .Y(new_new_n345_));
  NAi21      g323(.An(i_1_), .B(i_5_), .Y(new_new_n346_));
  NA2        g324(.A(new_new_n346_), .B(new_new_n345_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n347_), .B(new_new_n25_), .Y(new_new_n348_));
  OAI210     g326(.A0(new_new_n348_), .A1(new_new_n153_), .B0(new_new_n239_), .Y(new_new_n349_));
  NAi41      g327(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n350_));
  OAI220     g328(.A0(new_new_n350_), .A1(new_new_n346_), .B0(new_new_n214_), .B1(new_new_n153_), .Y(new_new_n351_));
  AOI210     g329(.A0(new_new_n350_), .A1(new_new_n153_), .B0(new_new_n151_), .Y(new_new_n352_));
  NOi32      g330(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n353_));
  NA2        g331(.A(new_new_n353_), .B(new_new_n46_), .Y(new_new_n354_));
  NO2        g332(.A(new_new_n354_), .B(i_0_), .Y(new_new_n355_));
  OR3        g333(.A(new_new_n355_), .B(new_new_n352_), .C(new_new_n351_), .Y(new_new_n356_));
  NO2        g334(.A(i_1_), .B(new_new_n95_), .Y(new_new_n357_));
  NAi21      g335(.An(i_3_), .B(i_4_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n358_), .B(i_9_), .Y(new_new_n359_));
  AN2        g337(.A(i_6_), .B(i_7_), .Y(new_new_n360_));
  OAI210     g338(.A0(new_new_n360_), .A1(new_new_n357_), .B0(new_new_n359_), .Y(new_new_n361_));
  NA2        g339(.A(i_2_), .B(i_7_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n358_), .B(i_10_), .Y(new_new_n363_));
  AOI220     g341(.A0(new_new_n363_), .A1(new_new_n328_), .B0(new_new_n232_), .B1(new_new_n180_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n356_), .B(new_new_n349_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n365_), .B(new_new_n344_), .Y(new_new_n366_));
  NO2        g344(.A(new_new_n56_), .B(new_new_n25_), .Y(new_new_n367_));
  AN2        g345(.A(i_12_), .B(i_5_), .Y(new_new_n368_));
  NO2        g346(.A(i_4_), .B(new_new_n26_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n369_), .B(new_new_n368_), .Y(new_new_n370_));
  NO2        g348(.A(i_11_), .B(i_6_), .Y(new_new_n371_));
  NA3        g349(.A(new_new_n371_), .B(new_new_n315_), .C(new_new_n219_), .Y(new_new_n372_));
  NO2        g350(.A(new_new_n372_), .B(new_new_n370_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n236_), .B(i_5_), .Y(new_new_n374_));
  NO2        g352(.A(i_5_), .B(i_10_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n137_), .B(new_new_n45_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n376_), .B(new_new_n236_), .Y(new_new_n377_));
  OAI210     g355(.A0(new_new_n377_), .A1(new_new_n373_), .B0(new_new_n367_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n379_));
  INV        g357(.A(new_new_n143_), .Y(new_new_n380_));
  OAI210     g358(.A0(new_new_n380_), .A1(new_new_n373_), .B0(new_new_n379_), .Y(new_new_n381_));
  NO3        g359(.A(new_new_n79_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n382_));
  NO2        g360(.A(i_3_), .B(new_new_n95_), .Y(new_new_n383_));
  NA2        g361(.A(new_new_n290_), .B(new_new_n70_), .Y(new_new_n384_));
  NO2        g362(.A(i_11_), .B(i_12_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n385_), .B(new_new_n36_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n384_), .B(new_new_n386_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n375_), .B(new_new_n231_), .Y(new_new_n388_));
  NA3        g366(.A(new_new_n107_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(new_new_n214_), .Y(new_new_n390_));
  NAi21      g368(.An(i_13_), .B(i_0_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n391_), .B(new_new_n233_), .Y(new_new_n392_));
  OAI210     g370(.A0(new_new_n390_), .A1(new_new_n387_), .B0(new_new_n392_), .Y(new_new_n393_));
  NA3        g371(.A(new_new_n393_), .B(new_new_n381_), .C(new_new_n378_), .Y(new_new_n394_));
  NO3        g372(.A(i_1_), .B(i_12_), .C(new_new_n79_), .Y(new_new_n395_));
  NO2        g373(.A(i_0_), .B(i_11_), .Y(new_new_n396_));
  AN2        g374(.A(i_1_), .B(i_6_), .Y(new_new_n397_));
  NOi21      g375(.An(i_2_), .B(i_12_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n398_), .B(new_new_n397_), .Y(new_new_n399_));
  INV        g377(.A(new_new_n399_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n135_), .B(i_9_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n401_), .B(i_4_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n400_), .B(new_new_n402_), .Y(new_new_n403_));
  OR2        g381(.A(i_13_), .B(i_10_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n165_), .B(new_new_n117_), .Y(new_new_n405_));
  OR2        g383(.A(new_new_n209_), .B(new_new_n208_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n95_), .B(new_new_n25_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n276_), .B(new_new_n407_), .Y(new_new_n408_));
  OAI220     g386(.A0(new_new_n60_), .A1(new_new_n406_), .B0(new_new_n408_), .B1(new_new_n97_), .Y(new_new_n409_));
  INV        g387(.A(new_new_n409_), .Y(new_new_n410_));
  AOI210     g388(.A0(new_new_n410_), .A1(new_new_n403_), .B0(new_new_n26_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n312_), .B(new_new_n311_), .Y(new_new_n412_));
  AOI220     g390(.A0(new_new_n288_), .A1(new_new_n279_), .B0(new_new_n282_), .B1(new_new_n303_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n413_), .B(i_5_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n174_), .B(new_new_n79_), .Y(new_new_n415_));
  AOI220     g393(.A0(new_new_n415_), .A1(new_new_n287_), .B0(new_new_n271_), .B1(new_new_n203_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n416_), .B(i_7_), .Y(new_new_n417_));
  NO3        g395(.A(new_new_n417_), .B(new_new_n414_), .C(new_new_n412_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n188_), .B(new_new_n90_), .Y(new_new_n419_));
  AOI210     g397(.A0(new_new_n151_), .A1(new_new_n419_), .B0(new_new_n313_), .Y(new_new_n420_));
  NA3        g398(.A(new_new_n249_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n288_), .B(new_new_n229_), .Y(new_new_n422_));
  OAI220     g400(.A0(new_new_n422_), .A1(new_new_n174_), .B0(new_new_n421_), .B1(new_new_n978_), .Y(new_new_n423_));
  NO2        g401(.A(i_3_), .B(new_new_n48_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n327_), .B(new_new_n424_), .Y(new_new_n425_));
  NA2        g403(.A(new_new_n305_), .B(new_new_n310_), .Y(new_new_n426_));
  OAI210     g404(.A0(new_new_n426_), .A1(new_new_n181_), .B0(new_new_n425_), .Y(new_new_n427_));
  NO3        g405(.A(new_new_n427_), .B(new_new_n423_), .C(new_new_n420_), .Y(new_new_n428_));
  AOI210     g406(.A0(new_new_n428_), .A1(new_new_n418_), .B0(new_new_n265_), .Y(new_new_n429_));
  NO4        g407(.A(new_new_n429_), .B(new_new_n411_), .C(new_new_n394_), .D(new_new_n366_), .Y(new_new_n430_));
  NO2        g408(.A(new_new_n68_), .B(i_13_), .Y(new_new_n431_));
  NO2        g409(.A(i_10_), .B(i_9_), .Y(new_new_n432_));
  NAi21      g410(.An(i_12_), .B(i_8_), .Y(new_new_n433_));
  NO2        g411(.A(new_new_n433_), .B(i_3_), .Y(new_new_n434_));
  NO2        g412(.A(new_new_n46_), .B(i_4_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n435_), .B(new_new_n98_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n197_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n298_), .B(i_0_), .Y(new_new_n438_));
  NO3        g416(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n260_), .B(new_new_n91_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n440_), .B(new_new_n439_), .Y(new_new_n441_));
  NA2        g419(.A(i_8_), .B(i_9_), .Y(new_new_n442_));
  NO2        g420(.A(new_new_n441_), .B(new_new_n438_), .Y(new_new_n443_));
  NO3        g421(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n444_));
  NA3        g422(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n443_), .B(new_new_n437_), .Y(new_new_n446_));
  NA2        g424(.A(new_new_n287_), .B(new_new_n102_), .Y(new_new_n447_));
  OA220      g425(.A0(new_new_n339_), .A1(new_new_n156_), .B0(new_new_n447_), .B1(new_new_n226_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n90_), .B(i_13_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n415_), .B(new_new_n367_), .Y(new_new_n450_));
  NO2        g428(.A(i_2_), .B(i_13_), .Y(new_new_n451_));
  NA3        g429(.A(new_new_n451_), .B(new_new_n155_), .C(new_new_n93_), .Y(new_new_n452_));
  OAI220     g430(.A0(new_new_n452_), .A1(new_new_n231_), .B0(new_new_n450_), .B1(new_new_n449_), .Y(new_new_n453_));
  NO3        g431(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n454_));
  NO2        g432(.A(i_6_), .B(i_7_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n455_), .B(new_new_n454_), .Y(new_new_n456_));
  NO2        g434(.A(i_11_), .B(i_1_), .Y(new_new_n457_));
  OR2        g435(.A(i_11_), .B(i_8_), .Y(new_new_n458_));
  NOi21      g436(.An(i_2_), .B(i_7_), .Y(new_new_n459_));
  NAi31      g437(.An(new_new_n458_), .B(new_new_n459_), .C(i_0_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n404_), .B(i_6_), .Y(new_new_n461_));
  NA3        g439(.A(new_new_n461_), .B(i_1_), .C(new_new_n70_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n462_), .B(new_new_n460_), .Y(new_new_n463_));
  NO2        g441(.A(i_3_), .B(new_new_n185_), .Y(new_new_n464_));
  NO2        g442(.A(i_6_), .B(i_10_), .Y(new_new_n465_));
  NA4        g443(.A(new_new_n465_), .B(new_new_n302_), .C(new_new_n464_), .D(new_new_n231_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n466_), .B(new_new_n149_), .Y(new_new_n467_));
  NA3        g445(.A(new_new_n238_), .B(new_new_n164_), .C(new_new_n126_), .Y(new_new_n468_));
  NA2        g446(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n469_));
  NO2        g447(.A(new_new_n151_), .B(i_3_), .Y(new_new_n470_));
  NAi31      g448(.An(new_new_n469_), .B(new_new_n470_), .C(new_new_n220_), .Y(new_new_n471_));
  NA3        g449(.A(new_new_n379_), .B(new_new_n171_), .C(new_new_n142_), .Y(new_new_n472_));
  NA3        g450(.A(new_new_n472_), .B(new_new_n471_), .C(new_new_n468_), .Y(new_new_n473_));
  NO4        g451(.A(new_new_n473_), .B(new_new_n467_), .C(new_new_n463_), .D(new_new_n453_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n439_), .B(new_new_n368_), .Y(new_new_n475_));
  NAi21      g453(.An(new_new_n209_), .B(new_new_n385_), .Y(new_new_n476_));
  NO2        g454(.A(new_new_n26_), .B(i_5_), .Y(new_new_n477_));
  NO2        g455(.A(i_0_), .B(new_new_n79_), .Y(new_new_n478_));
  NA3        g456(.A(new_new_n478_), .B(new_new_n477_), .C(new_new_n135_), .Y(new_new_n479_));
  NO2        g457(.A(new_new_n38_), .B(new_new_n479_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n302_), .B(new_new_n232_), .Y(new_new_n481_));
  NO2        g459(.A(new_new_n481_), .B(new_new_n421_), .Y(new_new_n482_));
  NA4        g460(.A(new_new_n296_), .B(new_new_n217_), .C(new_new_n68_), .D(new_new_n231_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n483_), .B(new_new_n456_), .Y(new_new_n484_));
  NO3        g462(.A(new_new_n484_), .B(new_new_n482_), .C(new_new_n480_), .Y(new_new_n485_));
  NA4        g463(.A(new_new_n485_), .B(new_new_n474_), .C(new_new_n448_), .D(new_new_n446_), .Y(new_new_n486_));
  NA3        g464(.A(new_new_n296_), .B(new_new_n168_), .C(new_new_n166_), .Y(new_new_n487_));
  OAI210     g465(.A0(new_new_n291_), .A1(new_new_n172_), .B0(new_new_n487_), .Y(new_new_n488_));
  AN2        g466(.A(new_new_n279_), .B(new_new_n228_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n116_), .B(new_new_n106_), .Y(new_new_n491_));
  AN2        g469(.A(new_new_n491_), .B(new_new_n439_), .Y(new_new_n492_));
  OAI210     g470(.A0(i_2_), .A1(new_new_n226_), .B0(new_new_n297_), .Y(new_new_n493_));
  AOI220     g471(.A0(new_new_n493_), .A1(new_new_n314_), .B0(new_new_n492_), .B1(new_new_n298_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n368_), .B(new_new_n219_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n343_), .B(new_new_n68_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n360_), .B(new_new_n353_), .Y(new_new_n497_));
  OR2        g475(.A(new_new_n495_), .B(new_new_n497_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n36_), .B(i_8_), .Y(new_new_n499_));
  INV        g477(.A(new_new_n498_), .Y(new_new_n500_));
  OAI210     g478(.A0(i_8_), .A1(new_new_n60_), .B0(new_new_n128_), .Y(new_new_n501_));
  INV        g479(.A(new_new_n259_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n502_), .B(new_new_n191_), .Y(new_new_n503_));
  AOI220     g481(.A0(i_6_), .A1(new_new_n503_), .B0(new_new_n501_), .B1(new_new_n405_), .Y(new_new_n504_));
  NA4        g482(.A(new_new_n504_), .B(new_new_n498_), .C(new_new_n494_), .D(new_new_n490_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n374_), .B(new_new_n287_), .Y(new_new_n506_));
  OAI210     g484(.A0(new_new_n370_), .A1(new_new_n162_), .B0(new_new_n506_), .Y(new_new_n507_));
  NO2        g485(.A(i_12_), .B(new_new_n185_), .Y(new_new_n508_));
  NA2        g486(.A(new_new_n508_), .B(new_new_n219_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n404_), .B(new_new_n38_), .Y(new_new_n510_));
  NA2        g488(.A(new_new_n510_), .B(new_new_n507_), .Y(new_new_n511_));
  NO2        g489(.A(i_8_), .B(i_7_), .Y(new_new_n512_));
  AOI220     g490(.A0(new_new_n315_), .A1(new_new_n39_), .B0(new_new_n229_), .B1(new_new_n200_), .Y(new_new_n513_));
  OAI220     g491(.A0(new_new_n513_), .A1(new_new_n174_), .B0(i_5_), .B1(new_new_n236_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n44_), .B(i_10_), .Y(new_new_n515_));
  NO2        g493(.A(new_new_n515_), .B(i_6_), .Y(new_new_n516_));
  NA3        g494(.A(new_new_n516_), .B(new_new_n514_), .C(new_new_n512_), .Y(new_new_n517_));
  AOI220     g495(.A0(new_new_n415_), .A1(new_new_n315_), .B0(new_new_n240_), .B1(new_new_n237_), .Y(new_new_n518_));
  OAI220     g496(.A0(new_new_n518_), .A1(new_new_n256_), .B0(new_new_n449_), .B1(new_new_n127_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n519_), .B(new_new_n259_), .Y(new_new_n520_));
  NOi31      g498(.An(new_new_n282_), .B(new_new_n291_), .C(new_new_n172_), .Y(new_new_n521_));
  NA3        g499(.A(new_new_n296_), .B(new_new_n166_), .C(new_new_n90_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n151_), .B(i_5_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n523_), .B(new_new_n308_), .Y(new_new_n524_));
  NA2        g502(.A(new_new_n524_), .B(new_new_n522_), .Y(new_new_n525_));
  OAI210     g503(.A0(new_new_n525_), .A1(new_new_n521_), .B0(new_new_n444_), .Y(new_new_n526_));
  NA4        g504(.A(new_new_n526_), .B(new_new_n520_), .C(new_new_n517_), .D(new_new_n511_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n276_), .B(new_new_n78_), .Y(new_new_n528_));
  NO2        g506(.A(new_new_n335_), .B(new_new_n528_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n288_), .B(new_new_n279_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n530_), .B(new_new_n165_), .Y(new_new_n531_));
  NA2        g509(.A(new_new_n217_), .B(new_new_n216_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n432_), .B(new_new_n215_), .Y(new_new_n533_));
  NO2        g511(.A(new_new_n532_), .B(new_new_n533_), .Y(new_new_n534_));
  NA3        g512(.A(new_new_n508_), .B(new_new_n267_), .C(i_5_), .Y(new_new_n535_));
  NO2        g513(.A(i_1_), .B(new_new_n535_), .Y(new_new_n536_));
  NO4        g514(.A(new_new_n536_), .B(new_new_n534_), .C(new_new_n531_), .D(new_new_n529_), .Y(new_new_n537_));
  NO4        g515(.A(new_new_n245_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n538_));
  NO3        g516(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n227_), .B(new_new_n36_), .Y(new_new_n540_));
  AN2        g518(.A(new_new_n540_), .B(new_new_n539_), .Y(new_new_n541_));
  OA210      g519(.A0(new_new_n541_), .A1(new_new_n538_), .B0(new_new_n343_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n404_), .B(i_1_), .Y(new_new_n543_));
  NOi31      g521(.An(new_new_n543_), .B(new_new_n440_), .C(new_new_n68_), .Y(new_new_n544_));
  AN3        g522(.A(new_new_n544_), .B(new_new_n402_), .C(new_new_n477_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n413_), .B(new_new_n169_), .Y(new_new_n546_));
  NO3        g524(.A(new_new_n546_), .B(new_new_n545_), .C(new_new_n542_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n79_), .B(new_new_n25_), .Y(new_new_n548_));
  NA2        g526(.A(new_new_n276_), .B(new_new_n548_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n549_), .B(new_new_n438_), .Y(new_new_n550_));
  NO2        g528(.A(new_new_n109_), .B(new_new_n23_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n305_), .Y(new_new_n552_));
  AOI220     g530(.A0(new_new_n552_), .A1(new_new_n422_), .B0(new_new_n175_), .B1(new_new_n173_), .Y(new_new_n553_));
  NOi21      g531(.An(new_new_n139_), .B(new_new_n323_), .Y(new_new_n554_));
  NO3        g532(.A(new_new_n554_), .B(new_new_n553_), .C(new_new_n550_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n496_), .B(new_new_n364_), .Y(new_new_n556_));
  NO2        g534(.A(i_12_), .B(new_new_n79_), .Y(new_new_n557_));
  NA3        g535(.A(new_new_n557_), .B(new_new_n267_), .C(i_5_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n558_), .B(i_3_), .Y(new_new_n559_));
  NA2        g537(.A(new_new_n166_), .B(i_0_), .Y(new_new_n560_));
  NO3        g538(.A(new_new_n560_), .B(new_new_n977_), .C(new_new_n291_), .Y(new_new_n561_));
  OR2        g539(.A(i_2_), .B(i_5_), .Y(new_new_n562_));
  OR2        g540(.A(new_new_n562_), .B(new_new_n397_), .Y(new_new_n563_));
  AOI210     g541(.A0(new_new_n362_), .A1(new_new_n237_), .B0(new_new_n190_), .Y(new_new_n564_));
  AOI210     g542(.A0(new_new_n564_), .A1(new_new_n563_), .B0(new_new_n476_), .Y(new_new_n565_));
  NO4        g543(.A(new_new_n565_), .B(new_new_n561_), .C(new_new_n559_), .D(new_new_n556_), .Y(new_new_n566_));
  NA4        g544(.A(new_new_n566_), .B(new_new_n555_), .C(new_new_n547_), .D(new_new_n537_), .Y(new_new_n567_));
  NO4        g545(.A(new_new_n567_), .B(new_new_n527_), .C(new_new_n505_), .D(new_new_n486_), .Y(new_new_n568_));
  NA4        g546(.A(new_new_n568_), .B(new_new_n430_), .C(new_new_n342_), .D(new_new_n301_), .Y(men7));
  NO2        g547(.A(new_new_n86_), .B(new_new_n52_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n102_), .B(new_new_n83_), .Y(new_new_n571_));
  NA2        g549(.A(new_new_n369_), .B(new_new_n571_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n465_), .B(new_new_n78_), .Y(new_new_n573_));
  NA2        g551(.A(new_new_n137_), .B(i_8_), .Y(new_new_n574_));
  OAI210     g552(.A0(new_new_n574_), .A1(new_new_n573_), .B0(new_new_n572_), .Y(new_new_n575_));
  NA3        g553(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n576_));
  NO2        g554(.A(new_new_n231_), .B(i_4_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n577_), .B(i_8_), .Y(new_new_n578_));
  NA2        g556(.A(i_2_), .B(new_new_n79_), .Y(new_new_n579_));
  OAI210     g557(.A0(new_new_n82_), .A1(new_new_n195_), .B0(new_new_n196_), .Y(new_new_n580_));
  NA2        g558(.A(i_4_), .B(i_8_), .Y(new_new_n581_));
  NA2        g559(.A(new_new_n581_), .B(new_new_n296_), .Y(new_new_n582_));
  OAI220     g560(.A0(new_new_n582_), .A1(new_new_n579_), .B0(new_new_n580_), .B1(i_13_), .Y(new_new_n583_));
  NO3        g561(.A(new_new_n583_), .B(new_new_n575_), .C(new_new_n570_), .Y(new_new_n584_));
  AOI210     g562(.A0(new_new_n122_), .A1(new_new_n59_), .B0(i_10_), .Y(new_new_n585_));
  AOI210     g563(.A0(new_new_n585_), .A1(new_new_n231_), .B0(new_new_n155_), .Y(new_new_n586_));
  OR2        g564(.A(i_6_), .B(i_10_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n587_), .B(new_new_n23_), .Y(new_new_n588_));
  OR3        g566(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n589_));
  NO3        g567(.A(new_new_n589_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n590_));
  INV        g568(.A(new_new_n192_), .Y(new_new_n591_));
  INV        g569(.A(new_new_n590_), .Y(new_new_n592_));
  OA220      g570(.A0(new_new_n592_), .A1(i_3_), .B0(new_new_n586_), .B1(new_new_n261_), .Y(new_new_n593_));
  AOI210     g571(.A0(new_new_n593_), .A1(new_new_n584_), .B0(new_new_n60_), .Y(new_new_n594_));
  NOi21      g572(.An(i_11_), .B(i_7_), .Y(new_new_n595_));
  AO210      g573(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n596_));
  NO2        g574(.A(new_new_n596_), .B(new_new_n595_), .Y(new_new_n597_));
  NA3        g575(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n598_));
  NAi31      g576(.An(new_new_n598_), .B(new_new_n208_), .C(i_11_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n599_), .B(new_new_n60_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n81_), .B(new_new_n60_), .Y(new_new_n601_));
  AO210      g579(.A0(new_new_n601_), .A1(new_new_n364_), .B0(new_new_n40_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n60_), .B(i_9_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n60_), .B(new_new_n985_), .Y(new_new_n604_));
  NO2        g582(.A(i_1_), .B(i_12_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n604_), .B(new_new_n602_), .Y(new_new_n606_));
  OAI210     g584(.A0(new_new_n606_), .A1(new_new_n600_), .B0(i_6_), .Y(new_new_n607_));
  NO2        g585(.A(i_6_), .B(i_11_), .Y(new_new_n608_));
  INV        g586(.A(new_new_n441_), .Y(new_new_n609_));
  NO4        g587(.A(new_new_n208_), .B(new_new_n122_), .C(i_13_), .D(new_new_n79_), .Y(new_new_n610_));
  NA2        g588(.A(new_new_n610_), .B(new_new_n603_), .Y(new_new_n611_));
  NO3        g589(.A(new_new_n587_), .B(new_new_n227_), .C(new_new_n23_), .Y(new_new_n612_));
  AOI210     g590(.A0(i_1_), .A1(new_new_n252_), .B0(new_new_n612_), .Y(new_new_n613_));
  OAI210     g591(.A0(new_new_n613_), .A1(new_new_n44_), .B0(new_new_n611_), .Y(new_new_n614_));
  NA3        g592(.A(new_new_n512_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n615_));
  NA2        g593(.A(new_new_n132_), .B(i_9_), .Y(new_new_n616_));
  NA3        g594(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n46_), .B(i_1_), .Y(new_new_n618_));
  NA3        g596(.A(new_new_n618_), .B(new_new_n260_), .C(new_new_n44_), .Y(new_new_n619_));
  OAI220     g597(.A0(new_new_n619_), .A1(new_new_n617_), .B0(new_new_n616_), .B1(new_new_n974_), .Y(new_new_n620_));
  NA3        g598(.A(new_new_n603_), .B(new_new_n308_), .C(i_6_), .Y(new_new_n621_));
  NO2        g599(.A(new_new_n621_), .B(new_new_n23_), .Y(new_new_n622_));
  AOI210     g600(.A0(new_new_n457_), .A1(new_new_n407_), .B0(new_new_n235_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n623_), .B(new_new_n579_), .Y(new_new_n624_));
  NAi21      g602(.An(new_new_n615_), .B(new_new_n85_), .Y(new_new_n625_));
  NA2        g603(.A(new_new_n618_), .B(new_new_n260_), .Y(new_new_n626_));
  NO2        g604(.A(i_11_), .B(new_new_n37_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n627_), .B(new_new_n24_), .Y(new_new_n628_));
  OAI210     g606(.A0(new_new_n628_), .A1(new_new_n626_), .B0(new_new_n625_), .Y(new_new_n629_));
  OR4        g607(.A(new_new_n629_), .B(new_new_n624_), .C(new_new_n622_), .D(new_new_n620_), .Y(new_new_n630_));
  NO3        g608(.A(new_new_n630_), .B(new_new_n614_), .C(new_new_n609_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n231_), .B(new_new_n95_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n632_), .B(new_new_n595_), .Y(new_new_n633_));
  NA2        g611(.A(new_new_n633_), .B(i_1_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n634_), .B(new_new_n589_), .Y(new_new_n635_));
  NA2        g613(.A(new_new_n635_), .B(new_new_n46_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n980_), .B(new_new_n109_), .Y(new_new_n637_));
  AN2        g615(.A(new_new_n637_), .B(new_new_n516_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n227_), .B(new_new_n44_), .Y(new_new_n639_));
  NO3        g617(.A(new_new_n639_), .B(new_new_n298_), .C(i_11_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n111_), .B(new_new_n37_), .Y(new_new_n641_));
  NO2        g619(.A(new_new_n641_), .B(i_6_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n79_), .B(i_9_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n643_), .B(new_new_n60_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n644_), .B(new_new_n605_), .Y(new_new_n645_));
  NO4        g623(.A(new_new_n645_), .B(new_new_n642_), .C(new_new_n640_), .D(i_4_), .Y(new_new_n646_));
  NA2        g624(.A(i_1_), .B(i_3_), .Y(new_new_n647_));
  NO2        g625(.A(new_new_n442_), .B(new_new_n86_), .Y(new_new_n648_));
  AOI210     g626(.A0(new_new_n639_), .A1(i_10_), .B0(new_new_n648_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n649_), .B(new_new_n647_), .Y(new_new_n650_));
  NO3        g628(.A(new_new_n650_), .B(new_new_n646_), .C(new_new_n638_), .Y(new_new_n651_));
  NA4        g629(.A(new_new_n651_), .B(new_new_n636_), .C(new_new_n631_), .D(new_new_n607_), .Y(new_new_n652_));
  NO3        g630(.A(new_new_n458_), .B(i_3_), .C(i_7_), .Y(new_new_n653_));
  NOi21      g631(.An(new_new_n653_), .B(i_10_), .Y(new_new_n654_));
  AN2        g632(.A(new_new_n238_), .B(new_new_n79_), .Y(new_new_n655_));
  NA2        g633(.A(new_new_n360_), .B(new_new_n359_), .Y(new_new_n656_));
  NA3        g634(.A(new_new_n465_), .B(new_new_n499_), .C(new_new_n46_), .Y(new_new_n657_));
  NO3        g635(.A(new_new_n459_), .B(new_new_n581_), .C(new_new_n79_), .Y(new_new_n658_));
  NA2        g636(.A(new_new_n658_), .B(new_new_n25_), .Y(new_new_n659_));
  NA3        g637(.A(new_new_n155_), .B(new_new_n78_), .C(new_new_n79_), .Y(new_new_n660_));
  NA4        g638(.A(new_new_n660_), .B(new_new_n659_), .C(new_new_n657_), .D(new_new_n656_), .Y(new_new_n661_));
  OAI210     g639(.A0(new_new_n661_), .A1(new_new_n655_), .B0(i_1_), .Y(new_new_n662_));
  AOI210     g640(.A0(new_new_n260_), .A1(new_new_n91_), .B0(i_1_), .Y(new_new_n663_));
  NO2        g641(.A(new_new_n358_), .B(i_2_), .Y(new_new_n664_));
  NA2        g642(.A(new_new_n664_), .B(new_new_n663_), .Y(new_new_n665_));
  OAI210     g643(.A0(new_new_n621_), .A1(new_new_n433_), .B0(new_new_n665_), .Y(new_new_n666_));
  INV        g644(.A(new_new_n666_), .Y(new_new_n667_));
  AOI210     g645(.A0(new_new_n667_), .A1(new_new_n662_), .B0(i_13_), .Y(new_new_n668_));
  OR2        g646(.A(i_11_), .B(i_7_), .Y(new_new_n669_));
  NA3        g647(.A(new_new_n669_), .B(new_new_n100_), .C(new_new_n132_), .Y(new_new_n670_));
  AOI220     g648(.A0(new_new_n451_), .A1(new_new_n155_), .B0(new_new_n435_), .B1(new_new_n132_), .Y(new_new_n671_));
  OAI210     g649(.A0(new_new_n671_), .A1(new_new_n44_), .B0(new_new_n670_), .Y(new_new_n672_));
  NA2        g650(.A(new_new_n238_), .B(new_new_n125_), .Y(new_new_n673_));
  NO2        g651(.A(new_new_n673_), .B(new_new_n40_), .Y(new_new_n674_));
  AOI210     g652(.A0(new_new_n672_), .A1(new_new_n325_), .B0(new_new_n674_), .Y(new_new_n675_));
  AOI220     g653(.A0(i_7_), .A1(new_new_n67_), .B0(new_new_n371_), .B1(new_new_n618_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n676_), .B(new_new_n236_), .Y(new_new_n677_));
  NA2        g655(.A(new_new_n121_), .B(i_13_), .Y(new_new_n678_));
  NO2        g656(.A(new_new_n617_), .B(new_new_n109_), .Y(new_new_n679_));
  INV        g657(.A(new_new_n679_), .Y(new_new_n680_));
  OAI220     g658(.A0(new_new_n680_), .A1(new_new_n66_), .B0(new_new_n678_), .B1(new_new_n663_), .Y(new_new_n681_));
  NO3        g659(.A(new_new_n66_), .B(new_new_n32_), .C(new_new_n95_), .Y(new_new_n682_));
  NA2        g660(.A(new_new_n26_), .B(new_new_n185_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n683_), .B(i_7_), .Y(new_new_n684_));
  NO3        g662(.A(new_new_n459_), .B(new_new_n231_), .C(new_new_n79_), .Y(new_new_n685_));
  AOI210     g663(.A0(new_new_n685_), .A1(new_new_n684_), .B0(new_new_n682_), .Y(new_new_n686_));
  NO2        g664(.A(new_new_n686_), .B(new_new_n591_), .Y(new_new_n687_));
  NO3        g665(.A(new_new_n687_), .B(new_new_n681_), .C(new_new_n677_), .Y(new_new_n688_));
  OR2        g666(.A(i_11_), .B(i_6_), .Y(new_new_n689_));
  NA3        g667(.A(new_new_n577_), .B(new_new_n683_), .C(i_7_), .Y(new_new_n690_));
  AOI210     g668(.A0(new_new_n690_), .A1(new_new_n680_), .B0(new_new_n689_), .Y(new_new_n691_));
  NA2        g669(.A(new_new_n608_), .B(i_13_), .Y(new_new_n692_));
  NA2        g670(.A(new_new_n96_), .B(new_new_n683_), .Y(new_new_n693_));
  NAi21      g671(.An(i_11_), .B(i_12_), .Y(new_new_n694_));
  NOi41      g672(.An(new_new_n105_), .B(new_new_n694_), .C(i_13_), .D(new_new_n79_), .Y(new_new_n695_));
  NO2        g673(.A(new_new_n459_), .B(new_new_n581_), .Y(new_new_n696_));
  AOI220     g674(.A0(new_new_n696_), .A1(new_new_n302_), .B0(new_new_n695_), .B1(new_new_n693_), .Y(new_new_n697_));
  NA2        g675(.A(new_new_n697_), .B(new_new_n692_), .Y(new_new_n698_));
  OAI210     g676(.A0(new_new_n698_), .A1(new_new_n691_), .B0(new_new_n60_), .Y(new_new_n699_));
  NO2        g677(.A(i_2_), .B(i_12_), .Y(new_new_n700_));
  NA2        g678(.A(new_new_n357_), .B(new_new_n700_), .Y(new_new_n701_));
  OAI210     g679(.A0(i_8_), .A1(new_new_n359_), .B0(new_new_n357_), .Y(new_new_n702_));
  NO2        g680(.A(new_new_n122_), .B(i_2_), .Y(new_new_n703_));
  NA2        g681(.A(new_new_n703_), .B(new_new_n605_), .Y(new_new_n704_));
  NA3        g682(.A(new_new_n704_), .B(new_new_n702_), .C(new_new_n701_), .Y(new_new_n705_));
  NA3        g683(.A(new_new_n705_), .B(new_new_n45_), .C(new_new_n219_), .Y(new_new_n706_));
  NA4        g684(.A(new_new_n706_), .B(new_new_n699_), .C(new_new_n688_), .D(new_new_n675_), .Y(new_new_n707_));
  OR4        g685(.A(new_new_n707_), .B(new_new_n668_), .C(new_new_n652_), .D(new_new_n594_), .Y(men5));
  AOI210     g686(.A0(new_new_n633_), .A1(new_new_n263_), .B0(new_new_n405_), .Y(new_new_n709_));
  NO2        g687(.A(new_new_n578_), .B(i_11_), .Y(new_new_n710_));
  NA2        g688(.A(new_new_n82_), .B(new_new_n710_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n711_), .B(new_new_n709_), .Y(new_new_n712_));
  NO3        g690(.A(i_11_), .B(new_new_n231_), .C(i_13_), .Y(new_new_n713_));
  NO2        g691(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n714_));
  NA2        g692(.A(i_12_), .B(i_8_), .Y(new_new_n715_));
  INV        g693(.A(new_new_n715_), .Y(new_new_n716_));
  INV        g694(.A(new_new_n432_), .Y(new_new_n717_));
  AOI220     g695(.A0(new_new_n308_), .A1(new_new_n551_), .B0(new_new_n716_), .B1(new_new_n714_), .Y(new_new_n718_));
  INV        g696(.A(new_new_n718_), .Y(new_new_n719_));
  NO2        g697(.A(new_new_n719_), .B(new_new_n712_), .Y(new_new_n720_));
  INV        g698(.A(new_new_n164_), .Y(new_new_n721_));
  OAI210     g699(.A0(new_new_n664_), .A1(new_new_n434_), .B0(new_new_n105_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n722_), .B(new_new_n721_), .Y(new_new_n723_));
  NO2        g701(.A(new_new_n442_), .B(new_new_n26_), .Y(new_new_n724_));
  NO2        g702(.A(new_new_n724_), .B(new_new_n407_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n725_), .B(i_2_), .Y(new_new_n726_));
  INV        g704(.A(new_new_n726_), .Y(new_new_n727_));
  AOI210     g705(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n404_), .Y(new_new_n728_));
  AOI210     g706(.A0(new_new_n728_), .A1(new_new_n727_), .B0(new_new_n723_), .Y(new_new_n729_));
  OA210      g707(.A0(new_new_n597_), .A1(new_new_n120_), .B0(i_13_), .Y(new_new_n730_));
  NA2        g708(.A(new_new_n192_), .B(new_new_n195_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n145_), .B(i_8_), .Y(new_new_n732_));
  AOI210     g710(.A0(new_new_n732_), .A1(new_new_n731_), .B0(new_new_n362_), .Y(new_new_n733_));
  AOI210     g711(.A0(new_new_n201_), .A1(new_new_n141_), .B0(new_new_n499_), .Y(new_new_n734_));
  NA2        g712(.A(new_new_n734_), .B(new_new_n407_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n96_), .B(new_new_n44_), .Y(new_new_n736_));
  INV        g714(.A(new_new_n292_), .Y(new_new_n737_));
  NA4        g715(.A(new_new_n737_), .B(new_new_n296_), .C(new_new_n118_), .D(new_new_n42_), .Y(new_new_n738_));
  OAI210     g716(.A0(new_new_n738_), .A1(new_new_n736_), .B0(new_new_n735_), .Y(new_new_n739_));
  NO3        g717(.A(new_new_n739_), .B(new_new_n733_), .C(new_new_n730_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n551_), .B(new_new_n28_), .Y(new_new_n741_));
  NA2        g719(.A(new_new_n713_), .B(new_new_n268_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n742_), .B(new_new_n741_), .Y(new_new_n743_));
  AOI220     g721(.A0(new_new_n120_), .A1(new_new_n36_), .B0(new_new_n743_), .B1(new_new_n46_), .Y(new_new_n744_));
  NA4        g722(.A(new_new_n744_), .B(new_new_n740_), .C(new_new_n729_), .D(new_new_n720_), .Y(men6));
  NA2        g723(.A(new_new_n981_), .B(new_new_n703_), .Y(new_new_n746_));
  NA4        g724(.A(new_new_n375_), .B(new_new_n464_), .C(new_new_n66_), .D(new_new_n95_), .Y(new_new_n747_));
  INV        g725(.A(new_new_n747_), .Y(new_new_n748_));
  NO2        g726(.A(new_new_n214_), .B(new_new_n469_), .Y(new_new_n749_));
  INV        g727(.A(i_9_), .Y(new_new_n750_));
  NO2        g728(.A(new_new_n748_), .B(new_new_n320_), .Y(new_new_n751_));
  AO210      g729(.A0(new_new_n751_), .A1(new_new_n746_), .B0(i_12_), .Y(new_new_n752_));
  NA2        g730(.A(new_new_n363_), .B(new_new_n328_), .Y(new_new_n753_));
  NA2        g731(.A(new_new_n557_), .B(new_new_n60_), .Y(new_new_n754_));
  NA2        g732(.A(new_new_n654_), .B(new_new_n66_), .Y(new_new_n755_));
  NA4        g733(.A(new_new_n601_), .B(new_new_n755_), .C(new_new_n754_), .D(new_new_n753_), .Y(new_new_n756_));
  INV        g734(.A(new_new_n189_), .Y(new_new_n757_));
  AOI220     g735(.A0(new_new_n757_), .A1(new_new_n750_), .B0(new_new_n756_), .B1(new_new_n68_), .Y(new_new_n758_));
  INV        g736(.A(new_new_n319_), .Y(new_new_n759_));
  NA2        g737(.A(new_new_n70_), .B(new_new_n125_), .Y(new_new_n760_));
  AOI210     g738(.A0(new_new_n118_), .A1(new_new_n760_), .B0(new_new_n759_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n497_), .B(new_new_n177_), .Y(new_new_n762_));
  INV        g740(.A(i_11_), .Y(new_new_n763_));
  NA3        g741(.A(new_new_n763_), .B(new_new_n455_), .C(new_new_n375_), .Y(new_new_n764_));
  NAi32      g742(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n765_));
  NO2        g743(.A(new_new_n689_), .B(new_new_n765_), .Y(new_new_n766_));
  OAI210     g744(.A0(new_new_n653_), .A1(new_new_n540_), .B0(new_new_n539_), .Y(new_new_n767_));
  NAi31      g745(.An(new_new_n766_), .B(new_new_n767_), .C(new_new_n764_), .Y(new_new_n768_));
  OR3        g746(.A(new_new_n768_), .B(new_new_n762_), .C(new_new_n761_), .Y(new_new_n769_));
  NA3        g747(.A(new_new_n338_), .B(new_new_n248_), .C(i_7_), .Y(new_new_n770_));
  OR2        g748(.A(new_new_n597_), .B(new_new_n434_), .Y(new_new_n771_));
  NA2        g749(.A(new_new_n771_), .B(new_new_n140_), .Y(new_new_n772_));
  OR2        g750(.A(new_new_n717_), .B(new_new_n36_), .Y(new_new_n773_));
  NA3        g751(.A(new_new_n773_), .B(new_new_n772_), .C(new_new_n770_), .Y(new_new_n774_));
  AOI220     g752(.A0(new_new_n979_), .A1(new_new_n539_), .B0(new_new_n749_), .B1(new_new_n684_), .Y(new_new_n775_));
  NA3        g753(.A(new_new_n362_), .B(new_new_n232_), .C(new_new_n140_), .Y(new_new_n776_));
  NA2        g754(.A(new_new_n382_), .B(new_new_n65_), .Y(new_new_n777_));
  NA4        g755(.A(new_new_n777_), .B(new_new_n776_), .C(new_new_n775_), .D(new_new_n580_), .Y(new_new_n778_));
  AO210      g756(.A0(new_new_n499_), .A1(new_new_n46_), .B0(new_new_n81_), .Y(new_new_n779_));
  NA3        g757(.A(new_new_n779_), .B(new_new_n465_), .C(new_new_n211_), .Y(new_new_n780_));
  AOI210     g758(.A0(new_new_n434_), .A1(new_new_n432_), .B0(new_new_n538_), .Y(new_new_n781_));
  NO2        g759(.A(new_new_n587_), .B(new_new_n96_), .Y(new_new_n782_));
  OAI210     g760(.A0(new_new_n782_), .A1(new_new_n106_), .B0(new_new_n396_), .Y(new_new_n783_));
  NA2        g761(.A(new_new_n237_), .B(new_new_n46_), .Y(new_new_n784_));
  INV        g762(.A(new_new_n563_), .Y(new_new_n785_));
  NA3        g763(.A(new_new_n785_), .B(new_new_n319_), .C(i_7_), .Y(new_new_n786_));
  NA4        g764(.A(new_new_n786_), .B(new_new_n783_), .C(new_new_n781_), .D(new_new_n780_), .Y(new_new_n787_));
  NO4        g765(.A(new_new_n787_), .B(new_new_n778_), .C(new_new_n774_), .D(new_new_n769_), .Y(new_new_n788_));
  NA4        g766(.A(new_new_n788_), .B(new_new_n758_), .C(new_new_n752_), .D(new_new_n365_), .Y(men3));
  NA2        g767(.A(i_12_), .B(i_10_), .Y(new_new_n790_));
  NA2        g768(.A(i_6_), .B(i_7_), .Y(new_new_n791_));
  NO2        g769(.A(new_new_n791_), .B(i_0_), .Y(new_new_n792_));
  NO2        g770(.A(i_11_), .B(new_new_n231_), .Y(new_new_n793_));
  NO3        g771(.A(new_new_n438_), .B(new_new_n83_), .C(new_new_n44_), .Y(new_new_n794_));
  AN2        g772(.A(new_new_n794_), .B(new_new_n166_), .Y(new_new_n795_));
  NA3        g773(.A(new_new_n776_), .B(new_new_n580_), .C(new_new_n361_), .Y(new_new_n796_));
  NA2        g774(.A(new_new_n796_), .B(new_new_n39_), .Y(new_new_n797_));
  NO3        g775(.A(new_new_n201_), .B(new_new_n442_), .C(new_new_n125_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n398_), .B(new_new_n45_), .Y(new_new_n799_));
  AN2        g777(.A(new_new_n440_), .B(new_new_n53_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n800_), .B(new_new_n798_), .Y(new_new_n801_));
  AOI210     g779(.A0(new_new_n801_), .A1(new_new_n797_), .B0(new_new_n48_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n984_), .B(new_new_n643_), .Y(new_new_n803_));
  NA2        g781(.A(new_new_n326_), .B(new_new_n424_), .Y(new_new_n804_));
  NO2        g782(.A(new_new_n804_), .B(new_new_n803_), .Y(new_new_n805_));
  NOi21      g783(.An(i_5_), .B(i_9_), .Y(new_new_n806_));
  NA2        g784(.A(new_new_n806_), .B(new_new_n431_), .Y(new_new_n807_));
  AOI210     g785(.A0(new_new_n260_), .A1(new_new_n457_), .B0(new_new_n658_), .Y(new_new_n808_));
  NO2        g786(.A(new_new_n808_), .B(new_new_n807_), .Y(new_new_n809_));
  NO4        g787(.A(new_new_n809_), .B(new_new_n805_), .C(new_new_n802_), .D(new_new_n795_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n177_), .B(new_new_n24_), .Y(new_new_n811_));
  INV        g789(.A(new_new_n641_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n812_), .B(new_new_n811_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n302_), .B(new_new_n123_), .Y(new_new_n814_));
  NAi21      g792(.An(new_new_n156_), .B(new_new_n424_), .Y(new_new_n815_));
  OAI220     g793(.A0(new_new_n815_), .A1(new_new_n784_), .B0(new_new_n814_), .B1(new_new_n388_), .Y(new_new_n816_));
  NO2        g794(.A(new_new_n816_), .B(new_new_n813_), .Y(new_new_n817_));
  NA2        g795(.A(new_new_n548_), .B(i_0_), .Y(new_new_n818_));
  NO3        g796(.A(new_new_n818_), .B(new_new_n370_), .C(new_new_n82_), .Y(new_new_n819_));
  NO4        g797(.A(new_new_n562_), .B(new_new_n208_), .C(new_new_n404_), .D(new_new_n397_), .Y(new_new_n820_));
  AOI210     g798(.A0(new_new_n820_), .A1(i_11_), .B0(new_new_n819_), .Y(new_new_n821_));
  NA2        g799(.A(new_new_n713_), .B(new_new_n320_), .Y(new_new_n822_));
  AOI210     g800(.A0(new_new_n465_), .A1(new_new_n82_), .B0(new_new_n55_), .Y(new_new_n823_));
  OAI220     g801(.A0(new_new_n823_), .A1(new_new_n822_), .B0(new_new_n628_), .B1(i_5_), .Y(new_new_n824_));
  NA2        g802(.A(i_0_), .B(i_10_), .Y(new_new_n825_));
  AOI220     g803(.A0(new_new_n326_), .A1(new_new_n92_), .B0(new_new_n177_), .B1(new_new_n78_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n543_), .B(i_4_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n180_), .B(new_new_n195_), .Y(new_new_n828_));
  OAI220     g806(.A0(new_new_n828_), .A1(new_new_n822_), .B0(new_new_n827_), .B1(new_new_n826_), .Y(new_new_n829_));
  NO2        g807(.A(new_new_n829_), .B(new_new_n824_), .Y(new_new_n830_));
  NA3        g808(.A(new_new_n830_), .B(new_new_n821_), .C(new_new_n817_), .Y(new_new_n831_));
  NO2        g809(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n832_));
  NA2        g810(.A(i_11_), .B(i_9_), .Y(new_new_n833_));
  NO3        g811(.A(i_12_), .B(new_new_n833_), .C(new_new_n579_), .Y(new_new_n834_));
  AN2        g812(.A(new_new_n834_), .B(new_new_n832_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n379_), .B(new_new_n171_), .Y(new_new_n836_));
  NA2        g814(.A(new_new_n836_), .B(new_new_n154_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n833_), .B(new_new_n68_), .Y(new_new_n838_));
  NO2        g816(.A(new_new_n167_), .B(i_0_), .Y(new_new_n839_));
  AOI210     g817(.A0(new_new_n360_), .A1(new_new_n41_), .B0(new_new_n395_), .Y(new_new_n840_));
  NO2        g818(.A(new_new_n840_), .B(new_new_n807_), .Y(new_new_n841_));
  NO3        g819(.A(new_new_n841_), .B(new_new_n837_), .C(new_new_n835_), .Y(new_new_n842_));
  NA2        g820(.A(new_new_n627_), .B(new_new_n115_), .Y(new_new_n843_));
  NO2        g821(.A(i_6_), .B(new_new_n843_), .Y(new_new_n844_));
  AOI210     g822(.A0(new_new_n433_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n845_));
  NA2        g823(.A(new_new_n164_), .B(new_new_n97_), .Y(new_new_n846_));
  NOi32      g824(.An(new_new_n845_), .Bn(new_new_n180_), .C(new_new_n846_), .Y(new_new_n847_));
  NO2        g825(.A(new_new_n976_), .B(new_new_n799_), .Y(new_new_n848_));
  NO3        g826(.A(new_new_n848_), .B(new_new_n847_), .C(new_new_n844_), .Y(new_new_n849_));
  NOi21      g827(.An(i_7_), .B(i_5_), .Y(new_new_n850_));
  NOi31      g828(.An(new_new_n850_), .B(i_0_), .C(new_new_n694_), .Y(new_new_n851_));
  NA3        g829(.A(new_new_n851_), .B(new_new_n369_), .C(i_6_), .Y(new_new_n852_));
  OA210      g830(.A0(new_new_n846_), .A1(new_new_n497_), .B0(new_new_n852_), .Y(new_new_n853_));
  NO3        g831(.A(new_new_n391_), .B(new_new_n350_), .C(new_new_n346_), .Y(new_new_n854_));
  INV        g832(.A(new_new_n309_), .Y(new_new_n855_));
  NO2        g833(.A(new_new_n694_), .B(new_new_n250_), .Y(new_new_n856_));
  AOI210     g834(.A0(new_new_n856_), .A1(new_new_n855_), .B0(new_new_n854_), .Y(new_new_n857_));
  NA4        g835(.A(new_new_n857_), .B(new_new_n853_), .C(new_new_n849_), .D(new_new_n842_), .Y(new_new_n858_));
  AN2        g836(.A(new_new_n325_), .B(new_new_n320_), .Y(new_new_n859_));
  NO2        g837(.A(new_new_n790_), .B(new_new_n308_), .Y(new_new_n860_));
  BUFFER     g838(.A(new_new_n454_), .Y(new_new_n861_));
  NA2        g839(.A(new_new_n860_), .B(new_new_n838_), .Y(new_new_n862_));
  NO2        g840(.A(new_new_n815_), .B(i_6_), .Y(new_new_n863_));
  NA2        g841(.A(new_new_n838_), .B(new_new_n296_), .Y(new_new_n864_));
  NA2        g842(.A(new_new_n179_), .B(new_new_n864_), .Y(new_new_n865_));
  AOI220     g843(.A0(new_new_n865_), .A1(new_new_n455_), .B0(new_new_n863_), .B1(new_new_n68_), .Y(new_new_n866_));
  NO2        g844(.A(new_new_n70_), .B(new_new_n715_), .Y(new_new_n867_));
  INV        g845(.A(new_new_n867_), .Y(new_new_n868_));
  NO2        g846(.A(new_new_n868_), .B(new_new_n47_), .Y(new_new_n869_));
  NO3        g847(.A(new_new_n562_), .B(new_new_n345_), .C(new_new_n24_), .Y(new_new_n870_));
  INV        g848(.A(new_new_n870_), .Y(new_new_n871_));
  NAi21      g849(.An(i_9_), .B(i_5_), .Y(new_new_n872_));
  NO2        g850(.A(new_new_n872_), .B(new_new_n391_), .Y(new_new_n873_));
  NO2        g851(.A(new_new_n576_), .B(new_new_n99_), .Y(new_new_n874_));
  AOI220     g852(.A0(new_new_n874_), .A1(i_0_), .B0(new_new_n873_), .B1(new_new_n597_), .Y(new_new_n875_));
  OAI220     g853(.A0(new_new_n875_), .A1(new_new_n79_), .B0(new_new_n871_), .B1(new_new_n165_), .Y(new_new_n876_));
  NO3        g854(.A(new_new_n876_), .B(new_new_n869_), .C(new_new_n500_), .Y(new_new_n877_));
  NA3        g855(.A(new_new_n877_), .B(new_new_n866_), .C(new_new_n862_), .Y(new_new_n878_));
  NO3        g856(.A(new_new_n878_), .B(new_new_n858_), .C(new_new_n831_), .Y(new_new_n879_));
  NO2        g857(.A(i_0_), .B(new_new_n694_), .Y(new_new_n880_));
  NA2        g858(.A(new_new_n68_), .B(new_new_n44_), .Y(new_new_n881_));
  AN2        g859(.A(new_new_n880_), .B(new_new_n166_), .Y(new_new_n882_));
  NO2        g860(.A(new_new_n754_), .B(new_new_n846_), .Y(new_new_n883_));
  AOI210     g861(.A0(new_new_n882_), .A1(i_8_), .B0(new_new_n883_), .Y(new_new_n884_));
  NA2        g862(.A(new_new_n703_), .B(new_new_n139_), .Y(new_new_n885_));
  INV        g863(.A(new_new_n885_), .Y(new_new_n886_));
  NA2        g864(.A(new_new_n886_), .B(new_new_n643_), .Y(new_new_n887_));
  NO2        g865(.A(new_new_n767_), .B(new_new_n391_), .Y(new_new_n888_));
  NA3        g866(.A(new_new_n792_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n889_));
  NA2        g867(.A(new_new_n793_), .B(i_9_), .Y(new_new_n890_));
  AOI210     g868(.A0(new_new_n889_), .A1(new_new_n479_), .B0(new_new_n890_), .Y(new_new_n891_));
  OAI210     g869(.A0(new_new_n237_), .A1(i_9_), .B0(new_new_n224_), .Y(new_new_n892_));
  AOI210     g870(.A0(new_new_n892_), .A1(new_new_n818_), .B0(new_new_n147_), .Y(new_new_n893_));
  NO3        g871(.A(new_new_n893_), .B(new_new_n891_), .C(new_new_n888_), .Y(new_new_n894_));
  NA3        g872(.A(new_new_n894_), .B(new_new_n887_), .C(new_new_n884_), .Y(new_new_n895_));
  INV        g873(.A(new_new_n859_), .Y(new_new_n896_));
  AOI210     g874(.A0(new_new_n291_), .A1(new_new_n156_), .B0(new_new_n896_), .Y(new_new_n897_));
  NA3        g875(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n898_));
  NA2        g876(.A(i_5_), .B(new_new_n470_), .Y(new_new_n899_));
  AOI210     g877(.A0(new_new_n898_), .A1(new_new_n156_), .B0(new_new_n899_), .Y(new_new_n900_));
  NO2        g878(.A(new_new_n900_), .B(new_new_n897_), .Y(new_new_n901_));
  NO3        g879(.A(new_new_n825_), .B(new_new_n806_), .C(new_new_n182_), .Y(new_new_n902_));
  AOI220     g880(.A0(new_new_n902_), .A1(i_11_), .B0(new_new_n544_), .B1(new_new_n70_), .Y(new_new_n903_));
  NO3        g881(.A(new_new_n202_), .B(new_new_n368_), .C(i_0_), .Y(new_new_n904_));
  OAI210     g882(.A0(new_new_n904_), .A1(new_new_n71_), .B0(i_13_), .Y(new_new_n905_));
  OAI220     g883(.A0(new_new_n509_), .A1(new_new_n982_), .B0(i_12_), .B1(new_new_n591_), .Y(new_new_n906_));
  NA3        g884(.A(new_new_n906_), .B(new_new_n383_), .C(i_0_), .Y(new_new_n907_));
  NA4        g885(.A(new_new_n907_), .B(new_new_n905_), .C(new_new_n903_), .D(new_new_n901_), .Y(new_new_n908_));
  NO2        g886(.A(new_new_n236_), .B(new_new_n86_), .Y(new_new_n909_));
  AOI210     g887(.A0(new_new_n909_), .A1(new_new_n880_), .B0(new_new_n103_), .Y(new_new_n910_));
  AOI210     g888(.A0(new_new_n792_), .A1(new_new_n157_), .B0(new_new_n470_), .Y(new_new_n911_));
  NA2        g889(.A(new_new_n338_), .B(new_new_n168_), .Y(new_new_n912_));
  OA220      g890(.A0(new_new_n912_), .A1(new_new_n911_), .B0(new_new_n910_), .B1(i_5_), .Y(new_new_n913_));
  AOI210     g891(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n167_), .Y(new_new_n914_));
  NA2        g892(.A(new_new_n914_), .B(new_new_n861_), .Y(new_new_n915_));
  NA3        g893(.A(new_new_n475_), .B(new_new_n468_), .C(new_new_n452_), .Y(new_new_n916_));
  INV        g894(.A(new_new_n916_), .Y(new_new_n917_));
  NA3        g895(.A(new_new_n375_), .B(new_new_n164_), .C(new_new_n163_), .Y(new_new_n918_));
  NA3        g896(.A(new_new_n375_), .B(new_new_n327_), .C(new_new_n215_), .Y(new_new_n919_));
  INV        g897(.A(new_new_n919_), .Y(new_new_n920_));
  NOi31      g898(.An(new_new_n374_), .B(new_new_n881_), .C(new_new_n233_), .Y(new_new_n921_));
  NO3        g899(.A(new_new_n921_), .B(new_new_n920_), .C(new_new_n975_), .Y(new_new_n922_));
  NA4        g900(.A(new_new_n922_), .B(new_new_n917_), .C(new_new_n915_), .D(new_new_n913_), .Y(new_new_n923_));
  INV        g901(.A(i_5_), .Y(new_new_n924_));
  NA3        g902(.A(new_new_n793_), .B(new_new_n104_), .C(new_new_n118_), .Y(new_new_n925_));
  INV        g903(.A(new_new_n925_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n926_), .B(new_new_n924_), .Y(new_new_n927_));
  NO4        g905(.A(new_new_n233_), .B(new_new_n202_), .C(i_0_), .D(i_12_), .Y(new_new_n928_));
  AOI220     g906(.A0(new_new_n928_), .A1(i_10_), .B0(new_new_n748_), .B1(new_new_n168_), .Y(new_new_n929_));
  BUFFER     g907(.A(new_new_n825_), .Y(new_new_n930_));
  NO3        g908(.A(new_new_n930_), .B(i_12_), .C(new_new_n125_), .Y(new_new_n931_));
  NA2        g909(.A(new_new_n931_), .B(new_new_n211_), .Y(new_new_n932_));
  NA2        g910(.A(new_new_n850_), .B(new_new_n451_), .Y(new_new_n933_));
  OAI220     g911(.A0(i_7_), .A1(new_new_n983_), .B0(new_new_n933_), .B1(new_new_n644_), .Y(new_new_n934_));
  NA2        g912(.A(new_new_n934_), .B(new_new_n839_), .Y(new_new_n935_));
  NA4        g913(.A(new_new_n935_), .B(new_new_n932_), .C(new_new_n929_), .D(new_new_n927_), .Y(new_new_n936_));
  NO4        g914(.A(new_new_n936_), .B(new_new_n923_), .C(new_new_n908_), .D(new_new_n895_), .Y(new_new_n937_));
  NA3        g915(.A(new_new_n845_), .B(new_new_n357_), .C(i_5_), .Y(new_new_n938_));
  NA2        g916(.A(new_new_n938_), .B(new_new_n586_), .Y(new_new_n939_));
  NA2        g917(.A(new_new_n939_), .B(new_new_n200_), .Y(new_new_n940_));
  AN2        g918(.A(new_new_n669_), .B(new_new_n358_), .Y(new_new_n941_));
  NA2        g919(.A(new_new_n178_), .B(new_new_n180_), .Y(new_new_n942_));
  AO210      g920(.A0(new_new_n941_), .A1(new_new_n33_), .B0(new_new_n942_), .Y(new_new_n943_));
  OAI210     g921(.A0(new_new_n590_), .A1(new_new_n588_), .B0(new_new_n308_), .Y(new_new_n944_));
  NA2        g922(.A(new_new_n944_), .B(new_new_n943_), .Y(new_new_n945_));
  NO2        g923(.A(new_new_n445_), .B(new_new_n260_), .Y(new_new_n946_));
  NO2        g924(.A(new_new_n946_), .B(new_new_n820_), .Y(new_new_n947_));
  INV        g925(.A(new_new_n947_), .Y(new_new_n948_));
  AOI210     g926(.A0(new_new_n945_), .A1(new_new_n48_), .B0(new_new_n948_), .Y(new_new_n949_));
  AOI210     g927(.A0(new_new_n949_), .A1(new_new_n940_), .B0(new_new_n68_), .Y(new_new_n950_));
  INV        g928(.A(new_new_n71_), .Y(new_new_n951_));
  INV        g929(.A(new_new_n851_), .Y(new_new_n952_));
  AOI210     g930(.A0(new_new_n952_), .A1(new_new_n951_), .B0(new_new_n647_), .Y(new_new_n953_));
  NA2        g931(.A(i_8_), .B(new_new_n71_), .Y(new_new_n954_));
  NO2        g932(.A(new_new_n954_), .B(new_new_n231_), .Y(new_new_n955_));
  NO2        g933(.A(new_new_n955_), .B(new_new_n953_), .Y(new_new_n956_));
  OAI210     g934(.A0(new_new_n262_), .A1(new_new_n152_), .B0(new_new_n82_), .Y(new_new_n957_));
  NA3        g935(.A(new_new_n724_), .B(new_new_n282_), .C(new_new_n75_), .Y(new_new_n958_));
  AOI210     g936(.A0(new_new_n958_), .A1(new_new_n957_), .B0(i_11_), .Y(new_new_n959_));
  NA2        g937(.A(new_new_n581_), .B(new_new_n208_), .Y(new_new_n960_));
  OAI210     g938(.A0(new_new_n960_), .A1(new_new_n845_), .B0(new_new_n200_), .Y(new_new_n961_));
  NA2        g939(.A(new_new_n158_), .B(i_5_), .Y(new_new_n962_));
  AOI210     g940(.A0(new_new_n961_), .A1(new_new_n731_), .B0(new_new_n962_), .Y(new_new_n963_));
  NO4        g941(.A(new_new_n872_), .B(new_new_n458_), .C(new_new_n246_), .D(new_new_n245_), .Y(new_new_n964_));
  NO2        g942(.A(new_new_n964_), .B(new_new_n538_), .Y(new_new_n965_));
  INV        g943(.A(new_new_n351_), .Y(new_new_n966_));
  AOI210     g944(.A0(new_new_n966_), .A1(new_new_n965_), .B0(new_new_n40_), .Y(new_new_n967_));
  NO3        g945(.A(new_new_n967_), .B(new_new_n963_), .C(new_new_n959_), .Y(new_new_n968_));
  OAI210     g946(.A0(new_new_n956_), .A1(i_4_), .B0(new_new_n968_), .Y(new_new_n969_));
  NO3        g947(.A(new_new_n969_), .B(new_new_n541_), .C(new_new_n950_), .Y(new_new_n970_));
  NA4        g948(.A(new_new_n970_), .B(new_new_n937_), .C(new_new_n879_), .D(new_new_n810_), .Y(men4));
  INV        g949(.A(i_2_), .Y(new_new_n974_));
  INV        g950(.A(new_new_n918_), .Y(new_new_n975_));
  INV        g951(.A(new_new_n320_), .Y(new_new_n976_));
  INV        g952(.A(i_6_), .Y(new_new_n977_));
  INV        g953(.A(i_10_), .Y(new_new_n978_));
  INV        g954(.A(i_11_), .Y(new_new_n979_));
  INV        g955(.A(i_3_), .Y(new_new_n980_));
  INV        g956(.A(i_9_), .Y(new_new_n981_));
  INV        g957(.A(i_6_), .Y(new_new_n982_));
  INV        g958(.A(i_5_), .Y(new_new_n983_));
  INV        g959(.A(i_12_), .Y(new_new_n984_));
  INV        g960(.A(new_new_n201_), .Y(new_new_n985_));
endmodule


