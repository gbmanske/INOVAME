// Benchmark "top" written by ABC on Thu Jun 20 14:00:11 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n127_,
    new_new_n128_, new_new_n129_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n637_, new_new_n638_,
    new_new_n639_, new_new_n640_, new_new_n641_, new_new_n642_,
    new_new_n643_, new_new_n644_, new_new_n645_, new_new_n646_,
    new_new_n647_, new_new_n648_, new_new_n649_, new_new_n650_,
    new_new_n651_, new_new_n652_, new_new_n653_, new_new_n654_,
    new_new_n655_, new_new_n656_, new_new_n657_, new_new_n658_,
    new_new_n659_, new_new_n660_, new_new_n661_, new_new_n662_,
    new_new_n663_, new_new_n664_, new_new_n665_, new_new_n666_,
    new_new_n667_, new_new_n668_, new_new_n669_, new_new_n670_,
    new_new_n671_, new_new_n672_, new_new_n673_, new_new_n675_,
    new_new_n676_, new_new_n677_, new_new_n678_, new_new_n679_,
    new_new_n680_, new_new_n681_, new_new_n682_, new_new_n683_,
    new_new_n684_, new_new_n685_, new_new_n686_, new_new_n687_,
    new_new_n688_, new_new_n689_, new_new_n690_, new_new_n691_,
    new_new_n692_, new_new_n693_, new_new_n694_, new_new_n695_,
    new_new_n696_, new_new_n697_, new_new_n698_, new_new_n699_,
    new_new_n700_, new_new_n701_, new_new_n702_, new_new_n703_,
    new_new_n704_, new_new_n705_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n709_, new_new_n710_, new_new_n711_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n874_, new_new_n875_,
    new_new_n876_, new_new_n877_, new_new_n878_, new_new_n879_,
    new_new_n880_, new_new_n881_, new_new_n882_, new_new_n883_,
    new_new_n884_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n55_));
  NA3        g033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  OAI210     g036(.A0(new_new_n58_), .A1(new_new_n57_), .B0(new_new_n56_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g039(.A(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_10_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NAi21      g042(.An(new_new_n64_), .B(new_new_n60_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n50_), .B(i_2_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_6_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(new_new_n25_), .Y(new_new_n68_));
  INV        g046(.A(i_0_), .Y(new_new_n69_));
  NAi21      g047(.An(i_5_), .B(i_10_), .Y(new_new_n70_));
  NA2        g048(.A(i_5_), .B(i_9_), .Y(new_new_n71_));
  AOI210     g049(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n69_), .Y(new_new_n72_));
  INV        g050(.A(new_new_n72_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n72_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n74_));
  NA2        g052(.A(i_12_), .B(i_5_), .Y(new_new_n75_));
  NA2        g053(.A(i_2_), .B(i_8_), .Y(new_new_n76_));
  NO2        g054(.A(i_3_), .B(i_9_), .Y(new_new_n77_));
  NO2        g055(.A(i_3_), .B(i_7_), .Y(new_new_n78_));
  NO3        g056(.A(new_new_n78_), .B(new_new_n77_), .C(new_new_n62_), .Y(new_new_n79_));
  INV        g057(.A(i_6_), .Y(new_new_n80_));
  OR4        g058(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n81_));
  INV        g059(.A(new_new_n81_), .Y(new_new_n82_));
  NO2        g060(.A(i_2_), .B(i_7_), .Y(new_new_n83_));
  NA2        g061(.A(new_new_n79_), .B(i_2_), .Y(new_new_n84_));
  NAi21      g062(.An(i_6_), .B(i_10_), .Y(new_new_n85_));
  NA2        g063(.A(i_2_), .B(i_6_), .Y(new_new_n86_));
  NO2        g064(.A(new_new_n84_), .B(new_new_n75_), .Y(new_new_n87_));
  AN3        g065(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_11_), .Y(new_new_n89_));
  NO2        g067(.A(i_5_), .B(i_8_), .Y(new_new_n90_));
  NOi21      g068(.An(new_new_n90_), .B(new_new_n89_), .Y(new_new_n91_));
  AOI220     g069(.A0(new_new_n91_), .A1(new_new_n61_), .B0(new_new_n88_), .B1(new_new_n32_), .Y(new_new_n92_));
  INV        g070(.A(i_7_), .Y(new_new_n93_));
  NO2        g071(.A(i_0_), .B(i_5_), .Y(new_new_n94_));
  NA2        g072(.A(i_12_), .B(i_3_), .Y(new_new_n95_));
  INV        g073(.A(new_new_n95_), .Y(new_new_n96_));
  NAi21      g074(.An(i_7_), .B(i_11_), .Y(new_new_n97_));
  NO3        g075(.A(new_new_n97_), .B(new_new_n85_), .C(new_new_n53_), .Y(new_new_n98_));
  AN2        g076(.A(i_2_), .B(i_10_), .Y(new_new_n99_));
  NO2        g077(.A(new_new_n99_), .B(i_7_), .Y(new_new_n100_));
  OR2        g078(.A(new_new_n75_), .B(new_new_n57_), .Y(new_new_n101_));
  NO2        g079(.A(i_8_), .B(new_new_n93_), .Y(new_new_n102_));
  NO3        g080(.A(new_new_n102_), .B(new_new_n101_), .C(new_new_n100_), .Y(new_new_n103_));
  NA2        g081(.A(i_12_), .B(i_7_), .Y(new_new_n104_));
  NO2        g082(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n105_));
  NA2        g083(.A(new_new_n105_), .B(i_0_), .Y(new_new_n106_));
  NA2        g084(.A(i_11_), .B(i_12_), .Y(new_new_n107_));
  OAI210     g085(.A0(new_new_n106_), .A1(new_new_n104_), .B0(new_new_n107_), .Y(new_new_n108_));
  NO2        g086(.A(new_new_n108_), .B(new_new_n103_), .Y(new_new_n109_));
  NAi31      g087(.An(new_new_n98_), .B(new_new_n109_), .C(new_new_n92_), .Y(new_new_n110_));
  NOi21      g088(.An(i_1_), .B(i_5_), .Y(new_new_n111_));
  NA2        g089(.A(new_new_n111_), .B(i_11_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n93_), .B(new_new_n37_), .Y(new_new_n113_));
  NA2        g091(.A(i_7_), .B(new_new_n25_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n114_), .B(new_new_n113_), .Y(new_new_n115_));
  NO2        g093(.A(new_new_n115_), .B(new_new_n46_), .Y(new_new_n116_));
  NAi21      g094(.An(i_3_), .B(i_8_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(new_new_n61_), .Y(new_new_n118_));
  BUFFER     g096(.A(new_new_n118_), .Y(new_new_n119_));
  NO2        g097(.A(i_1_), .B(new_new_n80_), .Y(new_new_n120_));
  NO2        g098(.A(i_6_), .B(i_5_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n121_), .B(i_3_), .Y(new_new_n122_));
  AO210      g100(.A0(new_new_n122_), .A1(new_new_n47_), .B0(new_new_n120_), .Y(new_new_n123_));
  OAI220     g101(.A0(new_new_n123_), .A1(new_new_n97_), .B0(new_new_n119_), .B1(new_new_n112_), .Y(new_new_n124_));
  NO3        g102(.A(new_new_n124_), .B(new_new_n110_), .C(new_new_n87_), .Y(new_new_n125_));
  NA3        g103(.A(new_new_n125_), .B(new_new_n74_), .C(new_new_n55_), .Y(mai2));
  NO2        g104(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n127_));
  NA2        g105(.A(i_6_), .B(new_new_n25_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(new_new_n127_), .Y(new_new_n129_));
  NA4        g107(.A(new_new_n129_), .B(new_new_n73_), .C(new_new_n66_), .D(new_new_n30_), .Y(mai0));
  AN2        g108(.A(i_8_), .B(i_7_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(i_6_), .Y(new_new_n132_));
  NO2        g110(.A(i_12_), .B(i_13_), .Y(new_new_n133_));
  NAi21      g111(.An(i_5_), .B(i_11_), .Y(new_new_n134_));
  NOi21      g112(.An(new_new_n133_), .B(new_new_n134_), .Y(new_new_n135_));
  NO2        g113(.A(i_0_), .B(i_1_), .Y(new_new_n136_));
  NA2        g114(.A(i_2_), .B(i_3_), .Y(new_new_n137_));
  NO2        g115(.A(new_new_n137_), .B(i_4_), .Y(new_new_n138_));
  NA3        g116(.A(new_new_n138_), .B(new_new_n136_), .C(new_new_n135_), .Y(new_new_n139_));
  NA2        g117(.A(i_1_), .B(i_5_), .Y(new_new_n140_));
  NO2        g118(.A(new_new_n69_), .B(new_new_n46_), .Y(new_new_n141_));
  NA2        g119(.A(new_new_n141_), .B(new_new_n36_), .Y(new_new_n142_));
  NO3        g120(.A(new_new_n142_), .B(new_new_n140_), .C(i_13_), .Y(new_new_n143_));
  OR2        g121(.A(i_0_), .B(i_1_), .Y(new_new_n144_));
  NO3        g122(.A(new_new_n144_), .B(new_new_n75_), .C(i_13_), .Y(new_new_n145_));
  NAi32      g123(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n146_));
  NAi21      g124(.An(new_new_n146_), .B(new_new_n145_), .Y(new_new_n147_));
  NOi21      g125(.An(i_4_), .B(i_10_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n40_), .Y(new_new_n149_));
  NO2        g127(.A(i_3_), .B(i_5_), .Y(new_new_n150_));
  NO3        g128(.A(new_new_n69_), .B(i_2_), .C(i_1_), .Y(new_new_n151_));
  NA2        g129(.A(new_new_n151_), .B(new_new_n150_), .Y(new_new_n152_));
  OAI210     g130(.A0(new_new_n152_), .A1(new_new_n149_), .B0(new_new_n147_), .Y(new_new_n153_));
  NO2        g131(.A(new_new_n153_), .B(new_new_n143_), .Y(new_new_n154_));
  NO2        g132(.A(new_new_n154_), .B(new_new_n132_), .Y(new_new_n155_));
  NA2        g133(.A(i_3_), .B(new_new_n48_), .Y(new_new_n156_));
  NOi21      g134(.An(i_4_), .B(i_9_), .Y(new_new_n157_));
  NOi21      g135(.An(i_11_), .B(i_13_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n157_), .Y(new_new_n159_));
  OR2        g137(.A(new_new_n159_), .B(new_new_n156_), .Y(new_new_n160_));
  NO2        g138(.A(i_4_), .B(i_5_), .Y(new_new_n161_));
  NAi21      g139(.An(i_12_), .B(i_11_), .Y(new_new_n162_));
  NA3        g140(.A(new_new_n883_), .B(new_new_n161_), .C(new_new_n77_), .Y(new_new_n163_));
  NA2        g141(.A(new_new_n163_), .B(new_new_n160_), .Y(new_new_n164_));
  NO2        g142(.A(new_new_n69_), .B(new_new_n62_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n46_), .Y(new_new_n166_));
  NA2        g144(.A(new_new_n36_), .B(i_5_), .Y(new_new_n167_));
  NAi31      g145(.An(new_new_n167_), .B(new_new_n77_), .C(i_11_), .Y(new_new_n168_));
  NA2        g146(.A(i_3_), .B(i_5_), .Y(new_new_n169_));
  AOI210     g147(.A0(new_new_n159_), .A1(new_new_n168_), .B0(new_new_n166_), .Y(new_new_n170_));
  NO2        g148(.A(new_new_n69_), .B(i_5_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n171_), .B(new_new_n44_), .Y(new_new_n172_));
  NO2        g150(.A(i_2_), .B(i_1_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(i_3_), .Y(new_new_n174_));
  NAi21      g152(.An(i_4_), .B(i_12_), .Y(new_new_n175_));
  NO3        g153(.A(new_new_n175_), .B(new_new_n174_), .C(new_new_n172_), .Y(new_new_n176_));
  NO3        g154(.A(new_new_n176_), .B(new_new_n170_), .C(new_new_n164_), .Y(new_new_n177_));
  INV        g155(.A(i_8_), .Y(new_new_n178_));
  NO2        g156(.A(new_new_n178_), .B(i_7_), .Y(new_new_n179_));
  NA2        g157(.A(new_new_n179_), .B(i_6_), .Y(new_new_n180_));
  NO3        g158(.A(i_3_), .B(new_new_n80_), .C(new_new_n48_), .Y(new_new_n181_));
  NA2        g159(.A(new_new_n181_), .B(new_new_n102_), .Y(new_new_n182_));
  NO3        g160(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n183_));
  NA3        g161(.A(new_new_n183_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n184_));
  NO2        g162(.A(i_11_), .B(new_new_n182_), .Y(new_new_n185_));
  NO2        g163(.A(i_3_), .B(i_8_), .Y(new_new_n186_));
  NO3        g164(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n187_));
  NA3        g165(.A(new_new_n187_), .B(new_new_n186_), .C(new_new_n40_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n94_), .B(new_new_n57_), .Y(new_new_n189_));
  NO2        g167(.A(i_13_), .B(i_9_), .Y(new_new_n190_));
  NA3        g168(.A(new_new_n190_), .B(i_6_), .C(new_new_n178_), .Y(new_new_n191_));
  BUFFER     g169(.A(new_new_n191_), .Y(new_new_n192_));
  NO2        g170(.A(new_new_n44_), .B(i_5_), .Y(new_new_n193_));
  NO3        g171(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n194_));
  NA3        g172(.A(new_new_n194_), .B(new_new_n193_), .C(i_10_), .Y(new_new_n195_));
  OAI220     g173(.A0(new_new_n195_), .A1(new_new_n192_), .B0(new_new_n57_), .B1(new_new_n188_), .Y(new_new_n196_));
  AOI210     g174(.A0(new_new_n196_), .A1(i_7_), .B0(new_new_n185_), .Y(new_new_n197_));
  OAI220     g175(.A0(new_new_n197_), .A1(i_4_), .B0(new_new_n180_), .B1(new_new_n177_), .Y(new_new_n198_));
  NA3        g176(.A(i_13_), .B(new_new_n178_), .C(i_10_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n199_), .B(i_12_), .Y(new_new_n200_));
  NA2        g178(.A(i_0_), .B(i_5_), .Y(new_new_n201_));
  OAI220     g179(.A0(new_new_n80_), .A1(new_new_n174_), .B0(new_new_n166_), .B1(new_new_n122_), .Y(new_new_n202_));
  NAi31      g180(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n203_));
  INV        g181(.A(i_13_), .Y(new_new_n204_));
  NO2        g182(.A(i_12_), .B(new_new_n204_), .Y(new_new_n205_));
  NA3        g183(.A(new_new_n205_), .B(new_new_n183_), .C(new_new_n181_), .Y(new_new_n206_));
  INV        g184(.A(new_new_n206_), .Y(new_new_n207_));
  AOI220     g185(.A0(new_new_n207_), .A1(new_new_n131_), .B0(new_new_n202_), .B1(new_new_n200_), .Y(new_new_n208_));
  NO2        g186(.A(i_12_), .B(new_new_n37_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n169_), .B(i_4_), .Y(new_new_n210_));
  NA2        g188(.A(new_new_n210_), .B(new_new_n209_), .Y(new_new_n211_));
  OR2        g189(.A(i_8_), .B(i_7_), .Y(new_new_n212_));
  NO2        g190(.A(new_new_n212_), .B(new_new_n80_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n53_), .B(i_1_), .Y(new_new_n214_));
  NA2        g192(.A(new_new_n214_), .B(new_new_n213_), .Y(new_new_n215_));
  INV        g193(.A(i_12_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n44_), .B(new_new_n216_), .Y(new_new_n217_));
  NO3        g195(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n218_));
  NA2        g196(.A(i_2_), .B(i_1_), .Y(new_new_n219_));
  NO2        g197(.A(new_new_n215_), .B(new_new_n211_), .Y(new_new_n220_));
  NO3        g198(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n221_));
  NAi21      g199(.An(i_4_), .B(i_3_), .Y(new_new_n222_));
  NO2        g200(.A(i_0_), .B(i_6_), .Y(new_new_n223_));
  NOi41      g201(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n219_), .B(new_new_n169_), .Y(new_new_n226_));
  NAi21      g204(.An(new_new_n225_), .B(new_new_n226_), .Y(new_new_n227_));
  INV        g205(.A(new_new_n227_), .Y(new_new_n228_));
  AOI210     g206(.A0(new_new_n228_), .A1(new_new_n40_), .B0(new_new_n220_), .Y(new_new_n229_));
  NO2        g207(.A(i_11_), .B(new_new_n204_), .Y(new_new_n230_));
  NOi21      g208(.An(i_1_), .B(i_6_), .Y(new_new_n231_));
  NAi21      g209(.An(i_3_), .B(i_7_), .Y(new_new_n232_));
  NA2        g210(.A(new_new_n216_), .B(i_9_), .Y(new_new_n233_));
  NA2        g211(.A(new_new_n69_), .B(i_5_), .Y(new_new_n234_));
  NA3        g212(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n235_));
  INV        g213(.A(new_new_n132_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n216_), .B(i_13_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n237_), .B(new_new_n71_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n238_), .B(new_new_n236_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n212_), .B(new_new_n37_), .Y(new_new_n240_));
  NA2        g218(.A(i_12_), .B(i_6_), .Y(new_new_n241_));
  OR2        g219(.A(i_13_), .B(i_9_), .Y(new_new_n242_));
  NO3        g220(.A(new_new_n242_), .B(new_new_n241_), .C(new_new_n48_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n222_), .B(i_2_), .Y(new_new_n244_));
  NA3        g222(.A(new_new_n244_), .B(new_new_n243_), .C(new_new_n44_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n230_), .B(i_9_), .Y(new_new_n246_));
  OAI210     g224(.A0(new_new_n62_), .A1(new_new_n246_), .B0(new_new_n245_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n141_), .B(new_new_n62_), .Y(new_new_n248_));
  NO3        g226(.A(i_11_), .B(new_new_n204_), .C(new_new_n25_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n232_), .B(i_8_), .Y(new_new_n250_));
  NO2        g228(.A(i_6_), .B(new_new_n48_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n250_), .B(new_new_n249_), .Y(new_new_n252_));
  NA3        g230(.A(i_6_), .B(new_new_n240_), .C(new_new_n205_), .Y(new_new_n253_));
  AOI210     g231(.A0(new_new_n253_), .A1(new_new_n252_), .B0(new_new_n248_), .Y(new_new_n254_));
  AOI210     g232(.A0(new_new_n247_), .A1(new_new_n240_), .B0(new_new_n254_), .Y(new_new_n255_));
  NA4        g233(.A(new_new_n255_), .B(new_new_n239_), .C(new_new_n229_), .D(new_new_n208_), .Y(new_new_n256_));
  NO3        g234(.A(i_12_), .B(new_new_n204_), .C(new_new_n37_), .Y(new_new_n257_));
  INV        g235(.A(new_new_n257_), .Y(new_new_n258_));
  NO3        g236(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n259_));
  NO3        g237(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n219_), .B(i_0_), .Y(new_new_n261_));
  AOI220     g239(.A0(new_new_n261_), .A1(new_new_n179_), .B0(new_new_n260_), .B1(new_new_n131_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n251_), .B(new_new_n26_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n263_), .B(new_new_n262_), .Y(new_new_n264_));
  NA2        g242(.A(i_0_), .B(i_1_), .Y(new_new_n265_));
  NO2        g243(.A(new_new_n265_), .B(i_2_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n58_), .B(i_6_), .Y(new_new_n267_));
  NA3        g245(.A(new_new_n267_), .B(new_new_n266_), .C(new_new_n150_), .Y(new_new_n268_));
  OAI210     g246(.A0(new_new_n152_), .A1(new_new_n132_), .B0(new_new_n268_), .Y(new_new_n269_));
  NO2        g247(.A(new_new_n269_), .B(new_new_n264_), .Y(new_new_n270_));
  NO2        g248(.A(i_3_), .B(i_10_), .Y(new_new_n271_));
  NA3        g249(.A(new_new_n271_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n272_));
  NO2        g250(.A(i_2_), .B(new_new_n93_), .Y(new_new_n273_));
  NA2        g251(.A(i_1_), .B(new_new_n36_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n274_), .B(i_8_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n275_), .B(new_new_n273_), .Y(new_new_n276_));
  AN2        g254(.A(i_3_), .B(i_10_), .Y(new_new_n277_));
  NA3        g255(.A(new_new_n183_), .B(new_new_n883_), .C(new_new_n161_), .Y(new_new_n278_));
  NO2        g256(.A(i_5_), .B(new_new_n37_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n280_));
  OR2        g258(.A(new_new_n276_), .B(new_new_n272_), .Y(new_new_n281_));
  OAI220     g259(.A0(new_new_n281_), .A1(i_6_), .B0(new_new_n270_), .B1(new_new_n258_), .Y(new_new_n282_));
  NO4        g260(.A(new_new_n282_), .B(new_new_n256_), .C(new_new_n198_), .D(new_new_n155_), .Y(new_new_n283_));
  NO3        g261(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n284_));
  NO3        g262(.A(i_6_), .B(new_new_n178_), .C(i_7_), .Y(new_new_n285_));
  AOI210     g263(.A0(i_1_), .A1(new_new_n219_), .B0(new_new_n156_), .Y(new_new_n286_));
  NO2        g264(.A(i_2_), .B(i_3_), .Y(new_new_n287_));
  OR2        g265(.A(i_0_), .B(i_5_), .Y(new_new_n288_));
  NA2        g266(.A(new_new_n201_), .B(new_new_n288_), .Y(new_new_n289_));
  NA4        g267(.A(new_new_n289_), .B(new_new_n213_), .C(new_new_n287_), .D(i_1_), .Y(new_new_n290_));
  NA3        g268(.A(new_new_n261_), .B(new_new_n150_), .C(new_new_n102_), .Y(new_new_n291_));
  NAi21      g269(.An(i_8_), .B(i_7_), .Y(new_new_n292_));
  NO2        g270(.A(new_new_n292_), .B(i_6_), .Y(new_new_n293_));
  NA3        g271(.A(i_2_), .B(new_new_n293_), .C(new_new_n150_), .Y(new_new_n294_));
  NA3        g272(.A(new_new_n294_), .B(new_new_n291_), .C(new_new_n290_), .Y(new_new_n295_));
  OAI210     g273(.A0(new_new_n295_), .A1(new_new_n286_), .B0(i_4_), .Y(new_new_n296_));
  NO2        g274(.A(i_12_), .B(i_10_), .Y(new_new_n297_));
  NOi21      g275(.An(i_5_), .B(i_0_), .Y(new_new_n298_));
  NO3        g276(.A(new_new_n274_), .B(new_new_n298_), .C(new_new_n117_), .Y(new_new_n299_));
  NA4        g277(.A(new_new_n78_), .B(new_new_n36_), .C(new_new_n80_), .D(i_8_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n299_), .B(new_new_n297_), .Y(new_new_n301_));
  NO2        g279(.A(i_6_), .B(i_8_), .Y(new_new_n302_));
  NOi21      g280(.An(i_0_), .B(i_2_), .Y(new_new_n303_));
  AN2        g281(.A(new_new_n303_), .B(new_new_n302_), .Y(new_new_n304_));
  NO2        g282(.A(i_1_), .B(i_7_), .Y(new_new_n305_));
  AO220      g283(.A0(new_new_n305_), .A1(new_new_n304_), .B0(new_new_n293_), .B1(new_new_n214_), .Y(new_new_n306_));
  NA2        g284(.A(new_new_n306_), .B(i_4_), .Y(new_new_n307_));
  NA3        g285(.A(new_new_n307_), .B(new_new_n301_), .C(new_new_n296_), .Y(new_new_n308_));
  NO3        g286(.A(new_new_n212_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n309_));
  NO3        g287(.A(new_new_n292_), .B(i_2_), .C(i_1_), .Y(new_new_n310_));
  OAI210     g288(.A0(new_new_n310_), .A1(new_new_n309_), .B0(i_6_), .Y(new_new_n311_));
  NA2        g289(.A(new_new_n231_), .B(new_new_n273_), .Y(new_new_n312_));
  AOI210     g290(.A0(new_new_n312_), .A1(new_new_n311_), .B0(new_new_n289_), .Y(new_new_n313_));
  NA2        g291(.A(new_new_n313_), .B(i_3_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n86_), .B(new_new_n178_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n315_), .B(new_new_n62_), .Y(new_new_n316_));
  NO2        g294(.A(new_new_n316_), .B(i_7_), .Y(new_new_n317_));
  NO2        g295(.A(new_new_n178_), .B(i_9_), .Y(new_new_n318_));
  NA2        g296(.A(new_new_n318_), .B(new_new_n189_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n317_), .B(new_new_n264_), .Y(new_new_n320_));
  AOI210     g298(.A0(new_new_n320_), .A1(new_new_n314_), .B0(new_new_n149_), .Y(new_new_n321_));
  AOI210     g299(.A0(new_new_n308_), .A1(new_new_n284_), .B0(new_new_n321_), .Y(new_new_n322_));
  NOi32      g300(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n323_));
  INV        g301(.A(new_new_n323_), .Y(new_new_n324_));
  NAi21      g302(.An(i_0_), .B(i_6_), .Y(new_new_n325_));
  NAi21      g303(.An(i_1_), .B(i_5_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n326_), .B(new_new_n325_), .Y(new_new_n327_));
  NA2        g305(.A(new_new_n327_), .B(new_new_n25_), .Y(new_new_n328_));
  OAI210     g306(.A0(new_new_n328_), .A1(new_new_n146_), .B0(new_new_n225_), .Y(new_new_n329_));
  NAi41      g307(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n330_));
  OAI220     g308(.A0(new_new_n330_), .A1(new_new_n326_), .B0(new_new_n203_), .B1(new_new_n146_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n146_), .B(new_new_n144_), .Y(new_new_n332_));
  OR2        g310(.A(new_new_n332_), .B(new_new_n331_), .Y(new_new_n333_));
  NO2        g311(.A(i_1_), .B(new_new_n93_), .Y(new_new_n334_));
  NAi21      g312(.An(i_3_), .B(i_4_), .Y(new_new_n335_));
  NA2        g313(.A(i_2_), .B(i_7_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n335_), .B(i_10_), .Y(new_new_n337_));
  AOI210     g315(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n338_));
  OAI210     g316(.A0(new_new_n338_), .A1(new_new_n173_), .B0(new_new_n337_), .Y(new_new_n339_));
  AOI220     g317(.A0(new_new_n337_), .A1(new_new_n305_), .B0(new_new_n218_), .B1(new_new_n173_), .Y(new_new_n340_));
  AOI210     g318(.A0(new_new_n340_), .A1(new_new_n339_), .B0(i_5_), .Y(new_new_n341_));
  NO3        g319(.A(new_new_n341_), .B(new_new_n333_), .C(new_new_n329_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n342_), .B(new_new_n324_), .Y(new_new_n343_));
  NO2        g321(.A(new_new_n58_), .B(new_new_n25_), .Y(new_new_n344_));
  AN2        g322(.A(i_12_), .B(i_5_), .Y(new_new_n345_));
  NO2        g323(.A(i_4_), .B(new_new_n26_), .Y(new_new_n346_));
  NA2        g324(.A(new_new_n346_), .B(new_new_n345_), .Y(new_new_n347_));
  NO2        g325(.A(i_11_), .B(i_6_), .Y(new_new_n348_));
  NA3        g326(.A(new_new_n348_), .B(i_2_), .C(new_new_n204_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(new_new_n347_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n222_), .B(i_5_), .Y(new_new_n351_));
  NO2        g329(.A(i_5_), .B(i_10_), .Y(new_new_n352_));
  AOI220     g330(.A0(new_new_n352_), .A1(new_new_n244_), .B0(new_new_n351_), .B1(new_new_n183_), .Y(new_new_n353_));
  NA2        g331(.A(new_new_n133_), .B(new_new_n45_), .Y(new_new_n354_));
  NO2        g332(.A(new_new_n354_), .B(new_new_n353_), .Y(new_new_n355_));
  OAI210     g333(.A0(new_new_n355_), .A1(new_new_n350_), .B0(new_new_n344_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n139_), .B(new_new_n80_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n358_), .B(new_new_n350_), .Y(new_new_n359_));
  NO2        g337(.A(i_11_), .B(i_12_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n352_), .B(new_new_n216_), .Y(new_new_n361_));
  NAi21      g339(.An(i_13_), .B(i_0_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n362_), .B(new_new_n219_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n877_), .B(new_new_n363_), .Y(new_new_n364_));
  NA3        g342(.A(new_new_n364_), .B(new_new_n359_), .C(new_new_n356_), .Y(new_new_n365_));
  NA2        g343(.A(new_new_n44_), .B(new_new_n204_), .Y(new_new_n366_));
  NO2        g344(.A(i_0_), .B(i_11_), .Y(new_new_n367_));
  AN2        g345(.A(i_1_), .B(i_6_), .Y(new_new_n368_));
  NOi21      g346(.An(i_2_), .B(i_12_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n369_), .B(new_new_n368_), .Y(new_new_n370_));
  INV        g348(.A(new_new_n370_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n881_), .B(i_4_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n371_), .B(new_new_n372_), .Y(new_new_n373_));
  OR2        g351(.A(i_13_), .B(i_10_), .Y(new_new_n374_));
  NO3        g352(.A(new_new_n374_), .B(new_new_n107_), .C(i_9_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n159_), .B(new_new_n113_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n93_), .B(new_new_n25_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n251_), .B(new_new_n194_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n378_), .B(new_new_n199_), .Y(new_new_n379_));
  INV        g357(.A(new_new_n379_), .Y(new_new_n380_));
  AOI210     g358(.A0(new_new_n380_), .A1(new_new_n373_), .B0(new_new_n26_), .Y(new_new_n381_));
  NA2        g359(.A(new_new_n291_), .B(new_new_n290_), .Y(new_new_n382_));
  AOI220     g360(.A0(new_new_n267_), .A1(new_new_n259_), .B0(new_new_n261_), .B1(i_6_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n156_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n169_), .B(new_new_n80_), .Y(new_new_n385_));
  AOI220     g363(.A0(new_new_n385_), .A1(new_new_n266_), .B0(i_6_), .B1(new_new_n194_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n386_), .B(i_7_), .Y(new_new_n387_));
  NO3        g365(.A(new_new_n387_), .B(new_new_n384_), .C(new_new_n382_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n181_), .B(new_new_n88_), .Y(new_new_n389_));
  NA3        g367(.A(i_2_), .B(new_new_n150_), .C(new_new_n80_), .Y(new_new_n390_));
  AOI210     g368(.A0(new_new_n390_), .A1(new_new_n389_), .B0(new_new_n292_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n267_), .B(new_new_n214_), .Y(new_new_n392_));
  NO2        g370(.A(new_new_n392_), .B(new_new_n169_), .Y(new_new_n393_));
  NA3        g371(.A(new_new_n305_), .B(new_new_n304_), .C(i_5_), .Y(new_new_n394_));
  INV        g372(.A(new_new_n285_), .Y(new_new_n395_));
  OAI210     g373(.A0(new_new_n395_), .A1(new_new_n174_), .B0(new_new_n394_), .Y(new_new_n396_));
  NO3        g374(.A(new_new_n396_), .B(new_new_n393_), .C(new_new_n391_), .Y(new_new_n397_));
  AOI210     g375(.A0(new_new_n397_), .A1(new_new_n388_), .B0(new_new_n246_), .Y(new_new_n398_));
  NO4        g376(.A(new_new_n398_), .B(new_new_n381_), .C(new_new_n365_), .D(new_new_n343_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n69_), .B(i_13_), .Y(new_new_n400_));
  NA3        g378(.A(new_new_n400_), .B(i_1_), .C(i_2_), .Y(new_new_n401_));
  NO2        g379(.A(i_10_), .B(i_9_), .Y(new_new_n402_));
  NAi21      g380(.An(i_12_), .B(i_8_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n403_), .B(i_3_), .Y(new_new_n404_));
  NA2        g382(.A(i_2_), .B(i_6_), .Y(new_new_n405_));
  OAI220     g383(.A0(new_new_n405_), .A1(new_new_n188_), .B0(new_new_n880_), .B1(new_new_n401_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n280_), .B(i_0_), .Y(new_new_n407_));
  NO3        g385(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n241_), .B(new_new_n89_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n409_), .B(new_new_n408_), .Y(new_new_n410_));
  NA2        g388(.A(i_8_), .B(i_9_), .Y(new_new_n411_));
  NO2        g389(.A(i_7_), .B(i_2_), .Y(new_new_n412_));
  OR2        g390(.A(new_new_n412_), .B(new_new_n411_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n257_), .B(new_new_n189_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n414_), .B(new_new_n413_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n230_), .B(new_new_n279_), .Y(new_new_n416_));
  NO3        g394(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n417_));
  INV        g395(.A(new_new_n417_), .Y(new_new_n418_));
  NA3        g396(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n419_));
  NA3        g397(.A(new_new_n134_), .B(new_new_n105_), .C(new_new_n23_), .Y(new_new_n420_));
  OAI220     g398(.A0(new_new_n420_), .A1(new_new_n419_), .B0(new_new_n418_), .B1(new_new_n416_), .Y(new_new_n421_));
  NO3        g399(.A(new_new_n421_), .B(new_new_n415_), .C(new_new_n406_), .Y(new_new_n422_));
  OR2        g400(.A(new_new_n265_), .B(new_new_n191_), .Y(new_new_n423_));
  OA210      g401(.A0(new_new_n319_), .A1(new_new_n93_), .B0(new_new_n268_), .Y(new_new_n424_));
  OA220      g402(.A0(new_new_n424_), .A1(new_new_n149_), .B0(new_new_n423_), .B1(new_new_n211_), .Y(new_new_n425_));
  NA2        g403(.A(new_new_n88_), .B(i_13_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n385_), .B(new_new_n344_), .Y(new_new_n427_));
  NO2        g405(.A(i_2_), .B(i_13_), .Y(new_new_n428_));
  NO2        g406(.A(new_new_n427_), .B(new_new_n426_), .Y(new_new_n429_));
  NO3        g407(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n430_));
  NO2        g408(.A(i_6_), .B(i_7_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n431_), .B(new_new_n430_), .Y(new_new_n432_));
  NO2        g410(.A(i_11_), .B(i_1_), .Y(new_new_n433_));
  NOi21      g411(.An(i_2_), .B(i_7_), .Y(new_new_n434_));
  NAi31      g412(.An(i_11_), .B(new_new_n434_), .C(i_0_), .Y(new_new_n435_));
  NO2        g413(.A(new_new_n374_), .B(i_6_), .Y(new_new_n436_));
  NA3        g414(.A(new_new_n436_), .B(i_1_), .C(new_new_n71_), .Y(new_new_n437_));
  NO2        g415(.A(new_new_n437_), .B(new_new_n435_), .Y(new_new_n438_));
  NO2        g416(.A(i_3_), .B(new_new_n178_), .Y(new_new_n439_));
  NO2        g417(.A(i_6_), .B(i_10_), .Y(new_new_n440_));
  NA3        g418(.A(new_new_n440_), .B(new_new_n284_), .C(new_new_n439_), .Y(new_new_n441_));
  NO2        g419(.A(new_new_n441_), .B(new_new_n142_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n443_));
  NO2        g421(.A(new_new_n144_), .B(i_3_), .Y(new_new_n444_));
  NAi31      g422(.An(new_new_n443_), .B(new_new_n444_), .C(new_new_n205_), .Y(new_new_n445_));
  NA3        g423(.A(new_new_n357_), .B(new_new_n165_), .C(new_new_n138_), .Y(new_new_n446_));
  NA2        g424(.A(new_new_n446_), .B(new_new_n445_), .Y(new_new_n447_));
  NO4        g425(.A(new_new_n447_), .B(new_new_n442_), .C(new_new_n438_), .D(new_new_n429_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n408_), .B(new_new_n345_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n417_), .B(new_new_n352_), .Y(new_new_n450_));
  NAi21      g428(.An(new_new_n199_), .B(new_new_n360_), .Y(new_new_n451_));
  INV        g429(.A(new_new_n305_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n26_), .B(i_5_), .Y(new_new_n453_));
  NA3        g431(.A(i_6_), .B(new_new_n453_), .C(new_new_n131_), .Y(new_new_n454_));
  OR3        g432(.A(new_new_n274_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n455_));
  OAI220     g433(.A0(new_new_n455_), .A1(new_new_n454_), .B0(new_new_n452_), .B1(new_new_n451_), .Y(new_new_n456_));
  NA3        g434(.A(new_new_n277_), .B(i_1_), .C(new_new_n69_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n457_), .B(new_new_n432_), .Y(new_new_n458_));
  NO2        g436(.A(new_new_n458_), .B(new_new_n456_), .Y(new_new_n459_));
  NA4        g437(.A(new_new_n459_), .B(new_new_n448_), .C(new_new_n425_), .D(new_new_n422_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n112_), .B(new_new_n101_), .Y(new_new_n461_));
  AN2        g439(.A(new_new_n461_), .B(new_new_n408_), .Y(new_new_n462_));
  INV        g440(.A(new_new_n151_), .Y(new_new_n463_));
  OAI210     g441(.A0(new_new_n463_), .A1(new_new_n211_), .B0(new_new_n278_), .Y(new_new_n464_));
  AOI220     g442(.A0(new_new_n464_), .A1(new_new_n293_), .B0(new_new_n462_), .B1(new_new_n280_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n323_), .B(new_new_n69_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n36_), .B(i_8_), .Y(new_new_n467_));
  NAi41      g445(.An(new_new_n466_), .B(new_new_n440_), .C(new_new_n467_), .D(new_new_n46_), .Y(new_new_n468_));
  AOI210     g446(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n375_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n469_), .B(new_new_n468_), .Y(new_new_n470_));
  INV        g448(.A(new_new_n470_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n234_), .B(i_1_), .Y(new_new_n472_));
  OAI210     g450(.A0(i_8_), .A1(new_new_n472_), .B0(new_new_n123_), .Y(new_new_n473_));
  INV        g451(.A(new_new_n184_), .Y(new_new_n474_));
  OR2        g452(.A(new_new_n169_), .B(i_4_), .Y(new_new_n475_));
  INV        g453(.A(new_new_n475_), .Y(new_new_n476_));
  AOI220     g454(.A0(new_new_n476_), .A1(new_new_n474_), .B0(new_new_n473_), .B1(new_new_n376_), .Y(new_new_n477_));
  NA3        g455(.A(new_new_n477_), .B(new_new_n471_), .C(new_new_n465_), .Y(new_new_n478_));
  NA2        g456(.A(new_new_n351_), .B(new_new_n266_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n347_), .B(new_new_n479_), .Y(new_new_n480_));
  NO2        g458(.A(new_new_n374_), .B(new_new_n38_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n481_), .B(new_new_n480_), .Y(new_new_n482_));
  NO2        g460(.A(i_8_), .B(i_7_), .Y(new_new_n483_));
  OAI220     g461(.A0(new_new_n46_), .A1(new_new_n475_), .B0(i_5_), .B1(new_new_n222_), .Y(new_new_n484_));
  NO2        g462(.A(i_11_), .B(i_6_), .Y(new_new_n485_));
  NA3        g463(.A(new_new_n485_), .B(new_new_n484_), .C(new_new_n483_), .Y(new_new_n486_));
  AOI220     g464(.A0(new_new_n385_), .A1(i_2_), .B0(new_new_n226_), .B1(new_new_n223_), .Y(new_new_n487_));
  OAI220     g465(.A0(new_new_n487_), .A1(new_new_n237_), .B0(new_new_n426_), .B1(new_new_n122_), .Y(new_new_n488_));
  NA2        g466(.A(new_new_n488_), .B(new_new_n240_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n272_), .B(new_new_n167_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n161_), .B(new_new_n88_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n144_), .B(i_5_), .Y(new_new_n492_));
  NA3        g470(.A(new_new_n492_), .B(new_new_n366_), .C(new_new_n287_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n493_), .B(new_new_n491_), .Y(new_new_n494_));
  OAI210     g472(.A0(new_new_n494_), .A1(new_new_n490_), .B0(new_new_n417_), .Y(new_new_n495_));
  NA4        g473(.A(new_new_n495_), .B(new_new_n489_), .C(new_new_n486_), .D(new_new_n482_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n257_), .B(new_new_n78_), .Y(new_new_n497_));
  NO2        g475(.A(new_new_n76_), .B(new_new_n497_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n46_), .B(new_new_n160_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n499_), .B(new_new_n498_), .Y(new_new_n500_));
  NO4        g478(.A(new_new_n231_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n501_));
  NO3        g479(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n212_), .B(new_new_n36_), .Y(new_new_n503_));
  AN2        g481(.A(new_new_n503_), .B(new_new_n502_), .Y(new_new_n504_));
  OA210      g482(.A0(new_new_n504_), .A1(new_new_n501_), .B0(new_new_n323_), .Y(new_new_n505_));
  NO2        g483(.A(new_new_n374_), .B(i_1_), .Y(new_new_n506_));
  NOi31      g484(.An(new_new_n506_), .B(new_new_n409_), .C(new_new_n69_), .Y(new_new_n507_));
  AN4        g485(.A(new_new_n507_), .B(new_new_n372_), .C(new_new_n453_), .D(i_2_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n383_), .B(new_new_n163_), .Y(new_new_n509_));
  NO3        g487(.A(new_new_n509_), .B(new_new_n508_), .C(new_new_n505_), .Y(new_new_n510_));
  NOi21      g488(.An(i_10_), .B(i_6_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n249_), .B(new_new_n511_), .Y(new_new_n512_));
  NO2        g490(.A(new_new_n512_), .B(new_new_n407_), .Y(new_new_n513_));
  NO2        g491(.A(new_new_n104_), .B(new_new_n23_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n285_), .B(new_new_n151_), .Y(new_new_n515_));
  AOI220     g493(.A0(new_new_n515_), .A1(new_new_n392_), .B0(new_new_n159_), .B1(new_new_n168_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n183_), .B(new_new_n37_), .Y(new_new_n517_));
  NOi31      g495(.An(new_new_n135_), .B(new_new_n517_), .C(new_new_n300_), .Y(new_new_n518_));
  NO3        g496(.A(new_new_n518_), .B(new_new_n516_), .C(new_new_n513_), .Y(new_new_n519_));
  NO2        g497(.A(new_new_n466_), .B(new_new_n340_), .Y(new_new_n520_));
  INV        g498(.A(new_new_n287_), .Y(new_new_n521_));
  NO2        g499(.A(i_12_), .B(new_new_n80_), .Y(new_new_n522_));
  NA3        g500(.A(new_new_n522_), .B(new_new_n249_), .C(i_5_), .Y(new_new_n523_));
  NA3        g501(.A(new_new_n348_), .B(new_new_n257_), .C(new_new_n201_), .Y(new_new_n524_));
  AOI210     g502(.A0(new_new_n524_), .A1(new_new_n523_), .B0(new_new_n521_), .Y(new_new_n525_));
  NO3        g503(.A(i_4_), .B(new_new_n311_), .C(new_new_n272_), .Y(new_new_n526_));
  NO3        g504(.A(new_new_n526_), .B(new_new_n525_), .C(new_new_n520_), .Y(new_new_n527_));
  NA4        g505(.A(new_new_n527_), .B(new_new_n519_), .C(new_new_n510_), .D(new_new_n500_), .Y(new_new_n528_));
  NO4        g506(.A(new_new_n528_), .B(new_new_n496_), .C(new_new_n478_), .D(new_new_n460_), .Y(new_new_n529_));
  NA4        g507(.A(new_new_n529_), .B(new_new_n399_), .C(new_new_n322_), .D(new_new_n283_), .Y(mai7));
  NO2        g508(.A(new_new_n86_), .B(new_new_n54_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n97_), .B(new_new_n85_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n440_), .B(new_new_n78_), .Y(new_new_n533_));
  NA2        g511(.A(i_11_), .B(new_new_n178_), .Y(new_new_n534_));
  NA3        g512(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n216_), .B(i_4_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n95_), .B(new_new_n535_), .Y(new_new_n537_));
  NA2        g515(.A(i_2_), .B(new_new_n80_), .Y(new_new_n538_));
  NO2        g516(.A(i_7_), .B(new_new_n37_), .Y(new_new_n539_));
  NA2        g517(.A(i_4_), .B(i_8_), .Y(new_new_n540_));
  NO4        g518(.A(new_new_n187_), .B(new_new_n537_), .C(new_new_n532_), .D(new_new_n531_), .Y(new_new_n541_));
  AOI210     g519(.A0(new_new_n117_), .A1(new_new_n61_), .B0(i_10_), .Y(new_new_n542_));
  AOI210     g520(.A0(new_new_n542_), .A1(new_new_n216_), .B0(new_new_n148_), .Y(new_new_n543_));
  OR2        g521(.A(i_6_), .B(i_10_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n544_), .B(new_new_n23_), .Y(new_new_n545_));
  NO3        g523(.A(i_10_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n546_), .B(new_new_n545_), .Y(new_new_n547_));
  OA220      g525(.A0(new_new_n547_), .A1(new_new_n521_), .B0(new_new_n543_), .B1(new_new_n242_), .Y(new_new_n548_));
  AOI210     g526(.A0(new_new_n548_), .A1(new_new_n541_), .B0(new_new_n62_), .Y(new_new_n549_));
  NOi21      g527(.An(i_11_), .B(i_7_), .Y(new_new_n550_));
  NO2        g528(.A(i_2_), .B(new_new_n550_), .Y(new_new_n551_));
  NA3        g529(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n552_));
  NAi21      g530(.An(new_new_n552_), .B(i_11_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n553_), .B(new_new_n62_), .Y(new_new_n554_));
  NA2        g532(.A(new_new_n82_), .B(new_new_n62_), .Y(new_new_n555_));
  AO210      g533(.A0(new_new_n555_), .A1(new_new_n340_), .B0(new_new_n41_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n205_), .B(new_new_n62_), .Y(new_new_n557_));
  NO2        g535(.A(new_new_n62_), .B(i_9_), .Y(new_new_n558_));
  NO2        g536(.A(i_1_), .B(i_12_), .Y(new_new_n559_));
  NA2        g537(.A(new_new_n557_), .B(new_new_n556_), .Y(new_new_n560_));
  OAI210     g538(.A0(new_new_n560_), .A1(new_new_n554_), .B0(i_6_), .Y(new_new_n561_));
  NO2        g539(.A(i_6_), .B(i_11_), .Y(new_new_n562_));
  INV        g540(.A(new_new_n410_), .Y(new_new_n563_));
  NO4        g541(.A(i_12_), .B(new_new_n117_), .C(i_13_), .D(new_new_n80_), .Y(new_new_n564_));
  NA2        g542(.A(new_new_n564_), .B(new_new_n558_), .Y(new_new_n565_));
  INV        g543(.A(new_new_n565_), .Y(new_new_n566_));
  NA3        g544(.A(new_new_n483_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n127_), .B(i_9_), .Y(new_new_n568_));
  NA3        g546(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n569_));
  NO2        g547(.A(new_new_n568_), .B(new_new_n875_), .Y(new_new_n570_));
  NA3        g548(.A(new_new_n558_), .B(new_new_n287_), .C(i_6_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n571_), .B(new_new_n23_), .Y(new_new_n572_));
  AOI210     g550(.A0(new_new_n433_), .A1(new_new_n377_), .B0(new_new_n221_), .Y(new_new_n573_));
  NO2        g551(.A(new_new_n573_), .B(new_new_n538_), .Y(new_new_n574_));
  NO2        g552(.A(i_11_), .B(new_new_n37_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n575_), .B(new_new_n24_), .Y(new_new_n576_));
  NO2        g554(.A(new_new_n576_), .B(i_6_), .Y(new_new_n577_));
  OR4        g555(.A(new_new_n577_), .B(new_new_n574_), .C(new_new_n572_), .D(new_new_n570_), .Y(new_new_n578_));
  NO3        g556(.A(new_new_n578_), .B(new_new_n566_), .C(new_new_n563_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n212_), .B(new_new_n44_), .Y(new_new_n580_));
  NO3        g558(.A(new_new_n580_), .B(new_new_n280_), .C(new_new_n217_), .Y(new_new_n581_));
  NO2        g559(.A(i_10_), .B(i_6_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n80_), .B(i_9_), .Y(new_new_n583_));
  NO2        g561(.A(new_new_n583_), .B(new_new_n62_), .Y(new_new_n584_));
  NO2        g562(.A(new_new_n584_), .B(new_new_n559_), .Y(new_new_n585_));
  NO4        g563(.A(new_new_n585_), .B(new_new_n582_), .C(new_new_n581_), .D(i_4_), .Y(new_new_n586_));
  NA2        g564(.A(i_1_), .B(i_3_), .Y(new_new_n587_));
  INV        g565(.A(new_new_n586_), .Y(new_new_n588_));
  NA3        g566(.A(new_new_n588_), .B(new_new_n579_), .C(new_new_n561_), .Y(new_new_n589_));
  NO3        g567(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n590_));
  NOi21      g568(.An(new_new_n590_), .B(i_10_), .Y(new_new_n591_));
  OA210      g569(.A0(new_new_n591_), .A1(new_new_n224_), .B0(new_new_n80_), .Y(new_new_n592_));
  NA3        g570(.A(new_new_n440_), .B(new_new_n467_), .C(new_new_n46_), .Y(new_new_n593_));
  NO3        g571(.A(new_new_n434_), .B(new_new_n540_), .C(new_new_n80_), .Y(new_new_n594_));
  NA2        g572(.A(new_new_n594_), .B(new_new_n25_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n595_), .B(new_new_n593_), .Y(new_new_n596_));
  OAI210     g574(.A0(new_new_n596_), .A1(new_new_n592_), .B0(i_1_), .Y(new_new_n597_));
  AOI210     g575(.A0(new_new_n241_), .A1(new_new_n89_), .B0(i_1_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n335_), .B(i_2_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n599_), .B(new_new_n598_), .Y(new_new_n600_));
  AOI210     g578(.A0(new_new_n600_), .A1(new_new_n597_), .B0(i_13_), .Y(new_new_n601_));
  NA2        g579(.A(new_new_n96_), .B(new_new_n127_), .Y(new_new_n602_));
  AOI220     g580(.A0(new_new_n428_), .A1(new_new_n148_), .B0(i_2_), .B1(new_new_n127_), .Y(new_new_n603_));
  OAI210     g581(.A0(new_new_n603_), .A1(new_new_n44_), .B0(new_new_n602_), .Y(new_new_n604_));
  NO2        g582(.A(new_new_n54_), .B(i_12_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n224_), .B(new_new_n120_), .Y(new_new_n606_));
  OAI220     g584(.A0(new_new_n606_), .A1(new_new_n41_), .B0(new_new_n874_), .B1(new_new_n86_), .Y(new_new_n607_));
  AOI210     g585(.A0(new_new_n604_), .A1(new_new_n302_), .B0(new_new_n607_), .Y(new_new_n608_));
  AOI220     g586(.A0(i_7_), .A1(new_new_n68_), .B0(new_new_n348_), .B1(i_2_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n609_), .B(new_new_n222_), .Y(new_new_n610_));
  AOI210     g588(.A0(new_new_n403_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n611_));
  NOi31      g589(.An(new_new_n611_), .B(new_new_n533_), .C(new_new_n44_), .Y(new_new_n612_));
  NO3        g590(.A(new_new_n67_), .B(new_new_n32_), .C(new_new_n93_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n26_), .B(new_new_n178_), .Y(new_new_n614_));
  NO3        g592(.A(new_new_n434_), .B(new_new_n216_), .C(new_new_n80_), .Y(new_new_n615_));
  AOI210     g593(.A0(new_new_n615_), .A1(new_new_n26_), .B0(new_new_n613_), .Y(new_new_n616_));
  NO2        g594(.A(new_new_n616_), .B(i_9_), .Y(new_new_n617_));
  NO3        g595(.A(new_new_n617_), .B(new_new_n612_), .C(new_new_n610_), .Y(new_new_n618_));
  OR2        g596(.A(i_11_), .B(i_6_), .Y(new_new_n619_));
  NA3        g597(.A(new_new_n536_), .B(new_new_n614_), .C(i_7_), .Y(new_new_n620_));
  AOI210     g598(.A0(new_new_n620_), .A1(new_new_n569_), .B0(new_new_n619_), .Y(new_new_n621_));
  NA3        g599(.A(new_new_n369_), .B(new_new_n539_), .C(new_new_n89_), .Y(new_new_n622_));
  NA2        g600(.A(new_new_n562_), .B(i_13_), .Y(new_new_n623_));
  NA2        g601(.A(i_2_), .B(new_new_n614_), .Y(new_new_n624_));
  NAi21      g602(.An(i_11_), .B(i_12_), .Y(new_new_n625_));
  NOi41      g603(.An(new_new_n100_), .B(new_new_n625_), .C(i_13_), .D(new_new_n80_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n626_), .B(new_new_n624_), .Y(new_new_n627_));
  NA3        g605(.A(new_new_n627_), .B(new_new_n623_), .C(new_new_n622_), .Y(new_new_n628_));
  OAI210     g606(.A0(new_new_n628_), .A1(new_new_n621_), .B0(new_new_n62_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n216_), .B(new_new_n334_), .Y(new_new_n630_));
  NO2        g608(.A(new_new_n117_), .B(i_2_), .Y(new_new_n631_));
  NA2        g609(.A(new_new_n631_), .B(new_new_n559_), .Y(new_new_n632_));
  NA2        g610(.A(new_new_n632_), .B(new_new_n630_), .Y(new_new_n633_));
  NA3        g611(.A(new_new_n633_), .B(new_new_n45_), .C(new_new_n204_), .Y(new_new_n634_));
  NA4        g612(.A(new_new_n634_), .B(new_new_n629_), .C(new_new_n618_), .D(new_new_n608_), .Y(new_new_n635_));
  OR4        g613(.A(new_new_n635_), .B(new_new_n601_), .C(new_new_n589_), .D(new_new_n549_), .Y(mai5));
  NO2        g614(.A(i_4_), .B(i_11_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n83_), .B(new_new_n637_), .Y(new_new_n638_));
  INV        g616(.A(new_new_n638_), .Y(new_new_n639_));
  NO3        g617(.A(i_11_), .B(new_new_n216_), .C(i_13_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n114_), .B(new_new_n23_), .Y(new_new_n641_));
  NA2        g619(.A(i_12_), .B(i_8_), .Y(new_new_n642_));
  INV        g620(.A(new_new_n402_), .Y(new_new_n643_));
  NA2        g621(.A(new_new_n287_), .B(new_new_n514_), .Y(new_new_n644_));
  INV        g622(.A(new_new_n644_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n639_), .Y(new_new_n646_));
  INV        g624(.A(new_new_n158_), .Y(new_new_n647_));
  OAI210     g625(.A0(new_new_n599_), .A1(new_new_n404_), .B0(new_new_n100_), .Y(new_new_n648_));
  NO2        g626(.A(new_new_n648_), .B(new_new_n647_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n411_), .B(new_new_n26_), .Y(new_new_n650_));
  INV        g628(.A(new_new_n377_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n651_), .B(i_2_), .Y(new_new_n652_));
  INV        g630(.A(new_new_n652_), .Y(new_new_n653_));
  INV        g631(.A(new_new_n374_), .Y(new_new_n654_));
  AOI210     g632(.A0(new_new_n654_), .A1(new_new_n653_), .B0(new_new_n649_), .Y(new_new_n655_));
  OAI210     g633(.A0(new_new_n884_), .A1(new_new_n641_), .B0(i_2_), .Y(new_new_n656_));
  NO2        g634(.A(new_new_n38_), .B(new_new_n26_), .Y(new_new_n657_));
  AOI210     g635(.A0(new_new_n876_), .A1(new_new_n656_), .B0(new_new_n178_), .Y(new_new_n658_));
  OA210      g636(.A0(new_new_n551_), .A1(new_new_n116_), .B0(i_13_), .Y(new_new_n659_));
  INV        g637(.A(new_new_n77_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n660_), .B(new_new_n336_), .Y(new_new_n661_));
  NO2        g639(.A(new_new_n137_), .B(new_new_n467_), .Y(new_new_n662_));
  NA2        g640(.A(new_new_n662_), .B(new_new_n377_), .Y(new_new_n663_));
  NO2        g641(.A(i_2_), .B(new_new_n44_), .Y(new_new_n664_));
  NA3        g642(.A(new_new_n277_), .B(new_new_n114_), .C(new_new_n42_), .Y(new_new_n665_));
  OAI210     g643(.A0(new_new_n665_), .A1(new_new_n664_), .B0(new_new_n663_), .Y(new_new_n666_));
  NO4        g644(.A(new_new_n666_), .B(new_new_n661_), .C(new_new_n659_), .D(new_new_n658_), .Y(new_new_n667_));
  NA2        g645(.A(new_new_n514_), .B(new_new_n28_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n640_), .B(new_new_n250_), .Y(new_new_n669_));
  NA2        g647(.A(new_new_n669_), .B(new_new_n668_), .Y(new_new_n670_));
  NO2        g648(.A(i_7_), .B(new_new_n116_), .Y(new_new_n671_));
  NO2        g649(.A(new_new_n671_), .B(new_new_n534_), .Y(new_new_n672_));
  AOI220     g650(.A0(new_new_n672_), .A1(new_new_n36_), .B0(new_new_n670_), .B1(new_new_n46_), .Y(new_new_n673_));
  NA4        g651(.A(new_new_n673_), .B(new_new_n667_), .C(new_new_n655_), .D(new_new_n646_), .Y(mai6));
  NO2        g652(.A(new_new_n279_), .B(i_1_), .Y(new_new_n675_));
  NO2        g653(.A(new_new_n171_), .B(new_new_n128_), .Y(new_new_n676_));
  OAI210     g654(.A0(new_new_n676_), .A1(new_new_n675_), .B0(new_new_n631_), .Y(new_new_n677_));
  NA4        g655(.A(new_new_n352_), .B(new_new_n439_), .C(new_new_n67_), .D(new_new_n93_), .Y(new_new_n678_));
  INV        g656(.A(new_new_n678_), .Y(new_new_n679_));
  NO2        g657(.A(new_new_n679_), .B(new_new_n298_), .Y(new_new_n680_));
  AO210      g658(.A0(new_new_n680_), .A1(new_new_n677_), .B0(i_12_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n337_), .B(new_new_n305_), .Y(new_new_n682_));
  NA2        g660(.A(new_new_n522_), .B(new_new_n62_), .Y(new_new_n683_));
  INV        g661(.A(new_new_n591_), .Y(new_new_n684_));
  NA3        g662(.A(new_new_n684_), .B(new_new_n683_), .C(new_new_n682_), .Y(new_new_n685_));
  NA2        g663(.A(new_new_n685_), .B(new_new_n69_), .Y(new_new_n686_));
  INV        g664(.A(new_new_n297_), .Y(new_new_n687_));
  NA2        g665(.A(new_new_n71_), .B(new_new_n120_), .Y(new_new_n688_));
  AOI210     g666(.A0(new_new_n114_), .A1(new_new_n688_), .B0(new_new_n687_), .Y(new_new_n689_));
  NO2        g667(.A(new_new_n231_), .B(i_9_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n690_), .B(i_7_), .Y(new_new_n691_));
  NO2        g669(.A(new_new_n691_), .B(new_new_n171_), .Y(new_new_n692_));
  NA3        g670(.A(new_new_n879_), .B(new_new_n431_), .C(new_new_n352_), .Y(new_new_n693_));
  NAi32      g671(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n694_));
  AOI210     g672(.A0(new_new_n619_), .A1(new_new_n81_), .B0(new_new_n694_), .Y(new_new_n695_));
  NA2        g673(.A(new_new_n503_), .B(new_new_n502_), .Y(new_new_n696_));
  NAi31      g674(.An(new_new_n695_), .B(new_new_n696_), .C(new_new_n693_), .Y(new_new_n697_));
  OR3        g675(.A(new_new_n697_), .B(new_new_n692_), .C(new_new_n689_), .Y(new_new_n698_));
  OR2        g676(.A(new_new_n551_), .B(new_new_n404_), .Y(new_new_n699_));
  NA3        g677(.A(new_new_n699_), .B(new_new_n136_), .C(new_new_n66_), .Y(new_new_n700_));
  AO210      g678(.A0(new_new_n450_), .A1(new_new_n643_), .B0(new_new_n36_), .Y(new_new_n701_));
  NA2        g679(.A(new_new_n701_), .B(new_new_n700_), .Y(new_new_n702_));
  NA2        g680(.A(new_new_n878_), .B(new_new_n502_), .Y(new_new_n703_));
  INV        g681(.A(new_new_n703_), .Y(new_new_n704_));
  AO210      g682(.A0(new_new_n467_), .A1(new_new_n46_), .B0(new_new_n82_), .Y(new_new_n705_));
  NA2        g683(.A(new_new_n705_), .B(new_new_n440_), .Y(new_new_n706_));
  AOI210     g684(.A0(new_new_n404_), .A1(new_new_n402_), .B0(new_new_n501_), .Y(new_new_n707_));
  NA2        g685(.A(new_new_n101_), .B(new_new_n367_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n223_), .B(new_new_n46_), .Y(new_new_n709_));
  NA3        g687(.A(new_new_n708_), .B(new_new_n707_), .C(new_new_n706_), .Y(new_new_n710_));
  NO4        g688(.A(new_new_n710_), .B(new_new_n704_), .C(new_new_n702_), .D(new_new_n698_), .Y(new_new_n711_));
  NA4        g689(.A(new_new_n711_), .B(new_new_n686_), .C(new_new_n681_), .D(new_new_n342_), .Y(mai3));
  NO2        g690(.A(i_11_), .B(new_new_n216_), .Y(new_new_n713_));
  OAI210     g691(.A0(i_6_), .A1(new_new_n261_), .B0(new_new_n713_), .Y(new_new_n714_));
  NO2        g692(.A(new_new_n714_), .B(new_new_n178_), .Y(new_new_n715_));
  NO2        g693(.A(new_new_n407_), .B(new_new_n44_), .Y(new_new_n716_));
  OA210      g694(.A0(new_new_n716_), .A1(new_new_n715_), .B0(new_new_n161_), .Y(new_new_n717_));
  NA2        g695(.A(new_new_n369_), .B(new_new_n45_), .Y(new_new_n718_));
  NO4        g696(.A(new_new_n338_), .B(new_new_n345_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n171_), .B(new_new_n511_), .Y(new_new_n720_));
  NOi21      g698(.An(new_new_n720_), .B(new_new_n719_), .Y(new_new_n721_));
  NA2        g699(.A(new_new_n611_), .B(new_new_n583_), .Y(new_new_n722_));
  NA2        g700(.A(new_new_n303_), .B(i_5_), .Y(new_new_n723_));
  OAI220     g701(.A0(new_new_n723_), .A1(new_new_n722_), .B0(new_new_n721_), .B1(new_new_n62_), .Y(new_new_n724_));
  NOi21      g702(.An(i_5_), .B(i_9_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n725_), .B(new_new_n400_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n162_), .B(new_new_n137_), .Y(new_new_n727_));
  NA2        g705(.A(new_new_n727_), .B(new_new_n223_), .Y(new_new_n728_));
  OAI220     g706(.A0(new_new_n728_), .A1(new_new_n167_), .B0(i_1_), .B1(new_new_n726_), .Y(new_new_n729_));
  NO3        g707(.A(new_new_n729_), .B(new_new_n724_), .C(new_new_n717_), .Y(new_new_n730_));
  NA2        g708(.A(new_new_n171_), .B(new_new_n24_), .Y(new_new_n731_));
  NO2        g709(.A(new_new_n37_), .B(new_new_n731_), .Y(new_new_n732_));
  NA2        g710(.A(new_new_n284_), .B(new_new_n118_), .Y(new_new_n733_));
  NAi21      g711(.An(new_new_n149_), .B(i_5_), .Y(new_new_n734_));
  OAI220     g712(.A0(new_new_n734_), .A1(new_new_n709_), .B0(new_new_n733_), .B1(new_new_n361_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n735_), .B(new_new_n732_), .Y(new_new_n736_));
  NA2        g714(.A(i_9_), .B(i_0_), .Y(new_new_n737_));
  NO3        g715(.A(new_new_n737_), .B(new_new_n347_), .C(new_new_n83_), .Y(new_new_n738_));
  INV        g716(.A(new_new_n738_), .Y(new_new_n739_));
  INV        g717(.A(new_new_n431_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n640_), .B(new_new_n298_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n576_), .B(i_5_), .Y(new_new_n742_));
  NO2        g720(.A(new_new_n233_), .B(new_new_n140_), .Y(new_new_n743_));
  NA2        g721(.A(i_0_), .B(i_10_), .Y(new_new_n744_));
  AN2        g722(.A(new_new_n743_), .B(i_6_), .Y(new_new_n745_));
  NO2        g723(.A(i_1_), .B(new_new_n741_), .Y(new_new_n746_));
  NO3        g724(.A(new_new_n746_), .B(new_new_n745_), .C(new_new_n742_), .Y(new_new_n747_));
  NA3        g725(.A(new_new_n747_), .B(new_new_n739_), .C(new_new_n736_), .Y(new_new_n748_));
  NA2        g726(.A(i_11_), .B(i_9_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n48_), .B(i_7_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n357_), .B(new_new_n165_), .Y(new_new_n751_));
  NA2        g729(.A(new_new_n751_), .B(new_new_n147_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n162_), .B(i_0_), .Y(new_new_n753_));
  NA2        g731(.A(new_new_n431_), .B(new_new_n210_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n754_), .B(new_new_n162_), .Y(new_new_n755_));
  NO2        g733(.A(new_new_n755_), .B(new_new_n752_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n575_), .B(new_new_n111_), .Y(new_new_n757_));
  NO2        g735(.A(i_6_), .B(new_new_n757_), .Y(new_new_n758_));
  AOI210     g736(.A0(new_new_n403_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n759_));
  INV        g737(.A(new_new_n94_), .Y(new_new_n760_));
  NOi32      g738(.An(new_new_n759_), .Bn(new_new_n173_), .C(new_new_n760_), .Y(new_new_n761_));
  NA2        g739(.A(new_new_n539_), .B(new_new_n298_), .Y(new_new_n762_));
  NO2        g740(.A(new_new_n762_), .B(new_new_n718_), .Y(new_new_n763_));
  NO3        g741(.A(new_new_n763_), .B(new_new_n761_), .C(new_new_n758_), .Y(new_new_n764_));
  NOi21      g742(.An(i_7_), .B(i_5_), .Y(new_new_n765_));
  NOi31      g743(.An(new_new_n765_), .B(i_0_), .C(new_new_n625_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n235_), .B(new_new_n288_), .Y(new_new_n767_));
  INV        g745(.A(new_new_n625_), .Y(new_new_n768_));
  NA2        g746(.A(new_new_n768_), .B(new_new_n767_), .Y(new_new_n769_));
  NA3        g747(.A(new_new_n769_), .B(new_new_n764_), .C(new_new_n756_), .Y(new_new_n770_));
  NO2        g748(.A(new_new_n731_), .B(new_new_n219_), .Y(new_new_n771_));
  AN2        g749(.A(new_new_n302_), .B(new_new_n298_), .Y(new_new_n772_));
  AN2        g750(.A(new_new_n772_), .B(new_new_n727_), .Y(new_new_n773_));
  OAI210     g751(.A0(new_new_n773_), .A1(new_new_n771_), .B0(i_10_), .Y(new_new_n774_));
  NA3        g752(.A(new_new_n430_), .B(new_new_n369_), .C(new_new_n45_), .Y(new_new_n775_));
  OAI210     g753(.A0(new_new_n734_), .A1(new_new_n740_), .B0(new_new_n775_), .Y(new_new_n776_));
  NA2        g754(.A(i_0_), .B(new_new_n277_), .Y(new_new_n777_));
  NA2        g755(.A(new_new_n172_), .B(new_new_n777_), .Y(new_new_n778_));
  AOI220     g756(.A0(new_new_n778_), .A1(new_new_n431_), .B0(new_new_n776_), .B1(new_new_n69_), .Y(new_new_n779_));
  NO2        g757(.A(new_new_n71_), .B(new_new_n642_), .Y(new_new_n780_));
  AOI210     g758(.A0(new_new_n161_), .A1(new_new_n532_), .B0(new_new_n780_), .Y(new_new_n781_));
  NO2        g759(.A(new_new_n781_), .B(new_new_n47_), .Y(new_new_n782_));
  NO3        g760(.A(i_5_), .B(new_new_n325_), .C(new_new_n24_), .Y(new_new_n783_));
  INV        g761(.A(new_new_n783_), .Y(new_new_n784_));
  NO2        g762(.A(new_new_n535_), .B(new_new_n95_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n785_), .B(i_0_), .Y(new_new_n786_));
  OAI220     g764(.A0(new_new_n786_), .A1(new_new_n80_), .B0(new_new_n784_), .B1(new_new_n159_), .Y(new_new_n787_));
  NO3        g765(.A(new_new_n787_), .B(new_new_n782_), .C(new_new_n470_), .Y(new_new_n788_));
  NA3        g766(.A(new_new_n788_), .B(new_new_n779_), .C(new_new_n774_), .Y(new_new_n789_));
  NO3        g767(.A(new_new_n789_), .B(new_new_n770_), .C(new_new_n748_), .Y(new_new_n790_));
  NO2        g768(.A(i_0_), .B(new_new_n625_), .Y(new_new_n791_));
  NO2        g769(.A(new_new_n683_), .B(new_new_n760_), .Y(new_new_n792_));
  INV        g770(.A(new_new_n792_), .Y(new_new_n793_));
  NA3        g771(.A(new_new_n135_), .B(new_new_n583_), .C(new_new_n69_), .Y(new_new_n794_));
  NA3        g772(.A(i_6_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n795_));
  NA2        g773(.A(new_new_n713_), .B(i_9_), .Y(new_new_n796_));
  AOI210     g774(.A0(new_new_n795_), .A1(new_new_n454_), .B0(new_new_n796_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n223_), .B(new_new_n209_), .Y(new_new_n798_));
  AOI210     g776(.A0(new_new_n798_), .A1(new_new_n737_), .B0(new_new_n140_), .Y(new_new_n799_));
  NO2        g777(.A(new_new_n799_), .B(new_new_n797_), .Y(new_new_n800_));
  NA3        g778(.A(new_new_n800_), .B(new_new_n794_), .C(new_new_n793_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n772_), .B(new_new_n336_), .Y(new_new_n802_));
  AOI210     g780(.A0(new_new_n272_), .A1(new_new_n149_), .B0(new_new_n802_), .Y(new_new_n803_));
  NA2        g781(.A(new_new_n750_), .B(new_new_n444_), .Y(new_new_n804_));
  NO2        g782(.A(new_new_n149_), .B(new_new_n804_), .Y(new_new_n805_));
  NO2        g783(.A(new_new_n805_), .B(new_new_n803_), .Y(new_new_n806_));
  NO2        g784(.A(new_new_n744_), .B(new_new_n175_), .Y(new_new_n807_));
  AOI220     g785(.A0(new_new_n807_), .A1(i_11_), .B0(new_new_n507_), .B1(new_new_n71_), .Y(new_new_n808_));
  NO3        g786(.A(new_new_n193_), .B(new_new_n345_), .C(i_0_), .Y(new_new_n809_));
  OAI210     g787(.A0(new_new_n809_), .A1(new_new_n72_), .B0(i_13_), .Y(new_new_n810_));
  INV        g788(.A(new_new_n201_), .Y(new_new_n811_));
  NO2        g789(.A(i_13_), .B(new_new_n128_), .Y(new_new_n812_));
  NA3        g790(.A(new_new_n812_), .B(i_7_), .C(new_new_n811_), .Y(new_new_n813_));
  NA4        g791(.A(new_new_n813_), .B(new_new_n810_), .C(new_new_n808_), .D(new_new_n806_), .Y(new_new_n814_));
  AOI210     g792(.A0(i_6_), .A1(new_new_n791_), .B0(new_new_n98_), .Y(new_new_n815_));
  NA2        g793(.A(new_new_n765_), .B(new_new_n444_), .Y(new_new_n816_));
  OA220      g794(.A0(new_new_n162_), .A1(new_new_n816_), .B0(new_new_n815_), .B1(i_5_), .Y(new_new_n817_));
  NO2        g795(.A(i_0_), .B(new_new_n162_), .Y(new_new_n818_));
  NO3        g796(.A(new_new_n718_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n819_));
  INV        g797(.A(new_new_n449_), .Y(new_new_n820_));
  NO2        g798(.A(new_new_n820_), .B(new_new_n819_), .Y(new_new_n821_));
  NA3        g799(.A(new_new_n750_), .B(new_new_n261_), .C(new_new_n209_), .Y(new_new_n822_));
  INV        g800(.A(new_new_n822_), .Y(new_new_n823_));
  NA3        g801(.A(new_new_n352_), .B(new_new_n304_), .C(i_4_), .Y(new_new_n824_));
  INV        g802(.A(new_new_n824_), .Y(new_new_n825_));
  NOi31      g803(.An(new_new_n351_), .B(i_11_), .C(new_new_n219_), .Y(new_new_n826_));
  NO3        g804(.A(new_new_n749_), .B(new_new_n201_), .C(new_new_n175_), .Y(new_new_n827_));
  NO4        g805(.A(new_new_n827_), .B(new_new_n826_), .C(new_new_n825_), .D(new_new_n823_), .Y(new_new_n828_));
  NA3        g806(.A(new_new_n828_), .B(new_new_n821_), .C(new_new_n817_), .Y(new_new_n829_));
  NA3        g807(.A(new_new_n277_), .B(i_5_), .C(new_new_n178_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n830_), .B(new_new_n222_), .Y(new_new_n831_));
  NO3        g809(.A(new_new_n219_), .B(i_0_), .C(i_12_), .Y(new_new_n832_));
  AOI210     g810(.A0(new_new_n832_), .A1(new_new_n831_), .B0(new_new_n679_), .Y(new_new_n833_));
  AN2        g811(.A(new_new_n744_), .B(new_new_n140_), .Y(new_new_n834_));
  NO3        g812(.A(new_new_n834_), .B(i_12_), .C(new_new_n567_), .Y(new_new_n835_));
  INV        g813(.A(new_new_n835_), .Y(new_new_n836_));
  NA3        g814(.A(new_new_n90_), .B(new_new_n511_), .C(i_11_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n837_), .B(new_new_n142_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n765_), .B(new_new_n428_), .Y(new_new_n839_));
  OAI220     g817(.A0(i_7_), .A1(new_new_n830_), .B0(new_new_n839_), .B1(new_new_n584_), .Y(new_new_n840_));
  AOI210     g818(.A0(new_new_n840_), .A1(new_new_n753_), .B0(new_new_n838_), .Y(new_new_n841_));
  NA3        g819(.A(new_new_n841_), .B(new_new_n836_), .C(new_new_n833_), .Y(new_new_n842_));
  NO4        g820(.A(new_new_n842_), .B(new_new_n829_), .C(new_new_n814_), .D(new_new_n801_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n879_), .B(new_new_n37_), .Y(new_new_n844_));
  NA2        g822(.A(new_new_n844_), .B(new_new_n543_), .Y(new_new_n845_));
  NA2        g823(.A(new_new_n845_), .B(new_new_n190_), .Y(new_new_n846_));
  OR2        g824(.A(i_11_), .B(i_2_), .Y(new_new_n847_));
  NO2        g825(.A(new_new_n419_), .B(new_new_n241_), .Y(new_new_n848_));
  AOI210     g826(.A0(new_new_n882_), .A1(new_new_n48_), .B0(new_new_n848_), .Y(new_new_n849_));
  AOI210     g827(.A0(new_new_n849_), .A1(new_new_n846_), .B0(new_new_n69_), .Y(new_new_n850_));
  NO2        g828(.A(new_new_n504_), .B(new_new_n341_), .Y(new_new_n851_));
  NO2        g829(.A(new_new_n851_), .B(new_new_n647_), .Y(new_new_n852_));
  INV        g830(.A(new_new_n72_), .Y(new_new_n853_));
  AOI210     g831(.A0(new_new_n818_), .A1(new_new_n750_), .B0(new_new_n766_), .Y(new_new_n854_));
  AOI210     g832(.A0(new_new_n854_), .A1(new_new_n853_), .B0(new_new_n587_), .Y(new_new_n855_));
  NA2        g833(.A(i_8_), .B(new_new_n72_), .Y(new_new_n856_));
  NO2        g834(.A(new_new_n856_), .B(new_new_n216_), .Y(new_new_n857_));
  NA2        g835(.A(new_new_n88_), .B(new_new_n279_), .Y(new_new_n858_));
  INV        g836(.A(new_new_n858_), .Y(new_new_n859_));
  NO3        g837(.A(new_new_n859_), .B(new_new_n857_), .C(new_new_n855_), .Y(new_new_n860_));
  OAI210     g838(.A0(new_new_n243_), .A1(new_new_n145_), .B0(new_new_n83_), .Y(new_new_n861_));
  NA2        g839(.A(new_new_n650_), .B(new_new_n261_), .Y(new_new_n862_));
  AOI210     g840(.A0(new_new_n862_), .A1(new_new_n861_), .B0(i_11_), .Y(new_new_n863_));
  NO4        g841(.A(i_9_), .B(i_11_), .C(new_new_n232_), .D(new_new_n231_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n864_), .B(new_new_n501_), .Y(new_new_n865_));
  INV        g843(.A(new_new_n331_), .Y(new_new_n866_));
  AOI210     g844(.A0(new_new_n866_), .A1(new_new_n865_), .B0(new_new_n41_), .Y(new_new_n867_));
  NO2        g845(.A(new_new_n867_), .B(new_new_n863_), .Y(new_new_n868_));
  OAI210     g846(.A0(new_new_n860_), .A1(i_4_), .B0(new_new_n868_), .Y(new_new_n869_));
  NO3        g847(.A(new_new_n869_), .B(new_new_n852_), .C(new_new_n850_), .Y(new_new_n870_));
  NA4        g848(.A(new_new_n870_), .B(new_new_n843_), .C(new_new_n790_), .D(new_new_n730_), .Y(mai4));
  INV        g849(.A(new_new_n605_), .Y(new_new_n874_));
  INV        g850(.A(i_2_), .Y(new_new_n875_));
  INV        g851(.A(new_new_n657_), .Y(new_new_n876_));
  INV        g852(.A(new_new_n203_), .Y(new_new_n877_));
  INV        g853(.A(i_11_), .Y(new_new_n878_));
  INV        g854(.A(i_11_), .Y(new_new_n879_));
  INV        g855(.A(new_new_n402_), .Y(new_new_n880_));
  INV        g856(.A(i_7_), .Y(new_new_n881_));
  INV        g857(.A(new_new_n847_), .Y(new_new_n882_));
  INV        g858(.A(i_13_), .Y(new_new_n883_));
  INV        g859(.A(new_new_n175_), .Y(new_new_n884_));
endmodule


