library verilog;
use verilog.vl_types.all;
entity ContadorDe1_vlg_vec_tst is
end ContadorDe1_vlg_vec_tst;
