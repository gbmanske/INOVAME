//Benchmark atmr_9sym_175_0.5

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, ori00, mai00, men00;
  ONE        o0(.Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NA3        m013(.A(i_6_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_8_), .B(i_6_), .Y(mai_mai_n25_));
  NO2        m015(.A(mai_mai_n24_), .B(mai_mai_n22_), .Y(mai_mai_n26_));
  AOI210     m016(.A0(mai_mai_n26_), .A1(mai_mai_n11_), .B0(mai_mai_n20_), .Y(mai_mai_n27_));
  INV        m017(.A(i_2_), .Y(mai_mai_n28_));
  NOi21      m018(.An(i_5_), .B(i_0_), .Y(mai_mai_n29_));
  NOi21      m019(.An(i_6_), .B(i_8_), .Y(mai_mai_n30_));
  NOi21      m020(.An(i_7_), .B(i_1_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_5_), .B(i_6_), .Y(mai_mai_n32_));
  AOI220     m022(.A0(mai_mai_n32_), .A1(mai_mai_n31_), .B0(mai_mai_n30_), .B1(mai_mai_n29_), .Y(mai_mai_n33_));
  NO3        m023(.A(mai_mai_n33_), .B(mai_mai_n28_), .C(i_4_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_0_), .B(i_4_), .Y(mai_mai_n35_));
  XO2        m025(.A(i_1_), .B(i_3_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_7_), .B(i_5_), .Y(mai_mai_n37_));
  AN3        m027(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(mai_mai_n35_), .Y(mai_mai_n38_));
  INV        m028(.A(i_1_), .Y(mai_mai_n39_));
  NOi21      m029(.An(i_3_), .B(i_0_), .Y(mai_mai_n40_));
  NA2        m030(.A(mai_mai_n40_), .B(mai_mai_n39_), .Y(mai_mai_n41_));
  NA3        m031(.A(i_6_), .B(mai_mai_n14_), .C(i_7_), .Y(mai_mai_n42_));
  AOI210     m032(.A0(mai_mai_n42_), .A1(mai_mai_n24_), .B0(mai_mai_n41_), .Y(mai_mai_n43_));
  NO3        m033(.A(mai_mai_n43_), .B(mai_mai_n38_), .C(mai_mai_n34_), .Y(mai_mai_n44_));
  NOi21      m034(.An(i_4_), .B(i_0_), .Y(mai_mai_n45_));
  NA2        m035(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n46_));
  NOi21      m036(.An(i_2_), .B(i_8_), .Y(mai_mai_n47_));
  NOi31      m037(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n48_));
  NA2        m038(.A(mai_mai_n48_), .B(i_0_), .Y(mai_mai_n49_));
  NOi21      m039(.An(i_4_), .B(i_3_), .Y(mai_mai_n50_));
  NOi21      m040(.An(i_1_), .B(i_4_), .Y(mai_mai_n51_));
  OAI210     m041(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n52_));
  NA2        m042(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  AN2        m043(.A(i_8_), .B(i_7_), .Y(mai_mai_n54_));
  NA2        m044(.A(mai_mai_n54_), .B(mai_mai_n12_), .Y(mai_mai_n55_));
  NOi21      m045(.An(i_8_), .B(i_7_), .Y(mai_mai_n56_));
  NA3        m046(.A(mai_mai_n56_), .B(mai_mai_n50_), .C(i_6_), .Y(mai_mai_n57_));
  OAI210     m047(.A0(mai_mai_n55_), .A1(mai_mai_n46_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  AOI220     m048(.A0(mai_mai_n58_), .A1(mai_mai_n28_), .B0(mai_mai_n53_), .B1(mai_mai_n32_), .Y(mai_mai_n59_));
  NA3        m049(.A(mai_mai_n59_), .B(mai_mai_n44_), .C(mai_mai_n27_), .Y(mai_mai_n60_));
  NA2        m050(.A(i_8_), .B(i_7_), .Y(mai_mai_n61_));
  NO3        m051(.A(mai_mai_n61_), .B(mai_mai_n13_), .C(i_1_), .Y(mai_mai_n62_));
  NA2        m052(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n63_));
  AOI220     m053(.A0(mai_mai_n40_), .A1(i_1_), .B0(mai_mai_n36_), .B1(i_2_), .Y(mai_mai_n64_));
  NOi21      m054(.An(i_1_), .B(i_2_), .Y(mai_mai_n65_));
  NA3        m055(.A(mai_mai_n65_), .B(mai_mai_n45_), .C(i_6_), .Y(mai_mai_n66_));
  OAI210     m056(.A0(mai_mai_n64_), .A1(mai_mai_n63_), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  OAI210     m057(.A0(mai_mai_n67_), .A1(mai_mai_n62_), .B0(mai_mai_n14_), .Y(mai_mai_n68_));
  INV        m058(.A(mai_mai_n68_), .Y(mai_mai_n69_));
  NA2        m059(.A(mai_mai_n30_), .B(mai_mai_n29_), .Y(mai_mai_n70_));
  NOi21      m060(.An(i_7_), .B(i_8_), .Y(mai_mai_n71_));
  INV        m061(.A(mai_mai_n70_), .Y(mai_mai_n72_));
  NA2        m062(.A(mai_mai_n72_), .B(mai_mai_n65_), .Y(mai_mai_n73_));
  AOI220     m063(.A0(mai_mai_n40_), .A1(mai_mai_n39_), .B0(mai_mai_n18_), .B1(mai_mai_n28_), .Y(mai_mai_n74_));
  NA3        m064(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n75_));
  NO2        m065(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n76_));
  INV        m066(.A(mai_mai_n76_), .Y(mai_mai_n77_));
  NA3        m067(.A(mai_mai_n56_), .B(mai_mai_n28_), .C(i_3_), .Y(mai_mai_n78_));
  NA2        m068(.A(mai_mai_n39_), .B(i_6_), .Y(mai_mai_n79_));
  AOI210     m069(.A0(mai_mai_n79_), .A1(mai_mai_n22_), .B0(mai_mai_n78_), .Y(mai_mai_n80_));
  NAi21      m070(.An(i_6_), .B(i_0_), .Y(mai_mai_n81_));
  NA3        m071(.A(mai_mai_n51_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n82_));
  NOi21      m072(.An(i_4_), .B(i_6_), .Y(mai_mai_n83_));
  NOi21      m073(.An(i_5_), .B(i_3_), .Y(mai_mai_n84_));
  NA3        m074(.A(mai_mai_n84_), .B(mai_mai_n65_), .C(mai_mai_n83_), .Y(mai_mai_n85_));
  OAI210     m075(.A0(mai_mai_n82_), .A1(mai_mai_n81_), .B0(mai_mai_n85_), .Y(mai_mai_n86_));
  NO2        m076(.A(mai_mai_n86_), .B(mai_mai_n80_), .Y(mai_mai_n87_));
  NOi21      m077(.An(i_6_), .B(i_1_), .Y(mai_mai_n88_));
  AOI220     m078(.A0(mai_mai_n88_), .A1(i_7_), .B0(mai_mai_n25_), .B1(i_5_), .Y(mai_mai_n89_));
  NOi31      m079(.An(mai_mai_n45_), .B(mai_mai_n89_), .C(i_2_), .Y(mai_mai_n90_));
  INV        m080(.A(mai_mai_n90_), .Y(mai_mai_n91_));
  NA4        m081(.A(mai_mai_n91_), .B(mai_mai_n87_), .C(mai_mai_n77_), .D(mai_mai_n73_), .Y(mai_mai_n92_));
  NA2        m082(.A(mai_mai_n47_), .B(mai_mai_n15_), .Y(mai_mai_n93_));
  NA3        m083(.A(mai_mai_n30_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n94_));
  NA2        m084(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n95_));
  NA2        m085(.A(mai_mai_n95_), .B(mai_mai_n35_), .Y(mai_mai_n96_));
  NA3        m086(.A(mai_mai_n56_), .B(mai_mai_n48_), .C(i_6_), .Y(mai_mai_n97_));
  INV        m087(.A(mai_mai_n97_), .Y(mai_mai_n98_));
  NOi21      m088(.An(i_0_), .B(i_2_), .Y(mai_mai_n99_));
  NA3        m089(.A(mai_mai_n99_), .B(mai_mai_n31_), .C(mai_mai_n83_), .Y(mai_mai_n100_));
  NA3        m090(.A(mai_mai_n99_), .B(mai_mai_n50_), .C(mai_mai_n30_), .Y(mai_mai_n101_));
  NA2        m091(.A(mai_mai_n101_), .B(mai_mai_n100_), .Y(mai_mai_n102_));
  NA4        m092(.A(mai_mai_n48_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n103_));
  NA4        m093(.A(mai_mai_n51_), .B(mai_mai_n32_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n104_));
  NA2        m094(.A(mai_mai_n104_), .B(mai_mai_n103_), .Y(mai_mai_n105_));
  NO3        m095(.A(mai_mai_n105_), .B(mai_mai_n102_), .C(mai_mai_n98_), .Y(mai_mai_n106_));
  NO2        m096(.A(mai_mai_n93_), .B(mai_mai_n79_), .Y(mai_mai_n107_));
  INV        m097(.A(mai_mai_n107_), .Y(mai_mai_n108_));
  NA2        m098(.A(mai_mai_n71_), .B(mai_mai_n12_), .Y(mai_mai_n109_));
  NA3        m099(.A(i_2_), .B(i_1_), .C(mai_mai_n14_), .Y(mai_mai_n110_));
  NA2        m100(.A(mai_mai_n45_), .B(i_3_), .Y(mai_mai_n111_));
  AOI210     m101(.A0(mai_mai_n111_), .A1(mai_mai_n110_), .B0(mai_mai_n109_), .Y(mai_mai_n112_));
  NA3        m102(.A(mai_mai_n99_), .B(mai_mai_n56_), .C(mai_mai_n83_), .Y(mai_mai_n113_));
  INV        m103(.A(mai_mai_n113_), .Y(mai_mai_n114_));
  NA4        m104(.A(mai_mai_n84_), .B(mai_mai_n54_), .C(mai_mai_n39_), .D(mai_mai_n21_), .Y(mai_mai_n115_));
  NA3        m105(.A(mai_mai_n47_), .B(mai_mai_n29_), .C(mai_mai_n15_), .Y(mai_mai_n116_));
  NA2        m106(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NO3        m107(.A(mai_mai_n117_), .B(mai_mai_n114_), .C(mai_mai_n112_), .Y(mai_mai_n118_));
  NA4        m108(.A(mai_mai_n118_), .B(mai_mai_n108_), .C(mai_mai_n106_), .D(mai_mai_n96_), .Y(mai_mai_n119_));
  OR4        m109(.A(mai_mai_n119_), .B(mai_mai_n92_), .C(mai_mai_n69_), .D(mai_mai_n60_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  INV        u002(.A(i_5_), .Y(men_men_n13_));
  NOi21      u003(.An(i_3_), .B(i_7_), .Y(men_men_n14_));
  INV        u004(.A(i_0_), .Y(men_men_n15_));
  NOi21      u005(.An(i_1_), .B(i_3_), .Y(men_men_n16_));
  INV        u006(.A(i_4_), .Y(men_men_n17_));
  NA2        u007(.A(i_0_), .B(men_men_n17_), .Y(men_men_n18_));
  INV        u008(.A(i_7_), .Y(men_men_n19_));
  NOi21      u009(.An(i_8_), .B(i_6_), .Y(men_men_n20_));
  NOi21      u010(.An(i_1_), .B(i_8_), .Y(men_men_n21_));
  AOI220     u011(.A0(men_men_n21_), .A1(i_2_), .B0(men_men_n20_), .B1(i_5_), .Y(men_men_n22_));
  NO2        u012(.A(men_men_n22_), .B(men_men_n18_), .Y(men_men_n23_));
  NA2        u013(.A(men_men_n23_), .B(men_men_n11_), .Y(men_men_n24_));
  NA2        u014(.A(i_0_), .B(men_men_n13_), .Y(men_men_n25_));
  NA2        u015(.A(men_men_n15_), .B(i_5_), .Y(men_men_n26_));
  NO2        u016(.A(i_2_), .B(i_4_), .Y(men_men_n27_));
  NA3        u017(.A(men_men_n27_), .B(i_6_), .C(i_8_), .Y(men_men_n28_));
  AOI210     u018(.A0(men_men_n26_), .A1(men_men_n25_), .B0(men_men_n28_), .Y(men_men_n29_));
  INV        u019(.A(i_2_), .Y(men_men_n30_));
  NOi21      u020(.An(i_6_), .B(i_8_), .Y(men_men_n31_));
  NOi21      u021(.An(i_7_), .B(i_1_), .Y(men_men_n32_));
  NOi21      u022(.An(i_0_), .B(i_4_), .Y(men_men_n33_));
  NOi21      u023(.An(i_7_), .B(i_5_), .Y(men_men_n34_));
  INV        u024(.A(i_1_), .Y(men_men_n35_));
  NOi21      u025(.An(i_3_), .B(i_0_), .Y(men_men_n36_));
  INV        u026(.A(men_men_n29_), .Y(men_men_n37_));
  INV        u027(.A(i_8_), .Y(men_men_n38_));
  NA2        u028(.A(i_1_), .B(men_men_n11_), .Y(men_men_n39_));
  NO4        u029(.A(men_men_n39_), .B(men_men_n25_), .C(i_2_), .D(men_men_n38_), .Y(men_men_n40_));
  NOi21      u030(.An(i_4_), .B(i_0_), .Y(men_men_n41_));
  AOI210     u031(.A0(men_men_n41_), .A1(men_men_n20_), .B0(men_men_n14_), .Y(men_men_n42_));
  NA2        u032(.A(i_1_), .B(men_men_n13_), .Y(men_men_n43_));
  NOi21      u033(.An(i_2_), .B(i_8_), .Y(men_men_n44_));
  NO3        u034(.A(men_men_n44_), .B(men_men_n41_), .C(men_men_n33_), .Y(men_men_n45_));
  NO3        u035(.A(men_men_n45_), .B(men_men_n43_), .C(men_men_n42_), .Y(men_men_n46_));
  NO2        u036(.A(men_men_n46_), .B(men_men_n40_), .Y(men_men_n47_));
  NOi21      u037(.An(i_4_), .B(i_3_), .Y(men_men_n48_));
  NOi21      u038(.An(i_1_), .B(i_4_), .Y(men_men_n49_));
  AN2        u039(.A(i_8_), .B(i_7_), .Y(men_men_n50_));
  NOi21      u040(.An(i_8_), .B(i_7_), .Y(men_men_n51_));
  NA3        u041(.A(men_men_n47_), .B(men_men_n37_), .C(men_men_n24_), .Y(men_men_n52_));
  NA2        u042(.A(i_8_), .B(i_7_), .Y(men_men_n53_));
  NOi21      u043(.An(i_1_), .B(i_2_), .Y(men_men_n54_));
  NA3        u044(.A(men_men_n51_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n55_));
  NA3        u045(.A(men_men_n21_), .B(i_0_), .C(men_men_n13_), .Y(men_men_n56_));
  NA2        u046(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  NOi32      u047(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n58_), .B(i_3_), .Y(men_men_n59_));
  NA3        u049(.A(men_men_n16_), .B(i_2_), .C(i_6_), .Y(men_men_n60_));
  NA2        u050(.A(men_men_n60_), .B(men_men_n59_), .Y(men_men_n61_));
  NO2        u051(.A(i_0_), .B(i_4_), .Y(men_men_n62_));
  AOI220     u052(.A0(men_men_n62_), .A1(men_men_n61_), .B0(men_men_n57_), .B1(men_men_n48_), .Y(men_men_n63_));
  INV        u053(.A(men_men_n63_), .Y(men_men_n64_));
  NAi21      u054(.An(i_3_), .B(i_6_), .Y(men_men_n65_));
  NO3        u055(.A(men_men_n65_), .B(i_0_), .C(men_men_n38_), .Y(men_men_n66_));
  NOi21      u056(.An(i_7_), .B(i_8_), .Y(men_men_n67_));
  NOi31      u057(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n68_));
  AOI210     u058(.A0(men_men_n67_), .A1(men_men_n12_), .B0(men_men_n68_), .Y(men_men_n69_));
  NO2        u059(.A(men_men_n69_), .B(men_men_n11_), .Y(men_men_n70_));
  OAI210     u060(.A0(men_men_n70_), .A1(men_men_n66_), .B0(men_men_n54_), .Y(men_men_n71_));
  NA3        u061(.A(men_men_n20_), .B(i_2_), .C(men_men_n13_), .Y(men_men_n72_));
  AOI210     u062(.A0(men_men_n18_), .A1(men_men_n39_), .B0(men_men_n72_), .Y(men_men_n73_));
  OAI210     u063(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n74_));
  NA3        u064(.A(men_men_n53_), .B(men_men_n16_), .C(men_men_n15_), .Y(men_men_n75_));
  NO2        u065(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  NO2        u066(.A(men_men_n76_), .B(men_men_n73_), .Y(men_men_n77_));
  NA3        u067(.A(men_men_n51_), .B(men_men_n30_), .C(i_3_), .Y(men_men_n78_));
  NA2        u068(.A(men_men_n35_), .B(i_6_), .Y(men_men_n79_));
  NOi21      u069(.An(i_2_), .B(i_1_), .Y(men_men_n80_));
  AN3        u070(.A(men_men_n67_), .B(men_men_n80_), .C(men_men_n41_), .Y(men_men_n81_));
  NAi21      u071(.An(i_6_), .B(i_0_), .Y(men_men_n82_));
  NOi21      u072(.An(i_4_), .B(i_6_), .Y(men_men_n83_));
  NA2        u073(.A(men_men_n54_), .B(men_men_n31_), .Y(men_men_n84_));
  NOi21      u074(.An(men_men_n34_), .B(men_men_n84_), .Y(men_men_n85_));
  NO2        u075(.A(men_men_n85_), .B(men_men_n81_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n51_), .B(men_men_n12_), .Y(men_men_n87_));
  NA2        u077(.A(men_men_n31_), .B(men_men_n13_), .Y(men_men_n88_));
  NOi21      u078(.An(i_3_), .B(i_1_), .Y(men_men_n89_));
  NA2        u079(.A(men_men_n89_), .B(i_4_), .Y(men_men_n90_));
  AOI210     u080(.A0(men_men_n88_), .A1(men_men_n87_), .B0(men_men_n90_), .Y(men_men_n91_));
  AOI220     u081(.A0(men_men_n67_), .A1(men_men_n13_), .B0(men_men_n83_), .B1(men_men_n19_), .Y(men_men_n92_));
  NOi31      u082(.An(men_men_n36_), .B(men_men_n92_), .C(men_men_n30_), .Y(men_men_n93_));
  NO2        u083(.A(men_men_n93_), .B(men_men_n91_), .Y(men_men_n94_));
  NA4        u084(.A(men_men_n94_), .B(men_men_n86_), .C(men_men_n77_), .D(men_men_n71_), .Y(men_men_n95_));
  NOi31      u085(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n96_));
  NOi31      u086(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n97_));
  OAI210     u087(.A0(men_men_n97_), .A1(men_men_n96_), .B0(i_7_), .Y(men_men_n98_));
  NA2        u088(.A(men_men_n98_), .B(men_men_n84_), .Y(men_men_n99_));
  NA2        u089(.A(men_men_n99_), .B(men_men_n33_), .Y(men_men_n100_));
  NA2        u090(.A(men_men_n48_), .B(men_men_n32_), .Y(men_men_n101_));
  AOI210     u091(.A0(men_men_n101_), .A1(men_men_n55_), .B0(men_men_n26_), .Y(men_men_n102_));
  NA4        u092(.A(men_men_n50_), .B(men_men_n80_), .C(men_men_n15_), .D(men_men_n12_), .Y(men_men_n103_));
  NAi31      u093(.An(men_men_n82_), .B(men_men_n67_), .C(men_men_n80_), .Y(men_men_n104_));
  NA2        u094(.A(men_men_n104_), .B(men_men_n103_), .Y(men_men_n105_));
  NA3        u095(.A(men_men_n41_), .B(men_men_n34_), .C(men_men_n16_), .Y(men_men_n106_));
  NOi32      u096(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n107_));
  NA2        u097(.A(men_men_n107_), .B(men_men_n96_), .Y(men_men_n108_));
  NA2        u098(.A(men_men_n108_), .B(men_men_n106_), .Y(men_men_n109_));
  NA4        u099(.A(men_men_n49_), .B(men_men_n36_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n110_));
  INV        u100(.A(men_men_n110_), .Y(men_men_n111_));
  NO4        u101(.A(men_men_n111_), .B(men_men_n109_), .C(men_men_n105_), .D(men_men_n102_), .Y(men_men_n112_));
  NOi21      u102(.An(i_5_), .B(i_2_), .Y(men_men_n113_));
  AOI220     u103(.A0(men_men_n113_), .A1(men_men_n67_), .B0(men_men_n50_), .B1(men_men_n27_), .Y(men_men_n114_));
  NO2        u104(.A(men_men_n114_), .B(men_men_n79_), .Y(men_men_n115_));
  NO4        u105(.A(i_2_), .B(men_men_n17_), .C(men_men_n11_), .D(men_men_n13_), .Y(men_men_n116_));
  NA2        u106(.A(i_2_), .B(i_4_), .Y(men_men_n117_));
  AOI210     u107(.A0(men_men_n82_), .A1(men_men_n65_), .B0(men_men_n117_), .Y(men_men_n118_));
  NO2        u108(.A(i_8_), .B(i_7_), .Y(men_men_n119_));
  OA210      u109(.A0(men_men_n118_), .A1(men_men_n116_), .B0(men_men_n119_), .Y(men_men_n120_));
  NA4        u110(.A(men_men_n89_), .B(i_0_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n121_));
  NO2        u111(.A(men_men_n121_), .B(i_4_), .Y(men_men_n122_));
  NO3        u112(.A(men_men_n122_), .B(men_men_n120_), .C(men_men_n115_), .Y(men_men_n123_));
  NO2        u113(.A(men_men_n78_), .B(men_men_n26_), .Y(men_men_n124_));
  NA3        u114(.A(men_men_n68_), .B(men_men_n89_), .C(i_0_), .Y(men_men_n125_));
  NOi31      u115(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n126_));
  OAI210     u116(.A0(men_men_n107_), .A1(men_men_n58_), .B0(men_men_n126_), .Y(men_men_n127_));
  NA2        u117(.A(men_men_n127_), .B(men_men_n125_), .Y(men_men_n128_));
  NO2        u118(.A(men_men_n128_), .B(men_men_n124_), .Y(men_men_n129_));
  NA4        u119(.A(men_men_n129_), .B(men_men_n123_), .C(men_men_n112_), .D(men_men_n100_), .Y(men_men_n130_));
  OR4        u120(.A(men_men_n130_), .B(men_men_n95_), .C(men_men_n64_), .D(men_men_n52_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule