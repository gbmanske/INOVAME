// Benchmark "top" written by ABC on Fri Jun 21 17:49:26 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n124_, new_new_n125_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n384_, new_new_n385_,
    new_new_n386_, new_new_n387_, new_new_n388_, new_new_n389_,
    new_new_n390_, new_new_n391_, new_new_n392_, new_new_n393_,
    new_new_n394_, new_new_n395_, new_new_n396_, new_new_n397_,
    new_new_n398_, new_new_n399_, new_new_n400_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n406_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n499_, new_new_n500_, new_new_n501_, new_new_n502_,
    new_new_n503_, new_new_n504_, new_new_n505_, new_new_n506_,
    new_new_n507_, new_new_n508_, new_new_n509_, new_new_n510_,
    new_new_n511_, new_new_n512_, new_new_n513_, new_new_n514_,
    new_new_n515_, new_new_n516_, new_new_n517_, new_new_n518_,
    new_new_n519_, new_new_n520_, new_new_n521_, new_new_n522_,
    new_new_n523_, new_new_n524_, new_new_n525_, new_new_n526_,
    new_new_n527_, new_new_n528_, new_new_n529_, new_new_n530_,
    new_new_n531_, new_new_n532_, new_new_n533_, new_new_n534_,
    new_new_n535_, new_new_n536_, new_new_n537_, new_new_n538_,
    new_new_n539_, new_new_n540_, new_new_n541_, new_new_n543_,
    new_new_n544_, new_new_n545_, new_new_n546_, new_new_n547_,
    new_new_n548_, new_new_n549_, new_new_n550_, new_new_n551_,
    new_new_n552_, new_new_n553_, new_new_n554_, new_new_n555_,
    new_new_n556_, new_new_n557_, new_new_n558_, new_new_n559_,
    new_new_n560_, new_new_n561_, new_new_n562_, new_new_n563_,
    new_new_n564_, new_new_n565_, new_new_n566_, new_new_n567_,
    new_new_n568_, new_new_n569_, new_new_n570_, new_new_n571_,
    new_new_n572_, new_new_n573_, new_new_n574_, new_new_n575_,
    new_new_n576_, new_new_n577_, new_new_n578_, new_new_n579_,
    new_new_n580_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n653_, new_new_n654_, new_new_n655_, new_new_n656_,
    new_new_n657_, new_new_n658_, new_new_n659_, new_new_n660_,
    new_new_n661_, new_new_n662_, new_new_n663_, new_new_n664_,
    new_new_n665_, new_new_n666_, new_new_n667_, new_new_n668_,
    new_new_n669_, new_new_n670_, new_new_n671_, new_new_n672_,
    new_new_n673_, new_new_n674_, new_new_n675_, new_new_n676_,
    new_new_n677_, new_new_n678_, new_new_n679_, new_new_n680_,
    new_new_n681_, new_new_n682_, new_new_n683_, new_new_n684_,
    new_new_n685_, new_new_n686_, new_new_n687_, new_new_n688_,
    new_new_n689_, new_new_n690_, new_new_n691_, new_new_n692_,
    new_new_n693_, new_new_n694_, new_new_n695_, new_new_n696_,
    new_new_n697_, new_new_n698_, new_new_n699_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n709_, new_new_n710_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NAi31      g018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(ori1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_5_), .A1(new_new_n46_), .B0(new_new_n45_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA2        g031(.A(new_new_n50_), .B(new_new_n44_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  NAi21      g034(.An(i_2_), .B(i_7_), .Y(new_new_n57_));
  INV        g035(.A(i_1_), .Y(new_new_n58_));
  NA2        g036(.A(new_new_n58_), .B(i_6_), .Y(new_new_n59_));
  NA3        g037(.A(new_new_n59_), .B(new_new_n57_), .C(new_new_n31_), .Y(new_new_n60_));
  INV        g038(.A(new_new_n60_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n49_), .B(i_2_), .Y(new_new_n62_));
  AOI210     g040(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(i_1_), .B(i_6_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(new_new_n25_), .Y(new_new_n65_));
  INV        g043(.A(i_0_), .Y(new_new_n66_));
  NAi21      g044(.An(i_5_), .B(i_10_), .Y(new_new_n67_));
  NA2        g045(.A(i_5_), .B(i_9_), .Y(new_new_n68_));
  AOI210     g046(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n66_), .Y(new_new_n69_));
  NO2        g047(.A(new_new_n69_), .B(new_new_n65_), .Y(new_new_n70_));
  OAI210     g048(.A0(new_new_n63_), .A1(new_new_n62_), .B0(new_new_n70_), .Y(new_new_n71_));
  OAI210     g049(.A0(new_new_n71_), .A1(new_new_n61_), .B0(i_0_), .Y(new_new_n72_));
  NA2        g050(.A(i_12_), .B(i_5_), .Y(new_new_n73_));
  NO2        g051(.A(i_3_), .B(i_7_), .Y(new_new_n74_));
  INV        g052(.A(i_6_), .Y(new_new_n75_));
  OR4        g053(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n76_));
  INV        g054(.A(new_new_n76_), .Y(new_new_n77_));
  NO2        g055(.A(i_2_), .B(i_7_), .Y(new_new_n78_));
  NO2        g056(.A(new_new_n77_), .B(new_new_n78_), .Y(new_new_n79_));
  OAI210     g057(.A0(i_1_), .A1(i_6_), .B0(new_new_n79_), .Y(new_new_n80_));
  NAi21      g058(.An(i_6_), .B(i_10_), .Y(new_new_n81_));
  NA2        g059(.A(i_6_), .B(i_9_), .Y(new_new_n82_));
  AOI210     g060(.A0(new_new_n82_), .A1(new_new_n81_), .B0(new_new_n58_), .Y(new_new_n83_));
  NA2        g061(.A(i_2_), .B(i_6_), .Y(new_new_n84_));
  INV        g062(.A(new_new_n83_), .Y(new_new_n85_));
  AOI210     g063(.A0(new_new_n85_), .A1(new_new_n80_), .B0(new_new_n73_), .Y(new_new_n86_));
  AN3        g064(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n87_));
  NAi21      g065(.An(i_6_), .B(i_11_), .Y(new_new_n88_));
  NA2        g066(.A(new_new_n87_), .B(new_new_n32_), .Y(new_new_n89_));
  INV        g067(.A(i_7_), .Y(new_new_n90_));
  NA2        g068(.A(new_new_n45_), .B(new_new_n90_), .Y(new_new_n91_));
  NO2        g069(.A(i_0_), .B(i_5_), .Y(new_new_n92_));
  NO2        g070(.A(new_new_n92_), .B(new_new_n75_), .Y(new_new_n93_));
  NA2        g071(.A(i_12_), .B(i_3_), .Y(new_new_n94_));
  INV        g072(.A(new_new_n94_), .Y(new_new_n95_));
  NAi21      g073(.An(i_7_), .B(i_11_), .Y(new_new_n96_));
  NO3        g074(.A(new_new_n96_), .B(new_new_n81_), .C(new_new_n51_), .Y(new_new_n97_));
  NO2        g075(.A(i_2_), .B(i_7_), .Y(new_new_n98_));
  OR2        g076(.A(new_new_n73_), .B(new_new_n55_), .Y(new_new_n99_));
  NA2        g077(.A(i_12_), .B(i_7_), .Y(new_new_n100_));
  NO2        g078(.A(new_new_n58_), .B(new_new_n26_), .Y(new_new_n101_));
  NA2        g079(.A(new_new_n101_), .B(i_0_), .Y(new_new_n102_));
  NA2        g080(.A(i_11_), .B(i_12_), .Y(new_new_n103_));
  OAI210     g081(.A0(new_new_n102_), .A1(new_new_n100_), .B0(new_new_n103_), .Y(new_new_n104_));
  INV        g082(.A(new_new_n104_), .Y(new_new_n105_));
  NAi31      g083(.An(new_new_n97_), .B(new_new_n105_), .C(new_new_n89_), .Y(new_new_n106_));
  NOi21      g084(.An(i_1_), .B(i_5_), .Y(new_new_n107_));
  NA2        g085(.A(new_new_n107_), .B(i_11_), .Y(new_new_n108_));
  NA2        g086(.A(new_new_n90_), .B(new_new_n37_), .Y(new_new_n109_));
  NA2        g087(.A(i_7_), .B(new_new_n25_), .Y(new_new_n110_));
  NA2        g088(.A(new_new_n110_), .B(new_new_n109_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(new_new_n45_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n82_), .B(new_new_n81_), .Y(new_new_n113_));
  NAi21      g091(.An(i_3_), .B(i_8_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n114_), .B(new_new_n57_), .Y(new_new_n115_));
  NOi31      g093(.An(new_new_n115_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n116_));
  NO2        g094(.A(i_1_), .B(new_new_n75_), .Y(new_new_n117_));
  NO2        g095(.A(i_6_), .B(i_5_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n118_), .B(i_3_), .Y(new_new_n119_));
  AO210      g097(.A0(new_new_n119_), .A1(new_new_n46_), .B0(new_new_n117_), .Y(new_new_n120_));
  OAI220     g098(.A0(new_new_n120_), .A1(new_new_n96_), .B0(new_new_n116_), .B1(new_new_n108_), .Y(new_new_n121_));
  NO3        g099(.A(new_new_n121_), .B(new_new_n106_), .C(new_new_n86_), .Y(new_new_n122_));
  NA3        g100(.A(new_new_n122_), .B(new_new_n72_), .C(new_new_n54_), .Y(ori2));
  NO2        g101(.A(new_new_n58_), .B(new_new_n37_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n707_), .B(new_new_n124_), .Y(new_new_n125_));
  NA4        g103(.A(new_new_n125_), .B(new_new_n70_), .C(new_new_n62_), .D(new_new_n30_), .Y(ori0));
  NO2        g104(.A(i_12_), .B(i_13_), .Y(new_new_n127_));
  NAi21      g105(.An(i_5_), .B(i_11_), .Y(new_new_n128_));
  NO2        g106(.A(i_0_), .B(i_1_), .Y(new_new_n129_));
  NA2        g107(.A(i_2_), .B(i_3_), .Y(new_new_n130_));
  NA2        g108(.A(i_1_), .B(i_5_), .Y(new_new_n131_));
  OR2        g109(.A(i_0_), .B(i_1_), .Y(new_new_n132_));
  NO3        g110(.A(new_new_n132_), .B(new_new_n73_), .C(i_13_), .Y(new_new_n133_));
  NAi32      g111(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n134_));
  NOi21      g112(.An(i_4_), .B(i_10_), .Y(new_new_n135_));
  NA2        g113(.A(new_new_n135_), .B(new_new_n39_), .Y(new_new_n136_));
  NOi21      g114(.An(i_4_), .B(i_9_), .Y(new_new_n137_));
  NOi21      g115(.An(i_11_), .B(i_13_), .Y(new_new_n138_));
  NA2        g116(.A(new_new_n138_), .B(new_new_n137_), .Y(new_new_n139_));
  NO2        g117(.A(i_4_), .B(i_5_), .Y(new_new_n140_));
  NAi21      g118(.An(i_12_), .B(i_11_), .Y(new_new_n141_));
  NO2        g119(.A(new_new_n141_), .B(i_13_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n66_), .B(new_new_n58_), .Y(new_new_n143_));
  NO2        g121(.A(new_new_n66_), .B(i_5_), .Y(new_new_n144_));
  NO2        g122(.A(i_13_), .B(i_10_), .Y(new_new_n145_));
  NO2        g123(.A(i_2_), .B(i_1_), .Y(new_new_n146_));
  NAi21      g124(.An(i_4_), .B(i_12_), .Y(new_new_n147_));
  INV        g125(.A(i_8_), .Y(new_new_n148_));
  NO3        g126(.A(i_3_), .B(new_new_n75_), .C(new_new_n47_), .Y(new_new_n149_));
  NA2        g127(.A(new_new_n149_), .B(i_7_), .Y(new_new_n150_));
  NO3        g128(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n151_));
  NO2        g129(.A(i_3_), .B(i_8_), .Y(new_new_n152_));
  NO3        g130(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n153_));
  NA3        g131(.A(new_new_n153_), .B(new_new_n152_), .C(new_new_n39_), .Y(new_new_n154_));
  NO2        g132(.A(new_new_n92_), .B(new_new_n55_), .Y(new_new_n155_));
  INV        g133(.A(new_new_n155_), .Y(new_new_n156_));
  NO2        g134(.A(i_13_), .B(i_9_), .Y(new_new_n157_));
  NAi21      g135(.An(i_12_), .B(i_3_), .Y(new_new_n158_));
  NO2        g136(.A(new_new_n43_), .B(i_5_), .Y(new_new_n159_));
  NO2        g137(.A(new_new_n156_), .B(new_new_n154_), .Y(new_new_n160_));
  NA2        g138(.A(new_new_n160_), .B(i_7_), .Y(new_new_n161_));
  NO2        g139(.A(new_new_n161_), .B(i_4_), .Y(new_new_n162_));
  NA3        g140(.A(i_13_), .B(new_new_n148_), .C(i_10_), .Y(new_new_n163_));
  NA2        g141(.A(i_0_), .B(i_5_), .Y(new_new_n164_));
  NAi31      g142(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n165_));
  NO2        g143(.A(new_new_n36_), .B(i_13_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n66_), .B(new_new_n26_), .Y(new_new_n167_));
  NO2        g145(.A(new_new_n45_), .B(new_new_n58_), .Y(new_new_n168_));
  INV        g146(.A(i_13_), .Y(new_new_n169_));
  NO2        g147(.A(i_12_), .B(new_new_n169_), .Y(new_new_n170_));
  NO2        g148(.A(i_12_), .B(new_new_n37_), .Y(new_new_n171_));
  OR2        g149(.A(i_8_), .B(i_7_), .Y(new_new_n172_));
  INV        g150(.A(i_12_), .Y(new_new_n173_));
  NO3        g151(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n174_));
  NA2        g152(.A(i_2_), .B(i_1_), .Y(new_new_n175_));
  NO3        g153(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n176_));
  NAi21      g154(.An(i_4_), .B(i_3_), .Y(new_new_n177_));
  NO2        g155(.A(i_0_), .B(i_6_), .Y(new_new_n178_));
  NOi41      g156(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n179_));
  NO2        g157(.A(i_11_), .B(new_new_n169_), .Y(new_new_n180_));
  NOi21      g158(.An(i_1_), .B(i_6_), .Y(new_new_n181_));
  NAi21      g159(.An(i_3_), .B(i_7_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n173_), .B(i_9_), .Y(new_new_n183_));
  OR4        g161(.A(new_new_n183_), .B(new_new_n182_), .C(new_new_n181_), .D(new_new_n144_), .Y(new_new_n184_));
  NA2        g162(.A(new_new_n66_), .B(i_5_), .Y(new_new_n185_));
  NA2        g163(.A(i_3_), .B(i_9_), .Y(new_new_n186_));
  NAi21      g164(.An(i_7_), .B(i_10_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n187_), .B(new_new_n186_), .Y(new_new_n188_));
  NA3        g166(.A(new_new_n188_), .B(new_new_n185_), .C(new_new_n59_), .Y(new_new_n189_));
  NA2        g167(.A(new_new_n189_), .B(new_new_n184_), .Y(new_new_n190_));
  NA2        g168(.A(new_new_n190_), .B(new_new_n180_), .Y(new_new_n191_));
  NO2        g169(.A(new_new_n172_), .B(new_new_n37_), .Y(new_new_n192_));
  NA2        g170(.A(i_12_), .B(i_6_), .Y(new_new_n193_));
  OR2        g171(.A(i_13_), .B(i_9_), .Y(new_new_n194_));
  NO3        g172(.A(new_new_n194_), .B(new_new_n193_), .C(new_new_n47_), .Y(new_new_n195_));
  NO2        g173(.A(new_new_n177_), .B(i_2_), .Y(new_new_n196_));
  NA3        g174(.A(new_new_n196_), .B(new_new_n195_), .C(new_new_n43_), .Y(new_new_n197_));
  NA2        g175(.A(new_new_n180_), .B(i_9_), .Y(new_new_n198_));
  OAI210     g176(.A0(new_new_n66_), .A1(new_new_n198_), .B0(new_new_n197_), .Y(new_new_n199_));
  NO3        g177(.A(i_11_), .B(new_new_n169_), .C(new_new_n25_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n182_), .B(i_8_), .Y(new_new_n201_));
  NA2        g179(.A(new_new_n199_), .B(new_new_n192_), .Y(new_new_n202_));
  NA2        g180(.A(new_new_n202_), .B(new_new_n191_), .Y(new_new_n203_));
  NO3        g181(.A(i_12_), .B(new_new_n169_), .C(new_new_n37_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n175_), .B(i_0_), .Y(new_new_n205_));
  NO2        g183(.A(i_3_), .B(i_10_), .Y(new_new_n206_));
  NO2        g184(.A(i_2_), .B(new_new_n90_), .Y(new_new_n207_));
  AN2        g185(.A(i_3_), .B(i_10_), .Y(new_new_n208_));
  NO2        g186(.A(i_5_), .B(new_new_n37_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n45_), .B(new_new_n26_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n203_), .B(new_new_n162_), .Y(new_new_n211_));
  NO3        g189(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n212_));
  NO2        g190(.A(i_2_), .B(i_3_), .Y(new_new_n213_));
  OR2        g191(.A(i_0_), .B(i_5_), .Y(new_new_n214_));
  NO2        g192(.A(i_12_), .B(i_10_), .Y(new_new_n215_));
  NOi21      g193(.An(i_5_), .B(i_0_), .Y(new_new_n216_));
  NO2        g194(.A(i_2_), .B(new_new_n90_), .Y(new_new_n217_));
  NO4        g195(.A(new_new_n217_), .B(i_4_), .C(new_new_n216_), .D(new_new_n114_), .Y(new_new_n218_));
  NA2        g196(.A(new_new_n218_), .B(new_new_n215_), .Y(new_new_n219_));
  INV        g197(.A(i_6_), .Y(new_new_n220_));
  NO2        g198(.A(i_1_), .B(i_7_), .Y(new_new_n221_));
  INV        g199(.A(new_new_n219_), .Y(new_new_n222_));
  NOi21      g200(.An(new_new_n131_), .B(new_new_n93_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n223_), .B(new_new_n110_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n224_), .B(i_3_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n148_), .B(i_9_), .Y(new_new_n226_));
  NA2        g204(.A(new_new_n226_), .B(new_new_n155_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n45_), .Y(new_new_n228_));
  INV        g206(.A(new_new_n228_), .Y(new_new_n229_));
  AOI210     g207(.A0(new_new_n229_), .A1(new_new_n225_), .B0(new_new_n136_), .Y(new_new_n230_));
  AOI210     g208(.A0(new_new_n222_), .A1(new_new_n212_), .B0(new_new_n230_), .Y(new_new_n231_));
  NOi32      g209(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n232_));
  INV        g210(.A(new_new_n232_), .Y(new_new_n233_));
  NAi21      g211(.An(i_0_), .B(i_6_), .Y(new_new_n234_));
  NAi21      g212(.An(i_1_), .B(i_5_), .Y(new_new_n235_));
  NA2        g213(.A(new_new_n235_), .B(new_new_n234_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n236_), .B(new_new_n25_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n237_), .B(new_new_n134_), .Y(new_new_n238_));
  NAi41      g216(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n239_));
  OAI220     g217(.A0(new_new_n239_), .A1(new_new_n235_), .B0(new_new_n165_), .B1(new_new_n134_), .Y(new_new_n240_));
  AOI210     g218(.A0(new_new_n239_), .A1(new_new_n134_), .B0(new_new_n132_), .Y(new_new_n241_));
  NOi32      g219(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n242_));
  NAi21      g220(.An(i_6_), .B(i_1_), .Y(new_new_n243_));
  NA3        g221(.A(new_new_n243_), .B(new_new_n242_), .C(new_new_n45_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n244_), .B(i_0_), .Y(new_new_n245_));
  OR3        g223(.A(new_new_n245_), .B(new_new_n241_), .C(new_new_n240_), .Y(new_new_n246_));
  NAi21      g224(.An(i_3_), .B(i_4_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n247_), .B(i_9_), .Y(new_new_n248_));
  AN2        g226(.A(i_6_), .B(i_7_), .Y(new_new_n249_));
  NA2        g227(.A(i_2_), .B(i_7_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n247_), .B(i_10_), .Y(new_new_n251_));
  AOI210     g229(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n252_));
  OAI210     g230(.A0(new_new_n252_), .A1(new_new_n146_), .B0(new_new_n251_), .Y(new_new_n253_));
  AOI220     g231(.A0(new_new_n251_), .A1(new_new_n221_), .B0(new_new_n174_), .B1(new_new_n146_), .Y(new_new_n254_));
  AOI210     g232(.A0(new_new_n254_), .A1(new_new_n253_), .B0(i_5_), .Y(new_new_n255_));
  NO3        g233(.A(new_new_n255_), .B(new_new_n246_), .C(new_new_n238_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n256_), .B(new_new_n233_), .Y(new_new_n257_));
  AN2        g235(.A(i_12_), .B(i_5_), .Y(new_new_n258_));
  NA2        g236(.A(i_3_), .B(new_new_n258_), .Y(new_new_n259_));
  NO2        g237(.A(i_11_), .B(i_6_), .Y(new_new_n260_));
  NO2        g238(.A(i_5_), .B(i_10_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n262_));
  NA4        g240(.A(new_new_n206_), .B(new_new_n82_), .C(new_new_n68_), .D(new_new_n52_), .Y(new_new_n263_));
  NO2        g241(.A(i_11_), .B(i_12_), .Y(new_new_n264_));
  NA2        g242(.A(new_new_n264_), .B(new_new_n36_), .Y(new_new_n265_));
  NO2        g243(.A(new_new_n263_), .B(new_new_n265_), .Y(new_new_n266_));
  NAi21      g244(.An(i_13_), .B(i_0_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n267_), .B(new_new_n175_), .Y(new_new_n268_));
  NA2        g246(.A(new_new_n266_), .B(new_new_n268_), .Y(new_new_n269_));
  NO2        g247(.A(i_0_), .B(i_11_), .Y(new_new_n270_));
  NOi21      g248(.An(i_2_), .B(i_12_), .Y(new_new_n271_));
  NAi21      g249(.An(i_9_), .B(i_4_), .Y(new_new_n272_));
  OR2        g250(.A(i_13_), .B(i_10_), .Y(new_new_n273_));
  NO3        g251(.A(new_new_n273_), .B(new_new_n103_), .C(new_new_n272_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n139_), .B(new_new_n109_), .Y(new_new_n275_));
  NO2        g253(.A(new_new_n90_), .B(new_new_n25_), .Y(new_new_n276_));
  NA2        g254(.A(new_new_n204_), .B(new_new_n276_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n277_), .B(new_new_n223_), .Y(new_new_n278_));
  NA2        g256(.A(new_new_n148_), .B(i_10_), .Y(new_new_n279_));
  NA3        g257(.A(new_new_n185_), .B(new_new_n59_), .C(i_2_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(new_new_n279_), .Y(new_new_n281_));
  INV        g259(.A(new_new_n281_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n282_), .B(new_new_n198_), .Y(new_new_n283_));
  NO4        g261(.A(new_new_n283_), .B(new_new_n278_), .C(new_new_n708_), .D(new_new_n257_), .Y(new_new_n284_));
  NO2        g262(.A(new_new_n66_), .B(i_13_), .Y(new_new_n285_));
  NO2        g263(.A(i_10_), .B(i_9_), .Y(new_new_n286_));
  NAi21      g264(.An(i_12_), .B(i_8_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n287_), .B(i_3_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n45_), .B(i_4_), .Y(new_new_n289_));
  NA2        g267(.A(new_new_n289_), .B(new_new_n93_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n290_), .B(new_new_n154_), .Y(new_new_n291_));
  NA2        g269(.A(new_new_n210_), .B(i_0_), .Y(new_new_n292_));
  NO3        g270(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n293_));
  NA2        g271(.A(new_new_n193_), .B(new_new_n88_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n294_), .B(new_new_n293_), .Y(new_new_n295_));
  NA2        g273(.A(i_8_), .B(i_9_), .Y(new_new_n296_));
  NO2        g274(.A(i_7_), .B(i_2_), .Y(new_new_n297_));
  OR2        g275(.A(new_new_n297_), .B(new_new_n296_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n204_), .B(new_new_n155_), .Y(new_new_n299_));
  OAI220     g277(.A0(new_new_n299_), .A1(new_new_n298_), .B0(new_new_n295_), .B1(new_new_n292_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n180_), .B(new_new_n209_), .Y(new_new_n301_));
  NO3        g279(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n302_));
  INV        g280(.A(new_new_n302_), .Y(new_new_n303_));
  NA3        g281(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n304_));
  NA4        g282(.A(new_new_n128_), .B(new_new_n101_), .C(new_new_n73_), .D(new_new_n23_), .Y(new_new_n305_));
  OAI220     g283(.A0(new_new_n305_), .A1(new_new_n304_), .B0(new_new_n303_), .B1(new_new_n301_), .Y(new_new_n306_));
  NO3        g284(.A(new_new_n306_), .B(new_new_n300_), .C(new_new_n291_), .Y(new_new_n307_));
  OR2        g285(.A(new_new_n227_), .B(new_new_n90_), .Y(new_new_n308_));
  OR2        g286(.A(new_new_n308_), .B(new_new_n136_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n87_), .B(i_13_), .Y(new_new_n310_));
  NO2        g288(.A(i_2_), .B(i_13_), .Y(new_new_n311_));
  NO3        g289(.A(i_4_), .B(new_new_n47_), .C(i_8_), .Y(new_new_n312_));
  NO2        g290(.A(i_6_), .B(i_7_), .Y(new_new_n313_));
  NO2        g291(.A(i_11_), .B(i_1_), .Y(new_new_n314_));
  NOi21      g292(.An(i_2_), .B(i_7_), .Y(new_new_n315_));
  NO2        g293(.A(i_3_), .B(new_new_n148_), .Y(new_new_n316_));
  NO2        g294(.A(i_6_), .B(i_10_), .Y(new_new_n317_));
  NA3        g295(.A(new_new_n179_), .B(new_new_n138_), .C(new_new_n118_), .Y(new_new_n318_));
  NA2        g296(.A(new_new_n45_), .B(new_new_n43_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n132_), .B(i_3_), .Y(new_new_n320_));
  NAi31      g298(.An(new_new_n319_), .B(new_new_n320_), .C(new_new_n170_), .Y(new_new_n321_));
  NA2        g299(.A(new_new_n293_), .B(new_new_n258_), .Y(new_new_n322_));
  NAi21      g300(.An(new_new_n163_), .B(new_new_n264_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n221_), .B(new_new_n164_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n324_), .B(new_new_n323_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n27_), .B(i_10_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n212_), .B(new_new_n174_), .Y(new_new_n327_));
  OAI220     g305(.A0(new_new_n327_), .A1(new_new_n280_), .B0(new_new_n326_), .B1(new_new_n310_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n328_), .B(new_new_n325_), .Y(new_new_n329_));
  NA4        g307(.A(new_new_n329_), .B(new_new_n321_), .C(new_new_n309_), .D(new_new_n307_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n108_), .B(new_new_n99_), .Y(new_new_n331_));
  AN2        g309(.A(new_new_n331_), .B(new_new_n293_), .Y(new_new_n332_));
  NA2        g310(.A(new_new_n332_), .B(new_new_n210_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n258_), .B(new_new_n169_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n232_), .B(new_new_n66_), .Y(new_new_n335_));
  NA2        g313(.A(new_new_n249_), .B(new_new_n242_), .Y(new_new_n336_));
  OR2        g314(.A(new_new_n334_), .B(new_new_n336_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n36_), .B(i_8_), .Y(new_new_n338_));
  INV        g316(.A(new_new_n274_), .Y(new_new_n339_));
  NA2        g317(.A(new_new_n339_), .B(new_new_n337_), .Y(new_new_n340_));
  INV        g318(.A(new_new_n340_), .Y(new_new_n341_));
  INV        g319(.A(new_new_n185_), .Y(new_new_n342_));
  OAI210     g320(.A0(i_8_), .A1(new_new_n342_), .B0(new_new_n120_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n343_), .B(new_new_n275_), .Y(new_new_n344_));
  NA3        g322(.A(new_new_n344_), .B(new_new_n341_), .C(new_new_n333_), .Y(new_new_n345_));
  NO2        g323(.A(i_12_), .B(new_new_n148_), .Y(new_new_n346_));
  NO2        g324(.A(i_8_), .B(i_7_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n43_), .B(i_10_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(i_6_), .Y(new_new_n349_));
  NA3        g327(.A(new_new_n208_), .B(new_new_n140_), .C(new_new_n87_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n132_), .B(i_5_), .Y(new_new_n351_));
  INV        g329(.A(new_new_n350_), .Y(new_new_n352_));
  NA2        g330(.A(new_new_n352_), .B(new_new_n302_), .Y(new_new_n353_));
  INV        g331(.A(new_new_n353_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n355_));
  NA2        g333(.A(new_new_n286_), .B(new_new_n166_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n355_), .B(new_new_n356_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n45_), .B(i_7_), .Y(new_new_n358_));
  NA2        g336(.A(i_0_), .B(new_new_n47_), .Y(new_new_n359_));
  NA3        g337(.A(new_new_n346_), .B(new_new_n200_), .C(new_new_n359_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n358_), .B(new_new_n360_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n361_), .B(new_new_n357_), .Y(new_new_n362_));
  NO4        g340(.A(new_new_n181_), .B(new_new_n41_), .C(i_2_), .D(new_new_n47_), .Y(new_new_n363_));
  NO3        g341(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n364_));
  NOi21      g342(.An(i_10_), .B(i_6_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n75_), .B(new_new_n25_), .Y(new_new_n366_));
  AOI220     g344(.A0(new_new_n204_), .A1(new_new_n366_), .B0(new_new_n200_), .B1(new_new_n365_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(new_new_n292_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n100_), .B(new_new_n23_), .Y(new_new_n369_));
  INV        g347(.A(new_new_n368_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n335_), .B(new_new_n254_), .Y(new_new_n371_));
  INV        g349(.A(new_new_n213_), .Y(new_new_n372_));
  NO2        g350(.A(i_12_), .B(new_new_n75_), .Y(new_new_n373_));
  NA2        g351(.A(new_new_n373_), .B(new_new_n200_), .Y(new_new_n374_));
  NA3        g352(.A(new_new_n260_), .B(new_new_n204_), .C(new_new_n164_), .Y(new_new_n375_));
  AOI210     g353(.A0(new_new_n375_), .A1(new_new_n374_), .B0(new_new_n372_), .Y(new_new_n376_));
  OR2        g354(.A(i_2_), .B(i_5_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n250_), .B(new_new_n178_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n378_), .B(new_new_n323_), .Y(new_new_n379_));
  NO3        g357(.A(new_new_n379_), .B(new_new_n376_), .C(new_new_n371_), .Y(new_new_n380_));
  NA3        g358(.A(new_new_n380_), .B(new_new_n370_), .C(new_new_n362_), .Y(new_new_n381_));
  NO4        g359(.A(new_new_n381_), .B(new_new_n354_), .C(new_new_n345_), .D(new_new_n330_), .Y(new_new_n382_));
  NA4        g360(.A(new_new_n382_), .B(new_new_n284_), .C(new_new_n231_), .D(new_new_n211_), .Y(ori7));
  NO2        g361(.A(new_new_n84_), .B(new_new_n52_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n96_), .B(new_new_n81_), .Y(new_new_n385_));
  NA2        g363(.A(i_3_), .B(new_new_n385_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n317_), .B(new_new_n74_), .Y(new_new_n387_));
  NA2        g365(.A(i_11_), .B(new_new_n148_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n127_), .B(new_new_n388_), .Y(new_new_n389_));
  OAI210     g367(.A0(new_new_n389_), .A1(new_new_n387_), .B0(new_new_n386_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n173_), .B(i_4_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n391_), .B(i_8_), .Y(new_new_n392_));
  NA2        g370(.A(i_2_), .B(new_new_n75_), .Y(new_new_n393_));
  OAI210     g371(.A0(new_new_n78_), .A1(new_new_n152_), .B0(new_new_n153_), .Y(new_new_n394_));
  NO2        g372(.A(i_7_), .B(new_new_n37_), .Y(new_new_n395_));
  NA2        g373(.A(i_4_), .B(i_8_), .Y(new_new_n396_));
  NO2        g374(.A(new_new_n394_), .B(i_13_), .Y(new_new_n397_));
  NO3        g375(.A(new_new_n397_), .B(new_new_n390_), .C(new_new_n384_), .Y(new_new_n398_));
  AOI210     g376(.A0(new_new_n114_), .A1(new_new_n57_), .B0(i_10_), .Y(new_new_n399_));
  AOI210     g377(.A0(new_new_n399_), .A1(new_new_n173_), .B0(new_new_n135_), .Y(new_new_n400_));
  OR2        g378(.A(i_6_), .B(i_10_), .Y(new_new_n401_));
  INV        g379(.A(new_new_n151_), .Y(new_new_n402_));
  OR2        g380(.A(new_new_n400_), .B(new_new_n194_), .Y(new_new_n403_));
  AOI210     g381(.A0(new_new_n403_), .A1(new_new_n398_), .B0(new_new_n58_), .Y(new_new_n404_));
  NOi21      g382(.An(i_11_), .B(i_7_), .Y(new_new_n405_));
  AO210      g383(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n406_), .B(new_new_n405_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n407_), .B(new_new_n157_), .Y(new_new_n408_));
  NA3        g386(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n409_));
  NAi31      g387(.An(new_new_n409_), .B(i_12_), .C(i_11_), .Y(new_new_n410_));
  AOI210     g388(.A0(new_new_n410_), .A1(new_new_n408_), .B0(new_new_n58_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n77_), .B(new_new_n58_), .Y(new_new_n412_));
  AO210      g390(.A0(new_new_n412_), .A1(new_new_n254_), .B0(new_new_n40_), .Y(new_new_n413_));
  NO3        g391(.A(new_new_n187_), .B(new_new_n158_), .C(new_new_n388_), .Y(new_new_n414_));
  OAI210     g392(.A0(new_new_n414_), .A1(new_new_n170_), .B0(new_new_n58_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n271_), .B(new_new_n31_), .Y(new_new_n416_));
  OR2        g394(.A(new_new_n158_), .B(new_new_n96_), .Y(new_new_n417_));
  NA2        g395(.A(new_new_n417_), .B(new_new_n416_), .Y(new_new_n418_));
  NO2        g396(.A(i_1_), .B(i_4_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n419_), .B(new_new_n418_), .Y(new_new_n420_));
  NO2        g398(.A(i_1_), .B(i_12_), .Y(new_new_n421_));
  NA3        g399(.A(new_new_n421_), .B(i_2_), .C(new_new_n24_), .Y(new_new_n422_));
  BUFFER     g400(.A(new_new_n422_), .Y(new_new_n423_));
  NA4        g401(.A(new_new_n423_), .B(new_new_n420_), .C(new_new_n415_), .D(new_new_n413_), .Y(new_new_n424_));
  OAI210     g402(.A0(new_new_n424_), .A1(new_new_n411_), .B0(i_6_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n409_), .B(new_new_n96_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n426_), .B(new_new_n373_), .Y(new_new_n427_));
  NO2        g405(.A(i_6_), .B(i_11_), .Y(new_new_n428_));
  NA2        g406(.A(new_new_n427_), .B(new_new_n295_), .Y(new_new_n429_));
  NO3        g407(.A(new_new_n401_), .B(new_new_n172_), .C(new_new_n23_), .Y(new_new_n430_));
  AOI210     g408(.A0(i_1_), .A1(new_new_n188_), .B0(new_new_n430_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n431_), .B(new_new_n43_), .Y(new_new_n432_));
  NA3        g410(.A(new_new_n347_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n433_));
  INV        g411(.A(i_2_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n124_), .B(i_9_), .Y(new_new_n435_));
  NA3        g413(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n45_), .B(i_1_), .Y(new_new_n437_));
  NA3        g415(.A(new_new_n437_), .B(new_new_n193_), .C(new_new_n43_), .Y(new_new_n438_));
  OAI220     g416(.A0(new_new_n438_), .A1(new_new_n436_), .B0(new_new_n435_), .B1(new_new_n434_), .Y(new_new_n439_));
  AOI210     g417(.A0(new_new_n314_), .A1(new_new_n276_), .B0(new_new_n176_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n440_), .B(new_new_n393_), .Y(new_new_n441_));
  NAi21      g419(.An(new_new_n433_), .B(new_new_n83_), .Y(new_new_n442_));
  INV        g420(.A(new_new_n442_), .Y(new_new_n443_));
  OR3        g421(.A(new_new_n443_), .B(new_new_n441_), .C(new_new_n439_), .Y(new_new_n444_));
  NO3        g422(.A(new_new_n444_), .B(new_new_n432_), .C(new_new_n429_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n173_), .B(new_new_n90_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n446_), .B(new_new_n405_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n709_), .B(new_new_n100_), .Y(new_new_n448_));
  AN2        g426(.A(new_new_n448_), .B(new_new_n349_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n450_));
  NA2        g428(.A(i_1_), .B(i_3_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n296_), .B(new_new_n84_), .Y(new_new_n452_));
  INV        g430(.A(new_new_n452_), .Y(new_new_n453_));
  NO2        g431(.A(new_new_n453_), .B(new_new_n451_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n454_), .B(new_new_n449_), .Y(new_new_n455_));
  NA3        g433(.A(new_new_n455_), .B(new_new_n445_), .C(new_new_n425_), .Y(new_new_n456_));
  NA2        g434(.A(new_new_n249_), .B(new_new_n248_), .Y(new_new_n457_));
  NO3        g435(.A(new_new_n315_), .B(new_new_n396_), .C(new_new_n75_), .Y(new_new_n458_));
  NA2        g436(.A(new_new_n458_), .B(new_new_n25_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n459_), .B(new_new_n457_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n460_), .B(i_1_), .Y(new_new_n461_));
  AOI210     g439(.A0(new_new_n193_), .A1(new_new_n88_), .B0(i_1_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n247_), .B(i_2_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n463_), .B(new_new_n462_), .Y(new_new_n464_));
  AOI210     g442(.A0(new_new_n464_), .A1(new_new_n461_), .B0(i_13_), .Y(new_new_n465_));
  OR2        g443(.A(i_11_), .B(i_7_), .Y(new_new_n466_));
  NA3        g444(.A(new_new_n466_), .B(new_new_n95_), .C(new_new_n124_), .Y(new_new_n467_));
  AOI220     g445(.A0(new_new_n311_), .A1(new_new_n135_), .B0(new_new_n289_), .B1(new_new_n124_), .Y(new_new_n468_));
  OAI210     g446(.A0(new_new_n468_), .A1(new_new_n43_), .B0(new_new_n467_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n469_), .B(new_new_n220_), .Y(new_new_n470_));
  INV        g448(.A(new_new_n100_), .Y(new_new_n471_));
  AOI220     g449(.A0(new_new_n471_), .A1(new_new_n65_), .B0(new_new_n260_), .B1(new_new_n437_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n177_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n113_), .B(i_13_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n436_), .B(new_new_n100_), .Y(new_new_n475_));
  INV        g453(.A(new_new_n475_), .Y(new_new_n476_));
  OAI220     g454(.A0(new_new_n476_), .A1(new_new_n64_), .B0(new_new_n474_), .B1(new_new_n462_), .Y(new_new_n477_));
  NO3        g455(.A(new_new_n64_), .B(new_new_n32_), .C(new_new_n90_), .Y(new_new_n478_));
  NA2        g456(.A(i_3_), .B(i_7_), .Y(new_new_n479_));
  NO3        g457(.A(new_new_n315_), .B(new_new_n173_), .C(new_new_n75_), .Y(new_new_n480_));
  AOI210     g458(.A0(new_new_n480_), .A1(new_new_n479_), .B0(new_new_n478_), .Y(new_new_n481_));
  AOI220     g459(.A0(new_new_n260_), .A1(new_new_n437_), .B0(new_new_n83_), .B1(new_new_n91_), .Y(new_new_n482_));
  OAI220     g460(.A0(new_new_n482_), .A1(new_new_n392_), .B0(new_new_n481_), .B1(new_new_n402_), .Y(new_new_n483_));
  NO3        g461(.A(new_new_n483_), .B(new_new_n477_), .C(new_new_n473_), .Y(new_new_n484_));
  OR2        g462(.A(i_11_), .B(i_6_), .Y(new_new_n485_));
  NO2        g463(.A(new_new_n476_), .B(new_new_n485_), .Y(new_new_n486_));
  NA3        g464(.A(new_new_n271_), .B(new_new_n395_), .C(new_new_n88_), .Y(new_new_n487_));
  NA2        g465(.A(new_new_n428_), .B(i_13_), .Y(new_new_n488_));
  NAi21      g466(.An(i_11_), .B(i_12_), .Y(new_new_n489_));
  NO3        g467(.A(new_new_n315_), .B(new_new_n373_), .C(new_new_n396_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n490_), .B(new_new_n212_), .Y(new_new_n491_));
  NA3        g469(.A(new_new_n491_), .B(new_new_n488_), .C(new_new_n487_), .Y(new_new_n492_));
  OAI210     g470(.A0(new_new_n492_), .A1(new_new_n486_), .B0(new_new_n58_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n710_), .B(new_new_n421_), .Y(new_new_n494_));
  INV        g472(.A(new_new_n494_), .Y(new_new_n495_));
  NA3        g473(.A(new_new_n495_), .B(new_new_n44_), .C(new_new_n169_), .Y(new_new_n496_));
  NA4        g474(.A(new_new_n496_), .B(new_new_n493_), .C(new_new_n484_), .D(new_new_n470_), .Y(new_new_n497_));
  OR4        g475(.A(new_new_n497_), .B(new_new_n465_), .C(new_new_n456_), .D(new_new_n404_), .Y(ori5));
  NA2        g476(.A(new_new_n447_), .B(new_new_n196_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n392_), .B(i_11_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n78_), .B(new_new_n500_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n501_), .B(new_new_n499_), .Y(new_new_n502_));
  NO3        g480(.A(i_11_), .B(new_new_n173_), .C(i_13_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n110_), .B(new_new_n23_), .Y(new_new_n504_));
  INV        g482(.A(new_new_n286_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n213_), .B(new_new_n369_), .Y(new_new_n506_));
  INV        g484(.A(new_new_n506_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(new_new_n502_), .Y(new_new_n508_));
  INV        g486(.A(new_new_n138_), .Y(new_new_n509_));
  INV        g487(.A(new_new_n179_), .Y(new_new_n510_));
  OAI210     g488(.A0(new_new_n463_), .A1(new_new_n288_), .B0(new_new_n98_), .Y(new_new_n511_));
  AOI210     g489(.A0(new_new_n511_), .A1(new_new_n510_), .B0(new_new_n509_), .Y(new_new_n512_));
  NO2        g490(.A(new_new_n296_), .B(new_new_n26_), .Y(new_new_n513_));
  NO2        g491(.A(new_new_n513_), .B(new_new_n276_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n514_), .B(i_2_), .Y(new_new_n515_));
  INV        g493(.A(new_new_n515_), .Y(new_new_n516_));
  AOI210     g494(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n273_), .Y(new_new_n517_));
  AOI210     g495(.A0(new_new_n517_), .A1(new_new_n516_), .B0(new_new_n512_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n147_), .B(new_new_n111_), .Y(new_new_n519_));
  OAI210     g497(.A0(new_new_n519_), .A1(new_new_n504_), .B0(i_2_), .Y(new_new_n520_));
  INV        g498(.A(new_new_n139_), .Y(new_new_n521_));
  NO3        g499(.A(new_new_n406_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n522_));
  AOI210     g500(.A0(new_new_n521_), .A1(new_new_n78_), .B0(new_new_n522_), .Y(new_new_n523_));
  AOI210     g501(.A0(new_new_n523_), .A1(new_new_n520_), .B0(new_new_n148_), .Y(new_new_n524_));
  OA210      g502(.A0(new_new_n407_), .A1(new_new_n112_), .B0(i_13_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n151_), .B(new_new_n152_), .Y(new_new_n526_));
  NO2        g504(.A(new_new_n526_), .B(new_new_n250_), .Y(new_new_n527_));
  AOI210     g505(.A0(new_new_n158_), .A1(new_new_n130_), .B0(new_new_n338_), .Y(new_new_n528_));
  NA2        g506(.A(new_new_n528_), .B(new_new_n276_), .Y(new_new_n529_));
  NO2        g507(.A(new_new_n91_), .B(new_new_n43_), .Y(new_new_n530_));
  INV        g508(.A(new_new_n207_), .Y(new_new_n531_));
  NA4        g509(.A(new_new_n531_), .B(new_new_n208_), .C(new_new_n110_), .D(new_new_n41_), .Y(new_new_n532_));
  OAI210     g510(.A0(new_new_n532_), .A1(new_new_n530_), .B0(new_new_n529_), .Y(new_new_n533_));
  NO4        g511(.A(new_new_n533_), .B(new_new_n527_), .C(new_new_n525_), .D(new_new_n524_), .Y(new_new_n534_));
  NA2        g512(.A(new_new_n369_), .B(new_new_n28_), .Y(new_new_n535_));
  NA2        g513(.A(new_new_n503_), .B(new_new_n201_), .Y(new_new_n536_));
  NA2        g514(.A(new_new_n536_), .B(new_new_n535_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n57_), .B(i_12_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n538_), .B(new_new_n112_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n539_), .B(new_new_n388_), .Y(new_new_n540_));
  AOI220     g518(.A0(new_new_n540_), .A1(new_new_n36_), .B0(new_new_n537_), .B1(new_new_n45_), .Y(new_new_n541_));
  NA4        g519(.A(new_new_n541_), .B(new_new_n534_), .C(new_new_n518_), .D(new_new_n508_), .Y(ori6));
  NA4        g520(.A(new_new_n261_), .B(new_new_n316_), .C(new_new_n64_), .D(new_new_n90_), .Y(new_new_n543_));
  INV        g521(.A(new_new_n543_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n165_), .B(new_new_n319_), .Y(new_new_n545_));
  NO2        g523(.A(i_11_), .B(i_9_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n544_), .B(new_new_n216_), .Y(new_new_n547_));
  OR2        g525(.A(new_new_n547_), .B(i_12_), .Y(new_new_n548_));
  NA2        g526(.A(new_new_n373_), .B(new_new_n58_), .Y(new_new_n549_));
  BUFFER     g527(.A(new_new_n412_), .Y(new_new_n550_));
  NA2        g528(.A(new_new_n550_), .B(new_new_n549_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n150_), .Y(new_new_n552_));
  AOI220     g530(.A0(new_new_n552_), .A1(new_new_n546_), .B0(new_new_n551_), .B1(new_new_n66_), .Y(new_new_n553_));
  INV        g531(.A(new_new_n215_), .Y(new_new_n554_));
  NA2        g532(.A(new_new_n68_), .B(new_new_n117_), .Y(new_new_n555_));
  INV        g533(.A(new_new_n110_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n556_), .B(new_new_n45_), .Y(new_new_n557_));
  AOI210     g535(.A0(new_new_n557_), .A1(new_new_n555_), .B0(new_new_n554_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n181_), .B(i_9_), .Y(new_new_n559_));
  NA2        g537(.A(new_new_n559_), .B(new_new_n538_), .Y(new_new_n560_));
  AOI210     g538(.A0(new_new_n560_), .A1(new_new_n336_), .B0(new_new_n144_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n32_), .B(i_11_), .Y(new_new_n562_));
  NAi32      g540(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n563_));
  NO2        g541(.A(new_new_n485_), .B(new_new_n563_), .Y(new_new_n564_));
  OR3        g542(.A(new_new_n564_), .B(new_new_n561_), .C(new_new_n558_), .Y(new_new_n565_));
  NO2        g543(.A(new_new_n466_), .B(i_2_), .Y(new_new_n566_));
  NA3        g544(.A(new_new_n288_), .B(new_new_n129_), .C(new_new_n62_), .Y(new_new_n567_));
  OR2        g545(.A(new_new_n505_), .B(new_new_n36_), .Y(new_new_n568_));
  NA2        g546(.A(new_new_n568_), .B(new_new_n567_), .Y(new_new_n569_));
  OAI210     g547(.A0(i_6_), .A1(i_11_), .B0(new_new_n76_), .Y(new_new_n570_));
  AOI220     g548(.A0(new_new_n570_), .A1(new_new_n364_), .B0(new_new_n545_), .B1(new_new_n479_), .Y(new_new_n571_));
  NA3        g549(.A(new_new_n250_), .B(new_new_n174_), .C(new_new_n129_), .Y(new_new_n572_));
  NA3        g550(.A(new_new_n572_), .B(new_new_n571_), .C(new_new_n394_), .Y(new_new_n573_));
  AO210      g551(.A0(new_new_n338_), .A1(new_new_n45_), .B0(new_new_n77_), .Y(new_new_n574_));
  NA3        g552(.A(new_new_n574_), .B(new_new_n317_), .C(new_new_n164_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n288_), .B(new_new_n286_), .Y(new_new_n576_));
  NO2        g554(.A(new_new_n401_), .B(new_new_n91_), .Y(new_new_n577_));
  OAI210     g555(.A0(new_new_n577_), .A1(new_new_n99_), .B0(new_new_n270_), .Y(new_new_n578_));
  NA3        g556(.A(new_new_n578_), .B(new_new_n576_), .C(new_new_n575_), .Y(new_new_n579_));
  NO4        g557(.A(new_new_n579_), .B(new_new_n573_), .C(new_new_n569_), .D(new_new_n565_), .Y(new_new_n580_));
  NA4        g558(.A(new_new_n580_), .B(new_new_n553_), .C(new_new_n548_), .D(new_new_n256_), .Y(ori3));
  NA2        g559(.A(i_12_), .B(i_10_), .Y(new_new_n582_));
  NA2        g560(.A(new_new_n572_), .B(new_new_n394_), .Y(new_new_n583_));
  NA2        g561(.A(new_new_n583_), .B(new_new_n39_), .Y(new_new_n584_));
  NOi21      g562(.An(new_new_n87_), .B(new_new_n514_), .Y(new_new_n585_));
  NO3        g563(.A(new_new_n417_), .B(new_new_n296_), .C(new_new_n117_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n271_), .B(new_new_n44_), .Y(new_new_n587_));
  AN2        g565(.A(new_new_n294_), .B(new_new_n53_), .Y(new_new_n588_));
  NO3        g566(.A(new_new_n588_), .B(new_new_n586_), .C(new_new_n585_), .Y(new_new_n589_));
  AOI210     g567(.A0(new_new_n589_), .A1(new_new_n584_), .B0(new_new_n47_), .Y(new_new_n590_));
  NO3        g568(.A(new_new_n258_), .B(new_new_n38_), .C(i_0_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n144_), .B(new_new_n365_), .Y(new_new_n592_));
  NOi21      g570(.An(new_new_n592_), .B(new_new_n591_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n593_), .B(new_new_n58_), .Y(new_new_n594_));
  NOi21      g572(.An(i_5_), .B(i_9_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n595_), .B(new_new_n285_), .Y(new_new_n596_));
  BUFFER     g574(.A(new_new_n193_), .Y(new_new_n597_));
  AOI210     g575(.A0(new_new_n597_), .A1(new_new_n314_), .B0(new_new_n458_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n598_), .B(new_new_n596_), .Y(new_new_n599_));
  NO3        g577(.A(new_new_n599_), .B(new_new_n594_), .C(new_new_n590_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n144_), .B(new_new_n24_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n450_), .B(new_new_n385_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n602_), .B(new_new_n601_), .Y(new_new_n603_));
  INV        g581(.A(new_new_n603_), .Y(new_new_n604_));
  NA2        g582(.A(new_new_n366_), .B(i_0_), .Y(new_new_n605_));
  NO3        g583(.A(new_new_n605_), .B(new_new_n259_), .C(new_new_n78_), .Y(new_new_n606_));
  NO4        g584(.A(new_new_n377_), .B(i_12_), .C(new_new_n273_), .D(i_6_), .Y(new_new_n607_));
  AOI210     g585(.A0(new_new_n607_), .A1(i_11_), .B0(new_new_n606_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n503_), .B(new_new_n216_), .Y(new_new_n609_));
  AOI210     g587(.A0(new_new_n317_), .A1(new_new_n78_), .B0(new_new_n55_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n610_), .B(new_new_n609_), .Y(new_new_n611_));
  NO2        g589(.A(new_new_n183_), .B(new_new_n131_), .Y(new_new_n612_));
  INV        g590(.A(new_new_n348_), .Y(new_new_n613_));
  NO4        g591(.A(new_new_n100_), .B(new_new_n55_), .C(new_new_n709_), .D(i_5_), .Y(new_new_n614_));
  AO220      g592(.A0(new_new_n614_), .A1(new_new_n613_), .B0(new_new_n612_), .B1(i_6_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n615_), .B(new_new_n611_), .Y(new_new_n616_));
  NA3        g594(.A(new_new_n616_), .B(new_new_n608_), .C(new_new_n604_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n92_), .B(new_new_n37_), .Y(new_new_n618_));
  NA2        g596(.A(i_11_), .B(i_9_), .Y(new_new_n619_));
  NO3        g597(.A(i_12_), .B(new_new_n619_), .C(new_new_n393_), .Y(new_new_n620_));
  AN2        g598(.A(new_new_n620_), .B(new_new_n618_), .Y(new_new_n621_));
  NA2        g599(.A(new_new_n262_), .B(new_new_n143_), .Y(new_new_n622_));
  INV        g600(.A(new_new_n622_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n619_), .B(new_new_n66_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n623_), .B(new_new_n621_), .Y(new_new_n625_));
  NA2        g603(.A(new_new_n138_), .B(new_new_n92_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n395_), .B(new_new_n216_), .Y(new_new_n627_));
  NO2        g605(.A(new_new_n627_), .B(new_new_n587_), .Y(new_new_n628_));
  INV        g606(.A(new_new_n628_), .Y(new_new_n629_));
  INV        g607(.A(new_new_n214_), .Y(new_new_n630_));
  NA2        g608(.A(new_new_n629_), .B(new_new_n625_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n582_), .B(new_new_n213_), .Y(new_new_n632_));
  OA210      g610(.A0(new_new_n313_), .A1(new_new_n168_), .B0(new_new_n312_), .Y(new_new_n633_));
  NA2        g611(.A(new_new_n632_), .B(new_new_n624_), .Y(new_new_n634_));
  NA2        g612(.A(new_new_n624_), .B(new_new_n208_), .Y(new_new_n635_));
  INV        g613(.A(new_new_n635_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n636_), .B(new_new_n313_), .Y(new_new_n637_));
  NO3        g615(.A(new_new_n377_), .B(new_new_n234_), .C(new_new_n24_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n351_), .B(new_new_n638_), .Y(new_new_n639_));
  NAi21      g617(.An(i_9_), .B(i_5_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n640_), .B(new_new_n267_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n641_), .B(new_new_n407_), .Y(new_new_n642_));
  OAI220     g620(.A0(new_new_n642_), .A1(new_new_n75_), .B0(new_new_n639_), .B1(new_new_n139_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n643_), .B(new_new_n340_), .Y(new_new_n644_));
  NA3        g622(.A(new_new_n644_), .B(new_new_n637_), .C(new_new_n634_), .Y(new_new_n645_));
  NO3        g623(.A(new_new_n645_), .B(new_new_n631_), .C(new_new_n617_), .Y(new_new_n646_));
  NO2        g624(.A(i_0_), .B(new_new_n489_), .Y(new_new_n647_));
  AOI210     g625(.A0(new_new_n549_), .A1(new_new_n457_), .B0(new_new_n626_), .Y(new_new_n648_));
  INV        g626(.A(new_new_n648_), .Y(new_new_n649_));
  NA2        g627(.A(new_new_n178_), .B(new_new_n171_), .Y(new_new_n650_));
  AOI210     g628(.A0(new_new_n650_), .A1(new_new_n605_), .B0(new_new_n131_), .Y(new_new_n651_));
  INV        g629(.A(new_new_n651_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n652_), .B(new_new_n649_), .Y(new_new_n653_));
  NO3        g631(.A(new_new_n159_), .B(new_new_n258_), .C(i_0_), .Y(new_new_n654_));
  OAI210     g632(.A0(new_new_n654_), .A1(new_new_n69_), .B0(i_13_), .Y(new_new_n655_));
  INV        g633(.A(new_new_n655_), .Y(new_new_n656_));
  INV        g634(.A(new_new_n84_), .Y(new_new_n657_));
  AOI210     g635(.A0(new_new_n657_), .A1(new_new_n647_), .B0(new_new_n97_), .Y(new_new_n658_));
  OR2        g636(.A(new_new_n658_), .B(i_5_), .Y(new_new_n659_));
  AOI210     g637(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n141_), .Y(new_new_n660_));
  NA2        g638(.A(new_new_n660_), .B(new_new_n633_), .Y(new_new_n661_));
  NO3        g639(.A(new_new_n587_), .B(new_new_n52_), .C(new_new_n47_), .Y(new_new_n662_));
  NA2        g640(.A(new_new_n322_), .B(new_new_n318_), .Y(new_new_n663_));
  NO3        g641(.A(new_new_n663_), .B(new_new_n662_), .C(new_new_n706_), .Y(new_new_n664_));
  NA3        g642(.A(new_new_n261_), .B(new_new_n138_), .C(new_new_n137_), .Y(new_new_n665_));
  NA3        g643(.A(i_5_), .B(new_new_n205_), .C(new_new_n171_), .Y(new_new_n666_));
  NA2        g644(.A(new_new_n666_), .B(new_new_n665_), .Y(new_new_n667_));
  NO3        g645(.A(new_new_n619_), .B(new_new_n164_), .C(new_new_n147_), .Y(new_new_n668_));
  NO2        g646(.A(new_new_n668_), .B(new_new_n667_), .Y(new_new_n669_));
  NA4        g647(.A(new_new_n669_), .B(new_new_n664_), .C(new_new_n661_), .D(new_new_n659_), .Y(new_new_n670_));
  BUFFER     g648(.A(new_new_n176_), .Y(new_new_n671_));
  NO3        g649(.A(new_new_n175_), .B(i_0_), .C(i_12_), .Y(new_new_n672_));
  AOI220     g650(.A0(new_new_n672_), .A1(new_new_n671_), .B0(new_new_n544_), .B1(new_new_n142_), .Y(new_new_n673_));
  INV        g651(.A(new_new_n673_), .Y(new_new_n674_));
  NO4        g652(.A(new_new_n674_), .B(new_new_n670_), .C(new_new_n656_), .D(new_new_n653_), .Y(new_new_n675_));
  OAI210     g653(.A0(new_new_n566_), .A1(new_new_n562_), .B0(new_new_n37_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n676_), .B(new_new_n400_), .Y(new_new_n677_));
  NA2        g655(.A(new_new_n677_), .B(new_new_n157_), .Y(new_new_n678_));
  BUFFER     g656(.A(new_new_n466_), .Y(new_new_n679_));
  NA2        g657(.A(new_new_n145_), .B(new_new_n146_), .Y(new_new_n680_));
  AO210      g658(.A0(new_new_n679_), .A1(new_new_n33_), .B0(new_new_n680_), .Y(new_new_n681_));
  NAi31      g659(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n682_));
  NO2        g660(.A(new_new_n63_), .B(new_new_n682_), .Y(new_new_n683_));
  NO2        g661(.A(new_new_n683_), .B(new_new_n430_), .Y(new_new_n684_));
  NA2        g662(.A(new_new_n684_), .B(new_new_n681_), .Y(new_new_n685_));
  NO2        g663(.A(new_new_n304_), .B(new_new_n193_), .Y(new_new_n686_));
  AOI210     g664(.A0(new_new_n685_), .A1(new_new_n47_), .B0(new_new_n686_), .Y(new_new_n687_));
  AOI210     g665(.A0(new_new_n687_), .A1(new_new_n678_), .B0(new_new_n66_), .Y(new_new_n688_));
  INV        g666(.A(new_new_n255_), .Y(new_new_n689_));
  NO2        g667(.A(new_new_n689_), .B(new_new_n509_), .Y(new_new_n690_));
  OAI210     g668(.A0(new_new_n195_), .A1(new_new_n133_), .B0(new_new_n78_), .Y(new_new_n691_));
  NO2        g669(.A(new_new_n691_), .B(i_11_), .Y(new_new_n692_));
  NO3        g670(.A(new_new_n56_), .B(new_new_n55_), .C(i_4_), .Y(new_new_n693_));
  OAI210     g671(.A0(new_new_n630_), .A1(new_new_n209_), .B0(new_new_n693_), .Y(new_new_n694_));
  NO2        g672(.A(new_new_n694_), .B(new_new_n489_), .Y(new_new_n695_));
  NO4        g673(.A(new_new_n640_), .B(i_11_), .C(new_new_n182_), .D(new_new_n181_), .Y(new_new_n696_));
  NO2        g674(.A(new_new_n696_), .B(new_new_n363_), .Y(new_new_n697_));
  INV        g675(.A(new_new_n240_), .Y(new_new_n698_));
  AOI210     g676(.A0(new_new_n698_), .A1(new_new_n697_), .B0(new_new_n40_), .Y(new_new_n699_));
  NO3        g677(.A(new_new_n699_), .B(new_new_n695_), .C(new_new_n692_), .Y(new_new_n700_));
  INV        g678(.A(new_new_n700_), .Y(new_new_n701_));
  NO3        g679(.A(new_new_n701_), .B(new_new_n690_), .C(new_new_n688_), .Y(new_new_n702_));
  NA4        g680(.A(new_new_n702_), .B(new_new_n675_), .C(new_new_n646_), .D(new_new_n600_), .Y(ori4));
  INV        g681(.A(new_new_n350_), .Y(new_new_n706_));
  INV        g682(.A(i_6_), .Y(new_new_n707_));
  INV        g683(.A(new_new_n269_), .Y(new_new_n708_));
  INV        g684(.A(i_3_), .Y(new_new_n709_));
  INV        g685(.A(i_2_), .Y(new_new_n710_));
endmodule


