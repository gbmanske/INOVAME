//Benchmark atmr_alu4_1266_0.0156

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n142_, ori_ori_n143_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n894_, ori_ori_n895_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  OAI210     o033(.A0(ori_ori_n55_), .A1(ori_ori_n52_), .B0(ori_ori_n45_), .Y(ori_ori_n56_));
  NA3        o034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(ori_ori_n57_));
  NO2        o035(.A(i_1_), .B(i_6_), .Y(ori_ori_n58_));
  NA2        o036(.A(i_8_), .B(i_7_), .Y(ori_ori_n59_));
  OAI210     o037(.A0(ori_ori_n59_), .A1(ori_ori_n58_), .B0(ori_ori_n57_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(i_12_), .Y(ori_ori_n61_));
  NAi21      o039(.An(i_2_), .B(i_7_), .Y(ori_ori_n62_));
  INV        o040(.A(i_1_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n63_), .B(i_6_), .Y(ori_ori_n64_));
  NA3        o042(.A(ori_ori_n64_), .B(ori_ori_n62_), .C(ori_ori_n31_), .Y(ori_ori_n65_));
  NA2        o043(.A(i_1_), .B(i_10_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n66_), .B(i_6_), .Y(ori_ori_n67_));
  NAi31      o045(.An(ori_ori_n67_), .B(ori_ori_n65_), .C(ori_ori_n61_), .Y(ori_ori_n68_));
  NA2        o046(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_1_), .B(i_6_), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n71_), .B(ori_ori_n25_), .Y(ori_ori_n72_));
  INV        o050(.A(i_0_), .Y(ori_ori_n73_));
  NAi21      o051(.An(i_5_), .B(i_10_), .Y(ori_ori_n74_));
  NA2        o052(.A(i_5_), .B(i_9_), .Y(ori_ori_n75_));
  AOI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n73_), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n70_), .A1(ori_ori_n69_), .B0(ori_ori_n77_), .Y(ori_ori_n78_));
  OAI210     o056(.A0(ori_ori_n78_), .A1(ori_ori_n68_), .B0(i_0_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_12_), .B(i_5_), .Y(ori_ori_n80_));
  NA2        o058(.A(i_2_), .B(i_8_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n81_), .B(ori_ori_n58_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_3_), .B(i_9_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_3_), .B(i_7_), .Y(ori_ori_n84_));
  NO3        o062(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(ori_ori_n63_), .Y(ori_ori_n85_));
  INV        o063(.A(i_6_), .Y(ori_ori_n86_));
  OR4        o064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  NO2        o066(.A(i_2_), .B(i_7_), .Y(ori_ori_n89_));
  AOI210     o067(.A0(ori_ori_n88_), .A1(ori_ori_n86_), .B0(ori_ori_n89_), .Y(ori_ori_n90_));
  OAI210     o068(.A0(ori_ori_n85_), .A1(ori_ori_n82_), .B0(ori_ori_n90_), .Y(ori_ori_n91_));
  NAi21      o069(.An(i_6_), .B(i_10_), .Y(ori_ori_n92_));
  NA2        o070(.A(i_6_), .B(i_9_), .Y(ori_ori_n93_));
  AOI210     o071(.A0(ori_ori_n93_), .A1(ori_ori_n92_), .B0(ori_ori_n63_), .Y(ori_ori_n94_));
  NA2        o072(.A(i_2_), .B(i_6_), .Y(ori_ori_n95_));
  NO3        o073(.A(ori_ori_n95_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n96_));
  NO2        o074(.A(ori_ori_n96_), .B(ori_ori_n94_), .Y(ori_ori_n97_));
  AOI210     o075(.A0(ori_ori_n97_), .A1(ori_ori_n91_), .B0(ori_ori_n80_), .Y(ori_ori_n98_));
  AN3        o076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n99_));
  NAi21      o077(.An(i_6_), .B(i_11_), .Y(ori_ori_n100_));
  NO2        o078(.A(i_5_), .B(i_8_), .Y(ori_ori_n101_));
  NOi21      o079(.An(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  AOI220     o080(.A0(ori_ori_n102_), .A1(ori_ori_n62_), .B0(ori_ori_n99_), .B1(ori_ori_n32_), .Y(ori_ori_n103_));
  INV        o081(.A(i_7_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n46_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  NO2        o083(.A(i_0_), .B(i_5_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(ori_ori_n86_), .Y(ori_ori_n107_));
  NA2        o085(.A(i_12_), .B(i_3_), .Y(ori_ori_n108_));
  INV        o086(.A(ori_ori_n108_), .Y(ori_ori_n109_));
  NA3        o087(.A(ori_ori_n109_), .B(ori_ori_n107_), .C(ori_ori_n105_), .Y(ori_ori_n110_));
  NAi21      o088(.An(i_7_), .B(i_11_), .Y(ori_ori_n111_));
  NO3        o089(.A(ori_ori_n111_), .B(ori_ori_n92_), .C(ori_ori_n53_), .Y(ori_ori_n112_));
  AN2        o090(.A(i_2_), .B(i_10_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n113_), .B(i_7_), .Y(ori_ori_n114_));
  OR2        o092(.A(ori_ori_n80_), .B(ori_ori_n58_), .Y(ori_ori_n115_));
  NO2        o093(.A(i_8_), .B(ori_ori_n104_), .Y(ori_ori_n116_));
  NO3        o094(.A(ori_ori_n116_), .B(ori_ori_n115_), .C(ori_ori_n114_), .Y(ori_ori_n117_));
  NA2        o095(.A(i_12_), .B(i_7_), .Y(ori_ori_n118_));
  NO2        o096(.A(ori_ori_n63_), .B(ori_ori_n26_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(i_0_), .Y(ori_ori_n120_));
  NA2        o098(.A(i_11_), .B(i_12_), .Y(ori_ori_n121_));
  OAI210     o099(.A0(ori_ori_n120_), .A1(ori_ori_n118_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n122_), .B(ori_ori_n117_), .Y(ori_ori_n123_));
  NAi41      o101(.An(ori_ori_n112_), .B(ori_ori_n123_), .C(ori_ori_n110_), .D(ori_ori_n103_), .Y(ori_ori_n124_));
  NOi21      o102(.An(i_1_), .B(i_5_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n125_), .B(i_11_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n104_), .B(ori_ori_n37_), .Y(ori_ori_n127_));
  NA2        o105(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n127_), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n129_), .B(ori_ori_n46_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n93_), .B(ori_ori_n92_), .Y(ori_ori_n131_));
  NAi21      o109(.An(i_3_), .B(i_8_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n132_), .B(ori_ori_n62_), .Y(ori_ori_n133_));
  NOi31      o111(.An(ori_ori_n133_), .B(ori_ori_n131_), .C(ori_ori_n130_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_1_), .B(ori_ori_n86_), .Y(ori_ori_n135_));
  NO2        o113(.A(i_6_), .B(i_5_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n136_), .B(i_3_), .Y(ori_ori_n137_));
  AO210      o115(.A0(ori_ori_n137_), .A1(ori_ori_n47_), .B0(ori_ori_n135_), .Y(ori_ori_n138_));
  OAI220     o116(.A0(ori_ori_n138_), .A1(ori_ori_n111_), .B0(ori_ori_n134_), .B1(ori_ori_n126_), .Y(ori_ori_n139_));
  NO3        o117(.A(ori_ori_n139_), .B(ori_ori_n124_), .C(ori_ori_n98_), .Y(ori_ori_n140_));
  NA3        o118(.A(ori_ori_n140_), .B(ori_ori_n79_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o119(.A(ori_ori_n63_), .B(ori_ori_n37_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n895_), .B(ori_ori_n142_), .Y(ori_ori_n143_));
  NA4        o121(.A(ori_ori_n143_), .B(ori_ori_n77_), .C(ori_ori_n69_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o122(.A(i_8_), .B(i_7_), .Y(ori_ori_n145_));
  NA2        o123(.A(ori_ori_n145_), .B(i_6_), .Y(ori_ori_n146_));
  NO2        o124(.A(i_12_), .B(i_13_), .Y(ori_ori_n147_));
  NAi21      o125(.An(i_5_), .B(i_11_), .Y(ori_ori_n148_));
  NOi21      o126(.An(ori_ori_n147_), .B(ori_ori_n148_), .Y(ori_ori_n149_));
  NO2        o127(.A(i_0_), .B(i_1_), .Y(ori_ori_n150_));
  NA2        o128(.A(i_2_), .B(i_3_), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n151_), .B(i_4_), .Y(ori_ori_n152_));
  NA3        o130(.A(ori_ori_n152_), .B(ori_ori_n150_), .C(ori_ori_n149_), .Y(ori_ori_n153_));
  AN2        o131(.A(ori_ori_n147_), .B(ori_ori_n83_), .Y(ori_ori_n154_));
  NA2        o132(.A(i_1_), .B(i_5_), .Y(ori_ori_n155_));
  OR2        o133(.A(i_0_), .B(i_1_), .Y(ori_ori_n156_));
  NO3        o134(.A(ori_ori_n156_), .B(ori_ori_n80_), .C(i_13_), .Y(ori_ori_n157_));
  NAi32      o135(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n158_));
  NAi21      o136(.An(ori_ori_n158_), .B(ori_ori_n157_), .Y(ori_ori_n159_));
  NOi21      o137(.An(i_4_), .B(i_10_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(ori_ori_n40_), .Y(ori_ori_n161_));
  NO3        o139(.A(ori_ori_n73_), .B(i_2_), .C(i_1_), .Y(ori_ori_n162_));
  NO2        o140(.A(ori_ori_n159_), .B(ori_ori_n146_), .Y(ori_ori_n163_));
  NOi21      o141(.An(i_4_), .B(i_9_), .Y(ori_ori_n164_));
  NOi21      o142(.An(i_11_), .B(i_13_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n165_), .B(ori_ori_n164_), .Y(ori_ori_n166_));
  NO2        o144(.A(i_4_), .B(i_5_), .Y(ori_ori_n167_));
  NAi21      o145(.An(i_12_), .B(i_11_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n168_), .B(i_13_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n73_), .B(ori_ori_n63_), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n170_), .B(ori_ori_n46_), .Y(ori_ori_n171_));
  NA2        o149(.A(i_3_), .B(i_5_), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n173_));
  NO2        o151(.A(i_13_), .B(i_10_), .Y(ori_ori_n174_));
  NA3        o152(.A(ori_ori_n174_), .B(ori_ori_n173_), .C(ori_ori_n44_), .Y(ori_ori_n175_));
  NO2        o153(.A(i_2_), .B(i_1_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(i_3_), .Y(ori_ori_n177_));
  NAi21      o155(.An(i_4_), .B(i_12_), .Y(ori_ori_n178_));
  INV        o156(.A(i_8_), .Y(ori_ori_n179_));
  NO3        o157(.A(i_3_), .B(ori_ori_n86_), .C(ori_ori_n48_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n180_), .B(ori_ori_n116_), .Y(ori_ori_n181_));
  NO3        o159(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n182_));
  NO3        o160(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n183_));
  NA2        o161(.A(i_12_), .B(ori_ori_n183_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n184_), .B(ori_ori_n181_), .Y(ori_ori_n185_));
  NO2        o163(.A(i_3_), .B(i_8_), .Y(ori_ori_n186_));
  NO3        o164(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n187_));
  NA3        o165(.A(ori_ori_n187_), .B(ori_ori_n186_), .C(ori_ori_n40_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n106_), .B(ori_ori_n58_), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n189_), .B(ori_ori_n156_), .Y(ori_ori_n190_));
  NO2        o168(.A(i_13_), .B(i_9_), .Y(ori_ori_n191_));
  NAi21      o169(.An(i_12_), .B(i_3_), .Y(ori_ori_n192_));
  NO2        o170(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n190_), .B(ori_ori_n188_), .Y(ori_ori_n194_));
  AOI210     o172(.A0(ori_ori_n194_), .A1(i_7_), .B0(ori_ori_n185_), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n195_), .B(i_4_), .Y(ori_ori_n196_));
  NAi21      o174(.An(i_12_), .B(i_7_), .Y(ori_ori_n197_));
  NA3        o175(.A(i_13_), .B(ori_ori_n179_), .C(i_10_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n198_), .B(ori_ori_n197_), .Y(ori_ori_n199_));
  NA2        o177(.A(i_0_), .B(i_5_), .Y(ori_ori_n200_));
  NA2        o178(.A(ori_ori_n200_), .B(ori_ori_n107_), .Y(ori_ori_n201_));
  OAI220     o179(.A0(ori_ori_n201_), .A1(ori_ori_n177_), .B0(ori_ori_n171_), .B1(ori_ori_n137_), .Y(ori_ori_n202_));
  NAi31      o180(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n73_), .B(ori_ori_n26_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n46_), .B(ori_ori_n63_), .Y(ori_ori_n206_));
  INV        o184(.A(i_13_), .Y(ori_ori_n207_));
  NO2        o185(.A(i_12_), .B(ori_ori_n207_), .Y(ori_ori_n208_));
  NA3        o186(.A(ori_ori_n208_), .B(ori_ori_n182_), .C(ori_ori_n180_), .Y(ori_ori_n209_));
  INV        o187(.A(ori_ori_n209_), .Y(ori_ori_n210_));
  AOI220     o188(.A0(ori_ori_n210_), .A1(ori_ori_n145_), .B0(ori_ori_n202_), .B1(ori_ori_n199_), .Y(ori_ori_n211_));
  NO2        o189(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n212_));
  OR2        o190(.A(i_8_), .B(i_7_), .Y(ori_ori_n213_));
  INV        o191(.A(i_12_), .Y(ori_ori_n214_));
  NO2        o192(.A(ori_ori_n44_), .B(ori_ori_n214_), .Y(ori_ori_n215_));
  NO3        o193(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n216_));
  NA2        o194(.A(i_2_), .B(i_1_), .Y(ori_ori_n217_));
  NO3        o195(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n218_));
  NAi21      o196(.An(i_4_), .B(i_3_), .Y(ori_ori_n219_));
  NO2        o197(.A(i_0_), .B(i_6_), .Y(ori_ori_n220_));
  NOi41      o198(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n221_));
  NA2        o199(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n217_), .B(ori_ori_n172_), .Y(ori_ori_n223_));
  NO2        o201(.A(i_11_), .B(ori_ori_n207_), .Y(ori_ori_n224_));
  NOi21      o202(.An(i_1_), .B(i_6_), .Y(ori_ori_n225_));
  NAi21      o203(.An(i_3_), .B(i_7_), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n214_), .B(i_9_), .Y(ori_ori_n227_));
  OR4        o205(.A(ori_ori_n227_), .B(ori_ori_n226_), .C(ori_ori_n225_), .D(ori_ori_n173_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n229_));
  NA2        o207(.A(i_3_), .B(i_9_), .Y(ori_ori_n230_));
  NAi21      o208(.An(i_7_), .B(i_10_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NA3        o210(.A(ori_ori_n232_), .B(ori_ori_n229_), .C(ori_ori_n64_), .Y(ori_ori_n233_));
  NA2        o211(.A(ori_ori_n233_), .B(ori_ori_n228_), .Y(ori_ori_n234_));
  INV        o212(.A(ori_ori_n146_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n214_), .B(i_13_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(ori_ori_n75_), .Y(ori_ori_n237_));
  AOI220     o215(.A0(ori_ori_n237_), .A1(ori_ori_n235_), .B0(ori_ori_n234_), .B1(ori_ori_n224_), .Y(ori_ori_n238_));
  NO2        o216(.A(ori_ori_n213_), .B(ori_ori_n37_), .Y(ori_ori_n239_));
  NA2        o217(.A(i_12_), .B(i_6_), .Y(ori_ori_n240_));
  OR2        o218(.A(i_13_), .B(i_9_), .Y(ori_ori_n241_));
  NO3        o219(.A(ori_ori_n241_), .B(ori_ori_n240_), .C(ori_ori_n48_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n219_), .B(i_2_), .Y(ori_ori_n243_));
  NA3        o221(.A(ori_ori_n243_), .B(ori_ori_n242_), .C(ori_ori_n44_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n224_), .B(i_9_), .Y(ori_ori_n245_));
  NA3        o223(.A(ori_ori_n229_), .B(ori_ori_n156_), .C(ori_ori_n64_), .Y(ori_ori_n246_));
  OAI210     o224(.A0(ori_ori_n246_), .A1(ori_ori_n245_), .B0(ori_ori_n244_), .Y(ori_ori_n247_));
  NO3        o225(.A(i_11_), .B(ori_ori_n207_), .C(ori_ori_n25_), .Y(ori_ori_n248_));
  NO2        o226(.A(ori_ori_n226_), .B(i_8_), .Y(ori_ori_n249_));
  NA2        o227(.A(ori_ori_n247_), .B(ori_ori_n239_), .Y(ori_ori_n250_));
  NA3        o228(.A(ori_ori_n250_), .B(ori_ori_n238_), .C(ori_ori_n211_), .Y(ori_ori_n251_));
  NO3        o229(.A(i_12_), .B(ori_ori_n207_), .C(ori_ori_n37_), .Y(ori_ori_n252_));
  NO2        o230(.A(ori_ori_n217_), .B(i_0_), .Y(ori_ori_n253_));
  NO2        o231(.A(i_2_), .B(ori_ori_n104_), .Y(ori_ori_n254_));
  AN2        o232(.A(i_3_), .B(i_10_), .Y(ori_ori_n255_));
  NO2        o233(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n256_));
  NO2        o234(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n257_));
  NO3        o235(.A(ori_ori_n251_), .B(ori_ori_n196_), .C(ori_ori_n163_), .Y(ori_ori_n258_));
  NO3        o236(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n259_));
  NO2        o237(.A(i_2_), .B(i_3_), .Y(ori_ori_n260_));
  OR2        o238(.A(i_0_), .B(i_5_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n156_), .B(ori_ori_n46_), .Y(ori_ori_n262_));
  NO2        o240(.A(i_12_), .B(i_10_), .Y(ori_ori_n263_));
  NOi21      o241(.An(i_5_), .B(i_0_), .Y(ori_ori_n264_));
  NA4        o242(.A(ori_ori_n84_), .B(ori_ori_n36_), .C(ori_ori_n86_), .D(i_8_), .Y(ori_ori_n265_));
  NO2        o243(.A(i_6_), .B(i_8_), .Y(ori_ori_n266_));
  NO2        o244(.A(i_1_), .B(i_7_), .Y(ori_ori_n267_));
  NOi21      o245(.An(ori_ori_n155_), .B(ori_ori_n107_), .Y(ori_ori_n268_));
  NO2        o246(.A(ori_ori_n268_), .B(ori_ori_n128_), .Y(ori_ori_n269_));
  NA2        o247(.A(ori_ori_n269_), .B(i_3_), .Y(ori_ori_n270_));
  NO2        o248(.A(ori_ori_n179_), .B(i_9_), .Y(ori_ori_n271_));
  NA3        o249(.A(ori_ori_n271_), .B(ori_ori_n189_), .C(ori_ori_n156_), .Y(ori_ori_n272_));
  NO2        o250(.A(ori_ori_n272_), .B(ori_ori_n46_), .Y(ori_ori_n273_));
  INV        o251(.A(ori_ori_n273_), .Y(ori_ori_n274_));
  AOI210     o252(.A0(ori_ori_n274_), .A1(ori_ori_n270_), .B0(ori_ori_n161_), .Y(ori_ori_n275_));
  INV        o253(.A(ori_ori_n275_), .Y(ori_ori_n276_));
  NOi32      o254(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n277_));
  INV        o255(.A(ori_ori_n277_), .Y(ori_ori_n278_));
  NAi21      o256(.An(i_0_), .B(i_6_), .Y(ori_ori_n279_));
  NAi21      o257(.An(i_1_), .B(i_5_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n280_), .B(ori_ori_n279_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n281_), .B(ori_ori_n25_), .Y(ori_ori_n282_));
  OAI210     o260(.A0(ori_ori_n282_), .A1(ori_ori_n158_), .B0(ori_ori_n222_), .Y(ori_ori_n283_));
  NAi41      o261(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n284_));
  OAI220     o262(.A0(ori_ori_n284_), .A1(ori_ori_n280_), .B0(ori_ori_n203_), .B1(ori_ori_n158_), .Y(ori_ori_n285_));
  AOI210     o263(.A0(ori_ori_n284_), .A1(ori_ori_n158_), .B0(ori_ori_n156_), .Y(ori_ori_n286_));
  NOi32      o264(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n287_));
  NAi21      o265(.An(i_6_), .B(i_1_), .Y(ori_ori_n288_));
  NA3        o266(.A(ori_ori_n288_), .B(ori_ori_n287_), .C(ori_ori_n46_), .Y(ori_ori_n289_));
  NO2        o267(.A(ori_ori_n289_), .B(i_0_), .Y(ori_ori_n290_));
  OR3        o268(.A(ori_ori_n290_), .B(ori_ori_n286_), .C(ori_ori_n285_), .Y(ori_ori_n291_));
  NO2        o269(.A(i_1_), .B(ori_ori_n104_), .Y(ori_ori_n292_));
  NAi21      o270(.An(i_3_), .B(i_4_), .Y(ori_ori_n293_));
  NO2        o271(.A(ori_ori_n293_), .B(i_9_), .Y(ori_ori_n294_));
  AN2        o272(.A(i_6_), .B(i_7_), .Y(ori_ori_n295_));
  OAI210     o273(.A0(ori_ori_n295_), .A1(ori_ori_n292_), .B0(ori_ori_n294_), .Y(ori_ori_n296_));
  NA2        o274(.A(i_2_), .B(i_7_), .Y(ori_ori_n297_));
  NO2        o275(.A(ori_ori_n293_), .B(i_10_), .Y(ori_ori_n298_));
  NA3        o276(.A(ori_ori_n298_), .B(ori_ori_n297_), .C(ori_ori_n220_), .Y(ori_ori_n299_));
  AOI210     o277(.A0(ori_ori_n299_), .A1(ori_ori_n296_), .B0(ori_ori_n173_), .Y(ori_ori_n300_));
  AOI210     o278(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n301_));
  OAI210     o279(.A0(ori_ori_n301_), .A1(ori_ori_n176_), .B0(ori_ori_n298_), .Y(ori_ori_n302_));
  AOI220     o280(.A0(ori_ori_n298_), .A1(ori_ori_n267_), .B0(ori_ori_n216_), .B1(ori_ori_n176_), .Y(ori_ori_n303_));
  AOI210     o281(.A0(ori_ori_n303_), .A1(ori_ori_n302_), .B0(i_5_), .Y(ori_ori_n304_));
  NO4        o282(.A(ori_ori_n304_), .B(ori_ori_n300_), .C(ori_ori_n291_), .D(ori_ori_n283_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n305_), .B(ori_ori_n278_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n59_), .B(ori_ori_n25_), .Y(ori_ori_n307_));
  AN2        o285(.A(i_12_), .B(i_5_), .Y(ori_ori_n308_));
  NO2        o286(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n309_));
  NA2        o287(.A(ori_ori_n309_), .B(ori_ori_n308_), .Y(ori_ori_n310_));
  NO2        o288(.A(i_11_), .B(i_6_), .Y(ori_ori_n311_));
  NA3        o289(.A(ori_ori_n311_), .B(ori_ori_n262_), .C(ori_ori_n207_), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n312_), .B(ori_ori_n310_), .Y(ori_ori_n313_));
  NO2        o291(.A(i_5_), .B(i_10_), .Y(ori_ori_n314_));
  NO2        o292(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n315_));
  NO2        o293(.A(ori_ori_n153_), .B(ori_ori_n86_), .Y(ori_ori_n316_));
  OAI210     o294(.A0(ori_ori_n316_), .A1(ori_ori_n313_), .B0(ori_ori_n315_), .Y(ori_ori_n317_));
  NO3        o295(.A(ori_ori_n86_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n318_));
  NO2        o296(.A(i_11_), .B(i_12_), .Y(ori_ori_n319_));
  NAi21      o297(.An(i_13_), .B(i_0_), .Y(ori_ori_n320_));
  INV        o298(.A(ori_ori_n317_), .Y(ori_ori_n321_));
  NA2        o299(.A(ori_ori_n44_), .B(ori_ori_n207_), .Y(ori_ori_n322_));
  NO3        o300(.A(i_1_), .B(i_12_), .C(ori_ori_n86_), .Y(ori_ori_n323_));
  NO2        o301(.A(i_0_), .B(i_11_), .Y(ori_ori_n324_));
  AN2        o302(.A(i_1_), .B(i_6_), .Y(ori_ori_n325_));
  NOi21      o303(.An(i_2_), .B(i_12_), .Y(ori_ori_n326_));
  NAi21      o304(.An(i_9_), .B(i_4_), .Y(ori_ori_n327_));
  OR2        o305(.A(i_13_), .B(i_10_), .Y(ori_ori_n328_));
  NO3        o306(.A(ori_ori_n328_), .B(ori_ori_n121_), .C(ori_ori_n327_), .Y(ori_ori_n329_));
  NO2        o307(.A(ori_ori_n166_), .B(ori_ori_n127_), .Y(ori_ori_n330_));
  NO2        o308(.A(ori_ori_n104_), .B(ori_ori_n25_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n252_), .B(ori_ori_n331_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n332_), .B(ori_ori_n268_), .Y(ori_ori_n333_));
  INV        o311(.A(ori_ori_n333_), .Y(ori_ori_n334_));
  NO2        o312(.A(ori_ori_n334_), .B(ori_ori_n26_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n172_), .B(ori_ori_n86_), .Y(ori_ori_n336_));
  NA2        o314(.A(ori_ori_n179_), .B(i_10_), .Y(ori_ori_n337_));
  NA3        o315(.A(ori_ori_n229_), .B(ori_ori_n64_), .C(i_2_), .Y(ori_ori_n338_));
  NO2        o316(.A(ori_ori_n338_), .B(ori_ori_n337_), .Y(ori_ori_n339_));
  NO2        o317(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n340_));
  INV        o318(.A(ori_ori_n339_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n341_), .B(ori_ori_n245_), .Y(ori_ori_n342_));
  NO4        o320(.A(ori_ori_n342_), .B(ori_ori_n335_), .C(ori_ori_n321_), .D(ori_ori_n306_), .Y(ori_ori_n343_));
  NO2        o321(.A(ori_ori_n63_), .B(i_4_), .Y(ori_ori_n344_));
  NO2        o322(.A(ori_ori_n73_), .B(i_13_), .Y(ori_ori_n345_));
  NA3        o323(.A(ori_ori_n345_), .B(ori_ori_n344_), .C(i_2_), .Y(ori_ori_n346_));
  NO2        o324(.A(i_10_), .B(i_9_), .Y(ori_ori_n347_));
  NAi21      o325(.An(i_12_), .B(i_8_), .Y(ori_ori_n348_));
  NO2        o326(.A(ori_ori_n348_), .B(i_3_), .Y(ori_ori_n349_));
  NA2        o327(.A(ori_ori_n349_), .B(ori_ori_n347_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n351_));
  NA2        o329(.A(ori_ori_n351_), .B(ori_ori_n107_), .Y(ori_ori_n352_));
  OAI220     o330(.A0(ori_ori_n352_), .A1(ori_ori_n188_), .B0(ori_ori_n350_), .B1(ori_ori_n346_), .Y(ori_ori_n353_));
  NA2        o331(.A(ori_ori_n257_), .B(i_0_), .Y(ori_ori_n354_));
  NO3        o332(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n355_));
  NA2        o333(.A(ori_ori_n240_), .B(ori_ori_n100_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n356_), .B(ori_ori_n355_), .Y(ori_ori_n357_));
  NA2        o335(.A(i_8_), .B(i_9_), .Y(ori_ori_n358_));
  AOI210     o336(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n359_));
  OR2        o337(.A(ori_ori_n359_), .B(ori_ori_n358_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n252_), .B(ori_ori_n189_), .Y(ori_ori_n361_));
  OAI220     o339(.A0(ori_ori_n361_), .A1(ori_ori_n360_), .B0(ori_ori_n357_), .B1(ori_ori_n354_), .Y(ori_ori_n362_));
  NA2        o340(.A(ori_ori_n224_), .B(ori_ori_n256_), .Y(ori_ori_n363_));
  NO3        o341(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n364_));
  INV        o342(.A(ori_ori_n364_), .Y(ori_ori_n365_));
  NA3        o343(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n366_));
  NA4        o344(.A(ori_ori_n148_), .B(ori_ori_n119_), .C(ori_ori_n80_), .D(ori_ori_n23_), .Y(ori_ori_n367_));
  OAI220     o345(.A0(ori_ori_n367_), .A1(ori_ori_n366_), .B0(ori_ori_n365_), .B1(ori_ori_n363_), .Y(ori_ori_n368_));
  NO3        o346(.A(ori_ori_n368_), .B(ori_ori_n362_), .C(ori_ori_n353_), .Y(ori_ori_n369_));
  OR2        o347(.A(ori_ori_n272_), .B(ori_ori_n104_), .Y(ori_ori_n370_));
  OR2        o348(.A(ori_ori_n370_), .B(ori_ori_n161_), .Y(ori_ori_n371_));
  NA2        o349(.A(ori_ori_n99_), .B(i_13_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n336_), .B(ori_ori_n307_), .Y(ori_ori_n373_));
  NO2        o351(.A(i_2_), .B(i_13_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n373_), .B(ori_ori_n372_), .Y(ori_ori_n375_));
  NO3        o353(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n376_));
  NO2        o354(.A(i_6_), .B(i_7_), .Y(ori_ori_n377_));
  NO2        o355(.A(i_11_), .B(i_1_), .Y(ori_ori_n378_));
  OR2        o356(.A(i_11_), .B(i_8_), .Y(ori_ori_n379_));
  NOi21      o357(.An(i_2_), .B(i_7_), .Y(ori_ori_n380_));
  NO2        o358(.A(i_3_), .B(ori_ori_n179_), .Y(ori_ori_n381_));
  NO2        o359(.A(i_6_), .B(i_10_), .Y(ori_ori_n382_));
  NA3        o360(.A(ori_ori_n221_), .B(ori_ori_n165_), .C(ori_ori_n136_), .Y(ori_ori_n383_));
  NA2        o361(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n384_));
  NO2        o362(.A(ori_ori_n156_), .B(i_3_), .Y(ori_ori_n385_));
  NAi31      o363(.An(ori_ori_n384_), .B(ori_ori_n385_), .C(ori_ori_n208_), .Y(ori_ori_n386_));
  NA3        o364(.A(ori_ori_n315_), .B(ori_ori_n170_), .C(ori_ori_n152_), .Y(ori_ori_n387_));
  NA3        o365(.A(ori_ori_n387_), .B(ori_ori_n386_), .C(ori_ori_n383_), .Y(ori_ori_n388_));
  NO2        o366(.A(ori_ori_n388_), .B(ori_ori_n375_), .Y(ori_ori_n389_));
  NA2        o367(.A(ori_ori_n355_), .B(ori_ori_n308_), .Y(ori_ori_n390_));
  NA2        o368(.A(ori_ori_n364_), .B(ori_ori_n314_), .Y(ori_ori_n391_));
  NAi21      o369(.An(ori_ori_n198_), .B(ori_ori_n319_), .Y(ori_ori_n392_));
  NA2        o370(.A(ori_ori_n267_), .B(ori_ori_n200_), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n393_), .B(ori_ori_n392_), .Y(ori_ori_n394_));
  NA2        o372(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n395_));
  NA2        o373(.A(ori_ori_n259_), .B(ori_ori_n216_), .Y(ori_ori_n396_));
  OAI220     o374(.A0(ori_ori_n396_), .A1(ori_ori_n338_), .B0(ori_ori_n395_), .B1(ori_ori_n372_), .Y(ori_ori_n397_));
  NO2        o375(.A(ori_ori_n397_), .B(ori_ori_n394_), .Y(ori_ori_n398_));
  NA4        o376(.A(ori_ori_n398_), .B(ori_ori_n389_), .C(ori_ori_n371_), .D(ori_ori_n369_), .Y(ori_ori_n399_));
  NA2        o377(.A(ori_ori_n126_), .B(ori_ori_n115_), .Y(ori_ori_n400_));
  AN2        o378(.A(ori_ori_n400_), .B(ori_ori_n355_), .Y(ori_ori_n401_));
  NA2        o379(.A(ori_ori_n401_), .B(ori_ori_n257_), .Y(ori_ori_n402_));
  NA4        o380(.A(ori_ori_n345_), .B(ori_ori_n344_), .C(ori_ori_n186_), .D(i_2_), .Y(ori_ori_n403_));
  INV        o381(.A(ori_ori_n403_), .Y(ori_ori_n404_));
  NA2        o382(.A(ori_ori_n308_), .B(ori_ori_n207_), .Y(ori_ori_n405_));
  NA2        o383(.A(ori_ori_n277_), .B(ori_ori_n73_), .Y(ori_ori_n406_));
  NA2        o384(.A(ori_ori_n295_), .B(ori_ori_n287_), .Y(ori_ori_n407_));
  OR2        o385(.A(ori_ori_n405_), .B(ori_ori_n407_), .Y(ori_ori_n408_));
  NO2        o386(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n409_));
  AOI210     o387(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n329_), .Y(ori_ori_n410_));
  NA2        o388(.A(ori_ori_n410_), .B(ori_ori_n408_), .Y(ori_ori_n411_));
  AOI210     o389(.A0(ori_ori_n404_), .A1(ori_ori_n187_), .B0(ori_ori_n411_), .Y(ori_ori_n412_));
  NA2        o390(.A(ori_ori_n229_), .B(ori_ori_n64_), .Y(ori_ori_n413_));
  OAI210     o391(.A0(i_8_), .A1(ori_ori_n413_), .B0(ori_ori_n138_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n414_), .B(ori_ori_n330_), .Y(ori_ori_n415_));
  NA3        o393(.A(ori_ori_n415_), .B(ori_ori_n412_), .C(ori_ori_n402_), .Y(ori_ori_n416_));
  NO2        o394(.A(i_12_), .B(ori_ori_n179_), .Y(ori_ori_n417_));
  NO2        o395(.A(i_8_), .B(i_7_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n419_));
  NO2        o397(.A(ori_ori_n419_), .B(i_6_), .Y(ori_ori_n420_));
  AOI220     o398(.A0(ori_ori_n336_), .A1(ori_ori_n262_), .B0(ori_ori_n223_), .B1(ori_ori_n220_), .Y(ori_ori_n421_));
  OAI220     o399(.A0(ori_ori_n421_), .A1(ori_ori_n236_), .B0(ori_ori_n372_), .B1(ori_ori_n137_), .Y(ori_ori_n422_));
  NA2        o400(.A(ori_ori_n422_), .B(ori_ori_n239_), .Y(ori_ori_n423_));
  NA3        o401(.A(ori_ori_n255_), .B(ori_ori_n167_), .C(ori_ori_n99_), .Y(ori_ori_n424_));
  NO2        o402(.A(ori_ori_n204_), .B(ori_ori_n44_), .Y(ori_ori_n425_));
  NO2        o403(.A(ori_ori_n156_), .B(i_5_), .Y(ori_ori_n426_));
  NA3        o404(.A(ori_ori_n426_), .B(ori_ori_n322_), .C(ori_ori_n260_), .Y(ori_ori_n427_));
  OAI210     o405(.A0(ori_ori_n427_), .A1(ori_ori_n425_), .B0(ori_ori_n424_), .Y(ori_ori_n428_));
  NA2        o406(.A(ori_ori_n428_), .B(ori_ori_n364_), .Y(ori_ori_n429_));
  NA2        o407(.A(ori_ori_n429_), .B(ori_ori_n423_), .Y(ori_ori_n430_));
  NA3        o408(.A(ori_ori_n200_), .B(ori_ori_n71_), .C(ori_ori_n44_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n252_), .B(ori_ori_n84_), .Y(ori_ori_n432_));
  NO2        o410(.A(ori_ori_n431_), .B(ori_ori_n432_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n206_), .B(ori_ori_n205_), .Y(ori_ori_n434_));
  NA2        o412(.A(ori_ori_n347_), .B(ori_ori_n204_), .Y(ori_ori_n435_));
  NO2        o413(.A(ori_ori_n434_), .B(ori_ori_n435_), .Y(ori_ori_n436_));
  AOI210     o414(.A0(ori_ori_n288_), .A1(ori_ori_n46_), .B0(ori_ori_n292_), .Y(ori_ori_n437_));
  NA2        o415(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n438_));
  NA3        o416(.A(ori_ori_n417_), .B(ori_ori_n248_), .C(ori_ori_n438_), .Y(ori_ori_n439_));
  NO2        o417(.A(ori_ori_n437_), .B(ori_ori_n439_), .Y(ori_ori_n440_));
  NO3        o418(.A(ori_ori_n440_), .B(ori_ori_n436_), .C(ori_ori_n433_), .Y(ori_ori_n441_));
  NO4        o419(.A(ori_ori_n225_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n442_));
  NO3        o420(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n443_));
  NO2        o421(.A(ori_ori_n328_), .B(i_1_), .Y(ori_ori_n444_));
  NOi31      o422(.An(ori_ori_n444_), .B(ori_ori_n356_), .C(ori_ori_n73_), .Y(ori_ori_n445_));
  NOi21      o423(.An(i_10_), .B(i_6_), .Y(ori_ori_n446_));
  NO2        o424(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n447_));
  AOI220     o425(.A0(ori_ori_n252_), .A1(ori_ori_n447_), .B0(ori_ori_n248_), .B1(ori_ori_n446_), .Y(ori_ori_n448_));
  NO2        o426(.A(ori_ori_n448_), .B(ori_ori_n354_), .Y(ori_ori_n449_));
  NO2        o427(.A(ori_ori_n118_), .B(ori_ori_n23_), .Y(ori_ori_n450_));
  NO2        o428(.A(ori_ori_n182_), .B(ori_ori_n37_), .Y(ori_ori_n451_));
  NOi31      o429(.An(ori_ori_n149_), .B(ori_ori_n451_), .C(ori_ori_n265_), .Y(ori_ori_n452_));
  NO2        o430(.A(ori_ori_n452_), .B(ori_ori_n449_), .Y(ori_ori_n453_));
  NO2        o431(.A(ori_ori_n406_), .B(ori_ori_n303_), .Y(ori_ori_n454_));
  INV        o432(.A(ori_ori_n260_), .Y(ori_ori_n455_));
  NO2        o433(.A(i_12_), .B(ori_ori_n86_), .Y(ori_ori_n456_));
  NA3        o434(.A(ori_ori_n456_), .B(ori_ori_n248_), .C(ori_ori_n438_), .Y(ori_ori_n457_));
  NA3        o435(.A(ori_ori_n311_), .B(ori_ori_n252_), .C(ori_ori_n200_), .Y(ori_ori_n458_));
  AOI210     o436(.A0(ori_ori_n458_), .A1(ori_ori_n457_), .B0(ori_ori_n455_), .Y(ori_ori_n459_));
  OR2        o437(.A(i_2_), .B(i_5_), .Y(ori_ori_n460_));
  OR2        o438(.A(ori_ori_n460_), .B(ori_ori_n325_), .Y(ori_ori_n461_));
  AOI210     o439(.A0(ori_ori_n297_), .A1(ori_ori_n220_), .B0(ori_ori_n182_), .Y(ori_ori_n462_));
  AOI210     o440(.A0(ori_ori_n462_), .A1(ori_ori_n461_), .B0(ori_ori_n392_), .Y(ori_ori_n463_));
  NO3        o441(.A(ori_ori_n463_), .B(ori_ori_n459_), .C(ori_ori_n454_), .Y(ori_ori_n464_));
  NA3        o442(.A(ori_ori_n464_), .B(ori_ori_n453_), .C(ori_ori_n441_), .Y(ori_ori_n465_));
  NO4        o443(.A(ori_ori_n465_), .B(ori_ori_n430_), .C(ori_ori_n416_), .D(ori_ori_n399_), .Y(ori_ori_n466_));
  NA4        o444(.A(ori_ori_n466_), .B(ori_ori_n343_), .C(ori_ori_n276_), .D(ori_ori_n258_), .Y(ori7));
  NO2        o445(.A(ori_ori_n95_), .B(ori_ori_n54_), .Y(ori_ori_n468_));
  NO2        o446(.A(ori_ori_n111_), .B(ori_ori_n92_), .Y(ori_ori_n469_));
  NA2        o447(.A(ori_ori_n309_), .B(ori_ori_n469_), .Y(ori_ori_n470_));
  NA2        o448(.A(ori_ori_n382_), .B(ori_ori_n84_), .Y(ori_ori_n471_));
  NA2        o449(.A(i_11_), .B(ori_ori_n179_), .Y(ori_ori_n472_));
  NA2        o450(.A(ori_ori_n147_), .B(ori_ori_n472_), .Y(ori_ori_n473_));
  OAI210     o451(.A0(ori_ori_n473_), .A1(ori_ori_n471_), .B0(ori_ori_n470_), .Y(ori_ori_n474_));
  NA3        o452(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n475_));
  NO2        o453(.A(ori_ori_n214_), .B(i_4_), .Y(ori_ori_n476_));
  NA2        o454(.A(ori_ori_n476_), .B(i_8_), .Y(ori_ori_n477_));
  NO2        o455(.A(ori_ori_n108_), .B(ori_ori_n475_), .Y(ori_ori_n478_));
  NA2        o456(.A(i_2_), .B(ori_ori_n86_), .Y(ori_ori_n479_));
  OAI210     o457(.A0(ori_ori_n89_), .A1(ori_ori_n186_), .B0(ori_ori_n187_), .Y(ori_ori_n480_));
  NO2        o458(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n481_));
  NA2        o459(.A(i_4_), .B(i_8_), .Y(ori_ori_n482_));
  AOI210     o460(.A0(ori_ori_n482_), .A1(ori_ori_n255_), .B0(ori_ori_n481_), .Y(ori_ori_n483_));
  OAI220     o461(.A0(ori_ori_n483_), .A1(ori_ori_n479_), .B0(ori_ori_n480_), .B1(i_13_), .Y(ori_ori_n484_));
  NO4        o462(.A(ori_ori_n484_), .B(ori_ori_n478_), .C(ori_ori_n474_), .D(ori_ori_n468_), .Y(ori_ori_n485_));
  AOI210     o463(.A0(ori_ori_n132_), .A1(ori_ori_n62_), .B0(i_10_), .Y(ori_ori_n486_));
  AOI210     o464(.A0(ori_ori_n486_), .A1(ori_ori_n214_), .B0(ori_ori_n160_), .Y(ori_ori_n487_));
  OR2        o465(.A(i_6_), .B(i_10_), .Y(ori_ori_n488_));
  NO2        o466(.A(ori_ori_n488_), .B(ori_ori_n23_), .Y(ori_ori_n489_));
  OR3        o467(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n490_));
  NO3        o468(.A(ori_ori_n490_), .B(i_8_), .C(ori_ori_n31_), .Y(ori_ori_n491_));
  INV        o469(.A(ori_ori_n183_), .Y(ori_ori_n492_));
  NO2        o470(.A(ori_ori_n491_), .B(ori_ori_n489_), .Y(ori_ori_n493_));
  OA220      o471(.A0(ori_ori_n493_), .A1(ori_ori_n455_), .B0(ori_ori_n487_), .B1(ori_ori_n241_), .Y(ori_ori_n494_));
  AOI210     o472(.A0(ori_ori_n494_), .A1(ori_ori_n485_), .B0(ori_ori_n63_), .Y(ori_ori_n495_));
  NOi21      o473(.An(i_11_), .B(i_7_), .Y(ori_ori_n496_));
  AO210      o474(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n497_));
  NO2        o475(.A(ori_ori_n497_), .B(ori_ori_n496_), .Y(ori_ori_n498_));
  NA2        o476(.A(ori_ori_n498_), .B(ori_ori_n191_), .Y(ori_ori_n499_));
  NA3        o477(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n500_));
  NAi31      o478(.An(ori_ori_n500_), .B(ori_ori_n197_), .C(i_11_), .Y(ori_ori_n501_));
  AOI210     o479(.A0(ori_ori_n501_), .A1(ori_ori_n499_), .B0(ori_ori_n63_), .Y(ori_ori_n502_));
  NA2        o480(.A(ori_ori_n88_), .B(ori_ori_n63_), .Y(ori_ori_n503_));
  AO210      o481(.A0(ori_ori_n503_), .A1(ori_ori_n303_), .B0(ori_ori_n41_), .Y(ori_ori_n504_));
  NO3        o482(.A(ori_ori_n231_), .B(ori_ori_n192_), .C(ori_ori_n472_), .Y(ori_ori_n505_));
  OAI210     o483(.A0(ori_ori_n505_), .A1(ori_ori_n208_), .B0(ori_ori_n63_), .Y(ori_ori_n506_));
  NA2        o484(.A(ori_ori_n326_), .B(ori_ori_n31_), .Y(ori_ori_n507_));
  OR2        o485(.A(ori_ori_n192_), .B(ori_ori_n111_), .Y(ori_ori_n508_));
  NA2        o486(.A(ori_ori_n508_), .B(ori_ori_n507_), .Y(ori_ori_n509_));
  NO2        o487(.A(ori_ori_n63_), .B(i_9_), .Y(ori_ori_n510_));
  NO2        o488(.A(ori_ori_n510_), .B(i_4_), .Y(ori_ori_n511_));
  NA2        o489(.A(ori_ori_n511_), .B(ori_ori_n509_), .Y(ori_ori_n512_));
  NO2        o490(.A(i_1_), .B(i_12_), .Y(ori_ori_n513_));
  NA3        o491(.A(ori_ori_n513_), .B(ori_ori_n113_), .C(ori_ori_n24_), .Y(ori_ori_n514_));
  BUFFER     o492(.A(ori_ori_n514_), .Y(ori_ori_n515_));
  NA4        o493(.A(ori_ori_n515_), .B(ori_ori_n512_), .C(ori_ori_n506_), .D(ori_ori_n504_), .Y(ori_ori_n516_));
  OAI210     o494(.A0(ori_ori_n516_), .A1(ori_ori_n502_), .B0(i_6_), .Y(ori_ori_n517_));
  NO2        o495(.A(ori_ori_n500_), .B(ori_ori_n111_), .Y(ori_ori_n518_));
  NA2        o496(.A(ori_ori_n518_), .B(ori_ori_n456_), .Y(ori_ori_n519_));
  NO2        o497(.A(ori_ori_n214_), .B(ori_ori_n86_), .Y(ori_ori_n520_));
  NO2        o498(.A(ori_ori_n520_), .B(i_11_), .Y(ori_ori_n521_));
  NA2        o499(.A(ori_ori_n519_), .B(ori_ori_n357_), .Y(ori_ori_n522_));
  NO3        o500(.A(ori_ori_n488_), .B(ori_ori_n213_), .C(ori_ori_n23_), .Y(ori_ori_n523_));
  AOI210     o501(.A0(i_1_), .A1(ori_ori_n232_), .B0(ori_ori_n523_), .Y(ori_ori_n524_));
  NO2        o502(.A(ori_ori_n524_), .B(ori_ori_n44_), .Y(ori_ori_n525_));
  NA3        o503(.A(ori_ori_n418_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n526_));
  INV        o504(.A(i_2_), .Y(ori_ori_n527_));
  NA2        o505(.A(ori_ori_n142_), .B(i_9_), .Y(ori_ori_n528_));
  NA3        o506(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n529_));
  NO2        o507(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n530_));
  NA3        o508(.A(ori_ori_n530_), .B(ori_ori_n240_), .C(ori_ori_n44_), .Y(ori_ori_n531_));
  OAI220     o509(.A0(ori_ori_n531_), .A1(ori_ori_n529_), .B0(ori_ori_n528_), .B1(ori_ori_n527_), .Y(ori_ori_n532_));
  AOI210     o510(.A0(ori_ori_n378_), .A1(ori_ori_n331_), .B0(ori_ori_n218_), .Y(ori_ori_n533_));
  NO2        o511(.A(ori_ori_n533_), .B(ori_ori_n479_), .Y(ori_ori_n534_));
  NAi21      o512(.An(ori_ori_n526_), .B(ori_ori_n94_), .Y(ori_ori_n535_));
  NA2        o513(.A(ori_ori_n530_), .B(ori_ori_n240_), .Y(ori_ori_n536_));
  NO2        o514(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n537_));
  NA2        o515(.A(ori_ori_n537_), .B(ori_ori_n24_), .Y(ori_ori_n538_));
  OAI210     o516(.A0(ori_ori_n538_), .A1(ori_ori_n536_), .B0(ori_ori_n535_), .Y(ori_ori_n539_));
  OR3        o517(.A(ori_ori_n539_), .B(ori_ori_n534_), .C(ori_ori_n532_), .Y(ori_ori_n540_));
  NO3        o518(.A(ori_ori_n540_), .B(ori_ori_n525_), .C(ori_ori_n522_), .Y(ori_ori_n541_));
  NO2        o519(.A(ori_ori_n214_), .B(ori_ori_n104_), .Y(ori_ori_n542_));
  NO2        o520(.A(ori_ori_n542_), .B(ori_ori_n496_), .Y(ori_ori_n543_));
  NA2        o521(.A(ori_ori_n543_), .B(i_1_), .Y(ori_ori_n544_));
  NO2        o522(.A(ori_ori_n544_), .B(ori_ori_n490_), .Y(ori_ori_n545_));
  NO2        o523(.A(ori_ori_n327_), .B(ori_ori_n86_), .Y(ori_ori_n546_));
  NA2        o524(.A(ori_ori_n545_), .B(ori_ori_n46_), .Y(ori_ori_n547_));
  NA2        o525(.A(i_3_), .B(ori_ori_n179_), .Y(ori_ori_n548_));
  NO2        o526(.A(ori_ori_n548_), .B(ori_ori_n118_), .Y(ori_ori_n549_));
  AN2        o527(.A(ori_ori_n549_), .B(ori_ori_n420_), .Y(ori_ori_n550_));
  NO2        o528(.A(ori_ori_n213_), .B(ori_ori_n44_), .Y(ori_ori_n551_));
  NO3        o529(.A(ori_ori_n551_), .B(ori_ori_n257_), .C(ori_ori_n215_), .Y(ori_ori_n552_));
  NO2        o530(.A(ori_ori_n121_), .B(ori_ori_n37_), .Y(ori_ori_n553_));
  NO2        o531(.A(ori_ori_n553_), .B(i_6_), .Y(ori_ori_n554_));
  NO2        o532(.A(ori_ori_n86_), .B(i_9_), .Y(ori_ori_n555_));
  NO2        o533(.A(ori_ori_n555_), .B(ori_ori_n63_), .Y(ori_ori_n556_));
  NO2        o534(.A(ori_ori_n556_), .B(ori_ori_n513_), .Y(ori_ori_n557_));
  NO4        o535(.A(ori_ori_n557_), .B(ori_ori_n554_), .C(ori_ori_n552_), .D(i_4_), .Y(ori_ori_n558_));
  NA2        o536(.A(i_1_), .B(i_3_), .Y(ori_ori_n559_));
  NO2        o537(.A(ori_ori_n358_), .B(ori_ori_n95_), .Y(ori_ori_n560_));
  AOI210     o538(.A0(ori_ori_n551_), .A1(ori_ori_n446_), .B0(ori_ori_n560_), .Y(ori_ori_n561_));
  NO2        o539(.A(ori_ori_n561_), .B(ori_ori_n559_), .Y(ori_ori_n562_));
  NO3        o540(.A(ori_ori_n562_), .B(ori_ori_n558_), .C(ori_ori_n550_), .Y(ori_ori_n563_));
  NA4        o541(.A(ori_ori_n563_), .B(ori_ori_n547_), .C(ori_ori_n541_), .D(ori_ori_n517_), .Y(ori_ori_n564_));
  AN2        o542(.A(ori_ori_n221_), .B(ori_ori_n86_), .Y(ori_ori_n565_));
  NA2        o543(.A(ori_ori_n295_), .B(ori_ori_n294_), .Y(ori_ori_n566_));
  NA3        o544(.A(ori_ori_n382_), .B(ori_ori_n409_), .C(ori_ori_n46_), .Y(ori_ori_n567_));
  NO3        o545(.A(ori_ori_n380_), .B(ori_ori_n482_), .C(ori_ori_n86_), .Y(ori_ori_n568_));
  NA2        o546(.A(ori_ori_n568_), .B(ori_ori_n25_), .Y(ori_ori_n569_));
  NA3        o547(.A(ori_ori_n160_), .B(ori_ori_n84_), .C(ori_ori_n86_), .Y(ori_ori_n570_));
  NA4        o548(.A(ori_ori_n570_), .B(ori_ori_n569_), .C(ori_ori_n567_), .D(ori_ori_n566_), .Y(ori_ori_n571_));
  OAI210     o549(.A0(ori_ori_n571_), .A1(ori_ori_n565_), .B0(i_1_), .Y(ori_ori_n572_));
  AOI210     o550(.A0(ori_ori_n240_), .A1(ori_ori_n100_), .B0(i_1_), .Y(ori_ori_n573_));
  NO2        o551(.A(ori_ori_n293_), .B(i_2_), .Y(ori_ori_n574_));
  NA2        o552(.A(ori_ori_n574_), .B(ori_ori_n573_), .Y(ori_ori_n575_));
  AOI210     o553(.A0(ori_ori_n575_), .A1(ori_ori_n572_), .B0(i_13_), .Y(ori_ori_n576_));
  OR2        o554(.A(i_11_), .B(i_7_), .Y(ori_ori_n577_));
  NA3        o555(.A(ori_ori_n577_), .B(ori_ori_n109_), .C(ori_ori_n142_), .Y(ori_ori_n578_));
  AOI220     o556(.A0(ori_ori_n374_), .A1(ori_ori_n160_), .B0(ori_ori_n351_), .B1(ori_ori_n142_), .Y(ori_ori_n579_));
  OAI210     o557(.A0(ori_ori_n579_), .A1(ori_ori_n44_), .B0(ori_ori_n578_), .Y(ori_ori_n580_));
  AOI210     o558(.A0(ori_ori_n529_), .A1(ori_ori_n54_), .B0(i_12_), .Y(ori_ori_n581_));
  NO2        o559(.A(ori_ori_n380_), .B(ori_ori_n24_), .Y(ori_ori_n582_));
  AOI220     o560(.A0(ori_ori_n582_), .A1(ori_ori_n546_), .B0(ori_ori_n221_), .B1(ori_ori_n135_), .Y(ori_ori_n583_));
  OAI220     o561(.A0(ori_ori_n583_), .A1(ori_ori_n41_), .B0(ori_ori_n894_), .B1(ori_ori_n95_), .Y(ori_ori_n584_));
  AOI210     o562(.A0(ori_ori_n580_), .A1(ori_ori_n266_), .B0(ori_ori_n584_), .Y(ori_ori_n585_));
  INV        o563(.A(ori_ori_n118_), .Y(ori_ori_n586_));
  AOI220     o564(.A0(ori_ori_n586_), .A1(ori_ori_n72_), .B0(ori_ori_n311_), .B1(ori_ori_n530_), .Y(ori_ori_n587_));
  NO2        o565(.A(ori_ori_n587_), .B(ori_ori_n219_), .Y(ori_ori_n588_));
  AOI210     o566(.A0(ori_ori_n348_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n589_));
  NOi31      o567(.An(ori_ori_n589_), .B(ori_ori_n471_), .C(ori_ori_n44_), .Y(ori_ori_n590_));
  NA2        o568(.A(ori_ori_n131_), .B(i_13_), .Y(ori_ori_n591_));
  NO2        o569(.A(ori_ori_n529_), .B(ori_ori_n118_), .Y(ori_ori_n592_));
  INV        o570(.A(ori_ori_n592_), .Y(ori_ori_n593_));
  OAI220     o571(.A0(ori_ori_n593_), .A1(ori_ori_n71_), .B0(ori_ori_n591_), .B1(ori_ori_n573_), .Y(ori_ori_n594_));
  NO3        o572(.A(ori_ori_n71_), .B(ori_ori_n32_), .C(ori_ori_n104_), .Y(ori_ori_n595_));
  NA2        o573(.A(ori_ori_n26_), .B(ori_ori_n179_), .Y(ori_ori_n596_));
  NA2        o574(.A(ori_ori_n596_), .B(i_7_), .Y(ori_ori_n597_));
  NO3        o575(.A(ori_ori_n380_), .B(ori_ori_n214_), .C(ori_ori_n86_), .Y(ori_ori_n598_));
  AOI210     o576(.A0(ori_ori_n598_), .A1(ori_ori_n597_), .B0(ori_ori_n595_), .Y(ori_ori_n599_));
  AOI220     o577(.A0(ori_ori_n311_), .A1(ori_ori_n530_), .B0(ori_ori_n94_), .B1(ori_ori_n105_), .Y(ori_ori_n600_));
  OAI220     o578(.A0(ori_ori_n600_), .A1(ori_ori_n477_), .B0(ori_ori_n599_), .B1(ori_ori_n492_), .Y(ori_ori_n601_));
  NO4        o579(.A(ori_ori_n601_), .B(ori_ori_n594_), .C(ori_ori_n590_), .D(ori_ori_n588_), .Y(ori_ori_n602_));
  OR2        o580(.A(i_11_), .B(i_6_), .Y(ori_ori_n603_));
  NA3        o581(.A(ori_ori_n476_), .B(ori_ori_n596_), .C(i_7_), .Y(ori_ori_n604_));
  AOI210     o582(.A0(ori_ori_n604_), .A1(ori_ori_n593_), .B0(ori_ori_n603_), .Y(ori_ori_n605_));
  NA3        o583(.A(ori_ori_n326_), .B(ori_ori_n481_), .C(ori_ori_n100_), .Y(ori_ori_n606_));
  NA2        o584(.A(ori_ori_n521_), .B(i_13_), .Y(ori_ori_n607_));
  NA2        o585(.A(ori_ori_n105_), .B(ori_ori_n596_), .Y(ori_ori_n608_));
  NAi21      o586(.An(i_11_), .B(i_12_), .Y(ori_ori_n609_));
  NOi41      o587(.An(ori_ori_n114_), .B(ori_ori_n609_), .C(i_13_), .D(ori_ori_n86_), .Y(ori_ori_n610_));
  NO3        o588(.A(ori_ori_n380_), .B(ori_ori_n456_), .C(ori_ori_n482_), .Y(ori_ori_n611_));
  AOI220     o589(.A0(ori_ori_n611_), .A1(ori_ori_n259_), .B0(ori_ori_n610_), .B1(ori_ori_n608_), .Y(ori_ori_n612_));
  NA3        o590(.A(ori_ori_n612_), .B(ori_ori_n607_), .C(ori_ori_n606_), .Y(ori_ori_n613_));
  OAI210     o591(.A0(ori_ori_n613_), .A1(ori_ori_n605_), .B0(ori_ori_n63_), .Y(ori_ori_n614_));
  NO2        o592(.A(i_2_), .B(i_12_), .Y(ori_ori_n615_));
  NA2        o593(.A(ori_ori_n292_), .B(ori_ori_n615_), .Y(ori_ori_n616_));
  NA2        o594(.A(i_8_), .B(ori_ori_n25_), .Y(ori_ori_n617_));
  NO3        o595(.A(ori_ori_n617_), .B(ori_ori_n309_), .C(ori_ori_n476_), .Y(ori_ori_n618_));
  OAI210     o596(.A0(ori_ori_n618_), .A1(ori_ori_n294_), .B0(ori_ori_n292_), .Y(ori_ori_n619_));
  NO2        o597(.A(ori_ori_n132_), .B(i_2_), .Y(ori_ori_n620_));
  NA2        o598(.A(ori_ori_n620_), .B(ori_ori_n513_), .Y(ori_ori_n621_));
  NA3        o599(.A(ori_ori_n621_), .B(ori_ori_n619_), .C(ori_ori_n616_), .Y(ori_ori_n622_));
  NA3        o600(.A(ori_ori_n622_), .B(ori_ori_n45_), .C(ori_ori_n207_), .Y(ori_ori_n623_));
  NA4        o601(.A(ori_ori_n623_), .B(ori_ori_n614_), .C(ori_ori_n602_), .D(ori_ori_n585_), .Y(ori_ori_n624_));
  OR4        o602(.A(ori_ori_n624_), .B(ori_ori_n576_), .C(ori_ori_n564_), .D(ori_ori_n495_), .Y(ori5));
  NA2        o603(.A(ori_ori_n543_), .B(ori_ori_n243_), .Y(ori_ori_n626_));
  AN2        o604(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n627_));
  NA3        o605(.A(ori_ori_n627_), .B(ori_ori_n615_), .C(ori_ori_n111_), .Y(ori_ori_n628_));
  NO2        o606(.A(ori_ori_n477_), .B(i_11_), .Y(ori_ori_n629_));
  OAI210     o607(.A0(ori_ori_n481_), .A1(ori_ori_n89_), .B0(ori_ori_n629_), .Y(ori_ori_n630_));
  NA3        o608(.A(ori_ori_n630_), .B(ori_ori_n628_), .C(ori_ori_n626_), .Y(ori_ori_n631_));
  NO3        o609(.A(i_11_), .B(ori_ori_n214_), .C(i_13_), .Y(ori_ori_n632_));
  NO2        o610(.A(ori_ori_n128_), .B(ori_ori_n23_), .Y(ori_ori_n633_));
  NA2        o611(.A(i_12_), .B(i_8_), .Y(ori_ori_n634_));
  OAI210     o612(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n634_), .Y(ori_ori_n635_));
  INV        o613(.A(ori_ori_n347_), .Y(ori_ori_n636_));
  AOI220     o614(.A0(ori_ori_n260_), .A1(ori_ori_n450_), .B0(ori_ori_n635_), .B1(ori_ori_n633_), .Y(ori_ori_n637_));
  INV        o615(.A(ori_ori_n637_), .Y(ori_ori_n638_));
  NO2        o616(.A(ori_ori_n638_), .B(ori_ori_n631_), .Y(ori_ori_n639_));
  INV        o617(.A(ori_ori_n165_), .Y(ori_ori_n640_));
  INV        o618(.A(ori_ori_n221_), .Y(ori_ori_n641_));
  OAI210     o619(.A0(ori_ori_n574_), .A1(ori_ori_n349_), .B0(ori_ori_n114_), .Y(ori_ori_n642_));
  AOI210     o620(.A0(ori_ori_n642_), .A1(ori_ori_n641_), .B0(ori_ori_n640_), .Y(ori_ori_n643_));
  NO2        o621(.A(ori_ori_n358_), .B(ori_ori_n26_), .Y(ori_ori_n644_));
  NO2        o622(.A(ori_ori_n644_), .B(ori_ori_n331_), .Y(ori_ori_n645_));
  NA2        o623(.A(ori_ori_n645_), .B(i_2_), .Y(ori_ori_n646_));
  INV        o624(.A(ori_ori_n646_), .Y(ori_ori_n647_));
  AOI210     o625(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n328_), .Y(ori_ori_n648_));
  AOI210     o626(.A0(ori_ori_n648_), .A1(ori_ori_n647_), .B0(ori_ori_n643_), .Y(ori_ori_n649_));
  NO2        o627(.A(ori_ori_n178_), .B(ori_ori_n129_), .Y(ori_ori_n650_));
  OAI210     o628(.A0(ori_ori_n650_), .A1(ori_ori_n633_), .B0(i_2_), .Y(ori_ori_n651_));
  INV        o629(.A(ori_ori_n166_), .Y(ori_ori_n652_));
  NO3        o630(.A(ori_ori_n497_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n653_));
  AOI210     o631(.A0(ori_ori_n652_), .A1(ori_ori_n89_), .B0(ori_ori_n653_), .Y(ori_ori_n654_));
  AOI210     o632(.A0(ori_ori_n654_), .A1(ori_ori_n651_), .B0(ori_ori_n179_), .Y(ori_ori_n655_));
  OA210      o633(.A0(ori_ori_n498_), .A1(ori_ori_n130_), .B0(i_13_), .Y(ori_ori_n656_));
  NA2        o634(.A(ori_ori_n183_), .B(ori_ori_n186_), .Y(ori_ori_n657_));
  NA2        o635(.A(ori_ori_n154_), .B(ori_ori_n472_), .Y(ori_ori_n658_));
  AOI210     o636(.A0(ori_ori_n658_), .A1(ori_ori_n657_), .B0(ori_ori_n297_), .Y(ori_ori_n659_));
  AOI210     o637(.A0(ori_ori_n192_), .A1(ori_ori_n151_), .B0(ori_ori_n409_), .Y(ori_ori_n660_));
  OAI210     o638(.A0(ori_ori_n660_), .A1(ori_ori_n208_), .B0(ori_ori_n331_), .Y(ori_ori_n661_));
  NO2        o639(.A(ori_ori_n105_), .B(ori_ori_n44_), .Y(ori_ori_n662_));
  INV        o640(.A(ori_ori_n254_), .Y(ori_ori_n663_));
  NA4        o641(.A(ori_ori_n663_), .B(ori_ori_n255_), .C(ori_ori_n128_), .D(ori_ori_n42_), .Y(ori_ori_n664_));
  OAI210     o642(.A0(ori_ori_n664_), .A1(ori_ori_n662_), .B0(ori_ori_n661_), .Y(ori_ori_n665_));
  NO4        o643(.A(ori_ori_n665_), .B(ori_ori_n659_), .C(ori_ori_n656_), .D(ori_ori_n655_), .Y(ori_ori_n666_));
  NA2        o644(.A(ori_ori_n450_), .B(ori_ori_n28_), .Y(ori_ori_n667_));
  NA2        o645(.A(ori_ori_n632_), .B(ori_ori_n249_), .Y(ori_ori_n668_));
  NA2        o646(.A(ori_ori_n668_), .B(ori_ori_n667_), .Y(ori_ori_n669_));
  NO2        o647(.A(ori_ori_n62_), .B(i_12_), .Y(ori_ori_n670_));
  NO2        o648(.A(ori_ori_n670_), .B(ori_ori_n130_), .Y(ori_ori_n671_));
  NO2        o649(.A(ori_ori_n671_), .B(ori_ori_n472_), .Y(ori_ori_n672_));
  AOI220     o650(.A0(ori_ori_n672_), .A1(ori_ori_n36_), .B0(ori_ori_n669_), .B1(ori_ori_n46_), .Y(ori_ori_n673_));
  NA4        o651(.A(ori_ori_n673_), .B(ori_ori_n666_), .C(ori_ori_n649_), .D(ori_ori_n639_), .Y(ori6));
  NA4        o652(.A(ori_ori_n314_), .B(ori_ori_n381_), .C(ori_ori_n71_), .D(ori_ori_n104_), .Y(ori_ori_n675_));
  INV        o653(.A(ori_ori_n675_), .Y(ori_ori_n676_));
  NO2        o654(.A(ori_ori_n203_), .B(ori_ori_n384_), .Y(ori_ori_n677_));
  NO2        o655(.A(i_11_), .B(i_9_), .Y(ori_ori_n678_));
  NO2        o656(.A(ori_ori_n676_), .B(ori_ori_n264_), .Y(ori_ori_n679_));
  OR2        o657(.A(ori_ori_n679_), .B(i_12_), .Y(ori_ori_n680_));
  NA2        o658(.A(ori_ori_n298_), .B(ori_ori_n267_), .Y(ori_ori_n681_));
  NA2        o659(.A(ori_ori_n456_), .B(ori_ori_n63_), .Y(ori_ori_n682_));
  BUFFER     o660(.A(ori_ori_n503_), .Y(ori_ori_n683_));
  NA3        o661(.A(ori_ori_n683_), .B(ori_ori_n682_), .C(ori_ori_n681_), .Y(ori_ori_n684_));
  INV        o662(.A(ori_ori_n181_), .Y(ori_ori_n685_));
  AOI220     o663(.A0(ori_ori_n685_), .A1(ori_ori_n678_), .B0(ori_ori_n684_), .B1(ori_ori_n73_), .Y(ori_ori_n686_));
  INV        o664(.A(ori_ori_n263_), .Y(ori_ori_n687_));
  NA2        o665(.A(ori_ori_n75_), .B(ori_ori_n135_), .Y(ori_ori_n688_));
  INV        o666(.A(ori_ori_n128_), .Y(ori_ori_n689_));
  NA2        o667(.A(ori_ori_n689_), .B(ori_ori_n46_), .Y(ori_ori_n690_));
  AOI210     o668(.A0(ori_ori_n690_), .A1(ori_ori_n688_), .B0(ori_ori_n687_), .Y(ori_ori_n691_));
  NO3        o669(.A(ori_ori_n225_), .B(ori_ori_n136_), .C(i_9_), .Y(ori_ori_n692_));
  NA2        o670(.A(ori_ori_n692_), .B(ori_ori_n670_), .Y(ori_ori_n693_));
  AOI210     o671(.A0(ori_ori_n693_), .A1(ori_ori_n407_), .B0(ori_ori_n173_), .Y(ori_ori_n694_));
  NO2        o672(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n695_));
  NAi32      o673(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n696_));
  AOI210     o674(.A0(ori_ori_n603_), .A1(ori_ori_n87_), .B0(ori_ori_n696_), .Y(ori_ori_n697_));
  OR3        o675(.A(ori_ori_n697_), .B(ori_ori_n694_), .C(ori_ori_n691_), .Y(ori_ori_n698_));
  NO2        o676(.A(ori_ori_n577_), .B(i_2_), .Y(ori_ori_n699_));
  NA2        o677(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n700_));
  OAI210     o678(.A0(ori_ori_n700_), .A1(ori_ori_n325_), .B0(ori_ori_n282_), .Y(ori_ori_n701_));
  NA2        o679(.A(ori_ori_n701_), .B(ori_ori_n699_), .Y(ori_ori_n702_));
  OR2        o680(.A(ori_ori_n498_), .B(ori_ori_n349_), .Y(ori_ori_n703_));
  NA3        o681(.A(ori_ori_n703_), .B(ori_ori_n150_), .C(ori_ori_n69_), .Y(ori_ori_n704_));
  AO210      o682(.A0(ori_ori_n391_), .A1(ori_ori_n636_), .B0(ori_ori_n36_), .Y(ori_ori_n705_));
  NA3        o683(.A(ori_ori_n705_), .B(ori_ori_n704_), .C(ori_ori_n702_), .Y(ori_ori_n706_));
  OAI210     o684(.A0(ori_ori_n520_), .A1(i_11_), .B0(ori_ori_n87_), .Y(ori_ori_n707_));
  AOI220     o685(.A0(ori_ori_n707_), .A1(ori_ori_n443_), .B0(ori_ori_n677_), .B1(ori_ori_n597_), .Y(ori_ori_n708_));
  NA3        o686(.A(ori_ori_n297_), .B(ori_ori_n216_), .C(ori_ori_n150_), .Y(ori_ori_n709_));
  NA2        o687(.A(ori_ori_n318_), .B(ori_ori_n70_), .Y(ori_ori_n710_));
  NA4        o688(.A(ori_ori_n710_), .B(ori_ori_n709_), .C(ori_ori_n708_), .D(ori_ori_n480_), .Y(ori_ori_n711_));
  AO210      o689(.A0(ori_ori_n409_), .A1(ori_ori_n46_), .B0(ori_ori_n88_), .Y(ori_ori_n712_));
  NA3        o690(.A(ori_ori_n712_), .B(ori_ori_n382_), .C(ori_ori_n200_), .Y(ori_ori_n713_));
  AOI210     o691(.A0(ori_ori_n349_), .A1(ori_ori_n347_), .B0(ori_ori_n442_), .Y(ori_ori_n714_));
  NO2        o692(.A(ori_ori_n488_), .B(ori_ori_n105_), .Y(ori_ori_n715_));
  OAI210     o693(.A0(ori_ori_n715_), .A1(ori_ori_n115_), .B0(ori_ori_n324_), .Y(ori_ori_n716_));
  NA2        o694(.A(ori_ori_n220_), .B(ori_ori_n46_), .Y(ori_ori_n717_));
  INV        o695(.A(ori_ori_n461_), .Y(ori_ori_n718_));
  NA3        o696(.A(ori_ori_n718_), .B(ori_ori_n263_), .C(i_7_), .Y(ori_ori_n719_));
  NA4        o697(.A(ori_ori_n719_), .B(ori_ori_n716_), .C(ori_ori_n714_), .D(ori_ori_n713_), .Y(ori_ori_n720_));
  NO4        o698(.A(ori_ori_n720_), .B(ori_ori_n711_), .C(ori_ori_n706_), .D(ori_ori_n698_), .Y(ori_ori_n721_));
  NA4        o699(.A(ori_ori_n721_), .B(ori_ori_n686_), .C(ori_ori_n680_), .D(ori_ori_n305_), .Y(ori3));
  NA2        o700(.A(i_12_), .B(i_10_), .Y(ori_ori_n723_));
  NO2        o701(.A(i_11_), .B(ori_ori_n214_), .Y(ori_ori_n724_));
  NA3        o702(.A(ori_ori_n709_), .B(ori_ori_n480_), .C(ori_ori_n296_), .Y(ori_ori_n725_));
  NA2        o703(.A(ori_ori_n725_), .B(ori_ori_n40_), .Y(ori_ori_n726_));
  NOi21      o704(.An(ori_ori_n99_), .B(ori_ori_n645_), .Y(ori_ori_n727_));
  NO3        o705(.A(ori_ori_n508_), .B(ori_ori_n358_), .C(ori_ori_n135_), .Y(ori_ori_n728_));
  NA2        o706(.A(ori_ori_n326_), .B(ori_ori_n45_), .Y(ori_ori_n729_));
  AN2        o707(.A(ori_ori_n356_), .B(ori_ori_n55_), .Y(ori_ori_n730_));
  NO3        o708(.A(ori_ori_n730_), .B(ori_ori_n728_), .C(ori_ori_n727_), .Y(ori_ori_n731_));
  AOI210     o709(.A0(ori_ori_n731_), .A1(ori_ori_n726_), .B0(ori_ori_n48_), .Y(ori_ori_n732_));
  NO4        o710(.A(ori_ori_n301_), .B(ori_ori_n308_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n733_));
  NA2        o711(.A(ori_ori_n173_), .B(ori_ori_n446_), .Y(ori_ori_n734_));
  NOi31      o712(.An(ori_ori_n734_), .B(ori_ori_n733_), .C(ori_ori_n39_), .Y(ori_ori_n735_));
  NO2        o713(.A(ori_ori_n735_), .B(ori_ori_n63_), .Y(ori_ori_n736_));
  NOi21      o714(.An(i_5_), .B(i_9_), .Y(ori_ori_n737_));
  NA2        o715(.A(ori_ori_n737_), .B(ori_ori_n345_), .Y(ori_ori_n738_));
  BUFFER     o716(.A(ori_ori_n240_), .Y(ori_ori_n739_));
  AOI210     o717(.A0(ori_ori_n739_), .A1(ori_ori_n378_), .B0(ori_ori_n568_), .Y(ori_ori_n740_));
  NO2        o718(.A(ori_ori_n740_), .B(ori_ori_n738_), .Y(ori_ori_n741_));
  NO3        o719(.A(ori_ori_n741_), .B(ori_ori_n736_), .C(ori_ori_n732_), .Y(ori_ori_n742_));
  NA2        o720(.A(ori_ori_n173_), .B(ori_ori_n24_), .Y(ori_ori_n743_));
  NO2        o721(.A(ori_ori_n553_), .B(ori_ori_n469_), .Y(ori_ori_n744_));
  NO2        o722(.A(ori_ori_n744_), .B(ori_ori_n743_), .Y(ori_ori_n745_));
  NAi21      o723(.An(ori_ori_n161_), .B(ori_ori_n340_), .Y(ori_ori_n746_));
  NO2        o724(.A(ori_ori_n746_), .B(ori_ori_n717_), .Y(ori_ori_n747_));
  NO2        o725(.A(ori_ori_n747_), .B(ori_ori_n745_), .Y(ori_ori_n748_));
  NA2        o726(.A(ori_ori_n447_), .B(i_0_), .Y(ori_ori_n749_));
  NO3        o727(.A(ori_ori_n749_), .B(ori_ori_n310_), .C(ori_ori_n89_), .Y(ori_ori_n750_));
  NO4        o728(.A(ori_ori_n460_), .B(ori_ori_n197_), .C(ori_ori_n328_), .D(ori_ori_n325_), .Y(ori_ori_n751_));
  AOI210     o729(.A0(ori_ori_n751_), .A1(i_11_), .B0(ori_ori_n750_), .Y(ori_ori_n752_));
  INV        o730(.A(ori_ori_n377_), .Y(ori_ori_n753_));
  NA2        o731(.A(ori_ori_n632_), .B(ori_ori_n264_), .Y(ori_ori_n754_));
  AOI210     o732(.A0(ori_ori_n382_), .A1(ori_ori_n89_), .B0(ori_ori_n58_), .Y(ori_ori_n755_));
  NO2        o733(.A(ori_ori_n755_), .B(ori_ori_n754_), .Y(ori_ori_n756_));
  NO2        o734(.A(ori_ori_n227_), .B(ori_ori_n155_), .Y(ori_ori_n757_));
  NA2        o735(.A(i_0_), .B(i_10_), .Y(ori_ori_n758_));
  INV        o736(.A(ori_ori_n419_), .Y(ori_ori_n759_));
  NO4        o737(.A(ori_ori_n118_), .B(ori_ori_n58_), .C(ori_ori_n548_), .D(i_5_), .Y(ori_ori_n760_));
  AO220      o738(.A0(ori_ori_n760_), .A1(ori_ori_n759_), .B0(ori_ori_n757_), .B1(i_6_), .Y(ori_ori_n761_));
  NO2        o739(.A(ori_ori_n761_), .B(ori_ori_n756_), .Y(ori_ori_n762_));
  NA3        o740(.A(ori_ori_n762_), .B(ori_ori_n752_), .C(ori_ori_n748_), .Y(ori_ori_n763_));
  NO2        o741(.A(ori_ori_n106_), .B(ori_ori_n37_), .Y(ori_ori_n764_));
  NA2        o742(.A(i_11_), .B(i_9_), .Y(ori_ori_n765_));
  NO3        o743(.A(i_12_), .B(ori_ori_n765_), .C(ori_ori_n479_), .Y(ori_ori_n766_));
  AN2        o744(.A(ori_ori_n766_), .B(ori_ori_n764_), .Y(ori_ori_n767_));
  NO2        o745(.A(ori_ori_n48_), .B(i_7_), .Y(ori_ori_n768_));
  NA2        o746(.A(ori_ori_n315_), .B(ori_ori_n170_), .Y(ori_ori_n769_));
  NA3        o747(.A(ori_ori_n769_), .B(ori_ori_n363_), .C(ori_ori_n159_), .Y(ori_ori_n770_));
  NO2        o748(.A(ori_ori_n765_), .B(ori_ori_n73_), .Y(ori_ori_n771_));
  NO2        o749(.A(ori_ori_n168_), .B(i_0_), .Y(ori_ori_n772_));
  INV        o750(.A(ori_ori_n323_), .Y(ori_ori_n773_));
  NO2        o751(.A(ori_ori_n773_), .B(ori_ori_n738_), .Y(ori_ori_n774_));
  NO3        o752(.A(ori_ori_n774_), .B(ori_ori_n770_), .C(ori_ori_n767_), .Y(ori_ori_n775_));
  NA2        o753(.A(ori_ori_n537_), .B(ori_ori_n125_), .Y(ori_ori_n776_));
  NO2        o754(.A(i_6_), .B(ori_ori_n776_), .Y(ori_ori_n777_));
  AOI210     o755(.A0(ori_ori_n348_), .A1(ori_ori_n36_), .B0(i_3_), .Y(ori_ori_n778_));
  NA2        o756(.A(ori_ori_n165_), .B(ori_ori_n106_), .Y(ori_ori_n779_));
  NOi32      o757(.An(ori_ori_n778_), .Bn(ori_ori_n176_), .C(ori_ori_n779_), .Y(ori_ori_n780_));
  NA2        o758(.A(ori_ori_n481_), .B(ori_ori_n264_), .Y(ori_ori_n781_));
  NO2        o759(.A(ori_ori_n781_), .B(ori_ori_n729_), .Y(ori_ori_n782_));
  NO3        o760(.A(ori_ori_n782_), .B(ori_ori_n780_), .C(ori_ori_n777_), .Y(ori_ori_n783_));
  NOi21      o761(.An(i_7_), .B(i_5_), .Y(ori_ori_n784_));
  NOi31      o762(.An(ori_ori_n784_), .B(i_0_), .C(ori_ori_n609_), .Y(ori_ori_n785_));
  NA3        o763(.A(ori_ori_n785_), .B(ori_ori_n309_), .C(i_6_), .Y(ori_ori_n786_));
  BUFFER     o764(.A(ori_ori_n786_), .Y(ori_ori_n787_));
  INV        o765(.A(ori_ori_n261_), .Y(ori_ori_n788_));
  NA3        o766(.A(ori_ori_n787_), .B(ori_ori_n783_), .C(ori_ori_n775_), .Y(ori_ori_n789_));
  NO2        o767(.A(ori_ori_n723_), .B(ori_ori_n260_), .Y(ori_ori_n790_));
  OA210      o768(.A0(ori_ori_n377_), .A1(ori_ori_n206_), .B0(ori_ori_n376_), .Y(ori_ori_n791_));
  NA2        o769(.A(ori_ori_n790_), .B(ori_ori_n771_), .Y(ori_ori_n792_));
  NA3        o770(.A(ori_ori_n376_), .B(ori_ori_n326_), .C(ori_ori_n45_), .Y(ori_ori_n793_));
  OAI210     o771(.A0(ori_ori_n746_), .A1(ori_ori_n753_), .B0(ori_ori_n793_), .Y(ori_ori_n794_));
  NA2        o772(.A(ori_ori_n771_), .B(ori_ori_n255_), .Y(ori_ori_n795_));
  OAI210     o773(.A0(i_2_), .A1(ori_ori_n175_), .B0(ori_ori_n795_), .Y(ori_ori_n796_));
  AOI220     o774(.A0(ori_ori_n796_), .A1(ori_ori_n377_), .B0(ori_ori_n794_), .B1(ori_ori_n73_), .Y(ori_ori_n797_));
  NA3        o775(.A(ori_ori_n700_), .B(ori_ori_n307_), .C(ori_ori_n520_), .Y(ori_ori_n798_));
  NA2        o776(.A(ori_ori_n95_), .B(ori_ori_n44_), .Y(ori_ori_n799_));
  NO2        o777(.A(ori_ori_n75_), .B(ori_ori_n634_), .Y(ori_ori_n800_));
  AOI220     o778(.A0(ori_ori_n800_), .A1(ori_ori_n799_), .B0(ori_ori_n167_), .B1(ori_ori_n469_), .Y(ori_ori_n801_));
  AOI210     o779(.A0(ori_ori_n801_), .A1(ori_ori_n798_), .B0(ori_ori_n47_), .Y(ori_ori_n802_));
  NO3        o780(.A(ori_ori_n460_), .B(ori_ori_n279_), .C(ori_ori_n24_), .Y(ori_ori_n803_));
  AOI210     o781(.A0(ori_ori_n582_), .A1(ori_ori_n426_), .B0(ori_ori_n803_), .Y(ori_ori_n804_));
  NAi21      o782(.An(i_9_), .B(i_5_), .Y(ori_ori_n805_));
  NO2        o783(.A(ori_ori_n805_), .B(ori_ori_n320_), .Y(ori_ori_n806_));
  NA2        o784(.A(ori_ori_n806_), .B(ori_ori_n498_), .Y(ori_ori_n807_));
  OAI220     o785(.A0(ori_ori_n807_), .A1(ori_ori_n86_), .B0(ori_ori_n804_), .B1(ori_ori_n166_), .Y(ori_ori_n808_));
  NO3        o786(.A(ori_ori_n808_), .B(ori_ori_n802_), .C(ori_ori_n411_), .Y(ori_ori_n809_));
  NA3        o787(.A(ori_ori_n809_), .B(ori_ori_n797_), .C(ori_ori_n792_), .Y(ori_ori_n810_));
  NO3        o788(.A(ori_ori_n810_), .B(ori_ori_n789_), .C(ori_ori_n763_), .Y(ori_ori_n811_));
  NO2        o789(.A(i_0_), .B(ori_ori_n609_), .Y(ori_ori_n812_));
  AOI210     o790(.A0(ori_ori_n682_), .A1(ori_ori_n566_), .B0(ori_ori_n779_), .Y(ori_ori_n813_));
  INV        o791(.A(ori_ori_n813_), .Y(ori_ori_n814_));
  OAI210     o792(.A0(ori_ori_n220_), .A1(i_9_), .B0(ori_ori_n212_), .Y(ori_ori_n815_));
  AOI210     o793(.A0(ori_ori_n815_), .A1(ori_ori_n749_), .B0(ori_ori_n155_), .Y(ori_ori_n816_));
  INV        o794(.A(ori_ori_n816_), .Y(ori_ori_n817_));
  NA2        o795(.A(ori_ori_n817_), .B(ori_ori_n814_), .Y(ori_ori_n818_));
  NO3        o796(.A(ori_ori_n758_), .B(ori_ori_n737_), .C(ori_ori_n178_), .Y(ori_ori_n819_));
  AOI220     o797(.A0(ori_ori_n819_), .A1(i_11_), .B0(ori_ori_n445_), .B1(ori_ori_n75_), .Y(ori_ori_n820_));
  NO3        o798(.A(ori_ori_n193_), .B(ori_ori_n308_), .C(i_0_), .Y(ori_ori_n821_));
  OAI210     o799(.A0(ori_ori_n821_), .A1(ori_ori_n76_), .B0(i_13_), .Y(ori_ori_n822_));
  NA2        o800(.A(ori_ori_n822_), .B(ori_ori_n820_), .Y(ori_ori_n823_));
  NO2        o801(.A(ori_ori_n219_), .B(ori_ori_n95_), .Y(ori_ori_n824_));
  AOI210     o802(.A0(ori_ori_n824_), .A1(ori_ori_n812_), .B0(ori_ori_n112_), .Y(ori_ori_n825_));
  OR2        o803(.A(ori_ori_n825_), .B(i_5_), .Y(ori_ori_n826_));
  AOI210     o804(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n168_), .Y(ori_ori_n827_));
  NA2        o805(.A(ori_ori_n827_), .B(ori_ori_n791_), .Y(ori_ori_n828_));
  INV        o806(.A(ori_ori_n424_), .Y(ori_ori_n829_));
  NO3        o807(.A(ori_ori_n729_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n830_));
  NA2        o808(.A(ori_ori_n390_), .B(ori_ori_n383_), .Y(ori_ori_n831_));
  NO3        o809(.A(ori_ori_n831_), .B(ori_ori_n830_), .C(ori_ori_n829_), .Y(ori_ori_n832_));
  NA3        o810(.A(ori_ori_n314_), .B(ori_ori_n165_), .C(ori_ori_n164_), .Y(ori_ori_n833_));
  NA3        o811(.A(ori_ori_n768_), .B(ori_ori_n253_), .C(ori_ori_n212_), .Y(ori_ori_n834_));
  NA2        o812(.A(ori_ori_n834_), .B(ori_ori_n833_), .Y(ori_ori_n835_));
  NO3        o813(.A(ori_ori_n765_), .B(ori_ori_n200_), .C(ori_ori_n178_), .Y(ori_ori_n836_));
  NO2        o814(.A(ori_ori_n836_), .B(ori_ori_n835_), .Y(ori_ori_n837_));
  NA4        o815(.A(ori_ori_n837_), .B(ori_ori_n832_), .C(ori_ori_n828_), .D(ori_ori_n826_), .Y(ori_ori_n838_));
  NO2        o816(.A(ori_ori_n86_), .B(i_5_), .Y(ori_ori_n839_));
  NA3        o817(.A(ori_ori_n724_), .B(ori_ori_n113_), .C(ori_ori_n128_), .Y(ori_ori_n840_));
  INV        o818(.A(ori_ori_n840_), .Y(ori_ori_n841_));
  NA2        o819(.A(ori_ori_n841_), .B(ori_ori_n839_), .Y(ori_ori_n842_));
  NA3        o820(.A(ori_ori_n255_), .B(i_5_), .C(ori_ori_n179_), .Y(ori_ori_n843_));
  NAi31      o821(.An(ori_ori_n218_), .B(ori_ori_n843_), .C(ori_ori_n219_), .Y(ori_ori_n844_));
  NO4        o822(.A(ori_ori_n217_), .B(ori_ori_n193_), .C(i_0_), .D(i_12_), .Y(ori_ori_n845_));
  AOI220     o823(.A0(ori_ori_n845_), .A1(ori_ori_n844_), .B0(ori_ori_n676_), .B1(ori_ori_n169_), .Y(ori_ori_n846_));
  NA2        o824(.A(ori_ori_n784_), .B(ori_ori_n374_), .Y(ori_ori_n847_));
  NA2        o825(.A(ori_ori_n64_), .B(ori_ori_n104_), .Y(ori_ori_n848_));
  OAI220     o826(.A0(ori_ori_n848_), .A1(ori_ori_n843_), .B0(ori_ori_n847_), .B1(ori_ori_n556_), .Y(ori_ori_n849_));
  NA2        o827(.A(ori_ori_n849_), .B(ori_ori_n772_), .Y(ori_ori_n850_));
  NA3        o828(.A(ori_ori_n850_), .B(ori_ori_n846_), .C(ori_ori_n842_), .Y(ori_ori_n851_));
  NO4        o829(.A(ori_ori_n851_), .B(ori_ori_n838_), .C(ori_ori_n823_), .D(ori_ori_n818_), .Y(ori_ori_n852_));
  OAI210     o830(.A0(ori_ori_n699_), .A1(ori_ori_n695_), .B0(ori_ori_n37_), .Y(ori_ori_n853_));
  NA2        o831(.A(ori_ori_n853_), .B(ori_ori_n487_), .Y(ori_ori_n854_));
  NA2        o832(.A(ori_ori_n854_), .B(ori_ori_n191_), .Y(ori_ori_n855_));
  NA2        o833(.A(ori_ori_n174_), .B(ori_ori_n176_), .Y(ori_ori_n856_));
  AO210      o834(.A0(ori_ori_n577_), .A1(ori_ori_n33_), .B0(ori_ori_n856_), .Y(ori_ori_n857_));
  NAi31      o835(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n858_));
  AOI210     o836(.A0(ori_ori_n121_), .A1(ori_ori_n70_), .B0(ori_ori_n858_), .Y(ori_ori_n859_));
  NO2        o837(.A(ori_ori_n859_), .B(ori_ori_n523_), .Y(ori_ori_n860_));
  NA2        o838(.A(ori_ori_n860_), .B(ori_ori_n857_), .Y(ori_ori_n861_));
  NO2        o839(.A(ori_ori_n366_), .B(ori_ori_n240_), .Y(ori_ori_n862_));
  NO2        o840(.A(ori_ori_n862_), .B(ori_ori_n751_), .Y(ori_ori_n863_));
  INV        o841(.A(ori_ori_n863_), .Y(ori_ori_n864_));
  AOI210     o842(.A0(ori_ori_n861_), .A1(ori_ori_n48_), .B0(ori_ori_n864_), .Y(ori_ori_n865_));
  AOI210     o843(.A0(ori_ori_n865_), .A1(ori_ori_n855_), .B0(ori_ori_n73_), .Y(ori_ori_n866_));
  INV        o844(.A(ori_ori_n304_), .Y(ori_ori_n867_));
  NO2        o845(.A(ori_ori_n867_), .B(ori_ori_n640_), .Y(ori_ori_n868_));
  OAI210     o846(.A0(ori_ori_n80_), .A1(ori_ori_n54_), .B0(ori_ori_n111_), .Y(ori_ori_n869_));
  NA2        o847(.A(ori_ori_n869_), .B(ori_ori_n76_), .Y(ori_ori_n870_));
  AOI210     o848(.A0(ori_ori_n827_), .A1(ori_ori_n768_), .B0(ori_ori_n785_), .Y(ori_ori_n871_));
  AOI210     o849(.A0(ori_ori_n871_), .A1(ori_ori_n870_), .B0(ori_ori_n559_), .Y(ori_ori_n872_));
  INV        o850(.A(ori_ori_n872_), .Y(ori_ori_n873_));
  OAI210     o851(.A0(ori_ori_n242_), .A1(ori_ori_n157_), .B0(ori_ori_n89_), .Y(ori_ori_n874_));
  NA3        o852(.A(ori_ori_n644_), .B(ori_ori_n253_), .C(ori_ori_n80_), .Y(ori_ori_n875_));
  AOI210     o853(.A0(ori_ori_n875_), .A1(ori_ori_n874_), .B0(i_11_), .Y(ori_ori_n876_));
  NA2        o854(.A(ori_ori_n482_), .B(ori_ori_n197_), .Y(ori_ori_n877_));
  OAI210     o855(.A0(ori_ori_n877_), .A1(ori_ori_n778_), .B0(ori_ori_n191_), .Y(ori_ori_n878_));
  NA2        o856(.A(ori_ori_n162_), .B(i_5_), .Y(ori_ori_n879_));
  NO2        o857(.A(ori_ori_n878_), .B(ori_ori_n879_), .Y(ori_ori_n880_));
  NO3        o858(.A(ori_ori_n59_), .B(ori_ori_n58_), .C(i_4_), .Y(ori_ori_n881_));
  OAI210     o859(.A0(ori_ori_n788_), .A1(ori_ori_n256_), .B0(ori_ori_n881_), .Y(ori_ori_n882_));
  NO2        o860(.A(ori_ori_n882_), .B(ori_ori_n609_), .Y(ori_ori_n883_));
  NO4        o861(.A(ori_ori_n805_), .B(ori_ori_n379_), .C(ori_ori_n226_), .D(ori_ori_n225_), .Y(ori_ori_n884_));
  NO2        o862(.A(ori_ori_n884_), .B(ori_ori_n442_), .Y(ori_ori_n885_));
  NO2        o863(.A(ori_ori_n697_), .B(ori_ori_n285_), .Y(ori_ori_n886_));
  AOI210     o864(.A0(ori_ori_n886_), .A1(ori_ori_n885_), .B0(ori_ori_n41_), .Y(ori_ori_n887_));
  NO4        o865(.A(ori_ori_n887_), .B(ori_ori_n883_), .C(ori_ori_n880_), .D(ori_ori_n876_), .Y(ori_ori_n888_));
  OAI210     o866(.A0(ori_ori_n873_), .A1(i_4_), .B0(ori_ori_n888_), .Y(ori_ori_n889_));
  NO3        o867(.A(ori_ori_n889_), .B(ori_ori_n868_), .C(ori_ori_n866_), .Y(ori_ori_n890_));
  NA4        o868(.A(ori_ori_n890_), .B(ori_ori_n852_), .C(ori_ori_n811_), .D(ori_ori_n742_), .Y(ori4));
  INV        o869(.A(ori_ori_n581_), .Y(ori_ori_n894_));
  INV        o870(.A(i_6_), .Y(ori_ori_n895_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m0019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m0021(.A(mai_mai_n35_), .Y(mai1));
  INV        m0022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m0023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m0024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m0025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m0026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m0027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m0028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m0029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m0030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m0032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NO2        m0033(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  OAI210     m0034(.A0(mai_mai_n56_), .A1(mai_mai_n53_), .B0(mai_mai_n46_), .Y(mai_mai_n57_));
  NA3        m0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n58_));
  NO2        m0036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NA2        m0037(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  OAI210     m0038(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m0039(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n62_));
  NAi21      m0040(.An(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  INV        m0041(.A(i_1_), .Y(mai_mai_n64_));
  NA2        m0042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NA3        m0043(.A(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m0044(.A(i_1_), .B(i_10_), .Y(mai_mai_n67_));
  NO2        m0045(.A(mai_mai_n67_), .B(i_6_), .Y(mai_mai_n68_));
  NAi31      m0046(.An(mai_mai_n68_), .B(mai_mai_n66_), .C(mai_mai_n62_), .Y(mai_mai_n69_));
  NA2        m0047(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n70_));
  AOI210     m0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n71_));
  NA2        m0049(.A(i_1_), .B(i_6_), .Y(mai_mai_n72_));
  NO2        m0050(.A(mai_mai_n72_), .B(mai_mai_n25_), .Y(mai_mai_n73_));
  INV        m0051(.A(i_0_), .Y(mai_mai_n74_));
  NAi21      m0052(.An(i_5_), .B(i_10_), .Y(mai_mai_n75_));
  NA2        m0053(.A(i_5_), .B(i_9_), .Y(mai_mai_n76_));
  AOI210     m0054(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .Y(mai_mai_n77_));
  NO2        m0055(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OAI210     m0056(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m0057(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(i_0_), .Y(mai_mai_n80_));
  NA2        m0058(.A(i_12_), .B(i_5_), .Y(mai_mai_n81_));
  NA2        m0059(.A(i_2_), .B(i_8_), .Y(mai_mai_n82_));
  NO2        m0060(.A(mai_mai_n82_), .B(mai_mai_n59_), .Y(mai_mai_n83_));
  NO2        m0061(.A(i_3_), .B(i_9_), .Y(mai_mai_n84_));
  NO2        m0062(.A(i_3_), .B(i_7_), .Y(mai_mai_n85_));
  NO3        m0063(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n64_), .Y(mai_mai_n86_));
  INV        m0064(.A(i_6_), .Y(mai_mai_n87_));
  NO2        m0065(.A(i_2_), .B(i_7_), .Y(mai_mai_n88_));
  INV        m0066(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  OAI210     m0067(.A0(mai_mai_n86_), .A1(mai_mai_n83_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NAi21      m0068(.An(i_6_), .B(i_10_), .Y(mai_mai_n91_));
  NA2        m0069(.A(i_6_), .B(i_9_), .Y(mai_mai_n92_));
  AOI210     m0070(.A0(mai_mai_n92_), .A1(mai_mai_n91_), .B0(mai_mai_n64_), .Y(mai_mai_n93_));
  NA2        m0071(.A(i_2_), .B(i_6_), .Y(mai_mai_n94_));
  NO3        m0072(.A(mai_mai_n94_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n95_));
  NO2        m0073(.A(mai_mai_n95_), .B(mai_mai_n93_), .Y(mai_mai_n96_));
  AOI210     m0074(.A0(mai_mai_n96_), .A1(mai_mai_n90_), .B0(mai_mai_n81_), .Y(mai_mai_n97_));
  AN3        m0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n98_));
  NAi21      m0076(.An(i_6_), .B(i_11_), .Y(mai_mai_n99_));
  NO2        m0077(.A(i_5_), .B(i_8_), .Y(mai_mai_n100_));
  NOi21      m0078(.An(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  AOI220     m0079(.A0(mai_mai_n101_), .A1(mai_mai_n63_), .B0(mai_mai_n98_), .B1(mai_mai_n32_), .Y(mai_mai_n102_));
  INV        m0080(.A(i_7_), .Y(mai_mai_n103_));
  NA2        m0081(.A(mai_mai_n47_), .B(mai_mai_n103_), .Y(mai_mai_n104_));
  NO2        m0082(.A(i_0_), .B(i_5_), .Y(mai_mai_n105_));
  NO2        m0083(.A(mai_mai_n105_), .B(mai_mai_n87_), .Y(mai_mai_n106_));
  NA2        m0084(.A(i_12_), .B(i_3_), .Y(mai_mai_n107_));
  INV        m0085(.A(mai_mai_n107_), .Y(mai_mai_n108_));
  NA3        m0086(.A(mai_mai_n108_), .B(mai_mai_n106_), .C(mai_mai_n104_), .Y(mai_mai_n109_));
  NAi21      m0087(.An(i_7_), .B(i_11_), .Y(mai_mai_n110_));
  AN2        m0088(.A(i_2_), .B(i_10_), .Y(mai_mai_n111_));
  NO2        m0089(.A(mai_mai_n111_), .B(i_7_), .Y(mai_mai_n112_));
  OR2        m0090(.A(mai_mai_n81_), .B(mai_mai_n59_), .Y(mai_mai_n113_));
  NO2        m0091(.A(i_8_), .B(mai_mai_n103_), .Y(mai_mai_n114_));
  NO3        m0092(.A(mai_mai_n114_), .B(mai_mai_n113_), .C(mai_mai_n112_), .Y(mai_mai_n115_));
  NA2        m0093(.A(i_12_), .B(i_7_), .Y(mai_mai_n116_));
  NO2        m0094(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n117_));
  NA2        m0095(.A(mai_mai_n117_), .B(i_0_), .Y(mai_mai_n118_));
  NA2        m0096(.A(i_11_), .B(i_12_), .Y(mai_mai_n119_));
  OAI210     m0097(.A0(mai_mai_n118_), .A1(mai_mai_n116_), .B0(mai_mai_n119_), .Y(mai_mai_n120_));
  NO2        m0098(.A(mai_mai_n120_), .B(mai_mai_n115_), .Y(mai_mai_n121_));
  NA3        m0099(.A(mai_mai_n121_), .B(mai_mai_n109_), .C(mai_mai_n102_), .Y(mai_mai_n122_));
  NOi21      m0100(.An(i_1_), .B(i_5_), .Y(mai_mai_n123_));
  NA2        m0101(.A(mai_mai_n123_), .B(i_11_), .Y(mai_mai_n124_));
  NA2        m0102(.A(mai_mai_n103_), .B(mai_mai_n37_), .Y(mai_mai_n125_));
  NA2        m0103(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n126_));
  NA2        m0104(.A(mai_mai_n126_), .B(mai_mai_n125_), .Y(mai_mai_n127_));
  NO2        m0105(.A(mai_mai_n127_), .B(mai_mai_n47_), .Y(mai_mai_n128_));
  NA2        m0106(.A(mai_mai_n92_), .B(mai_mai_n91_), .Y(mai_mai_n129_));
  NAi21      m0107(.An(i_3_), .B(i_8_), .Y(mai_mai_n130_));
  NA2        m0108(.A(mai_mai_n130_), .B(mai_mai_n63_), .Y(mai_mai_n131_));
  NOi31      m0109(.An(mai_mai_n131_), .B(mai_mai_n129_), .C(mai_mai_n128_), .Y(mai_mai_n132_));
  NO2        m0110(.A(i_1_), .B(mai_mai_n87_), .Y(mai_mai_n133_));
  NO2        m0111(.A(i_6_), .B(i_5_), .Y(mai_mai_n134_));
  NA2        m0112(.A(mai_mai_n134_), .B(i_3_), .Y(mai_mai_n135_));
  AO210      m0113(.A0(mai_mai_n135_), .A1(mai_mai_n48_), .B0(mai_mai_n133_), .Y(mai_mai_n136_));
  OAI220     m0114(.A0(mai_mai_n136_), .A1(mai_mai_n110_), .B0(mai_mai_n132_), .B1(mai_mai_n124_), .Y(mai_mai_n137_));
  NO3        m0115(.A(mai_mai_n137_), .B(mai_mai_n122_), .C(mai_mai_n97_), .Y(mai_mai_n138_));
  NA3        m0116(.A(mai_mai_n138_), .B(mai_mai_n80_), .C(mai_mai_n57_), .Y(mai2));
  NO2        m0117(.A(mai_mai_n64_), .B(mai_mai_n37_), .Y(mai_mai_n140_));
  NA2        m0118(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n141_));
  NA2        m0119(.A(mai_mai_n141_), .B(mai_mai_n140_), .Y(mai_mai_n142_));
  NA4        m0120(.A(mai_mai_n142_), .B(mai_mai_n78_), .C(mai_mai_n70_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0121(.A(i_8_), .B(i_7_), .Y(mai_mai_n144_));
  NA2        m0122(.A(mai_mai_n144_), .B(i_6_), .Y(mai_mai_n145_));
  NO2        m0123(.A(i_12_), .B(i_13_), .Y(mai_mai_n146_));
  NAi21      m0124(.An(i_5_), .B(i_11_), .Y(mai_mai_n147_));
  NOi21      m0125(.An(mai_mai_n146_), .B(mai_mai_n147_), .Y(mai_mai_n148_));
  NO2        m0126(.A(i_0_), .B(i_1_), .Y(mai_mai_n149_));
  NA2        m0127(.A(i_2_), .B(i_3_), .Y(mai_mai_n150_));
  NO2        m0128(.A(mai_mai_n150_), .B(i_4_), .Y(mai_mai_n151_));
  NA3        m0129(.A(mai_mai_n151_), .B(mai_mai_n149_), .C(mai_mai_n148_), .Y(mai_mai_n152_));
  AN2        m0130(.A(mai_mai_n146_), .B(mai_mai_n84_), .Y(mai_mai_n153_));
  NO2        m0131(.A(mai_mai_n153_), .B(mai_mai_n27_), .Y(mai_mai_n154_));
  NA2        m0132(.A(i_1_), .B(i_5_), .Y(mai_mai_n155_));
  NO2        m0133(.A(mai_mai_n74_), .B(mai_mai_n47_), .Y(mai_mai_n156_));
  NA2        m0134(.A(mai_mai_n156_), .B(mai_mai_n36_), .Y(mai_mai_n157_));
  NO3        m0135(.A(mai_mai_n157_), .B(mai_mai_n155_), .C(mai_mai_n154_), .Y(mai_mai_n158_));
  OR2        m0136(.A(i_0_), .B(i_1_), .Y(mai_mai_n159_));
  NO3        m0137(.A(mai_mai_n159_), .B(mai_mai_n81_), .C(i_13_), .Y(mai_mai_n160_));
  NAi32      m0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n161_));
  NAi21      m0139(.An(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  NOi21      m0140(.An(i_4_), .B(i_10_), .Y(mai_mai_n163_));
  NA2        m0141(.A(mai_mai_n163_), .B(mai_mai_n40_), .Y(mai_mai_n164_));
  NO2        m0142(.A(i_3_), .B(i_5_), .Y(mai_mai_n165_));
  NO3        m0143(.A(mai_mai_n74_), .B(i_2_), .C(i_1_), .Y(mai_mai_n166_));
  NA2        m0144(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  OAI210     m0145(.A0(mai_mai_n167_), .A1(mai_mai_n164_), .B0(mai_mai_n162_), .Y(mai_mai_n168_));
  NO2        m0146(.A(mai_mai_n168_), .B(mai_mai_n158_), .Y(mai_mai_n169_));
  AOI210     m0147(.A0(mai_mai_n169_), .A1(mai_mai_n152_), .B0(mai_mai_n145_), .Y(mai_mai_n170_));
  NA3        m0148(.A(mai_mai_n74_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n171_));
  NA2        m0149(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n172_));
  NOi21      m0150(.An(i_4_), .B(i_9_), .Y(mai_mai_n173_));
  NOi21      m0151(.An(i_11_), .B(i_13_), .Y(mai_mai_n174_));
  NA2        m0152(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  OR2        m0153(.A(mai_mai_n175_), .B(mai_mai_n172_), .Y(mai_mai_n176_));
  NO2        m0154(.A(i_4_), .B(i_5_), .Y(mai_mai_n177_));
  NAi21      m0155(.An(i_12_), .B(i_11_), .Y(mai_mai_n178_));
  NO2        m0156(.A(mai_mai_n178_), .B(i_13_), .Y(mai_mai_n179_));
  NA3        m0157(.A(mai_mai_n179_), .B(mai_mai_n177_), .C(mai_mai_n84_), .Y(mai_mai_n180_));
  AOI210     m0158(.A0(mai_mai_n180_), .A1(mai_mai_n176_), .B0(mai_mai_n171_), .Y(mai_mai_n181_));
  NO2        m0159(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n182_));
  NA2        m0160(.A(mai_mai_n182_), .B(mai_mai_n47_), .Y(mai_mai_n183_));
  NA2        m0161(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n184_));
  NAi31      m0162(.An(mai_mai_n184_), .B(mai_mai_n153_), .C(i_11_), .Y(mai_mai_n185_));
  NA2        m0163(.A(i_3_), .B(i_5_), .Y(mai_mai_n186_));
  OR2        m0164(.A(mai_mai_n186_), .B(mai_mai_n175_), .Y(mai_mai_n187_));
  AOI210     m0165(.A0(mai_mai_n187_), .A1(mai_mai_n185_), .B0(mai_mai_n183_), .Y(mai_mai_n188_));
  NO2        m0166(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n189_));
  NO2        m0167(.A(i_13_), .B(i_10_), .Y(mai_mai_n190_));
  NA3        m0168(.A(mai_mai_n190_), .B(mai_mai_n189_), .C(mai_mai_n45_), .Y(mai_mai_n191_));
  NO2        m0169(.A(i_2_), .B(i_1_), .Y(mai_mai_n192_));
  NA2        m0170(.A(mai_mai_n192_), .B(i_3_), .Y(mai_mai_n193_));
  NAi21      m0171(.An(i_4_), .B(i_12_), .Y(mai_mai_n194_));
  NO4        m0172(.A(mai_mai_n194_), .B(mai_mai_n193_), .C(mai_mai_n191_), .D(mai_mai_n25_), .Y(mai_mai_n195_));
  NO3        m0173(.A(mai_mai_n195_), .B(mai_mai_n188_), .C(mai_mai_n181_), .Y(mai_mai_n196_));
  INV        m0174(.A(i_8_), .Y(mai_mai_n197_));
  NO2        m0175(.A(mai_mai_n197_), .B(i_7_), .Y(mai_mai_n198_));
  NA2        m0176(.A(mai_mai_n198_), .B(i_6_), .Y(mai_mai_n199_));
  NO3        m0177(.A(i_3_), .B(mai_mai_n87_), .C(mai_mai_n49_), .Y(mai_mai_n200_));
  NA2        m0178(.A(mai_mai_n200_), .B(mai_mai_n114_), .Y(mai_mai_n201_));
  NO3        m0179(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n202_));
  NA3        m0180(.A(mai_mai_n202_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n203_));
  NO3        m0181(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n204_));
  OAI210     m0182(.A0(mai_mai_n98_), .A1(i_12_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  AOI210     m0183(.A0(mai_mai_n205_), .A1(mai_mai_n203_), .B0(mai_mai_n201_), .Y(mai_mai_n206_));
  NO2        m0184(.A(i_3_), .B(i_8_), .Y(mai_mai_n207_));
  NO3        m0185(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n208_));
  NO2        m0186(.A(mai_mai_n105_), .B(mai_mai_n59_), .Y(mai_mai_n209_));
  NO2        m0187(.A(i_13_), .B(i_9_), .Y(mai_mai_n210_));
  NA3        m0188(.A(mai_mai_n210_), .B(i_6_), .C(mai_mai_n197_), .Y(mai_mai_n211_));
  NAi21      m0189(.An(i_12_), .B(i_3_), .Y(mai_mai_n212_));
  NO2        m0190(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n213_));
  NO3        m0191(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n214_));
  NA3        m0192(.A(mai_mai_n214_), .B(mai_mai_n213_), .C(i_10_), .Y(mai_mai_n215_));
  NO2        m0193(.A(mai_mai_n215_), .B(mai_mai_n211_), .Y(mai_mai_n216_));
  AOI210     m0194(.A0(mai_mai_n216_), .A1(i_7_), .B0(mai_mai_n206_), .Y(mai_mai_n217_));
  OAI220     m0195(.A0(mai_mai_n217_), .A1(i_4_), .B0(mai_mai_n199_), .B1(mai_mai_n196_), .Y(mai_mai_n218_));
  NAi21      m0196(.An(i_12_), .B(i_7_), .Y(mai_mai_n219_));
  NA3        m0197(.A(i_13_), .B(mai_mai_n197_), .C(i_10_), .Y(mai_mai_n220_));
  NA2        m0198(.A(i_0_), .B(i_5_), .Y(mai_mai_n221_));
  NAi31      m0199(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n222_));
  NO2        m0200(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n223_));
  NO2        m0201(.A(mai_mai_n74_), .B(mai_mai_n26_), .Y(mai_mai_n224_));
  NO2        m0202(.A(mai_mai_n47_), .B(mai_mai_n64_), .Y(mai_mai_n225_));
  NA3        m0203(.A(mai_mai_n225_), .B(mai_mai_n224_), .C(mai_mai_n223_), .Y(mai_mai_n226_));
  INV        m0204(.A(i_13_), .Y(mai_mai_n227_));
  NO2        m0205(.A(i_12_), .B(mai_mai_n227_), .Y(mai_mai_n228_));
  NO2        m0206(.A(mai_mai_n226_), .B(mai_mai_n222_), .Y(mai_mai_n229_));
  NA2        m0207(.A(mai_mai_n229_), .B(mai_mai_n144_), .Y(mai_mai_n230_));
  NO2        m0208(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n231_));
  NO2        m0209(.A(mai_mai_n186_), .B(i_4_), .Y(mai_mai_n232_));
  NA2        m0210(.A(mai_mai_n232_), .B(mai_mai_n231_), .Y(mai_mai_n233_));
  OR2        m0211(.A(i_8_), .B(i_7_), .Y(mai_mai_n234_));
  NO2        m0212(.A(mai_mai_n234_), .B(mai_mai_n87_), .Y(mai_mai_n235_));
  NO2        m0213(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n236_));
  NA2        m0214(.A(mai_mai_n236_), .B(mai_mai_n235_), .Y(mai_mai_n237_));
  INV        m0215(.A(i_12_), .Y(mai_mai_n238_));
  NO2        m0216(.A(mai_mai_n45_), .B(mai_mai_n238_), .Y(mai_mai_n239_));
  NO3        m0217(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n240_));
  NA2        m0218(.A(i_2_), .B(i_1_), .Y(mai_mai_n241_));
  NO2        m0219(.A(mai_mai_n237_), .B(mai_mai_n233_), .Y(mai_mai_n242_));
  NO3        m0220(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n243_));
  NAi21      m0221(.An(i_4_), .B(i_3_), .Y(mai_mai_n244_));
  NO2        m0222(.A(mai_mai_n244_), .B(mai_mai_n76_), .Y(mai_mai_n245_));
  NO2        m0223(.A(i_0_), .B(i_6_), .Y(mai_mai_n246_));
  NOi41      m0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n247_));
  NA2        m0225(.A(mai_mai_n247_), .B(mai_mai_n246_), .Y(mai_mai_n248_));
  NO2        m0226(.A(mai_mai_n241_), .B(mai_mai_n186_), .Y(mai_mai_n249_));
  NAi21      m0227(.An(mai_mai_n248_), .B(mai_mai_n249_), .Y(mai_mai_n250_));
  INV        m0228(.A(mai_mai_n250_), .Y(mai_mai_n251_));
  AOI220     m0229(.A0(mai_mai_n251_), .A1(mai_mai_n40_), .B0(mai_mai_n242_), .B1(mai_mai_n210_), .Y(mai_mai_n252_));
  NO2        m0230(.A(i_11_), .B(mai_mai_n227_), .Y(mai_mai_n253_));
  NOi21      m0231(.An(i_1_), .B(i_6_), .Y(mai_mai_n254_));
  NAi21      m0232(.An(i_3_), .B(i_7_), .Y(mai_mai_n255_));
  NA2        m0233(.A(mai_mai_n238_), .B(i_9_), .Y(mai_mai_n256_));
  OR4        m0234(.A(mai_mai_n256_), .B(mai_mai_n255_), .C(mai_mai_n254_), .D(mai_mai_n189_), .Y(mai_mai_n257_));
  NO2        m0235(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n258_));
  NO2        m0236(.A(i_12_), .B(i_3_), .Y(mai_mai_n259_));
  NA2        m0237(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n260_));
  NA2        m0238(.A(i_3_), .B(i_9_), .Y(mai_mai_n261_));
  NAi21      m0239(.An(i_7_), .B(i_10_), .Y(mai_mai_n262_));
  NO2        m0240(.A(mai_mai_n262_), .B(mai_mai_n261_), .Y(mai_mai_n263_));
  NA3        m0241(.A(mai_mai_n263_), .B(mai_mai_n260_), .C(mai_mai_n65_), .Y(mai_mai_n264_));
  NA2        m0242(.A(mai_mai_n264_), .B(mai_mai_n257_), .Y(mai_mai_n265_));
  NA3        m0243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n266_));
  INV        m0244(.A(mai_mai_n145_), .Y(mai_mai_n267_));
  NA2        m0245(.A(mai_mai_n238_), .B(i_13_), .Y(mai_mai_n268_));
  NO2        m0246(.A(mai_mai_n268_), .B(mai_mai_n76_), .Y(mai_mai_n269_));
  AOI220     m0247(.A0(mai_mai_n269_), .A1(mai_mai_n267_), .B0(mai_mai_n265_), .B1(mai_mai_n253_), .Y(mai_mai_n270_));
  NO2        m0248(.A(mai_mai_n234_), .B(mai_mai_n37_), .Y(mai_mai_n271_));
  NA2        m0249(.A(i_12_), .B(i_6_), .Y(mai_mai_n272_));
  OR2        m0250(.A(i_13_), .B(i_9_), .Y(mai_mai_n273_));
  NO3        m0251(.A(mai_mai_n273_), .B(mai_mai_n272_), .C(mai_mai_n49_), .Y(mai_mai_n274_));
  NO2        m0252(.A(mai_mai_n244_), .B(i_2_), .Y(mai_mai_n275_));
  NA2        m0253(.A(mai_mai_n253_), .B(i_9_), .Y(mai_mai_n276_));
  NA2        m0254(.A(mai_mai_n156_), .B(mai_mai_n64_), .Y(mai_mai_n277_));
  NO3        m0255(.A(i_11_), .B(mai_mai_n227_), .C(mai_mai_n25_), .Y(mai_mai_n278_));
  NO2        m0256(.A(mai_mai_n255_), .B(i_8_), .Y(mai_mai_n279_));
  NO2        m0257(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n280_));
  NA3        m0258(.A(mai_mai_n280_), .B(mai_mai_n279_), .C(mai_mai_n278_), .Y(mai_mai_n281_));
  NO3        m0259(.A(mai_mai_n26_), .B(mai_mai_n87_), .C(i_5_), .Y(mai_mai_n282_));
  NA3        m0260(.A(mai_mai_n282_), .B(mai_mai_n271_), .C(mai_mai_n228_), .Y(mai_mai_n283_));
  AOI210     m0261(.A0(mai_mai_n283_), .A1(mai_mai_n281_), .B0(mai_mai_n277_), .Y(mai_mai_n284_));
  INV        m0262(.A(mai_mai_n284_), .Y(mai_mai_n285_));
  NA4        m0263(.A(mai_mai_n285_), .B(mai_mai_n270_), .C(mai_mai_n252_), .D(mai_mai_n230_), .Y(mai_mai_n286_));
  NO3        m0264(.A(i_12_), .B(mai_mai_n227_), .C(mai_mai_n37_), .Y(mai_mai_n287_));
  INV        m0265(.A(mai_mai_n287_), .Y(mai_mai_n288_));
  NA2        m0266(.A(i_8_), .B(mai_mai_n103_), .Y(mai_mai_n289_));
  NOi21      m0267(.An(mai_mai_n165_), .B(mai_mai_n87_), .Y(mai_mai_n290_));
  NO3        m0268(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n291_));
  AOI220     m0269(.A0(mai_mai_n291_), .A1(mai_mai_n200_), .B0(mai_mai_n290_), .B1(mai_mai_n236_), .Y(mai_mai_n292_));
  NO2        m0270(.A(mai_mai_n292_), .B(mai_mai_n289_), .Y(mai_mai_n293_));
  NO3        m0271(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n294_));
  NO2        m0272(.A(mai_mai_n241_), .B(i_0_), .Y(mai_mai_n295_));
  AOI220     m0273(.A0(mai_mai_n295_), .A1(mai_mai_n198_), .B0(mai_mai_n294_), .B1(mai_mai_n144_), .Y(mai_mai_n296_));
  NA2        m0274(.A(mai_mai_n280_), .B(mai_mai_n26_), .Y(mai_mai_n297_));
  NO2        m0275(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n298_));
  NA2        m0276(.A(i_0_), .B(i_1_), .Y(mai_mai_n299_));
  NO2        m0277(.A(mai_mai_n299_), .B(i_2_), .Y(mai_mai_n300_));
  NO2        m0278(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n301_));
  NA3        m0279(.A(mai_mai_n301_), .B(mai_mai_n300_), .C(mai_mai_n165_), .Y(mai_mai_n302_));
  OAI210     m0280(.A0(mai_mai_n167_), .A1(mai_mai_n145_), .B0(mai_mai_n302_), .Y(mai_mai_n303_));
  NO3        m0281(.A(mai_mai_n303_), .B(mai_mai_n298_), .C(mai_mai_n293_), .Y(mai_mai_n304_));
  NO2        m0282(.A(i_3_), .B(i_10_), .Y(mai_mai_n305_));
  NA3        m0283(.A(mai_mai_n305_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n306_));
  NO2        m0284(.A(i_2_), .B(mai_mai_n103_), .Y(mai_mai_n307_));
  NA2        m0285(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n308_));
  NO2        m0286(.A(mai_mai_n308_), .B(i_8_), .Y(mai_mai_n309_));
  NA2        m0287(.A(mai_mai_n309_), .B(mai_mai_n307_), .Y(mai_mai_n310_));
  AN2        m0288(.A(i_3_), .B(i_10_), .Y(mai_mai_n311_));
  NA4        m0289(.A(mai_mai_n311_), .B(mai_mai_n202_), .C(mai_mai_n179_), .D(mai_mai_n177_), .Y(mai_mai_n312_));
  NO2        m0290(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n313_));
  NO2        m0291(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n314_));
  OR2        m0292(.A(mai_mai_n310_), .B(mai_mai_n306_), .Y(mai_mai_n315_));
  OAI220     m0293(.A0(mai_mai_n315_), .A1(i_6_), .B0(mai_mai_n304_), .B1(mai_mai_n288_), .Y(mai_mai_n316_));
  NO4        m0294(.A(mai_mai_n316_), .B(mai_mai_n286_), .C(mai_mai_n218_), .D(mai_mai_n170_), .Y(mai_mai_n317_));
  NO3        m0295(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n318_));
  NO2        m0296(.A(mai_mai_n60_), .B(mai_mai_n87_), .Y(mai_mai_n319_));
  NA2        m0297(.A(mai_mai_n295_), .B(mai_mai_n319_), .Y(mai_mai_n320_));
  NO3        m0298(.A(i_6_), .B(mai_mai_n197_), .C(i_7_), .Y(mai_mai_n321_));
  NA2        m0299(.A(mai_mai_n321_), .B(mai_mai_n202_), .Y(mai_mai_n322_));
  AOI210     m0300(.A0(mai_mai_n322_), .A1(mai_mai_n320_), .B0(mai_mai_n172_), .Y(mai_mai_n323_));
  NO2        m0301(.A(i_2_), .B(i_3_), .Y(mai_mai_n324_));
  OR2        m0302(.A(i_0_), .B(i_5_), .Y(mai_mai_n325_));
  NA2        m0303(.A(mai_mai_n221_), .B(mai_mai_n325_), .Y(mai_mai_n326_));
  NA4        m0304(.A(mai_mai_n326_), .B(mai_mai_n235_), .C(mai_mai_n324_), .D(i_1_), .Y(mai_mai_n327_));
  NA3        m0305(.A(mai_mai_n295_), .B(mai_mai_n290_), .C(mai_mai_n114_), .Y(mai_mai_n328_));
  NAi21      m0306(.An(i_8_), .B(i_7_), .Y(mai_mai_n329_));
  NO2        m0307(.A(mai_mai_n329_), .B(i_6_), .Y(mai_mai_n330_));
  NO2        m0308(.A(mai_mai_n159_), .B(mai_mai_n47_), .Y(mai_mai_n331_));
  NA3        m0309(.A(mai_mai_n331_), .B(mai_mai_n330_), .C(mai_mai_n165_), .Y(mai_mai_n332_));
  NA3        m0310(.A(mai_mai_n332_), .B(mai_mai_n328_), .C(mai_mai_n327_), .Y(mai_mai_n333_));
  OAI210     m0311(.A0(mai_mai_n333_), .A1(mai_mai_n323_), .B0(i_4_), .Y(mai_mai_n334_));
  NO2        m0312(.A(i_12_), .B(i_10_), .Y(mai_mai_n335_));
  NOi21      m0313(.An(i_5_), .B(i_0_), .Y(mai_mai_n336_));
  AOI210     m0314(.A0(i_2_), .A1(mai_mai_n49_), .B0(mai_mai_n103_), .Y(mai_mai_n337_));
  NO4        m0315(.A(mai_mai_n337_), .B(mai_mai_n308_), .C(mai_mai_n336_), .D(mai_mai_n130_), .Y(mai_mai_n338_));
  NA4        m0316(.A(mai_mai_n85_), .B(mai_mai_n36_), .C(mai_mai_n87_), .D(i_8_), .Y(mai_mai_n339_));
  NA2        m0317(.A(mai_mai_n338_), .B(mai_mai_n335_), .Y(mai_mai_n340_));
  NO2        m0318(.A(i_6_), .B(i_8_), .Y(mai_mai_n341_));
  NOi21      m0319(.An(i_0_), .B(i_2_), .Y(mai_mai_n342_));
  AN2        m0320(.A(mai_mai_n342_), .B(mai_mai_n341_), .Y(mai_mai_n343_));
  NO2        m0321(.A(i_1_), .B(i_7_), .Y(mai_mai_n344_));
  AO220      m0322(.A0(mai_mai_n344_), .A1(mai_mai_n343_), .B0(mai_mai_n330_), .B1(mai_mai_n236_), .Y(mai_mai_n345_));
  NA3        m0323(.A(mai_mai_n345_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n346_));
  NA3        m0324(.A(mai_mai_n346_), .B(mai_mai_n340_), .C(mai_mai_n334_), .Y(mai_mai_n347_));
  NO3        m0325(.A(mai_mai_n234_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n348_));
  NO3        m0326(.A(mai_mai_n329_), .B(i_2_), .C(i_1_), .Y(mai_mai_n349_));
  OAI210     m0327(.A0(mai_mai_n349_), .A1(mai_mai_n348_), .B0(i_6_), .Y(mai_mai_n350_));
  NA3        m0328(.A(mai_mai_n254_), .B(mai_mai_n307_), .C(mai_mai_n197_), .Y(mai_mai_n351_));
  AOI210     m0329(.A0(mai_mai_n351_), .A1(mai_mai_n350_), .B0(mai_mai_n326_), .Y(mai_mai_n352_));
  NOi21      m0330(.An(mai_mai_n155_), .B(mai_mai_n106_), .Y(mai_mai_n353_));
  NO2        m0331(.A(mai_mai_n353_), .B(mai_mai_n126_), .Y(mai_mai_n354_));
  OAI210     m0332(.A0(mai_mai_n354_), .A1(mai_mai_n352_), .B0(i_3_), .Y(mai_mai_n355_));
  INV        m0333(.A(mai_mai_n85_), .Y(mai_mai_n356_));
  NO2        m0334(.A(mai_mai_n299_), .B(mai_mai_n82_), .Y(mai_mai_n357_));
  NA2        m0335(.A(mai_mai_n357_), .B(mai_mai_n134_), .Y(mai_mai_n358_));
  NO2        m0336(.A(mai_mai_n94_), .B(mai_mai_n197_), .Y(mai_mai_n359_));
  NA2        m0337(.A(mai_mai_n359_), .B(mai_mai_n64_), .Y(mai_mai_n360_));
  AOI210     m0338(.A0(mai_mai_n360_), .A1(mai_mai_n358_), .B0(mai_mai_n356_), .Y(mai_mai_n361_));
  NO2        m0339(.A(mai_mai_n197_), .B(i_9_), .Y(mai_mai_n362_));
  NA3        m0340(.A(mai_mai_n362_), .B(mai_mai_n209_), .C(mai_mai_n159_), .Y(mai_mai_n363_));
  NO2        m0341(.A(mai_mai_n363_), .B(mai_mai_n47_), .Y(mai_mai_n364_));
  NO3        m0342(.A(mai_mai_n364_), .B(mai_mai_n361_), .C(mai_mai_n298_), .Y(mai_mai_n365_));
  AOI210     m0343(.A0(mai_mai_n365_), .A1(mai_mai_n355_), .B0(mai_mai_n164_), .Y(mai_mai_n366_));
  AOI210     m0344(.A0(mai_mai_n347_), .A1(mai_mai_n318_), .B0(mai_mai_n366_), .Y(mai_mai_n367_));
  NOi32      m0345(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n368_));
  INV        m0346(.A(mai_mai_n368_), .Y(mai_mai_n369_));
  NAi21      m0347(.An(i_0_), .B(i_6_), .Y(mai_mai_n370_));
  NAi21      m0348(.An(i_1_), .B(i_5_), .Y(mai_mai_n371_));
  NA2        m0349(.A(mai_mai_n371_), .B(mai_mai_n370_), .Y(mai_mai_n372_));
  INV        m0350(.A(mai_mai_n248_), .Y(mai_mai_n373_));
  NAi41      m0351(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n374_));
  OAI220     m0352(.A0(mai_mai_n374_), .A1(mai_mai_n371_), .B0(mai_mai_n222_), .B1(mai_mai_n161_), .Y(mai_mai_n375_));
  AOI210     m0353(.A0(mai_mai_n374_), .A1(mai_mai_n161_), .B0(mai_mai_n159_), .Y(mai_mai_n376_));
  NOi32      m0354(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n377_));
  NAi21      m0355(.An(i_6_), .B(i_1_), .Y(mai_mai_n378_));
  NA3        m0356(.A(mai_mai_n378_), .B(mai_mai_n377_), .C(mai_mai_n47_), .Y(mai_mai_n379_));
  NO2        m0357(.A(mai_mai_n379_), .B(i_0_), .Y(mai_mai_n380_));
  OR3        m0358(.A(mai_mai_n380_), .B(mai_mai_n376_), .C(mai_mai_n375_), .Y(mai_mai_n381_));
  NO2        m0359(.A(i_1_), .B(mai_mai_n103_), .Y(mai_mai_n382_));
  NAi21      m0360(.An(i_3_), .B(i_4_), .Y(mai_mai_n383_));
  NO2        m0361(.A(mai_mai_n383_), .B(i_9_), .Y(mai_mai_n384_));
  AN2        m0362(.A(i_6_), .B(i_7_), .Y(mai_mai_n385_));
  OAI210     m0363(.A0(mai_mai_n385_), .A1(mai_mai_n382_), .B0(mai_mai_n384_), .Y(mai_mai_n386_));
  NA2        m0364(.A(i_2_), .B(i_7_), .Y(mai_mai_n387_));
  NO2        m0365(.A(mai_mai_n383_), .B(i_10_), .Y(mai_mai_n388_));
  NA3        m0366(.A(mai_mai_n388_), .B(mai_mai_n387_), .C(mai_mai_n246_), .Y(mai_mai_n389_));
  AOI210     m0367(.A0(mai_mai_n389_), .A1(mai_mai_n386_), .B0(mai_mai_n189_), .Y(mai_mai_n390_));
  AOI210     m0368(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n391_));
  OAI210     m0369(.A0(mai_mai_n391_), .A1(mai_mai_n192_), .B0(mai_mai_n388_), .Y(mai_mai_n392_));
  AOI220     m0370(.A0(mai_mai_n388_), .A1(mai_mai_n344_), .B0(mai_mai_n240_), .B1(mai_mai_n192_), .Y(mai_mai_n393_));
  AOI210     m0371(.A0(mai_mai_n393_), .A1(mai_mai_n392_), .B0(i_5_), .Y(mai_mai_n394_));
  NO4        m0372(.A(mai_mai_n394_), .B(mai_mai_n390_), .C(mai_mai_n381_), .D(mai_mai_n373_), .Y(mai_mai_n395_));
  NO2        m0373(.A(mai_mai_n395_), .B(mai_mai_n369_), .Y(mai_mai_n396_));
  NO2        m0374(.A(mai_mai_n60_), .B(mai_mai_n25_), .Y(mai_mai_n397_));
  AN2        m0375(.A(i_12_), .B(i_5_), .Y(mai_mai_n398_));
  NA2        m0376(.A(i_3_), .B(mai_mai_n398_), .Y(mai_mai_n399_));
  NO2        m0377(.A(i_11_), .B(i_6_), .Y(mai_mai_n400_));
  NA3        m0378(.A(mai_mai_n400_), .B(mai_mai_n331_), .C(mai_mai_n227_), .Y(mai_mai_n401_));
  NO2        m0379(.A(mai_mai_n401_), .B(mai_mai_n399_), .Y(mai_mai_n402_));
  NO2        m0380(.A(mai_mai_n244_), .B(i_5_), .Y(mai_mai_n403_));
  NO2        m0381(.A(i_5_), .B(i_10_), .Y(mai_mai_n404_));
  AOI220     m0382(.A0(mai_mai_n404_), .A1(mai_mai_n275_), .B0(mai_mai_n403_), .B1(mai_mai_n202_), .Y(mai_mai_n405_));
  NA2        m0383(.A(mai_mai_n146_), .B(mai_mai_n46_), .Y(mai_mai_n406_));
  NO2        m0384(.A(mai_mai_n406_), .B(mai_mai_n405_), .Y(mai_mai_n407_));
  OAI210     m0385(.A0(mai_mai_n407_), .A1(mai_mai_n402_), .B0(mai_mai_n397_), .Y(mai_mai_n408_));
  NO2        m0386(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n409_));
  NO3        m0387(.A(mai_mai_n87_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n410_));
  NO2        m0388(.A(i_3_), .B(mai_mai_n103_), .Y(mai_mai_n411_));
  NO2        m0389(.A(i_11_), .B(i_12_), .Y(mai_mai_n412_));
  NA2        m0390(.A(mai_mai_n404_), .B(mai_mai_n238_), .Y(mai_mai_n413_));
  NA3        m0391(.A(mai_mai_n114_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n414_));
  OAI220     m0392(.A0(mai_mai_n414_), .A1(mai_mai_n222_), .B0(mai_mai_n413_), .B1(mai_mai_n339_), .Y(mai_mai_n415_));
  NAi21      m0393(.An(i_13_), .B(i_0_), .Y(mai_mai_n416_));
  NO2        m0394(.A(mai_mai_n416_), .B(mai_mai_n241_), .Y(mai_mai_n417_));
  NA2        m0395(.A(mai_mai_n415_), .B(mai_mai_n417_), .Y(mai_mai_n418_));
  NA2        m0396(.A(mai_mai_n418_), .B(mai_mai_n408_), .Y(mai_mai_n419_));
  NO3        m0397(.A(i_1_), .B(i_12_), .C(mai_mai_n87_), .Y(mai_mai_n420_));
  NO2        m0398(.A(i_0_), .B(i_11_), .Y(mai_mai_n421_));
  INV        m0399(.A(i_5_), .Y(mai_mai_n422_));
  AN2        m0400(.A(i_1_), .B(i_6_), .Y(mai_mai_n423_));
  NOi21      m0401(.An(i_2_), .B(i_12_), .Y(mai_mai_n424_));
  NA2        m0402(.A(mai_mai_n424_), .B(mai_mai_n423_), .Y(mai_mai_n425_));
  NO2        m0403(.A(mai_mai_n425_), .B(mai_mai_n422_), .Y(mai_mai_n426_));
  NA2        m0404(.A(mai_mai_n144_), .B(i_9_), .Y(mai_mai_n427_));
  NO2        m0405(.A(mai_mai_n427_), .B(i_4_), .Y(mai_mai_n428_));
  NA2        m0406(.A(mai_mai_n426_), .B(mai_mai_n428_), .Y(mai_mai_n429_));
  NAi21      m0407(.An(i_9_), .B(i_4_), .Y(mai_mai_n430_));
  OR2        m0408(.A(i_13_), .B(i_10_), .Y(mai_mai_n431_));
  NO3        m0409(.A(mai_mai_n431_), .B(mai_mai_n119_), .C(mai_mai_n430_), .Y(mai_mai_n432_));
  NO2        m0410(.A(mai_mai_n175_), .B(mai_mai_n125_), .Y(mai_mai_n433_));
  OR2        m0411(.A(mai_mai_n220_), .B(mai_mai_n219_), .Y(mai_mai_n434_));
  NO2        m0412(.A(mai_mai_n103_), .B(mai_mai_n25_), .Y(mai_mai_n435_));
  NA2        m0413(.A(mai_mai_n287_), .B(mai_mai_n435_), .Y(mai_mai_n436_));
  NA2        m0414(.A(mai_mai_n280_), .B(mai_mai_n214_), .Y(mai_mai_n437_));
  OAI220     m0415(.A0(mai_mai_n437_), .A1(mai_mai_n434_), .B0(mai_mai_n436_), .B1(mai_mai_n353_), .Y(mai_mai_n438_));
  INV        m0416(.A(mai_mai_n438_), .Y(mai_mai_n439_));
  AOI210     m0417(.A0(mai_mai_n439_), .A1(mai_mai_n429_), .B0(mai_mai_n26_), .Y(mai_mai_n440_));
  NA2        m0418(.A(mai_mai_n328_), .B(mai_mai_n327_), .Y(mai_mai_n441_));
  AOI220     m0419(.A0(mai_mai_n301_), .A1(mai_mai_n291_), .B0(mai_mai_n295_), .B1(mai_mai_n319_), .Y(mai_mai_n442_));
  NO2        m0420(.A(mai_mai_n442_), .B(mai_mai_n172_), .Y(mai_mai_n443_));
  NO2        m0421(.A(mai_mai_n186_), .B(mai_mai_n87_), .Y(mai_mai_n444_));
  AOI220     m0422(.A0(mai_mai_n444_), .A1(mai_mai_n300_), .B0(mai_mai_n282_), .B1(mai_mai_n214_), .Y(mai_mai_n445_));
  NO2        m0423(.A(mai_mai_n445_), .B(mai_mai_n289_), .Y(mai_mai_n446_));
  NO3        m0424(.A(mai_mai_n446_), .B(mai_mai_n443_), .C(mai_mai_n441_), .Y(mai_mai_n447_));
  NA2        m0425(.A(mai_mai_n200_), .B(mai_mai_n98_), .Y(mai_mai_n448_));
  NA3        m0426(.A(mai_mai_n331_), .B(mai_mai_n165_), .C(mai_mai_n87_), .Y(mai_mai_n449_));
  AOI210     m0427(.A0(mai_mai_n449_), .A1(mai_mai_n448_), .B0(mai_mai_n329_), .Y(mai_mai_n450_));
  NA2        m0428(.A(mai_mai_n197_), .B(i_10_), .Y(mai_mai_n451_));
  NA3        m0429(.A(mai_mai_n260_), .B(mai_mai_n65_), .C(i_2_), .Y(mai_mai_n452_));
  NA2        m0430(.A(mai_mai_n301_), .B(mai_mai_n236_), .Y(mai_mai_n453_));
  OAI220     m0431(.A0(mai_mai_n453_), .A1(mai_mai_n186_), .B0(mai_mai_n452_), .B1(mai_mai_n451_), .Y(mai_mai_n454_));
  NO2        m0432(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n455_));
  NA3        m0433(.A(mai_mai_n344_), .B(mai_mai_n343_), .C(mai_mai_n455_), .Y(mai_mai_n456_));
  NA2        m0434(.A(mai_mai_n321_), .B(mai_mai_n326_), .Y(mai_mai_n457_));
  OAI210     m0435(.A0(mai_mai_n457_), .A1(mai_mai_n193_), .B0(mai_mai_n456_), .Y(mai_mai_n458_));
  NO3        m0436(.A(mai_mai_n458_), .B(mai_mai_n454_), .C(mai_mai_n450_), .Y(mai_mai_n459_));
  AOI210     m0437(.A0(mai_mai_n459_), .A1(mai_mai_n447_), .B0(mai_mai_n276_), .Y(mai_mai_n460_));
  NO4        m0438(.A(mai_mai_n460_), .B(mai_mai_n440_), .C(mai_mai_n419_), .D(mai_mai_n396_), .Y(mai_mai_n461_));
  NO2        m0439(.A(mai_mai_n64_), .B(i_4_), .Y(mai_mai_n462_));
  NO2        m0440(.A(mai_mai_n74_), .B(i_13_), .Y(mai_mai_n463_));
  NO2        m0441(.A(i_10_), .B(i_9_), .Y(mai_mai_n464_));
  NAi21      m0442(.An(i_12_), .B(i_8_), .Y(mai_mai_n465_));
  NO2        m0443(.A(mai_mai_n465_), .B(i_3_), .Y(mai_mai_n466_));
  NA2        m0444(.A(mai_mai_n314_), .B(i_0_), .Y(mai_mai_n467_));
  NO3        m0445(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n468_));
  NA2        m0446(.A(mai_mai_n272_), .B(mai_mai_n99_), .Y(mai_mai_n469_));
  NA2        m0447(.A(mai_mai_n469_), .B(mai_mai_n468_), .Y(mai_mai_n470_));
  NA2        m0448(.A(i_8_), .B(i_9_), .Y(mai_mai_n471_));
  AOI210     m0449(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n472_));
  OR2        m0450(.A(mai_mai_n472_), .B(mai_mai_n471_), .Y(mai_mai_n473_));
  NA2        m0451(.A(mai_mai_n287_), .B(mai_mai_n209_), .Y(mai_mai_n474_));
  NO2        m0452(.A(mai_mai_n474_), .B(mai_mai_n473_), .Y(mai_mai_n475_));
  NA2        m0453(.A(mai_mai_n253_), .B(mai_mai_n313_), .Y(mai_mai_n476_));
  NO3        m0454(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n477_));
  AOI210     m0455(.A0(mai_mai_n259_), .A1(mai_mai_n192_), .B0(mai_mai_n477_), .Y(mai_mai_n478_));
  NA3        m0456(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n479_));
  NA4        m0457(.A(mai_mai_n147_), .B(mai_mai_n117_), .C(mai_mai_n81_), .D(mai_mai_n23_), .Y(mai_mai_n480_));
  OAI220     m0458(.A0(mai_mai_n480_), .A1(mai_mai_n479_), .B0(mai_mai_n478_), .B1(mai_mai_n476_), .Y(mai_mai_n481_));
  NO2        m0459(.A(mai_mai_n481_), .B(mai_mai_n475_), .Y(mai_mai_n482_));
  NA2        m0460(.A(mai_mai_n300_), .B(mai_mai_n110_), .Y(mai_mai_n483_));
  OR2        m0461(.A(mai_mai_n483_), .B(mai_mai_n211_), .Y(mai_mai_n484_));
  OA220      m0462(.A0(mai_mai_n302_), .A1(mai_mai_n164_), .B0(mai_mai_n484_), .B1(mai_mai_n233_), .Y(mai_mai_n485_));
  NA2        m0463(.A(mai_mai_n98_), .B(i_13_), .Y(mai_mai_n486_));
  NO2        m0464(.A(i_2_), .B(i_13_), .Y(mai_mai_n487_));
  NO3        m0465(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n488_));
  NO2        m0466(.A(i_6_), .B(i_7_), .Y(mai_mai_n489_));
  NA2        m0467(.A(mai_mai_n489_), .B(mai_mai_n488_), .Y(mai_mai_n490_));
  NO2        m0468(.A(i_11_), .B(i_1_), .Y(mai_mai_n491_));
  NO2        m0469(.A(mai_mai_n74_), .B(i_3_), .Y(mai_mai_n492_));
  OR2        m0470(.A(i_11_), .B(i_8_), .Y(mai_mai_n493_));
  NOi21      m0471(.An(i_2_), .B(i_7_), .Y(mai_mai_n494_));
  NAi31      m0472(.An(mai_mai_n493_), .B(mai_mai_n494_), .C(mai_mai_n492_), .Y(mai_mai_n495_));
  NO2        m0473(.A(mai_mai_n431_), .B(i_6_), .Y(mai_mai_n496_));
  NA3        m0474(.A(mai_mai_n496_), .B(mai_mai_n462_), .C(mai_mai_n76_), .Y(mai_mai_n497_));
  NO2        m0475(.A(mai_mai_n497_), .B(mai_mai_n495_), .Y(mai_mai_n498_));
  NO2        m0476(.A(i_3_), .B(mai_mai_n197_), .Y(mai_mai_n499_));
  NO2        m0477(.A(i_6_), .B(i_10_), .Y(mai_mai_n500_));
  NA4        m0478(.A(mai_mai_n500_), .B(mai_mai_n318_), .C(mai_mai_n499_), .D(mai_mai_n238_), .Y(mai_mai_n501_));
  NO2        m0479(.A(mai_mai_n501_), .B(mai_mai_n157_), .Y(mai_mai_n502_));
  NA3        m0480(.A(mai_mai_n247_), .B(mai_mai_n174_), .C(mai_mai_n134_), .Y(mai_mai_n503_));
  NA2        m0481(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n504_));
  NO2        m0482(.A(mai_mai_n159_), .B(i_3_), .Y(mai_mai_n505_));
  NAi31      m0483(.An(mai_mai_n504_), .B(mai_mai_n505_), .C(mai_mai_n228_), .Y(mai_mai_n506_));
  NA3        m0484(.A(mai_mai_n409_), .B(mai_mai_n182_), .C(mai_mai_n151_), .Y(mai_mai_n507_));
  NA3        m0485(.A(mai_mai_n507_), .B(mai_mai_n506_), .C(mai_mai_n503_), .Y(mai_mai_n508_));
  NO3        m0486(.A(mai_mai_n508_), .B(mai_mai_n502_), .C(mai_mai_n498_), .Y(mai_mai_n509_));
  NA2        m0487(.A(mai_mai_n468_), .B(mai_mai_n398_), .Y(mai_mai_n510_));
  NA2        m0488(.A(mai_mai_n477_), .B(mai_mai_n404_), .Y(mai_mai_n511_));
  NO2        m0489(.A(mai_mai_n511_), .B(mai_mai_n226_), .Y(mai_mai_n512_));
  NAi21      m0490(.An(mai_mai_n220_), .B(mai_mai_n412_), .Y(mai_mai_n513_));
  NO2        m0491(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n514_));
  NO2        m0492(.A(i_0_), .B(mai_mai_n87_), .Y(mai_mai_n515_));
  NA3        m0493(.A(mai_mai_n515_), .B(mai_mai_n514_), .C(mai_mai_n144_), .Y(mai_mai_n516_));
  OR3        m0494(.A(mai_mai_n308_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n517_));
  NO2        m0495(.A(mai_mai_n517_), .B(mai_mai_n516_), .Y(mai_mai_n518_));
  NA2        m0496(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n519_));
  NA2        m0497(.A(mai_mai_n318_), .B(mai_mai_n240_), .Y(mai_mai_n520_));
  OAI220     m0498(.A0(mai_mai_n520_), .A1(mai_mai_n452_), .B0(mai_mai_n519_), .B1(mai_mai_n486_), .Y(mai_mai_n521_));
  NA4        m0499(.A(mai_mai_n311_), .B(mai_mai_n225_), .C(mai_mai_n74_), .D(mai_mai_n238_), .Y(mai_mai_n522_));
  NO2        m0500(.A(mai_mai_n522_), .B(mai_mai_n490_), .Y(mai_mai_n523_));
  NO4        m0501(.A(mai_mai_n523_), .B(mai_mai_n521_), .C(mai_mai_n518_), .D(mai_mai_n512_), .Y(mai_mai_n524_));
  NA4        m0502(.A(mai_mai_n524_), .B(mai_mai_n509_), .C(mai_mai_n485_), .D(mai_mai_n482_), .Y(mai_mai_n525_));
  NA3        m0503(.A(mai_mai_n311_), .B(mai_mai_n179_), .C(mai_mai_n177_), .Y(mai_mai_n526_));
  OAI210     m0504(.A0(mai_mai_n306_), .A1(mai_mai_n184_), .B0(mai_mai_n526_), .Y(mai_mai_n527_));
  AN2        m0505(.A(mai_mai_n291_), .B(mai_mai_n235_), .Y(mai_mai_n528_));
  NA2        m0506(.A(mai_mai_n528_), .B(mai_mai_n527_), .Y(mai_mai_n529_));
  NA2        m0507(.A(mai_mai_n318_), .B(mai_mai_n166_), .Y(mai_mai_n530_));
  OAI210     m0508(.A0(mai_mai_n530_), .A1(mai_mai_n233_), .B0(mai_mai_n312_), .Y(mai_mai_n531_));
  NA2        m0509(.A(mai_mai_n531_), .B(mai_mai_n330_), .Y(mai_mai_n532_));
  NA4        m0510(.A(mai_mai_n463_), .B(mai_mai_n462_), .C(mai_mai_n207_), .D(i_2_), .Y(mai_mai_n533_));
  INV        m0511(.A(mai_mai_n533_), .Y(mai_mai_n534_));
  NA2        m0512(.A(mai_mai_n398_), .B(mai_mai_n227_), .Y(mai_mai_n535_));
  NA2        m0513(.A(mai_mai_n368_), .B(mai_mai_n74_), .Y(mai_mai_n536_));
  NA2        m0514(.A(mai_mai_n385_), .B(mai_mai_n377_), .Y(mai_mai_n537_));
  AO210      m0515(.A0(mai_mai_n536_), .A1(mai_mai_n535_), .B0(mai_mai_n537_), .Y(mai_mai_n538_));
  NO2        m0516(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n539_));
  NAi41      m0517(.An(mai_mai_n536_), .B(mai_mai_n500_), .C(mai_mai_n539_), .D(mai_mai_n47_), .Y(mai_mai_n540_));
  AOI210     m0518(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n432_), .Y(mai_mai_n541_));
  NA3        m0519(.A(mai_mai_n541_), .B(mai_mai_n540_), .C(mai_mai_n538_), .Y(mai_mai_n542_));
  AOI210     m0520(.A0(mai_mai_n534_), .A1(mai_mai_n208_), .B0(mai_mai_n542_), .Y(mai_mai_n543_));
  INV        m0521(.A(mai_mai_n136_), .Y(mai_mai_n544_));
  AOI210     m0522(.A0(mai_mai_n198_), .A1(i_9_), .B0(mai_mai_n271_), .Y(mai_mai_n545_));
  NO2        m0523(.A(mai_mai_n545_), .B(mai_mai_n203_), .Y(mai_mai_n546_));
  OR2        m0524(.A(mai_mai_n186_), .B(i_4_), .Y(mai_mai_n547_));
  NO2        m0525(.A(mai_mai_n547_), .B(mai_mai_n87_), .Y(mai_mai_n548_));
  AOI220     m0526(.A0(mai_mai_n548_), .A1(mai_mai_n546_), .B0(mai_mai_n544_), .B1(mai_mai_n433_), .Y(mai_mai_n549_));
  NA4        m0527(.A(mai_mai_n549_), .B(mai_mai_n543_), .C(mai_mai_n532_), .D(mai_mai_n529_), .Y(mai_mai_n550_));
  NA2        m0528(.A(mai_mai_n403_), .B(mai_mai_n300_), .Y(mai_mai_n551_));
  OAI210     m0529(.A0(mai_mai_n399_), .A1(mai_mai_n171_), .B0(mai_mai_n551_), .Y(mai_mai_n552_));
  NO2        m0530(.A(i_12_), .B(mai_mai_n197_), .Y(mai_mai_n553_));
  NA2        m0531(.A(mai_mai_n553_), .B(mai_mai_n227_), .Y(mai_mai_n554_));
  NA3        m0532(.A(mai_mai_n500_), .B(mai_mai_n177_), .C(mai_mai_n27_), .Y(mai_mai_n555_));
  NO2        m0533(.A(mai_mai_n555_), .B(mai_mai_n554_), .Y(mai_mai_n556_));
  NOi31      m0534(.An(mai_mai_n321_), .B(mai_mai_n431_), .C(mai_mai_n38_), .Y(mai_mai_n557_));
  OAI210     m0535(.A0(mai_mai_n557_), .A1(mai_mai_n556_), .B0(mai_mai_n552_), .Y(mai_mai_n558_));
  NO2        m0536(.A(i_8_), .B(i_7_), .Y(mai_mai_n559_));
  OAI210     m0537(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n560_));
  NA2        m0538(.A(mai_mai_n560_), .B(mai_mai_n225_), .Y(mai_mai_n561_));
  AOI220     m0539(.A0(mai_mai_n331_), .A1(mai_mai_n40_), .B0(mai_mai_n236_), .B1(mai_mai_n210_), .Y(mai_mai_n562_));
  OAI220     m0540(.A0(mai_mai_n562_), .A1(mai_mai_n547_), .B0(mai_mai_n561_), .B1(mai_mai_n244_), .Y(mai_mai_n563_));
  NA2        m0541(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n564_));
  NO2        m0542(.A(mai_mai_n564_), .B(i_6_), .Y(mai_mai_n565_));
  NA3        m0543(.A(mai_mai_n565_), .B(mai_mai_n563_), .C(mai_mai_n559_), .Y(mai_mai_n566_));
  NOi31      m0544(.An(mai_mai_n295_), .B(mai_mai_n306_), .C(mai_mai_n184_), .Y(mai_mai_n567_));
  NO2        m0545(.A(mai_mai_n159_), .B(i_5_), .Y(mai_mai_n568_));
  NA2        m0546(.A(mai_mai_n567_), .B(mai_mai_n477_), .Y(mai_mai_n569_));
  NA3        m0547(.A(mai_mai_n569_), .B(mai_mai_n566_), .C(mai_mai_n558_), .Y(mai_mai_n570_));
  NA3        m0548(.A(mai_mai_n221_), .B(mai_mai_n72_), .C(mai_mai_n45_), .Y(mai_mai_n571_));
  NA2        m0549(.A(mai_mai_n287_), .B(mai_mai_n85_), .Y(mai_mai_n572_));
  AOI210     m0550(.A0(mai_mai_n571_), .A1(mai_mai_n358_), .B0(mai_mai_n572_), .Y(mai_mai_n573_));
  NA2        m0551(.A(mai_mai_n301_), .B(mai_mai_n291_), .Y(mai_mai_n574_));
  NO2        m0552(.A(mai_mai_n574_), .B(mai_mai_n176_), .Y(mai_mai_n575_));
  NA2        m0553(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n576_));
  NA2        m0554(.A(mai_mai_n464_), .B(mai_mai_n223_), .Y(mai_mai_n577_));
  NO2        m0555(.A(mai_mai_n576_), .B(mai_mai_n577_), .Y(mai_mai_n578_));
  AOI210     m0556(.A0(mai_mai_n378_), .A1(mai_mai_n47_), .B0(mai_mai_n382_), .Y(mai_mai_n579_));
  NA2        m0557(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n580_));
  NA3        m0558(.A(mai_mai_n553_), .B(mai_mai_n278_), .C(mai_mai_n580_), .Y(mai_mai_n581_));
  NO2        m0559(.A(mai_mai_n579_), .B(mai_mai_n581_), .Y(mai_mai_n582_));
  NO4        m0560(.A(mai_mai_n582_), .B(mai_mai_n578_), .C(mai_mai_n575_), .D(mai_mai_n573_), .Y(mai_mai_n583_));
  NO4        m0561(.A(mai_mai_n254_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n584_));
  NO3        m0562(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n585_));
  NO2        m0563(.A(mai_mai_n234_), .B(mai_mai_n36_), .Y(mai_mai_n586_));
  AN2        m0564(.A(mai_mai_n586_), .B(mai_mai_n585_), .Y(mai_mai_n587_));
  OA210      m0565(.A0(mai_mai_n587_), .A1(mai_mai_n584_), .B0(mai_mai_n368_), .Y(mai_mai_n588_));
  NO2        m0566(.A(mai_mai_n431_), .B(i_1_), .Y(mai_mai_n589_));
  NOi31      m0567(.An(mai_mai_n589_), .B(mai_mai_n469_), .C(mai_mai_n74_), .Y(mai_mai_n590_));
  AN4        m0568(.A(mai_mai_n590_), .B(mai_mai_n428_), .C(mai_mai_n514_), .D(i_2_), .Y(mai_mai_n591_));
  NO2        m0569(.A(mai_mai_n442_), .B(mai_mai_n180_), .Y(mai_mai_n592_));
  NO3        m0570(.A(mai_mai_n592_), .B(mai_mai_n591_), .C(mai_mai_n588_), .Y(mai_mai_n593_));
  NOi21      m0571(.An(i_10_), .B(i_6_), .Y(mai_mai_n594_));
  NO2        m0572(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n595_));
  NO2        m0573(.A(mai_mai_n116_), .B(mai_mai_n23_), .Y(mai_mai_n596_));
  NA2        m0574(.A(mai_mai_n321_), .B(mai_mai_n166_), .Y(mai_mai_n597_));
  AOI220     m0575(.A0(mai_mai_n597_), .A1(mai_mai_n453_), .B0(mai_mai_n187_), .B1(mai_mai_n185_), .Y(mai_mai_n598_));
  NOi31      m0576(.An(mai_mai_n148_), .B(i_10_), .C(mai_mai_n339_), .Y(mai_mai_n599_));
  NO2        m0577(.A(mai_mai_n599_), .B(mai_mai_n598_), .Y(mai_mai_n600_));
  NO2        m0578(.A(i_12_), .B(mai_mai_n87_), .Y(mai_mai_n601_));
  NA2        m0579(.A(mai_mai_n177_), .B(i_0_), .Y(mai_mai_n602_));
  NO3        m0580(.A(mai_mai_n602_), .B(mai_mai_n350_), .C(mai_mai_n306_), .Y(mai_mai_n603_));
  OR2        m0581(.A(i_2_), .B(i_5_), .Y(mai_mai_n604_));
  OR2        m0582(.A(mai_mai_n604_), .B(mai_mai_n423_), .Y(mai_mai_n605_));
  AOI210     m0583(.A0(mai_mai_n387_), .A1(mai_mai_n246_), .B0(mai_mai_n202_), .Y(mai_mai_n606_));
  AOI210     m0584(.A0(mai_mai_n606_), .A1(mai_mai_n605_), .B0(mai_mai_n513_), .Y(mai_mai_n607_));
  NO2        m0585(.A(mai_mai_n607_), .B(mai_mai_n603_), .Y(mai_mai_n608_));
  NA4        m0586(.A(mai_mai_n608_), .B(mai_mai_n600_), .C(mai_mai_n593_), .D(mai_mai_n583_), .Y(mai_mai_n609_));
  NO4        m0587(.A(mai_mai_n609_), .B(mai_mai_n570_), .C(mai_mai_n550_), .D(mai_mai_n525_), .Y(mai_mai_n610_));
  NA4        m0588(.A(mai_mai_n610_), .B(mai_mai_n461_), .C(mai_mai_n367_), .D(mai_mai_n317_), .Y(mai7));
  NO2        m0589(.A(mai_mai_n94_), .B(mai_mai_n55_), .Y(mai_mai_n612_));
  NA2        m0590(.A(mai_mai_n500_), .B(mai_mai_n85_), .Y(mai_mai_n613_));
  NA2        m0591(.A(i_11_), .B(mai_mai_n197_), .Y(mai_mai_n614_));
  NA2        m0592(.A(mai_mai_n146_), .B(mai_mai_n614_), .Y(mai_mai_n615_));
  NO2        m0593(.A(mai_mai_n615_), .B(mai_mai_n613_), .Y(mai_mai_n616_));
  NA3        m0594(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n617_));
  NO2        m0595(.A(mai_mai_n238_), .B(i_4_), .Y(mai_mai_n618_));
  NA2        m0596(.A(mai_mai_n618_), .B(i_8_), .Y(mai_mai_n619_));
  NO2        m0597(.A(mai_mai_n107_), .B(mai_mai_n617_), .Y(mai_mai_n620_));
  NA2        m0598(.A(i_2_), .B(mai_mai_n87_), .Y(mai_mai_n621_));
  OAI210     m0599(.A0(mai_mai_n88_), .A1(mai_mai_n207_), .B0(mai_mai_n208_), .Y(mai_mai_n622_));
  NO2        m0600(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n623_));
  NA2        m0601(.A(i_4_), .B(i_8_), .Y(mai_mai_n624_));
  AOI210     m0602(.A0(mai_mai_n624_), .A1(mai_mai_n311_), .B0(mai_mai_n623_), .Y(mai_mai_n625_));
  OAI220     m0603(.A0(mai_mai_n625_), .A1(mai_mai_n621_), .B0(mai_mai_n622_), .B1(i_13_), .Y(mai_mai_n626_));
  NO4        m0604(.A(mai_mai_n626_), .B(mai_mai_n620_), .C(mai_mai_n616_), .D(mai_mai_n612_), .Y(mai_mai_n627_));
  AOI210     m0605(.A0(mai_mai_n130_), .A1(mai_mai_n63_), .B0(i_10_), .Y(mai_mai_n628_));
  AOI210     m0606(.A0(mai_mai_n628_), .A1(mai_mai_n238_), .B0(mai_mai_n163_), .Y(mai_mai_n629_));
  OR2        m0607(.A(i_6_), .B(i_10_), .Y(mai_mai_n630_));
  NO2        m0608(.A(mai_mai_n630_), .B(mai_mai_n23_), .Y(mai_mai_n631_));
  OR3        m0609(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n632_));
  NO3        m0610(.A(mai_mai_n632_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n633_));
  INV        m0611(.A(mai_mai_n204_), .Y(mai_mai_n634_));
  OR2        m0612(.A(mai_mai_n629_), .B(mai_mai_n273_), .Y(mai_mai_n635_));
  AOI210     m0613(.A0(mai_mai_n635_), .A1(mai_mai_n627_), .B0(mai_mai_n64_), .Y(mai_mai_n636_));
  NOi21      m0614(.An(i_11_), .B(i_7_), .Y(mai_mai_n637_));
  AO210      m0615(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n638_));
  NO2        m0616(.A(mai_mai_n638_), .B(mai_mai_n637_), .Y(mai_mai_n639_));
  NA2        m0617(.A(mai_mai_n639_), .B(mai_mai_n210_), .Y(mai_mai_n640_));
  NA3        m0618(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n641_));
  NO2        m0619(.A(mai_mai_n640_), .B(mai_mai_n64_), .Y(mai_mai_n642_));
  OR2        m0620(.A(mai_mai_n393_), .B(mai_mai_n41_), .Y(mai_mai_n643_));
  NO3        m0621(.A(mai_mai_n262_), .B(mai_mai_n212_), .C(mai_mai_n614_), .Y(mai_mai_n644_));
  OAI210     m0622(.A0(mai_mai_n644_), .A1(mai_mai_n228_), .B0(mai_mai_n64_), .Y(mai_mai_n645_));
  NA2        m0623(.A(mai_mai_n424_), .B(mai_mai_n31_), .Y(mai_mai_n646_));
  OR2        m0624(.A(mai_mai_n212_), .B(mai_mai_n110_), .Y(mai_mai_n647_));
  NA2        m0625(.A(mai_mai_n647_), .B(mai_mai_n646_), .Y(mai_mai_n648_));
  NO2        m0626(.A(mai_mai_n64_), .B(i_9_), .Y(mai_mai_n649_));
  NO2        m0627(.A(mai_mai_n649_), .B(i_4_), .Y(mai_mai_n650_));
  NA2        m0628(.A(mai_mai_n650_), .B(mai_mai_n648_), .Y(mai_mai_n651_));
  NO2        m0629(.A(i_1_), .B(i_12_), .Y(mai_mai_n652_));
  NA3        m0630(.A(mai_mai_n651_), .B(mai_mai_n645_), .C(mai_mai_n643_), .Y(mai_mai_n653_));
  OAI210     m0631(.A0(mai_mai_n653_), .A1(mai_mai_n642_), .B0(i_6_), .Y(mai_mai_n654_));
  NO2        m0632(.A(mai_mai_n641_), .B(mai_mai_n110_), .Y(mai_mai_n655_));
  NA2        m0633(.A(mai_mai_n655_), .B(mai_mai_n601_), .Y(mai_mai_n656_));
  NO2        m0634(.A(i_6_), .B(i_11_), .Y(mai_mai_n657_));
  NA2        m0635(.A(mai_mai_n656_), .B(mai_mai_n470_), .Y(mai_mai_n658_));
  NO4        m0636(.A(mai_mai_n219_), .B(mai_mai_n130_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n659_));
  NA2        m0637(.A(mai_mai_n659_), .B(mai_mai_n649_), .Y(mai_mai_n660_));
  NA2        m0638(.A(mai_mai_n238_), .B(i_6_), .Y(mai_mai_n661_));
  NO3        m0639(.A(mai_mai_n630_), .B(mai_mai_n234_), .C(mai_mai_n23_), .Y(mai_mai_n662_));
  AOI210     m0640(.A0(i_1_), .A1(mai_mai_n263_), .B0(mai_mai_n662_), .Y(mai_mai_n663_));
  OAI210     m0641(.A0(mai_mai_n663_), .A1(mai_mai_n45_), .B0(mai_mai_n660_), .Y(mai_mai_n664_));
  NA3        m0642(.A(mai_mai_n559_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n665_));
  NA2        m0643(.A(mai_mai_n140_), .B(i_9_), .Y(mai_mai_n666_));
  NA3        m0644(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n667_));
  NO2        m0645(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n668_));
  NA3        m0646(.A(mai_mai_n668_), .B(mai_mai_n272_), .C(mai_mai_n45_), .Y(mai_mai_n669_));
  OAI220     m0647(.A0(mai_mai_n669_), .A1(mai_mai_n667_), .B0(mai_mai_n666_), .B1(mai_mai_n1073_), .Y(mai_mai_n670_));
  NA3        m0648(.A(mai_mai_n649_), .B(mai_mai_n324_), .C(i_6_), .Y(mai_mai_n671_));
  NO2        m0649(.A(mai_mai_n671_), .B(mai_mai_n23_), .Y(mai_mai_n672_));
  AOI210     m0650(.A0(mai_mai_n491_), .A1(mai_mai_n435_), .B0(mai_mai_n243_), .Y(mai_mai_n673_));
  NO2        m0651(.A(mai_mai_n673_), .B(mai_mai_n621_), .Y(mai_mai_n674_));
  NAi21      m0652(.An(mai_mai_n665_), .B(mai_mai_n93_), .Y(mai_mai_n675_));
  NA2        m0653(.A(mai_mai_n668_), .B(mai_mai_n272_), .Y(mai_mai_n676_));
  NO2        m0654(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n677_));
  NA2        m0655(.A(mai_mai_n677_), .B(mai_mai_n24_), .Y(mai_mai_n678_));
  OAI210     m0656(.A0(mai_mai_n678_), .A1(mai_mai_n676_), .B0(mai_mai_n675_), .Y(mai_mai_n679_));
  OR4        m0657(.A(mai_mai_n679_), .B(mai_mai_n674_), .C(mai_mai_n672_), .D(mai_mai_n670_), .Y(mai_mai_n680_));
  NO3        m0658(.A(mai_mai_n680_), .B(mai_mai_n664_), .C(mai_mai_n658_), .Y(mai_mai_n681_));
  NO2        m0659(.A(mai_mai_n238_), .B(mai_mai_n103_), .Y(mai_mai_n682_));
  NO2        m0660(.A(mai_mai_n682_), .B(mai_mai_n637_), .Y(mai_mai_n683_));
  NA2        m0661(.A(mai_mai_n683_), .B(i_1_), .Y(mai_mai_n684_));
  NO2        m0662(.A(mai_mai_n684_), .B(mai_mai_n632_), .Y(mai_mai_n685_));
  NO2        m0663(.A(mai_mai_n430_), .B(mai_mai_n87_), .Y(mai_mai_n686_));
  NA2        m0664(.A(mai_mai_n685_), .B(mai_mai_n47_), .Y(mai_mai_n687_));
  NA2        m0665(.A(i_3_), .B(mai_mai_n197_), .Y(mai_mai_n688_));
  NO2        m0666(.A(mai_mai_n688_), .B(mai_mai_n116_), .Y(mai_mai_n689_));
  AN2        m0667(.A(mai_mai_n689_), .B(mai_mai_n565_), .Y(mai_mai_n690_));
  NO2        m0668(.A(mai_mai_n234_), .B(mai_mai_n45_), .Y(mai_mai_n691_));
  NO3        m0669(.A(mai_mai_n691_), .B(mai_mai_n314_), .C(mai_mai_n239_), .Y(mai_mai_n692_));
  NO2        m0670(.A(mai_mai_n119_), .B(mai_mai_n37_), .Y(mai_mai_n693_));
  NO2        m0671(.A(mai_mai_n693_), .B(i_6_), .Y(mai_mai_n694_));
  NO2        m0672(.A(mai_mai_n87_), .B(i_9_), .Y(mai_mai_n695_));
  NO2        m0673(.A(mai_mai_n695_), .B(mai_mai_n64_), .Y(mai_mai_n696_));
  NO2        m0674(.A(mai_mai_n696_), .B(mai_mai_n652_), .Y(mai_mai_n697_));
  NO4        m0675(.A(mai_mai_n697_), .B(mai_mai_n694_), .C(mai_mai_n692_), .D(i_4_), .Y(mai_mai_n698_));
  NA2        m0676(.A(i_1_), .B(i_3_), .Y(mai_mai_n699_));
  NO2        m0677(.A(mai_mai_n471_), .B(mai_mai_n94_), .Y(mai_mai_n700_));
  AOI210     m0678(.A0(mai_mai_n691_), .A1(mai_mai_n594_), .B0(mai_mai_n700_), .Y(mai_mai_n701_));
  NO2        m0679(.A(mai_mai_n701_), .B(mai_mai_n699_), .Y(mai_mai_n702_));
  NO3        m0680(.A(mai_mai_n702_), .B(mai_mai_n698_), .C(mai_mai_n690_), .Y(mai_mai_n703_));
  NA4        m0681(.A(mai_mai_n703_), .B(mai_mai_n687_), .C(mai_mai_n681_), .D(mai_mai_n654_), .Y(mai_mai_n704_));
  NO3        m0682(.A(mai_mai_n493_), .B(i_3_), .C(i_7_), .Y(mai_mai_n705_));
  NOi21      m0683(.An(mai_mai_n705_), .B(i_10_), .Y(mai_mai_n706_));
  OA210      m0684(.A0(mai_mai_n706_), .A1(mai_mai_n247_), .B0(mai_mai_n87_), .Y(mai_mai_n707_));
  NA2        m0685(.A(mai_mai_n385_), .B(mai_mai_n384_), .Y(mai_mai_n708_));
  NA3        m0686(.A(mai_mai_n500_), .B(mai_mai_n539_), .C(mai_mai_n47_), .Y(mai_mai_n709_));
  NO3        m0687(.A(mai_mai_n494_), .B(mai_mai_n624_), .C(mai_mai_n87_), .Y(mai_mai_n710_));
  NA2        m0688(.A(mai_mai_n710_), .B(mai_mai_n25_), .Y(mai_mai_n711_));
  NA3        m0689(.A(mai_mai_n711_), .B(mai_mai_n709_), .C(mai_mai_n708_), .Y(mai_mai_n712_));
  OAI210     m0690(.A0(mai_mai_n712_), .A1(mai_mai_n707_), .B0(i_1_), .Y(mai_mai_n713_));
  AOI210     m0691(.A0(mai_mai_n272_), .A1(mai_mai_n99_), .B0(i_1_), .Y(mai_mai_n714_));
  NO2        m0692(.A(mai_mai_n383_), .B(i_2_), .Y(mai_mai_n715_));
  NA2        m0693(.A(mai_mai_n715_), .B(mai_mai_n714_), .Y(mai_mai_n716_));
  OAI210     m0694(.A0(mai_mai_n671_), .A1(mai_mai_n465_), .B0(mai_mai_n716_), .Y(mai_mai_n717_));
  INV        m0695(.A(mai_mai_n717_), .Y(mai_mai_n718_));
  AOI210     m0696(.A0(mai_mai_n718_), .A1(mai_mai_n713_), .B0(i_13_), .Y(mai_mai_n719_));
  OR2        m0697(.A(i_11_), .B(i_7_), .Y(mai_mai_n720_));
  AOI210     m0698(.A0(mai_mai_n667_), .A1(mai_mai_n55_), .B0(i_12_), .Y(mai_mai_n721_));
  NO2        m0699(.A(mai_mai_n494_), .B(mai_mai_n24_), .Y(mai_mai_n722_));
  AOI220     m0700(.A0(mai_mai_n722_), .A1(mai_mai_n686_), .B0(mai_mai_n247_), .B1(mai_mai_n133_), .Y(mai_mai_n723_));
  OAI220     m0701(.A0(mai_mai_n723_), .A1(mai_mai_n41_), .B0(mai_mai_n1072_), .B1(mai_mai_n94_), .Y(mai_mai_n724_));
  INV        m0702(.A(mai_mai_n724_), .Y(mai_mai_n725_));
  INV        m0703(.A(mai_mai_n116_), .Y(mai_mai_n726_));
  AOI220     m0704(.A0(mai_mai_n726_), .A1(mai_mai_n73_), .B0(mai_mai_n400_), .B1(mai_mai_n668_), .Y(mai_mai_n727_));
  NO2        m0705(.A(mai_mai_n727_), .B(mai_mai_n244_), .Y(mai_mai_n728_));
  AOI210     m0706(.A0(mai_mai_n465_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n729_));
  NOi31      m0707(.An(mai_mai_n729_), .B(mai_mai_n613_), .C(mai_mai_n45_), .Y(mai_mai_n730_));
  NA2        m0708(.A(mai_mai_n129_), .B(i_13_), .Y(mai_mai_n731_));
  NO2        m0709(.A(mai_mai_n667_), .B(mai_mai_n116_), .Y(mai_mai_n732_));
  INV        m0710(.A(mai_mai_n732_), .Y(mai_mai_n733_));
  OAI220     m0711(.A0(mai_mai_n733_), .A1(mai_mai_n72_), .B0(mai_mai_n731_), .B1(mai_mai_n714_), .Y(mai_mai_n734_));
  NA2        m0712(.A(mai_mai_n26_), .B(mai_mai_n197_), .Y(mai_mai_n735_));
  NA2        m0713(.A(mai_mai_n735_), .B(i_7_), .Y(mai_mai_n736_));
  NO3        m0714(.A(mai_mai_n494_), .B(mai_mai_n238_), .C(mai_mai_n87_), .Y(mai_mai_n737_));
  NA2        m0715(.A(mai_mai_n737_), .B(mai_mai_n736_), .Y(mai_mai_n738_));
  AOI220     m0716(.A0(mai_mai_n400_), .A1(mai_mai_n668_), .B0(mai_mai_n93_), .B1(mai_mai_n104_), .Y(mai_mai_n739_));
  OAI220     m0717(.A0(mai_mai_n739_), .A1(mai_mai_n619_), .B0(mai_mai_n738_), .B1(mai_mai_n634_), .Y(mai_mai_n740_));
  NO4        m0718(.A(mai_mai_n740_), .B(mai_mai_n734_), .C(mai_mai_n730_), .D(mai_mai_n728_), .Y(mai_mai_n741_));
  OR2        m0719(.A(i_11_), .B(i_6_), .Y(mai_mai_n742_));
  NA3        m0720(.A(mai_mai_n618_), .B(mai_mai_n735_), .C(i_7_), .Y(mai_mai_n743_));
  AOI210     m0721(.A0(mai_mai_n743_), .A1(mai_mai_n733_), .B0(mai_mai_n742_), .Y(mai_mai_n744_));
  NA3        m0722(.A(mai_mai_n424_), .B(mai_mai_n623_), .C(mai_mai_n99_), .Y(mai_mai_n745_));
  NA2        m0723(.A(mai_mai_n657_), .B(i_13_), .Y(mai_mai_n746_));
  NA2        m0724(.A(mai_mai_n104_), .B(mai_mai_n735_), .Y(mai_mai_n747_));
  NAi21      m0725(.An(i_11_), .B(i_12_), .Y(mai_mai_n748_));
  NOi41      m0726(.An(mai_mai_n112_), .B(mai_mai_n748_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n749_));
  NO3        m0727(.A(mai_mai_n494_), .B(mai_mai_n601_), .C(mai_mai_n624_), .Y(mai_mai_n750_));
  AOI220     m0728(.A0(mai_mai_n750_), .A1(mai_mai_n318_), .B0(mai_mai_n749_), .B1(mai_mai_n747_), .Y(mai_mai_n751_));
  NA3        m0729(.A(mai_mai_n751_), .B(mai_mai_n746_), .C(mai_mai_n745_), .Y(mai_mai_n752_));
  OAI210     m0730(.A0(mai_mai_n752_), .A1(mai_mai_n744_), .B0(mai_mai_n64_), .Y(mai_mai_n753_));
  NO2        m0731(.A(i_2_), .B(i_12_), .Y(mai_mai_n754_));
  NA2        m0732(.A(mai_mai_n382_), .B(mai_mai_n754_), .Y(mai_mai_n755_));
  NA2        m0733(.A(mai_mai_n384_), .B(mai_mai_n382_), .Y(mai_mai_n756_));
  NO2        m0734(.A(mai_mai_n130_), .B(i_2_), .Y(mai_mai_n757_));
  NA2        m0735(.A(mai_mai_n757_), .B(mai_mai_n652_), .Y(mai_mai_n758_));
  NA3        m0736(.A(mai_mai_n758_), .B(mai_mai_n756_), .C(mai_mai_n755_), .Y(mai_mai_n759_));
  NA3        m0737(.A(mai_mai_n759_), .B(mai_mai_n46_), .C(mai_mai_n227_), .Y(mai_mai_n760_));
  NA4        m0738(.A(mai_mai_n760_), .B(mai_mai_n753_), .C(mai_mai_n741_), .D(mai_mai_n725_), .Y(mai_mai_n761_));
  OR4        m0739(.A(mai_mai_n761_), .B(mai_mai_n719_), .C(mai_mai_n704_), .D(mai_mai_n636_), .Y(mai5));
  NA2        m0740(.A(mai_mai_n683_), .B(mai_mai_n275_), .Y(mai_mai_n763_));
  AN2        m0741(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n764_));
  NA3        m0742(.A(mai_mai_n764_), .B(mai_mai_n754_), .C(mai_mai_n110_), .Y(mai_mai_n765_));
  NO2        m0743(.A(mai_mai_n619_), .B(i_11_), .Y(mai_mai_n766_));
  OAI210     m0744(.A0(mai_mai_n623_), .A1(mai_mai_n88_), .B0(mai_mai_n766_), .Y(mai_mai_n767_));
  NA3        m0745(.A(mai_mai_n767_), .B(mai_mai_n765_), .C(mai_mai_n763_), .Y(mai_mai_n768_));
  NO3        m0746(.A(i_11_), .B(mai_mai_n238_), .C(i_13_), .Y(mai_mai_n769_));
  NO2        m0747(.A(mai_mai_n126_), .B(mai_mai_n23_), .Y(mai_mai_n770_));
  NA2        m0748(.A(i_12_), .B(i_8_), .Y(mai_mai_n771_));
  OAI210     m0749(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n771_), .Y(mai_mai_n772_));
  INV        m0750(.A(mai_mai_n464_), .Y(mai_mai_n773_));
  AOI220     m0751(.A0(mai_mai_n324_), .A1(mai_mai_n596_), .B0(mai_mai_n772_), .B1(mai_mai_n770_), .Y(mai_mai_n774_));
  INV        m0752(.A(mai_mai_n774_), .Y(mai_mai_n775_));
  NO2        m0753(.A(mai_mai_n775_), .B(mai_mai_n768_), .Y(mai_mai_n776_));
  INV        m0754(.A(mai_mai_n174_), .Y(mai_mai_n777_));
  INV        m0755(.A(mai_mai_n247_), .Y(mai_mai_n778_));
  OAI210     m0756(.A0(mai_mai_n715_), .A1(mai_mai_n466_), .B0(mai_mai_n112_), .Y(mai_mai_n779_));
  AOI210     m0757(.A0(mai_mai_n779_), .A1(mai_mai_n778_), .B0(mai_mai_n777_), .Y(mai_mai_n780_));
  NO2        m0758(.A(mai_mai_n471_), .B(mai_mai_n26_), .Y(mai_mai_n781_));
  NO2        m0759(.A(mai_mai_n781_), .B(mai_mai_n435_), .Y(mai_mai_n782_));
  NA2        m0760(.A(mai_mai_n782_), .B(i_2_), .Y(mai_mai_n783_));
  INV        m0761(.A(mai_mai_n783_), .Y(mai_mai_n784_));
  AOI210     m0762(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n431_), .Y(mai_mai_n785_));
  AOI210     m0763(.A0(mai_mai_n785_), .A1(mai_mai_n784_), .B0(mai_mai_n780_), .Y(mai_mai_n786_));
  NO2        m0764(.A(mai_mai_n194_), .B(mai_mai_n127_), .Y(mai_mai_n787_));
  OAI210     m0765(.A0(mai_mai_n787_), .A1(mai_mai_n770_), .B0(i_2_), .Y(mai_mai_n788_));
  INV        m0766(.A(mai_mai_n175_), .Y(mai_mai_n789_));
  NO3        m0767(.A(mai_mai_n638_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n790_));
  AOI210     m0768(.A0(mai_mai_n789_), .A1(mai_mai_n88_), .B0(mai_mai_n790_), .Y(mai_mai_n791_));
  AOI210     m0769(.A0(mai_mai_n791_), .A1(mai_mai_n788_), .B0(mai_mai_n197_), .Y(mai_mai_n792_));
  OA210      m0770(.A0(mai_mai_n639_), .A1(mai_mai_n128_), .B0(i_13_), .Y(mai_mai_n793_));
  NA2        m0771(.A(mai_mai_n204_), .B(mai_mai_n207_), .Y(mai_mai_n794_));
  NA2        m0772(.A(mai_mai_n153_), .B(mai_mai_n614_), .Y(mai_mai_n795_));
  AOI210     m0773(.A0(mai_mai_n795_), .A1(mai_mai_n794_), .B0(mai_mai_n387_), .Y(mai_mai_n796_));
  AOI210     m0774(.A0(mai_mai_n212_), .A1(mai_mai_n150_), .B0(mai_mai_n539_), .Y(mai_mai_n797_));
  OAI210     m0775(.A0(mai_mai_n797_), .A1(mai_mai_n228_), .B0(mai_mai_n435_), .Y(mai_mai_n798_));
  NO2        m0776(.A(mai_mai_n104_), .B(mai_mai_n45_), .Y(mai_mai_n799_));
  INV        m0777(.A(mai_mai_n307_), .Y(mai_mai_n800_));
  NA4        m0778(.A(mai_mai_n800_), .B(mai_mai_n311_), .C(mai_mai_n126_), .D(mai_mai_n43_), .Y(mai_mai_n801_));
  OAI210     m0779(.A0(mai_mai_n801_), .A1(mai_mai_n799_), .B0(mai_mai_n798_), .Y(mai_mai_n802_));
  NO4        m0780(.A(mai_mai_n802_), .B(mai_mai_n796_), .C(mai_mai_n793_), .D(mai_mai_n792_), .Y(mai_mai_n803_));
  NA2        m0781(.A(mai_mai_n596_), .B(mai_mai_n28_), .Y(mai_mai_n804_));
  NA2        m0782(.A(mai_mai_n769_), .B(mai_mai_n279_), .Y(mai_mai_n805_));
  NA2        m0783(.A(mai_mai_n805_), .B(mai_mai_n804_), .Y(mai_mai_n806_));
  NO2        m0784(.A(mai_mai_n63_), .B(i_12_), .Y(mai_mai_n807_));
  NO2        m0785(.A(mai_mai_n807_), .B(mai_mai_n128_), .Y(mai_mai_n808_));
  NO2        m0786(.A(mai_mai_n808_), .B(mai_mai_n614_), .Y(mai_mai_n809_));
  AOI220     m0787(.A0(mai_mai_n809_), .A1(mai_mai_n36_), .B0(mai_mai_n806_), .B1(mai_mai_n47_), .Y(mai_mai_n810_));
  NA4        m0788(.A(mai_mai_n810_), .B(mai_mai_n803_), .C(mai_mai_n786_), .D(mai_mai_n776_), .Y(mai6));
  NO3        m0789(.A(mai_mai_n258_), .B(mai_mai_n313_), .C(i_1_), .Y(mai_mai_n812_));
  NO2        m0790(.A(mai_mai_n189_), .B(mai_mai_n141_), .Y(mai_mai_n813_));
  OAI210     m0791(.A0(mai_mai_n813_), .A1(mai_mai_n812_), .B0(mai_mai_n757_), .Y(mai_mai_n814_));
  NA4        m0792(.A(mai_mai_n404_), .B(mai_mai_n499_), .C(mai_mai_n72_), .D(mai_mai_n103_), .Y(mai_mai_n815_));
  INV        m0793(.A(mai_mai_n815_), .Y(mai_mai_n816_));
  NO2        m0794(.A(mai_mai_n222_), .B(mai_mai_n504_), .Y(mai_mai_n817_));
  NO2        m0795(.A(i_11_), .B(i_9_), .Y(mai_mai_n818_));
  NO2        m0796(.A(mai_mai_n816_), .B(mai_mai_n336_), .Y(mai_mai_n819_));
  AO210      m0797(.A0(mai_mai_n819_), .A1(mai_mai_n814_), .B0(i_12_), .Y(mai_mai_n820_));
  NA2        m0798(.A(mai_mai_n388_), .B(mai_mai_n344_), .Y(mai_mai_n821_));
  NA2        m0799(.A(mai_mai_n601_), .B(mai_mai_n64_), .Y(mai_mai_n822_));
  NA2        m0800(.A(mai_mai_n706_), .B(mai_mai_n72_), .Y(mai_mai_n823_));
  NA3        m0801(.A(mai_mai_n823_), .B(mai_mai_n822_), .C(mai_mai_n821_), .Y(mai_mai_n824_));
  INV        m0802(.A(mai_mai_n201_), .Y(mai_mai_n825_));
  AOI220     m0803(.A0(mai_mai_n825_), .A1(mai_mai_n818_), .B0(mai_mai_n824_), .B1(mai_mai_n74_), .Y(mai_mai_n826_));
  INV        m0804(.A(mai_mai_n335_), .Y(mai_mai_n827_));
  NA2        m0805(.A(mai_mai_n76_), .B(mai_mai_n133_), .Y(mai_mai_n828_));
  INV        m0806(.A(mai_mai_n126_), .Y(mai_mai_n829_));
  NA2        m0807(.A(mai_mai_n829_), .B(mai_mai_n47_), .Y(mai_mai_n830_));
  AOI210     m0808(.A0(mai_mai_n830_), .A1(mai_mai_n828_), .B0(mai_mai_n827_), .Y(mai_mai_n831_));
  NO3        m0809(.A(mai_mai_n254_), .B(mai_mai_n134_), .C(i_9_), .Y(mai_mai_n832_));
  NA2        m0810(.A(mai_mai_n832_), .B(mai_mai_n807_), .Y(mai_mai_n833_));
  AOI210     m0811(.A0(mai_mai_n833_), .A1(mai_mai_n537_), .B0(mai_mai_n189_), .Y(mai_mai_n834_));
  NO2        m0812(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n835_));
  NA3        m0813(.A(mai_mai_n835_), .B(mai_mai_n489_), .C(mai_mai_n404_), .Y(mai_mai_n836_));
  NAi32      m0814(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n837_));
  NO2        m0815(.A(mai_mai_n742_), .B(mai_mai_n837_), .Y(mai_mai_n838_));
  OAI210     m0816(.A0(mai_mai_n705_), .A1(mai_mai_n586_), .B0(mai_mai_n585_), .Y(mai_mai_n839_));
  NAi31      m0817(.An(mai_mai_n838_), .B(mai_mai_n839_), .C(mai_mai_n836_), .Y(mai_mai_n840_));
  OR3        m0818(.A(mai_mai_n840_), .B(mai_mai_n834_), .C(mai_mai_n831_), .Y(mai_mai_n841_));
  NO2        m0819(.A(mai_mai_n720_), .B(i_2_), .Y(mai_mai_n842_));
  NA2        m0820(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n843_));
  NO2        m0821(.A(mai_mai_n843_), .B(mai_mai_n423_), .Y(mai_mai_n844_));
  NA2        m0822(.A(mai_mai_n844_), .B(mai_mai_n842_), .Y(mai_mai_n845_));
  AO220      m0823(.A0(mai_mai_n372_), .A1(mai_mai_n362_), .B0(mai_mai_n410_), .B1(mai_mai_n614_), .Y(mai_mai_n846_));
  NA3        m0824(.A(mai_mai_n846_), .B(mai_mai_n259_), .C(i_7_), .Y(mai_mai_n847_));
  NA3        m0825(.A(mai_mai_n639_), .B(mai_mai_n149_), .C(mai_mai_n70_), .Y(mai_mai_n848_));
  AO210      m0826(.A0(mai_mai_n511_), .A1(mai_mai_n773_), .B0(mai_mai_n36_), .Y(mai_mai_n849_));
  NA4        m0827(.A(mai_mai_n849_), .B(mai_mai_n848_), .C(mai_mai_n847_), .D(mai_mai_n845_), .Y(mai_mai_n850_));
  NO2        m0828(.A(i_6_), .B(i_11_), .Y(mai_mai_n851_));
  AOI220     m0829(.A0(mai_mai_n851_), .A1(mai_mai_n585_), .B0(mai_mai_n817_), .B1(mai_mai_n736_), .Y(mai_mai_n852_));
  NA3        m0830(.A(mai_mai_n387_), .B(mai_mai_n240_), .C(mai_mai_n149_), .Y(mai_mai_n853_));
  NA2        m0831(.A(mai_mai_n410_), .B(mai_mai_n71_), .Y(mai_mai_n854_));
  NA4        m0832(.A(mai_mai_n854_), .B(mai_mai_n853_), .C(mai_mai_n852_), .D(mai_mai_n622_), .Y(mai_mai_n855_));
  AN2        m0833(.A(mai_mai_n539_), .B(mai_mai_n47_), .Y(mai_mai_n856_));
  NA3        m0834(.A(mai_mai_n856_), .B(mai_mai_n500_), .C(mai_mai_n221_), .Y(mai_mai_n857_));
  AOI210     m0835(.A0(mai_mai_n466_), .A1(mai_mai_n464_), .B0(mai_mai_n584_), .Y(mai_mai_n858_));
  NO2        m0836(.A(mai_mai_n630_), .B(mai_mai_n104_), .Y(mai_mai_n859_));
  OAI210     m0837(.A0(mai_mai_n859_), .A1(mai_mai_n113_), .B0(mai_mai_n421_), .Y(mai_mai_n860_));
  INV        m0838(.A(mai_mai_n605_), .Y(mai_mai_n861_));
  NA3        m0839(.A(mai_mai_n861_), .B(mai_mai_n335_), .C(i_7_), .Y(mai_mai_n862_));
  NA4        m0840(.A(mai_mai_n862_), .B(mai_mai_n860_), .C(mai_mai_n858_), .D(mai_mai_n857_), .Y(mai_mai_n863_));
  NO4        m0841(.A(mai_mai_n863_), .B(mai_mai_n855_), .C(mai_mai_n850_), .D(mai_mai_n841_), .Y(mai_mai_n864_));
  NA4        m0842(.A(mai_mai_n864_), .B(mai_mai_n826_), .C(mai_mai_n820_), .D(mai_mai_n395_), .Y(mai3));
  NA2        m0843(.A(i_12_), .B(i_10_), .Y(mai_mai_n866_));
  NA2        m0844(.A(i_6_), .B(i_7_), .Y(mai_mai_n867_));
  NO2        m0845(.A(mai_mai_n867_), .B(i_0_), .Y(mai_mai_n868_));
  NO2        m0846(.A(i_11_), .B(mai_mai_n238_), .Y(mai_mai_n869_));
  OAI210     m0847(.A0(mai_mai_n868_), .A1(mai_mai_n295_), .B0(mai_mai_n869_), .Y(mai_mai_n870_));
  NO2        m0848(.A(mai_mai_n870_), .B(mai_mai_n197_), .Y(mai_mai_n871_));
  NO3        m0849(.A(mai_mai_n467_), .B(mai_mai_n91_), .C(mai_mai_n45_), .Y(mai_mai_n872_));
  OA210      m0850(.A0(mai_mai_n872_), .A1(mai_mai_n871_), .B0(mai_mai_n177_), .Y(mai_mai_n873_));
  NA2        m0851(.A(mai_mai_n853_), .B(mai_mai_n386_), .Y(mai_mai_n874_));
  NA2        m0852(.A(mai_mai_n874_), .B(mai_mai_n40_), .Y(mai_mai_n875_));
  NOi21      m0853(.An(mai_mai_n98_), .B(mai_mai_n782_), .Y(mai_mai_n876_));
  NO3        m0854(.A(mai_mai_n647_), .B(mai_mai_n471_), .C(mai_mai_n133_), .Y(mai_mai_n877_));
  NA2        m0855(.A(mai_mai_n424_), .B(mai_mai_n46_), .Y(mai_mai_n878_));
  AN2        m0856(.A(mai_mai_n469_), .B(mai_mai_n56_), .Y(mai_mai_n879_));
  NO3        m0857(.A(mai_mai_n879_), .B(mai_mai_n877_), .C(mai_mai_n876_), .Y(mai_mai_n880_));
  AOI210     m0858(.A0(mai_mai_n880_), .A1(mai_mai_n875_), .B0(mai_mai_n49_), .Y(mai_mai_n881_));
  NO4        m0859(.A(mai_mai_n391_), .B(mai_mai_n398_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n882_));
  NA2        m0860(.A(mai_mai_n189_), .B(mai_mai_n594_), .Y(mai_mai_n883_));
  NOi31      m0861(.An(mai_mai_n883_), .B(mai_mai_n882_), .C(mai_mai_n39_), .Y(mai_mai_n884_));
  NA2        m0862(.A(mai_mai_n729_), .B(mai_mai_n695_), .Y(mai_mai_n885_));
  NA2        m0863(.A(mai_mai_n342_), .B(mai_mai_n455_), .Y(mai_mai_n886_));
  OAI220     m0864(.A0(mai_mai_n886_), .A1(mai_mai_n885_), .B0(mai_mai_n884_), .B1(mai_mai_n64_), .Y(mai_mai_n887_));
  NOi21      m0865(.An(i_5_), .B(i_9_), .Y(mai_mai_n888_));
  NA2        m0866(.A(mai_mai_n888_), .B(mai_mai_n463_), .Y(mai_mai_n889_));
  BUFFER     m0867(.A(mai_mai_n272_), .Y(mai_mai_n890_));
  AOI210     m0868(.A0(mai_mai_n890_), .A1(mai_mai_n491_), .B0(mai_mai_n710_), .Y(mai_mai_n891_));
  NO3        m0869(.A(mai_mai_n427_), .B(mai_mai_n272_), .C(mai_mai_n74_), .Y(mai_mai_n892_));
  NO2        m0870(.A(mai_mai_n178_), .B(mai_mai_n150_), .Y(mai_mai_n893_));
  AOI210     m0871(.A0(mai_mai_n893_), .A1(mai_mai_n246_), .B0(mai_mai_n892_), .Y(mai_mai_n894_));
  OAI220     m0872(.A0(mai_mai_n894_), .A1(mai_mai_n184_), .B0(mai_mai_n891_), .B1(mai_mai_n889_), .Y(mai_mai_n895_));
  NO4        m0873(.A(mai_mai_n895_), .B(mai_mai_n887_), .C(mai_mai_n881_), .D(mai_mai_n873_), .Y(mai_mai_n896_));
  NA2        m0874(.A(mai_mai_n189_), .B(mai_mai_n24_), .Y(mai_mai_n897_));
  NA2        m0875(.A(mai_mai_n318_), .B(mai_mai_n131_), .Y(mai_mai_n898_));
  NO2        m0876(.A(mai_mai_n898_), .B(mai_mai_n413_), .Y(mai_mai_n899_));
  INV        m0877(.A(mai_mai_n899_), .Y(mai_mai_n900_));
  NO2        m0878(.A(mai_mai_n404_), .B(mai_mai_n299_), .Y(mai_mai_n901_));
  NA2        m0879(.A(mai_mai_n901_), .B(mai_mai_n732_), .Y(mai_mai_n902_));
  NA2        m0880(.A(mai_mai_n595_), .B(i_0_), .Y(mai_mai_n903_));
  NO4        m0881(.A(mai_mai_n604_), .B(mai_mai_n219_), .C(mai_mai_n431_), .D(mai_mai_n423_), .Y(mai_mai_n904_));
  NA2        m0882(.A(mai_mai_n904_), .B(i_11_), .Y(mai_mai_n905_));
  AN2        m0883(.A(mai_mai_n98_), .B(mai_mai_n245_), .Y(mai_mai_n906_));
  NA2        m0884(.A(mai_mai_n769_), .B(mai_mai_n336_), .Y(mai_mai_n907_));
  AOI210     m0885(.A0(mai_mai_n500_), .A1(mai_mai_n88_), .B0(mai_mai_n59_), .Y(mai_mai_n908_));
  OAI220     m0886(.A0(mai_mai_n908_), .A1(mai_mai_n907_), .B0(mai_mai_n678_), .B1(mai_mai_n561_), .Y(mai_mai_n909_));
  NO2        m0887(.A(mai_mai_n256_), .B(mai_mai_n155_), .Y(mai_mai_n910_));
  NA2        m0888(.A(i_0_), .B(i_10_), .Y(mai_mai_n911_));
  OAI210     m0889(.A0(mai_mai_n911_), .A1(mai_mai_n87_), .B0(mai_mai_n564_), .Y(mai_mai_n912_));
  NO4        m0890(.A(mai_mai_n116_), .B(mai_mai_n59_), .C(mai_mai_n688_), .D(i_5_), .Y(mai_mai_n913_));
  AO220      m0891(.A0(mai_mai_n913_), .A1(mai_mai_n912_), .B0(mai_mai_n910_), .B1(i_6_), .Y(mai_mai_n914_));
  AOI220     m0892(.A0(mai_mai_n342_), .A1(mai_mai_n100_), .B0(mai_mai_n189_), .B1(mai_mai_n85_), .Y(mai_mai_n915_));
  NA2        m0893(.A(mai_mai_n589_), .B(i_4_), .Y(mai_mai_n916_));
  NA2        m0894(.A(mai_mai_n192_), .B(mai_mai_n207_), .Y(mai_mai_n917_));
  OAI220     m0895(.A0(mai_mai_n917_), .A1(mai_mai_n907_), .B0(mai_mai_n916_), .B1(mai_mai_n915_), .Y(mai_mai_n918_));
  NO4        m0896(.A(mai_mai_n918_), .B(mai_mai_n914_), .C(mai_mai_n909_), .D(mai_mai_n906_), .Y(mai_mai_n919_));
  NA4        m0897(.A(mai_mai_n919_), .B(mai_mai_n905_), .C(mai_mai_n902_), .D(mai_mai_n900_), .Y(mai_mai_n920_));
  NO2        m0898(.A(mai_mai_n105_), .B(mai_mai_n37_), .Y(mai_mai_n921_));
  NA2        m0899(.A(i_11_), .B(i_9_), .Y(mai_mai_n922_));
  NO3        m0900(.A(i_12_), .B(mai_mai_n922_), .C(mai_mai_n621_), .Y(mai_mai_n923_));
  AN2        m0901(.A(mai_mai_n923_), .B(mai_mai_n921_), .Y(mai_mai_n924_));
  NO2        m0902(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n925_));
  NA2        m0903(.A(mai_mai_n409_), .B(mai_mai_n182_), .Y(mai_mai_n926_));
  NA3        m0904(.A(mai_mai_n926_), .B(mai_mai_n476_), .C(mai_mai_n162_), .Y(mai_mai_n927_));
  NO2        m0905(.A(mai_mai_n922_), .B(mai_mai_n74_), .Y(mai_mai_n928_));
  NO2        m0906(.A(mai_mai_n178_), .B(i_0_), .Y(mai_mai_n929_));
  INV        m0907(.A(mai_mai_n929_), .Y(mai_mai_n930_));
  NA2        m0908(.A(mai_mai_n489_), .B(mai_mai_n232_), .Y(mai_mai_n931_));
  AOI210     m0909(.A0(mai_mai_n385_), .A1(mai_mai_n42_), .B0(mai_mai_n420_), .Y(mai_mai_n932_));
  OAI220     m0910(.A0(mai_mai_n932_), .A1(mai_mai_n889_), .B0(mai_mai_n931_), .B1(mai_mai_n930_), .Y(mai_mai_n933_));
  NO3        m0911(.A(mai_mai_n933_), .B(mai_mai_n927_), .C(mai_mai_n924_), .Y(mai_mai_n934_));
  NA2        m0912(.A(mai_mai_n677_), .B(mai_mai_n123_), .Y(mai_mai_n935_));
  NO2        m0913(.A(i_6_), .B(mai_mai_n935_), .Y(mai_mai_n936_));
  AOI210     m0914(.A0(mai_mai_n465_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n937_));
  NA2        m0915(.A(mai_mai_n174_), .B(mai_mai_n105_), .Y(mai_mai_n938_));
  NOi32      m0916(.An(mai_mai_n937_), .Bn(mai_mai_n192_), .C(mai_mai_n938_), .Y(mai_mai_n939_));
  NO2        m0917(.A(mai_mai_n939_), .B(mai_mai_n936_), .Y(mai_mai_n940_));
  NOi21      m0918(.An(i_7_), .B(i_5_), .Y(mai_mai_n941_));
  OR2        m0919(.A(mai_mai_n938_), .B(mai_mai_n537_), .Y(mai_mai_n942_));
  NO3        m0920(.A(mai_mai_n416_), .B(mai_mai_n374_), .C(mai_mai_n371_), .Y(mai_mai_n943_));
  NO2        m0921(.A(mai_mai_n266_), .B(mai_mai_n325_), .Y(mai_mai_n944_));
  NO2        m0922(.A(mai_mai_n748_), .B(mai_mai_n261_), .Y(mai_mai_n945_));
  AOI210     m0923(.A0(mai_mai_n945_), .A1(mai_mai_n944_), .B0(mai_mai_n943_), .Y(mai_mai_n946_));
  NA4        m0924(.A(mai_mai_n946_), .B(mai_mai_n942_), .C(mai_mai_n940_), .D(mai_mai_n934_), .Y(mai_mai_n947_));
  NO2        m0925(.A(mai_mai_n897_), .B(mai_mai_n241_), .Y(mai_mai_n948_));
  AN2        m0926(.A(mai_mai_n341_), .B(mai_mai_n336_), .Y(mai_mai_n949_));
  AO220      m0927(.A0(mai_mai_n949_), .A1(mai_mai_n893_), .B0(mai_mai_n357_), .B1(mai_mai_n27_), .Y(mai_mai_n950_));
  OAI210     m0928(.A0(mai_mai_n950_), .A1(mai_mai_n948_), .B0(i_10_), .Y(mai_mai_n951_));
  NO2        m0929(.A(mai_mai_n866_), .B(mai_mai_n324_), .Y(mai_mai_n952_));
  OA210      m0930(.A0(mai_mai_n489_), .A1(mai_mai_n225_), .B0(mai_mai_n488_), .Y(mai_mai_n953_));
  NA2        m0931(.A(mai_mai_n952_), .B(mai_mai_n928_), .Y(mai_mai_n954_));
  NO2        m0932(.A(mai_mai_n259_), .B(mai_mai_n47_), .Y(mai_mai_n955_));
  NO2        m0933(.A(mai_mai_n955_), .B(mai_mai_n191_), .Y(mai_mai_n956_));
  NA2        m0934(.A(mai_mai_n956_), .B(mai_mai_n489_), .Y(mai_mai_n957_));
  NA2        m0935(.A(mai_mai_n722_), .B(mai_mai_n568_), .Y(mai_mai_n958_));
  NAi21      m0936(.An(i_9_), .B(i_5_), .Y(mai_mai_n959_));
  NO2        m0937(.A(mai_mai_n959_), .B(mai_mai_n416_), .Y(mai_mai_n960_));
  NO2        m0938(.A(mai_mai_n617_), .B(mai_mai_n107_), .Y(mai_mai_n961_));
  AOI220     m0939(.A0(mai_mai_n961_), .A1(i_0_), .B0(mai_mai_n960_), .B1(mai_mai_n639_), .Y(mai_mai_n962_));
  OAI220     m0940(.A0(mai_mai_n962_), .A1(mai_mai_n87_), .B0(mai_mai_n958_), .B1(mai_mai_n175_), .Y(mai_mai_n963_));
  NO2        m0941(.A(mai_mai_n963_), .B(mai_mai_n542_), .Y(mai_mai_n964_));
  NA4        m0942(.A(mai_mai_n964_), .B(mai_mai_n957_), .C(mai_mai_n954_), .D(mai_mai_n951_), .Y(mai_mai_n965_));
  NO3        m0943(.A(mai_mai_n965_), .B(mai_mai_n947_), .C(mai_mai_n920_), .Y(mai_mai_n966_));
  NO2        m0944(.A(i_0_), .B(mai_mai_n748_), .Y(mai_mai_n967_));
  NA2        m0945(.A(mai_mai_n74_), .B(mai_mai_n45_), .Y(mai_mai_n968_));
  NA2        m0946(.A(mai_mai_n911_), .B(mai_mai_n968_), .Y(mai_mai_n969_));
  NO3        m0947(.A(mai_mai_n107_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n970_));
  AO220      m0948(.A0(mai_mai_n970_), .A1(mai_mai_n969_), .B0(mai_mai_n967_), .B1(mai_mai_n177_), .Y(mai_mai_n971_));
  AOI210     m0949(.A0(mai_mai_n822_), .A1(mai_mai_n708_), .B0(mai_mai_n938_), .Y(mai_mai_n972_));
  AOI210     m0950(.A0(mai_mai_n971_), .A1(mai_mai_n359_), .B0(mai_mai_n972_), .Y(mai_mai_n973_));
  NA2        m0951(.A(mai_mai_n757_), .B(mai_mai_n148_), .Y(mai_mai_n974_));
  INV        m0952(.A(mai_mai_n974_), .Y(mai_mai_n975_));
  NA3        m0953(.A(mai_mai_n975_), .B(mai_mai_n695_), .C(mai_mai_n74_), .Y(mai_mai_n976_));
  NO2        m0954(.A(mai_mai_n839_), .B(mai_mai_n416_), .Y(mai_mai_n977_));
  NA3        m0955(.A(mai_mai_n868_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n978_));
  NA2        m0956(.A(mai_mai_n869_), .B(i_9_), .Y(mai_mai_n979_));
  AOI210     m0957(.A0(mai_mai_n978_), .A1(mai_mai_n516_), .B0(mai_mai_n979_), .Y(mai_mai_n980_));
  OAI210     m0958(.A0(mai_mai_n246_), .A1(i_9_), .B0(mai_mai_n231_), .Y(mai_mai_n981_));
  AOI210     m0959(.A0(mai_mai_n981_), .A1(mai_mai_n903_), .B0(mai_mai_n155_), .Y(mai_mai_n982_));
  NO3        m0960(.A(mai_mai_n982_), .B(mai_mai_n980_), .C(mai_mai_n977_), .Y(mai_mai_n983_));
  NA3        m0961(.A(mai_mai_n983_), .B(mai_mai_n976_), .C(mai_mai_n973_), .Y(mai_mai_n984_));
  NA2        m0962(.A(mai_mai_n949_), .B(mai_mai_n387_), .Y(mai_mai_n985_));
  AOI210     m0963(.A0(mai_mai_n306_), .A1(mai_mai_n164_), .B0(mai_mai_n985_), .Y(mai_mai_n986_));
  NA3        m0964(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n987_));
  NA2        m0965(.A(mai_mai_n925_), .B(mai_mai_n505_), .Y(mai_mai_n988_));
  AOI210     m0966(.A0(mai_mai_n987_), .A1(mai_mai_n164_), .B0(mai_mai_n988_), .Y(mai_mai_n989_));
  NO2        m0967(.A(mai_mai_n989_), .B(mai_mai_n986_), .Y(mai_mai_n990_));
  NO3        m0968(.A(mai_mai_n911_), .B(mai_mai_n888_), .C(mai_mai_n194_), .Y(mai_mai_n991_));
  AOI220     m0969(.A0(mai_mai_n991_), .A1(i_11_), .B0(mai_mai_n590_), .B1(mai_mai_n76_), .Y(mai_mai_n992_));
  NO3        m0970(.A(mai_mai_n213_), .B(mai_mai_n398_), .C(i_0_), .Y(mai_mai_n993_));
  OAI210     m0971(.A0(mai_mai_n993_), .A1(mai_mai_n77_), .B0(i_13_), .Y(mai_mai_n994_));
  INV        m0972(.A(mai_mai_n221_), .Y(mai_mai_n995_));
  OAI220     m0973(.A0(mai_mai_n554_), .A1(mai_mai_n141_), .B0(mai_mai_n661_), .B1(mai_mai_n634_), .Y(mai_mai_n996_));
  NA3        m0974(.A(mai_mai_n996_), .B(mai_mai_n411_), .C(mai_mai_n995_), .Y(mai_mai_n997_));
  NA4        m0975(.A(mai_mai_n997_), .B(mai_mai_n994_), .C(mai_mai_n992_), .D(mai_mai_n990_), .Y(mai_mai_n998_));
  AOI220     m0976(.A0(mai_mai_n941_), .A1(mai_mai_n505_), .B0(mai_mai_n868_), .B1(mai_mai_n165_), .Y(mai_mai_n999_));
  NA2        m0977(.A(mai_mai_n362_), .B(mai_mai_n179_), .Y(mai_mai_n1000_));
  OR2        m0978(.A(mai_mai_n1000_), .B(mai_mai_n999_), .Y(mai_mai_n1001_));
  AOI210     m0979(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n178_), .Y(mai_mai_n1002_));
  NA2        m0980(.A(mai_mai_n1002_), .B(mai_mai_n953_), .Y(mai_mai_n1003_));
  NA3        m0981(.A(mai_mai_n631_), .B(mai_mai_n189_), .C(mai_mai_n85_), .Y(mai_mai_n1004_));
  INV        m0982(.A(mai_mai_n1004_), .Y(mai_mai_n1005_));
  NO3        m0983(.A(mai_mai_n878_), .B(mai_mai_n55_), .C(mai_mai_n49_), .Y(mai_mai_n1006_));
  NA2        m0984(.A(mai_mai_n510_), .B(mai_mai_n503_), .Y(mai_mai_n1007_));
  NO3        m0985(.A(mai_mai_n1007_), .B(mai_mai_n1006_), .C(mai_mai_n1005_), .Y(mai_mai_n1008_));
  NA3        m0986(.A(mai_mai_n404_), .B(mai_mai_n174_), .C(mai_mai_n173_), .Y(mai_mai_n1009_));
  NA3        m0987(.A(mai_mai_n404_), .B(mai_mai_n343_), .C(mai_mai_n223_), .Y(mai_mai_n1010_));
  OAI210     m0988(.A0(mai_mai_n883_), .A1(mai_mai_n665_), .B0(mai_mai_n1010_), .Y(mai_mai_n1011_));
  NOi31      m0989(.An(mai_mai_n403_), .B(mai_mai_n968_), .C(mai_mai_n241_), .Y(mai_mai_n1012_));
  NO3        m0990(.A(mai_mai_n922_), .B(mai_mai_n221_), .C(mai_mai_n194_), .Y(mai_mai_n1013_));
  NO4        m0991(.A(mai_mai_n1013_), .B(mai_mai_n1012_), .C(mai_mai_n1011_), .D(mai_mai_n1074_), .Y(mai_mai_n1014_));
  NA4        m0992(.A(mai_mai_n1014_), .B(mai_mai_n1008_), .C(mai_mai_n1003_), .D(mai_mai_n1001_), .Y(mai_mai_n1015_));
  INV        m0993(.A(mai_mai_n633_), .Y(mai_mai_n1016_));
  NO3        m0994(.A(mai_mai_n1016_), .B(mai_mai_n580_), .C(mai_mai_n356_), .Y(mai_mai_n1017_));
  NO2        m0995(.A(mai_mai_n87_), .B(i_5_), .Y(mai_mai_n1018_));
  NA3        m0996(.A(mai_mai_n869_), .B(mai_mai_n111_), .C(mai_mai_n126_), .Y(mai_mai_n1019_));
  INV        m0997(.A(mai_mai_n1019_), .Y(mai_mai_n1020_));
  AOI210     m0998(.A0(mai_mai_n1020_), .A1(mai_mai_n1018_), .B0(mai_mai_n1017_), .Y(mai_mai_n1021_));
  NAi21      m0999(.An(mai_mai_n243_), .B(mai_mai_n244_), .Y(mai_mai_n1022_));
  NO4        m1000(.A(mai_mai_n241_), .B(mai_mai_n213_), .C(i_0_), .D(i_12_), .Y(mai_mai_n1023_));
  AOI220     m1001(.A0(mai_mai_n1023_), .A1(mai_mai_n1022_), .B0(mai_mai_n816_), .B1(mai_mai_n179_), .Y(mai_mai_n1024_));
  AN2        m1002(.A(mai_mai_n911_), .B(mai_mai_n155_), .Y(mai_mai_n1025_));
  NO4        m1003(.A(mai_mai_n1025_), .B(i_12_), .C(mai_mai_n665_), .D(mai_mai_n133_), .Y(mai_mai_n1026_));
  NA2        m1004(.A(mai_mai_n1026_), .B(mai_mai_n221_), .Y(mai_mai_n1027_));
  NA3        m1005(.A(mai_mai_n100_), .B(mai_mai_n594_), .C(i_11_), .Y(mai_mai_n1028_));
  NO2        m1006(.A(mai_mai_n1028_), .B(mai_mai_n157_), .Y(mai_mai_n1029_));
  NA2        m1007(.A(mai_mai_n941_), .B(mai_mai_n487_), .Y(mai_mai_n1030_));
  NO2        m1008(.A(mai_mai_n1030_), .B(mai_mai_n696_), .Y(mai_mai_n1031_));
  AOI210     m1009(.A0(mai_mai_n1031_), .A1(mai_mai_n929_), .B0(mai_mai_n1029_), .Y(mai_mai_n1032_));
  NA4        m1010(.A(mai_mai_n1032_), .B(mai_mai_n1027_), .C(mai_mai_n1024_), .D(mai_mai_n1021_), .Y(mai_mai_n1033_));
  NO4        m1011(.A(mai_mai_n1033_), .B(mai_mai_n1015_), .C(mai_mai_n998_), .D(mai_mai_n984_), .Y(mai_mai_n1034_));
  OAI210     m1012(.A0(mai_mai_n842_), .A1(mai_mai_n835_), .B0(mai_mai_n37_), .Y(mai_mai_n1035_));
  NA3        m1013(.A(mai_mai_n937_), .B(mai_mai_n382_), .C(i_5_), .Y(mai_mai_n1036_));
  NA3        m1014(.A(mai_mai_n1036_), .B(mai_mai_n1035_), .C(mai_mai_n629_), .Y(mai_mai_n1037_));
  NA2        m1015(.A(mai_mai_n1037_), .B(mai_mai_n210_), .Y(mai_mai_n1038_));
  AN2        m1016(.A(mai_mai_n720_), .B(mai_mai_n383_), .Y(mai_mai_n1039_));
  NA2        m1017(.A(mai_mai_n190_), .B(mai_mai_n192_), .Y(mai_mai_n1040_));
  AO210      m1018(.A0(mai_mai_n1039_), .A1(mai_mai_n33_), .B0(mai_mai_n1040_), .Y(mai_mai_n1041_));
  OAI210     m1019(.A0(mai_mai_n633_), .A1(mai_mai_n631_), .B0(mai_mai_n324_), .Y(mai_mai_n1042_));
  NAi31      m1020(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n1043_));
  AOI210     m1021(.A0(mai_mai_n119_), .A1(mai_mai_n71_), .B0(mai_mai_n1043_), .Y(mai_mai_n1044_));
  NO2        m1022(.A(mai_mai_n1044_), .B(mai_mai_n662_), .Y(mai_mai_n1045_));
  NA3        m1023(.A(mai_mai_n1045_), .B(mai_mai_n1042_), .C(mai_mai_n1041_), .Y(mai_mai_n1046_));
  NO2        m1024(.A(mai_mai_n479_), .B(mai_mai_n272_), .Y(mai_mai_n1047_));
  NO4        m1025(.A(mai_mai_n234_), .B(mai_mai_n147_), .C(mai_mai_n699_), .D(mai_mai_n37_), .Y(mai_mai_n1048_));
  NO3        m1026(.A(mai_mai_n1048_), .B(mai_mai_n1047_), .C(mai_mai_n904_), .Y(mai_mai_n1049_));
  OAI210     m1027(.A0(mai_mai_n1028_), .A1(mai_mai_n150_), .B0(mai_mai_n1049_), .Y(mai_mai_n1050_));
  AOI210     m1028(.A0(mai_mai_n1046_), .A1(mai_mai_n49_), .B0(mai_mai_n1050_), .Y(mai_mai_n1051_));
  AOI210     m1029(.A0(mai_mai_n1051_), .A1(mai_mai_n1038_), .B0(mai_mai_n74_), .Y(mai_mai_n1052_));
  NO2        m1030(.A(mai_mai_n587_), .B(mai_mai_n394_), .Y(mai_mai_n1053_));
  NO2        m1031(.A(mai_mai_n1053_), .B(mai_mai_n777_), .Y(mai_mai_n1054_));
  NA2        m1032(.A(mai_mai_n266_), .B(mai_mai_n58_), .Y(mai_mai_n1055_));
  AOI220     m1033(.A0(mai_mai_n1055_), .A1(mai_mai_n77_), .B0(mai_mai_n357_), .B1(mai_mai_n258_), .Y(mai_mai_n1056_));
  NO2        m1034(.A(mai_mai_n1056_), .B(mai_mai_n238_), .Y(mai_mai_n1057_));
  NA3        m1035(.A(mai_mai_n98_), .B(mai_mai_n313_), .C(mai_mai_n31_), .Y(mai_mai_n1058_));
  INV        m1036(.A(mai_mai_n1058_), .Y(mai_mai_n1059_));
  NO2        m1037(.A(mai_mai_n1059_), .B(mai_mai_n1057_), .Y(mai_mai_n1060_));
  OAI210     m1038(.A0(mai_mai_n274_), .A1(mai_mai_n160_), .B0(mai_mai_n88_), .Y(mai_mai_n1061_));
  NO2        m1039(.A(mai_mai_n1061_), .B(i_11_), .Y(mai_mai_n1062_));
  NO4        m1040(.A(mai_mai_n959_), .B(mai_mai_n493_), .C(mai_mai_n255_), .D(mai_mai_n254_), .Y(mai_mai_n1063_));
  NO2        m1041(.A(mai_mai_n1063_), .B(mai_mai_n584_), .Y(mai_mai_n1064_));
  NO2        m1042(.A(mai_mai_n1064_), .B(mai_mai_n41_), .Y(mai_mai_n1065_));
  NO2        m1043(.A(mai_mai_n1065_), .B(mai_mai_n1062_), .Y(mai_mai_n1066_));
  OAI210     m1044(.A0(mai_mai_n1060_), .A1(i_4_), .B0(mai_mai_n1066_), .Y(mai_mai_n1067_));
  NO3        m1045(.A(mai_mai_n1067_), .B(mai_mai_n1054_), .C(mai_mai_n1052_), .Y(mai_mai_n1068_));
  NA4        m1046(.A(mai_mai_n1068_), .B(mai_mai_n1034_), .C(mai_mai_n966_), .D(mai_mai_n896_), .Y(mai4));
  INV        m1047(.A(mai_mai_n721_), .Y(mai_mai_n1072_));
  INV        m1048(.A(i_2_), .Y(mai_mai_n1073_));
  INV        m1049(.A(mai_mai_n1009_), .Y(mai_mai_n1074_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n51_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(men_men_n81_), .B(men_men_n58_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_9_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_7_), .Y(men_men_n84_));
  NO3        u0062(.A(men_men_n84_), .B(men_men_n83_), .C(men_men_n63_), .Y(men_men_n85_));
  INV        u0063(.A(i_6_), .Y(men_men_n86_));
  OR4        u0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n87_));
  INV        u0065(.A(men_men_n87_), .Y(men_men_n88_));
  NO2        u0066(.A(i_2_), .B(i_7_), .Y(men_men_n89_));
  AOI210     u0067(.A0(men_men_n88_), .A1(men_men_n86_), .B0(men_men_n89_), .Y(men_men_n90_));
  OAI210     u0068(.A0(men_men_n85_), .A1(men_men_n82_), .B0(men_men_n90_), .Y(men_men_n91_));
  NAi21      u0069(.An(i_6_), .B(i_10_), .Y(men_men_n92_));
  NA2        u0070(.A(i_6_), .B(i_9_), .Y(men_men_n93_));
  AOI210     u0071(.A0(men_men_n93_), .A1(men_men_n92_), .B0(men_men_n63_), .Y(men_men_n94_));
  NA2        u0072(.A(i_2_), .B(i_6_), .Y(men_men_n95_));
  NO3        u0073(.A(men_men_n95_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n96_));
  NO2        u0074(.A(men_men_n96_), .B(men_men_n94_), .Y(men_men_n97_));
  AOI210     u0075(.A0(men_men_n97_), .A1(men_men_n91_), .B0(men_men_n80_), .Y(men_men_n98_));
  AN3        u0076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n99_));
  NAi21      u0077(.An(i_6_), .B(i_11_), .Y(men_men_n100_));
  NO2        u0078(.A(i_5_), .B(i_8_), .Y(men_men_n101_));
  NOi21      u0079(.An(men_men_n101_), .B(men_men_n100_), .Y(men_men_n102_));
  AOI220     u0080(.A0(men_men_n102_), .A1(men_men_n62_), .B0(men_men_n99_), .B1(men_men_n32_), .Y(men_men_n103_));
  INV        u0081(.A(i_7_), .Y(men_men_n104_));
  NA2        u0082(.A(men_men_n47_), .B(men_men_n104_), .Y(men_men_n105_));
  NO2        u0083(.A(i_0_), .B(i_5_), .Y(men_men_n106_));
  NO2        u0084(.A(men_men_n106_), .B(men_men_n86_), .Y(men_men_n107_));
  NA2        u0085(.A(i_12_), .B(i_3_), .Y(men_men_n108_));
  INV        u0086(.A(men_men_n108_), .Y(men_men_n109_));
  NA3        u0087(.A(men_men_n109_), .B(men_men_n107_), .C(men_men_n105_), .Y(men_men_n110_));
  NAi21      u0088(.An(i_7_), .B(i_11_), .Y(men_men_n111_));
  NO3        u0089(.A(men_men_n111_), .B(men_men_n92_), .C(men_men_n54_), .Y(men_men_n112_));
  AN2        u0090(.A(i_2_), .B(i_10_), .Y(men_men_n113_));
  NO2        u0091(.A(men_men_n113_), .B(i_7_), .Y(men_men_n114_));
  OR2        u0092(.A(men_men_n80_), .B(men_men_n58_), .Y(men_men_n115_));
  NO2        u0093(.A(i_8_), .B(men_men_n104_), .Y(men_men_n116_));
  NO3        u0094(.A(men_men_n116_), .B(men_men_n115_), .C(men_men_n114_), .Y(men_men_n117_));
  NA2        u0095(.A(i_12_), .B(i_7_), .Y(men_men_n118_));
  NO2        u0096(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n119_));
  NA2        u0097(.A(i_11_), .B(i_12_), .Y(men_men_n120_));
  INV        u0098(.A(men_men_n120_), .Y(men_men_n121_));
  NO2        u0099(.A(men_men_n121_), .B(men_men_n117_), .Y(men_men_n122_));
  NAi41      u0100(.An(men_men_n112_), .B(men_men_n122_), .C(men_men_n110_), .D(men_men_n103_), .Y(men_men_n123_));
  NOi21      u0101(.An(i_1_), .B(i_5_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(i_11_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n104_), .B(men_men_n37_), .Y(men_men_n126_));
  NA2        u0104(.A(i_7_), .B(men_men_n25_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n128_));
  NO2        u0106(.A(men_men_n128_), .B(men_men_n47_), .Y(men_men_n129_));
  NA2        u0107(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n130_));
  NAi21      u0108(.An(i_3_), .B(i_8_), .Y(men_men_n131_));
  NA2        u0109(.A(men_men_n131_), .B(men_men_n62_), .Y(men_men_n132_));
  NOi31      u0110(.An(men_men_n132_), .B(men_men_n130_), .C(men_men_n129_), .Y(men_men_n133_));
  NO2        u0111(.A(i_1_), .B(men_men_n86_), .Y(men_men_n134_));
  NO2        u0112(.A(i_6_), .B(i_5_), .Y(men_men_n135_));
  NA2        u0113(.A(men_men_n135_), .B(i_3_), .Y(men_men_n136_));
  AO210      u0114(.A0(men_men_n136_), .A1(men_men_n48_), .B0(men_men_n134_), .Y(men_men_n137_));
  OAI220     u0115(.A0(men_men_n137_), .A1(men_men_n111_), .B0(men_men_n133_), .B1(men_men_n125_), .Y(men_men_n138_));
  NO3        u0116(.A(men_men_n138_), .B(men_men_n123_), .C(men_men_n98_), .Y(men_men_n139_));
  NA3        u0117(.A(men_men_n139_), .B(men_men_n79_), .C(men_men_n56_), .Y(men2));
  NO2        u0118(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n141_));
  NA2        u0119(.A(i_6_), .B(men_men_n25_), .Y(men_men_n142_));
  NA2        u0120(.A(men_men_n142_), .B(men_men_n141_), .Y(men_men_n143_));
  NA4        u0121(.A(men_men_n143_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n30_), .Y(men0));
  AN2        u0122(.A(i_8_), .B(i_7_), .Y(men_men_n145_));
  NA2        u0123(.A(men_men_n145_), .B(i_6_), .Y(men_men_n146_));
  NO2        u0124(.A(i_12_), .B(i_13_), .Y(men_men_n147_));
  NAi21      u0125(.An(i_5_), .B(i_11_), .Y(men_men_n148_));
  NOi21      u0126(.An(men_men_n147_), .B(men_men_n148_), .Y(men_men_n149_));
  NO2        u0127(.A(i_0_), .B(i_1_), .Y(men_men_n150_));
  NA2        u0128(.A(i_2_), .B(i_3_), .Y(men_men_n151_));
  NO2        u0129(.A(men_men_n151_), .B(i_4_), .Y(men_men_n152_));
  NA3        u0130(.A(men_men_n152_), .B(men_men_n150_), .C(men_men_n149_), .Y(men_men_n153_));
  OR2        u0131(.A(men_men_n153_), .B(men_men_n25_), .Y(men_men_n154_));
  AN2        u0132(.A(men_men_n147_), .B(men_men_n83_), .Y(men_men_n155_));
  NO2        u0133(.A(men_men_n155_), .B(men_men_n27_), .Y(men_men_n156_));
  NA2        u0134(.A(i_1_), .B(i_5_), .Y(men_men_n157_));
  NO2        u0135(.A(men_men_n73_), .B(men_men_n47_), .Y(men_men_n158_));
  NA2        u0136(.A(men_men_n158_), .B(men_men_n36_), .Y(men_men_n159_));
  NO3        u0137(.A(men_men_n159_), .B(men_men_n157_), .C(men_men_n156_), .Y(men_men_n160_));
  OR2        u0138(.A(i_0_), .B(i_1_), .Y(men_men_n161_));
  NO3        u0139(.A(men_men_n161_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n162_));
  NAi32      u0140(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n163_));
  NAi21      u0141(.An(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  NOi21      u0142(.An(i_4_), .B(i_10_), .Y(men_men_n165_));
  NA2        u0143(.A(men_men_n165_), .B(men_men_n40_), .Y(men_men_n166_));
  NO2        u0144(.A(i_3_), .B(i_5_), .Y(men_men_n167_));
  NO3        u0145(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n168_));
  NA2        u0146(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  OAI210     u0147(.A0(men_men_n169_), .A1(men_men_n166_), .B0(men_men_n164_), .Y(men_men_n170_));
  NO2        u0148(.A(men_men_n170_), .B(men_men_n160_), .Y(men_men_n171_));
  AOI210     u0149(.A0(men_men_n171_), .A1(men_men_n154_), .B0(men_men_n146_), .Y(men_men_n172_));
  NA3        u0150(.A(men_men_n73_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n173_));
  NA2        u0151(.A(i_3_), .B(men_men_n49_), .Y(men_men_n174_));
  NOi21      u0152(.An(i_4_), .B(i_9_), .Y(men_men_n175_));
  NOi21      u0153(.An(i_11_), .B(i_13_), .Y(men_men_n176_));
  NA2        u0154(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  OR2        u0155(.A(men_men_n177_), .B(men_men_n174_), .Y(men_men_n178_));
  NO2        u0156(.A(i_4_), .B(i_5_), .Y(men_men_n179_));
  NAi21      u0157(.An(i_12_), .B(i_11_), .Y(men_men_n180_));
  NO2        u0158(.A(men_men_n180_), .B(i_13_), .Y(men_men_n181_));
  NA3        u0159(.A(men_men_n181_), .B(men_men_n179_), .C(men_men_n83_), .Y(men_men_n182_));
  AOI210     u0160(.A0(men_men_n182_), .A1(men_men_n178_), .B0(men_men_n173_), .Y(men_men_n183_));
  NO2        u0161(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n184_));
  NA2        u0162(.A(men_men_n184_), .B(men_men_n47_), .Y(men_men_n185_));
  NA2        u0163(.A(men_men_n36_), .B(i_5_), .Y(men_men_n186_));
  NAi31      u0164(.An(men_men_n186_), .B(men_men_n155_), .C(i_11_), .Y(men_men_n187_));
  NA2        u0165(.A(i_3_), .B(i_5_), .Y(men_men_n188_));
  OR2        u0166(.A(men_men_n188_), .B(men_men_n177_), .Y(men_men_n189_));
  AOI210     u0167(.A0(men_men_n189_), .A1(men_men_n187_), .B0(men_men_n185_), .Y(men_men_n190_));
  NO2        u0168(.A(men_men_n73_), .B(i_5_), .Y(men_men_n191_));
  NO2        u0169(.A(i_13_), .B(i_10_), .Y(men_men_n192_));
  NA3        u0170(.A(men_men_n192_), .B(men_men_n191_), .C(men_men_n45_), .Y(men_men_n193_));
  NO2        u0171(.A(i_2_), .B(i_1_), .Y(men_men_n194_));
  NA2        u0172(.A(men_men_n194_), .B(i_3_), .Y(men_men_n195_));
  NAi21      u0173(.An(i_4_), .B(i_12_), .Y(men_men_n196_));
  NO4        u0174(.A(men_men_n196_), .B(men_men_n195_), .C(men_men_n193_), .D(men_men_n25_), .Y(men_men_n197_));
  NO3        u0175(.A(men_men_n197_), .B(men_men_n190_), .C(men_men_n183_), .Y(men_men_n198_));
  INV        u0176(.A(i_8_), .Y(men_men_n199_));
  NO2        u0177(.A(men_men_n199_), .B(i_7_), .Y(men_men_n200_));
  NA2        u0178(.A(men_men_n200_), .B(i_6_), .Y(men_men_n201_));
  NO3        u0179(.A(i_3_), .B(men_men_n86_), .C(men_men_n49_), .Y(men_men_n202_));
  NA2        u0180(.A(men_men_n202_), .B(men_men_n116_), .Y(men_men_n203_));
  NO3        u0181(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n204_));
  NA3        u0182(.A(men_men_n204_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n205_));
  NO3        u0183(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n206_));
  OAI210     u0184(.A0(men_men_n99_), .A1(i_12_), .B0(men_men_n206_), .Y(men_men_n207_));
  AOI210     u0185(.A0(men_men_n207_), .A1(men_men_n205_), .B0(men_men_n203_), .Y(men_men_n208_));
  NO2        u0186(.A(i_3_), .B(i_8_), .Y(men_men_n209_));
  NO3        u0187(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n210_));
  NA3        u0188(.A(men_men_n210_), .B(men_men_n209_), .C(men_men_n40_), .Y(men_men_n211_));
  NO2        u0189(.A(men_men_n106_), .B(men_men_n58_), .Y(men_men_n212_));
  NA2        u0190(.A(men_men_n212_), .B(men_men_n161_), .Y(men_men_n213_));
  NO2        u0191(.A(i_13_), .B(i_9_), .Y(men_men_n214_));
  NA3        u0192(.A(men_men_n214_), .B(i_6_), .C(men_men_n199_), .Y(men_men_n215_));
  NAi21      u0193(.An(i_12_), .B(i_3_), .Y(men_men_n216_));
  OR2        u0194(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NO2        u0195(.A(men_men_n45_), .B(i_5_), .Y(men_men_n218_));
  NO3        u0196(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n219_));
  NA3        u0197(.A(men_men_n219_), .B(men_men_n218_), .C(i_10_), .Y(men_men_n220_));
  OAI220     u0198(.A0(men_men_n220_), .A1(men_men_n217_), .B0(men_men_n213_), .B1(men_men_n211_), .Y(men_men_n221_));
  AOI210     u0199(.A0(men_men_n221_), .A1(i_7_), .B0(men_men_n208_), .Y(men_men_n222_));
  OAI220     u0200(.A0(men_men_n222_), .A1(i_4_), .B0(men_men_n201_), .B1(men_men_n198_), .Y(men_men_n223_));
  NAi21      u0201(.An(i_12_), .B(i_7_), .Y(men_men_n224_));
  NA3        u0202(.A(i_13_), .B(men_men_n199_), .C(i_10_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  NA2        u0204(.A(i_0_), .B(i_5_), .Y(men_men_n227_));
  NA2        u0205(.A(men_men_n227_), .B(men_men_n107_), .Y(men_men_n228_));
  OAI220     u0206(.A0(men_men_n228_), .A1(men_men_n195_), .B0(men_men_n185_), .B1(men_men_n136_), .Y(men_men_n229_));
  NAi31      u0207(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n36_), .B(i_13_), .Y(men_men_n231_));
  NO2        u0209(.A(men_men_n73_), .B(men_men_n26_), .Y(men_men_n232_));
  NO2        u0210(.A(men_men_n47_), .B(men_men_n63_), .Y(men_men_n233_));
  NA3        u0211(.A(men_men_n233_), .B(men_men_n232_), .C(men_men_n231_), .Y(men_men_n234_));
  INV        u0212(.A(i_13_), .Y(men_men_n235_));
  NO2        u0213(.A(i_12_), .B(men_men_n235_), .Y(men_men_n236_));
  NA3        u0214(.A(men_men_n236_), .B(men_men_n204_), .C(men_men_n202_), .Y(men_men_n237_));
  OAI210     u0215(.A0(men_men_n234_), .A1(men_men_n230_), .B0(men_men_n237_), .Y(men_men_n238_));
  AOI220     u0216(.A0(men_men_n238_), .A1(men_men_n145_), .B0(men_men_n229_), .B1(men_men_n226_), .Y(men_men_n239_));
  NO2        u0217(.A(i_12_), .B(men_men_n37_), .Y(men_men_n240_));
  NO2        u0218(.A(men_men_n188_), .B(i_4_), .Y(men_men_n241_));
  NA2        u0219(.A(men_men_n241_), .B(men_men_n240_), .Y(men_men_n242_));
  OR2        u0220(.A(i_8_), .B(i_7_), .Y(men_men_n243_));
  NO2        u0221(.A(men_men_n243_), .B(men_men_n86_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n54_), .B(i_1_), .Y(men_men_n245_));
  NA2        u0223(.A(men_men_n245_), .B(men_men_n244_), .Y(men_men_n246_));
  INV        u0224(.A(i_12_), .Y(men_men_n247_));
  NO2        u0225(.A(men_men_n45_), .B(men_men_n247_), .Y(men_men_n248_));
  NO3        u0226(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n249_));
  NA2        u0227(.A(i_2_), .B(i_1_), .Y(men_men_n250_));
  NO2        u0228(.A(men_men_n246_), .B(men_men_n242_), .Y(men_men_n251_));
  NO3        u0229(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n252_));
  NAi21      u0230(.An(i_4_), .B(i_3_), .Y(men_men_n253_));
  NO2        u0231(.A(men_men_n253_), .B(men_men_n75_), .Y(men_men_n254_));
  NO2        u0232(.A(i_0_), .B(i_6_), .Y(men_men_n255_));
  NOi41      u0233(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n256_));
  NA2        u0234(.A(men_men_n256_), .B(men_men_n255_), .Y(men_men_n257_));
  NO2        u0235(.A(men_men_n250_), .B(men_men_n188_), .Y(men_men_n258_));
  NAi21      u0236(.An(men_men_n257_), .B(men_men_n258_), .Y(men_men_n259_));
  INV        u0237(.A(men_men_n259_), .Y(men_men_n260_));
  AOI220     u0238(.A0(men_men_n260_), .A1(men_men_n40_), .B0(men_men_n251_), .B1(men_men_n214_), .Y(men_men_n261_));
  NO2        u0239(.A(i_11_), .B(men_men_n235_), .Y(men_men_n262_));
  NOi21      u0240(.An(i_1_), .B(i_6_), .Y(men_men_n263_));
  NAi21      u0241(.An(i_3_), .B(i_7_), .Y(men_men_n264_));
  NA2        u0242(.A(men_men_n247_), .B(i_9_), .Y(men_men_n265_));
  OR4        u0243(.A(men_men_n265_), .B(men_men_n264_), .C(men_men_n263_), .D(men_men_n191_), .Y(men_men_n266_));
  NO2        u0244(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n267_));
  NO2        u0245(.A(i_12_), .B(i_3_), .Y(men_men_n268_));
  NA2        u0246(.A(men_men_n73_), .B(i_5_), .Y(men_men_n269_));
  NA2        u0247(.A(i_3_), .B(i_9_), .Y(men_men_n270_));
  NAi21      u0248(.An(i_7_), .B(i_10_), .Y(men_men_n271_));
  NO2        u0249(.A(men_men_n271_), .B(men_men_n270_), .Y(men_men_n272_));
  NA3        u0250(.A(men_men_n272_), .B(men_men_n269_), .C(men_men_n64_), .Y(men_men_n273_));
  NA2        u0251(.A(men_men_n273_), .B(men_men_n266_), .Y(men_men_n274_));
  NA3        u0252(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n275_));
  INV        u0253(.A(men_men_n146_), .Y(men_men_n276_));
  NA2        u0254(.A(men_men_n247_), .B(i_13_), .Y(men_men_n277_));
  NO2        u0255(.A(men_men_n277_), .B(men_men_n75_), .Y(men_men_n278_));
  AOI220     u0256(.A0(men_men_n278_), .A1(men_men_n276_), .B0(men_men_n274_), .B1(men_men_n262_), .Y(men_men_n279_));
  NO2        u0257(.A(men_men_n243_), .B(men_men_n37_), .Y(men_men_n280_));
  NA2        u0258(.A(i_12_), .B(i_6_), .Y(men_men_n281_));
  OR2        u0259(.A(i_13_), .B(i_9_), .Y(men_men_n282_));
  NO3        u0260(.A(men_men_n282_), .B(men_men_n281_), .C(men_men_n49_), .Y(men_men_n283_));
  NO2        u0261(.A(men_men_n253_), .B(i_2_), .Y(men_men_n284_));
  NA3        u0262(.A(men_men_n284_), .B(men_men_n283_), .C(men_men_n45_), .Y(men_men_n285_));
  NA2        u0263(.A(men_men_n262_), .B(i_9_), .Y(men_men_n286_));
  NA3        u0264(.A(men_men_n269_), .B(men_men_n161_), .C(men_men_n64_), .Y(men_men_n287_));
  OAI210     u0265(.A0(men_men_n287_), .A1(men_men_n286_), .B0(men_men_n285_), .Y(men_men_n288_));
  NA2        u0266(.A(men_men_n158_), .B(men_men_n63_), .Y(men_men_n289_));
  NO3        u0267(.A(i_11_), .B(men_men_n235_), .C(men_men_n25_), .Y(men_men_n290_));
  NO2        u0268(.A(men_men_n264_), .B(i_8_), .Y(men_men_n291_));
  NO2        u0269(.A(i_6_), .B(men_men_n49_), .Y(men_men_n292_));
  NA3        u0270(.A(men_men_n292_), .B(men_men_n291_), .C(men_men_n290_), .Y(men_men_n293_));
  NO3        u0271(.A(men_men_n26_), .B(men_men_n86_), .C(i_5_), .Y(men_men_n294_));
  NA3        u0272(.A(men_men_n294_), .B(men_men_n280_), .C(men_men_n236_), .Y(men_men_n295_));
  AOI210     u0273(.A0(men_men_n295_), .A1(men_men_n293_), .B0(men_men_n289_), .Y(men_men_n296_));
  AOI210     u0274(.A0(men_men_n288_), .A1(men_men_n280_), .B0(men_men_n296_), .Y(men_men_n297_));
  NA4        u0275(.A(men_men_n297_), .B(men_men_n279_), .C(men_men_n261_), .D(men_men_n239_), .Y(men_men_n298_));
  NO3        u0276(.A(i_12_), .B(men_men_n235_), .C(men_men_n37_), .Y(men_men_n299_));
  INV        u0277(.A(men_men_n299_), .Y(men_men_n300_));
  NA2        u0278(.A(i_8_), .B(men_men_n104_), .Y(men_men_n301_));
  NOi21      u0279(.An(men_men_n167_), .B(men_men_n86_), .Y(men_men_n302_));
  NO3        u0280(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n303_));
  AOI220     u0281(.A0(men_men_n303_), .A1(men_men_n202_), .B0(men_men_n302_), .B1(men_men_n245_), .Y(men_men_n304_));
  NO2        u0282(.A(men_men_n304_), .B(men_men_n301_), .Y(men_men_n305_));
  NO3        u0283(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n306_));
  NO2        u0284(.A(men_men_n250_), .B(i_0_), .Y(men_men_n307_));
  AOI220     u0285(.A0(men_men_n307_), .A1(men_men_n200_), .B0(men_men_n306_), .B1(men_men_n145_), .Y(men_men_n308_));
  NA2        u0286(.A(men_men_n292_), .B(men_men_n26_), .Y(men_men_n309_));
  NO2        u0287(.A(men_men_n309_), .B(men_men_n308_), .Y(men_men_n310_));
  NA2        u0288(.A(i_0_), .B(i_1_), .Y(men_men_n311_));
  NO2        u0289(.A(men_men_n311_), .B(i_2_), .Y(men_men_n312_));
  NO2        u0290(.A(men_men_n59_), .B(i_6_), .Y(men_men_n313_));
  NA3        u0291(.A(men_men_n313_), .B(men_men_n312_), .C(men_men_n167_), .Y(men_men_n314_));
  OAI210     u0292(.A0(men_men_n169_), .A1(men_men_n146_), .B0(men_men_n314_), .Y(men_men_n315_));
  NO3        u0293(.A(men_men_n315_), .B(men_men_n310_), .C(men_men_n305_), .Y(men_men_n316_));
  NO2        u0294(.A(i_3_), .B(i_10_), .Y(men_men_n317_));
  NA3        u0295(.A(men_men_n317_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n318_));
  NO2        u0296(.A(i_2_), .B(men_men_n104_), .Y(men_men_n319_));
  NA2        u0297(.A(i_1_), .B(men_men_n36_), .Y(men_men_n320_));
  NO2        u0298(.A(men_men_n320_), .B(i_8_), .Y(men_men_n321_));
  NOi21      u0299(.An(men_men_n227_), .B(men_men_n106_), .Y(men_men_n322_));
  NA3        u0300(.A(men_men_n322_), .B(men_men_n321_), .C(men_men_n319_), .Y(men_men_n323_));
  AN2        u0301(.A(i_3_), .B(i_10_), .Y(men_men_n324_));
  NA4        u0302(.A(men_men_n324_), .B(men_men_n204_), .C(men_men_n181_), .D(men_men_n179_), .Y(men_men_n325_));
  NO2        u0303(.A(i_5_), .B(men_men_n37_), .Y(men_men_n326_));
  NO2        u0304(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n327_));
  OR2        u0305(.A(men_men_n323_), .B(men_men_n318_), .Y(men_men_n328_));
  OAI220     u0306(.A0(men_men_n328_), .A1(i_6_), .B0(men_men_n316_), .B1(men_men_n300_), .Y(men_men_n329_));
  NO4        u0307(.A(men_men_n329_), .B(men_men_n298_), .C(men_men_n223_), .D(men_men_n172_), .Y(men_men_n330_));
  NO3        u0308(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n331_));
  NO2        u0309(.A(men_men_n59_), .B(men_men_n86_), .Y(men_men_n332_));
  NA2        u0310(.A(men_men_n307_), .B(men_men_n332_), .Y(men_men_n333_));
  NO3        u0311(.A(i_6_), .B(men_men_n199_), .C(i_7_), .Y(men_men_n334_));
  NA2        u0312(.A(men_men_n334_), .B(men_men_n204_), .Y(men_men_n335_));
  AOI210     u0313(.A0(men_men_n335_), .A1(men_men_n333_), .B0(men_men_n174_), .Y(men_men_n336_));
  NO2        u0314(.A(i_2_), .B(i_3_), .Y(men_men_n337_));
  OR2        u0315(.A(i_0_), .B(i_5_), .Y(men_men_n338_));
  NA2        u0316(.A(men_men_n227_), .B(men_men_n338_), .Y(men_men_n339_));
  NA4        u0317(.A(men_men_n339_), .B(men_men_n244_), .C(men_men_n337_), .D(i_1_), .Y(men_men_n340_));
  NA3        u0318(.A(men_men_n307_), .B(men_men_n302_), .C(men_men_n116_), .Y(men_men_n341_));
  NAi21      u0319(.An(i_8_), .B(i_7_), .Y(men_men_n342_));
  NO2        u0320(.A(men_men_n342_), .B(i_6_), .Y(men_men_n343_));
  NO2        u0321(.A(men_men_n161_), .B(men_men_n47_), .Y(men_men_n344_));
  NA3        u0322(.A(men_men_n344_), .B(men_men_n343_), .C(men_men_n167_), .Y(men_men_n345_));
  NA3        u0323(.A(men_men_n345_), .B(men_men_n341_), .C(men_men_n340_), .Y(men_men_n346_));
  OAI210     u0324(.A0(men_men_n346_), .A1(men_men_n336_), .B0(i_4_), .Y(men_men_n347_));
  NO2        u0325(.A(i_12_), .B(i_10_), .Y(men_men_n348_));
  NOi21      u0326(.An(i_5_), .B(i_0_), .Y(men_men_n349_));
  NO3        u0327(.A(men_men_n320_), .B(men_men_n349_), .C(men_men_n131_), .Y(men_men_n350_));
  NA4        u0328(.A(men_men_n84_), .B(men_men_n36_), .C(men_men_n86_), .D(i_8_), .Y(men_men_n351_));
  NA2        u0329(.A(men_men_n350_), .B(men_men_n348_), .Y(men_men_n352_));
  NO2        u0330(.A(i_6_), .B(i_8_), .Y(men_men_n353_));
  NOi21      u0331(.An(i_0_), .B(i_2_), .Y(men_men_n354_));
  AN2        u0332(.A(men_men_n354_), .B(men_men_n353_), .Y(men_men_n355_));
  NO2        u0333(.A(i_1_), .B(i_7_), .Y(men_men_n356_));
  AO220      u0334(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n343_), .B1(men_men_n245_), .Y(men_men_n357_));
  NA3        u0335(.A(men_men_n357_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n358_));
  NA3        u0336(.A(men_men_n358_), .B(men_men_n352_), .C(men_men_n347_), .Y(men_men_n359_));
  NO3        u0337(.A(men_men_n243_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n360_));
  NO3        u0338(.A(men_men_n342_), .B(i_2_), .C(i_1_), .Y(men_men_n361_));
  OAI210     u0339(.A0(men_men_n361_), .A1(men_men_n360_), .B0(i_6_), .Y(men_men_n362_));
  NA3        u0340(.A(men_men_n263_), .B(men_men_n319_), .C(men_men_n199_), .Y(men_men_n363_));
  AOI210     u0341(.A0(men_men_n363_), .A1(men_men_n362_), .B0(men_men_n339_), .Y(men_men_n364_));
  NOi21      u0342(.An(men_men_n157_), .B(men_men_n107_), .Y(men_men_n365_));
  NA2        u0343(.A(men_men_n364_), .B(i_3_), .Y(men_men_n366_));
  INV        u0344(.A(men_men_n84_), .Y(men_men_n367_));
  NO2        u0345(.A(men_men_n311_), .B(men_men_n81_), .Y(men_men_n368_));
  NA2        u0346(.A(men_men_n368_), .B(men_men_n135_), .Y(men_men_n369_));
  NO2        u0347(.A(men_men_n95_), .B(men_men_n199_), .Y(men_men_n370_));
  NA3        u0348(.A(men_men_n322_), .B(men_men_n370_), .C(men_men_n63_), .Y(men_men_n371_));
  AOI210     u0349(.A0(men_men_n371_), .A1(men_men_n369_), .B0(men_men_n367_), .Y(men_men_n372_));
  NO2        u0350(.A(men_men_n199_), .B(i_9_), .Y(men_men_n373_));
  NA3        u0351(.A(men_men_n373_), .B(men_men_n212_), .C(men_men_n161_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n372_), .B(men_men_n310_), .Y(men_men_n375_));
  AOI210     u0353(.A0(men_men_n375_), .A1(men_men_n366_), .B0(men_men_n166_), .Y(men_men_n376_));
  AOI210     u0354(.A0(men_men_n359_), .A1(men_men_n331_), .B0(men_men_n376_), .Y(men_men_n377_));
  NOi32      u0355(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n378_));
  INV        u0356(.A(men_men_n378_), .Y(men_men_n379_));
  NAi21      u0357(.An(i_0_), .B(i_6_), .Y(men_men_n380_));
  NAi21      u0358(.An(i_1_), .B(i_5_), .Y(men_men_n381_));
  NA2        u0359(.A(men_men_n381_), .B(men_men_n380_), .Y(men_men_n382_));
  NA2        u0360(.A(men_men_n382_), .B(men_men_n25_), .Y(men_men_n383_));
  OAI210     u0361(.A0(men_men_n383_), .A1(men_men_n163_), .B0(men_men_n257_), .Y(men_men_n384_));
  NAi41      u0362(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n385_));
  OAI220     u0363(.A0(men_men_n385_), .A1(men_men_n381_), .B0(men_men_n230_), .B1(men_men_n163_), .Y(men_men_n386_));
  AOI210     u0364(.A0(men_men_n385_), .A1(men_men_n163_), .B0(men_men_n161_), .Y(men_men_n387_));
  NOi32      u0365(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n388_));
  OR2        u0366(.A(men_men_n387_), .B(men_men_n386_), .Y(men_men_n389_));
  NO2        u0367(.A(i_1_), .B(men_men_n104_), .Y(men_men_n390_));
  NAi21      u0368(.An(i_3_), .B(i_4_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n391_), .B(i_9_), .Y(men_men_n392_));
  AN2        u0370(.A(i_6_), .B(i_7_), .Y(men_men_n393_));
  OAI210     u0371(.A0(men_men_n393_), .A1(men_men_n390_), .B0(men_men_n392_), .Y(men_men_n394_));
  NA2        u0372(.A(i_2_), .B(i_7_), .Y(men_men_n395_));
  NO2        u0373(.A(men_men_n391_), .B(i_10_), .Y(men_men_n396_));
  NA3        u0374(.A(men_men_n396_), .B(men_men_n395_), .C(men_men_n255_), .Y(men_men_n397_));
  AOI210     u0375(.A0(men_men_n397_), .A1(men_men_n394_), .B0(men_men_n191_), .Y(men_men_n398_));
  AOI210     u0376(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n399_));
  OAI210     u0377(.A0(men_men_n399_), .A1(men_men_n194_), .B0(men_men_n396_), .Y(men_men_n400_));
  AOI220     u0378(.A0(men_men_n396_), .A1(men_men_n356_), .B0(men_men_n249_), .B1(men_men_n194_), .Y(men_men_n401_));
  AOI210     u0379(.A0(men_men_n401_), .A1(men_men_n400_), .B0(i_5_), .Y(men_men_n402_));
  NO4        u0380(.A(men_men_n402_), .B(men_men_n398_), .C(men_men_n389_), .D(men_men_n384_), .Y(men_men_n403_));
  NO2        u0381(.A(men_men_n403_), .B(men_men_n379_), .Y(men_men_n404_));
  NO2        u0382(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n405_));
  AN2        u0383(.A(i_12_), .B(i_5_), .Y(men_men_n406_));
  NO2        u0384(.A(i_4_), .B(men_men_n26_), .Y(men_men_n407_));
  NA2        u0385(.A(men_men_n407_), .B(men_men_n406_), .Y(men_men_n408_));
  NO2        u0386(.A(i_11_), .B(i_6_), .Y(men_men_n409_));
  NA3        u0387(.A(men_men_n409_), .B(men_men_n344_), .C(men_men_n235_), .Y(men_men_n410_));
  NO2        u0388(.A(men_men_n410_), .B(men_men_n408_), .Y(men_men_n411_));
  NO2        u0389(.A(men_men_n253_), .B(i_5_), .Y(men_men_n412_));
  NO2        u0390(.A(i_5_), .B(i_10_), .Y(men_men_n413_));
  AOI220     u0391(.A0(men_men_n413_), .A1(men_men_n284_), .B0(men_men_n412_), .B1(men_men_n204_), .Y(men_men_n414_));
  NA2        u0392(.A(men_men_n147_), .B(men_men_n46_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n415_), .B(men_men_n414_), .Y(men_men_n416_));
  OAI210     u0394(.A0(men_men_n416_), .A1(men_men_n411_), .B0(men_men_n405_), .Y(men_men_n417_));
  NO2        u0395(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n418_));
  NO2        u0396(.A(men_men_n153_), .B(men_men_n86_), .Y(men_men_n419_));
  OAI210     u0397(.A0(men_men_n419_), .A1(men_men_n411_), .B0(men_men_n418_), .Y(men_men_n420_));
  NO3        u0398(.A(men_men_n86_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n421_));
  NO2        u0399(.A(i_11_), .B(i_12_), .Y(men_men_n422_));
  NA2        u0400(.A(men_men_n413_), .B(men_men_n247_), .Y(men_men_n423_));
  NA3        u0401(.A(men_men_n116_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n424_));
  OAI220     u0402(.A0(men_men_n424_), .A1(men_men_n230_), .B0(men_men_n423_), .B1(men_men_n351_), .Y(men_men_n425_));
  NAi21      u0403(.An(i_13_), .B(i_0_), .Y(men_men_n426_));
  NO2        u0404(.A(men_men_n426_), .B(men_men_n250_), .Y(men_men_n427_));
  NA2        u0405(.A(men_men_n425_), .B(men_men_n427_), .Y(men_men_n428_));
  NA3        u0406(.A(men_men_n428_), .B(men_men_n420_), .C(men_men_n417_), .Y(men_men_n429_));
  NA2        u0407(.A(men_men_n45_), .B(men_men_n235_), .Y(men_men_n430_));
  NO3        u0408(.A(i_1_), .B(i_12_), .C(men_men_n86_), .Y(men_men_n431_));
  NO2        u0409(.A(i_0_), .B(i_11_), .Y(men_men_n432_));
  INV        u0410(.A(i_5_), .Y(men_men_n433_));
  AN2        u0411(.A(i_1_), .B(i_6_), .Y(men_men_n434_));
  NOi21      u0412(.An(i_2_), .B(i_12_), .Y(men_men_n435_));
  NA2        u0413(.A(men_men_n435_), .B(men_men_n434_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n436_), .B(men_men_n433_), .Y(men_men_n437_));
  NA2        u0415(.A(men_men_n145_), .B(i_9_), .Y(men_men_n438_));
  NO2        u0416(.A(men_men_n438_), .B(i_4_), .Y(men_men_n439_));
  NA2        u0417(.A(men_men_n437_), .B(men_men_n439_), .Y(men_men_n440_));
  NAi21      u0418(.An(i_9_), .B(i_4_), .Y(men_men_n441_));
  OR2        u0419(.A(i_13_), .B(i_10_), .Y(men_men_n442_));
  NO3        u0420(.A(men_men_n442_), .B(men_men_n120_), .C(men_men_n441_), .Y(men_men_n443_));
  NO2        u0421(.A(men_men_n177_), .B(men_men_n126_), .Y(men_men_n444_));
  OR2        u0422(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n445_));
  NO2        u0423(.A(men_men_n104_), .B(men_men_n25_), .Y(men_men_n446_));
  NA2        u0424(.A(men_men_n299_), .B(men_men_n446_), .Y(men_men_n447_));
  NA2        u0425(.A(men_men_n292_), .B(men_men_n219_), .Y(men_men_n448_));
  OAI220     u0426(.A0(men_men_n448_), .A1(men_men_n445_), .B0(men_men_n447_), .B1(men_men_n365_), .Y(men_men_n449_));
  INV        u0427(.A(men_men_n449_), .Y(men_men_n450_));
  AOI210     u0428(.A0(men_men_n450_), .A1(men_men_n440_), .B0(men_men_n26_), .Y(men_men_n451_));
  NA2        u0429(.A(men_men_n341_), .B(men_men_n340_), .Y(men_men_n452_));
  AOI220     u0430(.A0(men_men_n313_), .A1(men_men_n303_), .B0(men_men_n307_), .B1(men_men_n332_), .Y(men_men_n453_));
  NO2        u0431(.A(men_men_n453_), .B(men_men_n174_), .Y(men_men_n454_));
  NO2        u0432(.A(men_men_n188_), .B(men_men_n86_), .Y(men_men_n455_));
  AOI220     u0433(.A0(men_men_n455_), .A1(men_men_n312_), .B0(men_men_n294_), .B1(men_men_n219_), .Y(men_men_n456_));
  NO2        u0434(.A(men_men_n456_), .B(men_men_n301_), .Y(men_men_n457_));
  NO3        u0435(.A(men_men_n457_), .B(men_men_n454_), .C(men_men_n452_), .Y(men_men_n458_));
  NA2        u0436(.A(men_men_n202_), .B(men_men_n99_), .Y(men_men_n459_));
  NA3        u0437(.A(men_men_n344_), .B(men_men_n167_), .C(men_men_n86_), .Y(men_men_n460_));
  AOI210     u0438(.A0(men_men_n460_), .A1(men_men_n459_), .B0(men_men_n342_), .Y(men_men_n461_));
  NA2        u0439(.A(men_men_n313_), .B(men_men_n245_), .Y(men_men_n462_));
  NO2        u0440(.A(men_men_n462_), .B(men_men_n188_), .Y(men_men_n463_));
  NO2        u0441(.A(i_3_), .B(men_men_n49_), .Y(men_men_n464_));
  NA3        u0442(.A(men_men_n356_), .B(men_men_n355_), .C(men_men_n464_), .Y(men_men_n465_));
  NA2        u0443(.A(men_men_n334_), .B(men_men_n339_), .Y(men_men_n466_));
  OAI210     u0444(.A0(men_men_n466_), .A1(men_men_n195_), .B0(men_men_n465_), .Y(men_men_n467_));
  NO3        u0445(.A(men_men_n467_), .B(men_men_n463_), .C(men_men_n461_), .Y(men_men_n468_));
  AOI210     u0446(.A0(men_men_n468_), .A1(men_men_n458_), .B0(men_men_n286_), .Y(men_men_n469_));
  NO4        u0447(.A(men_men_n469_), .B(men_men_n451_), .C(men_men_n429_), .D(men_men_n404_), .Y(men_men_n470_));
  NO2        u0448(.A(men_men_n63_), .B(i_4_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n73_), .B(i_13_), .Y(men_men_n472_));
  NA3        u0450(.A(men_men_n472_), .B(men_men_n471_), .C(i_2_), .Y(men_men_n473_));
  NO2        u0451(.A(i_10_), .B(i_9_), .Y(men_men_n474_));
  NAi21      u0452(.An(i_12_), .B(i_8_), .Y(men_men_n475_));
  NO2        u0453(.A(men_men_n475_), .B(i_3_), .Y(men_men_n476_));
  NA2        u0454(.A(men_men_n476_), .B(men_men_n474_), .Y(men_men_n477_));
  NO2        u0455(.A(men_men_n47_), .B(i_4_), .Y(men_men_n478_));
  NA2        u0456(.A(men_men_n478_), .B(men_men_n107_), .Y(men_men_n479_));
  OAI220     u0457(.A0(men_men_n479_), .A1(men_men_n211_), .B0(men_men_n477_), .B1(men_men_n473_), .Y(men_men_n480_));
  NA2        u0458(.A(men_men_n327_), .B(i_0_), .Y(men_men_n481_));
  NO3        u0459(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n281_), .B(men_men_n100_), .Y(men_men_n483_));
  NA2        u0461(.A(men_men_n483_), .B(men_men_n482_), .Y(men_men_n484_));
  NA2        u0462(.A(i_8_), .B(i_9_), .Y(men_men_n485_));
  AOI210     u0463(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n486_));
  OR2        u0464(.A(men_men_n486_), .B(men_men_n485_), .Y(men_men_n487_));
  NA2        u0465(.A(men_men_n299_), .B(men_men_n212_), .Y(men_men_n488_));
  OAI220     u0466(.A0(men_men_n488_), .A1(men_men_n487_), .B0(men_men_n484_), .B1(men_men_n481_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n262_), .B(men_men_n326_), .Y(men_men_n490_));
  NO3        u0468(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n491_));
  INV        u0469(.A(men_men_n491_), .Y(men_men_n492_));
  NA3        u0470(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n493_));
  NA4        u0471(.A(men_men_n148_), .B(men_men_n119_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n494_));
  OAI220     u0472(.A0(men_men_n494_), .A1(men_men_n493_), .B0(men_men_n492_), .B1(men_men_n490_), .Y(men_men_n495_));
  NO3        u0473(.A(men_men_n495_), .B(men_men_n489_), .C(men_men_n480_), .Y(men_men_n496_));
  NA2        u0474(.A(men_men_n312_), .B(men_men_n111_), .Y(men_men_n497_));
  OR2        u0475(.A(men_men_n497_), .B(men_men_n215_), .Y(men_men_n498_));
  OA210      u0476(.A0(men_men_n374_), .A1(men_men_n104_), .B0(men_men_n314_), .Y(men_men_n499_));
  OA220      u0477(.A0(men_men_n499_), .A1(men_men_n166_), .B0(men_men_n498_), .B1(men_men_n242_), .Y(men_men_n500_));
  NA2        u0478(.A(men_men_n99_), .B(i_13_), .Y(men_men_n501_));
  NA2        u0479(.A(men_men_n455_), .B(men_men_n405_), .Y(men_men_n502_));
  NO2        u0480(.A(i_2_), .B(i_13_), .Y(men_men_n503_));
  NA3        u0481(.A(men_men_n503_), .B(men_men_n165_), .C(men_men_n102_), .Y(men_men_n504_));
  OAI220     u0482(.A0(men_men_n504_), .A1(men_men_n247_), .B0(men_men_n502_), .B1(men_men_n501_), .Y(men_men_n505_));
  NO3        u0483(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n506_));
  NO2        u0484(.A(i_6_), .B(i_7_), .Y(men_men_n507_));
  NA2        u0485(.A(men_men_n507_), .B(men_men_n506_), .Y(men_men_n508_));
  NO2        u0486(.A(i_11_), .B(i_1_), .Y(men_men_n509_));
  NO2        u0487(.A(men_men_n73_), .B(i_3_), .Y(men_men_n510_));
  OR2        u0488(.A(i_11_), .B(i_8_), .Y(men_men_n511_));
  NOi21      u0489(.An(i_2_), .B(i_7_), .Y(men_men_n512_));
  NAi31      u0490(.An(men_men_n511_), .B(men_men_n512_), .C(men_men_n510_), .Y(men_men_n513_));
  NO2        u0491(.A(men_men_n442_), .B(i_6_), .Y(men_men_n514_));
  NA3        u0492(.A(men_men_n514_), .B(men_men_n471_), .C(men_men_n75_), .Y(men_men_n515_));
  NO2        u0493(.A(men_men_n515_), .B(men_men_n513_), .Y(men_men_n516_));
  NO2        u0494(.A(i_3_), .B(men_men_n199_), .Y(men_men_n517_));
  NO2        u0495(.A(i_6_), .B(i_10_), .Y(men_men_n518_));
  NA4        u0496(.A(men_men_n518_), .B(men_men_n331_), .C(men_men_n517_), .D(men_men_n247_), .Y(men_men_n519_));
  NO2        u0497(.A(men_men_n519_), .B(men_men_n159_), .Y(men_men_n520_));
  NA3        u0498(.A(men_men_n256_), .B(men_men_n176_), .C(men_men_n135_), .Y(men_men_n521_));
  NA2        u0499(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n522_));
  NO2        u0500(.A(men_men_n161_), .B(i_3_), .Y(men_men_n523_));
  NAi31      u0501(.An(men_men_n522_), .B(men_men_n523_), .C(men_men_n236_), .Y(men_men_n524_));
  NA3        u0502(.A(men_men_n418_), .B(men_men_n184_), .C(men_men_n152_), .Y(men_men_n525_));
  NA3        u0503(.A(men_men_n525_), .B(men_men_n524_), .C(men_men_n521_), .Y(men_men_n526_));
  NO4        u0504(.A(men_men_n526_), .B(men_men_n520_), .C(men_men_n516_), .D(men_men_n505_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n482_), .B(men_men_n406_), .Y(men_men_n528_));
  NA2        u0506(.A(men_men_n491_), .B(men_men_n413_), .Y(men_men_n529_));
  NO2        u0507(.A(men_men_n529_), .B(men_men_n234_), .Y(men_men_n530_));
  NAi21      u0508(.An(men_men_n225_), .B(men_men_n422_), .Y(men_men_n531_));
  NA2        u0509(.A(men_men_n356_), .B(men_men_n227_), .Y(men_men_n532_));
  NO2        u0510(.A(men_men_n26_), .B(i_5_), .Y(men_men_n533_));
  NO2        u0511(.A(i_0_), .B(men_men_n86_), .Y(men_men_n534_));
  NA3        u0512(.A(men_men_n534_), .B(men_men_n533_), .C(men_men_n145_), .Y(men_men_n535_));
  OR3        u0513(.A(men_men_n320_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n536_));
  OAI220     u0514(.A0(men_men_n536_), .A1(men_men_n535_), .B0(men_men_n532_), .B1(men_men_n531_), .Y(men_men_n537_));
  NA2        u0515(.A(men_men_n27_), .B(i_10_), .Y(men_men_n538_));
  NO2        u0516(.A(men_men_n538_), .B(men_men_n501_), .Y(men_men_n539_));
  NA4        u0517(.A(men_men_n324_), .B(men_men_n233_), .C(men_men_n73_), .D(men_men_n247_), .Y(men_men_n540_));
  NO2        u0518(.A(men_men_n540_), .B(men_men_n508_), .Y(men_men_n541_));
  NO4        u0519(.A(men_men_n541_), .B(men_men_n539_), .C(men_men_n537_), .D(men_men_n530_), .Y(men_men_n542_));
  NA4        u0520(.A(men_men_n542_), .B(men_men_n527_), .C(men_men_n500_), .D(men_men_n496_), .Y(men_men_n543_));
  NA3        u0521(.A(men_men_n324_), .B(men_men_n181_), .C(men_men_n179_), .Y(men_men_n544_));
  OAI210     u0522(.A0(men_men_n318_), .A1(men_men_n186_), .B0(men_men_n544_), .Y(men_men_n545_));
  AN2        u0523(.A(men_men_n303_), .B(men_men_n244_), .Y(men_men_n546_));
  NA2        u0524(.A(men_men_n546_), .B(men_men_n545_), .Y(men_men_n547_));
  NA2        u0525(.A(men_men_n125_), .B(men_men_n115_), .Y(men_men_n548_));
  AO220      u0526(.A0(men_men_n548_), .A1(men_men_n482_), .B0(men_men_n443_), .B1(i_6_), .Y(men_men_n549_));
  NA2        u0527(.A(men_men_n331_), .B(men_men_n168_), .Y(men_men_n550_));
  OAI210     u0528(.A0(men_men_n550_), .A1(men_men_n242_), .B0(men_men_n325_), .Y(men_men_n551_));
  AOI220     u0529(.A0(men_men_n551_), .A1(men_men_n343_), .B0(men_men_n549_), .B1(men_men_n327_), .Y(men_men_n552_));
  NA2        u0530(.A(men_men_n406_), .B(men_men_n235_), .Y(men_men_n553_));
  NA2        u0531(.A(men_men_n378_), .B(men_men_n73_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n393_), .B(men_men_n388_), .Y(men_men_n555_));
  AO210      u0533(.A0(men_men_n554_), .A1(men_men_n553_), .B0(men_men_n555_), .Y(men_men_n556_));
  NO2        u0534(.A(men_men_n36_), .B(i_8_), .Y(men_men_n557_));
  AOI210     u0535(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n443_), .Y(men_men_n558_));
  NA2        u0536(.A(men_men_n558_), .B(men_men_n556_), .Y(men_men_n559_));
  INV        u0537(.A(men_men_n559_), .Y(men_men_n560_));
  NA2        u0538(.A(men_men_n269_), .B(men_men_n64_), .Y(men_men_n561_));
  OAI210     u0539(.A0(i_8_), .A1(men_men_n561_), .B0(men_men_n137_), .Y(men_men_n562_));
  NO2        u0540(.A(i_7_), .B(men_men_n205_), .Y(men_men_n563_));
  OR2        u0541(.A(men_men_n188_), .B(i_4_), .Y(men_men_n564_));
  NO2        u0542(.A(men_men_n564_), .B(men_men_n86_), .Y(men_men_n565_));
  AOI220     u0543(.A0(men_men_n565_), .A1(men_men_n563_), .B0(men_men_n562_), .B1(men_men_n444_), .Y(men_men_n566_));
  NA4        u0544(.A(men_men_n566_), .B(men_men_n560_), .C(men_men_n552_), .D(men_men_n547_), .Y(men_men_n567_));
  NA2        u0545(.A(men_men_n412_), .B(men_men_n312_), .Y(men_men_n568_));
  OAI210     u0546(.A0(men_men_n408_), .A1(men_men_n173_), .B0(men_men_n568_), .Y(men_men_n569_));
  NO2        u0547(.A(i_12_), .B(men_men_n199_), .Y(men_men_n570_));
  NA2        u0548(.A(men_men_n570_), .B(men_men_n235_), .Y(men_men_n571_));
  NO3        u0549(.A(men_men_n1116_), .B(men_men_n571_), .C(men_men_n497_), .Y(men_men_n572_));
  NOi31      u0550(.An(men_men_n334_), .B(men_men_n442_), .C(men_men_n38_), .Y(men_men_n573_));
  OAI210     u0551(.A0(men_men_n573_), .A1(men_men_n572_), .B0(men_men_n569_), .Y(men_men_n574_));
  NO2        u0552(.A(i_8_), .B(i_7_), .Y(men_men_n575_));
  OAI210     u0553(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n576_));
  NA2        u0554(.A(men_men_n576_), .B(men_men_n233_), .Y(men_men_n577_));
  AOI220     u0555(.A0(men_men_n344_), .A1(men_men_n40_), .B0(men_men_n245_), .B1(men_men_n214_), .Y(men_men_n578_));
  OAI220     u0556(.A0(men_men_n578_), .A1(men_men_n564_), .B0(men_men_n577_), .B1(men_men_n253_), .Y(men_men_n579_));
  NA2        u0557(.A(men_men_n45_), .B(i_10_), .Y(men_men_n580_));
  NO2        u0558(.A(men_men_n580_), .B(i_6_), .Y(men_men_n581_));
  NA3        u0559(.A(men_men_n581_), .B(men_men_n579_), .C(men_men_n575_), .Y(men_men_n582_));
  AOI220     u0560(.A0(men_men_n455_), .A1(men_men_n344_), .B0(men_men_n258_), .B1(men_men_n255_), .Y(men_men_n583_));
  OAI220     u0561(.A0(men_men_n583_), .A1(men_men_n277_), .B0(men_men_n501_), .B1(men_men_n136_), .Y(men_men_n584_));
  NA2        u0562(.A(men_men_n584_), .B(men_men_n280_), .Y(men_men_n585_));
  NOi31      u0563(.An(men_men_n307_), .B(men_men_n318_), .C(men_men_n186_), .Y(men_men_n586_));
  NA3        u0564(.A(men_men_n324_), .B(men_men_n179_), .C(men_men_n99_), .Y(men_men_n587_));
  NO2        u0565(.A(men_men_n231_), .B(men_men_n45_), .Y(men_men_n588_));
  NO2        u0566(.A(men_men_n161_), .B(i_5_), .Y(men_men_n589_));
  NA3        u0567(.A(men_men_n589_), .B(men_men_n430_), .C(men_men_n337_), .Y(men_men_n590_));
  OAI210     u0568(.A0(men_men_n590_), .A1(men_men_n588_), .B0(men_men_n587_), .Y(men_men_n591_));
  OAI210     u0569(.A0(men_men_n591_), .A1(men_men_n586_), .B0(men_men_n491_), .Y(men_men_n592_));
  NA4        u0570(.A(men_men_n592_), .B(men_men_n585_), .C(men_men_n582_), .D(men_men_n574_), .Y(men_men_n593_));
  NA3        u0571(.A(men_men_n227_), .B(men_men_n71_), .C(men_men_n45_), .Y(men_men_n594_));
  NA2        u0572(.A(men_men_n299_), .B(men_men_n84_), .Y(men_men_n595_));
  AOI210     u0573(.A0(men_men_n594_), .A1(men_men_n369_), .B0(men_men_n595_), .Y(men_men_n596_));
  NA2        u0574(.A(men_men_n313_), .B(men_men_n303_), .Y(men_men_n597_));
  NO2        u0575(.A(men_men_n597_), .B(men_men_n178_), .Y(men_men_n598_));
  NA2        u0576(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n599_));
  NA2        u0577(.A(men_men_n474_), .B(men_men_n231_), .Y(men_men_n600_));
  NO2        u0578(.A(men_men_n599_), .B(men_men_n600_), .Y(men_men_n601_));
  AOI210     u0579(.A0(i_6_), .A1(men_men_n47_), .B0(men_men_n390_), .Y(men_men_n602_));
  NA2        u0580(.A(i_0_), .B(men_men_n49_), .Y(men_men_n603_));
  NA3        u0581(.A(men_men_n570_), .B(men_men_n290_), .C(men_men_n603_), .Y(men_men_n604_));
  NO2        u0582(.A(men_men_n602_), .B(men_men_n604_), .Y(men_men_n605_));
  NO4        u0583(.A(men_men_n605_), .B(men_men_n601_), .C(men_men_n598_), .D(men_men_n596_), .Y(men_men_n606_));
  NO4        u0584(.A(men_men_n263_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n607_));
  NO3        u0585(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n608_));
  NO2        u0586(.A(men_men_n243_), .B(men_men_n36_), .Y(men_men_n609_));
  AN2        u0587(.A(men_men_n609_), .B(men_men_n608_), .Y(men_men_n610_));
  OA210      u0588(.A0(men_men_n610_), .A1(men_men_n607_), .B0(men_men_n378_), .Y(men_men_n611_));
  NO2        u0589(.A(men_men_n442_), .B(i_1_), .Y(men_men_n612_));
  NOi31      u0590(.An(men_men_n612_), .B(men_men_n483_), .C(men_men_n73_), .Y(men_men_n613_));
  AN4        u0591(.A(men_men_n613_), .B(men_men_n439_), .C(men_men_n533_), .D(i_2_), .Y(men_men_n614_));
  NO2        u0592(.A(men_men_n453_), .B(men_men_n182_), .Y(men_men_n615_));
  NO3        u0593(.A(men_men_n615_), .B(men_men_n614_), .C(men_men_n611_), .Y(men_men_n616_));
  NOi21      u0594(.An(i_10_), .B(i_6_), .Y(men_men_n617_));
  NO2        u0595(.A(men_men_n86_), .B(men_men_n25_), .Y(men_men_n618_));
  AOI220     u0596(.A0(men_men_n299_), .A1(men_men_n618_), .B0(men_men_n290_), .B1(men_men_n617_), .Y(men_men_n619_));
  NO2        u0597(.A(men_men_n619_), .B(men_men_n481_), .Y(men_men_n620_));
  NO2        u0598(.A(men_men_n118_), .B(men_men_n23_), .Y(men_men_n621_));
  NA2        u0599(.A(men_men_n334_), .B(men_men_n168_), .Y(men_men_n622_));
  AOI220     u0600(.A0(men_men_n622_), .A1(men_men_n462_), .B0(men_men_n189_), .B1(men_men_n187_), .Y(men_men_n623_));
  NO2        u0601(.A(men_men_n204_), .B(men_men_n37_), .Y(men_men_n624_));
  NOi31      u0602(.An(men_men_n149_), .B(men_men_n624_), .C(men_men_n351_), .Y(men_men_n625_));
  NO3        u0603(.A(men_men_n625_), .B(men_men_n623_), .C(men_men_n620_), .Y(men_men_n626_));
  NO2        u0604(.A(men_men_n554_), .B(men_men_n401_), .Y(men_men_n627_));
  INV        u0605(.A(men_men_n337_), .Y(men_men_n628_));
  NO2        u0606(.A(i_12_), .B(men_men_n86_), .Y(men_men_n629_));
  NA3        u0607(.A(men_men_n629_), .B(men_men_n290_), .C(men_men_n603_), .Y(men_men_n630_));
  NA3        u0608(.A(men_men_n409_), .B(men_men_n299_), .C(men_men_n227_), .Y(men_men_n631_));
  AOI210     u0609(.A0(men_men_n631_), .A1(men_men_n630_), .B0(men_men_n628_), .Y(men_men_n632_));
  NA2        u0610(.A(men_men_n179_), .B(i_0_), .Y(men_men_n633_));
  NO3        u0611(.A(men_men_n633_), .B(men_men_n362_), .C(men_men_n318_), .Y(men_men_n634_));
  OR2        u0612(.A(i_2_), .B(i_5_), .Y(men_men_n635_));
  OR2        u0613(.A(men_men_n635_), .B(men_men_n434_), .Y(men_men_n636_));
  NO2        u0614(.A(men_men_n636_), .B(men_men_n531_), .Y(men_men_n637_));
  NO4        u0615(.A(men_men_n637_), .B(men_men_n634_), .C(men_men_n632_), .D(men_men_n627_), .Y(men_men_n638_));
  NA4        u0616(.A(men_men_n638_), .B(men_men_n626_), .C(men_men_n616_), .D(men_men_n606_), .Y(men_men_n639_));
  NO4        u0617(.A(men_men_n639_), .B(men_men_n593_), .C(men_men_n567_), .D(men_men_n543_), .Y(men_men_n640_));
  NA4        u0618(.A(men_men_n640_), .B(men_men_n470_), .C(men_men_n377_), .D(men_men_n330_), .Y(men7));
  NO2        u0619(.A(men_men_n95_), .B(men_men_n55_), .Y(men_men_n642_));
  NO2        u0620(.A(men_men_n111_), .B(men_men_n92_), .Y(men_men_n643_));
  NA2        u0621(.A(men_men_n407_), .B(men_men_n643_), .Y(men_men_n644_));
  NA2        u0622(.A(men_men_n518_), .B(men_men_n84_), .Y(men_men_n645_));
  NA2        u0623(.A(i_11_), .B(men_men_n199_), .Y(men_men_n646_));
  INV        u0624(.A(men_men_n644_), .Y(men_men_n647_));
  NA3        u0625(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n648_));
  NO2        u0626(.A(men_men_n247_), .B(i_4_), .Y(men_men_n649_));
  NA2        u0627(.A(men_men_n649_), .B(i_8_), .Y(men_men_n650_));
  NO2        u0628(.A(men_men_n108_), .B(men_men_n648_), .Y(men_men_n651_));
  NA2        u0629(.A(i_2_), .B(men_men_n86_), .Y(men_men_n652_));
  OAI210     u0630(.A0(men_men_n89_), .A1(men_men_n209_), .B0(men_men_n210_), .Y(men_men_n653_));
  NO2        u0631(.A(i_7_), .B(men_men_n37_), .Y(men_men_n654_));
  NA2        u0632(.A(i_4_), .B(i_8_), .Y(men_men_n655_));
  AOI210     u0633(.A0(men_men_n655_), .A1(men_men_n324_), .B0(men_men_n654_), .Y(men_men_n656_));
  OAI220     u0634(.A0(men_men_n656_), .A1(men_men_n652_), .B0(men_men_n653_), .B1(i_13_), .Y(men_men_n657_));
  NO4        u0635(.A(men_men_n657_), .B(men_men_n651_), .C(men_men_n647_), .D(men_men_n642_), .Y(men_men_n658_));
  AOI210     u0636(.A0(men_men_n131_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n659_));
  AOI210     u0637(.A0(men_men_n659_), .A1(men_men_n247_), .B0(men_men_n165_), .Y(men_men_n660_));
  OR2        u0638(.A(i_6_), .B(i_10_), .Y(men_men_n661_));
  NO2        u0639(.A(men_men_n661_), .B(men_men_n23_), .Y(men_men_n662_));
  OR3        u0640(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n663_));
  NO3        u0641(.A(men_men_n663_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n664_));
  INV        u0642(.A(men_men_n206_), .Y(men_men_n665_));
  NO2        u0643(.A(men_men_n664_), .B(men_men_n662_), .Y(men_men_n666_));
  OA220      u0644(.A0(men_men_n666_), .A1(men_men_n628_), .B0(men_men_n660_), .B1(men_men_n282_), .Y(men_men_n667_));
  AOI210     u0645(.A0(men_men_n667_), .A1(men_men_n658_), .B0(men_men_n63_), .Y(men_men_n668_));
  NOi21      u0646(.An(i_11_), .B(i_7_), .Y(men_men_n669_));
  AO210      u0647(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n670_));
  NO2        u0648(.A(men_men_n670_), .B(men_men_n669_), .Y(men_men_n671_));
  NA2        u0649(.A(men_men_n671_), .B(men_men_n214_), .Y(men_men_n672_));
  NA3        u0650(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n673_));
  NAi31      u0651(.An(men_men_n673_), .B(men_men_n224_), .C(i_11_), .Y(men_men_n674_));
  AOI210     u0652(.A0(men_men_n674_), .A1(men_men_n672_), .B0(men_men_n63_), .Y(men_men_n675_));
  NA2        u0653(.A(men_men_n88_), .B(men_men_n63_), .Y(men_men_n676_));
  AO210      u0654(.A0(men_men_n676_), .A1(men_men_n401_), .B0(men_men_n41_), .Y(men_men_n677_));
  NO3        u0655(.A(men_men_n271_), .B(men_men_n216_), .C(men_men_n646_), .Y(men_men_n678_));
  OAI210     u0656(.A0(men_men_n678_), .A1(men_men_n236_), .B0(men_men_n63_), .Y(men_men_n679_));
  NA2        u0657(.A(men_men_n435_), .B(men_men_n31_), .Y(men_men_n680_));
  OR2        u0658(.A(men_men_n216_), .B(men_men_n111_), .Y(men_men_n681_));
  NA2        u0659(.A(men_men_n681_), .B(men_men_n680_), .Y(men_men_n682_));
  NO2        u0660(.A(men_men_n63_), .B(i_9_), .Y(men_men_n683_));
  NO2        u0661(.A(men_men_n683_), .B(i_4_), .Y(men_men_n684_));
  NA2        u0662(.A(men_men_n684_), .B(men_men_n682_), .Y(men_men_n685_));
  NO2        u0663(.A(i_1_), .B(i_12_), .Y(men_men_n686_));
  NA3        u0664(.A(men_men_n686_), .B(men_men_n113_), .C(men_men_n24_), .Y(men_men_n687_));
  NA4        u0665(.A(men_men_n687_), .B(men_men_n685_), .C(men_men_n679_), .D(men_men_n677_), .Y(men_men_n688_));
  OAI210     u0666(.A0(men_men_n688_), .A1(men_men_n675_), .B0(i_6_), .Y(men_men_n689_));
  NO2        u0667(.A(men_men_n247_), .B(men_men_n86_), .Y(men_men_n690_));
  NO2        u0668(.A(men_men_n690_), .B(i_11_), .Y(men_men_n691_));
  INV        u0669(.A(men_men_n484_), .Y(men_men_n692_));
  NO4        u0670(.A(men_men_n224_), .B(men_men_n131_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n693_));
  NA2        u0671(.A(men_men_n693_), .B(men_men_n683_), .Y(men_men_n694_));
  NA2        u0672(.A(men_men_n247_), .B(i_6_), .Y(men_men_n695_));
  NO3        u0673(.A(men_men_n661_), .B(men_men_n243_), .C(men_men_n23_), .Y(men_men_n696_));
  AOI210     u0674(.A0(i_1_), .A1(men_men_n272_), .B0(men_men_n696_), .Y(men_men_n697_));
  OAI210     u0675(.A0(men_men_n697_), .A1(men_men_n45_), .B0(men_men_n694_), .Y(men_men_n698_));
  NA3        u0676(.A(men_men_n575_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n699_));
  NA2        u0677(.A(men_men_n141_), .B(i_9_), .Y(men_men_n700_));
  NA3        u0678(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n701_));
  NO2        u0679(.A(men_men_n47_), .B(i_1_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n700_), .B(men_men_n1114_), .Y(men_men_n703_));
  NA3        u0681(.A(men_men_n683_), .B(men_men_n337_), .C(i_6_), .Y(men_men_n704_));
  NO2        u0682(.A(men_men_n704_), .B(men_men_n23_), .Y(men_men_n705_));
  AOI210     u0683(.A0(men_men_n509_), .A1(men_men_n446_), .B0(men_men_n252_), .Y(men_men_n706_));
  NO2        u0684(.A(men_men_n706_), .B(men_men_n652_), .Y(men_men_n707_));
  NO2        u0685(.A(i_11_), .B(men_men_n37_), .Y(men_men_n708_));
  NA2        u0686(.A(men_men_n708_), .B(men_men_n24_), .Y(men_men_n709_));
  OR3        u0687(.A(men_men_n707_), .B(men_men_n705_), .C(men_men_n703_), .Y(men_men_n710_));
  NO3        u0688(.A(men_men_n710_), .B(men_men_n698_), .C(men_men_n692_), .Y(men_men_n711_));
  NO2        u0689(.A(men_men_n247_), .B(men_men_n104_), .Y(men_men_n712_));
  NO2        u0690(.A(men_men_n712_), .B(men_men_n669_), .Y(men_men_n713_));
  NA2        u0691(.A(men_men_n713_), .B(i_1_), .Y(men_men_n714_));
  NO2        u0692(.A(men_men_n714_), .B(men_men_n663_), .Y(men_men_n715_));
  NO2        u0693(.A(men_men_n441_), .B(men_men_n86_), .Y(men_men_n716_));
  NA2        u0694(.A(men_men_n715_), .B(men_men_n47_), .Y(men_men_n717_));
  NO2        u0695(.A(men_men_n243_), .B(men_men_n45_), .Y(men_men_n718_));
  NO3        u0696(.A(men_men_n718_), .B(men_men_n327_), .C(men_men_n248_), .Y(men_men_n719_));
  NO2        u0697(.A(men_men_n120_), .B(men_men_n37_), .Y(men_men_n720_));
  NO2        u0698(.A(men_men_n720_), .B(i_6_), .Y(men_men_n721_));
  NO2        u0699(.A(men_men_n86_), .B(i_9_), .Y(men_men_n722_));
  NO2        u0700(.A(men_men_n722_), .B(men_men_n63_), .Y(men_men_n723_));
  NO2        u0701(.A(men_men_n723_), .B(men_men_n686_), .Y(men_men_n724_));
  NO4        u0702(.A(men_men_n724_), .B(men_men_n721_), .C(men_men_n719_), .D(i_4_), .Y(men_men_n725_));
  NA2        u0703(.A(i_1_), .B(i_3_), .Y(men_men_n726_));
  INV        u0704(.A(men_men_n725_), .Y(men_men_n727_));
  NA4        u0705(.A(men_men_n727_), .B(men_men_n717_), .C(men_men_n711_), .D(men_men_n689_), .Y(men_men_n728_));
  NO3        u0706(.A(men_men_n511_), .B(i_3_), .C(i_7_), .Y(men_men_n729_));
  NOi21      u0707(.An(men_men_n729_), .B(i_10_), .Y(men_men_n730_));
  OA210      u0708(.A0(men_men_n730_), .A1(men_men_n256_), .B0(men_men_n86_), .Y(men_men_n731_));
  NO3        u0709(.A(men_men_n512_), .B(men_men_n655_), .C(men_men_n86_), .Y(men_men_n732_));
  NA2        u0710(.A(men_men_n732_), .B(men_men_n25_), .Y(men_men_n733_));
  NA3        u0711(.A(men_men_n165_), .B(men_men_n84_), .C(men_men_n86_), .Y(men_men_n734_));
  NA2        u0712(.A(men_men_n734_), .B(men_men_n733_), .Y(men_men_n735_));
  OAI210     u0713(.A0(men_men_n735_), .A1(men_men_n731_), .B0(i_1_), .Y(men_men_n736_));
  AOI210     u0714(.A0(men_men_n281_), .A1(men_men_n100_), .B0(i_1_), .Y(men_men_n737_));
  NO2        u0715(.A(men_men_n391_), .B(i_2_), .Y(men_men_n738_));
  NA2        u0716(.A(men_men_n738_), .B(men_men_n737_), .Y(men_men_n739_));
  OAI210     u0717(.A0(men_men_n704_), .A1(men_men_n475_), .B0(men_men_n739_), .Y(men_men_n740_));
  INV        u0718(.A(men_men_n740_), .Y(men_men_n741_));
  AOI210     u0719(.A0(men_men_n741_), .A1(men_men_n736_), .B0(i_13_), .Y(men_men_n742_));
  OR2        u0720(.A(i_11_), .B(i_7_), .Y(men_men_n743_));
  NA3        u0721(.A(men_men_n743_), .B(men_men_n109_), .C(men_men_n141_), .Y(men_men_n744_));
  AOI220     u0722(.A0(men_men_n503_), .A1(men_men_n165_), .B0(men_men_n478_), .B1(men_men_n141_), .Y(men_men_n745_));
  OAI210     u0723(.A0(men_men_n745_), .A1(men_men_n45_), .B0(men_men_n744_), .Y(men_men_n746_));
  AOI210     u0724(.A0(men_men_n701_), .A1(men_men_n55_), .B0(i_12_), .Y(men_men_n747_));
  INV        u0725(.A(men_men_n747_), .Y(men_men_n748_));
  NO2        u0726(.A(men_men_n512_), .B(men_men_n24_), .Y(men_men_n749_));
  AOI220     u0727(.A0(men_men_n749_), .A1(men_men_n716_), .B0(men_men_n256_), .B1(men_men_n134_), .Y(men_men_n750_));
  OAI220     u0728(.A0(men_men_n750_), .A1(men_men_n41_), .B0(men_men_n748_), .B1(men_men_n95_), .Y(men_men_n751_));
  AOI210     u0729(.A0(men_men_n746_), .A1(men_men_n353_), .B0(men_men_n751_), .Y(men_men_n752_));
  NA2        u0730(.A(men_men_n409_), .B(men_men_n702_), .Y(men_men_n753_));
  NO2        u0731(.A(men_men_n753_), .B(men_men_n253_), .Y(men_men_n754_));
  AOI210     u0732(.A0(men_men_n475_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n755_));
  NOi31      u0733(.An(men_men_n755_), .B(men_men_n645_), .C(men_men_n45_), .Y(men_men_n756_));
  NA2        u0734(.A(men_men_n130_), .B(i_13_), .Y(men_men_n757_));
  NO2        u0735(.A(men_men_n701_), .B(men_men_n118_), .Y(men_men_n758_));
  INV        u0736(.A(men_men_n758_), .Y(men_men_n759_));
  OAI220     u0737(.A0(men_men_n759_), .A1(men_men_n71_), .B0(men_men_n757_), .B1(men_men_n737_), .Y(men_men_n760_));
  NO3        u0738(.A(men_men_n71_), .B(men_men_n32_), .C(men_men_n104_), .Y(men_men_n761_));
  NA2        u0739(.A(men_men_n26_), .B(men_men_n199_), .Y(men_men_n762_));
  AOI220     u0740(.A0(men_men_n409_), .A1(men_men_n702_), .B0(men_men_n94_), .B1(men_men_n105_), .Y(men_men_n763_));
  OAI220     u0741(.A0(men_men_n763_), .A1(men_men_n650_), .B0(men_men_n1115_), .B1(men_men_n665_), .Y(men_men_n764_));
  NO4        u0742(.A(men_men_n764_), .B(men_men_n760_), .C(men_men_n756_), .D(men_men_n754_), .Y(men_men_n765_));
  OR2        u0743(.A(i_11_), .B(i_6_), .Y(men_men_n766_));
  NA3        u0744(.A(men_men_n649_), .B(men_men_n762_), .C(i_7_), .Y(men_men_n767_));
  AOI210     u0745(.A0(men_men_n767_), .A1(men_men_n759_), .B0(men_men_n766_), .Y(men_men_n768_));
  NA3        u0746(.A(men_men_n435_), .B(men_men_n654_), .C(men_men_n100_), .Y(men_men_n769_));
  NA2        u0747(.A(men_men_n691_), .B(i_13_), .Y(men_men_n770_));
  NA2        u0748(.A(men_men_n105_), .B(men_men_n762_), .Y(men_men_n771_));
  NAi21      u0749(.An(i_11_), .B(i_12_), .Y(men_men_n772_));
  NOi41      u0750(.An(men_men_n114_), .B(men_men_n772_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n773_));
  NA2        u0751(.A(men_men_n773_), .B(men_men_n771_), .Y(men_men_n774_));
  NA3        u0752(.A(men_men_n774_), .B(men_men_n770_), .C(men_men_n769_), .Y(men_men_n775_));
  OAI210     u0753(.A0(men_men_n775_), .A1(men_men_n768_), .B0(men_men_n63_), .Y(men_men_n776_));
  NO2        u0754(.A(i_2_), .B(i_12_), .Y(men_men_n777_));
  NA2        u0755(.A(men_men_n390_), .B(men_men_n777_), .Y(men_men_n778_));
  NA2        u0756(.A(i_8_), .B(men_men_n25_), .Y(men_men_n779_));
  NO3        u0757(.A(men_men_n779_), .B(men_men_n407_), .C(men_men_n649_), .Y(men_men_n780_));
  OAI210     u0758(.A0(men_men_n780_), .A1(men_men_n392_), .B0(men_men_n390_), .Y(men_men_n781_));
  NO2        u0759(.A(men_men_n131_), .B(i_2_), .Y(men_men_n782_));
  NA2        u0760(.A(men_men_n782_), .B(men_men_n686_), .Y(men_men_n783_));
  NA3        u0761(.A(men_men_n783_), .B(men_men_n781_), .C(men_men_n778_), .Y(men_men_n784_));
  NA3        u0762(.A(men_men_n784_), .B(men_men_n46_), .C(men_men_n235_), .Y(men_men_n785_));
  NA4        u0763(.A(men_men_n785_), .B(men_men_n776_), .C(men_men_n765_), .D(men_men_n752_), .Y(men_men_n786_));
  OR4        u0764(.A(men_men_n786_), .B(men_men_n742_), .C(men_men_n728_), .D(men_men_n668_), .Y(men5));
  AOI210     u0765(.A0(men_men_n713_), .A1(men_men_n284_), .B0(men_men_n444_), .Y(men_men_n788_));
  AN2        u0766(.A(men_men_n24_), .B(i_10_), .Y(men_men_n789_));
  NA3        u0767(.A(men_men_n789_), .B(men_men_n777_), .C(men_men_n111_), .Y(men_men_n790_));
  NO2        u0768(.A(men_men_n650_), .B(i_11_), .Y(men_men_n791_));
  OAI210     u0769(.A0(men_men_n654_), .A1(men_men_n89_), .B0(men_men_n791_), .Y(men_men_n792_));
  NA3        u0770(.A(men_men_n792_), .B(men_men_n790_), .C(men_men_n788_), .Y(men_men_n793_));
  NO3        u0771(.A(i_11_), .B(men_men_n247_), .C(i_13_), .Y(men_men_n794_));
  NO2        u0772(.A(men_men_n127_), .B(men_men_n23_), .Y(men_men_n795_));
  NA2        u0773(.A(i_12_), .B(i_8_), .Y(men_men_n796_));
  OAI210     u0774(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n796_), .Y(men_men_n797_));
  INV        u0775(.A(men_men_n474_), .Y(men_men_n798_));
  AOI220     u0776(.A0(men_men_n337_), .A1(men_men_n621_), .B0(men_men_n797_), .B1(men_men_n795_), .Y(men_men_n799_));
  INV        u0777(.A(men_men_n799_), .Y(men_men_n800_));
  NO2        u0778(.A(men_men_n800_), .B(men_men_n793_), .Y(men_men_n801_));
  INV        u0779(.A(men_men_n176_), .Y(men_men_n802_));
  INV        u0780(.A(men_men_n256_), .Y(men_men_n803_));
  OAI210     u0781(.A0(men_men_n738_), .A1(men_men_n476_), .B0(men_men_n114_), .Y(men_men_n804_));
  AOI210     u0782(.A0(men_men_n804_), .A1(men_men_n803_), .B0(men_men_n802_), .Y(men_men_n805_));
  NO2        u0783(.A(men_men_n485_), .B(men_men_n26_), .Y(men_men_n806_));
  NO2        u0784(.A(men_men_n806_), .B(men_men_n446_), .Y(men_men_n807_));
  NA2        u0785(.A(men_men_n807_), .B(i_2_), .Y(men_men_n808_));
  INV        u0786(.A(men_men_n808_), .Y(men_men_n809_));
  AOI210     u0787(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n442_), .Y(men_men_n810_));
  AOI210     u0788(.A0(men_men_n810_), .A1(men_men_n809_), .B0(men_men_n805_), .Y(men_men_n811_));
  NO2        u0789(.A(men_men_n196_), .B(men_men_n128_), .Y(men_men_n812_));
  OAI210     u0790(.A0(men_men_n812_), .A1(men_men_n795_), .B0(i_2_), .Y(men_men_n813_));
  INV        u0791(.A(men_men_n177_), .Y(men_men_n814_));
  NO3        u0792(.A(men_men_n670_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n815_));
  AOI210     u0793(.A0(men_men_n814_), .A1(men_men_n89_), .B0(men_men_n815_), .Y(men_men_n816_));
  AOI210     u0794(.A0(men_men_n816_), .A1(men_men_n813_), .B0(men_men_n199_), .Y(men_men_n817_));
  OA210      u0795(.A0(men_men_n671_), .A1(men_men_n129_), .B0(i_13_), .Y(men_men_n818_));
  NA2        u0796(.A(men_men_n206_), .B(men_men_n209_), .Y(men_men_n819_));
  NA2        u0797(.A(men_men_n155_), .B(men_men_n646_), .Y(men_men_n820_));
  AOI210     u0798(.A0(men_men_n820_), .A1(men_men_n819_), .B0(men_men_n395_), .Y(men_men_n821_));
  AOI210     u0799(.A0(men_men_n216_), .A1(men_men_n151_), .B0(men_men_n557_), .Y(men_men_n822_));
  OAI210     u0800(.A0(men_men_n822_), .A1(men_men_n236_), .B0(men_men_n446_), .Y(men_men_n823_));
  NO2        u0801(.A(men_men_n105_), .B(men_men_n45_), .Y(men_men_n824_));
  INV        u0802(.A(men_men_n319_), .Y(men_men_n825_));
  NA4        u0803(.A(men_men_n825_), .B(men_men_n324_), .C(men_men_n127_), .D(men_men_n43_), .Y(men_men_n826_));
  OAI210     u0804(.A0(men_men_n826_), .A1(men_men_n824_), .B0(men_men_n823_), .Y(men_men_n827_));
  NO4        u0805(.A(men_men_n827_), .B(men_men_n821_), .C(men_men_n818_), .D(men_men_n817_), .Y(men_men_n828_));
  NA2        u0806(.A(men_men_n621_), .B(men_men_n28_), .Y(men_men_n829_));
  NA2        u0807(.A(men_men_n794_), .B(men_men_n291_), .Y(men_men_n830_));
  NA2        u0808(.A(men_men_n830_), .B(men_men_n829_), .Y(men_men_n831_));
  NO2        u0809(.A(men_men_n62_), .B(i_12_), .Y(men_men_n832_));
  NO2        u0810(.A(men_men_n832_), .B(men_men_n129_), .Y(men_men_n833_));
  NO2        u0811(.A(men_men_n833_), .B(men_men_n646_), .Y(men_men_n834_));
  AOI220     u0812(.A0(men_men_n834_), .A1(men_men_n36_), .B0(men_men_n831_), .B1(men_men_n47_), .Y(men_men_n835_));
  NA4        u0813(.A(men_men_n835_), .B(men_men_n828_), .C(men_men_n811_), .D(men_men_n801_), .Y(men6));
  NO3        u0814(.A(men_men_n267_), .B(men_men_n326_), .C(i_1_), .Y(men_men_n837_));
  NO2        u0815(.A(men_men_n191_), .B(men_men_n142_), .Y(men_men_n838_));
  OAI210     u0816(.A0(men_men_n838_), .A1(men_men_n837_), .B0(men_men_n782_), .Y(men_men_n839_));
  NO2        u0817(.A(men_men_n230_), .B(men_men_n522_), .Y(men_men_n840_));
  INV        u0818(.A(men_men_n349_), .Y(men_men_n841_));
  AO210      u0819(.A0(men_men_n841_), .A1(men_men_n839_), .B0(i_12_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n629_), .B(men_men_n63_), .Y(men_men_n843_));
  NA2        u0821(.A(men_men_n730_), .B(men_men_n71_), .Y(men_men_n844_));
  BUFFER     u0822(.A(men_men_n676_), .Y(men_men_n845_));
  NA3        u0823(.A(men_men_n845_), .B(men_men_n844_), .C(men_men_n843_), .Y(men_men_n846_));
  NA2        u0824(.A(men_men_n846_), .B(men_men_n73_), .Y(men_men_n847_));
  INV        u0825(.A(men_men_n348_), .Y(men_men_n848_));
  NA2        u0826(.A(men_men_n75_), .B(men_men_n134_), .Y(men_men_n849_));
  INV        u0827(.A(men_men_n127_), .Y(men_men_n850_));
  NA2        u0828(.A(men_men_n850_), .B(men_men_n47_), .Y(men_men_n851_));
  AOI210     u0829(.A0(men_men_n851_), .A1(men_men_n849_), .B0(men_men_n848_), .Y(men_men_n852_));
  NO3        u0830(.A(men_men_n263_), .B(men_men_n135_), .C(i_9_), .Y(men_men_n853_));
  NA2        u0831(.A(men_men_n853_), .B(men_men_n832_), .Y(men_men_n854_));
  AOI210     u0832(.A0(men_men_n854_), .A1(men_men_n555_), .B0(men_men_n191_), .Y(men_men_n855_));
  NO2        u0833(.A(men_men_n32_), .B(i_11_), .Y(men_men_n856_));
  NA3        u0834(.A(men_men_n856_), .B(men_men_n507_), .C(men_men_n413_), .Y(men_men_n857_));
  NAi32      u0835(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n858_));
  AOI210     u0836(.A0(men_men_n766_), .A1(men_men_n87_), .B0(men_men_n858_), .Y(men_men_n859_));
  OAI210     u0837(.A0(men_men_n729_), .A1(men_men_n609_), .B0(men_men_n608_), .Y(men_men_n860_));
  NAi31      u0838(.An(men_men_n859_), .B(men_men_n860_), .C(men_men_n857_), .Y(men_men_n861_));
  OR3        u0839(.A(men_men_n861_), .B(men_men_n855_), .C(men_men_n852_), .Y(men_men_n862_));
  NO2        u0840(.A(men_men_n743_), .B(i_2_), .Y(men_men_n863_));
  NA2        u0841(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n864_));
  OAI210     u0842(.A0(men_men_n864_), .A1(men_men_n434_), .B0(men_men_n383_), .Y(men_men_n865_));
  NA2        u0843(.A(men_men_n865_), .B(men_men_n863_), .Y(men_men_n866_));
  AO220      u0844(.A0(men_men_n382_), .A1(men_men_n373_), .B0(men_men_n421_), .B1(men_men_n646_), .Y(men_men_n867_));
  NA3        u0845(.A(men_men_n867_), .B(men_men_n268_), .C(i_7_), .Y(men_men_n868_));
  OR2        u0846(.A(men_men_n671_), .B(men_men_n476_), .Y(men_men_n869_));
  NA3        u0847(.A(men_men_n869_), .B(men_men_n150_), .C(men_men_n69_), .Y(men_men_n870_));
  AO210      u0848(.A0(men_men_n529_), .A1(men_men_n798_), .B0(men_men_n36_), .Y(men_men_n871_));
  NA4        u0849(.A(men_men_n871_), .B(men_men_n870_), .C(men_men_n868_), .D(men_men_n866_), .Y(men_men_n872_));
  OAI210     u0850(.A0(men_men_n690_), .A1(i_11_), .B0(men_men_n87_), .Y(men_men_n873_));
  AOI220     u0851(.A0(men_men_n873_), .A1(men_men_n608_), .B0(men_men_n840_), .B1(men_men_n1117_), .Y(men_men_n874_));
  NA3        u0852(.A(men_men_n395_), .B(men_men_n249_), .C(men_men_n150_), .Y(men_men_n875_));
  OAI210     u0853(.A0(men_men_n421_), .A1(men_men_n210_), .B0(men_men_n70_), .Y(men_men_n876_));
  NA4        u0854(.A(men_men_n876_), .B(men_men_n875_), .C(men_men_n874_), .D(men_men_n653_), .Y(men_men_n877_));
  NA3        u0855(.A(men_men_n88_), .B(men_men_n518_), .C(men_men_n227_), .Y(men_men_n878_));
  AOI210     u0856(.A0(men_men_n476_), .A1(men_men_n474_), .B0(men_men_n607_), .Y(men_men_n879_));
  NO2        u0857(.A(men_men_n661_), .B(men_men_n105_), .Y(men_men_n880_));
  OAI210     u0858(.A0(men_men_n880_), .A1(men_men_n115_), .B0(men_men_n432_), .Y(men_men_n881_));
  NA2        u0859(.A(men_men_n255_), .B(men_men_n47_), .Y(men_men_n882_));
  NA2        u0860(.A(men_men_n882_), .B(men_men_n636_), .Y(men_men_n883_));
  NA3        u0861(.A(men_men_n883_), .B(men_men_n348_), .C(i_7_), .Y(men_men_n884_));
  NA4        u0862(.A(men_men_n884_), .B(men_men_n881_), .C(men_men_n879_), .D(men_men_n878_), .Y(men_men_n885_));
  NO4        u0863(.A(men_men_n885_), .B(men_men_n877_), .C(men_men_n872_), .D(men_men_n862_), .Y(men_men_n886_));
  NA4        u0864(.A(men_men_n886_), .B(men_men_n847_), .C(men_men_n842_), .D(men_men_n403_), .Y(men3));
  NA2        u0865(.A(i_6_), .B(i_7_), .Y(men_men_n888_));
  NO2        u0866(.A(men_men_n888_), .B(i_0_), .Y(men_men_n889_));
  NO2        u0867(.A(i_11_), .B(men_men_n247_), .Y(men_men_n890_));
  OAI210     u0868(.A0(men_men_n889_), .A1(men_men_n307_), .B0(men_men_n890_), .Y(men_men_n891_));
  NO2        u0869(.A(men_men_n891_), .B(men_men_n199_), .Y(men_men_n892_));
  NO3        u0870(.A(men_men_n481_), .B(men_men_n92_), .C(men_men_n45_), .Y(men_men_n893_));
  OA210      u0871(.A0(men_men_n893_), .A1(men_men_n892_), .B0(men_men_n179_), .Y(men_men_n894_));
  NA3        u0872(.A(men_men_n875_), .B(men_men_n653_), .C(men_men_n394_), .Y(men_men_n895_));
  NA2        u0873(.A(men_men_n895_), .B(men_men_n40_), .Y(men_men_n896_));
  NOi21      u0874(.An(men_men_n99_), .B(men_men_n807_), .Y(men_men_n897_));
  NO3        u0875(.A(men_men_n681_), .B(men_men_n485_), .C(men_men_n134_), .Y(men_men_n898_));
  NA2        u0876(.A(men_men_n435_), .B(men_men_n46_), .Y(men_men_n899_));
  NO2        u0877(.A(men_men_n898_), .B(men_men_n897_), .Y(men_men_n900_));
  AOI210     u0878(.A0(men_men_n900_), .A1(men_men_n896_), .B0(men_men_n49_), .Y(men_men_n901_));
  NO4        u0879(.A(men_men_n399_), .B(men_men_n406_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n902_));
  NA2        u0880(.A(men_men_n191_), .B(men_men_n617_), .Y(men_men_n903_));
  NOi31      u0881(.An(men_men_n903_), .B(men_men_n902_), .C(men_men_n39_), .Y(men_men_n904_));
  NA2        u0882(.A(men_men_n755_), .B(men_men_n722_), .Y(men_men_n905_));
  NA2        u0883(.A(men_men_n354_), .B(men_men_n464_), .Y(men_men_n906_));
  OAI220     u0884(.A0(men_men_n906_), .A1(men_men_n905_), .B0(men_men_n904_), .B1(men_men_n63_), .Y(men_men_n907_));
  NOi21      u0885(.An(i_5_), .B(i_9_), .Y(men_men_n908_));
  NA2        u0886(.A(men_men_n908_), .B(men_men_n472_), .Y(men_men_n909_));
  AOI210     u0887(.A0(men_men_n281_), .A1(men_men_n509_), .B0(men_men_n732_), .Y(men_men_n910_));
  NO3        u0888(.A(men_men_n438_), .B(men_men_n281_), .C(men_men_n73_), .Y(men_men_n911_));
  NO2        u0889(.A(men_men_n180_), .B(men_men_n151_), .Y(men_men_n912_));
  AOI210     u0890(.A0(men_men_n912_), .A1(men_men_n255_), .B0(men_men_n911_), .Y(men_men_n913_));
  OAI220     u0891(.A0(men_men_n913_), .A1(men_men_n186_), .B0(men_men_n910_), .B1(men_men_n909_), .Y(men_men_n914_));
  NO4        u0892(.A(men_men_n914_), .B(men_men_n907_), .C(men_men_n901_), .D(men_men_n894_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n191_), .B(men_men_n24_), .Y(men_men_n916_));
  NO2        u0894(.A(men_men_n720_), .B(men_men_n643_), .Y(men_men_n917_));
  NO2        u0895(.A(men_men_n917_), .B(men_men_n916_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n331_), .B(men_men_n132_), .Y(men_men_n919_));
  NAi21      u0897(.An(men_men_n166_), .B(men_men_n464_), .Y(men_men_n920_));
  OAI220     u0898(.A0(men_men_n920_), .A1(men_men_n882_), .B0(men_men_n919_), .B1(men_men_n423_), .Y(men_men_n921_));
  NO2        u0899(.A(men_men_n921_), .B(men_men_n918_), .Y(men_men_n922_));
  NO2        u0900(.A(men_men_n413_), .B(men_men_n311_), .Y(men_men_n923_));
  NA2        u0901(.A(men_men_n923_), .B(men_men_n758_), .Y(men_men_n924_));
  NA2        u0902(.A(men_men_n618_), .B(i_0_), .Y(men_men_n925_));
  NO3        u0903(.A(men_men_n925_), .B(men_men_n408_), .C(men_men_n89_), .Y(men_men_n926_));
  NO4        u0904(.A(men_men_n635_), .B(men_men_n224_), .C(men_men_n442_), .D(men_men_n434_), .Y(men_men_n927_));
  AOI210     u0905(.A0(men_men_n927_), .A1(i_11_), .B0(men_men_n926_), .Y(men_men_n928_));
  INV        u0906(.A(men_men_n507_), .Y(men_men_n929_));
  AN2        u0907(.A(men_men_n99_), .B(men_men_n254_), .Y(men_men_n930_));
  NA2        u0908(.A(men_men_n794_), .B(men_men_n349_), .Y(men_men_n931_));
  AOI210     u0909(.A0(men_men_n518_), .A1(men_men_n89_), .B0(men_men_n58_), .Y(men_men_n932_));
  OAI220     u0910(.A0(men_men_n932_), .A1(men_men_n931_), .B0(men_men_n709_), .B1(men_men_n577_), .Y(men_men_n933_));
  NO2        u0911(.A(men_men_n265_), .B(men_men_n157_), .Y(men_men_n934_));
  NA2        u0912(.A(i_0_), .B(i_10_), .Y(men_men_n935_));
  AN2        u0913(.A(men_men_n934_), .B(i_6_), .Y(men_men_n936_));
  AOI220     u0914(.A0(men_men_n354_), .A1(men_men_n101_), .B0(men_men_n191_), .B1(men_men_n84_), .Y(men_men_n937_));
  NA2        u0915(.A(men_men_n612_), .B(i_4_), .Y(men_men_n938_));
  NA2        u0916(.A(men_men_n194_), .B(men_men_n209_), .Y(men_men_n939_));
  OAI220     u0917(.A0(men_men_n939_), .A1(men_men_n931_), .B0(men_men_n938_), .B1(men_men_n937_), .Y(men_men_n940_));
  NO4        u0918(.A(men_men_n940_), .B(men_men_n936_), .C(men_men_n933_), .D(men_men_n930_), .Y(men_men_n941_));
  NA4        u0919(.A(men_men_n941_), .B(men_men_n928_), .C(men_men_n924_), .D(men_men_n922_), .Y(men_men_n942_));
  NA2        u0920(.A(i_11_), .B(i_9_), .Y(men_men_n943_));
  NO2        u0921(.A(men_men_n49_), .B(i_7_), .Y(men_men_n944_));
  NA2        u0922(.A(men_men_n418_), .B(men_men_n184_), .Y(men_men_n945_));
  NA3        u0923(.A(men_men_n945_), .B(men_men_n490_), .C(men_men_n164_), .Y(men_men_n946_));
  NO2        u0924(.A(men_men_n943_), .B(men_men_n73_), .Y(men_men_n947_));
  NO2        u0925(.A(men_men_n180_), .B(i_0_), .Y(men_men_n948_));
  INV        u0926(.A(men_men_n948_), .Y(men_men_n949_));
  NA2        u0927(.A(men_men_n507_), .B(men_men_n241_), .Y(men_men_n950_));
  AOI210     u0928(.A0(men_men_n393_), .A1(men_men_n42_), .B0(men_men_n431_), .Y(men_men_n951_));
  OAI220     u0929(.A0(men_men_n951_), .A1(men_men_n909_), .B0(men_men_n950_), .B1(men_men_n949_), .Y(men_men_n952_));
  NO2        u0930(.A(men_men_n952_), .B(men_men_n946_), .Y(men_men_n953_));
  NA2        u0931(.A(men_men_n708_), .B(men_men_n124_), .Y(men_men_n954_));
  NO2        u0932(.A(i_6_), .B(men_men_n954_), .Y(men_men_n955_));
  AOI210     u0933(.A0(men_men_n475_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n956_));
  NA2        u0934(.A(men_men_n176_), .B(men_men_n106_), .Y(men_men_n957_));
  NOi32      u0935(.An(men_men_n956_), .Bn(men_men_n194_), .C(men_men_n957_), .Y(men_men_n958_));
  AOI210     u0936(.A0(men_men_n654_), .A1(men_men_n349_), .B0(men_men_n254_), .Y(men_men_n959_));
  NO2        u0937(.A(men_men_n959_), .B(men_men_n899_), .Y(men_men_n960_));
  NO3        u0938(.A(men_men_n960_), .B(men_men_n958_), .C(men_men_n955_), .Y(men_men_n961_));
  NOi21      u0939(.An(i_7_), .B(i_5_), .Y(men_men_n962_));
  NOi31      u0940(.An(men_men_n962_), .B(i_0_), .C(men_men_n772_), .Y(men_men_n963_));
  NA3        u0941(.A(men_men_n963_), .B(men_men_n407_), .C(i_6_), .Y(men_men_n964_));
  OA210      u0942(.A0(men_men_n957_), .A1(men_men_n555_), .B0(men_men_n964_), .Y(men_men_n965_));
  NO3        u0943(.A(men_men_n426_), .B(men_men_n385_), .C(men_men_n381_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n275_), .B(men_men_n338_), .Y(men_men_n967_));
  NO2        u0945(.A(men_men_n772_), .B(men_men_n270_), .Y(men_men_n968_));
  AOI210     u0946(.A0(men_men_n968_), .A1(men_men_n967_), .B0(men_men_n966_), .Y(men_men_n969_));
  NA4        u0947(.A(men_men_n969_), .B(men_men_n965_), .C(men_men_n961_), .D(men_men_n953_), .Y(men_men_n970_));
  NO2        u0948(.A(men_men_n916_), .B(men_men_n250_), .Y(men_men_n971_));
  AN2        u0949(.A(men_men_n353_), .B(men_men_n349_), .Y(men_men_n972_));
  AO220      u0950(.A0(men_men_n972_), .A1(men_men_n912_), .B0(men_men_n368_), .B1(men_men_n27_), .Y(men_men_n973_));
  OAI210     u0951(.A0(men_men_n973_), .A1(men_men_n971_), .B0(i_10_), .Y(men_men_n974_));
  OA210      u0952(.A0(men_men_n507_), .A1(men_men_n233_), .B0(men_men_n506_), .Y(men_men_n975_));
  NA3        u0953(.A(men_men_n506_), .B(men_men_n435_), .C(men_men_n46_), .Y(men_men_n976_));
  OAI210     u0954(.A0(men_men_n920_), .A1(men_men_n929_), .B0(men_men_n976_), .Y(men_men_n977_));
  NO2        u0955(.A(men_men_n268_), .B(men_men_n47_), .Y(men_men_n978_));
  NA2        u0956(.A(men_men_n947_), .B(men_men_n324_), .Y(men_men_n979_));
  OAI210     u0957(.A0(men_men_n978_), .A1(men_men_n193_), .B0(men_men_n979_), .Y(men_men_n980_));
  AOI220     u0958(.A0(men_men_n980_), .A1(men_men_n507_), .B0(men_men_n977_), .B1(men_men_n73_), .Y(men_men_n981_));
  NA3        u0959(.A(men_men_n864_), .B(men_men_n405_), .C(men_men_n690_), .Y(men_men_n982_));
  NA2        u0960(.A(men_men_n95_), .B(men_men_n45_), .Y(men_men_n983_));
  NO2        u0961(.A(men_men_n75_), .B(men_men_n796_), .Y(men_men_n984_));
  AOI220     u0962(.A0(men_men_n984_), .A1(men_men_n983_), .B0(men_men_n179_), .B1(men_men_n643_), .Y(men_men_n985_));
  AOI210     u0963(.A0(men_men_n985_), .A1(men_men_n982_), .B0(men_men_n48_), .Y(men_men_n986_));
  NO3        u0964(.A(men_men_n635_), .B(men_men_n380_), .C(men_men_n24_), .Y(men_men_n987_));
  AOI210     u0965(.A0(men_men_n749_), .A1(men_men_n589_), .B0(men_men_n987_), .Y(men_men_n988_));
  NO2        u0966(.A(men_men_n648_), .B(men_men_n108_), .Y(men_men_n989_));
  NA2        u0967(.A(men_men_n989_), .B(i_0_), .Y(men_men_n990_));
  OAI220     u0968(.A0(men_men_n990_), .A1(men_men_n86_), .B0(men_men_n988_), .B1(men_men_n177_), .Y(men_men_n991_));
  NO3        u0969(.A(men_men_n991_), .B(men_men_n986_), .C(men_men_n559_), .Y(men_men_n992_));
  NA3        u0970(.A(men_men_n992_), .B(men_men_n981_), .C(men_men_n974_), .Y(men_men_n993_));
  NO3        u0971(.A(men_men_n993_), .B(men_men_n970_), .C(men_men_n942_), .Y(men_men_n994_));
  NO2        u0972(.A(i_0_), .B(men_men_n772_), .Y(men_men_n995_));
  NA2        u0973(.A(men_men_n73_), .B(men_men_n45_), .Y(men_men_n996_));
  NA2        u0974(.A(men_men_n935_), .B(men_men_n996_), .Y(men_men_n997_));
  NO3        u0975(.A(men_men_n108_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n998_));
  AO220      u0976(.A0(men_men_n998_), .A1(men_men_n997_), .B0(men_men_n995_), .B1(men_men_n179_), .Y(men_men_n999_));
  NO2        u0977(.A(men_men_n843_), .B(men_men_n957_), .Y(men_men_n1000_));
  AOI210     u0978(.A0(men_men_n999_), .A1(men_men_n370_), .B0(men_men_n1000_), .Y(men_men_n1001_));
  NA2        u0979(.A(men_men_n782_), .B(men_men_n149_), .Y(men_men_n1002_));
  INV        u0980(.A(men_men_n1002_), .Y(men_men_n1003_));
  NA3        u0981(.A(men_men_n1003_), .B(men_men_n722_), .C(men_men_n73_), .Y(men_men_n1004_));
  NO2        u0982(.A(men_men_n860_), .B(men_men_n426_), .Y(men_men_n1005_));
  NA3        u0983(.A(men_men_n889_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n1006_));
  NA2        u0984(.A(men_men_n890_), .B(i_9_), .Y(men_men_n1007_));
  AOI210     u0985(.A0(men_men_n1006_), .A1(men_men_n535_), .B0(men_men_n1007_), .Y(men_men_n1008_));
  OAI210     u0986(.A0(men_men_n255_), .A1(i_9_), .B0(men_men_n240_), .Y(men_men_n1009_));
  AOI210     u0987(.A0(men_men_n1009_), .A1(men_men_n925_), .B0(men_men_n157_), .Y(men_men_n1010_));
  NO3        u0988(.A(men_men_n1010_), .B(men_men_n1008_), .C(men_men_n1005_), .Y(men_men_n1011_));
  NA3        u0989(.A(men_men_n1011_), .B(men_men_n1004_), .C(men_men_n1001_), .Y(men_men_n1012_));
  NA2        u0990(.A(men_men_n972_), .B(men_men_n395_), .Y(men_men_n1013_));
  AOI210     u0991(.A0(men_men_n318_), .A1(men_men_n166_), .B0(men_men_n1013_), .Y(men_men_n1014_));
  NA3        u0992(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n1015_));
  NA2        u0993(.A(men_men_n944_), .B(men_men_n523_), .Y(men_men_n1016_));
  AOI210     u0994(.A0(men_men_n1015_), .A1(men_men_n166_), .B0(men_men_n1016_), .Y(men_men_n1017_));
  NO2        u0995(.A(men_men_n1017_), .B(men_men_n1014_), .Y(men_men_n1018_));
  NO3        u0996(.A(men_men_n935_), .B(men_men_n908_), .C(men_men_n196_), .Y(men_men_n1019_));
  AOI220     u0997(.A0(men_men_n1019_), .A1(i_11_), .B0(men_men_n613_), .B1(men_men_n75_), .Y(men_men_n1020_));
  NO3        u0998(.A(men_men_n218_), .B(men_men_n406_), .C(i_0_), .Y(men_men_n1021_));
  OAI210     u0999(.A0(men_men_n1021_), .A1(men_men_n76_), .B0(i_13_), .Y(men_men_n1022_));
  INV        u1000(.A(men_men_n227_), .Y(men_men_n1023_));
  OAI220     u1001(.A0(men_men_n571_), .A1(men_men_n142_), .B0(men_men_n695_), .B1(men_men_n665_), .Y(men_men_n1024_));
  NA3        u1002(.A(men_men_n1024_), .B(i_7_), .C(men_men_n1023_), .Y(men_men_n1025_));
  NA4        u1003(.A(men_men_n1025_), .B(men_men_n1022_), .C(men_men_n1020_), .D(men_men_n1018_), .Y(men_men_n1026_));
  NO2        u1004(.A(men_men_n253_), .B(men_men_n95_), .Y(men_men_n1027_));
  AOI210     u1005(.A0(men_men_n1027_), .A1(men_men_n995_), .B0(men_men_n112_), .Y(men_men_n1028_));
  AOI220     u1006(.A0(men_men_n962_), .A1(men_men_n523_), .B0(men_men_n889_), .B1(men_men_n167_), .Y(men_men_n1029_));
  NA2        u1007(.A(men_men_n373_), .B(men_men_n181_), .Y(men_men_n1030_));
  OA220      u1008(.A0(men_men_n1030_), .A1(men_men_n1029_), .B0(men_men_n1028_), .B1(i_5_), .Y(men_men_n1031_));
  AOI210     u1009(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n180_), .Y(men_men_n1032_));
  NA2        u1010(.A(men_men_n1032_), .B(men_men_n975_), .Y(men_men_n1033_));
  NA3        u1011(.A(men_men_n662_), .B(men_men_n191_), .C(men_men_n84_), .Y(men_men_n1034_));
  NA2        u1012(.A(men_men_n1034_), .B(men_men_n587_), .Y(men_men_n1035_));
  NO3        u1013(.A(men_men_n899_), .B(men_men_n55_), .C(men_men_n49_), .Y(men_men_n1036_));
  NA3        u1014(.A(men_men_n528_), .B(men_men_n521_), .C(men_men_n504_), .Y(men_men_n1037_));
  NO3        u1015(.A(men_men_n1037_), .B(men_men_n1036_), .C(men_men_n1035_), .Y(men_men_n1038_));
  NA3        u1016(.A(men_men_n413_), .B(men_men_n176_), .C(men_men_n175_), .Y(men_men_n1039_));
  NA3        u1017(.A(men_men_n944_), .B(men_men_n307_), .C(men_men_n240_), .Y(men_men_n1040_));
  NA2        u1018(.A(men_men_n1040_), .B(men_men_n1039_), .Y(men_men_n1041_));
  NA3        u1019(.A(men_men_n413_), .B(men_men_n355_), .C(men_men_n231_), .Y(men_men_n1042_));
  OAI210     u1020(.A0(men_men_n903_), .A1(men_men_n699_), .B0(men_men_n1042_), .Y(men_men_n1043_));
  NOi31      u1021(.An(men_men_n412_), .B(men_men_n996_), .C(men_men_n250_), .Y(men_men_n1044_));
  NO3        u1022(.A(men_men_n943_), .B(men_men_n227_), .C(men_men_n196_), .Y(men_men_n1045_));
  NO4        u1023(.A(men_men_n1045_), .B(men_men_n1044_), .C(men_men_n1043_), .D(men_men_n1041_), .Y(men_men_n1046_));
  NA4        u1024(.A(men_men_n1046_), .B(men_men_n1038_), .C(men_men_n1033_), .D(men_men_n1031_), .Y(men_men_n1047_));
  INV        u1025(.A(men_men_n664_), .Y(men_men_n1048_));
  NO3        u1026(.A(men_men_n1048_), .B(men_men_n603_), .C(men_men_n367_), .Y(men_men_n1049_));
  INV        u1027(.A(men_men_n1049_), .Y(men_men_n1050_));
  NA3        u1028(.A(men_men_n324_), .B(i_5_), .C(men_men_n199_), .Y(men_men_n1051_));
  NAi31      u1029(.An(men_men_n252_), .B(men_men_n1051_), .C(men_men_n253_), .Y(men_men_n1052_));
  NO4        u1030(.A(men_men_n250_), .B(men_men_n218_), .C(i_0_), .D(i_12_), .Y(men_men_n1053_));
  NA2        u1031(.A(men_men_n1053_), .B(men_men_n1052_), .Y(men_men_n1054_));
  AN2        u1032(.A(men_men_n935_), .B(men_men_n157_), .Y(men_men_n1055_));
  NO4        u1033(.A(men_men_n1055_), .B(i_12_), .C(men_men_n699_), .D(men_men_n134_), .Y(men_men_n1056_));
  NA2        u1034(.A(men_men_n1056_), .B(men_men_n227_), .Y(men_men_n1057_));
  NA3        u1035(.A(men_men_n101_), .B(men_men_n617_), .C(i_11_), .Y(men_men_n1058_));
  NO2        u1036(.A(men_men_n1058_), .B(men_men_n159_), .Y(men_men_n1059_));
  NA2        u1037(.A(men_men_n962_), .B(men_men_n503_), .Y(men_men_n1060_));
  NA2        u1038(.A(men_men_n64_), .B(men_men_n104_), .Y(men_men_n1061_));
  OAI220     u1039(.A0(men_men_n1061_), .A1(men_men_n1051_), .B0(men_men_n1060_), .B1(men_men_n723_), .Y(men_men_n1062_));
  AOI210     u1040(.A0(men_men_n1062_), .A1(men_men_n948_), .B0(men_men_n1059_), .Y(men_men_n1063_));
  NA4        u1041(.A(men_men_n1063_), .B(men_men_n1057_), .C(men_men_n1054_), .D(men_men_n1050_), .Y(men_men_n1064_));
  NO4        u1042(.A(men_men_n1064_), .B(men_men_n1047_), .C(men_men_n1026_), .D(men_men_n1012_), .Y(men_men_n1065_));
  OAI210     u1043(.A0(men_men_n863_), .A1(men_men_n856_), .B0(men_men_n37_), .Y(men_men_n1066_));
  NA3        u1044(.A(men_men_n956_), .B(men_men_n390_), .C(i_5_), .Y(men_men_n1067_));
  NA3        u1045(.A(men_men_n1067_), .B(men_men_n1066_), .C(men_men_n660_), .Y(men_men_n1068_));
  NA2        u1046(.A(men_men_n1068_), .B(men_men_n214_), .Y(men_men_n1069_));
  BUFFER     u1047(.A(men_men_n391_), .Y(men_men_n1070_));
  NA2        u1048(.A(men_men_n192_), .B(men_men_n194_), .Y(men_men_n1071_));
  AO210      u1049(.A0(men_men_n1070_), .A1(men_men_n33_), .B0(men_men_n1071_), .Y(men_men_n1072_));
  OAI210     u1050(.A0(men_men_n664_), .A1(men_men_n662_), .B0(men_men_n337_), .Y(men_men_n1073_));
  NAi31      u1051(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1074_));
  AOI210     u1052(.A0(men_men_n120_), .A1(men_men_n70_), .B0(men_men_n1074_), .Y(men_men_n1075_));
  NO2        u1053(.A(men_men_n1075_), .B(men_men_n696_), .Y(men_men_n1076_));
  NA3        u1054(.A(men_men_n1076_), .B(men_men_n1073_), .C(men_men_n1072_), .Y(men_men_n1077_));
  NO2        u1055(.A(men_men_n493_), .B(men_men_n281_), .Y(men_men_n1078_));
  NO4        u1056(.A(men_men_n243_), .B(men_men_n148_), .C(men_men_n726_), .D(men_men_n37_), .Y(men_men_n1079_));
  NO3        u1057(.A(men_men_n1079_), .B(men_men_n1078_), .C(men_men_n927_), .Y(men_men_n1080_));
  OAI210     u1058(.A0(men_men_n1058_), .A1(men_men_n151_), .B0(men_men_n1080_), .Y(men_men_n1081_));
  AOI210     u1059(.A0(men_men_n1077_), .A1(men_men_n49_), .B0(men_men_n1081_), .Y(men_men_n1082_));
  AOI210     u1060(.A0(men_men_n1082_), .A1(men_men_n1069_), .B0(men_men_n73_), .Y(men_men_n1083_));
  NO2        u1061(.A(men_men_n610_), .B(men_men_n402_), .Y(men_men_n1084_));
  NO2        u1062(.A(men_men_n1084_), .B(men_men_n802_), .Y(men_men_n1085_));
  OAI210     u1063(.A0(men_men_n80_), .A1(men_men_n55_), .B0(men_men_n111_), .Y(men_men_n1086_));
  NA2        u1064(.A(men_men_n1086_), .B(men_men_n76_), .Y(men_men_n1087_));
  AOI210     u1065(.A0(men_men_n1032_), .A1(men_men_n944_), .B0(men_men_n963_), .Y(men_men_n1088_));
  AOI210     u1066(.A0(men_men_n1088_), .A1(men_men_n1087_), .B0(men_men_n726_), .Y(men_men_n1089_));
  NA2        u1067(.A(men_men_n275_), .B(men_men_n57_), .Y(men_men_n1090_));
  AOI220     u1068(.A0(men_men_n1090_), .A1(men_men_n76_), .B0(men_men_n368_), .B1(men_men_n267_), .Y(men_men_n1091_));
  NO2        u1069(.A(men_men_n1091_), .B(men_men_n247_), .Y(men_men_n1092_));
  NA3        u1070(.A(men_men_n99_), .B(men_men_n326_), .C(men_men_n31_), .Y(men_men_n1093_));
  INV        u1071(.A(men_men_n1093_), .Y(men_men_n1094_));
  NO3        u1072(.A(men_men_n1094_), .B(men_men_n1092_), .C(men_men_n1089_), .Y(men_men_n1095_));
  OAI210     u1073(.A0(men_men_n283_), .A1(men_men_n162_), .B0(men_men_n89_), .Y(men_men_n1096_));
  NA3        u1074(.A(men_men_n806_), .B(men_men_n307_), .C(men_men_n80_), .Y(men_men_n1097_));
  AOI210     u1075(.A0(men_men_n1097_), .A1(men_men_n1096_), .B0(i_11_), .Y(men_men_n1098_));
  NA2        u1076(.A(men_men_n655_), .B(men_men_n224_), .Y(men_men_n1099_));
  OAI210     u1077(.A0(men_men_n1099_), .A1(men_men_n956_), .B0(men_men_n214_), .Y(men_men_n1100_));
  NA2        u1078(.A(men_men_n168_), .B(i_5_), .Y(men_men_n1101_));
  NO2        u1079(.A(men_men_n1100_), .B(men_men_n1101_), .Y(men_men_n1102_));
  NO3        u1080(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1103_));
  OAI210     u1081(.A0(men_men_n967_), .A1(men_men_n326_), .B0(men_men_n1103_), .Y(men_men_n1104_));
  NO2        u1082(.A(men_men_n1104_), .B(men_men_n772_), .Y(men_men_n1105_));
  NO2        u1083(.A(men_men_n859_), .B(men_men_n386_), .Y(men_men_n1106_));
  NO2        u1084(.A(men_men_n1106_), .B(men_men_n41_), .Y(men_men_n1107_));
  NO4        u1085(.A(men_men_n1107_), .B(men_men_n1105_), .C(men_men_n1102_), .D(men_men_n1098_), .Y(men_men_n1108_));
  OAI210     u1086(.A0(men_men_n1095_), .A1(i_4_), .B0(men_men_n1108_), .Y(men_men_n1109_));
  NO3        u1087(.A(men_men_n1109_), .B(men_men_n1085_), .C(men_men_n1083_), .Y(men_men_n1110_));
  NA4        u1088(.A(men_men_n1110_), .B(men_men_n1065_), .C(men_men_n994_), .D(men_men_n915_), .Y(men4));
  INV        u1089(.A(i_2_), .Y(men_men_n1114_));
  INV        u1090(.A(men_men_n761_), .Y(men_men_n1115_));
  INV        u1091(.A(men_men_n518_), .Y(men_men_n1116_));
  INV        u1092(.A(i_7_), .Y(men_men_n1117_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule