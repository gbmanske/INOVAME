// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n137_, new_new_n138_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n537_, new_new_n538_,
    new_new_n539_, new_new_n540_, new_new_n541_, new_new_n542_,
    new_new_n543_, new_new_n544_, new_new_n545_, new_new_n546_,
    new_new_n547_, new_new_n548_, new_new_n549_, new_new_n550_,
    new_new_n551_, new_new_n552_, new_new_n553_, new_new_n554_,
    new_new_n555_, new_new_n556_, new_new_n557_, new_new_n558_,
    new_new_n559_, new_new_n560_, new_new_n561_, new_new_n562_,
    new_new_n563_, new_new_n564_, new_new_n565_, new_new_n566_,
    new_new_n567_, new_new_n568_, new_new_n569_, new_new_n570_,
    new_new_n571_, new_new_n572_, new_new_n573_, new_new_n574_,
    new_new_n575_, new_new_n576_, new_new_n577_, new_new_n578_,
    new_new_n579_, new_new_n580_, new_new_n581_, new_new_n582_,
    new_new_n583_, new_new_n585_, new_new_n586_, new_new_n587_,
    new_new_n588_, new_new_n589_, new_new_n590_, new_new_n591_,
    new_new_n592_, new_new_n593_, new_new_n594_, new_new_n595_,
    new_new_n596_, new_new_n597_, new_new_n598_, new_new_n599_,
    new_new_n600_, new_new_n601_, new_new_n602_, new_new_n603_,
    new_new_n604_, new_new_n605_, new_new_n606_, new_new_n607_,
    new_new_n608_, new_new_n609_, new_new_n610_, new_new_n611_,
    new_new_n612_, new_new_n613_, new_new_n614_, new_new_n615_,
    new_new_n616_, new_new_n617_, new_new_n618_, new_new_n619_,
    new_new_n620_, new_new_n621_, new_new_n622_, new_new_n623_,
    new_new_n624_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n653_, new_new_n654_, new_new_n655_, new_new_n656_,
    new_new_n657_, new_new_n658_, new_new_n659_, new_new_n660_,
    new_new_n661_, new_new_n662_, new_new_n663_, new_new_n664_,
    new_new_n665_, new_new_n666_, new_new_n667_, new_new_n668_,
    new_new_n669_, new_new_n670_, new_new_n671_, new_new_n672_,
    new_new_n673_, new_new_n674_, new_new_n675_, new_new_n676_,
    new_new_n677_, new_new_n678_, new_new_n679_, new_new_n680_,
    new_new_n681_, new_new_n682_, new_new_n683_, new_new_n684_,
    new_new_n685_, new_new_n686_, new_new_n687_, new_new_n688_,
    new_new_n689_, new_new_n690_, new_new_n691_, new_new_n692_,
    new_new_n693_, new_new_n694_, new_new_n695_, new_new_n696_,
    new_new_n697_, new_new_n698_, new_new_n699_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n703_, new_new_n704_,
    new_new_n705_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n752_, new_new_n753_, new_new_n754_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  NAi21      g036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g037(.A(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA3        g039(.A(new_new_n61_), .B(new_new_n59_), .C(new_new_n31_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_10_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NAi21      g042(.An(new_new_n64_), .B(new_new_n62_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n50_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NA2        g055(.A(i_2_), .B(i_8_), .Y(new_new_n78_));
  NO2        g056(.A(new_new_n78_), .B(new_new_n57_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_9_), .Y(new_new_n80_));
  NO2        g058(.A(i_3_), .B(i_7_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n80_), .B(new_new_n60_), .Y(new_new_n82_));
  INV        g060(.A(i_6_), .Y(new_new_n83_));
  OR4        g061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n84_));
  INV        g062(.A(new_new_n84_), .Y(new_new_n85_));
  NO2        g063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  NO2        g064(.A(new_new_n85_), .B(new_new_n86_), .Y(new_new_n87_));
  OAI210     g065(.A0(new_new_n82_), .A1(new_new_n79_), .B0(new_new_n87_), .Y(new_new_n88_));
  NAi21      g066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n60_), .Y(new_new_n91_));
  NA2        g069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g070(.A(new_new_n92_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g072(.A0(new_new_n94_), .A1(new_new_n88_), .B0(new_new_n77_), .Y(new_new_n95_));
  AN3        g073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n96_), .B(new_new_n32_), .Y(new_new_n98_));
  INV        g076(.A(i_7_), .Y(new_new_n99_));
  NA2        g077(.A(new_new_n46_), .B(new_new_n99_), .Y(new_new_n100_));
  NO2        g078(.A(i_0_), .B(i_5_), .Y(new_new_n101_));
  NO2        g079(.A(new_new_n101_), .B(new_new_n83_), .Y(new_new_n102_));
  NA2        g080(.A(i_12_), .B(i_3_), .Y(new_new_n103_));
  INV        g081(.A(new_new_n103_), .Y(new_new_n104_));
  NA3        g082(.A(new_new_n104_), .B(new_new_n102_), .C(new_new_n100_), .Y(new_new_n105_));
  NAi21      g083(.An(i_7_), .B(i_11_), .Y(new_new_n106_));
  NO3        g084(.A(new_new_n106_), .B(new_new_n89_), .C(new_new_n53_), .Y(new_new_n107_));
  AN2        g085(.A(i_2_), .B(i_10_), .Y(new_new_n108_));
  NO2        g086(.A(new_new_n108_), .B(i_7_), .Y(new_new_n109_));
  OR2        g087(.A(new_new_n77_), .B(new_new_n57_), .Y(new_new_n110_));
  NO2        g088(.A(i_8_), .B(new_new_n99_), .Y(new_new_n111_));
  NO3        g089(.A(new_new_n111_), .B(new_new_n110_), .C(new_new_n109_), .Y(new_new_n112_));
  NA2        g090(.A(i_12_), .B(i_7_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n60_), .B(new_new_n26_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n114_), .B(i_0_), .Y(new_new_n115_));
  NA2        g093(.A(i_11_), .B(i_12_), .Y(new_new_n116_));
  OAI210     g094(.A0(new_new_n115_), .A1(new_new_n113_), .B0(new_new_n116_), .Y(new_new_n117_));
  NO2        g095(.A(new_new_n117_), .B(new_new_n112_), .Y(new_new_n118_));
  NAi41      g096(.An(new_new_n107_), .B(new_new_n118_), .C(new_new_n105_), .D(new_new_n98_), .Y(new_new_n119_));
  NOi21      g097(.An(i_1_), .B(i_5_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(i_11_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n122_));
  NA2        g100(.A(i_7_), .B(new_new_n25_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n122_), .Y(new_new_n124_));
  NO2        g102(.A(new_new_n124_), .B(new_new_n46_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n126_));
  NAi21      g104(.An(i_3_), .B(i_8_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(new_new_n59_), .Y(new_new_n128_));
  NOi31      g106(.An(new_new_n128_), .B(new_new_n126_), .C(new_new_n125_), .Y(new_new_n129_));
  NO2        g107(.A(i_1_), .B(new_new_n83_), .Y(new_new_n130_));
  NO2        g108(.A(i_6_), .B(i_5_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(i_3_), .Y(new_new_n132_));
  AO210      g110(.A0(new_new_n132_), .A1(new_new_n47_), .B0(new_new_n130_), .Y(new_new_n133_));
  OAI220     g111(.A0(new_new_n133_), .A1(new_new_n106_), .B0(new_new_n129_), .B1(new_new_n121_), .Y(new_new_n134_));
  NO3        g112(.A(new_new_n134_), .B(new_new_n119_), .C(new_new_n95_), .Y(new_new_n135_));
  NA3        g113(.A(new_new_n135_), .B(new_new_n76_), .C(new_new_n56_), .Y(ori2));
  NO2        g114(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n137_));
  NA2        g115(.A(new_new_n754_), .B(new_new_n137_), .Y(new_new_n138_));
  NA4        g116(.A(new_new_n138_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(ori0));
  NO2        g117(.A(i_12_), .B(i_13_), .Y(new_new_n140_));
  NAi21      g118(.An(i_5_), .B(i_11_), .Y(new_new_n141_));
  NO2        g119(.A(i_0_), .B(i_1_), .Y(new_new_n142_));
  NA2        g120(.A(i_2_), .B(i_3_), .Y(new_new_n143_));
  NO2        g121(.A(new_new_n143_), .B(i_4_), .Y(new_new_n144_));
  NA2        g122(.A(i_1_), .B(i_5_), .Y(new_new_n145_));
  OR2        g123(.A(i_0_), .B(i_1_), .Y(new_new_n146_));
  NAi32      g124(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n147_));
  NOi21      g125(.An(i_4_), .B(i_10_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n40_), .Y(new_new_n149_));
  NOi21      g127(.An(i_4_), .B(i_9_), .Y(new_new_n150_));
  NOi21      g128(.An(i_11_), .B(i_13_), .Y(new_new_n151_));
  NA2        g129(.A(new_new_n151_), .B(new_new_n150_), .Y(new_new_n152_));
  NO2        g130(.A(i_4_), .B(i_5_), .Y(new_new_n153_));
  NAi21      g131(.An(i_12_), .B(i_11_), .Y(new_new_n154_));
  NO2        g132(.A(new_new_n154_), .B(i_13_), .Y(new_new_n155_));
  NO2        g133(.A(new_new_n70_), .B(new_new_n60_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n70_), .B(i_5_), .Y(new_new_n157_));
  NO2        g135(.A(i_13_), .B(i_10_), .Y(new_new_n158_));
  NO2        g136(.A(i_2_), .B(i_1_), .Y(new_new_n159_));
  NAi21      g137(.An(i_4_), .B(i_12_), .Y(new_new_n160_));
  INV        g138(.A(i_8_), .Y(new_new_n161_));
  NO3        g139(.A(i_3_), .B(new_new_n83_), .C(new_new_n48_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n162_), .B(new_new_n111_), .Y(new_new_n163_));
  NO3        g141(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n164_));
  NO2        g142(.A(i_3_), .B(i_8_), .Y(new_new_n165_));
  NO3        g143(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n166_));
  NA3        g144(.A(new_new_n166_), .B(new_new_n165_), .C(new_new_n40_), .Y(new_new_n167_));
  NO2        g145(.A(new_new_n101_), .B(new_new_n57_), .Y(new_new_n168_));
  INV        g146(.A(new_new_n168_), .Y(new_new_n169_));
  NO2        g147(.A(i_13_), .B(i_9_), .Y(new_new_n170_));
  NAi21      g148(.An(i_12_), .B(i_3_), .Y(new_new_n171_));
  NO2        g149(.A(new_new_n44_), .B(i_5_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n169_), .B(new_new_n167_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(i_7_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n174_), .B(i_4_), .Y(new_new_n175_));
  NAi21      g153(.An(i_12_), .B(i_7_), .Y(new_new_n176_));
  NA3        g154(.A(i_13_), .B(new_new_n161_), .C(i_10_), .Y(new_new_n177_));
  NA2        g155(.A(i_0_), .B(i_5_), .Y(new_new_n178_));
  NAi31      g156(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n36_), .B(i_13_), .Y(new_new_n180_));
  NO2        g158(.A(new_new_n70_), .B(new_new_n26_), .Y(new_new_n181_));
  NO2        g159(.A(new_new_n46_), .B(new_new_n60_), .Y(new_new_n182_));
  INV        g160(.A(i_13_), .Y(new_new_n183_));
  NO2        g161(.A(i_12_), .B(new_new_n183_), .Y(new_new_n184_));
  NO2        g162(.A(i_12_), .B(new_new_n37_), .Y(new_new_n185_));
  OR2        g163(.A(i_8_), .B(i_7_), .Y(new_new_n186_));
  INV        g164(.A(i_12_), .Y(new_new_n187_));
  NO3        g165(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n188_));
  NA2        g166(.A(i_2_), .B(i_1_), .Y(new_new_n189_));
  NO3        g167(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n190_));
  NAi21      g168(.An(i_4_), .B(i_3_), .Y(new_new_n191_));
  NO2        g169(.A(i_0_), .B(i_6_), .Y(new_new_n192_));
  NOi41      g170(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n193_));
  NA2        g171(.A(new_new_n193_), .B(new_new_n192_), .Y(new_new_n194_));
  NO2        g172(.A(i_11_), .B(new_new_n183_), .Y(new_new_n195_));
  NOi21      g173(.An(i_1_), .B(i_6_), .Y(new_new_n196_));
  NAi21      g174(.An(i_3_), .B(i_7_), .Y(new_new_n197_));
  NA2        g175(.A(new_new_n187_), .B(i_9_), .Y(new_new_n198_));
  OR4        g176(.A(new_new_n198_), .B(new_new_n197_), .C(new_new_n196_), .D(new_new_n157_), .Y(new_new_n199_));
  NA2        g177(.A(new_new_n70_), .B(i_5_), .Y(new_new_n200_));
  NA2        g178(.A(i_3_), .B(i_9_), .Y(new_new_n201_));
  NAi21      g179(.An(i_7_), .B(i_10_), .Y(new_new_n202_));
  NO2        g180(.A(new_new_n202_), .B(new_new_n201_), .Y(new_new_n203_));
  NA3        g181(.A(new_new_n203_), .B(new_new_n200_), .C(new_new_n61_), .Y(new_new_n204_));
  NA2        g182(.A(new_new_n204_), .B(new_new_n199_), .Y(new_new_n205_));
  NA2        g183(.A(new_new_n205_), .B(new_new_n195_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n186_), .B(new_new_n37_), .Y(new_new_n207_));
  NA2        g185(.A(i_12_), .B(i_6_), .Y(new_new_n208_));
  OR2        g186(.A(i_13_), .B(i_9_), .Y(new_new_n209_));
  NO3        g187(.A(new_new_n209_), .B(new_new_n208_), .C(new_new_n48_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n191_), .B(i_2_), .Y(new_new_n211_));
  NA3        g189(.A(new_new_n211_), .B(new_new_n210_), .C(new_new_n44_), .Y(new_new_n212_));
  NA2        g190(.A(new_new_n195_), .B(i_9_), .Y(new_new_n213_));
  NA2        g191(.A(new_new_n200_), .B(new_new_n61_), .Y(new_new_n214_));
  OAI210     g192(.A0(new_new_n214_), .A1(new_new_n213_), .B0(new_new_n212_), .Y(new_new_n215_));
  NO3        g193(.A(i_11_), .B(new_new_n183_), .C(new_new_n25_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n197_), .B(i_8_), .Y(new_new_n217_));
  NA2        g195(.A(new_new_n215_), .B(new_new_n207_), .Y(new_new_n218_));
  NA2        g196(.A(new_new_n218_), .B(new_new_n206_), .Y(new_new_n219_));
  NO3        g197(.A(i_12_), .B(new_new_n183_), .C(new_new_n37_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n189_), .B(i_0_), .Y(new_new_n221_));
  NO2        g199(.A(i_3_), .B(i_10_), .Y(new_new_n222_));
  NO2        g200(.A(i_2_), .B(new_new_n99_), .Y(new_new_n223_));
  AN2        g201(.A(i_3_), .B(i_10_), .Y(new_new_n224_));
  NO2        g202(.A(i_5_), .B(new_new_n37_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n219_), .B(new_new_n175_), .Y(new_new_n227_));
  NO3        g205(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n228_));
  NO2        g206(.A(i_2_), .B(i_3_), .Y(new_new_n229_));
  OR2        g207(.A(i_0_), .B(i_5_), .Y(new_new_n230_));
  NO2        g208(.A(i_12_), .B(i_10_), .Y(new_new_n231_));
  NOi21      g209(.An(i_5_), .B(i_0_), .Y(new_new_n232_));
  NO2        g210(.A(i_2_), .B(new_new_n99_), .Y(new_new_n233_));
  NO4        g211(.A(new_new_n233_), .B(i_4_), .C(new_new_n232_), .D(new_new_n127_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n234_), .B(new_new_n231_), .Y(new_new_n235_));
  NO2        g213(.A(i_6_), .B(i_8_), .Y(new_new_n236_));
  NO2        g214(.A(i_1_), .B(i_7_), .Y(new_new_n237_));
  INV        g215(.A(new_new_n235_), .Y(new_new_n238_));
  NOi21      g216(.An(new_new_n145_), .B(new_new_n102_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n239_), .B(new_new_n123_), .Y(new_new_n240_));
  NA2        g218(.A(new_new_n240_), .B(i_3_), .Y(new_new_n241_));
  NO2        g219(.A(new_new_n161_), .B(i_9_), .Y(new_new_n242_));
  NA2        g220(.A(new_new_n242_), .B(new_new_n168_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n243_), .B(new_new_n46_), .Y(new_new_n244_));
  INV        g222(.A(new_new_n244_), .Y(new_new_n245_));
  AOI210     g223(.A0(new_new_n245_), .A1(new_new_n241_), .B0(new_new_n149_), .Y(new_new_n246_));
  AOI210     g224(.A0(new_new_n238_), .A1(new_new_n228_), .B0(new_new_n246_), .Y(new_new_n247_));
  NOi32      g225(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n248_));
  INV        g226(.A(new_new_n248_), .Y(new_new_n249_));
  NAi21      g227(.An(i_0_), .B(i_6_), .Y(new_new_n250_));
  NAi21      g228(.An(i_1_), .B(i_5_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n251_), .B(new_new_n250_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n252_), .B(new_new_n25_), .Y(new_new_n253_));
  OAI210     g231(.A0(new_new_n253_), .A1(new_new_n147_), .B0(new_new_n194_), .Y(new_new_n254_));
  NAi41      g232(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n255_));
  OAI220     g233(.A0(new_new_n255_), .A1(new_new_n251_), .B0(new_new_n179_), .B1(new_new_n147_), .Y(new_new_n256_));
  AOI210     g234(.A0(new_new_n255_), .A1(new_new_n147_), .B0(new_new_n146_), .Y(new_new_n257_));
  NOi32      g235(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n258_));
  NAi21      g236(.An(i_6_), .B(i_1_), .Y(new_new_n259_));
  NA3        g237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n46_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n260_), .B(i_0_), .Y(new_new_n261_));
  OR3        g239(.A(new_new_n261_), .B(new_new_n257_), .C(new_new_n256_), .Y(new_new_n262_));
  NO2        g240(.A(i_1_), .B(new_new_n99_), .Y(new_new_n263_));
  NAi21      g241(.An(i_3_), .B(i_4_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n264_), .B(i_9_), .Y(new_new_n265_));
  AN2        g243(.A(i_6_), .B(i_7_), .Y(new_new_n266_));
  NA2        g244(.A(i_2_), .B(i_7_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n264_), .B(i_10_), .Y(new_new_n268_));
  AOI210     g246(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n269_));
  OAI210     g247(.A0(new_new_n269_), .A1(new_new_n159_), .B0(new_new_n268_), .Y(new_new_n270_));
  AOI220     g248(.A0(new_new_n268_), .A1(new_new_n237_), .B0(new_new_n188_), .B1(new_new_n159_), .Y(new_new_n271_));
  AOI210     g249(.A0(new_new_n271_), .A1(new_new_n270_), .B0(i_5_), .Y(new_new_n272_));
  NO3        g250(.A(new_new_n272_), .B(new_new_n262_), .C(new_new_n254_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n273_), .B(new_new_n249_), .Y(new_new_n274_));
  AN2        g252(.A(i_12_), .B(i_5_), .Y(new_new_n275_));
  NA2        g253(.A(i_3_), .B(new_new_n275_), .Y(new_new_n276_));
  NO2        g254(.A(i_11_), .B(i_6_), .Y(new_new_n277_));
  NO2        g255(.A(i_5_), .B(i_10_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n279_));
  NO3        g257(.A(new_new_n83_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n280_));
  NA3        g258(.A(new_new_n222_), .B(new_new_n90_), .C(new_new_n72_), .Y(new_new_n281_));
  NO2        g259(.A(i_11_), .B(i_12_), .Y(new_new_n282_));
  NA2        g260(.A(new_new_n282_), .B(new_new_n36_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n281_), .B(new_new_n283_), .Y(new_new_n284_));
  NAi21      g262(.An(i_13_), .B(i_0_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n285_), .B(new_new_n189_), .Y(new_new_n286_));
  NA2        g264(.A(new_new_n284_), .B(new_new_n286_), .Y(new_new_n287_));
  INV        g265(.A(new_new_n287_), .Y(new_new_n288_));
  NO2        g266(.A(i_0_), .B(i_11_), .Y(new_new_n289_));
  NOi21      g267(.An(i_2_), .B(i_12_), .Y(new_new_n290_));
  NAi21      g268(.An(i_9_), .B(i_4_), .Y(new_new_n291_));
  OR2        g269(.A(i_13_), .B(i_10_), .Y(new_new_n292_));
  NO3        g270(.A(new_new_n292_), .B(new_new_n116_), .C(new_new_n291_), .Y(new_new_n293_));
  NO2        g271(.A(new_new_n152_), .B(new_new_n122_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n99_), .B(new_new_n25_), .Y(new_new_n295_));
  NA2        g273(.A(new_new_n220_), .B(new_new_n295_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n296_), .B(new_new_n239_), .Y(new_new_n297_));
  INV        g275(.A(new_new_n297_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n298_), .B(new_new_n26_), .Y(new_new_n299_));
  NA2        g277(.A(new_new_n161_), .B(i_10_), .Y(new_new_n300_));
  NA3        g278(.A(new_new_n200_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n301_), .B(new_new_n300_), .Y(new_new_n302_));
  INV        g280(.A(new_new_n302_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n303_), .B(new_new_n213_), .Y(new_new_n304_));
  NO4        g282(.A(new_new_n304_), .B(new_new_n299_), .C(new_new_n288_), .D(new_new_n274_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n70_), .B(i_13_), .Y(new_new_n306_));
  NO2        g284(.A(i_10_), .B(i_9_), .Y(new_new_n307_));
  NAi21      g285(.An(i_12_), .B(i_8_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n308_), .B(i_3_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n46_), .B(i_4_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n310_), .B(new_new_n102_), .Y(new_new_n311_));
  NO2        g289(.A(new_new_n311_), .B(new_new_n167_), .Y(new_new_n312_));
  NA2        g290(.A(new_new_n226_), .B(i_0_), .Y(new_new_n313_));
  NO3        g291(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n314_));
  NA2        g292(.A(new_new_n208_), .B(new_new_n97_), .Y(new_new_n315_));
  NA2        g293(.A(new_new_n315_), .B(new_new_n314_), .Y(new_new_n316_));
  NA2        g294(.A(i_8_), .B(i_9_), .Y(new_new_n317_));
  NA2        g295(.A(new_new_n220_), .B(new_new_n168_), .Y(new_new_n318_));
  OAI220     g296(.A0(new_new_n318_), .A1(new_new_n317_), .B0(new_new_n316_), .B1(new_new_n313_), .Y(new_new_n319_));
  NA2        g297(.A(new_new_n195_), .B(new_new_n225_), .Y(new_new_n320_));
  NO3        g298(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n321_));
  INV        g299(.A(new_new_n321_), .Y(new_new_n322_));
  NA3        g300(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n323_));
  NA4        g301(.A(new_new_n141_), .B(new_new_n114_), .C(new_new_n77_), .D(new_new_n23_), .Y(new_new_n324_));
  OAI220     g302(.A0(new_new_n324_), .A1(new_new_n323_), .B0(new_new_n322_), .B1(new_new_n320_), .Y(new_new_n325_));
  NO3        g303(.A(new_new_n325_), .B(new_new_n319_), .C(new_new_n312_), .Y(new_new_n326_));
  OR2        g304(.A(new_new_n243_), .B(new_new_n99_), .Y(new_new_n327_));
  OR2        g305(.A(new_new_n327_), .B(new_new_n149_), .Y(new_new_n328_));
  NO2        g306(.A(i_2_), .B(i_13_), .Y(new_new_n329_));
  NO3        g307(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n330_));
  NO2        g308(.A(i_6_), .B(i_7_), .Y(new_new_n331_));
  NO2        g309(.A(i_11_), .B(i_1_), .Y(new_new_n332_));
  OR2        g310(.A(i_11_), .B(i_8_), .Y(new_new_n333_));
  NOi21      g311(.An(i_2_), .B(i_7_), .Y(new_new_n334_));
  NO2        g312(.A(i_3_), .B(new_new_n161_), .Y(new_new_n335_));
  NO2        g313(.A(i_6_), .B(i_10_), .Y(new_new_n336_));
  NA3        g314(.A(new_new_n193_), .B(new_new_n151_), .C(new_new_n131_), .Y(new_new_n337_));
  NA2        g315(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n146_), .B(i_3_), .Y(new_new_n339_));
  NAi31      g317(.An(new_new_n338_), .B(new_new_n339_), .C(new_new_n184_), .Y(new_new_n340_));
  NA3        g318(.A(new_new_n279_), .B(new_new_n156_), .C(new_new_n144_), .Y(new_new_n341_));
  NA3        g319(.A(new_new_n341_), .B(new_new_n340_), .C(new_new_n337_), .Y(new_new_n342_));
  INV        g320(.A(new_new_n342_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n314_), .B(new_new_n275_), .Y(new_new_n344_));
  NAi21      g322(.An(new_new_n177_), .B(new_new_n282_), .Y(new_new_n345_));
  NA2        g323(.A(new_new_n237_), .B(new_new_n178_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n346_), .B(new_new_n345_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n228_), .B(new_new_n188_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(new_new_n301_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(new_new_n347_), .Y(new_new_n350_));
  NA4        g328(.A(new_new_n350_), .B(new_new_n343_), .C(new_new_n328_), .D(new_new_n326_), .Y(new_new_n351_));
  NA2        g329(.A(new_new_n121_), .B(new_new_n110_), .Y(new_new_n352_));
  AN2        g330(.A(new_new_n352_), .B(new_new_n314_), .Y(new_new_n353_));
  NA2        g331(.A(new_new_n353_), .B(new_new_n226_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n275_), .B(new_new_n183_), .Y(new_new_n355_));
  NA2        g333(.A(new_new_n248_), .B(new_new_n70_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n266_), .B(new_new_n258_), .Y(new_new_n357_));
  OR2        g335(.A(new_new_n355_), .B(new_new_n357_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n36_), .B(i_8_), .Y(new_new_n359_));
  AOI210     g337(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n293_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n360_), .B(new_new_n358_), .Y(new_new_n361_));
  INV        g339(.A(new_new_n361_), .Y(new_new_n362_));
  NA2        g340(.A(new_new_n200_), .B(new_new_n61_), .Y(new_new_n363_));
  OAI210     g341(.A0(i_8_), .A1(new_new_n363_), .B0(new_new_n133_), .Y(new_new_n364_));
  NA2        g342(.A(new_new_n364_), .B(new_new_n294_), .Y(new_new_n365_));
  NA3        g343(.A(new_new_n365_), .B(new_new_n362_), .C(new_new_n354_), .Y(new_new_n366_));
  NO2        g344(.A(i_12_), .B(new_new_n161_), .Y(new_new_n367_));
  NO2        g345(.A(i_8_), .B(i_7_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n44_), .B(i_10_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n369_), .B(i_6_), .Y(new_new_n370_));
  NA3        g348(.A(new_new_n224_), .B(new_new_n153_), .C(new_new_n96_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n146_), .B(i_5_), .Y(new_new_n372_));
  INV        g350(.A(new_new_n371_), .Y(new_new_n373_));
  NA2        g351(.A(new_new_n373_), .B(new_new_n321_), .Y(new_new_n374_));
  INV        g352(.A(new_new_n374_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n182_), .B(new_new_n181_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n307_), .B(new_new_n180_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n376_), .B(new_new_n377_), .Y(new_new_n378_));
  AOI210     g356(.A0(new_new_n259_), .A1(new_new_n46_), .B0(new_new_n263_), .Y(new_new_n379_));
  NA2        g357(.A(i_0_), .B(new_new_n48_), .Y(new_new_n380_));
  NA3        g358(.A(new_new_n367_), .B(new_new_n216_), .C(new_new_n380_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n379_), .B(new_new_n381_), .Y(new_new_n382_));
  NO2        g360(.A(new_new_n382_), .B(new_new_n378_), .Y(new_new_n383_));
  NO4        g361(.A(new_new_n196_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n384_));
  NO3        g362(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n292_), .B(i_1_), .Y(new_new_n386_));
  NOi31      g364(.An(new_new_n386_), .B(new_new_n315_), .C(new_new_n70_), .Y(new_new_n387_));
  NOi21      g365(.An(i_10_), .B(i_6_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n83_), .B(new_new_n25_), .Y(new_new_n389_));
  AOI220     g367(.A0(new_new_n220_), .A1(new_new_n389_), .B0(new_new_n216_), .B1(new_new_n388_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n313_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n113_), .B(new_new_n23_), .Y(new_new_n392_));
  INV        g370(.A(new_new_n391_), .Y(new_new_n393_));
  NO2        g371(.A(new_new_n356_), .B(new_new_n271_), .Y(new_new_n394_));
  INV        g372(.A(new_new_n229_), .Y(new_new_n395_));
  NO2        g373(.A(i_12_), .B(new_new_n83_), .Y(new_new_n396_));
  NA3        g374(.A(new_new_n396_), .B(new_new_n216_), .C(new_new_n380_), .Y(new_new_n397_));
  NA3        g375(.A(new_new_n277_), .B(new_new_n220_), .C(new_new_n178_), .Y(new_new_n398_));
  AOI210     g376(.A0(new_new_n398_), .A1(new_new_n397_), .B0(new_new_n395_), .Y(new_new_n399_));
  OR2        g377(.A(i_2_), .B(i_5_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n267_), .B(new_new_n192_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n401_), .B(new_new_n345_), .Y(new_new_n402_));
  NO3        g380(.A(new_new_n402_), .B(new_new_n399_), .C(new_new_n394_), .Y(new_new_n403_));
  NA3        g381(.A(new_new_n403_), .B(new_new_n393_), .C(new_new_n383_), .Y(new_new_n404_));
  NO4        g382(.A(new_new_n404_), .B(new_new_n375_), .C(new_new_n366_), .D(new_new_n351_), .Y(new_new_n405_));
  NA4        g383(.A(new_new_n405_), .B(new_new_n305_), .C(new_new_n247_), .D(new_new_n227_), .Y(ori7));
  NO2        g384(.A(new_new_n92_), .B(new_new_n54_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n106_), .B(new_new_n89_), .Y(new_new_n408_));
  NA2        g386(.A(i_3_), .B(new_new_n408_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n336_), .B(new_new_n81_), .Y(new_new_n410_));
  NA2        g388(.A(i_11_), .B(new_new_n161_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n140_), .B(new_new_n411_), .Y(new_new_n412_));
  OAI210     g390(.A0(new_new_n412_), .A1(new_new_n410_), .B0(new_new_n409_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n187_), .B(i_4_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n414_), .B(i_8_), .Y(new_new_n415_));
  NA2        g393(.A(i_2_), .B(new_new_n83_), .Y(new_new_n416_));
  OAI210     g394(.A0(new_new_n86_), .A1(new_new_n165_), .B0(new_new_n166_), .Y(new_new_n417_));
  NO2        g395(.A(i_7_), .B(new_new_n37_), .Y(new_new_n418_));
  NA2        g396(.A(i_4_), .B(i_8_), .Y(new_new_n419_));
  AOI210     g397(.A0(new_new_n419_), .A1(new_new_n224_), .B0(new_new_n418_), .Y(new_new_n420_));
  OAI220     g398(.A0(new_new_n420_), .A1(new_new_n416_), .B0(new_new_n417_), .B1(i_13_), .Y(new_new_n421_));
  NO3        g399(.A(new_new_n421_), .B(new_new_n413_), .C(new_new_n407_), .Y(new_new_n422_));
  AOI210     g400(.A0(new_new_n127_), .A1(new_new_n59_), .B0(i_10_), .Y(new_new_n423_));
  AOI210     g401(.A0(new_new_n423_), .A1(new_new_n187_), .B0(new_new_n148_), .Y(new_new_n424_));
  OR2        g402(.A(i_6_), .B(i_10_), .Y(new_new_n425_));
  OR3        g403(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n426_));
  INV        g404(.A(new_new_n164_), .Y(new_new_n427_));
  OR2        g405(.A(new_new_n424_), .B(new_new_n209_), .Y(new_new_n428_));
  AOI210     g406(.A0(new_new_n428_), .A1(new_new_n422_), .B0(new_new_n60_), .Y(new_new_n429_));
  NOi21      g407(.An(i_11_), .B(i_7_), .Y(new_new_n430_));
  AO210      g408(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n431_), .B(new_new_n430_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n432_), .B(new_new_n170_), .Y(new_new_n433_));
  NA3        g411(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n434_));
  NAi31      g412(.An(new_new_n434_), .B(new_new_n176_), .C(i_11_), .Y(new_new_n435_));
  AOI210     g413(.A0(new_new_n435_), .A1(new_new_n433_), .B0(new_new_n60_), .Y(new_new_n436_));
  NA2        g414(.A(new_new_n85_), .B(new_new_n60_), .Y(new_new_n437_));
  AO210      g415(.A0(new_new_n437_), .A1(new_new_n271_), .B0(new_new_n41_), .Y(new_new_n438_));
  NO3        g416(.A(new_new_n202_), .B(new_new_n171_), .C(new_new_n411_), .Y(new_new_n439_));
  OAI210     g417(.A0(new_new_n439_), .A1(new_new_n184_), .B0(new_new_n60_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n290_), .B(new_new_n31_), .Y(new_new_n441_));
  OR2        g419(.A(new_new_n171_), .B(new_new_n106_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n442_), .B(new_new_n441_), .Y(new_new_n443_));
  NO2        g421(.A(i_1_), .B(i_4_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n444_), .B(new_new_n443_), .Y(new_new_n445_));
  NO2        g423(.A(i_1_), .B(i_12_), .Y(new_new_n446_));
  NA3        g424(.A(new_new_n446_), .B(new_new_n108_), .C(new_new_n24_), .Y(new_new_n447_));
  BUFFER     g425(.A(new_new_n447_), .Y(new_new_n448_));
  NA4        g426(.A(new_new_n448_), .B(new_new_n445_), .C(new_new_n440_), .D(new_new_n438_), .Y(new_new_n449_));
  OAI210     g427(.A0(new_new_n449_), .A1(new_new_n436_), .B0(i_6_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n434_), .B(new_new_n106_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n451_), .B(new_new_n396_), .Y(new_new_n452_));
  NO2        g430(.A(i_6_), .B(i_11_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n452_), .B(new_new_n316_), .Y(new_new_n454_));
  NO3        g432(.A(new_new_n425_), .B(new_new_n186_), .C(new_new_n23_), .Y(new_new_n455_));
  AOI210     g433(.A0(i_1_), .A1(new_new_n203_), .B0(new_new_n455_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n456_), .B(new_new_n44_), .Y(new_new_n457_));
  NA3        g435(.A(new_new_n368_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n458_));
  INV        g436(.A(i_2_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n137_), .B(i_9_), .Y(new_new_n460_));
  NA3        g438(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n461_));
  NO2        g439(.A(new_new_n46_), .B(i_1_), .Y(new_new_n462_));
  NA3        g440(.A(new_new_n462_), .B(new_new_n208_), .C(new_new_n44_), .Y(new_new_n463_));
  OAI220     g441(.A0(new_new_n463_), .A1(new_new_n461_), .B0(new_new_n460_), .B1(new_new_n459_), .Y(new_new_n464_));
  AOI210     g442(.A0(new_new_n332_), .A1(new_new_n295_), .B0(new_new_n190_), .Y(new_new_n465_));
  NO2        g443(.A(new_new_n465_), .B(new_new_n416_), .Y(new_new_n466_));
  NAi21      g444(.An(new_new_n458_), .B(new_new_n91_), .Y(new_new_n467_));
  NO2        g445(.A(i_11_), .B(new_new_n37_), .Y(new_new_n468_));
  INV        g446(.A(new_new_n467_), .Y(new_new_n469_));
  OR3        g447(.A(new_new_n469_), .B(new_new_n466_), .C(new_new_n464_), .Y(new_new_n470_));
  NO3        g448(.A(new_new_n470_), .B(new_new_n457_), .C(new_new_n454_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n187_), .B(new_new_n99_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n430_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n473_), .B(i_1_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n474_), .B(new_new_n426_), .Y(new_new_n475_));
  NA2        g453(.A(new_new_n475_), .B(new_new_n46_), .Y(new_new_n476_));
  NA2        g454(.A(i_3_), .B(new_new_n161_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n477_), .B(new_new_n113_), .Y(new_new_n478_));
  AN2        g456(.A(new_new_n478_), .B(new_new_n370_), .Y(new_new_n479_));
  NO2        g457(.A(new_new_n116_), .B(new_new_n37_), .Y(new_new_n480_));
  NA2        g458(.A(i_1_), .B(i_3_), .Y(new_new_n481_));
  NO2        g459(.A(new_new_n317_), .B(new_new_n92_), .Y(new_new_n482_));
  INV        g460(.A(new_new_n482_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n483_), .B(new_new_n481_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n484_), .B(new_new_n479_), .Y(new_new_n485_));
  NA4        g463(.A(new_new_n485_), .B(new_new_n476_), .C(new_new_n471_), .D(new_new_n450_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n266_), .B(new_new_n265_), .Y(new_new_n487_));
  NO3        g465(.A(new_new_n334_), .B(new_new_n419_), .C(new_new_n83_), .Y(new_new_n488_));
  NA2        g466(.A(new_new_n488_), .B(new_new_n25_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n489_), .B(new_new_n487_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n490_), .B(i_1_), .Y(new_new_n491_));
  AOI210     g469(.A0(new_new_n208_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n492_));
  NO2        g470(.A(new_new_n264_), .B(i_2_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n493_), .B(new_new_n492_), .Y(new_new_n494_));
  AOI210     g472(.A0(new_new_n494_), .A1(new_new_n491_), .B0(i_13_), .Y(new_new_n495_));
  OR2        g473(.A(i_11_), .B(i_7_), .Y(new_new_n496_));
  NA3        g474(.A(new_new_n496_), .B(new_new_n104_), .C(new_new_n137_), .Y(new_new_n497_));
  AOI220     g475(.A0(new_new_n329_), .A1(new_new_n148_), .B0(new_new_n310_), .B1(new_new_n137_), .Y(new_new_n498_));
  OAI210     g476(.A0(new_new_n498_), .A1(new_new_n44_), .B0(new_new_n497_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n54_), .B(i_12_), .Y(new_new_n500_));
  NO2        g478(.A(new_new_n334_), .B(new_new_n24_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n752_), .B(new_new_n92_), .Y(new_new_n502_));
  AOI210     g480(.A0(new_new_n499_), .A1(new_new_n236_), .B0(new_new_n502_), .Y(new_new_n503_));
  INV        g481(.A(new_new_n113_), .Y(new_new_n504_));
  AOI220     g482(.A0(new_new_n504_), .A1(new_new_n69_), .B0(new_new_n277_), .B1(new_new_n462_), .Y(new_new_n505_));
  NO2        g483(.A(new_new_n505_), .B(new_new_n191_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n126_), .B(i_13_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n461_), .B(new_new_n113_), .Y(new_new_n508_));
  INV        g486(.A(new_new_n508_), .Y(new_new_n509_));
  OAI220     g487(.A0(new_new_n509_), .A1(new_new_n68_), .B0(new_new_n507_), .B1(new_new_n492_), .Y(new_new_n510_));
  NO3        g488(.A(new_new_n68_), .B(new_new_n32_), .C(new_new_n99_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n26_), .B(new_new_n161_), .Y(new_new_n512_));
  NA2        g490(.A(new_new_n512_), .B(i_7_), .Y(new_new_n513_));
  NO3        g491(.A(new_new_n334_), .B(new_new_n187_), .C(new_new_n83_), .Y(new_new_n514_));
  AOI210     g492(.A0(new_new_n514_), .A1(new_new_n513_), .B0(new_new_n511_), .Y(new_new_n515_));
  AOI220     g493(.A0(new_new_n277_), .A1(new_new_n462_), .B0(new_new_n91_), .B1(new_new_n100_), .Y(new_new_n516_));
  OAI220     g494(.A0(new_new_n516_), .A1(new_new_n415_), .B0(new_new_n515_), .B1(new_new_n427_), .Y(new_new_n517_));
  NO3        g495(.A(new_new_n517_), .B(new_new_n510_), .C(new_new_n506_), .Y(new_new_n518_));
  OR2        g496(.A(i_11_), .B(i_6_), .Y(new_new_n519_));
  NA3        g497(.A(new_new_n414_), .B(new_new_n512_), .C(i_7_), .Y(new_new_n520_));
  AOI210     g498(.A0(new_new_n520_), .A1(new_new_n509_), .B0(new_new_n519_), .Y(new_new_n521_));
  NA3        g499(.A(new_new_n290_), .B(new_new_n418_), .C(new_new_n97_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n453_), .B(i_13_), .Y(new_new_n523_));
  NAi21      g501(.An(i_11_), .B(i_12_), .Y(new_new_n524_));
  NO3        g502(.A(new_new_n334_), .B(new_new_n396_), .C(new_new_n419_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n525_), .B(new_new_n228_), .Y(new_new_n526_));
  NA3        g504(.A(new_new_n526_), .B(new_new_n523_), .C(new_new_n522_), .Y(new_new_n527_));
  OAI210     g505(.A0(new_new_n527_), .A1(new_new_n521_), .B0(new_new_n60_), .Y(new_new_n528_));
  NO2        g506(.A(i_2_), .B(i_12_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n263_), .B(new_new_n529_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n127_), .B(i_2_), .Y(new_new_n531_));
  NA2        g509(.A(new_new_n531_), .B(new_new_n446_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n532_), .B(new_new_n530_), .Y(new_new_n533_));
  NA3        g511(.A(new_new_n533_), .B(new_new_n45_), .C(new_new_n183_), .Y(new_new_n534_));
  NA4        g512(.A(new_new_n534_), .B(new_new_n528_), .C(new_new_n518_), .D(new_new_n503_), .Y(new_new_n535_));
  OR4        g513(.A(new_new_n535_), .B(new_new_n495_), .C(new_new_n486_), .D(new_new_n429_), .Y(ori5));
  NA2        g514(.A(new_new_n473_), .B(new_new_n211_), .Y(new_new_n537_));
  AN2        g515(.A(new_new_n24_), .B(i_10_), .Y(new_new_n538_));
  NA3        g516(.A(new_new_n538_), .B(new_new_n529_), .C(new_new_n106_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n415_), .B(i_11_), .Y(new_new_n540_));
  NA2        g518(.A(new_new_n86_), .B(new_new_n540_), .Y(new_new_n541_));
  NA3        g519(.A(new_new_n541_), .B(new_new_n539_), .C(new_new_n537_), .Y(new_new_n542_));
  NO3        g520(.A(i_11_), .B(new_new_n187_), .C(i_13_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n123_), .B(new_new_n23_), .Y(new_new_n544_));
  NA2        g522(.A(i_12_), .B(i_8_), .Y(new_new_n545_));
  OAI210     g523(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n545_), .Y(new_new_n546_));
  INV        g524(.A(new_new_n307_), .Y(new_new_n547_));
  AOI220     g525(.A0(new_new_n229_), .A1(new_new_n392_), .B0(new_new_n546_), .B1(new_new_n544_), .Y(new_new_n548_));
  INV        g526(.A(new_new_n548_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n549_), .B(new_new_n542_), .Y(new_new_n550_));
  INV        g528(.A(new_new_n151_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n193_), .Y(new_new_n552_));
  OAI210     g530(.A0(new_new_n493_), .A1(new_new_n309_), .B0(new_new_n109_), .Y(new_new_n553_));
  AOI210     g531(.A0(new_new_n553_), .A1(new_new_n552_), .B0(new_new_n551_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n317_), .B(new_new_n26_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n555_), .B(new_new_n295_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n556_), .B(i_2_), .Y(new_new_n557_));
  INV        g535(.A(new_new_n557_), .Y(new_new_n558_));
  AOI210     g536(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n292_), .Y(new_new_n559_));
  AOI210     g537(.A0(new_new_n559_), .A1(new_new_n558_), .B0(new_new_n554_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n160_), .B(new_new_n124_), .Y(new_new_n561_));
  OAI210     g539(.A0(new_new_n561_), .A1(new_new_n544_), .B0(i_2_), .Y(new_new_n562_));
  INV        g540(.A(new_new_n152_), .Y(new_new_n563_));
  NO3        g541(.A(new_new_n431_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n564_));
  AOI210     g542(.A0(new_new_n563_), .A1(new_new_n86_), .B0(new_new_n564_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n565_), .A1(new_new_n562_), .B0(new_new_n161_), .Y(new_new_n566_));
  OA210      g544(.A0(new_new_n432_), .A1(new_new_n125_), .B0(i_13_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n164_), .B(new_new_n165_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n568_), .B(new_new_n267_), .Y(new_new_n569_));
  AOI210     g547(.A0(new_new_n171_), .A1(new_new_n143_), .B0(new_new_n359_), .Y(new_new_n570_));
  NA2        g548(.A(new_new_n570_), .B(new_new_n295_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n100_), .B(new_new_n44_), .Y(new_new_n572_));
  INV        g550(.A(new_new_n223_), .Y(new_new_n573_));
  NA4        g551(.A(new_new_n573_), .B(new_new_n224_), .C(new_new_n123_), .D(new_new_n42_), .Y(new_new_n574_));
  OAI210     g552(.A0(new_new_n574_), .A1(new_new_n572_), .B0(new_new_n571_), .Y(new_new_n575_));
  NO4        g553(.A(new_new_n575_), .B(new_new_n569_), .C(new_new_n567_), .D(new_new_n566_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n392_), .B(new_new_n28_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n543_), .B(new_new_n217_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n578_), .B(new_new_n577_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n59_), .B(i_12_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n580_), .B(new_new_n125_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n581_), .B(new_new_n411_), .Y(new_new_n582_));
  AOI220     g560(.A0(new_new_n582_), .A1(new_new_n36_), .B0(new_new_n579_), .B1(new_new_n46_), .Y(new_new_n583_));
  NA4        g561(.A(new_new_n583_), .B(new_new_n576_), .C(new_new_n560_), .D(new_new_n550_), .Y(ori6));
  NA4        g562(.A(new_new_n278_), .B(new_new_n335_), .C(new_new_n68_), .D(new_new_n99_), .Y(new_new_n585_));
  INV        g563(.A(new_new_n585_), .Y(new_new_n586_));
  NO2        g564(.A(new_new_n179_), .B(new_new_n338_), .Y(new_new_n587_));
  NO2        g565(.A(i_11_), .B(i_9_), .Y(new_new_n588_));
  NO2        g566(.A(new_new_n586_), .B(new_new_n232_), .Y(new_new_n589_));
  OR2        g567(.A(new_new_n589_), .B(i_12_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n396_), .B(new_new_n60_), .Y(new_new_n591_));
  BUFFER     g569(.A(new_new_n437_), .Y(new_new_n592_));
  NA2        g570(.A(new_new_n592_), .B(new_new_n591_), .Y(new_new_n593_));
  INV        g571(.A(new_new_n163_), .Y(new_new_n594_));
  AOI220     g572(.A0(new_new_n594_), .A1(new_new_n588_), .B0(new_new_n593_), .B1(new_new_n70_), .Y(new_new_n595_));
  INV        g573(.A(new_new_n231_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n72_), .B(new_new_n130_), .Y(new_new_n597_));
  INV        g575(.A(new_new_n123_), .Y(new_new_n598_));
  NA2        g576(.A(new_new_n598_), .B(new_new_n46_), .Y(new_new_n599_));
  AOI210     g577(.A0(new_new_n599_), .A1(new_new_n597_), .B0(new_new_n596_), .Y(new_new_n600_));
  NO2        g578(.A(new_new_n196_), .B(i_9_), .Y(new_new_n601_));
  NA2        g579(.A(new_new_n601_), .B(new_new_n580_), .Y(new_new_n602_));
  AOI210     g580(.A0(new_new_n602_), .A1(new_new_n357_), .B0(new_new_n157_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n32_), .B(i_11_), .Y(new_new_n604_));
  NAi32      g582(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n605_));
  NO2        g583(.A(new_new_n519_), .B(new_new_n605_), .Y(new_new_n606_));
  OR3        g584(.A(new_new_n606_), .B(new_new_n603_), .C(new_new_n600_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n496_), .B(i_2_), .Y(new_new_n608_));
  OR2        g586(.A(new_new_n432_), .B(new_new_n309_), .Y(new_new_n609_));
  NA3        g587(.A(new_new_n609_), .B(new_new_n142_), .C(new_new_n66_), .Y(new_new_n610_));
  OR2        g588(.A(new_new_n547_), .B(new_new_n36_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n611_), .B(new_new_n610_), .Y(new_new_n612_));
  OAI210     g590(.A0(i_6_), .A1(i_11_), .B0(new_new_n84_), .Y(new_new_n613_));
  AOI220     g591(.A0(new_new_n613_), .A1(new_new_n385_), .B0(new_new_n587_), .B1(new_new_n513_), .Y(new_new_n614_));
  NA3        g592(.A(new_new_n267_), .B(new_new_n188_), .C(new_new_n142_), .Y(new_new_n615_));
  NA2        g593(.A(new_new_n280_), .B(new_new_n67_), .Y(new_new_n616_));
  NA4        g594(.A(new_new_n616_), .B(new_new_n615_), .C(new_new_n614_), .D(new_new_n417_), .Y(new_new_n617_));
  AO210      g595(.A0(new_new_n359_), .A1(new_new_n46_), .B0(new_new_n85_), .Y(new_new_n618_));
  NA3        g596(.A(new_new_n618_), .B(new_new_n336_), .C(new_new_n178_), .Y(new_new_n619_));
  AOI210     g597(.A0(new_new_n309_), .A1(new_new_n307_), .B0(new_new_n384_), .Y(new_new_n620_));
  NO2        g598(.A(new_new_n425_), .B(new_new_n100_), .Y(new_new_n621_));
  OAI210     g599(.A0(new_new_n621_), .A1(new_new_n110_), .B0(new_new_n289_), .Y(new_new_n622_));
  NA3        g600(.A(new_new_n622_), .B(new_new_n620_), .C(new_new_n619_), .Y(new_new_n623_));
  NO4        g601(.A(new_new_n623_), .B(new_new_n617_), .C(new_new_n612_), .D(new_new_n607_), .Y(new_new_n624_));
  NA4        g602(.A(new_new_n624_), .B(new_new_n595_), .C(new_new_n590_), .D(new_new_n273_), .Y(ori3));
  NA2        g603(.A(i_12_), .B(i_10_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n615_), .B(new_new_n417_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n627_), .B(new_new_n40_), .Y(new_new_n628_));
  NOi21      g606(.An(new_new_n96_), .B(new_new_n556_), .Y(new_new_n629_));
  NO3        g607(.A(new_new_n442_), .B(new_new_n317_), .C(new_new_n130_), .Y(new_new_n630_));
  NA2        g608(.A(new_new_n290_), .B(new_new_n45_), .Y(new_new_n631_));
  AN2        g609(.A(new_new_n315_), .B(new_new_n55_), .Y(new_new_n632_));
  NO3        g610(.A(new_new_n632_), .B(new_new_n630_), .C(new_new_n629_), .Y(new_new_n633_));
  AOI210     g611(.A0(new_new_n633_), .A1(new_new_n628_), .B0(new_new_n48_), .Y(new_new_n634_));
  NO4        g612(.A(new_new_n269_), .B(new_new_n275_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n635_));
  NA2        g613(.A(new_new_n157_), .B(new_new_n388_), .Y(new_new_n636_));
  NOi21      g614(.An(new_new_n636_), .B(new_new_n635_), .Y(new_new_n637_));
  NO2        g615(.A(new_new_n637_), .B(new_new_n60_), .Y(new_new_n638_));
  NOi21      g616(.An(i_5_), .B(i_9_), .Y(new_new_n639_));
  NA2        g617(.A(new_new_n639_), .B(new_new_n306_), .Y(new_new_n640_));
  BUFFER     g618(.A(new_new_n208_), .Y(new_new_n641_));
  AOI210     g619(.A0(new_new_n641_), .A1(new_new_n332_), .B0(new_new_n488_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n642_), .B(new_new_n640_), .Y(new_new_n643_));
  NO3        g621(.A(new_new_n643_), .B(new_new_n638_), .C(new_new_n634_), .Y(new_new_n644_));
  NA2        g622(.A(new_new_n157_), .B(new_new_n24_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n480_), .B(new_new_n408_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n646_), .B(new_new_n645_), .Y(new_new_n647_));
  INV        g625(.A(new_new_n647_), .Y(new_new_n648_));
  NA2        g626(.A(new_new_n389_), .B(i_0_), .Y(new_new_n649_));
  NO3        g627(.A(new_new_n649_), .B(new_new_n276_), .C(new_new_n86_), .Y(new_new_n650_));
  NO4        g628(.A(new_new_n400_), .B(new_new_n176_), .C(new_new_n292_), .D(i_6_), .Y(new_new_n651_));
  AOI210     g629(.A0(new_new_n651_), .A1(i_11_), .B0(new_new_n650_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n543_), .B(new_new_n232_), .Y(new_new_n653_));
  AOI210     g631(.A0(new_new_n336_), .A1(new_new_n86_), .B0(new_new_n57_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n654_), .B(new_new_n653_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n198_), .B(new_new_n145_), .Y(new_new_n656_));
  NA2        g634(.A(i_0_), .B(i_10_), .Y(new_new_n657_));
  INV        g635(.A(new_new_n369_), .Y(new_new_n658_));
  NO4        g636(.A(new_new_n113_), .B(new_new_n57_), .C(new_new_n477_), .D(i_5_), .Y(new_new_n659_));
  AO220      g637(.A0(new_new_n659_), .A1(new_new_n658_), .B0(new_new_n656_), .B1(i_6_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n660_), .B(new_new_n655_), .Y(new_new_n661_));
  NA3        g639(.A(new_new_n661_), .B(new_new_n652_), .C(new_new_n648_), .Y(new_new_n662_));
  NO2        g640(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n663_));
  NA2        g641(.A(i_11_), .B(i_9_), .Y(new_new_n664_));
  NO3        g642(.A(i_12_), .B(new_new_n664_), .C(new_new_n416_), .Y(new_new_n665_));
  AN2        g643(.A(new_new_n665_), .B(new_new_n663_), .Y(new_new_n666_));
  NA2        g644(.A(new_new_n279_), .B(new_new_n156_), .Y(new_new_n667_));
  INV        g645(.A(new_new_n667_), .Y(new_new_n668_));
  NO2        g646(.A(new_new_n664_), .B(new_new_n70_), .Y(new_new_n669_));
  NO2        g647(.A(new_new_n668_), .B(new_new_n666_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n468_), .B(new_new_n120_), .Y(new_new_n671_));
  NO2        g649(.A(i_6_), .B(new_new_n671_), .Y(new_new_n672_));
  NA2        g650(.A(new_new_n151_), .B(new_new_n101_), .Y(new_new_n673_));
  NA2        g651(.A(new_new_n418_), .B(new_new_n232_), .Y(new_new_n674_));
  NO2        g652(.A(new_new_n674_), .B(new_new_n631_), .Y(new_new_n675_));
  NO2        g653(.A(new_new_n675_), .B(new_new_n672_), .Y(new_new_n676_));
  INV        g654(.A(new_new_n230_), .Y(new_new_n677_));
  NA2        g655(.A(new_new_n676_), .B(new_new_n670_), .Y(new_new_n678_));
  NO2        g656(.A(new_new_n626_), .B(new_new_n229_), .Y(new_new_n679_));
  OA210      g657(.A0(new_new_n331_), .A1(new_new_n182_), .B0(new_new_n330_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n679_), .B(new_new_n669_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n669_), .B(new_new_n224_), .Y(new_new_n682_));
  INV        g660(.A(new_new_n682_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n683_), .B(new_new_n331_), .Y(new_new_n684_));
  NO3        g662(.A(new_new_n400_), .B(new_new_n250_), .C(new_new_n24_), .Y(new_new_n685_));
  AOI210     g663(.A0(new_new_n501_), .A1(new_new_n372_), .B0(new_new_n685_), .Y(new_new_n686_));
  NAi21      g664(.An(i_9_), .B(i_5_), .Y(new_new_n687_));
  NO2        g665(.A(new_new_n687_), .B(new_new_n285_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n688_), .B(new_new_n432_), .Y(new_new_n689_));
  OAI220     g667(.A0(new_new_n689_), .A1(new_new_n83_), .B0(new_new_n686_), .B1(new_new_n152_), .Y(new_new_n690_));
  NO2        g668(.A(new_new_n690_), .B(new_new_n361_), .Y(new_new_n691_));
  NA3        g669(.A(new_new_n691_), .B(new_new_n684_), .C(new_new_n681_), .Y(new_new_n692_));
  NO3        g670(.A(new_new_n692_), .B(new_new_n678_), .C(new_new_n662_), .Y(new_new_n693_));
  NO2        g671(.A(i_0_), .B(new_new_n524_), .Y(new_new_n694_));
  AOI210     g672(.A0(new_new_n591_), .A1(new_new_n487_), .B0(new_new_n673_), .Y(new_new_n695_));
  INV        g673(.A(new_new_n695_), .Y(new_new_n696_));
  NA2        g674(.A(new_new_n192_), .B(new_new_n185_), .Y(new_new_n697_));
  AOI210     g675(.A0(new_new_n697_), .A1(new_new_n649_), .B0(new_new_n145_), .Y(new_new_n698_));
  INV        g676(.A(new_new_n698_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n699_), .B(new_new_n696_), .Y(new_new_n700_));
  NO3        g678(.A(new_new_n657_), .B(new_new_n639_), .C(new_new_n160_), .Y(new_new_n701_));
  AOI220     g679(.A0(new_new_n701_), .A1(i_11_), .B0(new_new_n387_), .B1(new_new_n72_), .Y(new_new_n702_));
  NO3        g680(.A(new_new_n172_), .B(new_new_n275_), .C(i_0_), .Y(new_new_n703_));
  OAI210     g681(.A0(new_new_n703_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n704_), .B(new_new_n702_), .Y(new_new_n705_));
  INV        g683(.A(new_new_n92_), .Y(new_new_n706_));
  AOI210     g684(.A0(new_new_n706_), .A1(new_new_n694_), .B0(new_new_n107_), .Y(new_new_n707_));
  OR2        g685(.A(new_new_n707_), .B(i_5_), .Y(new_new_n708_));
  AOI210     g686(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n154_), .Y(new_new_n709_));
  NA2        g687(.A(new_new_n709_), .B(new_new_n680_), .Y(new_new_n710_));
  NO3        g688(.A(new_new_n631_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n344_), .B(new_new_n337_), .Y(new_new_n712_));
  NO3        g690(.A(new_new_n712_), .B(new_new_n711_), .C(new_new_n753_), .Y(new_new_n713_));
  NA3        g691(.A(new_new_n278_), .B(new_new_n151_), .C(new_new_n150_), .Y(new_new_n714_));
  NA3        g692(.A(i_5_), .B(new_new_n221_), .C(new_new_n185_), .Y(new_new_n715_));
  NA2        g693(.A(new_new_n715_), .B(new_new_n714_), .Y(new_new_n716_));
  NO3        g694(.A(new_new_n664_), .B(new_new_n178_), .C(new_new_n160_), .Y(new_new_n717_));
  NO2        g695(.A(new_new_n717_), .B(new_new_n716_), .Y(new_new_n718_));
  NA4        g696(.A(new_new_n718_), .B(new_new_n713_), .C(new_new_n710_), .D(new_new_n708_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n586_), .B(new_new_n155_), .Y(new_new_n720_));
  INV        g698(.A(new_new_n720_), .Y(new_new_n721_));
  NO4        g699(.A(new_new_n721_), .B(new_new_n719_), .C(new_new_n705_), .D(new_new_n700_), .Y(new_new_n722_));
  OAI210     g700(.A0(new_new_n608_), .A1(new_new_n604_), .B0(new_new_n37_), .Y(new_new_n723_));
  NA2        g701(.A(new_new_n723_), .B(new_new_n424_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n724_), .B(new_new_n170_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n158_), .B(new_new_n159_), .Y(new_new_n726_));
  AO210      g704(.A0(new_new_n496_), .A1(new_new_n33_), .B0(new_new_n726_), .Y(new_new_n727_));
  NAi31      g705(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n728_));
  AOI210     g706(.A0(new_new_n116_), .A1(new_new_n67_), .B0(new_new_n728_), .Y(new_new_n729_));
  NO2        g707(.A(new_new_n729_), .B(new_new_n455_), .Y(new_new_n730_));
  NA2        g708(.A(new_new_n730_), .B(new_new_n727_), .Y(new_new_n731_));
  NO2        g709(.A(new_new_n323_), .B(new_new_n208_), .Y(new_new_n732_));
  AOI210     g710(.A0(new_new_n731_), .A1(new_new_n48_), .B0(new_new_n732_), .Y(new_new_n733_));
  AOI210     g711(.A0(new_new_n733_), .A1(new_new_n725_), .B0(new_new_n70_), .Y(new_new_n734_));
  INV        g712(.A(new_new_n272_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n735_), .B(new_new_n551_), .Y(new_new_n736_));
  NA3        g714(.A(new_new_n555_), .B(new_new_n221_), .C(new_new_n77_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n737_), .B(i_11_), .Y(new_new_n738_));
  NO3        g716(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n739_));
  OAI210     g717(.A0(new_new_n677_), .A1(new_new_n225_), .B0(new_new_n739_), .Y(new_new_n740_));
  NO2        g718(.A(new_new_n740_), .B(new_new_n524_), .Y(new_new_n741_));
  NO4        g719(.A(new_new_n687_), .B(new_new_n333_), .C(new_new_n197_), .D(new_new_n196_), .Y(new_new_n742_));
  NO2        g720(.A(new_new_n742_), .B(new_new_n384_), .Y(new_new_n743_));
  INV        g721(.A(new_new_n256_), .Y(new_new_n744_));
  AOI210     g722(.A0(new_new_n744_), .A1(new_new_n743_), .B0(new_new_n41_), .Y(new_new_n745_));
  NO3        g723(.A(new_new_n745_), .B(new_new_n741_), .C(new_new_n738_), .Y(new_new_n746_));
  INV        g724(.A(new_new_n746_), .Y(new_new_n747_));
  NO3        g725(.A(new_new_n747_), .B(new_new_n736_), .C(new_new_n734_), .Y(new_new_n748_));
  NA4        g726(.A(new_new_n748_), .B(new_new_n722_), .C(new_new_n693_), .D(new_new_n644_), .Y(ori4));
  INV        g727(.A(new_new_n500_), .Y(new_new_n752_));
  INV        g728(.A(new_new_n371_), .Y(new_new_n753_));
  INV        g729(.A(i_6_), .Y(new_new_n754_));
endmodule


