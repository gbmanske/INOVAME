//Benchmark atmr_9sym_175_0.0156

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  NA2        o002(.A(i_4_), .B(ori_ori_n12_), .Y(ori_ori_n13_));
  INV        o003(.A(i_5_), .Y(ori_ori_n14_));
  NOi21      o004(.An(i_3_), .B(i_7_), .Y(ori_ori_n15_));
  NA3        o005(.A(ori_ori_n15_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n16_));
  INV        o006(.A(i_0_), .Y(ori_ori_n17_));
  NOi21      o007(.An(i_1_), .B(i_3_), .Y(ori_ori_n18_));
  NA3        o008(.A(ori_ori_n18_), .B(ori_ori_n17_), .C(i_2_), .Y(ori_ori_n19_));
  AOI210     o009(.A0(ori_ori_n19_), .A1(ori_ori_n16_), .B0(ori_ori_n13_), .Y(ori_ori_n20_));
  INV        o010(.A(i_4_), .Y(ori_ori_n21_));
  NA2        o011(.A(i_0_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  INV        o012(.A(i_7_), .Y(ori_ori_n23_));
  NA3        o013(.A(i_6_), .B(i_5_), .C(ori_ori_n23_), .Y(ori_ori_n24_));
  NOi21      o014(.An(i_8_), .B(i_6_), .Y(ori_ori_n25_));
  NOi21      o015(.An(i_1_), .B(i_8_), .Y(ori_ori_n26_));
  AOI220     o016(.A0(ori_ori_n26_), .A1(i_2_), .B0(ori_ori_n25_), .B1(i_5_), .Y(ori_ori_n27_));
  AOI210     o017(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n22_), .Y(ori_ori_n28_));
  AOI210     o018(.A0(ori_ori_n28_), .A1(ori_ori_n11_), .B0(ori_ori_n20_), .Y(ori_ori_n29_));
  NA2        o019(.A(i_0_), .B(ori_ori_n14_), .Y(ori_ori_n30_));
  NA2        o020(.A(ori_ori_n17_), .B(i_5_), .Y(ori_ori_n31_));
  NO2        o021(.A(i_2_), .B(i_4_), .Y(ori_ori_n32_));
  NA3        o022(.A(ori_ori_n32_), .B(i_6_), .C(i_8_), .Y(ori_ori_n33_));
  AOI210     o023(.A0(ori_ori_n31_), .A1(ori_ori_n30_), .B0(ori_ori_n33_), .Y(ori_ori_n34_));
  INV        o024(.A(i_2_), .Y(ori_ori_n35_));
  NOi21      o025(.An(i_5_), .B(i_0_), .Y(ori_ori_n36_));
  NOi21      o026(.An(i_6_), .B(i_8_), .Y(ori_ori_n37_));
  NOi21      o027(.An(i_7_), .B(i_1_), .Y(ori_ori_n38_));
  NOi21      o028(.An(i_5_), .B(i_6_), .Y(ori_ori_n39_));
  AOI220     o029(.A0(ori_ori_n39_), .A1(ori_ori_n38_), .B0(ori_ori_n37_), .B1(ori_ori_n36_), .Y(ori_ori_n40_));
  NO3        o030(.A(ori_ori_n40_), .B(ori_ori_n35_), .C(i_4_), .Y(ori_ori_n41_));
  NOi21      o031(.An(i_0_), .B(i_4_), .Y(ori_ori_n42_));
  XO2        o032(.A(i_1_), .B(i_3_), .Y(ori_ori_n43_));
  NOi21      o033(.An(i_7_), .B(i_5_), .Y(ori_ori_n44_));
  AN3        o034(.A(ori_ori_n44_), .B(ori_ori_n43_), .C(ori_ori_n42_), .Y(ori_ori_n45_));
  INV        o035(.A(i_1_), .Y(ori_ori_n46_));
  NOi21      o036(.An(i_3_), .B(i_0_), .Y(ori_ori_n47_));
  NA2        o037(.A(ori_ori_n47_), .B(ori_ori_n46_), .Y(ori_ori_n48_));
  NA3        o038(.A(i_6_), .B(ori_ori_n14_), .C(i_7_), .Y(ori_ori_n49_));
  AOI210     o039(.A0(ori_ori_n49_), .A1(ori_ori_n24_), .B0(ori_ori_n48_), .Y(ori_ori_n50_));
  NO4        o040(.A(ori_ori_n50_), .B(ori_ori_n45_), .C(ori_ori_n41_), .D(ori_ori_n34_), .Y(ori_ori_n51_));
  INV        o041(.A(i_8_), .Y(ori_ori_n52_));
  NA2        o042(.A(i_1_), .B(ori_ori_n11_), .Y(ori_ori_n53_));
  NOi21      o043(.An(i_4_), .B(i_0_), .Y(ori_ori_n54_));
  NO2        o044(.A(ori_ori_n25_), .B(ori_ori_n15_), .Y(ori_ori_n55_));
  NA2        o045(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n56_));
  NOi21      o046(.An(i_2_), .B(i_8_), .Y(ori_ori_n57_));
  NO3        o047(.A(ori_ori_n57_), .B(ori_ori_n54_), .C(ori_ori_n42_), .Y(ori_ori_n58_));
  NO3        o048(.A(ori_ori_n58_), .B(ori_ori_n56_), .C(ori_ori_n55_), .Y(ori_ori_n59_));
  INV        o049(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  NOi31      o050(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n61_));
  NA2        o051(.A(ori_ori_n61_), .B(i_0_), .Y(ori_ori_n62_));
  NOi21      o052(.An(i_4_), .B(i_3_), .Y(ori_ori_n63_));
  NOi21      o053(.An(i_1_), .B(i_4_), .Y(ori_ori_n64_));
  OAI210     o054(.A0(ori_ori_n64_), .A1(ori_ori_n63_), .B0(ori_ori_n57_), .Y(ori_ori_n65_));
  NA2        o055(.A(ori_ori_n65_), .B(ori_ori_n62_), .Y(ori_ori_n66_));
  AN2        o056(.A(i_8_), .B(i_7_), .Y(ori_ori_n67_));
  NA2        o057(.A(ori_ori_n67_), .B(ori_ori_n12_), .Y(ori_ori_n68_));
  NOi21      o058(.An(i_8_), .B(i_7_), .Y(ori_ori_n69_));
  NA3        o059(.A(ori_ori_n69_), .B(ori_ori_n63_), .C(i_6_), .Y(ori_ori_n70_));
  OAI210     o060(.A0(ori_ori_n68_), .A1(ori_ori_n56_), .B0(ori_ori_n70_), .Y(ori_ori_n71_));
  AOI220     o061(.A0(ori_ori_n71_), .A1(ori_ori_n35_), .B0(ori_ori_n66_), .B1(ori_ori_n39_), .Y(ori_ori_n72_));
  NA4        o062(.A(ori_ori_n72_), .B(ori_ori_n60_), .C(ori_ori_n51_), .D(ori_ori_n29_), .Y(ori_ori_n73_));
  NA2        o063(.A(i_8_), .B(i_7_), .Y(ori_ori_n74_));
  NA2        o064(.A(i_8_), .B(ori_ori_n23_), .Y(ori_ori_n75_));
  AOI220     o065(.A0(ori_ori_n47_), .A1(i_1_), .B0(ori_ori_n43_), .B1(i_2_), .Y(ori_ori_n76_));
  NOi21      o066(.An(i_1_), .B(i_2_), .Y(ori_ori_n77_));
  NA3        o067(.A(ori_ori_n77_), .B(ori_ori_n54_), .C(i_6_), .Y(ori_ori_n78_));
  OAI210     o068(.A0(ori_ori_n76_), .A1(ori_ori_n75_), .B0(ori_ori_n78_), .Y(ori_ori_n79_));
  NA2        o069(.A(ori_ori_n79_), .B(ori_ori_n14_), .Y(ori_ori_n80_));
  NA3        o070(.A(ori_ori_n69_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n81_));
  NA3        o071(.A(ori_ori_n26_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n82_));
  NA2        o072(.A(ori_ori_n82_), .B(ori_ori_n81_), .Y(ori_ori_n83_));
  NOi32      o073(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(ori_ori_n84_));
  NA2        o074(.A(ori_ori_n84_), .B(i_3_), .Y(ori_ori_n85_));
  NA3        o075(.A(ori_ori_n18_), .B(i_2_), .C(i_6_), .Y(ori_ori_n86_));
  NA2        o076(.A(ori_ori_n86_), .B(ori_ori_n85_), .Y(ori_ori_n87_));
  NO2        o077(.A(i_0_), .B(i_4_), .Y(ori_ori_n88_));
  AOI220     o078(.A0(ori_ori_n88_), .A1(ori_ori_n87_), .B0(ori_ori_n83_), .B1(ori_ori_n63_), .Y(ori_ori_n89_));
  NA2        o079(.A(ori_ori_n89_), .B(ori_ori_n80_), .Y(ori_ori_n90_));
  NAi21      o080(.An(i_3_), .B(i_6_), .Y(ori_ori_n91_));
  NO2        o081(.A(ori_ori_n91_), .B(ori_ori_n52_), .Y(ori_ori_n92_));
  NA2        o082(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n93_));
  NOi21      o083(.An(i_7_), .B(i_8_), .Y(ori_ori_n94_));
  NOi31      o084(.An(i_6_), .B(i_5_), .C(i_7_), .Y(ori_ori_n95_));
  AOI210     o085(.A0(ori_ori_n94_), .A1(ori_ori_n12_), .B0(ori_ori_n95_), .Y(ori_ori_n96_));
  OAI210     o086(.A0(ori_ori_n96_), .A1(ori_ori_n11_), .B0(ori_ori_n93_), .Y(ori_ori_n97_));
  OAI210     o087(.A0(ori_ori_n97_), .A1(ori_ori_n92_), .B0(ori_ori_n77_), .Y(ori_ori_n98_));
  NA3        o088(.A(ori_ori_n25_), .B(i_2_), .C(ori_ori_n14_), .Y(ori_ori_n99_));
  AOI210     o089(.A0(ori_ori_n22_), .A1(ori_ori_n53_), .B0(ori_ori_n99_), .Y(ori_ori_n100_));
  NA2        o090(.A(ori_ori_n47_), .B(ori_ori_n46_), .Y(ori_ori_n101_));
  NA3        o091(.A(ori_ori_n21_), .B(i_5_), .C(i_7_), .Y(ori_ori_n102_));
  OAI210     o092(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(ori_ori_n103_));
  NA3        o093(.A(ori_ori_n74_), .B(ori_ori_n18_), .C(ori_ori_n17_), .Y(ori_ori_n104_));
  OAI220     o094(.A0(ori_ori_n104_), .A1(ori_ori_n103_), .B0(ori_ori_n102_), .B1(ori_ori_n101_), .Y(ori_ori_n105_));
  NO2        o095(.A(ori_ori_n105_), .B(ori_ori_n100_), .Y(ori_ori_n106_));
  NA3        o096(.A(ori_ori_n69_), .B(ori_ori_n35_), .C(i_3_), .Y(ori_ori_n107_));
  NA2        o097(.A(ori_ori_n46_), .B(i_6_), .Y(ori_ori_n108_));
  AOI210     o098(.A0(ori_ori_n108_), .A1(ori_ori_n22_), .B0(ori_ori_n107_), .Y(ori_ori_n109_));
  NAi21      o099(.An(i_6_), .B(i_0_), .Y(ori_ori_n110_));
  NA3        o100(.A(ori_ori_n64_), .B(i_5_), .C(ori_ori_n23_), .Y(ori_ori_n111_));
  NOi21      o101(.An(i_4_), .B(i_6_), .Y(ori_ori_n112_));
  NOi21      o102(.An(i_5_), .B(i_3_), .Y(ori_ori_n113_));
  NA3        o103(.A(ori_ori_n113_), .B(ori_ori_n77_), .C(ori_ori_n112_), .Y(ori_ori_n114_));
  OAI210     o104(.A0(ori_ori_n111_), .A1(ori_ori_n110_), .B0(ori_ori_n114_), .Y(ori_ori_n115_));
  NA2        o105(.A(ori_ori_n77_), .B(ori_ori_n37_), .Y(ori_ori_n116_));
  NOi21      o106(.An(ori_ori_n44_), .B(ori_ori_n116_), .Y(ori_ori_n117_));
  NO3        o107(.A(ori_ori_n117_), .B(ori_ori_n115_), .C(ori_ori_n109_), .Y(ori_ori_n118_));
  NOi21      o108(.An(i_6_), .B(i_1_), .Y(ori_ori_n119_));
  AOI220     o109(.A0(ori_ori_n119_), .A1(i_7_), .B0(ori_ori_n25_), .B1(i_5_), .Y(ori_ori_n120_));
  NOi31      o110(.An(ori_ori_n54_), .B(ori_ori_n120_), .C(i_2_), .Y(ori_ori_n121_));
  NOi21      o111(.An(i_3_), .B(i_1_), .Y(ori_ori_n122_));
  NA2        o112(.A(ori_ori_n122_), .B(i_4_), .Y(ori_ori_n123_));
  AOI210     o113(.A0(i_8_), .A1(i_6_), .B0(ori_ori_n123_), .Y(ori_ori_n124_));
  NA2        o114(.A(ori_ori_n94_), .B(ori_ori_n14_), .Y(ori_ori_n125_));
  NOi31      o115(.An(ori_ori_n47_), .B(ori_ori_n125_), .C(ori_ori_n35_), .Y(ori_ori_n126_));
  NO3        o116(.A(ori_ori_n126_), .B(ori_ori_n124_), .C(ori_ori_n121_), .Y(ori_ori_n127_));
  NA4        o117(.A(ori_ori_n127_), .B(ori_ori_n118_), .C(ori_ori_n106_), .D(ori_ori_n98_), .Y(ori_ori_n128_));
  NA2        o118(.A(ori_ori_n57_), .B(ori_ori_n15_), .Y(ori_ori_n129_));
  NOi31      o119(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n130_));
  NOi31      o120(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n131_));
  OAI210     o121(.A0(ori_ori_n131_), .A1(ori_ori_n130_), .B0(i_7_), .Y(ori_ori_n132_));
  NA3        o122(.A(ori_ori_n37_), .B(i_2_), .C(ori_ori_n14_), .Y(ori_ori_n133_));
  NA4        o123(.A(ori_ori_n133_), .B(ori_ori_n132_), .C(ori_ori_n129_), .D(ori_ori_n116_), .Y(ori_ori_n134_));
  NA2        o124(.A(ori_ori_n134_), .B(ori_ori_n42_), .Y(ori_ori_n135_));
  NA2        o125(.A(ori_ori_n63_), .B(ori_ori_n38_), .Y(ori_ori_n136_));
  AOI210     o126(.A0(ori_ori_n136_), .A1(ori_ori_n81_), .B0(ori_ori_n31_), .Y(ori_ori_n137_));
  NA3        o127(.A(ori_ori_n69_), .B(ori_ori_n61_), .C(i_6_), .Y(ori_ori_n138_));
  INV        o128(.A(ori_ori_n138_), .Y(ori_ori_n139_));
  NOi21      o129(.An(i_0_), .B(i_2_), .Y(ori_ori_n140_));
  NA3        o130(.A(ori_ori_n140_), .B(ori_ori_n38_), .C(ori_ori_n112_), .Y(ori_ori_n141_));
  NA3        o131(.A(ori_ori_n54_), .B(ori_ori_n44_), .C(ori_ori_n18_), .Y(ori_ori_n142_));
  NOi32      o132(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n143_));
  NA2        o133(.A(ori_ori_n143_), .B(ori_ori_n130_), .Y(ori_ori_n144_));
  NA3        o134(.A(ori_ori_n140_), .B(ori_ori_n63_), .C(ori_ori_n37_), .Y(ori_ori_n145_));
  NA4        o135(.A(ori_ori_n145_), .B(ori_ori_n144_), .C(ori_ori_n142_), .D(ori_ori_n141_), .Y(ori_ori_n146_));
  NA3        o136(.A(ori_ori_n61_), .B(ori_ori_n14_), .C(i_7_), .Y(ori_ori_n147_));
  NA4        o137(.A(ori_ori_n64_), .B(ori_ori_n39_), .C(ori_ori_n17_), .D(i_8_), .Y(ori_ori_n148_));
  NA4        o138(.A(ori_ori_n64_), .B(ori_ori_n47_), .C(i_5_), .D(ori_ori_n23_), .Y(ori_ori_n149_));
  NA3        o139(.A(ori_ori_n149_), .B(ori_ori_n148_), .C(ori_ori_n147_), .Y(ori_ori_n150_));
  NO4        o140(.A(ori_ori_n150_), .B(ori_ori_n146_), .C(ori_ori_n139_), .D(ori_ori_n137_), .Y(ori_ori_n151_));
  AOI220     o141(.A0(i_5_), .A1(ori_ori_n94_), .B0(ori_ori_n67_), .B1(ori_ori_n32_), .Y(ori_ori_n152_));
  AOI210     o142(.A0(ori_ori_n152_), .A1(ori_ori_n129_), .B0(ori_ori_n108_), .Y(ori_ori_n153_));
  NO3        o143(.A(i_2_), .B(ori_ori_n21_), .C(ori_ori_n11_), .Y(ori_ori_n154_));
  NA2        o144(.A(i_2_), .B(i_4_), .Y(ori_ori_n155_));
  AOI210     o145(.A0(ori_ori_n110_), .A1(ori_ori_n91_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NO2        o146(.A(i_8_), .B(i_7_), .Y(ori_ori_n157_));
  OA210      o147(.A0(ori_ori_n156_), .A1(ori_ori_n154_), .B0(ori_ori_n157_), .Y(ori_ori_n158_));
  NA3        o148(.A(ori_ori_n122_), .B(i_0_), .C(ori_ori_n23_), .Y(ori_ori_n159_));
  NO2        o149(.A(ori_ori_n159_), .B(i_4_), .Y(ori_ori_n160_));
  NO3        o150(.A(ori_ori_n160_), .B(ori_ori_n158_), .C(ori_ori_n153_), .Y(ori_ori_n161_));
  NA2        o151(.A(ori_ori_n94_), .B(ori_ori_n12_), .Y(ori_ori_n162_));
  NA2        o152(.A(i_2_), .B(ori_ori_n14_), .Y(ori_ori_n163_));
  NA2        o153(.A(ori_ori_n54_), .B(i_3_), .Y(ori_ori_n164_));
  AOI210     o154(.A0(ori_ori_n164_), .A1(ori_ori_n163_), .B0(ori_ori_n162_), .Y(ori_ori_n165_));
  NA3        o155(.A(ori_ori_n140_), .B(ori_ori_n69_), .C(ori_ori_n112_), .Y(ori_ori_n166_));
  OAI210     o156(.A0(ori_ori_n107_), .A1(ori_ori_n31_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  NA4        o157(.A(ori_ori_n113_), .B(ori_ori_n67_), .C(ori_ori_n46_), .D(ori_ori_n21_), .Y(ori_ori_n168_));
  NA3        o158(.A(ori_ori_n57_), .B(ori_ori_n36_), .C(ori_ori_n15_), .Y(ori_ori_n169_));
  NOi31      o159(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n170_));
  OAI210     o160(.A0(ori_ori_n143_), .A1(ori_ori_n84_), .B0(ori_ori_n170_), .Y(ori_ori_n171_));
  NA3        o161(.A(ori_ori_n171_), .B(ori_ori_n169_), .C(ori_ori_n168_), .Y(ori_ori_n172_));
  NO3        o162(.A(ori_ori_n172_), .B(ori_ori_n167_), .C(ori_ori_n165_), .Y(ori_ori_n173_));
  NA4        o163(.A(ori_ori_n173_), .B(ori_ori_n161_), .C(ori_ori_n151_), .D(ori_ori_n135_), .Y(ori_ori_n174_));
  OR4        o164(.A(ori_ori_n174_), .B(ori_ori_n128_), .C(ori_ori_n90_), .D(ori_ori_n73_), .Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NA3        m013(.A(i_6_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_8_), .B(i_6_), .Y(mai_mai_n25_));
  NOi21      m015(.An(i_1_), .B(i_8_), .Y(mai_mai_n26_));
  AOI220     m016(.A0(mai_mai_n26_), .A1(i_2_), .B0(mai_mai_n25_), .B1(i_5_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n22_), .Y(mai_mai_n28_));
  AOI210     m018(.A0(mai_mai_n28_), .A1(mai_mai_n11_), .B0(mai_mai_n20_), .Y(mai_mai_n29_));
  NA2        m019(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n30_));
  NA2        m020(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n31_));
  NO2        m021(.A(i_2_), .B(i_4_), .Y(mai_mai_n32_));
  NA3        m022(.A(mai_mai_n32_), .B(i_6_), .C(i_8_), .Y(mai_mai_n33_));
  AOI210     m023(.A0(mai_mai_n31_), .A1(mai_mai_n30_), .B0(mai_mai_n33_), .Y(mai_mai_n34_));
  INV        m024(.A(i_2_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_6_), .B(i_8_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_7_), .B(i_1_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_5_), .B(i_6_), .Y(mai_mai_n38_));
  AOI220     m028(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n36_), .B1(i_5_), .Y(mai_mai_n39_));
  NO3        m029(.A(mai_mai_n39_), .B(mai_mai_n35_), .C(i_4_), .Y(mai_mai_n40_));
  NOi21      m030(.An(i_0_), .B(i_4_), .Y(mai_mai_n41_));
  XO2        m031(.A(i_1_), .B(i_3_), .Y(mai_mai_n42_));
  NOi21      m032(.An(i_7_), .B(i_5_), .Y(mai_mai_n43_));
  AN3        m033(.A(mai_mai_n43_), .B(mai_mai_n42_), .C(mai_mai_n41_), .Y(mai_mai_n44_));
  INV        m034(.A(i_1_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_3_), .B(i_0_), .Y(mai_mai_n46_));
  NA2        m036(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NA3        m037(.A(i_6_), .B(mai_mai_n14_), .C(i_7_), .Y(mai_mai_n48_));
  AOI210     m038(.A0(mai_mai_n48_), .A1(mai_mai_n24_), .B0(mai_mai_n47_), .Y(mai_mai_n49_));
  NO4        m039(.A(mai_mai_n49_), .B(mai_mai_n44_), .C(mai_mai_n40_), .D(mai_mai_n34_), .Y(mai_mai_n50_));
  NA2        m040(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n51_));
  NOi21      m041(.An(i_4_), .B(i_0_), .Y(mai_mai_n52_));
  NO2        m042(.A(mai_mai_n25_), .B(mai_mai_n15_), .Y(mai_mai_n53_));
  NA2        m043(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n54_));
  NOi21      m044(.An(i_2_), .B(i_8_), .Y(mai_mai_n55_));
  NO3        m045(.A(mai_mai_n55_), .B(mai_mai_n52_), .C(mai_mai_n41_), .Y(mai_mai_n56_));
  NO3        m046(.A(mai_mai_n56_), .B(mai_mai_n54_), .C(mai_mai_n53_), .Y(mai_mai_n57_));
  INV        m047(.A(mai_mai_n57_), .Y(mai_mai_n58_));
  NOi31      m048(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n59_));
  NA2        m049(.A(mai_mai_n59_), .B(i_0_), .Y(mai_mai_n60_));
  NOi21      m050(.An(i_4_), .B(i_3_), .Y(mai_mai_n61_));
  NOi21      m051(.An(i_1_), .B(i_4_), .Y(mai_mai_n62_));
  OAI210     m052(.A0(mai_mai_n62_), .A1(mai_mai_n61_), .B0(mai_mai_n55_), .Y(mai_mai_n63_));
  NA2        m053(.A(mai_mai_n63_), .B(mai_mai_n60_), .Y(mai_mai_n64_));
  AN2        m054(.A(i_8_), .B(i_7_), .Y(mai_mai_n65_));
  INV        m055(.A(mai_mai_n65_), .Y(mai_mai_n66_));
  NOi21      m056(.An(i_8_), .B(i_7_), .Y(mai_mai_n67_));
  NA3        m057(.A(mai_mai_n67_), .B(mai_mai_n61_), .C(i_6_), .Y(mai_mai_n68_));
  OAI210     m058(.A0(mai_mai_n66_), .A1(mai_mai_n54_), .B0(mai_mai_n68_), .Y(mai_mai_n69_));
  AOI220     m059(.A0(mai_mai_n69_), .A1(mai_mai_n35_), .B0(mai_mai_n64_), .B1(mai_mai_n38_), .Y(mai_mai_n70_));
  NA4        m060(.A(mai_mai_n70_), .B(mai_mai_n58_), .C(mai_mai_n50_), .D(mai_mai_n29_), .Y(mai_mai_n71_));
  NA2        m061(.A(i_8_), .B(i_7_), .Y(mai_mai_n72_));
  NO3        m062(.A(mai_mai_n72_), .B(mai_mai_n13_), .C(i_1_), .Y(mai_mai_n73_));
  NA2        m063(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n74_));
  AOI220     m064(.A0(mai_mai_n46_), .A1(i_1_), .B0(mai_mai_n42_), .B1(i_2_), .Y(mai_mai_n75_));
  NOi21      m065(.An(i_1_), .B(i_2_), .Y(mai_mai_n76_));
  NO2        m066(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n77_));
  OAI210     m067(.A0(mai_mai_n77_), .A1(mai_mai_n73_), .B0(mai_mai_n14_), .Y(mai_mai_n78_));
  NA3        m068(.A(mai_mai_n67_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n79_));
  NA3        m069(.A(mai_mai_n26_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n80_));
  NA2        m070(.A(mai_mai_n80_), .B(mai_mai_n79_), .Y(mai_mai_n81_));
  NOi32      m071(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n82_), .B(i_3_), .Y(mai_mai_n83_));
  NA2        m073(.A(mai_mai_n18_), .B(i_6_), .Y(mai_mai_n84_));
  NA2        m074(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n85_));
  NO2        m075(.A(i_0_), .B(i_4_), .Y(mai_mai_n86_));
  AOI220     m076(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n81_), .B1(mai_mai_n61_), .Y(mai_mai_n87_));
  NA2        m077(.A(mai_mai_n87_), .B(mai_mai_n78_), .Y(mai_mai_n88_));
  INV        m078(.A(i_6_), .Y(mai_mai_n89_));
  NO2        m079(.A(mai_mai_n89_), .B(i_0_), .Y(mai_mai_n90_));
  NOi21      m080(.An(i_7_), .B(i_8_), .Y(mai_mai_n91_));
  NOi31      m081(.An(i_6_), .B(i_5_), .C(i_7_), .Y(mai_mai_n92_));
  NO2        m082(.A(mai_mai_n91_), .B(mai_mai_n92_), .Y(mai_mai_n93_));
  NO2        m083(.A(mai_mai_n93_), .B(mai_mai_n11_), .Y(mai_mai_n94_));
  OAI210     m084(.A0(mai_mai_n94_), .A1(mai_mai_n90_), .B0(mai_mai_n76_), .Y(mai_mai_n95_));
  NA3        m085(.A(mai_mai_n25_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n96_));
  AOI210     m086(.A0(mai_mai_n22_), .A1(mai_mai_n51_), .B0(mai_mai_n96_), .Y(mai_mai_n97_));
  AOI220     m087(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n18_), .B1(mai_mai_n35_), .Y(mai_mai_n98_));
  NA3        m088(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n99_));
  NA2        m089(.A(i_4_), .B(i_5_), .Y(mai_mai_n100_));
  NA3        m090(.A(mai_mai_n72_), .B(mai_mai_n18_), .C(mai_mai_n17_), .Y(mai_mai_n101_));
  OAI220     m091(.A0(mai_mai_n101_), .A1(mai_mai_n100_), .B0(mai_mai_n99_), .B1(mai_mai_n98_), .Y(mai_mai_n102_));
  NO2        m092(.A(mai_mai_n102_), .B(mai_mai_n97_), .Y(mai_mai_n103_));
  NA3        m093(.A(mai_mai_n67_), .B(mai_mai_n35_), .C(i_3_), .Y(mai_mai_n104_));
  NA2        m094(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n105_));
  AOI210     m095(.A0(mai_mai_n105_), .A1(mai_mai_n22_), .B0(mai_mai_n104_), .Y(mai_mai_n106_));
  NOi21      m096(.An(i_2_), .B(i_1_), .Y(mai_mai_n107_));
  AN3        m097(.A(mai_mai_n91_), .B(mai_mai_n107_), .C(mai_mai_n52_), .Y(mai_mai_n108_));
  NAi21      m098(.An(i_6_), .B(i_0_), .Y(mai_mai_n109_));
  NA3        m099(.A(mai_mai_n62_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n110_));
  NOi21      m100(.An(i_4_), .B(i_6_), .Y(mai_mai_n111_));
  NOi21      m101(.An(i_5_), .B(i_3_), .Y(mai_mai_n112_));
  NA3        m102(.A(mai_mai_n112_), .B(mai_mai_n76_), .C(mai_mai_n111_), .Y(mai_mai_n113_));
  OAI210     m103(.A0(mai_mai_n110_), .A1(mai_mai_n109_), .B0(mai_mai_n113_), .Y(mai_mai_n114_));
  NA2        m104(.A(mai_mai_n76_), .B(mai_mai_n36_), .Y(mai_mai_n115_));
  NO3        m105(.A(mai_mai_n114_), .B(mai_mai_n108_), .C(mai_mai_n106_), .Y(mai_mai_n116_));
  AOI220     m106(.A0(i_6_), .A1(i_7_), .B0(mai_mai_n25_), .B1(i_5_), .Y(mai_mai_n117_));
  NOi31      m107(.An(mai_mai_n52_), .B(mai_mai_n117_), .C(i_2_), .Y(mai_mai_n118_));
  NA2        m108(.A(mai_mai_n67_), .B(mai_mai_n12_), .Y(mai_mai_n119_));
  NA2        m109(.A(mai_mai_n36_), .B(mai_mai_n14_), .Y(mai_mai_n120_));
  NOi21      m110(.An(i_3_), .B(i_1_), .Y(mai_mai_n121_));
  NA2        m111(.A(mai_mai_n121_), .B(i_4_), .Y(mai_mai_n122_));
  AOI210     m112(.A0(mai_mai_n120_), .A1(mai_mai_n119_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  AOI220     m113(.A0(mai_mai_n91_), .A1(mai_mai_n14_), .B0(mai_mai_n111_), .B1(mai_mai_n23_), .Y(mai_mai_n124_));
  NOi31      m114(.An(mai_mai_n46_), .B(mai_mai_n124_), .C(mai_mai_n35_), .Y(mai_mai_n125_));
  NO3        m115(.A(mai_mai_n125_), .B(mai_mai_n123_), .C(mai_mai_n118_), .Y(mai_mai_n126_));
  NA4        m116(.A(mai_mai_n126_), .B(mai_mai_n116_), .C(mai_mai_n103_), .D(mai_mai_n95_), .Y(mai_mai_n127_));
  NA2        m117(.A(mai_mai_n55_), .B(mai_mai_n15_), .Y(mai_mai_n128_));
  NOi31      m118(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n129_));
  NOi31      m119(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n130_));
  OAI210     m120(.A0(mai_mai_n130_), .A1(mai_mai_n129_), .B0(i_7_), .Y(mai_mai_n131_));
  NA3        m121(.A(mai_mai_n36_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n132_));
  NA4        m122(.A(mai_mai_n132_), .B(mai_mai_n131_), .C(mai_mai_n128_), .D(mai_mai_n115_), .Y(mai_mai_n133_));
  NA2        m123(.A(mai_mai_n133_), .B(mai_mai_n41_), .Y(mai_mai_n134_));
  NA2        m124(.A(mai_mai_n61_), .B(mai_mai_n37_), .Y(mai_mai_n135_));
  AOI210     m125(.A0(mai_mai_n135_), .A1(mai_mai_n79_), .B0(mai_mai_n31_), .Y(mai_mai_n136_));
  NA4        m126(.A(mai_mai_n65_), .B(mai_mai_n107_), .C(mai_mai_n17_), .D(mai_mai_n12_), .Y(mai_mai_n137_));
  NAi31      m127(.An(mai_mai_n109_), .B(mai_mai_n91_), .C(mai_mai_n107_), .Y(mai_mai_n138_));
  NA3        m128(.A(mai_mai_n67_), .B(mai_mai_n59_), .C(i_6_), .Y(mai_mai_n139_));
  NA3        m129(.A(mai_mai_n139_), .B(mai_mai_n138_), .C(mai_mai_n137_), .Y(mai_mai_n140_));
  NOi21      m130(.An(i_0_), .B(i_2_), .Y(mai_mai_n141_));
  NA3        m131(.A(mai_mai_n141_), .B(mai_mai_n37_), .C(mai_mai_n111_), .Y(mai_mai_n142_));
  NA3        m132(.A(mai_mai_n52_), .B(mai_mai_n43_), .C(mai_mai_n18_), .Y(mai_mai_n143_));
  NOi32      m133(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(mai_mai_n144_));
  NA2        m134(.A(mai_mai_n144_), .B(mai_mai_n129_), .Y(mai_mai_n145_));
  NA3        m135(.A(mai_mai_n141_), .B(mai_mai_n61_), .C(mai_mai_n36_), .Y(mai_mai_n146_));
  NA4        m136(.A(mai_mai_n146_), .B(mai_mai_n145_), .C(mai_mai_n143_), .D(mai_mai_n142_), .Y(mai_mai_n147_));
  NA4        m137(.A(mai_mai_n59_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n148_));
  NA4        m138(.A(mai_mai_n62_), .B(mai_mai_n38_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n149_));
  NA4        m139(.A(mai_mai_n62_), .B(mai_mai_n46_), .C(i_5_), .D(mai_mai_n23_), .Y(mai_mai_n150_));
  NA3        m140(.A(mai_mai_n150_), .B(mai_mai_n149_), .C(mai_mai_n148_), .Y(mai_mai_n151_));
  NO4        m141(.A(mai_mai_n151_), .B(mai_mai_n147_), .C(mai_mai_n140_), .D(mai_mai_n136_), .Y(mai_mai_n152_));
  NOi21      m142(.An(i_5_), .B(i_2_), .Y(mai_mai_n153_));
  AOI220     m143(.A0(mai_mai_n153_), .A1(mai_mai_n91_), .B0(mai_mai_n65_), .B1(mai_mai_n32_), .Y(mai_mai_n154_));
  AOI210     m144(.A0(mai_mai_n154_), .A1(mai_mai_n128_), .B0(mai_mai_n105_), .Y(mai_mai_n155_));
  NO4        m145(.A(i_2_), .B(mai_mai_n21_), .C(mai_mai_n11_), .D(mai_mai_n14_), .Y(mai_mai_n156_));
  NA2        m146(.A(i_2_), .B(i_4_), .Y(mai_mai_n157_));
  AOI210     m147(.A0(mai_mai_n109_), .A1(mai_mai_n89_), .B0(mai_mai_n157_), .Y(mai_mai_n158_));
  NO2        m148(.A(i_8_), .B(i_7_), .Y(mai_mai_n159_));
  OA210      m149(.A0(mai_mai_n158_), .A1(mai_mai_n156_), .B0(mai_mai_n159_), .Y(mai_mai_n160_));
  NA4        m150(.A(mai_mai_n121_), .B(i_0_), .C(i_5_), .D(mai_mai_n23_), .Y(mai_mai_n161_));
  NO2        m151(.A(mai_mai_n161_), .B(i_4_), .Y(mai_mai_n162_));
  NO3        m152(.A(mai_mai_n162_), .B(mai_mai_n160_), .C(mai_mai_n155_), .Y(mai_mai_n163_));
  NA2        m153(.A(mai_mai_n91_), .B(mai_mai_n12_), .Y(mai_mai_n164_));
  NA3        m154(.A(i_2_), .B(i_1_), .C(mai_mai_n14_), .Y(mai_mai_n165_));
  NA2        m155(.A(mai_mai_n52_), .B(i_3_), .Y(mai_mai_n166_));
  AOI210     m156(.A0(mai_mai_n166_), .A1(mai_mai_n165_), .B0(mai_mai_n164_), .Y(mai_mai_n167_));
  NA3        m157(.A(mai_mai_n141_), .B(mai_mai_n67_), .C(mai_mai_n111_), .Y(mai_mai_n168_));
  OAI210     m158(.A0(mai_mai_n104_), .A1(mai_mai_n31_), .B0(mai_mai_n168_), .Y(mai_mai_n169_));
  NA4        m159(.A(mai_mai_n112_), .B(mai_mai_n65_), .C(mai_mai_n45_), .D(mai_mai_n21_), .Y(mai_mai_n170_));
  NA3        m160(.A(mai_mai_n92_), .B(mai_mai_n121_), .C(i_0_), .Y(mai_mai_n171_));
  NOi31      m161(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n172_));
  OAI210     m162(.A0(mai_mai_n144_), .A1(mai_mai_n82_), .B0(mai_mai_n172_), .Y(mai_mai_n173_));
  NA3        m163(.A(mai_mai_n173_), .B(mai_mai_n171_), .C(mai_mai_n170_), .Y(mai_mai_n174_));
  NO3        m164(.A(mai_mai_n174_), .B(mai_mai_n169_), .C(mai_mai_n167_), .Y(mai_mai_n175_));
  NA4        m165(.A(mai_mai_n175_), .B(mai_mai_n163_), .C(mai_mai_n152_), .D(mai_mai_n134_), .Y(mai_mai_n176_));
  OR4        m166(.A(mai_mai_n176_), .B(mai_mai_n127_), .C(mai_mai_n88_), .D(mai_mai_n71_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NA3        u013(.A(i_6_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n24_));
  NOi21      u014(.An(i_8_), .B(i_6_), .Y(men_men_n25_));
  NOi21      u015(.An(i_1_), .B(i_8_), .Y(men_men_n26_));
  AOI220     u016(.A0(men_men_n26_), .A1(i_2_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n22_), .Y(men_men_n28_));
  AOI210     u018(.A0(men_men_n28_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n29_));
  NA2        u019(.A(i_0_), .B(men_men_n14_), .Y(men_men_n30_));
  NA2        u020(.A(men_men_n17_), .B(i_5_), .Y(men_men_n31_));
  NO2        u021(.A(i_2_), .B(i_4_), .Y(men_men_n32_));
  NA3        u022(.A(men_men_n32_), .B(i_6_), .C(i_8_), .Y(men_men_n33_));
  AOI210     u023(.A0(men_men_n31_), .A1(men_men_n30_), .B0(men_men_n33_), .Y(men_men_n34_));
  INV        u024(.A(i_2_), .Y(men_men_n35_));
  NOi21      u025(.An(i_5_), .B(i_0_), .Y(men_men_n36_));
  NOi21      u026(.An(i_6_), .B(i_8_), .Y(men_men_n37_));
  NOi21      u027(.An(i_7_), .B(i_1_), .Y(men_men_n38_));
  NOi21      u028(.An(i_5_), .B(i_6_), .Y(men_men_n39_));
  AOI220     u029(.A0(men_men_n39_), .A1(men_men_n38_), .B0(men_men_n37_), .B1(men_men_n36_), .Y(men_men_n40_));
  NO3        u030(.A(men_men_n40_), .B(men_men_n35_), .C(i_4_), .Y(men_men_n41_));
  NOi21      u031(.An(i_0_), .B(i_4_), .Y(men_men_n42_));
  XO2        u032(.A(i_1_), .B(i_3_), .Y(men_men_n43_));
  NOi21      u033(.An(i_7_), .B(i_5_), .Y(men_men_n44_));
  AN3        u034(.A(men_men_n44_), .B(men_men_n43_), .C(men_men_n42_), .Y(men_men_n45_));
  INV        u035(.A(i_1_), .Y(men_men_n46_));
  NOi21      u036(.An(i_3_), .B(i_0_), .Y(men_men_n47_));
  NA2        u037(.A(men_men_n47_), .B(men_men_n46_), .Y(men_men_n48_));
  NO2        u038(.A(men_men_n24_), .B(men_men_n48_), .Y(men_men_n49_));
  NO4        u039(.A(men_men_n49_), .B(men_men_n45_), .C(men_men_n41_), .D(men_men_n34_), .Y(men_men_n50_));
  INV        u040(.A(i_8_), .Y(men_men_n51_));
  NA2        u041(.A(i_1_), .B(men_men_n11_), .Y(men_men_n52_));
  NO4        u042(.A(men_men_n52_), .B(men_men_n30_), .C(i_2_), .D(men_men_n51_), .Y(men_men_n53_));
  NOi21      u043(.An(i_4_), .B(i_0_), .Y(men_men_n54_));
  AOI210     u044(.A0(men_men_n54_), .A1(men_men_n25_), .B0(men_men_n15_), .Y(men_men_n55_));
  NA2        u045(.A(i_1_), .B(men_men_n14_), .Y(men_men_n56_));
  NOi21      u046(.An(i_2_), .B(i_8_), .Y(men_men_n57_));
  NO3        u047(.A(men_men_n57_), .B(men_men_n54_), .C(men_men_n42_), .Y(men_men_n58_));
  NO3        u048(.A(men_men_n58_), .B(men_men_n56_), .C(men_men_n55_), .Y(men_men_n59_));
  NO2        u049(.A(men_men_n59_), .B(men_men_n53_), .Y(men_men_n60_));
  NOi31      u050(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n61_));
  NA2        u051(.A(men_men_n61_), .B(i_0_), .Y(men_men_n62_));
  NOi21      u052(.An(i_4_), .B(i_3_), .Y(men_men_n63_));
  NOi21      u053(.An(i_1_), .B(i_4_), .Y(men_men_n64_));
  OAI210     u054(.A0(men_men_n64_), .A1(men_men_n63_), .B0(men_men_n57_), .Y(men_men_n65_));
  NA2        u055(.A(men_men_n65_), .B(men_men_n62_), .Y(men_men_n66_));
  AN2        u056(.A(i_8_), .B(i_7_), .Y(men_men_n67_));
  NA2        u057(.A(men_men_n67_), .B(men_men_n12_), .Y(men_men_n68_));
  NOi21      u058(.An(i_8_), .B(i_7_), .Y(men_men_n69_));
  NA3        u059(.A(men_men_n69_), .B(men_men_n63_), .C(i_6_), .Y(men_men_n70_));
  OAI210     u060(.A0(men_men_n68_), .A1(men_men_n56_), .B0(men_men_n70_), .Y(men_men_n71_));
  AOI220     u061(.A0(men_men_n71_), .A1(men_men_n35_), .B0(men_men_n66_), .B1(men_men_n39_), .Y(men_men_n72_));
  NA4        u062(.A(men_men_n72_), .B(men_men_n60_), .C(men_men_n50_), .D(men_men_n29_), .Y(men_men_n73_));
  NA2        u063(.A(i_8_), .B(i_7_), .Y(men_men_n74_));
  NO3        u064(.A(men_men_n74_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n75_));
  NA2        u065(.A(i_8_), .B(men_men_n23_), .Y(men_men_n76_));
  AOI220     u066(.A0(men_men_n47_), .A1(i_1_), .B0(men_men_n43_), .B1(i_2_), .Y(men_men_n77_));
  NOi21      u067(.An(i_1_), .B(i_2_), .Y(men_men_n78_));
  NA3        u068(.A(men_men_n78_), .B(men_men_n54_), .C(i_6_), .Y(men_men_n79_));
  OAI210     u069(.A0(men_men_n77_), .A1(men_men_n76_), .B0(men_men_n79_), .Y(men_men_n80_));
  OAI210     u070(.A0(men_men_n80_), .A1(men_men_n75_), .B0(men_men_n14_), .Y(men_men_n81_));
  NA3        u071(.A(men_men_n69_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n82_));
  NA3        u072(.A(men_men_n26_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n83_));
  NA2        u073(.A(men_men_n83_), .B(men_men_n82_), .Y(men_men_n84_));
  NOi32      u074(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n85_));
  NA2        u075(.A(men_men_n85_), .B(i_3_), .Y(men_men_n86_));
  NA3        u076(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n87_));
  NA2        u077(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u078(.A(i_0_), .Y(men_men_n89_));
  AOI220     u079(.A0(men_men_n89_), .A1(men_men_n88_), .B0(men_men_n84_), .B1(men_men_n63_), .Y(men_men_n90_));
  NA2        u080(.A(men_men_n90_), .B(men_men_n81_), .Y(men_men_n91_));
  NAi21      u081(.An(i_3_), .B(i_6_), .Y(men_men_n92_));
  NO3        u082(.A(men_men_n92_), .B(i_0_), .C(men_men_n51_), .Y(men_men_n93_));
  NA2        u083(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n94_));
  NOi21      u084(.An(i_7_), .B(i_8_), .Y(men_men_n95_));
  NOi31      u085(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n96_));
  AOI210     u086(.A0(men_men_n95_), .A1(men_men_n12_), .B0(men_men_n96_), .Y(men_men_n97_));
  OAI210     u087(.A0(men_men_n97_), .A1(men_men_n11_), .B0(men_men_n94_), .Y(men_men_n98_));
  OAI210     u088(.A0(men_men_n98_), .A1(men_men_n93_), .B0(men_men_n78_), .Y(men_men_n99_));
  NA3        u089(.A(men_men_n25_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n100_));
  AOI210     u090(.A0(men_men_n22_), .A1(men_men_n52_), .B0(men_men_n100_), .Y(men_men_n101_));
  AOI220     u091(.A0(men_men_n47_), .A1(men_men_n46_), .B0(men_men_n18_), .B1(men_men_n35_), .Y(men_men_n102_));
  NA3        u092(.A(men_men_n21_), .B(i_5_), .C(i_7_), .Y(men_men_n103_));
  NO2        u093(.A(men_men_n103_), .B(men_men_n102_), .Y(men_men_n104_));
  NO2        u094(.A(men_men_n104_), .B(men_men_n101_), .Y(men_men_n105_));
  NA3        u095(.A(men_men_n69_), .B(men_men_n35_), .C(i_3_), .Y(men_men_n106_));
  NA2        u096(.A(men_men_n46_), .B(i_6_), .Y(men_men_n107_));
  AOI210     u097(.A0(men_men_n107_), .A1(men_men_n22_), .B0(men_men_n106_), .Y(men_men_n108_));
  NOi21      u098(.An(i_2_), .B(i_1_), .Y(men_men_n109_));
  AN3        u099(.A(men_men_n95_), .B(men_men_n109_), .C(men_men_n54_), .Y(men_men_n110_));
  NAi21      u100(.An(i_6_), .B(i_0_), .Y(men_men_n111_));
  NA3        u101(.A(men_men_n64_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n112_));
  NOi21      u102(.An(i_4_), .B(i_6_), .Y(men_men_n113_));
  NOi21      u103(.An(i_5_), .B(i_3_), .Y(men_men_n114_));
  NA3        u104(.A(men_men_n114_), .B(men_men_n78_), .C(men_men_n113_), .Y(men_men_n115_));
  OAI210     u105(.A0(men_men_n112_), .A1(men_men_n111_), .B0(men_men_n115_), .Y(men_men_n116_));
  NA2        u106(.A(men_men_n78_), .B(men_men_n37_), .Y(men_men_n117_));
  NOi21      u107(.An(men_men_n44_), .B(men_men_n117_), .Y(men_men_n118_));
  NO4        u108(.A(men_men_n118_), .B(men_men_n116_), .C(men_men_n110_), .D(men_men_n108_), .Y(men_men_n119_));
  NOi21      u109(.An(i_6_), .B(i_1_), .Y(men_men_n120_));
  AOI220     u110(.A0(men_men_n120_), .A1(i_7_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n121_));
  NOi31      u111(.An(men_men_n54_), .B(men_men_n121_), .C(i_2_), .Y(men_men_n122_));
  NA2        u112(.A(men_men_n69_), .B(men_men_n12_), .Y(men_men_n123_));
  NA2        u113(.A(men_men_n37_), .B(men_men_n14_), .Y(men_men_n124_));
  NOi21      u114(.An(i_3_), .B(i_1_), .Y(men_men_n125_));
  NA2        u115(.A(men_men_n125_), .B(i_4_), .Y(men_men_n126_));
  AOI210     u116(.A0(men_men_n124_), .A1(men_men_n123_), .B0(men_men_n126_), .Y(men_men_n127_));
  NOi31      u117(.An(men_men_n47_), .B(i_5_), .C(men_men_n35_), .Y(men_men_n128_));
  NO3        u118(.A(men_men_n128_), .B(men_men_n127_), .C(men_men_n122_), .Y(men_men_n129_));
  NA4        u119(.A(men_men_n129_), .B(men_men_n119_), .C(men_men_n105_), .D(men_men_n99_), .Y(men_men_n130_));
  NA2        u120(.A(men_men_n57_), .B(men_men_n15_), .Y(men_men_n131_));
  NOi31      u121(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n132_));
  NOi31      u122(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n133_));
  OAI210     u123(.A0(men_men_n133_), .A1(men_men_n132_), .B0(i_7_), .Y(men_men_n134_));
  NA3        u124(.A(men_men_n37_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n135_));
  NA4        u125(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n131_), .D(men_men_n117_), .Y(men_men_n136_));
  NA2        u126(.A(men_men_n136_), .B(men_men_n42_), .Y(men_men_n137_));
  NA2        u127(.A(men_men_n63_), .B(men_men_n38_), .Y(men_men_n138_));
  AOI210     u128(.A0(men_men_n138_), .A1(men_men_n82_), .B0(men_men_n31_), .Y(men_men_n139_));
  NA4        u129(.A(men_men_n67_), .B(men_men_n109_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n140_));
  NAi31      u130(.An(men_men_n111_), .B(men_men_n95_), .C(men_men_n109_), .Y(men_men_n141_));
  NA3        u131(.A(men_men_n69_), .B(men_men_n61_), .C(i_6_), .Y(men_men_n142_));
  NA3        u132(.A(men_men_n142_), .B(men_men_n141_), .C(men_men_n140_), .Y(men_men_n143_));
  NOi21      u133(.An(i_0_), .B(i_2_), .Y(men_men_n144_));
  NA3        u134(.A(men_men_n144_), .B(men_men_n38_), .C(men_men_n113_), .Y(men_men_n145_));
  NOi32      u135(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n146_));
  NA2        u136(.A(men_men_n146_), .B(men_men_n132_), .Y(men_men_n147_));
  NA3        u137(.A(men_men_n144_), .B(men_men_n63_), .C(men_men_n37_), .Y(men_men_n148_));
  NA3        u138(.A(men_men_n148_), .B(men_men_n147_), .C(men_men_n145_), .Y(men_men_n149_));
  NA4        u139(.A(men_men_n61_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n150_));
  NA4        u140(.A(men_men_n64_), .B(men_men_n39_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n151_));
  NA4        u141(.A(men_men_n64_), .B(men_men_n47_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n152_));
  NA3        u142(.A(men_men_n152_), .B(men_men_n151_), .C(men_men_n150_), .Y(men_men_n153_));
  NO4        u143(.A(men_men_n153_), .B(men_men_n149_), .C(men_men_n143_), .D(men_men_n139_), .Y(men_men_n154_));
  NA2        u144(.A(men_men_n67_), .B(men_men_n32_), .Y(men_men_n155_));
  AOI210     u145(.A0(men_men_n155_), .A1(men_men_n131_), .B0(men_men_n107_), .Y(men_men_n156_));
  NO4        u146(.A(i_2_), .B(men_men_n21_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n157_));
  NA2        u147(.A(i_2_), .B(i_4_), .Y(men_men_n158_));
  AOI210     u148(.A0(men_men_n111_), .A1(men_men_n92_), .B0(men_men_n158_), .Y(men_men_n159_));
  NO2        u149(.A(i_8_), .B(i_7_), .Y(men_men_n160_));
  OA210      u150(.A0(men_men_n159_), .A1(men_men_n157_), .B0(men_men_n160_), .Y(men_men_n161_));
  NA4        u151(.A(men_men_n125_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n162_));
  NO2        u152(.A(men_men_n162_), .B(i_4_), .Y(men_men_n163_));
  NO3        u153(.A(men_men_n163_), .B(men_men_n161_), .C(men_men_n156_), .Y(men_men_n164_));
  NA2        u154(.A(men_men_n95_), .B(men_men_n12_), .Y(men_men_n165_));
  NA2        u155(.A(i_1_), .B(men_men_n14_), .Y(men_men_n166_));
  NA2        u156(.A(men_men_n54_), .B(i_3_), .Y(men_men_n167_));
  AOI210     u157(.A0(men_men_n167_), .A1(men_men_n166_), .B0(men_men_n165_), .Y(men_men_n168_));
  NA3        u158(.A(men_men_n144_), .B(men_men_n69_), .C(men_men_n113_), .Y(men_men_n169_));
  OAI210     u159(.A0(men_men_n106_), .A1(men_men_n31_), .B0(men_men_n169_), .Y(men_men_n170_));
  NA4        u160(.A(men_men_n114_), .B(men_men_n67_), .C(men_men_n46_), .D(men_men_n21_), .Y(men_men_n171_));
  NA3        u161(.A(men_men_n96_), .B(men_men_n125_), .C(i_0_), .Y(men_men_n172_));
  NA3        u162(.A(men_men_n57_), .B(men_men_n36_), .C(men_men_n15_), .Y(men_men_n173_));
  NOi31      u163(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n174_));
  OAI210     u164(.A0(men_men_n146_), .A1(men_men_n85_), .B0(men_men_n174_), .Y(men_men_n175_));
  NA4        u165(.A(men_men_n175_), .B(men_men_n173_), .C(men_men_n172_), .D(men_men_n171_), .Y(men_men_n176_));
  NO3        u166(.A(men_men_n176_), .B(men_men_n170_), .C(men_men_n168_), .Y(men_men_n177_));
  NA4        u167(.A(men_men_n177_), .B(men_men_n164_), .C(men_men_n154_), .D(men_men_n137_), .Y(men_men_n178_));
  OR4        u168(.A(men_men_n178_), .B(men_men_n130_), .C(men_men_n91_), .D(men_men_n73_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule