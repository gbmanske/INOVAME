//Benchmark atmr_misex3_1774_0.25

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  INV        o000(.A(b), .Y(ori_ori_n29_));
  NOi32      o001(.An(i), .Bn(o), .C(h), .Y(ori_ori_n30_));
  NOi32      o002(.An(j), .Bn(o), .C(k), .Y(ori_ori_n31_));
  NA2        o003(.A(ori_ori_n31_), .B(m), .Y(ori_ori_n32_));
  NO2        o004(.A(ori_ori_n32_), .B(n), .Y(ori_ori_n33_));
  INV        o005(.A(h), .Y(ori_ori_n34_));
  INV        o006(.A(i), .Y(ori_ori_n35_));
  AN2        o007(.A(h), .B(o), .Y(ori_ori_n36_));
  NA2        o008(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n37_));
  NAi21      o009(.An(n), .B(m), .Y(ori_ori_n38_));
  NOi32      o010(.An(k), .Bn(h), .C(l), .Y(ori_ori_n39_));
  NOi32      o011(.An(k), .Bn(h), .C(o), .Y(ori_ori_n40_));
  INV        o012(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o013(.A(ori_ori_n41_), .B(ori_ori_n38_), .Y(ori_ori_n42_));
  INV        o014(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  NO2        o015(.A(ori_ori_n43_), .B(ori_ori_n29_), .Y(ori_ori_n44_));
  INV        o016(.A(c), .Y(ori_ori_n45_));
  NA2        o017(.A(e), .B(b), .Y(ori_ori_n46_));
  INV        o018(.A(d), .Y(ori_ori_n47_));
  NA2        o019(.A(o), .B(f), .Y(ori_ori_n48_));
  NAi31      o020(.An(l), .B(m), .C(k), .Y(ori_ori_n49_));
  NAi21      o021(.An(e), .B(h), .Y(ori_ori_n50_));
  INV        o022(.A(m), .Y(ori_ori_n51_));
  NOi21      o023(.An(k), .B(l), .Y(ori_ori_n52_));
  NA2        o024(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  AN4        o025(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n54_));
  NA2        o026(.A(h), .B(ori_ori_n54_), .Y(ori_ori_n55_));
  NAi32      o027(.An(m), .Bn(k), .C(j), .Y(ori_ori_n56_));
  OR2        o028(.A(ori_ori_n55_), .B(ori_ori_n53_), .Y(ori_ori_n57_));
  INV        o029(.A(ori_ori_n57_), .Y(ori_ori_n58_));
  INV        o030(.A(n), .Y(ori_ori_n59_));
  NOi32      o031(.An(e), .Bn(b), .C(d), .Y(ori_ori_n60_));
  INV        o032(.A(ori_ori_n60_), .Y(ori_ori_n61_));
  INV        o033(.A(j), .Y(ori_ori_n62_));
  AN3        o034(.A(m), .B(k), .C(i), .Y(ori_ori_n63_));
  NA3        o035(.A(ori_ori_n63_), .B(ori_ori_n62_), .C(o), .Y(ori_ori_n64_));
  NO2        o036(.A(ori_ori_n64_), .B(f), .Y(ori_ori_n65_));
  NAi32      o037(.An(o), .Bn(f), .C(h), .Y(ori_ori_n66_));
  NA2        o038(.A(m), .B(l), .Y(ori_ori_n67_));
  NA2        o039(.A(m), .B(l), .Y(ori_ori_n68_));
  NOi21      o040(.An(o), .B(i), .Y(ori_ori_n69_));
  NAi41      o041(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n70_));
  AN2        o042(.A(e), .B(b), .Y(ori_ori_n71_));
  NOi31      o043(.An(c), .B(h), .C(f), .Y(ori_ori_n72_));
  NA2        o044(.A(ori_ori_n72_), .B(ori_ori_n71_), .Y(ori_ori_n73_));
  NO2        o045(.A(ori_ori_n73_), .B(ori_ori_n70_), .Y(ori_ori_n74_));
  NOi21      o046(.An(i), .B(h), .Y(ori_ori_n75_));
  INV        o047(.A(a), .Y(ori_ori_n76_));
  INV        o048(.A(ori_ori_n71_), .Y(ori_ori_n77_));
  INV        o049(.A(l), .Y(ori_ori_n78_));
  NOi21      o050(.An(m), .B(n), .Y(ori_ori_n79_));
  AN2        o051(.A(k), .B(h), .Y(ori_ori_n80_));
  INV        o052(.A(b), .Y(ori_ori_n81_));
  NA2        o053(.A(l), .B(j), .Y(ori_ori_n82_));
  INV        o054(.A(ori_ori_n82_), .Y(ori_ori_n83_));
  INV        o055(.A(ori_ori_n74_), .Y(ori_ori_n84_));
  OAI210     o056(.A0(ori_ori_n64_), .A1(ori_ori_n61_), .B0(ori_ori_n84_), .Y(ori_ori_n85_));
  NOi31      o057(.An(k), .B(m), .C(j), .Y(ori_ori_n86_));
  NA3        o058(.A(ori_ori_n86_), .B(h), .C(ori_ori_n54_), .Y(ori_ori_n87_));
  NOi31      o059(.An(k), .B(m), .C(i), .Y(ori_ori_n88_));
  INV        o060(.A(ori_ori_n87_), .Y(ori_ori_n89_));
  NAi21      o061(.An(o), .B(h), .Y(ori_ori_n90_));
  NAi21      o062(.An(m), .B(n), .Y(ori_ori_n91_));
  NAi21      o063(.An(j), .B(k), .Y(ori_ori_n92_));
  NO3        o064(.A(ori_ori_n92_), .B(ori_ori_n91_), .C(ori_ori_n90_), .Y(ori_ori_n93_));
  NAi31      o065(.An(j), .B(k), .C(h), .Y(ori_ori_n94_));
  NA2        o066(.A(ori_ori_n93_), .B(f), .Y(ori_ori_n95_));
  INV        o067(.A(ori_ori_n91_), .Y(ori_ori_n96_));
  AN2        o068(.A(k), .B(j), .Y(ori_ori_n97_));
  NAi21      o069(.An(c), .B(b), .Y(ori_ori_n98_));
  NA2        o070(.A(f), .B(d), .Y(ori_ori_n99_));
  NO4        o071(.A(ori_ori_n99_), .B(ori_ori_n98_), .C(ori_ori_n97_), .D(ori_ori_n90_), .Y(ori_ori_n100_));
  NAi31      o072(.An(f), .B(e), .C(b), .Y(ori_ori_n101_));
  NA2        o073(.A(ori_ori_n100_), .B(ori_ori_n96_), .Y(ori_ori_n102_));
  NA2        o074(.A(d), .B(b), .Y(ori_ori_n103_));
  NAi21      o075(.An(e), .B(f), .Y(ori_ori_n104_));
  NA2        o076(.A(b), .B(a), .Y(ori_ori_n105_));
  NAi21      o077(.An(e), .B(o), .Y(ori_ori_n106_));
  NAi21      o078(.An(c), .B(d), .Y(ori_ori_n107_));
  NAi31      o079(.An(l), .B(k), .C(h), .Y(ori_ori_n108_));
  NAi31      o080(.An(ori_ori_n89_), .B(ori_ori_n102_), .C(ori_ori_n95_), .Y(ori_ori_n109_));
  NAi31      o081(.An(e), .B(f), .C(b), .Y(ori_ori_n110_));
  NOi21      o082(.An(k), .B(m), .Y(ori_ori_n111_));
  NAi31      o083(.An(d), .B(f), .C(c), .Y(ori_ori_n112_));
  NAi31      o084(.An(e), .B(f), .C(c), .Y(ori_ori_n113_));
  NA2        o085(.A(ori_ori_n113_), .B(ori_ori_n112_), .Y(ori_ori_n114_));
  NA2        o086(.A(j), .B(h), .Y(ori_ori_n115_));
  OR3        o087(.A(n), .B(m), .C(k), .Y(ori_ori_n116_));
  NO2        o088(.A(ori_ori_n116_), .B(ori_ori_n115_), .Y(ori_ori_n117_));
  NAi32      o089(.An(m), .Bn(k), .C(n), .Y(ori_ori_n118_));
  NA2        o090(.A(ori_ori_n117_), .B(ori_ori_n114_), .Y(ori_ori_n119_));
  NO2        o091(.A(n), .B(m), .Y(ori_ori_n120_));
  NA2        o092(.A(ori_ori_n120_), .B(ori_ori_n39_), .Y(ori_ori_n121_));
  NAi21      o093(.An(f), .B(e), .Y(ori_ori_n122_));
  NA2        o094(.A(d), .B(c), .Y(ori_ori_n123_));
  NO2        o095(.A(ori_ori_n123_), .B(ori_ori_n122_), .Y(ori_ori_n124_));
  NOi21      o096(.An(ori_ori_n124_), .B(ori_ori_n121_), .Y(ori_ori_n125_));
  NAi31      o097(.An(m), .B(n), .C(b), .Y(ori_ori_n126_));
  NA2        o098(.A(k), .B(i), .Y(ori_ori_n127_));
  NAi21      o099(.An(h), .B(f), .Y(ori_ori_n128_));
  NO2        o100(.A(ori_ori_n128_), .B(ori_ori_n127_), .Y(ori_ori_n129_));
  NO2        o101(.A(ori_ori_n126_), .B(ori_ori_n107_), .Y(ori_ori_n130_));
  NA2        o102(.A(ori_ori_n130_), .B(ori_ori_n129_), .Y(ori_ori_n131_));
  NOi32      o103(.An(f), .Bn(c), .C(d), .Y(ori_ori_n132_));
  NOi32      o104(.An(f), .Bn(c), .C(e), .Y(ori_ori_n133_));
  NO2        o105(.A(ori_ori_n133_), .B(ori_ori_n132_), .Y(ori_ori_n134_));
  NO3        o106(.A(n), .B(m), .C(j), .Y(ori_ori_n135_));
  NA2        o107(.A(ori_ori_n135_), .B(ori_ori_n80_), .Y(ori_ori_n136_));
  AO210      o108(.A0(ori_ori_n136_), .A1(ori_ori_n121_), .B0(ori_ori_n134_), .Y(ori_ori_n137_));
  NAi41      o109(.An(ori_ori_n125_), .B(ori_ori_n137_), .C(ori_ori_n131_), .D(ori_ori_n119_), .Y(ori_ori_n138_));
  OR2        o110(.A(ori_ori_n138_), .B(ori_ori_n109_), .Y(ori_ori_n139_));
  NO4        o111(.A(ori_ori_n139_), .B(ori_ori_n85_), .C(ori_ori_n58_), .D(ori_ori_n44_), .Y(ori_ori_n140_));
  NAi31      o112(.An(n), .B(h), .C(o), .Y(ori_ori_n141_));
  NOi32      o113(.An(m), .Bn(k), .C(l), .Y(ori_ori_n142_));
  NA3        o114(.A(ori_ori_n142_), .B(ori_ori_n62_), .C(o), .Y(ori_ori_n143_));
  NO2        o115(.A(ori_ori_n143_), .B(n), .Y(ori_ori_n144_));
  NOi21      o116(.An(k), .B(j), .Y(ori_ori_n145_));
  NA4        o117(.A(ori_ori_n145_), .B(ori_ori_n79_), .C(i), .D(o), .Y(ori_ori_n146_));
  INV        o118(.A(ori_ori_n146_), .Y(ori_ori_n147_));
  NAi41      o119(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n148_));
  INV        o120(.A(f), .Y(ori_ori_n149_));
  INV        o121(.A(o), .Y(ori_ori_n150_));
  NOi31      o122(.An(i), .B(j), .C(h), .Y(ori_ori_n151_));
  NOi21      o123(.An(l), .B(m), .Y(ori_ori_n152_));
  NA2        o124(.A(ori_ori_n152_), .B(ori_ori_n151_), .Y(ori_ori_n153_));
  NO2        o125(.A(ori_ori_n153_), .B(ori_ori_n149_), .Y(ori_ori_n154_));
  NOi21      o126(.An(n), .B(m), .Y(ori_ori_n155_));
  OR2        o127(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n156_));
  NAi21      o128(.An(j), .B(h), .Y(ori_ori_n157_));
  XN2        o129(.A(i), .B(h), .Y(ori_ori_n158_));
  NA2        o130(.A(ori_ori_n158_), .B(ori_ori_n157_), .Y(ori_ori_n159_));
  NOi31      o131(.An(k), .B(n), .C(m), .Y(ori_ori_n160_));
  NOi31      o132(.An(ori_ori_n160_), .B(ori_ori_n123_), .C(ori_ori_n122_), .Y(ori_ori_n161_));
  NA2        o133(.A(ori_ori_n161_), .B(ori_ori_n159_), .Y(ori_ori_n162_));
  NAi31      o134(.An(f), .B(e), .C(c), .Y(ori_ori_n163_));
  NO4        o135(.A(ori_ori_n163_), .B(ori_ori_n116_), .C(ori_ori_n115_), .D(ori_ori_n47_), .Y(ori_ori_n164_));
  NA3        o136(.A(e), .B(c), .C(b), .Y(ori_ori_n165_));
  NAi32      o137(.An(m), .Bn(i), .C(k), .Y(ori_ori_n166_));
  INV        o138(.A(ori_ori_n164_), .Y(ori_ori_n167_));
  NAi21      o139(.An(n), .B(a), .Y(ori_ori_n168_));
  NO2        o140(.A(ori_ori_n168_), .B(ori_ori_n103_), .Y(ori_ori_n169_));
  NAi41      o141(.An(o), .B(m), .C(k), .D(h), .Y(ori_ori_n170_));
  NO2        o142(.A(ori_ori_n170_), .B(e), .Y(ori_ori_n171_));
  NA2        o143(.A(ori_ori_n171_), .B(ori_ori_n169_), .Y(ori_ori_n172_));
  AN4        o144(.A(ori_ori_n172_), .B(ori_ori_n167_), .C(ori_ori_n162_), .D(ori_ori_n156_), .Y(ori_ori_n173_));
  OR2        o145(.A(h), .B(o), .Y(ori_ori_n174_));
  NO2        o146(.A(ori_ori_n174_), .B(ori_ori_n70_), .Y(ori_ori_n175_));
  NA2        o147(.A(ori_ori_n175_), .B(f), .Y(ori_ori_n176_));
  NAi41      o148(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n177_));
  NO2        o149(.A(ori_ori_n177_), .B(ori_ori_n149_), .Y(ori_ori_n178_));
  NA2        o150(.A(ori_ori_n111_), .B(ori_ori_n75_), .Y(ori_ori_n179_));
  NAi21      o151(.An(ori_ori_n179_), .B(ori_ori_n178_), .Y(ori_ori_n180_));
  NO2        o152(.A(n), .B(a), .Y(ori_ori_n181_));
  NAi31      o153(.An(ori_ori_n170_), .B(ori_ori_n181_), .C(ori_ori_n71_), .Y(ori_ori_n182_));
  AN2        o154(.A(ori_ori_n182_), .B(ori_ori_n180_), .Y(ori_ori_n183_));
  NAi21      o155(.An(h), .B(i), .Y(ori_ori_n184_));
  NA2        o156(.A(ori_ori_n120_), .B(k), .Y(ori_ori_n185_));
  NO2        o157(.A(ori_ori_n185_), .B(ori_ori_n184_), .Y(ori_ori_n186_));
  NA2        o158(.A(ori_ori_n183_), .B(ori_ori_n176_), .Y(ori_ori_n187_));
  NOi21      o159(.An(o), .B(e), .Y(ori_ori_n188_));
  NOi21      o160(.An(ori_ori_n173_), .B(ori_ori_n187_), .Y(ori_ori_n189_));
  NA3        o161(.A(ori_ori_n47_), .B(c), .C(b), .Y(ori_ori_n190_));
  NO2        o162(.A(ori_ori_n179_), .B(f), .Y(ori_ori_n191_));
  NAi31      o163(.An(o), .B(k), .C(h), .Y(ori_ori_n192_));
  NA2        o164(.A(ori_ori_n111_), .B(h), .Y(ori_ori_n193_));
  NA3        o165(.A(e), .B(c), .C(b), .Y(ori_ori_n194_));
  NAi32      o166(.An(j), .Bn(h), .C(i), .Y(ori_ori_n195_));
  NAi21      o167(.An(m), .B(l), .Y(ori_ori_n196_));
  NA2        o168(.A(h), .B(o), .Y(ori_ori_n197_));
  NO2        o169(.A(ori_ori_n101_), .B(d), .Y(ori_ori_n198_));
  NO2        o170(.A(ori_ori_n73_), .B(ori_ori_n70_), .Y(ori_ori_n199_));
  NAi32      o171(.An(n), .Bn(m), .C(l), .Y(ori_ori_n200_));
  NO2        o172(.A(ori_ori_n200_), .B(ori_ori_n195_), .Y(ori_ori_n201_));
  NA2        o173(.A(ori_ori_n201_), .B(ori_ori_n124_), .Y(ori_ori_n202_));
  NA2        o174(.A(ori_ori_n186_), .B(ori_ori_n133_), .Y(ori_ori_n203_));
  NAi21      o175(.An(m), .B(k), .Y(ori_ori_n204_));
  NO2        o176(.A(ori_ori_n158_), .B(ori_ori_n204_), .Y(ori_ori_n205_));
  NAi41      o177(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n206_));
  NO2        o178(.A(ori_ori_n206_), .B(ori_ori_n106_), .Y(ori_ori_n207_));
  NA2        o179(.A(ori_ori_n207_), .B(ori_ori_n205_), .Y(ori_ori_n208_));
  NA2        o180(.A(e), .B(c), .Y(ori_ori_n209_));
  NO3        o181(.A(ori_ori_n209_), .B(n), .C(d), .Y(ori_ori_n210_));
  NOi21      o182(.An(f), .B(h), .Y(ori_ori_n211_));
  NA2        o183(.A(ori_ori_n211_), .B(k), .Y(ori_ori_n212_));
  NO2        o184(.A(ori_ori_n212_), .B(ori_ori_n150_), .Y(ori_ori_n213_));
  NAi31      o185(.An(d), .B(e), .C(b), .Y(ori_ori_n214_));
  NO2        o186(.A(ori_ori_n91_), .B(ori_ori_n214_), .Y(ori_ori_n215_));
  NA2        o187(.A(ori_ori_n215_), .B(ori_ori_n213_), .Y(ori_ori_n216_));
  NA3        o188(.A(ori_ori_n216_), .B(ori_ori_n208_), .C(ori_ori_n203_), .Y(ori_ori_n217_));
  NO3        o189(.A(ori_ori_n206_), .B(ori_ori_n56_), .C(ori_ori_n50_), .Y(ori_ori_n218_));
  NA2        o190(.A(ori_ori_n181_), .B(ori_ori_n71_), .Y(ori_ori_n219_));
  OR2        o191(.A(ori_ori_n219_), .B(ori_ori_n143_), .Y(ori_ori_n220_));
  NOi31      o192(.An(l), .B(n), .C(m), .Y(ori_ori_n221_));
  NA2        o193(.A(ori_ori_n221_), .B(ori_ori_n151_), .Y(ori_ori_n222_));
  NO2        o194(.A(ori_ori_n222_), .B(ori_ori_n134_), .Y(ori_ori_n223_));
  NAi32      o195(.An(ori_ori_n223_), .Bn(ori_ori_n218_), .C(ori_ori_n220_), .Y(ori_ori_n224_));
  NAi32      o196(.An(m), .Bn(j), .C(k), .Y(ori_ori_n225_));
  NAi41      o197(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n226_));
  NA2        o198(.A(ori_ori_n148_), .B(ori_ori_n226_), .Y(ori_ori_n227_));
  NOi31      o199(.An(j), .B(m), .C(k), .Y(ori_ori_n228_));
  NO2        o200(.A(ori_ori_n86_), .B(ori_ori_n228_), .Y(ori_ori_n229_));
  AN3        o201(.A(h), .B(o), .C(f), .Y(ori_ori_n230_));
  NAi31      o202(.An(ori_ori_n229_), .B(ori_ori_n230_), .C(ori_ori_n227_), .Y(ori_ori_n231_));
  INV        o203(.A(m), .Y(ori_ori_n232_));
  NAi32      o204(.An(ori_ori_n232_), .Bn(ori_ori_n141_), .C(ori_ori_n198_), .Y(ori_ori_n233_));
  NO2        o205(.A(ori_ori_n196_), .B(ori_ori_n195_), .Y(ori_ori_n234_));
  NO2        o206(.A(ori_ori_n153_), .B(o), .Y(ori_ori_n235_));
  AOI220     o207(.A0(f), .A1(ori_ori_n235_), .B0(ori_ori_n178_), .B1(ori_ori_n234_), .Y(ori_ori_n236_));
  NA3        o208(.A(ori_ori_n236_), .B(ori_ori_n233_), .C(ori_ori_n231_), .Y(ori_ori_n237_));
  NA3        o209(.A(h), .B(o), .C(f), .Y(ori_ori_n238_));
  NO2        o210(.A(ori_ori_n238_), .B(ori_ori_n53_), .Y(ori_ori_n239_));
  NA2        o211(.A(e), .B(ori_ori_n239_), .Y(ori_ori_n240_));
  NOi32      o212(.An(j), .Bn(o), .C(i), .Y(ori_ori_n241_));
  NOi32      o213(.An(e), .Bn(b), .C(a), .Y(ori_ori_n242_));
  INV        o214(.A(ori_ori_n204_), .Y(ori_ori_n243_));
  NO3        o215(.A(ori_ori_n206_), .B(ori_ori_n50_), .C(ori_ori_n150_), .Y(ori_ori_n244_));
  INV        o216(.A(ori_ori_n146_), .Y(ori_ori_n245_));
  AOI220     o217(.A0(ori_ori_n245_), .A1(ori_ori_n242_), .B0(ori_ori_n244_), .B1(ori_ori_n243_), .Y(ori_ori_n246_));
  NA4        o218(.A(ori_ori_n142_), .B(ori_ori_n62_), .C(o), .D(ori_ori_n149_), .Y(ori_ori_n247_));
  NA2        o219(.A(ori_ori_n40_), .B(ori_ori_n79_), .Y(ori_ori_n248_));
  NA2        o220(.A(ori_ori_n246_), .B(ori_ori_n240_), .Y(ori_ori_n249_));
  NO4        o221(.A(ori_ori_n249_), .B(ori_ori_n237_), .C(ori_ori_n224_), .D(ori_ori_n217_), .Y(ori_ori_n250_));
  NA4        o222(.A(ori_ori_n250_), .B(ori_ori_n202_), .C(ori_ori_n189_), .D(ori_ori_n140_), .Y(ori10));
  NA3        o223(.A(m), .B(k), .C(i), .Y(ori_ori_n252_));
  NOi21      o224(.An(e), .B(f), .Y(ori_ori_n253_));
  NO3        o225(.A(ori_ori_n107_), .B(n), .C(ori_ori_n76_), .Y(ori_ori_n254_));
  NOi32      o226(.An(k), .Bn(h), .C(j), .Y(ori_ori_n255_));
  NA2        o227(.A(ori_ori_n255_), .B(ori_ori_n155_), .Y(ori_ori_n256_));
  AN2        o228(.A(j), .B(h), .Y(ori_ori_n257_));
  NO3        o229(.A(n), .B(m), .C(k), .Y(ori_ori_n258_));
  NA2        o230(.A(ori_ori_n258_), .B(ori_ori_n257_), .Y(ori_ori_n259_));
  NO3        o231(.A(ori_ori_n259_), .B(ori_ori_n107_), .C(ori_ori_n149_), .Y(ori_ori_n260_));
  OR2        o232(.A(m), .B(k), .Y(ori_ori_n261_));
  NO2        o233(.A(ori_ori_n115_), .B(ori_ori_n261_), .Y(ori_ori_n262_));
  NA4        o234(.A(n), .B(f), .C(c), .D(ori_ori_n81_), .Y(ori_ori_n263_));
  NOi21      o235(.An(ori_ori_n262_), .B(ori_ori_n263_), .Y(ori_ori_n264_));
  NOi32      o236(.An(d), .Bn(a), .C(c), .Y(ori_ori_n265_));
  NA2        o237(.A(ori_ori_n265_), .B(ori_ori_n122_), .Y(ori_ori_n266_));
  NO2        o238(.A(ori_ori_n264_), .B(ori_ori_n260_), .Y(ori_ori_n267_));
  NO2        o239(.A(ori_ori_n263_), .B(ori_ori_n196_), .Y(ori_ori_n268_));
  NOi32      o240(.An(f), .Bn(d), .C(c), .Y(ori_ori_n269_));
  INV        o241(.A(ori_ori_n267_), .Y(ori_ori_n270_));
  NA2        o242(.A(ori_ori_n181_), .B(b), .Y(ori_ori_n271_));
  INV        o243(.A(e), .Y(ori_ori_n272_));
  NA3        o244(.A(m), .B(o), .C(e), .Y(ori_ori_n273_));
  AN3        o245(.A(h), .B(o), .C(e), .Y(ori_ori_n274_));
  NO2        o246(.A(ori_ori_n273_), .B(ori_ori_n271_), .Y(ori_ori_n275_));
  NA3        o247(.A(ori_ori_n265_), .B(ori_ori_n122_), .C(ori_ori_n59_), .Y(ori_ori_n276_));
  NAi31      o248(.An(b), .B(c), .C(a), .Y(ori_ori_n277_));
  NO2        o249(.A(ori_ori_n277_), .B(n), .Y(ori_ori_n278_));
  NA2        o250(.A(ori_ori_n40_), .B(m), .Y(ori_ori_n279_));
  NO2        o251(.A(ori_ori_n279_), .B(ori_ori_n104_), .Y(ori_ori_n280_));
  NA2        o252(.A(ori_ori_n280_), .B(ori_ori_n278_), .Y(ori_ori_n281_));
  INV        o253(.A(ori_ori_n281_), .Y(ori_ori_n282_));
  NO3        o254(.A(ori_ori_n282_), .B(ori_ori_n275_), .C(ori_ori_n270_), .Y(ori_ori_n283_));
  NA2        o255(.A(i), .B(o), .Y(ori_ori_n284_));
  NA3        o256(.A(i), .B(o), .C(f), .Y(ori_ori_n285_));
  OR2        o257(.A(n), .B(m), .Y(ori_ori_n286_));
  NO2        o258(.A(ori_ori_n286_), .B(ori_ori_n108_), .Y(ori_ori_n287_));
  NO2        o259(.A(ori_ori_n123_), .B(ori_ori_n104_), .Y(ori_ori_n288_));
  OAI210     o260(.A0(ori_ori_n287_), .A1(ori_ori_n117_), .B0(ori_ori_n288_), .Y(ori_ori_n289_));
  INV        o261(.A(ori_ori_n248_), .Y(ori_ori_n290_));
  NA2        o262(.A(ori_ori_n290_), .B(ori_ori_n242_), .Y(ori_ori_n291_));
  NO2        o263(.A(ori_ori_n277_), .B(ori_ori_n38_), .Y(ori_ori_n292_));
  NAi21      o264(.An(k), .B(j), .Y(ori_ori_n293_));
  NA2        o265(.A(ori_ori_n184_), .B(ori_ori_n293_), .Y(ori_ori_n294_));
  NA3        o266(.A(ori_ori_n294_), .B(o), .C(ori_ori_n292_), .Y(ori_ori_n295_));
  NAi21      o267(.An(e), .B(d), .Y(ori_ori_n296_));
  INV        o268(.A(ori_ori_n296_), .Y(ori_ori_n297_));
  NO2        o269(.A(ori_ori_n185_), .B(ori_ori_n149_), .Y(ori_ori_n298_));
  NA3        o270(.A(ori_ori_n298_), .B(ori_ori_n297_), .C(ori_ori_n159_), .Y(ori_ori_n299_));
  NA4        o271(.A(ori_ori_n299_), .B(ori_ori_n295_), .C(ori_ori_n291_), .D(ori_ori_n289_), .Y(ori_ori_n300_));
  NO2        o272(.A(ori_ori_n222_), .B(ori_ori_n149_), .Y(ori_ori_n301_));
  NA2        o273(.A(ori_ori_n301_), .B(ori_ori_n297_), .Y(ori_ori_n302_));
  NOi31      o274(.An(n), .B(m), .C(k), .Y(ori_ori_n303_));
  AOI220     o275(.A0(ori_ori_n303_), .A1(ori_ori_n257_), .B0(ori_ori_n155_), .B1(ori_ori_n39_), .Y(ori_ori_n304_));
  NAi31      o276(.An(o), .B(f), .C(c), .Y(ori_ori_n305_));
  OR2        o277(.A(ori_ori_n305_), .B(ori_ori_n304_), .Y(ori_ori_n306_));
  NA3        o278(.A(ori_ori_n306_), .B(ori_ori_n302_), .C(ori_ori_n202_), .Y(ori_ori_n307_));
  NO2        o279(.A(ori_ori_n307_), .B(ori_ori_n300_), .Y(ori_ori_n308_));
  NOi32      o280(.An(c), .Bn(a), .C(b), .Y(ori_ori_n309_));
  NA2        o281(.A(ori_ori_n309_), .B(ori_ori_n79_), .Y(ori_ori_n310_));
  INV        o282(.A(ori_ori_n192_), .Y(ori_ori_n311_));
  AN2        o283(.A(e), .B(d), .Y(ori_ori_n312_));
  NA2        o284(.A(ori_ori_n312_), .B(ori_ori_n311_), .Y(ori_ori_n313_));
  NO2        o285(.A(ori_ori_n48_), .B(e), .Y(ori_ori_n314_));
  NA2        o286(.A(ori_ori_n52_), .B(ori_ori_n314_), .Y(ori_ori_n315_));
  AOI210     o287(.A0(ori_ori_n315_), .A1(ori_ori_n313_), .B0(ori_ori_n310_), .Y(ori_ori_n316_));
  NO2        o288(.A(ori_ori_n147_), .B(ori_ori_n144_), .Y(ori_ori_n317_));
  NA3        o289(.A(e), .B(d), .C(c), .Y(ori_ori_n318_));
  BUFFER     o290(.A(ori_ori_n318_), .Y(ori_ori_n319_));
  NO2        o291(.A(ori_ori_n276_), .B(ori_ori_n143_), .Y(ori_ori_n320_));
  NOi21      o292(.An(ori_ori_n319_), .B(ori_ori_n320_), .Y(ori_ori_n321_));
  NO2        o293(.A(ori_ori_n317_), .B(ori_ori_n321_), .Y(ori_ori_n322_));
  NO4        o294(.A(ori_ori_n128_), .B(ori_ori_n70_), .C(ori_ori_n45_), .D(b), .Y(ori_ori_n323_));
  NA2        o295(.A(l), .B(k), .Y(ori_ori_n324_));
  AOI210     o296(.A0(ori_ori_n166_), .A1(ori_ori_n225_), .B0(ori_ori_n59_), .Y(ori_ori_n325_));
  INV        o297(.A(ori_ori_n87_), .Y(ori_ori_n326_));
  INV        o298(.A(ori_ori_n87_), .Y(ori_ori_n327_));
  NO4        o299(.A(ori_ori_n327_), .B(ori_ori_n323_), .C(ori_ori_n322_), .D(ori_ori_n316_), .Y(ori_ori_n328_));
  INV        o300(.A(e), .Y(ori_ori_n329_));
  INV        o301(.A(ori_ori_n128_), .Y(ori_ori_n330_));
  NAi31      o302(.An(j), .B(l), .C(i), .Y(ori_ori_n331_));
  OAI210     o303(.A0(ori_ori_n331_), .A1(ori_ori_n91_), .B0(ori_ori_n70_), .Y(ori_ori_n332_));
  NA3        o304(.A(ori_ori_n332_), .B(ori_ori_n330_), .C(ori_ori_n329_), .Y(ori_ori_n333_));
  NO2        o305(.A(ori_ori_n266_), .B(ori_ori_n248_), .Y(ori_ori_n334_));
  NO3        o306(.A(ori_ori_n334_), .B(ori_ori_n125_), .C(ori_ori_n199_), .Y(ori_ori_n335_));
  NA3        o307(.A(ori_ori_n335_), .B(ori_ori_n333_), .C(ori_ori_n173_), .Y(ori_ori_n336_));
  OAI210     o308(.A0(ori_ori_n88_), .A1(ori_ori_n86_), .B0(n), .Y(ori_ori_n337_));
  XO2        o309(.A(i), .B(h), .Y(ori_ori_n338_));
  NA3        o310(.A(ori_ori_n338_), .B(ori_ori_n111_), .C(n), .Y(ori_ori_n339_));
  NA3        o311(.A(ori_ori_n339_), .B(ori_ori_n304_), .C(ori_ori_n256_), .Y(ori_ori_n340_));
  AN2        o312(.A(ori_ori_n340_), .B(ori_ori_n314_), .Y(ori_ori_n341_));
  NAi31      o313(.An(c), .B(f), .C(d), .Y(ori_ori_n342_));
  BUFFER     o314(.A(ori_ori_n57_), .Y(ori_ori_n343_));
  NA2        o315(.A(ori_ori_n160_), .B(ori_ori_n75_), .Y(ori_ori_n344_));
  AOI210     o316(.A0(ori_ori_n344_), .A1(ori_ori_n121_), .B0(ori_ori_n342_), .Y(ori_ori_n345_));
  INV        o317(.A(ori_ori_n345_), .Y(ori_ori_n346_));
  NA3        o318(.A(ori_ori_n31_), .B(m), .C(f), .Y(ori_ori_n347_));
  NA2        o319(.A(ori_ori_n346_), .B(ori_ori_n343_), .Y(ori_ori_n348_));
  NO3        o320(.A(ori_ori_n348_), .B(ori_ori_n341_), .C(ori_ori_n336_), .Y(ori_ori_n349_));
  NA4        o321(.A(ori_ori_n349_), .B(ori_ori_n328_), .C(ori_ori_n308_), .D(ori_ori_n283_), .Y(ori11));
  NAi31      o322(.An(i), .B(m), .C(l), .Y(ori_ori_n351_));
  NA2        o323(.A(m), .B(k), .Y(ori_ori_n352_));
  NOi32      o324(.An(e), .Bn(b), .C(f), .Y(ori_ori_n353_));
  NA2        o325(.A(ori_ori_n36_), .B(j), .Y(ori_ori_n354_));
  NAi31      o326(.An(d), .B(e), .C(a), .Y(ori_ori_n355_));
  NO2        o327(.A(ori_ori_n355_), .B(n), .Y(ori_ori_n356_));
  NA2        o328(.A(j), .B(i), .Y(ori_ori_n357_));
  NAi31      o329(.An(n), .B(m), .C(k), .Y(ori_ori_n358_));
  NO3        o330(.A(n), .B(d), .C(ori_ori_n81_), .Y(ori_ori_n359_));
  OR2        o331(.A(n), .B(c), .Y(ori_ori_n360_));
  NO2        o332(.A(ori_ori_n360_), .B(ori_ori_n105_), .Y(ori_ori_n361_));
  NO2        o333(.A(ori_ori_n192_), .B(ori_ori_n38_), .Y(ori_ori_n362_));
  NA2        o334(.A(ori_ori_n97_), .B(ori_ori_n30_), .Y(ori_ori_n363_));
  OAI220     o335(.A0(ori_ori_n363_), .A1(m), .B0(ori_ori_n354_), .B1(ori_ori_n166_), .Y(ori_ori_n364_));
  NOi41      o336(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n365_));
  NAi32      o337(.An(e), .Bn(b), .C(c), .Y(ori_ori_n366_));
  OR2        o338(.A(ori_ori_n366_), .B(ori_ori_n59_), .Y(ori_ori_n367_));
  AN2        o339(.A(ori_ori_n226_), .B(ori_ori_n206_), .Y(ori_ori_n368_));
  NA2        o340(.A(ori_ori_n368_), .B(ori_ori_n367_), .Y(ori_ori_n369_));
  OA210      o341(.A0(ori_ori_n369_), .A1(ori_ori_n365_), .B0(ori_ori_n364_), .Y(ori_ori_n370_));
  NAi32      o342(.An(d), .Bn(a), .C(b), .Y(ori_ori_n371_));
  NO2        o343(.A(ori_ori_n371_), .B(ori_ori_n38_), .Y(ori_ori_n372_));
  NO3        o344(.A(ori_ori_n118_), .B(ori_ori_n115_), .C(o), .Y(ori_ori_n373_));
  AOI220     o345(.A0(ori_ori_n373_), .A1(b), .B0(ori_ori_n830_), .B1(ori_ori_n372_), .Y(ori_ori_n374_));
  INV        o346(.A(ori_ori_n374_), .Y(ori_ori_n375_));
  AN3        o347(.A(j), .B(h), .C(o), .Y(ori_ori_n376_));
  NO2        o348(.A(ori_ori_n103_), .B(c), .Y(ori_ori_n377_));
  NA3        o349(.A(ori_ori_n377_), .B(ori_ori_n376_), .C(ori_ori_n303_), .Y(ori_ori_n378_));
  NA3        o350(.A(f), .B(d), .C(b), .Y(ori_ori_n379_));
  NO4        o351(.A(ori_ori_n379_), .B(ori_ori_n118_), .C(ori_ori_n115_), .D(o), .Y(ori_ori_n380_));
  INV        o352(.A(ori_ori_n378_), .Y(ori_ori_n381_));
  NO3        o353(.A(ori_ori_n381_), .B(ori_ori_n375_), .C(ori_ori_n370_), .Y(ori_ori_n382_));
  NAi41      o354(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n383_));
  OAI210     o355(.A0(ori_ori_n355_), .A1(n), .B0(ori_ori_n383_), .Y(ori_ori_n384_));
  NAi31      o356(.An(h), .B(o), .C(f), .Y(ori_ori_n385_));
  NAi31      o357(.An(f), .B(h), .C(o), .Y(ori_ori_n386_));
  NO2        o358(.A(n), .B(c), .Y(ori_ori_n387_));
  NA2        o359(.A(ori_ori_n305_), .B(ori_ori_n163_), .Y(ori_ori_n388_));
  NA3        o360(.A(ori_ori_n365_), .B(ori_ori_n228_), .C(ori_ori_n36_), .Y(ori_ori_n389_));
  NOi32      o361(.An(e), .Bn(c), .C(f), .Y(ori_ori_n390_));
  INV        o362(.A(ori_ori_n148_), .Y(ori_ori_n391_));
  AOI220     o363(.A0(ori_ori_n391_), .A1(ori_ori_n262_), .B0(ori_ori_n390_), .B1(ori_ori_n117_), .Y(ori_ori_n392_));
  NA3        o364(.A(ori_ori_n392_), .B(ori_ori_n389_), .C(ori_ori_n119_), .Y(ori_ori_n393_));
  NA2        o365(.A(ori_ori_n75_), .B(m), .Y(ori_ori_n394_));
  INV        o366(.A(ori_ori_n242_), .Y(ori_ori_n395_));
  NO2        o367(.A(ori_ori_n395_), .B(n), .Y(ori_ori_n396_));
  NAi31      o368(.An(ori_ori_n394_), .B(ori_ori_n396_), .C(o), .Y(ori_ori_n397_));
  NO2        o369(.A(ori_ori_n354_), .B(ori_ori_n118_), .Y(ori_ori_n398_));
  NA3        o370(.A(ori_ori_n366_), .B(ori_ori_n190_), .C(ori_ori_n101_), .Y(ori_ori_n399_));
  NA2        o371(.A(ori_ori_n338_), .B(ori_ori_n111_), .Y(ori_ori_n400_));
  NO3        o372(.A(ori_ori_n263_), .B(ori_ori_n400_), .C(ori_ori_n62_), .Y(ori_ori_n401_));
  AOI210     o373(.A0(ori_ori_n399_), .A1(ori_ori_n398_), .B0(ori_ori_n401_), .Y(ori_ori_n402_));
  AN3        o374(.A(f), .B(d), .C(b), .Y(ori_ori_n403_));
  NAi31      o375(.An(m), .B(n), .C(k), .Y(ori_ori_n404_));
  NA3        o376(.A(ori_ori_n182_), .B(ori_ori_n402_), .C(ori_ori_n397_), .Y(ori_ori_n405_));
  NO2        o377(.A(ori_ori_n405_), .B(ori_ori_n393_), .Y(ori_ori_n406_));
  NA2        o378(.A(ori_ori_n254_), .B(h), .Y(ori_ori_n407_));
  NAi31      o379(.An(o), .B(h), .C(f), .Y(ori_ori_n408_));
  OA210      o380(.A0(ori_ori_n355_), .A1(n), .B0(ori_ori_n383_), .Y(ori_ori_n409_));
  NO2        o381(.A(ori_ori_n407_), .B(ori_ori_n352_), .Y(ori_ori_n410_));
  NO3        o382(.A(o), .B(ori_ori_n149_), .C(ori_ori_n45_), .Y(ori_ori_n411_));
  NO2        o383(.A(ori_ori_n344_), .B(ori_ori_n62_), .Y(ori_ori_n412_));
  OAI210     o384(.A0(ori_ori_n412_), .A1(ori_ori_n262_), .B0(ori_ori_n411_), .Y(ori_ori_n413_));
  AOI210     o385(.A0(ori_ori_n371_), .A1(ori_ori_n277_), .B0(ori_ori_n38_), .Y(ori_ori_n414_));
  NA2        o386(.A(ori_ori_n822_), .B(ori_ori_n414_), .Y(ori_ori_n415_));
  NA2        o387(.A(ori_ori_n415_), .B(ori_ori_n413_), .Y(ori_ori_n416_));
  INV        o388(.A(ori_ori_n215_), .Y(ori_ori_n417_));
  OR2        o389(.A(ori_ori_n829_), .B(ori_ori_n363_), .Y(ori_ori_n418_));
  OAI210     o390(.A0(ori_ori_n417_), .A1(ori_ori_n820_), .B0(ori_ori_n418_), .Y(ori_ori_n419_));
  NO2        o391(.A(ori_ori_n269_), .B(ori_ori_n133_), .Y(ori_ori_n420_));
  NO3        o392(.A(ori_ori_n305_), .B(ori_ori_n115_), .C(i), .Y(ori_ori_n421_));
  NA2        o393(.A(ori_ori_n309_), .B(ori_ori_n59_), .Y(ori_ori_n422_));
  NO3        o394(.A(ori_ori_n352_), .B(ori_ori_n422_), .C(ori_ori_n90_), .Y(ori_ori_n423_));
  INV        o395(.A(ori_ori_n423_), .Y(ori_ori_n424_));
  NA2        o396(.A(ori_ori_n424_), .B(ori_ori_n267_), .Y(ori_ori_n425_));
  NO4        o397(.A(ori_ori_n425_), .B(ori_ori_n419_), .C(ori_ori_n416_), .D(ori_ori_n410_), .Y(ori_ori_n426_));
  NA4        o398(.A(ori_ori_n426_), .B(ori_ori_n406_), .C(ori_ori_n180_), .D(ori_ori_n382_), .Y(ori08));
  NO2        o399(.A(k), .B(h), .Y(ori_ori_n428_));
  AO210      o400(.A0(ori_ori_n184_), .A1(ori_ori_n293_), .B0(ori_ori_n428_), .Y(ori_ori_n429_));
  NO2        o401(.A(ori_ori_n429_), .B(ori_ori_n196_), .Y(ori_ori_n430_));
  NA2        o402(.A(ori_ori_n390_), .B(ori_ori_n59_), .Y(ori_ori_n431_));
  NA2        o403(.A(ori_ori_n431_), .B(ori_ori_n305_), .Y(ori_ori_n432_));
  NA2        o404(.A(ori_ori_n432_), .B(ori_ori_n430_), .Y(ori_ori_n433_));
  NA2        o405(.A(ori_ori_n59_), .B(ori_ori_n76_), .Y(ori_ori_n434_));
  NO2        o406(.A(ori_ori_n434_), .B(ori_ori_n46_), .Y(ori_ori_n435_));
  NO2        o407(.A(ori_ori_n252_), .B(j), .Y(ori_ori_n436_));
  NA2        o408(.A(ori_ori_n436_), .B(ori_ori_n435_), .Y(ori_ori_n437_));
  AOI210     o409(.A0(ori_ori_n379_), .A1(ori_ori_n110_), .B0(ori_ori_n59_), .Y(ori_ori_n438_));
  NA4        o410(.A(ori_ori_n152_), .B(ori_ori_n97_), .C(ori_ori_n35_), .D(h), .Y(ori_ori_n439_));
  NA4        o411(.A(k), .B(ori_ori_n75_), .C(ori_ori_n51_), .D(ori_ori_n150_), .Y(ori_ori_n440_));
  OAI210     o412(.A0(ori_ori_n439_), .A1(o), .B0(ori_ori_n440_), .Y(ori_ori_n441_));
  NA2        o413(.A(ori_ori_n441_), .B(ori_ori_n438_), .Y(ori_ori_n442_));
  NA4        o414(.A(ori_ori_n442_), .B(ori_ori_n437_), .C(ori_ori_n433_), .D(ori_ori_n236_), .Y(ori_ori_n443_));
  NO4        o415(.A(ori_ori_n115_), .B(ori_ori_n261_), .C(ori_ori_n78_), .D(o), .Y(ori_ori_n444_));
  NA2        o416(.A(ori_ori_n444_), .B(e), .Y(ori_ori_n445_));
  NO2        o417(.A(ori_ori_n32_), .B(ori_ori_n149_), .Y(ori_ori_n446_));
  NA2        o418(.A(ori_ori_n391_), .B(ori_ori_n234_), .Y(ori_ori_n447_));
  NA2        o419(.A(ori_ori_n447_), .B(ori_ori_n445_), .Y(ori_ori_n448_));
  NO3        o420(.A(ori_ori_n204_), .B(ori_ori_n90_), .C(j), .Y(ori_ori_n449_));
  NAi21      o421(.An(ori_ori_n449_), .B(ori_ori_n440_), .Y(ori_ori_n450_));
  NA2        o422(.A(ori_ori_n429_), .B(ori_ori_n94_), .Y(ori_ori_n451_));
  AOI220     o423(.A0(ori_ori_n451_), .A1(ori_ori_n268_), .B0(ori_ori_n450_), .B1(ori_ori_n54_), .Y(ori_ori_n452_));
  INV        o424(.A(ori_ori_n452_), .Y(ori_ori_n453_));
  NA3        o425(.A(m), .B(l), .C(k), .Y(ori_ori_n454_));
  NO3        o426(.A(ori_ori_n453_), .B(ori_ori_n448_), .C(ori_ori_n443_), .Y(ori_ori_n455_));
  NA2        o427(.A(ori_ori_n391_), .B(ori_ori_n262_), .Y(ori_ori_n456_));
  INV        o428(.A(ori_ori_n334_), .Y(ori_ori_n457_));
  NA3        o429(.A(ori_ori_n457_), .B(ori_ori_n456_), .C(ori_ori_n183_), .Y(ori_ori_n458_));
  NO2        o430(.A(ori_ori_n821_), .B(m), .Y(ori_ori_n459_));
  NO2        o431(.A(ori_ori_n458_), .B(ori_ori_n459_), .Y(ori_ori_n460_));
  NO3        o432(.A(ori_ori_n324_), .B(ori_ori_n285_), .C(j), .Y(ori_ori_n461_));
  INV        o433(.A(j), .Y(ori_ori_n462_));
  NO3        o434(.A(ori_ori_n196_), .B(ori_ori_n462_), .C(ori_ori_n34_), .Y(ori_ori_n463_));
  AOI210     o435(.A0(ori_ori_n353_), .A1(n), .B0(ori_ori_n365_), .Y(ori_ori_n464_));
  NA2        o436(.A(ori_ori_n464_), .B(ori_ori_n368_), .Y(ori_ori_n465_));
  AN3        o437(.A(ori_ori_n465_), .B(ori_ori_n463_), .C(ori_ori_n69_), .Y(ori_ori_n466_));
  NA2        o438(.A(ori_ori_n388_), .B(ori_ori_n201_), .Y(ori_ori_n467_));
  INV        o439(.A(ori_ori_n467_), .Y(ori_ori_n468_));
  NO2        o440(.A(ori_ori_n196_), .B(ori_ori_n94_), .Y(ori_ori_n469_));
  AOI220     o441(.A0(ori_ori_n469_), .A1(ori_ori_n391_), .B0(ori_ori_n449_), .B1(ori_ori_n438_), .Y(ori_ori_n470_));
  NO2        o442(.A(ori_ori_n454_), .B(ori_ori_n66_), .Y(ori_ori_n471_));
  NA2        o443(.A(ori_ori_n471_), .B(ori_ori_n384_), .Y(ori_ori_n472_));
  NO2        o444(.A(ori_ori_n385_), .B(ori_ori_n82_), .Y(ori_ori_n473_));
  OAI210     o445(.A0(ori_ori_n473_), .A1(ori_ori_n461_), .B0(ori_ori_n414_), .Y(ori_ori_n474_));
  NA3        o446(.A(ori_ori_n474_), .B(ori_ori_n472_), .C(ori_ori_n470_), .Y(ori_ori_n475_));
  OR3        o447(.A(ori_ori_n475_), .B(ori_ori_n468_), .C(ori_ori_n466_), .Y(ori_ori_n476_));
  NA3        o448(.A(ori_ori_n464_), .B(ori_ori_n368_), .C(ori_ori_n367_), .Y(ori_ori_n477_));
  NA4        o449(.A(ori_ori_n477_), .B(ori_ori_n152_), .C(ori_ori_n293_), .D(ori_ori_n30_), .Y(ori_ori_n478_));
  NO4        o450(.A(ori_ori_n324_), .B(ori_ori_n284_), .C(j), .D(f), .Y(ori_ori_n479_));
  NO2        o451(.A(ori_ori_n67_), .B(ori_ori_n37_), .Y(ori_ori_n480_));
  NA2        o452(.A(ori_ori_n480_), .B(ori_ori_n396_), .Y(ori_ori_n481_));
  NA2        o453(.A(ori_ori_n481_), .B(ori_ori_n478_), .Y(ori_ori_n482_));
  BUFFER     o454(.A(ori_ori_n471_), .Y(ori_ori_n483_));
  NA2        o455(.A(ori_ori_n483_), .B(ori_ori_n169_), .Y(ori_ori_n484_));
  NO2        o456(.A(ori_ori_n409_), .B(ori_ori_n51_), .Y(ori_ori_n485_));
  AOI210     o457(.A0(ori_ori_n479_), .A1(ori_ori_n485_), .B0(ori_ori_n223_), .Y(ori_ori_n486_));
  OAI210     o458(.A0(ori_ori_n454_), .A1(ori_ori_n408_), .B0(ori_ori_n347_), .Y(ori_ori_n487_));
  NA3        o459(.A(ori_ori_n181_), .B(ori_ori_n47_), .C(b), .Y(ori_ori_n488_));
  AOI220     o460(.A0(ori_ori_n387_), .A1(b), .B0(ori_ori_n309_), .B1(ori_ori_n59_), .Y(ori_ori_n489_));
  NA2        o461(.A(ori_ori_n489_), .B(ori_ori_n488_), .Y(ori_ori_n490_));
  NA2        o462(.A(ori_ori_n490_), .B(ori_ori_n487_), .Y(ori_ori_n491_));
  NA3        o463(.A(ori_ori_n491_), .B(ori_ori_n486_), .C(ori_ori_n484_), .Y(ori_ori_n492_));
  NO3        o464(.A(ori_ori_n492_), .B(ori_ori_n482_), .C(ori_ori_n476_), .Y(ori_ori_n493_));
  NO3        o465(.A(ori_ori_n229_), .B(ori_ori_n197_), .C(ori_ori_n78_), .Y(ori_ori_n494_));
  NA2        o466(.A(ori_ori_n494_), .B(ori_ori_n465_), .Y(ori_ori_n495_));
  NO2        o467(.A(ori_ori_n68_), .B(h), .Y(ori_ori_n496_));
  NA2        o468(.A(ori_ori_n496_), .B(ori_ori_n435_), .Y(ori_ori_n497_));
  NA2        o469(.A(ori_ori_n497_), .B(ori_ori_n495_), .Y(ori_ori_n498_));
  NO2        o470(.A(ori_ori_n823_), .B(n), .Y(ori_ori_n499_));
  NO2        o471(.A(ori_ori_n366_), .B(ori_ori_n59_), .Y(ori_ori_n500_));
  NA2        o472(.A(ori_ori_n494_), .B(ori_ori_n500_), .Y(ori_ori_n501_));
  OAI210     o473(.A0(ori_ori_n439_), .A1(ori_ori_n263_), .B0(ori_ori_n501_), .Y(ori_ori_n502_));
  NO2        o474(.A(ori_ori_n420_), .B(n), .Y(ori_ori_n503_));
  BUFFER     o475(.A(ori_ori_n469_), .Y(ori_ori_n504_));
  AOI220     o476(.A0(ori_ori_n504_), .A1(ori_ori_n411_), .B0(ori_ori_n503_), .B1(ori_ori_n430_), .Y(ori_ori_n505_));
  INV        o477(.A(ori_ori_n505_), .Y(ori_ori_n506_));
  NO3        o478(.A(ori_ori_n506_), .B(ori_ori_n502_), .C(ori_ori_n498_), .Y(ori_ori_n507_));
  NA4        o479(.A(ori_ori_n507_), .B(ori_ori_n493_), .C(ori_ori_n460_), .D(ori_ori_n455_), .Y(ori09));
  NA2        o480(.A(ori_ori_n287_), .B(e), .Y(ori_ori_n509_));
  NO2        o481(.A(ori_ori_n509_), .B(ori_ori_n342_), .Y(ori_ori_n510_));
  INV        o482(.A(ori_ori_n510_), .Y(ori_ori_n511_));
  NA3        o483(.A(m), .B(l), .C(i), .Y(ori_ori_n512_));
  OAI220     o484(.A0(ori_ori_n385_), .A1(ori_ori_n512_), .B0(ori_ori_n238_), .B1(ori_ori_n351_), .Y(ori_ori_n513_));
  BUFFER     o485(.A(ori_ori_n513_), .Y(ori_ori_n514_));
  AN2        o486(.A(ori_ori_n514_), .B(ori_ori_n499_), .Y(ori_ori_n515_));
  INV        o487(.A(ori_ori_n226_), .Y(ori_ori_n516_));
  INV        o488(.A(ori_ori_n86_), .Y(ori_ori_n517_));
  NOi31      o489(.An(k), .B(m), .C(l), .Y(ori_ori_n518_));
  NO2        o490(.A(ori_ori_n228_), .B(ori_ori_n518_), .Y(ori_ori_n519_));
  AOI210     o491(.A0(ori_ori_n519_), .A1(ori_ori_n517_), .B0(ori_ori_n386_), .Y(ori_ori_n520_));
  NA2        o492(.A(ori_ori_n488_), .B(ori_ori_n219_), .Y(ori_ori_n521_));
  NA2        o493(.A(ori_ori_n230_), .B(m), .Y(ori_ori_n522_));
  OAI210     o494(.A0(ori_ori_n143_), .A1(ori_ori_n149_), .B0(ori_ori_n522_), .Y(ori_ori_n523_));
  AOI220     o495(.A0(ori_ori_n523_), .A1(ori_ori_n521_), .B0(ori_ori_n520_), .B1(ori_ori_n516_), .Y(ori_ori_n524_));
  NA2        o496(.A(ori_ori_n429_), .B(ori_ori_n94_), .Y(ori_ori_n525_));
  NA3        o497(.A(ori_ori_n525_), .B(ori_ori_n130_), .C(e), .Y(ori_ori_n526_));
  NA4        o498(.A(ori_ori_n526_), .B(ori_ori_n524_), .C(ori_ori_n392_), .D(ori_ori_n57_), .Y(ori_ori_n527_));
  NA2        o499(.A(f), .B(m), .Y(ori_ori_n528_));
  NO2        o500(.A(ori_ori_n528_), .B(ori_ori_n41_), .Y(ori_ori_n529_));
  NA2        o501(.A(ori_ori_n529_), .B(ori_ori_n361_), .Y(ori_ori_n530_));
  NA3        o502(.A(k), .B(i), .C(ori_ori_n83_), .Y(ori_ori_n531_));
  NA3        o503(.A(a), .B(d), .C(ori_ori_n59_), .Y(ori_ori_n532_));
  NO3        o504(.A(ori_ori_n532_), .B(ori_ori_n51_), .C(ori_ori_n150_), .Y(ori_ori_n533_));
  NA2        o505(.A(ori_ori_n531_), .B(ori_ori_n533_), .Y(ori_ori_n534_));
  NAi31      o506(.An(ori_ori_n326_), .B(ori_ori_n534_), .C(ori_ori_n530_), .Y(ori_ori_n535_));
  NO3        o507(.A(ori_ori_n91_), .B(ori_ori_n214_), .C(ori_ori_n108_), .Y(ori_ori_n536_));
  INV        o508(.A(ori_ori_n536_), .Y(ori_ori_n537_));
  NA3        o509(.A(ori_ori_n111_), .B(ori_ori_n75_), .C(o), .Y(ori_ori_n538_));
  OAI220     o510(.A0(ori_ori_n532_), .A1(ori_ori_n279_), .B0(ori_ori_n226_), .B1(ori_ori_n538_), .Y(ori_ori_n539_));
  NOi31      o511(.An(ori_ori_n156_), .B(ori_ori_n539_), .C(ori_ori_n199_), .Y(ori_ori_n540_));
  NA2        o512(.A(c), .B(ori_ori_n81_), .Y(ori_ori_n541_));
  NO2        o513(.A(ori_ori_n541_), .B(ori_ori_n272_), .Y(ori_ori_n542_));
  NA3        o514(.A(ori_ori_n542_), .B(ori_ori_n340_), .C(f), .Y(ori_ori_n543_));
  OR2        o515(.A(ori_ori_n408_), .B(ori_ori_n358_), .Y(ori_ori_n544_));
  INV        o516(.A(ori_ori_n544_), .Y(ori_ori_n545_));
  NA2        o517(.A(b), .B(ori_ori_n545_), .Y(ori_ori_n546_));
  NA4        o518(.A(ori_ori_n546_), .B(ori_ori_n543_), .C(ori_ori_n540_), .D(ori_ori_n537_), .Y(ori_ori_n547_));
  NO4        o519(.A(ori_ori_n547_), .B(ori_ori_n535_), .C(ori_ori_n527_), .D(ori_ori_n515_), .Y(ori_ori_n548_));
  NO2        o520(.A(ori_ori_n94_), .B(ori_ori_n91_), .Y(ori_ori_n549_));
  NO2        o521(.A(ori_ori_n163_), .B(ori_ori_n157_), .Y(ori_ori_n550_));
  AOI220     o522(.A0(ori_ori_n550_), .A1(ori_ori_n160_), .B0(ori_ori_n198_), .B1(ori_ori_n549_), .Y(ori_ori_n551_));
  INV        o523(.A(ori_ori_n279_), .Y(ori_ori_n552_));
  INV        o524(.A(ori_ori_n551_), .Y(ori_ori_n553_));
  NA2        o525(.A(e), .B(d), .Y(ori_ori_n554_));
  OAI220     o526(.A0(ori_ori_n554_), .A1(c), .B0(ori_ori_n209_), .B1(d), .Y(ori_ori_n555_));
  AOI210     o527(.A0(ori_ori_n344_), .A1(ori_ori_n121_), .B0(ori_ori_n163_), .Y(ori_ori_n556_));
  INV        o528(.A(ori_ori_n556_), .Y(ori_ori_n557_));
  NA3        o529(.A(k), .B(ori_ori_n60_), .C(ori_ori_n30_), .Y(ori_ori_n558_));
  NA2        o530(.A(ori_ori_n558_), .B(ori_ori_n557_), .Y(ori_ori_n559_));
  NO2        o531(.A(ori_ori_n559_), .B(ori_ori_n553_), .Y(ori_ori_n560_));
  OR2        o532(.A(ori_ori_n431_), .B(ori_ori_n153_), .Y(ori_ori_n561_));
  NO2        o533(.A(ori_ori_n509_), .B(ori_ori_n112_), .Y(ori_ori_n562_));
  AN2        o534(.A(ori_ori_n521_), .B(ori_ori_n513_), .Y(ori_ori_n563_));
  NO2        o535(.A(ori_ori_n563_), .B(ori_ori_n562_), .Y(ori_ori_n564_));
  OAI210     o536(.A0(ori_ori_n117_), .A1(ori_ori_n301_), .B0(ori_ori_n555_), .Y(ori_ori_n565_));
  NO2        o537(.A(ori_ori_n285_), .B(ori_ori_n49_), .Y(ori_ori_n566_));
  AN3        o538(.A(ori_ori_n565_), .B(ori_ori_n564_), .C(ori_ori_n561_), .Y(ori_ori_n567_));
  NA4        o539(.A(ori_ori_n567_), .B(ori_ori_n560_), .C(ori_ori_n548_), .D(ori_ori_n511_), .Y(ori12));
  NO2        o540(.A(ori_ori_n296_), .B(c), .Y(ori_ori_n569_));
  NO3        o541(.A(ori_ori_n286_), .B(ori_ori_n184_), .C(ori_ori_n150_), .Y(ori_ori_n570_));
  NA2        o542(.A(ori_ori_n570_), .B(ori_ori_n569_), .Y(ori_ori_n571_));
  NA2        o543(.A(ori_ori_n361_), .B(ori_ori_n566_), .Y(ori_ori_n572_));
  NO2        o544(.A(ori_ori_n296_), .B(ori_ori_n81_), .Y(ori_ori_n573_));
  NO2        o545(.A(ori_ori_n408_), .B(ori_ori_n252_), .Y(ori_ori_n574_));
  NA2        o546(.A(ori_ori_n574_), .B(ori_ori_n359_), .Y(ori_ori_n575_));
  NA3        o547(.A(ori_ori_n575_), .B(ori_ori_n572_), .C(ori_ori_n571_), .Y(ori_ori_n576_));
  AOI210     o548(.A0(ori_ori_n166_), .A1(ori_ori_n225_), .B0(ori_ori_n141_), .Y(ori_ori_n577_));
  BUFFER     o549(.A(ori_ori_n577_), .Y(ori_ori_n578_));
  AOI210     o550(.A0(ori_ori_n222_), .A1(ori_ori_n259_), .B0(ori_ori_n150_), .Y(ori_ori_n579_));
  OAI210     o551(.A0(ori_ori_n579_), .A1(ori_ori_n578_), .B0(ori_ori_n269_), .Y(ori_ori_n580_));
  NO2        o552(.A(ori_ori_n394_), .B(f), .Y(ori_ori_n581_));
  NO2        o553(.A(ori_ori_n385_), .B(ori_ori_n512_), .Y(ori_ori_n582_));
  NO2        o554(.A(ori_ori_n107_), .B(ori_ori_n168_), .Y(ori_ori_n583_));
  NA3        o555(.A(ori_ori_n583_), .B(ori_ori_n171_), .C(i), .Y(ori_ori_n584_));
  NA2        o556(.A(ori_ori_n584_), .B(ori_ori_n580_), .Y(ori_ori_n585_));
  OR2        o557(.A(ori_ori_n210_), .B(ori_ori_n573_), .Y(ori_ori_n586_));
  NA2        o558(.A(ori_ori_n586_), .B(ori_ori_n239_), .Y(ori_ori_n587_));
  NO3        o559(.A(ori_ori_n91_), .B(ori_ori_n108_), .C(ori_ori_n150_), .Y(ori_ori_n588_));
  NA2        o560(.A(ori_ori_n588_), .B(ori_ori_n353_), .Y(ori_ori_n589_));
  NA4        o561(.A(ori_ori_n287_), .B(d), .C(ori_ori_n122_), .D(o), .Y(ori_ori_n590_));
  NA3        o562(.A(ori_ori_n590_), .B(ori_ori_n589_), .C(ori_ori_n587_), .Y(ori_ori_n591_));
  NO3        o563(.A(ori_ori_n591_), .B(ori_ori_n585_), .C(ori_ori_n576_), .Y(ori_ori_n592_));
  NA2        o564(.A(ori_ori_n366_), .B(ori_ori_n101_), .Y(ori_ori_n593_));
  NOi21      o565(.An(ori_ori_n30_), .B(ori_ori_n404_), .Y(ori_ori_n594_));
  NA2        o566(.A(ori_ori_n594_), .B(ori_ori_n593_), .Y(ori_ori_n595_));
  NA2        o567(.A(ori_ori_n182_), .B(ori_ori_n595_), .Y(ori_ori_n596_));
  INV        o568(.A(ori_ori_n208_), .Y(ori_ori_n597_));
  NO2        o569(.A(ori_ori_n337_), .B(ori_ori_n197_), .Y(ori_ori_n598_));
  INV        o570(.A(ori_ori_n246_), .Y(ori_ori_n599_));
  NO3        o571(.A(ori_ori_n599_), .B(ori_ori_n597_), .C(ori_ori_n596_), .Y(ori_ori_n600_));
  NA2        o572(.A(ori_ori_n234_), .B(o), .Y(ori_ori_n601_));
  NA2        o573(.A(h), .B(i), .Y(ori_ori_n602_));
  NO2        o574(.A(ori_ori_n101_), .B(ori_ori_n59_), .Y(ori_ori_n603_));
  OR2        o575(.A(ori_ori_n603_), .B(ori_ori_n365_), .Y(ori_ori_n604_));
  INV        o576(.A(ori_ori_n604_), .Y(ori_ori_n605_));
  OAI220     o577(.A0(ori_ori_n605_), .A1(ori_ori_n601_), .B0(ori_ori_n826_), .B1(ori_ori_n219_), .Y(ori_ori_n606_));
  NO2        o578(.A(ori_ori_n252_), .B(ori_ori_n66_), .Y(ori_ori_n607_));
  OAI210     o579(.A0(ori_ori_n607_), .A1(ori_ori_n581_), .B0(ori_ori_n169_), .Y(ori_ori_n608_));
  NO2        o580(.A(ori_ori_n304_), .B(ori_ori_n150_), .Y(ori_ori_n609_));
  AOI220     o581(.A0(ori_ori_n609_), .A1(f), .B0(ori_ori_n586_), .B1(ori_ori_n154_), .Y(ori_ori_n610_));
  AOI220     o582(.A0(ori_ori_n574_), .A1(ori_ori_n583_), .B0(ori_ori_n384_), .B1(ori_ori_n65_), .Y(ori_ori_n611_));
  NA3        o583(.A(ori_ori_n611_), .B(ori_ori_n610_), .C(ori_ori_n608_), .Y(ori_ori_n612_));
  NA2        o584(.A(ori_ori_n398_), .B(ori_ori_n353_), .Y(ori_ori_n613_));
  INV        o585(.A(ori_ori_n613_), .Y(ori_ori_n614_));
  NO3        o586(.A(ori_ori_n614_), .B(ori_ori_n612_), .C(ori_ori_n606_), .Y(ori_ori_n615_));
  NAi31      o587(.An(ori_ori_n98_), .B(ori_ori_n274_), .C(n), .Y(ori_ori_n616_));
  NO3        o588(.A(ori_ori_n86_), .B(ori_ori_n228_), .C(ori_ori_n518_), .Y(ori_ori_n617_));
  NO2        o589(.A(ori_ori_n617_), .B(ori_ori_n616_), .Y(ori_ori_n618_));
  NO3        o590(.A(h), .B(ori_ori_n98_), .C(ori_ori_n272_), .Y(ori_ori_n619_));
  AOI210     o591(.A0(ori_ori_n619_), .A1(ori_ori_n332_), .B0(ori_ori_n618_), .Y(ori_ori_n620_));
  INV        o592(.A(ori_ori_n620_), .Y(ori_ori_n621_));
  NA2        o593(.A(ori_ori_n163_), .B(ori_ori_n113_), .Y(ori_ori_n622_));
  NO3        o594(.A(ori_ori_n201_), .B(ori_ori_n287_), .C(ori_ori_n117_), .Y(ori_ori_n623_));
  NOi31      o595(.An(ori_ori_n622_), .B(ori_ori_n623_), .C(ori_ori_n150_), .Y(ori_ori_n624_));
  NAi21      o596(.An(ori_ori_n366_), .B(ori_ori_n609_), .Y(ori_ori_n625_));
  NA2        o597(.A(ori_ori_n323_), .B(o), .Y(ori_ori_n626_));
  NA2        o598(.A(ori_ori_n626_), .B(ori_ori_n625_), .Y(ori_ori_n627_));
  NA2        o599(.A(ori_ori_n577_), .B(ori_ori_n569_), .Y(ori_ori_n628_));
  OAI220     o600(.A0(ori_ori_n574_), .A1(ori_ori_n582_), .B0(ori_ori_n361_), .B1(ori_ori_n278_), .Y(ori_ori_n629_));
  NA3        o601(.A(ori_ori_n629_), .B(ori_ori_n628_), .C(ori_ori_n389_), .Y(ori_ori_n630_));
  NA3        o602(.A(c), .B(ori_ori_n325_), .C(ori_ori_n36_), .Y(ori_ori_n631_));
  INV        o603(.A(ori_ori_n218_), .Y(ori_ori_n632_));
  NA2        o604(.A(ori_ori_n632_), .B(ori_ori_n631_), .Y(ori_ori_n633_));
  OR2        o605(.A(ori_ori_n633_), .B(ori_ori_n630_), .Y(ori_ori_n634_));
  NO4        o606(.A(ori_ori_n634_), .B(ori_ori_n627_), .C(ori_ori_n624_), .D(ori_ori_n621_), .Y(ori_ori_n635_));
  NA4        o607(.A(ori_ori_n635_), .B(ori_ori_n615_), .C(ori_ori_n600_), .D(ori_ori_n592_), .Y(ori13));
  AN2        o608(.A(d), .B(c), .Y(ori_ori_n637_));
  NA2        o609(.A(ori_ori_n637_), .B(ori_ori_n81_), .Y(ori_ori_n638_));
  NAi32      o610(.An(f), .Bn(e), .C(c), .Y(ori_ori_n639_));
  NA3        o611(.A(k), .B(j), .C(i), .Y(ori_ori_n640_));
  NO2        o612(.A(f), .B(c), .Y(ori_ori_n641_));
  NOi21      o613(.An(ori_ori_n641_), .B(ori_ori_n286_), .Y(ori_ori_n642_));
  OR2        o614(.A(m), .B(i), .Y(ori_ori_n643_));
  AN3        o615(.A(o), .B(f), .C(c), .Y(ori_ori_n644_));
  NA3        o616(.A(l), .B(k), .C(j), .Y(ori_ori_n645_));
  NA2        o617(.A(i), .B(h), .Y(ori_ori_n646_));
  NO3        o618(.A(ori_ori_n646_), .B(ori_ori_n645_), .C(ori_ori_n91_), .Y(ori_ori_n647_));
  NO2        o619(.A(ori_ori_n99_), .B(ori_ori_n194_), .Y(ori_ori_n648_));
  NO2        o620(.A(ori_ori_n351_), .B(ori_ori_n386_), .Y(ori_ori_n649_));
  NA4        o621(.A(ori_ori_n63_), .B(ori_ori_n62_), .C(o), .D(ori_ori_n149_), .Y(ori_ori_n650_));
  NA4        o622(.A(ori_ori_n376_), .B(m), .C(ori_ori_n78_), .D(ori_ori_n149_), .Y(ori_ori_n651_));
  NA3        o623(.A(ori_ori_n651_), .B(ori_ori_n247_), .C(ori_ori_n650_), .Y(ori_ori_n652_));
  NO2        o624(.A(ori_ori_n652_), .B(ori_ori_n649_), .Y(ori_ori_n653_));
  NO3        o625(.A(ori_ori_n523_), .B(ori_ori_n514_), .C(ori_ori_n446_), .Y(ori_ori_n654_));
  OAI220     o626(.A0(ori_ori_n654_), .A1(ori_ori_n422_), .B0(ori_ori_n653_), .B1(ori_ori_n383_), .Y(ori_ori_n655_));
  NOi31      o627(.An(m), .B(n), .C(f), .Y(ori_ori_n656_));
  NA2        o628(.A(ori_ori_n656_), .B(ori_ori_n40_), .Y(ori_ori_n657_));
  NA2        o629(.A(e), .B(a), .Y(ori_ori_n658_));
  OAI220     o630(.A0(ori_ori_n658_), .A1(ori_ori_n657_), .B0(ori_ori_n544_), .B1(ori_ori_n277_), .Y(ori_ori_n659_));
  NO2        o631(.A(ori_ori_n194_), .B(a), .Y(ori_ori_n660_));
  NO2        o632(.A(ori_ori_n659_), .B(ori_ori_n655_), .Y(ori_ori_n661_));
  NA2        o633(.A(c), .B(b), .Y(ori_ori_n662_));
  NO2        o634(.A(ori_ori_n434_), .B(ori_ori_n662_), .Y(ori_ori_n663_));
  NA2        o635(.A(ori_ori_n529_), .B(ori_ori_n663_), .Y(ori_ori_n664_));
  NAi21      o636(.An(ori_ori_n273_), .B(ori_ori_n663_), .Y(ori_ori_n665_));
  OAI210     o637(.A0(ori_ori_n362_), .A1(ori_ori_n33_), .B0(ori_ori_n660_), .Y(ori_ori_n666_));
  NA2        o638(.A(ori_ori_n666_), .B(ori_ori_n665_), .Y(ori_ori_n667_));
  INV        o639(.A(ori_ori_n667_), .Y(ori_ori_n668_));
  NA3        o640(.A(ori_ori_n668_), .B(ori_ori_n664_), .C(ori_ori_n661_), .Y(ori00));
  NA2        o641(.A(ori_ori_n552_), .B(ori_ori_n583_), .Y(ori_ori_n670_));
  INV        o642(.A(ori_ori_n670_), .Y(ori_ori_n671_));
  NA2        o643(.A(ori_ori_n340_), .B(f), .Y(ori_ori_n672_));
  OAI210     o644(.A0(ori_ori_n617_), .A1(ori_ori_n34_), .B0(ori_ori_n400_), .Y(ori_ori_n673_));
  NA3        o645(.A(ori_ori_n673_), .B(ori_ori_n188_), .C(n), .Y(ori_ori_n674_));
  AOI210     o646(.A0(ori_ori_n674_), .A1(ori_ori_n672_), .B0(ori_ori_n638_), .Y(ori_ori_n675_));
  NO2        o647(.A(ori_ori_n675_), .B(ori_ori_n671_), .Y(ori_ori_n676_));
  NA2        o648(.A(d), .B(b), .Y(ori_ori_n677_));
  NA3        o649(.A(ori_ori_n255_), .B(ori_ori_n155_), .C(o), .Y(ori_ori_n678_));
  OR2        o650(.A(ori_ori_n678_), .B(ori_ori_n677_), .Y(ori_ori_n679_));
  NO2        o651(.A(h), .B(o), .Y(ori_ori_n680_));
  NA4        o652(.A(ori_ori_n332_), .B(ori_ori_n312_), .C(ori_ori_n680_), .D(b), .Y(ori_ori_n681_));
  NO2        o653(.A(ori_ori_n351_), .B(ori_ori_n386_), .Y(ori_ori_n682_));
  AOI220     o654(.A0(ori_ori_n682_), .A1(ori_ori_n356_), .B0(ori_ori_n588_), .B1(ori_ori_n377_), .Y(ori_ori_n683_));
  NA2        o655(.A(ori_ori_n205_), .B(ori_ori_n178_), .Y(ori_ori_n684_));
  NA4        o656(.A(ori_ori_n684_), .B(ori_ori_n683_), .C(ori_ori_n681_), .D(ori_ori_n679_), .Y(ori_ori_n685_));
  INV        o657(.A(ori_ori_n685_), .Y(ori_ori_n686_));
  AOI210     o658(.A0(ori_ori_n178_), .A1(ori_ori_n234_), .B0(ori_ori_n380_), .Y(ori_ori_n687_));
  INV        o659(.A(ori_ori_n687_), .Y(ori_ori_n688_));
  NO2        o660(.A(ori_ori_n170_), .B(ori_ori_n122_), .Y(ori_ori_n689_));
  NA2        o661(.A(ori_ori_n689_), .B(ori_ori_n278_), .Y(ori_ori_n690_));
  INV        o662(.A(ori_ori_n690_), .Y(ori_ori_n691_));
  NO2        o663(.A(ori_ori_n691_), .B(ori_ori_n688_), .Y(ori_ori_n692_));
  AN3        o664(.A(ori_ori_n692_), .B(ori_ori_n686_), .C(ori_ori_n378_), .Y(ori_ori_n693_));
  NA3        o665(.A(ori_ori_n656_), .B(a), .C(ori_ori_n311_), .Y(ori_ori_n694_));
  NA2        o666(.A(ori_ori_n694_), .B(ori_ori_n172_), .Y(ori_ori_n695_));
  NA2        o667(.A(ori_ori_n652_), .B(ori_ori_n356_), .Y(ori_ori_n696_));
  NA4        o668(.A(ori_ori_n403_), .B(ori_ori_n145_), .C(ori_ori_n155_), .D(h), .Y(ori_ori_n697_));
  NA2        o669(.A(ori_ori_n697_), .B(ori_ori_n696_), .Y(ori_ori_n698_));
  NA2        o670(.A(n), .B(e), .Y(ori_ori_n699_));
  NO2        o671(.A(ori_ori_n699_), .B(ori_ori_n103_), .Y(ori_ori_n700_));
  NA2        o672(.A(ori_ori_n700_), .B(ori_ori_n191_), .Y(ori_ori_n701_));
  NA2        o673(.A(o), .B(ori_ori_n292_), .Y(ori_ori_n702_));
  NA2        o674(.A(ori_ori_n702_), .B(ori_ori_n701_), .Y(ori_ori_n703_));
  NA2        o675(.A(ori_ori_n700_), .B(ori_ori_n520_), .Y(ori_ori_n704_));
  AOI220     o676(.A0(ori_ori_n594_), .A1(ori_ori_n377_), .B0(ori_ori_n403_), .B1(ori_ori_n175_), .Y(ori_ori_n705_));
  NA3        o677(.A(ori_ori_n705_), .B(ori_ori_n704_), .C(ori_ori_n530_), .Y(ori_ori_n706_));
  NO4        o678(.A(ori_ori_n706_), .B(ori_ori_n703_), .C(ori_ori_n698_), .D(ori_ori_n695_), .Y(ori_ori_n707_));
  NA3        o679(.A(ori_ori_n707_), .B(ori_ori_n693_), .C(ori_ori_n676_), .Y(ori01));
  INV        o680(.A(ori_ori_n320_), .Y(ori_ori_n709_));
  NA2        o681(.A(ori_ori_n264_), .B(i), .Y(ori_ori_n710_));
  NA3        o682(.A(ori_ori_n710_), .B(ori_ori_n709_), .C(ori_ori_n628_), .Y(ori_ori_n711_));
  NA2        o683(.A(ori_ori_n384_), .B(ori_ori_n65_), .Y(ori_ori_n712_));
  NA2        o684(.A(ori_ori_n366_), .B(ori_ori_n190_), .Y(ori_ori_n713_));
  NA2        o685(.A(ori_ori_n598_), .B(ori_ori_n713_), .Y(ori_ori_n714_));
  NA3        o686(.A(ori_ori_n714_), .B(ori_ori_n712_), .C(ori_ori_n220_), .Y(ori_ori_n715_));
  NA2        o687(.A(ori_ori_n35_), .B(f), .Y(ori_ori_n716_));
  NA2        o688(.A(k), .B(o), .Y(ori_ori_n717_));
  NO2        o689(.A(ori_ori_n717_), .B(ori_ori_n716_), .Y(ori_ori_n718_));
  OR2        o690(.A(ori_ori_n409_), .B(ori_ori_n247_), .Y(ori_ori_n719_));
  NA3        o691(.A(ori_ori_n719_), .B(ori_ori_n697_), .C(ori_ori_n551_), .Y(ori_ori_n720_));
  OR2        o692(.A(ori_ori_n136_), .B(ori_ori_n134_), .Y(ori_ori_n721_));
  NA2        o693(.A(ori_ori_n721_), .B(ori_ori_n95_), .Y(ori_ori_n722_));
  NO4        o694(.A(ori_ori_n722_), .B(ori_ori_n720_), .C(ori_ori_n715_), .D(ori_ori_n711_), .Y(ori_ori_n723_));
  OAI210     o695(.A0(ori_ori_n241_), .A1(ori_ori_n30_), .B0(m), .Y(ori_ori_n724_));
  OR2        o696(.A(ori_ori_n724_), .B(ori_ori_n219_), .Y(ori_ori_n725_));
  INV        o697(.A(ori_ori_n725_), .Y(ori_ori_n726_));
  NA2        o698(.A(ori_ori_n193_), .B(ori_ori_n136_), .Y(ori_ori_n727_));
  NA2        o699(.A(ori_ori_n727_), .B(ori_ori_n411_), .Y(ori_ori_n728_));
  OAI210     o700(.A0(ori_ori_n718_), .A1(ori_ori_n213_), .B0(ori_ori_n414_), .Y(ori_ori_n729_));
  NA3        o701(.A(ori_ori_n729_), .B(ori_ori_n728_), .C(ori_ori_n481_), .Y(ori_ori_n730_));
  NO2        o702(.A(ori_ori_n730_), .B(ori_ori_n726_), .Y(ori_ori_n731_));
  NO2        o703(.A(ori_ori_n146_), .B(ori_ori_n77_), .Y(ori_ori_n732_));
  NO2        o704(.A(ori_ori_n602_), .B(ori_ori_n165_), .Y(ori_ori_n733_));
  NO2        o705(.A(ori_ori_n831_), .B(ori_ori_n368_), .Y(ori_ori_n734_));
  OAI210     o706(.A0(ori_ori_n734_), .A1(ori_ori_n733_), .B0(ori_ori_n228_), .Y(ori_ori_n735_));
  NA2        o707(.A(ori_ori_n830_), .B(ori_ori_n372_), .Y(ori_ori_n736_));
  NO3        o708(.A(ori_ori_n56_), .B(ori_ori_n197_), .C(ori_ori_n35_), .Y(ori_ori_n737_));
  NA2        o709(.A(ori_ori_n737_), .B(ori_ori_n365_), .Y(ori_ori_n738_));
  NA2        o710(.A(ori_ori_n738_), .B(ori_ori_n736_), .Y(ori_ori_n739_));
  OR2        o711(.A(ori_ori_n678_), .B(ori_ori_n677_), .Y(ori_ori_n740_));
  NA2        o712(.A(ori_ori_n737_), .B(ori_ori_n500_), .Y(ori_ori_n741_));
  NA2        o713(.A(ori_ori_n741_), .B(ori_ori_n740_), .Y(ori_ori_n742_));
  NOi41      o714(.An(ori_ori_n735_), .B(ori_ori_n742_), .C(ori_ori_n739_), .D(ori_ori_n732_), .Y(ori_ori_n743_));
  NO2        o715(.A(ori_ori_n90_), .B(ori_ori_n35_), .Y(ori_ori_n744_));
  AO220      o716(.A0(i), .A1(ori_ori_n391_), .B0(ori_ori_n744_), .B1(ori_ori_n438_), .Y(ori_ori_n745_));
  NA2        o717(.A(ori_ori_n745_), .B(ori_ori_n228_), .Y(ori_ori_n746_));
  NO3        o718(.A(ori_ori_n646_), .B(ori_ori_n118_), .C(ori_ori_n62_), .Y(ori_ori_n747_));
  NA4        o719(.A(ori_ori_n746_), .B(ori_ori_n743_), .C(ori_ori_n731_), .D(ori_ori_n723_), .Y(ori06));
  NO2        o720(.A(ori_ori_n157_), .B(ori_ori_n70_), .Y(ori_ori_n749_));
  OAI210     o721(.A0(ori_ori_n749_), .A1(ori_ori_n747_), .B0(f), .Y(ori_ori_n750_));
  NA2        o722(.A(ori_ori_n750_), .B(ori_ori_n735_), .Y(ori_ori_n751_));
  NO3        o723(.A(ori_ori_n751_), .B(ori_ori_n739_), .C(ori_ori_n187_), .Y(ori_ori_n752_));
  NO2        o724(.A(ori_ori_n197_), .B(ori_ori_n35_), .Y(ori_ori_n753_));
  NA2        o725(.A(ori_ori_n753_), .B(ori_ori_n604_), .Y(ori_ori_n754_));
  AOI210     o726(.A0(ori_ori_n753_), .A1(ori_ori_n369_), .B0(ori_ori_n745_), .Y(ori_ori_n755_));
  AOI210     o727(.A0(ori_ori_n755_), .A1(ori_ori_n754_), .B0(ori_ori_n225_), .Y(ori_ori_n756_));
  NA2        o728(.A(ori_ori_n63_), .B(ori_ori_n396_), .Y(ori_ori_n757_));
  NO2        o729(.A(ori_ori_n824_), .B(ori_ori_n657_), .Y(ori_ori_n758_));
  OAI210     o730(.A0(ori_ori_n305_), .A1(ori_ori_n179_), .B0(ori_ori_n558_), .Y(ori_ori_n759_));
  NO2        o731(.A(ori_ori_n759_), .B(ori_ori_n758_), .Y(ori_ori_n760_));
  NA2        o732(.A(ori_ori_n760_), .B(ori_ori_n757_), .Y(ori_ori_n761_));
  AN2        o733(.A(ori_ori_n594_), .B(ori_ori_n399_), .Y(ori_ori_n762_));
  NO3        o734(.A(ori_ori_n762_), .B(ori_ori_n761_), .C(ori_ori_n756_), .Y(ori_ori_n763_));
  NA2        o735(.A(ori_ori_n242_), .B(ori_ori_n79_), .Y(ori_ori_n764_));
  NO3        o736(.A(ori_ori_n174_), .B(ori_ori_n70_), .C(ori_ori_n194_), .Y(ori_ori_n765_));
  OAI220     o737(.A0(ori_ori_n431_), .A1(ori_ori_n179_), .B0(ori_ori_n342_), .B1(ori_ori_n344_), .Y(ori_ori_n766_));
  INV        o738(.A(k), .Y(ori_ori_n767_));
  NO3        o739(.A(ori_ori_n767_), .B(ori_ori_n386_), .C(j), .Y(ori_ori_n768_));
  NO3        o740(.A(ori_ori_n766_), .B(ori_ori_n765_), .C(ori_ori_n659_), .Y(ori_ori_n769_));
  INV        o741(.A(ori_ori_n488_), .Y(ori_ori_n770_));
  NA2        o742(.A(ori_ori_n770_), .B(ori_ori_n142_), .Y(ori_ori_n771_));
  NA4        o743(.A(ori_ori_n771_), .B(ori_ori_n769_), .C(ori_ori_n764_), .D(ori_ori_n705_), .Y(ori_ori_n772_));
  NA2        o744(.A(ori_ori_n768_), .B(ori_ori_n485_), .Y(ori_ori_n773_));
  INV        o745(.A(ori_ori_n773_), .Y(ori_ori_n774_));
  AN2        o746(.A(ori_ori_n570_), .B(ori_ori_n569_), .Y(ori_ori_n775_));
  NO3        o747(.A(ori_ori_n775_), .B(ori_ori_n334_), .C(ori_ori_n323_), .Y(ori_ori_n776_));
  NA2        o748(.A(ori_ori_n776_), .B(ori_ori_n741_), .Y(ori_ori_n777_));
  NO3        o749(.A(ori_ori_n777_), .B(ori_ori_n774_), .C(ori_ori_n772_), .Y(ori_ori_n778_));
  NA4        o750(.A(ori_ori_n778_), .B(ori_ori_n763_), .C(ori_ori_n752_), .D(ori_ori_n746_), .Y(ori07));
  NAi32      o751(.An(m), .Bn(b), .C(n), .Y(ori_ori_n780_));
  NO3        o752(.A(ori_ori_n780_), .B(o), .C(f), .Y(ori_ori_n781_));
  NOi31      o753(.An(n), .B(m), .C(b), .Y(ori_ori_n782_));
  NO3        o754(.A(ori_ori_n91_), .B(ori_ori_n293_), .C(h), .Y(ori_ori_n783_));
  NO2        o755(.A(m), .B(h), .Y(ori_ori_n784_));
  NO2        o756(.A(ori_ori_n639_), .B(ori_ori_n286_), .Y(ori_ori_n785_));
  NO2        o757(.A(ori_ori_n640_), .B(ori_ori_n200_), .Y(ori_ori_n786_));
  NO2        o758(.A(ori_ori_n785_), .B(ori_ori_n781_), .Y(ori_ori_n787_));
  NO2        o759(.A(l), .B(k), .Y(ori_ori_n788_));
  NO3        o760(.A(ori_ori_n286_), .B(d), .C(c), .Y(ori_ori_n789_));
  NA2        o761(.A(ori_ori_n644_), .B(ori_ori_n312_), .Y(ori_ori_n790_));
  NO2        o762(.A(ori_ori_n790_), .B(ori_ori_n286_), .Y(ori_ori_n791_));
  NA2        o763(.A(ori_ori_n782_), .B(ori_ori_n253_), .Y(ori_ori_n792_));
  INV        o764(.A(ori_ori_n792_), .Y(ori_ori_n793_));
  INV        o765(.A(ori_ori_n647_), .Y(ori_ori_n794_));
  NAi21      o766(.An(ori_ori_n793_), .B(ori_ori_n794_), .Y(ori_ori_n795_));
  NA2        o767(.A(ori_ori_n784_), .B(ori_ori_n788_), .Y(ori_ori_n796_));
  NO2        o768(.A(ori_ori_n825_), .B(ori_ori_n795_), .Y(ori_ori_n797_));
  NA3        o769(.A(ori_ori_n797_), .B(ori_ori_n828_), .C(ori_ori_n787_), .Y(ori_ori_n798_));
  NA2        o770(.A(ori_ori_n642_), .B(ori_ori_n106_), .Y(ori_ori_n799_));
  NO2        o771(.A(ori_ori_n157_), .B(ori_ori_n118_), .Y(ori_ori_n800_));
  NO2        o772(.A(ori_ori_n643_), .B(h), .Y(ori_ori_n801_));
  NO2        o773(.A(j), .B(ori_ori_n116_), .Y(ori_ori_n802_));
  NA2        o774(.A(h), .B(ori_ori_n802_), .Y(ori_ori_n803_));
  INV        o775(.A(ori_ori_n803_), .Y(ori_ori_n804_));
  NO3        o776(.A(ori_ori_n804_), .B(ori_ori_n79_), .C(ori_ori_n801_), .Y(ori_ori_n805_));
  NA3        o777(.A(ori_ori_n805_), .B(ori_ori_n827_), .C(ori_ori_n799_), .Y(ori_ori_n806_));
  NA2        o778(.A(h), .B(ori_ori_n786_), .Y(ori_ori_n807_));
  NA2        o779(.A(ori_ori_n782_), .B(ori_ori_n541_), .Y(ori_ori_n808_));
  NA2        o780(.A(ori_ori_n808_), .B(ori_ori_n807_), .Y(ori_ori_n809_));
  INV        o781(.A(ori_ori_n809_), .Y(ori_ori_n810_));
  OR2        o782(.A(h), .B(ori_ori_n357_), .Y(ori_ori_n811_));
  NO2        o783(.A(ori_ori_n811_), .B(ori_ori_n116_), .Y(ori_ori_n812_));
  NA2        o784(.A(ori_ori_n648_), .B(ori_ori_n155_), .Y(ori_ori_n813_));
  INV        o785(.A(ori_ori_n813_), .Y(ori_ori_n814_));
  NO3        o786(.A(ori_ori_n814_), .B(ori_ori_n812_), .C(ori_ori_n789_), .Y(ori_ori_n815_));
  NA2        o787(.A(ori_ori_n815_), .B(ori_ori_n810_), .Y(ori_ori_n816_));
  OR4        o788(.A(ori_ori_n783_), .B(ori_ori_n816_), .C(ori_ori_n806_), .D(ori_ori_n798_), .Y(ori04));
  INV        o789(.A(ori_ori_n30_), .Y(ori_ori_n820_));
  INV        o790(.A(ori_ori_n421_), .Y(ori_ori_n821_));
  INV        o791(.A(ori_ori_n385_), .Y(ori_ori_n822_));
  INV        o792(.A(a), .Y(ori_ori_n823_));
  INV        o793(.A(a), .Y(ori_ori_n824_));
  INV        o794(.A(ori_ori_n796_), .Y(ori_ori_n825_));
  INV        o795(.A(ori_ori_n31_), .Y(ori_ori_n826_));
  INV        o796(.A(ori_ori_n800_), .Y(ori_ori_n827_));
  INV        o797(.A(ori_ori_n791_), .Y(ori_ori_n828_));
  INV        o798(.A(ori_ori_n353_), .Y(ori_ori_n829_));
  INV        o799(.A(k), .Y(ori_ori_n830_));
  INV        o800(.A(h), .Y(ori_ori_n831_));
  ZERO       o801(.Y(ori02));
  ZERO       o802(.Y(ori03));
  ZERO       o803(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(m), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(m), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(m), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(m), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(m), .Y(mai_mai_n50_));
  INV        m0022(.A(c), .Y(mai_mai_n51_));
  NA2        m0023(.A(e), .B(b), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  INV        m0025(.A(d), .Y(mai_mai_n54_));
  NAi21      m0026(.An(i), .B(h), .Y(mai_mai_n55_));
  NAi31      m0027(.An(i), .B(l), .C(j), .Y(mai_mai_n56_));
  OAI220     m0028(.A0(mai_mai_n56_), .A1(mai_mai_n49_), .B0(mai_mai_n55_), .B1(mai_mai_n44_), .Y(mai_mai_n57_));
  NAi31      m0029(.An(mai_mai_n1279_), .B(mai_mai_n57_), .C(mai_mai_n53_), .Y(mai_mai_n58_));
  NA2        m0030(.A(m), .B(f), .Y(mai_mai_n59_));
  NAi32      m0031(.An(n), .Bn(k), .C(m), .Y(mai_mai_n60_));
  NAi31      m0032(.An(l), .B(m), .C(k), .Y(mai_mai_n61_));
  NAi41      m0033(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n62_));
  INV        m0034(.A(m), .Y(mai_mai_n63_));
  NOi21      m0035(.An(k), .B(l), .Y(mai_mai_n64_));
  NOi32      m0036(.An(h), .Bn(m), .C(f), .Y(mai_mai_n65_));
  INV        m0037(.A(mai_mai_n58_), .Y(mai_mai_n66_));
  INV        m0038(.A(n), .Y(mai_mai_n67_));
  NOi32      m0039(.An(e), .Bn(b), .C(d), .Y(mai_mai_n68_));
  NA2        m0040(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  INV        m0041(.A(j), .Y(mai_mai_n70_));
  AN3        m0042(.A(m), .B(k), .C(i), .Y(mai_mai_n71_));
  NA3        m0043(.A(mai_mai_n71_), .B(mai_mai_n70_), .C(m), .Y(mai_mai_n72_));
  NAi32      m0044(.An(m), .Bn(f), .C(h), .Y(mai_mai_n73_));
  NAi31      m0045(.An(j), .B(m), .C(l), .Y(mai_mai_n74_));
  NO2        m0046(.A(mai_mai_n74_), .B(mai_mai_n73_), .Y(mai_mai_n75_));
  NA2        m0047(.A(m), .B(l), .Y(mai_mai_n76_));
  NAi31      m0048(.An(k), .B(j), .C(m), .Y(mai_mai_n77_));
  NO3        m0049(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(f), .Y(mai_mai_n78_));
  AN2        m0050(.A(j), .B(m), .Y(mai_mai_n79_));
  NOi32      m0051(.An(m), .Bn(l), .C(i), .Y(mai_mai_n80_));
  NOi21      m0052(.An(m), .B(i), .Y(mai_mai_n81_));
  NOi32      m0053(.An(m), .Bn(j), .C(k), .Y(mai_mai_n82_));
  AOI220     m0054(.A0(mai_mai_n82_), .A1(mai_mai_n81_), .B0(mai_mai_n80_), .B1(mai_mai_n79_), .Y(mai_mai_n83_));
  NO2        m0055(.A(mai_mai_n83_), .B(f), .Y(mai_mai_n84_));
  NO3        m0056(.A(mai_mai_n84_), .B(mai_mai_n78_), .C(mai_mai_n75_), .Y(mai_mai_n85_));
  NAi41      m0057(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n86_));
  AN2        m0058(.A(e), .B(b), .Y(mai_mai_n87_));
  NOi31      m0059(.An(c), .B(h), .C(f), .Y(mai_mai_n88_));
  NA2        m0060(.A(mai_mai_n88_), .B(mai_mai_n87_), .Y(mai_mai_n89_));
  NOi21      m0061(.An(m), .B(f), .Y(mai_mai_n90_));
  NOi21      m0062(.An(i), .B(h), .Y(mai_mai_n91_));
  NA3        m0063(.A(mai_mai_n91_), .B(mai_mai_n90_), .C(mai_mai_n36_), .Y(mai_mai_n92_));
  INV        m0064(.A(a), .Y(mai_mai_n93_));
  NA2        m0065(.A(mai_mai_n87_), .B(mai_mai_n93_), .Y(mai_mai_n94_));
  INV        m0066(.A(l), .Y(mai_mai_n95_));
  NOi21      m0067(.An(m), .B(n), .Y(mai_mai_n96_));
  NO2        m0068(.A(mai_mai_n92_), .B(mai_mai_n69_), .Y(mai_mai_n97_));
  INV        m0069(.A(b), .Y(mai_mai_n98_));
  NA2        m0070(.A(l), .B(j), .Y(mai_mai_n99_));
  AN2        m0071(.A(k), .B(i), .Y(mai_mai_n100_));
  NA2        m0072(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  NA2        m0073(.A(m), .B(e), .Y(mai_mai_n102_));
  NOi32      m0074(.An(c), .Bn(a), .C(d), .Y(mai_mai_n103_));
  NA2        m0075(.A(mai_mai_n103_), .B(mai_mai_n96_), .Y(mai_mai_n104_));
  INV        m0076(.A(mai_mai_n97_), .Y(mai_mai_n105_));
  OAI210     m0077(.A0(mai_mai_n85_), .A1(mai_mai_n69_), .B0(mai_mai_n105_), .Y(mai_mai_n106_));
  NOi31      m0078(.An(k), .B(m), .C(j), .Y(mai_mai_n107_));
  NOi31      m0079(.An(k), .B(m), .C(i), .Y(mai_mai_n108_));
  NA3        m0080(.A(mai_mai_n108_), .B(mai_mai_n65_), .C(c), .Y(mai_mai_n109_));
  INV        m0081(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NOi32      m0082(.An(f), .Bn(b), .C(e), .Y(mai_mai_n111_));
  NAi21      m0083(.An(m), .B(h), .Y(mai_mai_n112_));
  NAi21      m0084(.An(m), .B(n), .Y(mai_mai_n113_));
  NAi21      m0085(.An(j), .B(k), .Y(mai_mai_n114_));
  NAi41      m0086(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n115_));
  NAi31      m0087(.An(j), .B(k), .C(h), .Y(mai_mai_n116_));
  NO3        m0088(.A(mai_mai_n116_), .B(mai_mai_n115_), .C(mai_mai_n113_), .Y(mai_mai_n117_));
  INV        m0089(.A(mai_mai_n117_), .Y(mai_mai_n118_));
  NO2        m0090(.A(k), .B(j), .Y(mai_mai_n119_));
  AN2        m0091(.A(k), .B(j), .Y(mai_mai_n120_));
  NAi21      m0092(.An(c), .B(b), .Y(mai_mai_n121_));
  NA2        m0093(.A(f), .B(d), .Y(mai_mai_n122_));
  NA2        m0094(.A(h), .B(c), .Y(mai_mai_n123_));
  NAi31      m0095(.An(f), .B(e), .C(b), .Y(mai_mai_n124_));
  NA2        m0096(.A(d), .B(b), .Y(mai_mai_n125_));
  NAi21      m0097(.An(e), .B(f), .Y(mai_mai_n126_));
  NO2        m0098(.A(mai_mai_n126_), .B(mai_mai_n125_), .Y(mai_mai_n127_));
  NA2        m0099(.A(b), .B(a), .Y(mai_mai_n128_));
  NAi21      m0100(.An(c), .B(d), .Y(mai_mai_n129_));
  NAi31      m0101(.An(l), .B(k), .C(h), .Y(mai_mai_n130_));
  NO2        m0102(.A(mai_mai_n113_), .B(mai_mai_n130_), .Y(mai_mai_n131_));
  NA2        m0103(.A(mai_mai_n131_), .B(mai_mai_n127_), .Y(mai_mai_n132_));
  NAi31      m0104(.An(mai_mai_n110_), .B(mai_mai_n132_), .C(mai_mai_n118_), .Y(mai_mai_n133_));
  NAi31      m0105(.An(e), .B(f), .C(b), .Y(mai_mai_n134_));
  INV        m0106(.A(mai_mai_n134_), .Y(mai_mai_n135_));
  NOi21      m0107(.An(h), .B(i), .Y(mai_mai_n136_));
  NOi21      m0108(.An(k), .B(m), .Y(mai_mai_n137_));
  NA3        m0109(.A(mai_mai_n137_), .B(mai_mai_n136_), .C(n), .Y(mai_mai_n138_));
  NOi21      m0110(.An(mai_mai_n135_), .B(mai_mai_n138_), .Y(mai_mai_n139_));
  NOi21      m0111(.An(h), .B(m), .Y(mai_mai_n140_));
  NO2        m0112(.A(mai_mai_n122_), .B(mai_mai_n121_), .Y(mai_mai_n141_));
  NAi31      m0113(.An(l), .B(j), .C(h), .Y(mai_mai_n142_));
  NOi32      m0114(.An(n), .Bn(k), .C(m), .Y(mai_mai_n143_));
  NA2        m0115(.A(l), .B(i), .Y(mai_mai_n144_));
  NAi31      m0116(.An(d), .B(f), .C(c), .Y(mai_mai_n145_));
  NAi31      m0117(.An(e), .B(f), .C(c), .Y(mai_mai_n146_));
  NA2        m0118(.A(mai_mai_n146_), .B(mai_mai_n145_), .Y(mai_mai_n147_));
  NA2        m0119(.A(j), .B(h), .Y(mai_mai_n148_));
  OR3        m0120(.A(n), .B(m), .C(k), .Y(mai_mai_n149_));
  NO2        m0121(.A(mai_mai_n149_), .B(mai_mai_n148_), .Y(mai_mai_n150_));
  NAi32      m0122(.An(m), .Bn(k), .C(n), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n151_), .B(mai_mai_n148_), .Y(mai_mai_n152_));
  AOI220     m0124(.A0(mai_mai_n152_), .A1(mai_mai_n135_), .B0(mai_mai_n150_), .B1(mai_mai_n147_), .Y(mai_mai_n153_));
  NO2        m0125(.A(n), .B(m), .Y(mai_mai_n154_));
  NA2        m0126(.A(mai_mai_n154_), .B(h), .Y(mai_mai_n155_));
  NAi21      m0127(.An(f), .B(e), .Y(mai_mai_n156_));
  NA2        m0128(.A(d), .B(c), .Y(mai_mai_n157_));
  NAi21      m0129(.An(d), .B(c), .Y(mai_mai_n158_));
  NAi31      m0130(.An(m), .B(n), .C(b), .Y(mai_mai_n159_));
  NA2        m0131(.A(k), .B(i), .Y(mai_mai_n160_));
  NAi21      m0132(.An(h), .B(f), .Y(mai_mai_n161_));
  NO2        m0133(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n159_), .B(mai_mai_n129_), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  NOi32      m0136(.An(f), .Bn(c), .C(d), .Y(mai_mai_n165_));
  NOi32      m0137(.An(f), .Bn(c), .C(e), .Y(mai_mai_n166_));
  NO2        m0138(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  NO3        m0139(.A(n), .B(m), .C(j), .Y(mai_mai_n168_));
  NA2        m0140(.A(mai_mai_n168_), .B(h), .Y(mai_mai_n169_));
  AO210      m0141(.A0(mai_mai_n169_), .A1(mai_mai_n155_), .B0(mai_mai_n167_), .Y(mai_mai_n170_));
  NA3        m0142(.A(mai_mai_n170_), .B(mai_mai_n164_), .C(mai_mai_n153_), .Y(mai_mai_n171_));
  OR3        m0143(.A(mai_mai_n171_), .B(mai_mai_n139_), .C(mai_mai_n133_), .Y(mai_mai_n172_));
  NO3        m0144(.A(mai_mai_n172_), .B(mai_mai_n106_), .C(mai_mai_n66_), .Y(mai_mai_n173_));
  NA3        m0145(.A(m), .B(mai_mai_n95_), .C(j), .Y(mai_mai_n174_));
  NAi31      m0146(.An(n), .B(h), .C(m), .Y(mai_mai_n175_));
  NO2        m0147(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  NOi32      m0148(.An(m), .Bn(k), .C(l), .Y(mai_mai_n177_));
  NA3        m0149(.A(mai_mai_n177_), .B(mai_mai_n70_), .C(m), .Y(mai_mai_n178_));
  AN2        m0150(.A(i), .B(m), .Y(mai_mai_n179_));
  NA3        m0151(.A(mai_mai_n64_), .B(mai_mai_n179_), .C(mai_mai_n96_), .Y(mai_mai_n180_));
  NAi41      m0152(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n181_));
  INV        m0153(.A(mai_mai_n181_), .Y(mai_mai_n182_));
  INV        m0154(.A(f), .Y(mai_mai_n183_));
  INV        m0155(.A(m), .Y(mai_mai_n184_));
  NOi31      m0156(.An(i), .B(j), .C(h), .Y(mai_mai_n185_));
  NOi21      m0157(.An(l), .B(m), .Y(mai_mai_n186_));
  NA2        m0158(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  NO2        m0159(.A(mai_mai_n187_), .B(mai_mai_n184_), .Y(mai_mai_n188_));
  NA2        m0160(.A(mai_mai_n188_), .B(mai_mai_n182_), .Y(mai_mai_n189_));
  OAI210     m0161(.A0(mai_mai_n1276_), .A1(mai_mai_n32_), .B0(mai_mai_n189_), .Y(mai_mai_n190_));
  NOi21      m0162(.An(n), .B(m), .Y(mai_mai_n191_));
  NOi32      m0163(.An(l), .Bn(i), .C(j), .Y(mai_mai_n192_));
  NA2        m0164(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  OR2        m0165(.A(mai_mai_n193_), .B(mai_mai_n89_), .Y(mai_mai_n194_));
  NAi21      m0166(.An(j), .B(h), .Y(mai_mai_n195_));
  XN2        m0167(.A(i), .B(h), .Y(mai_mai_n196_));
  NA2        m0168(.A(mai_mai_n196_), .B(mai_mai_n195_), .Y(mai_mai_n197_));
  NOi31      m0169(.An(k), .B(n), .C(m), .Y(mai_mai_n198_));
  NOi31      m0170(.An(mai_mai_n198_), .B(mai_mai_n157_), .C(mai_mai_n156_), .Y(mai_mai_n199_));
  NA2        m0171(.A(mai_mai_n199_), .B(mai_mai_n197_), .Y(mai_mai_n200_));
  NAi31      m0172(.An(f), .B(e), .C(c), .Y(mai_mai_n201_));
  NO4        m0173(.A(mai_mai_n201_), .B(mai_mai_n149_), .C(mai_mai_n148_), .D(mai_mai_n54_), .Y(mai_mai_n202_));
  NA4        m0174(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n203_));
  NAi32      m0175(.An(m), .Bn(i), .C(k), .Y(mai_mai_n204_));
  NO3        m0176(.A(mai_mai_n204_), .B(mai_mai_n73_), .C(mai_mai_n203_), .Y(mai_mai_n205_));
  INV        m0177(.A(k), .Y(mai_mai_n206_));
  NO2        m0178(.A(mai_mai_n205_), .B(mai_mai_n202_), .Y(mai_mai_n207_));
  NAi21      m0179(.An(n), .B(a), .Y(mai_mai_n208_));
  AN3        m0180(.A(mai_mai_n207_), .B(mai_mai_n200_), .C(mai_mai_n194_), .Y(mai_mai_n209_));
  NO2        m0181(.A(h), .B(mai_mai_n86_), .Y(mai_mai_n210_));
  NA2        m0182(.A(mai_mai_n210_), .B(mai_mai_n111_), .Y(mai_mai_n211_));
  NO2        m0183(.A(e), .B(mai_mai_n183_), .Y(mai_mai_n212_));
  NA2        m0184(.A(mai_mai_n137_), .B(mai_mai_n91_), .Y(mai_mai_n213_));
  NO2        m0185(.A(n), .B(a), .Y(mai_mai_n214_));
  NAi21      m0186(.An(h), .B(i), .Y(mai_mai_n215_));
  NA2        m0187(.A(mai_mai_n154_), .B(k), .Y(mai_mai_n216_));
  NO2        m0188(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n217_));
  NA2        m0189(.A(mai_mai_n217_), .B(mai_mai_n165_), .Y(mai_mai_n218_));
  NA2        m0190(.A(mai_mai_n218_), .B(mai_mai_n211_), .Y(mai_mai_n219_));
  NOi21      m0191(.An(m), .B(e), .Y(mai_mai_n220_));
  NO2        m0192(.A(mai_mai_n62_), .B(mai_mai_n63_), .Y(mai_mai_n221_));
  NOi32      m0193(.An(l), .Bn(j), .C(i), .Y(mai_mai_n222_));
  AOI210     m0194(.A0(mai_mai_n64_), .A1(mai_mai_n70_), .B0(mai_mai_n222_), .Y(mai_mai_n223_));
  NAi21      m0195(.An(f), .B(m), .Y(mai_mai_n224_));
  NO2        m0196(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n225_));
  NOi31      m0197(.An(mai_mai_n209_), .B(mai_mai_n219_), .C(mai_mai_n190_), .Y(mai_mai_n226_));
  NO4        m0198(.A(mai_mai_n176_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n227_));
  NO2        m0199(.A(mai_mai_n227_), .B(mai_mai_n94_), .Y(mai_mai_n228_));
  NAi21      m0200(.An(h), .B(m), .Y(mai_mai_n229_));
  OR3        m0201(.A(mai_mai_n229_), .B(mai_mai_n193_), .C(e), .Y(mai_mai_n230_));
  NAi31      m0202(.An(m), .B(k), .C(h), .Y(mai_mai_n231_));
  NO3        m0203(.A(mai_mai_n113_), .B(mai_mai_n231_), .C(l), .Y(mai_mai_n232_));
  NAi31      m0204(.An(e), .B(d), .C(a), .Y(mai_mai_n233_));
  NA2        m0205(.A(mai_mai_n232_), .B(mai_mai_n111_), .Y(mai_mai_n234_));
  NA2        m0206(.A(mai_mai_n234_), .B(mai_mai_n230_), .Y(mai_mai_n235_));
  NA3        m0207(.A(mai_mai_n137_), .B(mai_mai_n136_), .C(mai_mai_n67_), .Y(mai_mai_n236_));
  NO2        m0208(.A(mai_mai_n236_), .B(mai_mai_n167_), .Y(mai_mai_n237_));
  NA3        m0209(.A(e), .B(c), .C(b), .Y(mai_mai_n238_));
  NO2        m0210(.A(mai_mai_n1279_), .B(mai_mai_n238_), .Y(mai_mai_n239_));
  NAi32      m0211(.An(k), .Bn(i), .C(j), .Y(mai_mai_n240_));
  NAi31      m0212(.An(h), .B(l), .C(i), .Y(mai_mai_n241_));
  NA3        m0213(.A(mai_mai_n241_), .B(mai_mai_n240_), .C(mai_mai_n142_), .Y(mai_mai_n242_));
  NOi21      m0214(.An(mai_mai_n242_), .B(mai_mai_n49_), .Y(mai_mai_n243_));
  NA2        m0215(.A(mai_mai_n239_), .B(mai_mai_n243_), .Y(mai_mai_n244_));
  NAi21      m0216(.An(l), .B(k), .Y(mai_mai_n245_));
  NOi21      m0217(.An(l), .B(j), .Y(mai_mai_n246_));
  NA2        m0218(.A(mai_mai_n140_), .B(mai_mai_n246_), .Y(mai_mai_n247_));
  OR3        m0219(.A(mai_mai_n62_), .B(mai_mai_n63_), .C(e), .Y(mai_mai_n248_));
  AOI210     m0220(.A0(mai_mai_n1280_), .A1(mai_mai_n247_), .B0(mai_mai_n248_), .Y(mai_mai_n249_));
  INV        m0221(.A(mai_mai_n249_), .Y(mai_mai_n250_));
  NAi32      m0222(.An(j), .Bn(h), .C(i), .Y(mai_mai_n251_));
  NAi21      m0223(.An(m), .B(l), .Y(mai_mai_n252_));
  NO3        m0224(.A(mai_mai_n252_), .B(mai_mai_n251_), .C(mai_mai_n67_), .Y(mai_mai_n253_));
  NA2        m0225(.A(h), .B(m), .Y(mai_mai_n254_));
  OAI210     m0226(.A0(mai_mai_n143_), .A1(mai_mai_n253_), .B0(mai_mai_n141_), .Y(mai_mai_n255_));
  NA3        m0227(.A(mai_mai_n255_), .B(mai_mai_n250_), .C(mai_mai_n244_), .Y(mai_mai_n256_));
  NAi32      m0228(.An(n), .Bn(m), .C(l), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n257_), .B(mai_mai_n251_), .Y(mai_mai_n258_));
  INV        m0230(.A(mai_mai_n104_), .Y(mai_mai_n259_));
  NAi31      m0231(.An(k), .B(l), .C(j), .Y(mai_mai_n260_));
  NA2        m0232(.A(mai_mai_n245_), .B(mai_mai_n260_), .Y(mai_mai_n261_));
  NA2        m0233(.A(mai_mai_n1281_), .B(mai_mai_n259_), .Y(mai_mai_n262_));
  INV        m0234(.A(mai_mai_n262_), .Y(mai_mai_n263_));
  NO4        m0235(.A(mai_mai_n263_), .B(mai_mai_n256_), .C(mai_mai_n235_), .D(mai_mai_n228_), .Y(mai_mai_n264_));
  NA2        m0236(.A(mai_mai_n217_), .B(mai_mai_n166_), .Y(mai_mai_n265_));
  NAi21      m0237(.An(m), .B(k), .Y(mai_mai_n266_));
  NO2        m0238(.A(mai_mai_n196_), .B(mai_mai_n266_), .Y(mai_mai_n267_));
  NAi41      m0239(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n268_));
  NO2        m0240(.A(mai_mai_n268_), .B(e), .Y(mai_mai_n269_));
  NA2        m0241(.A(mai_mai_n269_), .B(mai_mai_n267_), .Y(mai_mai_n270_));
  NAi31      m0242(.An(i), .B(l), .C(h), .Y(mai_mai_n271_));
  NA2        m0243(.A(e), .B(c), .Y(mai_mai_n272_));
  NO3        m0244(.A(mai_mai_n272_), .B(n), .C(d), .Y(mai_mai_n273_));
  NA2        m0245(.A(f), .B(mai_mai_n100_), .Y(mai_mai_n274_));
  NO2        m0246(.A(mai_mai_n274_), .B(mai_mai_n184_), .Y(mai_mai_n275_));
  NAi31      m0247(.An(d), .B(e), .C(b), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n113_), .B(mai_mai_n276_), .Y(mai_mai_n277_));
  NA2        m0249(.A(mai_mai_n277_), .B(mai_mai_n275_), .Y(mai_mai_n278_));
  NA3        m0250(.A(mai_mai_n278_), .B(mai_mai_n270_), .C(mai_mai_n265_), .Y(mai_mai_n279_));
  NA2        m0251(.A(mai_mai_n214_), .B(mai_mai_n87_), .Y(mai_mai_n280_));
  OR2        m0252(.A(mai_mai_n280_), .B(mai_mai_n178_), .Y(mai_mai_n281_));
  NOi31      m0253(.An(l), .B(n), .C(m), .Y(mai_mai_n282_));
  NA2        m0254(.A(mai_mai_n282_), .B(mai_mai_n185_), .Y(mai_mai_n283_));
  NO2        m0255(.A(mai_mai_n283_), .B(mai_mai_n167_), .Y(mai_mai_n284_));
  NAi21      m0256(.An(mai_mai_n284_), .B(mai_mai_n281_), .Y(mai_mai_n285_));
  NAi32      m0257(.An(m), .Bn(j), .C(k), .Y(mai_mai_n286_));
  NAi41      m0258(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n287_));
  NOi21      m0259(.An(j), .B(m), .Y(mai_mai_n288_));
  AN3        m0260(.A(h), .B(m), .C(f), .Y(mai_mai_n289_));
  NO2        m0261(.A(mai_mai_n252_), .B(mai_mai_n251_), .Y(mai_mai_n290_));
  NO2        m0262(.A(mai_mai_n187_), .B(m), .Y(mai_mai_n291_));
  INV        m0263(.A(mai_mai_n204_), .Y(mai_mai_n292_));
  NA3        m0264(.A(mai_mai_n292_), .B(mai_mai_n289_), .C(mai_mai_n182_), .Y(mai_mai_n293_));
  INV        m0265(.A(mai_mai_n293_), .Y(mai_mai_n294_));
  NA3        m0266(.A(h), .B(m), .C(f), .Y(mai_mai_n295_));
  NA2        m0267(.A(mai_mai_n140_), .B(e), .Y(mai_mai_n296_));
  NO2        m0268(.A(mai_mai_n296_), .B(mai_mai_n41_), .Y(mai_mai_n297_));
  NA2        m0269(.A(mai_mai_n297_), .B(mai_mai_n259_), .Y(mai_mai_n298_));
  NOi32      m0270(.An(j), .Bn(m), .C(i), .Y(mai_mai_n299_));
  NA3        m0271(.A(mai_mai_n299_), .B(mai_mai_n245_), .C(mai_mai_n96_), .Y(mai_mai_n300_));
  AO210      m0272(.A0(mai_mai_n94_), .A1(mai_mai_n32_), .B0(mai_mai_n300_), .Y(mai_mai_n301_));
  NOi32      m0273(.An(e), .Bn(b), .C(a), .Y(mai_mai_n302_));
  NA2        m0274(.A(mai_mai_n180_), .B(mai_mai_n35_), .Y(mai_mai_n303_));
  NA2        m0275(.A(mai_mai_n303_), .B(mai_mai_n302_), .Y(mai_mai_n304_));
  NO2        m0276(.A(mai_mai_n276_), .B(n), .Y(mai_mai_n305_));
  NA2        m0277(.A(mai_mai_n179_), .B(k), .Y(mai_mai_n306_));
  NA3        m0278(.A(m), .B(mai_mai_n95_), .C(mai_mai_n183_), .Y(mai_mai_n307_));
  NA4        m0279(.A(mai_mai_n177_), .B(mai_mai_n70_), .C(m), .D(mai_mai_n183_), .Y(mai_mai_n308_));
  NAi41      m0280(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n309_));
  NA2        m0281(.A(mai_mai_n50_), .B(mai_mai_n96_), .Y(mai_mai_n310_));
  NO2        m0282(.A(mai_mai_n310_), .B(mai_mai_n309_), .Y(mai_mai_n311_));
  AOI220     m0283(.A0(mai_mai_n311_), .A1(b), .B0(mai_mai_n177_), .B1(mai_mai_n305_), .Y(mai_mai_n312_));
  NA4        m0284(.A(mai_mai_n312_), .B(mai_mai_n304_), .C(mai_mai_n301_), .D(mai_mai_n298_), .Y(mai_mai_n313_));
  NO4        m0285(.A(mai_mai_n313_), .B(mai_mai_n294_), .C(mai_mai_n285_), .D(mai_mai_n279_), .Y(mai_mai_n314_));
  NA4        m0286(.A(mai_mai_n314_), .B(mai_mai_n264_), .C(mai_mai_n226_), .D(mai_mai_n173_), .Y(mai10));
  NA3        m0287(.A(m), .B(k), .C(i), .Y(mai_mai_n316_));
  NO2        m0288(.A(mai_mai_n316_), .B(mai_mai_n184_), .Y(mai_mai_n317_));
  NOi21      m0289(.An(e), .B(f), .Y(mai_mai_n318_));
  NO4        m0290(.A(mai_mai_n129_), .B(mai_mai_n318_), .C(n), .D(mai_mai_n93_), .Y(mai_mai_n319_));
  NAi31      m0291(.An(b), .B(f), .C(c), .Y(mai_mai_n320_));
  INV        m0292(.A(mai_mai_n320_), .Y(mai_mai_n321_));
  NOi32      m0293(.An(k), .Bn(h), .C(j), .Y(mai_mai_n322_));
  NA2        m0294(.A(mai_mai_n322_), .B(mai_mai_n191_), .Y(mai_mai_n323_));
  NA2        m0295(.A(mai_mai_n138_), .B(mai_mai_n323_), .Y(mai_mai_n324_));
  AOI220     m0296(.A0(mai_mai_n324_), .A1(mai_mai_n321_), .B0(mai_mai_n319_), .B1(mai_mai_n317_), .Y(mai_mai_n325_));
  NO3        m0297(.A(n), .B(m), .C(k), .Y(mai_mai_n326_));
  NA2        m0298(.A(mai_mai_n326_), .B(h), .Y(mai_mai_n327_));
  NO3        m0299(.A(mai_mai_n327_), .B(mai_mai_n129_), .C(mai_mai_n183_), .Y(mai_mai_n328_));
  OR2        m0300(.A(m), .B(k), .Y(mai_mai_n329_));
  NO2        m0301(.A(mai_mai_n148_), .B(mai_mai_n329_), .Y(mai_mai_n330_));
  NA4        m0302(.A(n), .B(f), .C(c), .D(mai_mai_n98_), .Y(mai_mai_n331_));
  NOi21      m0303(.An(mai_mai_n330_), .B(mai_mai_n331_), .Y(mai_mai_n332_));
  NOi32      m0304(.An(d), .Bn(a), .C(c), .Y(mai_mai_n333_));
  NA2        m0305(.A(mai_mai_n333_), .B(mai_mai_n156_), .Y(mai_mai_n334_));
  NAi21      m0306(.An(i), .B(m), .Y(mai_mai_n335_));
  NAi31      m0307(.An(k), .B(m), .C(j), .Y(mai_mai_n336_));
  NO3        m0308(.A(mai_mai_n336_), .B(mai_mai_n335_), .C(n), .Y(mai_mai_n337_));
  NOi21      m0309(.An(mai_mai_n337_), .B(mai_mai_n334_), .Y(mai_mai_n338_));
  NO3        m0310(.A(mai_mai_n338_), .B(mai_mai_n332_), .C(mai_mai_n328_), .Y(mai_mai_n339_));
  NO2        m0311(.A(mai_mai_n331_), .B(mai_mai_n252_), .Y(mai_mai_n340_));
  NOi32      m0312(.An(f), .Bn(d), .C(c), .Y(mai_mai_n341_));
  AOI210     m0313(.A0(mai_mai_n341_), .A1(mai_mai_n258_), .B0(mai_mai_n340_), .Y(mai_mai_n342_));
  NA3        m0314(.A(mai_mai_n342_), .B(mai_mai_n339_), .C(mai_mai_n325_), .Y(mai_mai_n343_));
  NO2        m0315(.A(mai_mai_n54_), .B(mai_mai_n98_), .Y(mai_mai_n344_));
  NA2        m0316(.A(mai_mai_n214_), .B(mai_mai_n344_), .Y(mai_mai_n345_));
  INV        m0317(.A(e), .Y(mai_mai_n346_));
  NA2        m0318(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n347_));
  OAI220     m0319(.A0(mai_mai_n347_), .A1(mai_mai_n174_), .B0(mai_mai_n178_), .B1(mai_mai_n346_), .Y(mai_mai_n348_));
  NA3        m0320(.A(e), .B(mai_mai_n177_), .C(i), .Y(mai_mai_n349_));
  INV        m0321(.A(mai_mai_n349_), .Y(mai_mai_n350_));
  INV        m0322(.A(mai_mai_n83_), .Y(mai_mai_n351_));
  NO3        m0323(.A(mai_mai_n351_), .B(mai_mai_n350_), .C(mai_mai_n348_), .Y(mai_mai_n352_));
  NOi32      m0324(.An(h), .Bn(e), .C(m), .Y(mai_mai_n353_));
  NA3        m0325(.A(mai_mai_n353_), .B(mai_mai_n246_), .C(m), .Y(mai_mai_n354_));
  NOi21      m0326(.An(m), .B(h), .Y(mai_mai_n355_));
  AN3        m0327(.A(m), .B(l), .C(i), .Y(mai_mai_n356_));
  NA3        m0328(.A(mai_mai_n356_), .B(mai_mai_n355_), .C(e), .Y(mai_mai_n357_));
  AN3        m0329(.A(h), .B(m), .C(e), .Y(mai_mai_n358_));
  NA2        m0330(.A(mai_mai_n358_), .B(mai_mai_n80_), .Y(mai_mai_n359_));
  AN3        m0331(.A(mai_mai_n359_), .B(mai_mai_n357_), .C(mai_mai_n354_), .Y(mai_mai_n360_));
  AOI210     m0332(.A0(mai_mai_n360_), .A1(mai_mai_n352_), .B0(mai_mai_n345_), .Y(mai_mai_n361_));
  NA3        m0333(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n362_));
  NO2        m0334(.A(mai_mai_n362_), .B(mai_mai_n345_), .Y(mai_mai_n363_));
  NA3        m0335(.A(mai_mai_n333_), .B(mai_mai_n156_), .C(mai_mai_n67_), .Y(mai_mai_n364_));
  NAi31      m0336(.An(b), .B(c), .C(a), .Y(mai_mai_n365_));
  NO2        m0337(.A(mai_mai_n365_), .B(n), .Y(mai_mai_n366_));
  NO3        m0338(.A(mai_mai_n363_), .B(mai_mai_n361_), .C(mai_mai_n343_), .Y(mai_mai_n367_));
  NO2        m0339(.A(mai_mai_n233_), .B(c), .Y(mai_mai_n368_));
  NOi21      m0340(.An(a), .B(n), .Y(mai_mai_n369_));
  NOi21      m0341(.An(d), .B(c), .Y(mai_mai_n370_));
  NA2        m0342(.A(mai_mai_n370_), .B(mai_mai_n369_), .Y(mai_mai_n371_));
  NA3        m0343(.A(i), .B(m), .C(f), .Y(mai_mai_n372_));
  OR2        m0344(.A(mai_mai_n372_), .B(mai_mai_n61_), .Y(mai_mai_n373_));
  NA3        m0345(.A(mai_mai_n356_), .B(mai_mai_n355_), .C(mai_mai_n156_), .Y(mai_mai_n374_));
  AOI210     m0346(.A0(mai_mai_n374_), .A1(mai_mai_n373_), .B0(mai_mai_n371_), .Y(mai_mai_n375_));
  INV        m0347(.A(mai_mai_n375_), .Y(mai_mai_n376_));
  OR2        m0348(.A(n), .B(m), .Y(mai_mai_n377_));
  NO2        m0349(.A(mai_mai_n377_), .B(mai_mai_n130_), .Y(mai_mai_n378_));
  NO2        m0350(.A(mai_mai_n157_), .B(mai_mai_n126_), .Y(mai_mai_n379_));
  OAI210     m0351(.A0(mai_mai_n378_), .A1(mai_mai_n150_), .B0(mai_mai_n379_), .Y(mai_mai_n380_));
  NO2        m0352(.A(mai_mai_n365_), .B(mai_mai_n49_), .Y(mai_mai_n381_));
  NAi21      m0353(.An(k), .B(j), .Y(mai_mai_n382_));
  NAi21      m0354(.An(e), .B(d), .Y(mai_mai_n383_));
  INV        m0355(.A(mai_mai_n383_), .Y(mai_mai_n384_));
  NO2        m0356(.A(mai_mai_n216_), .B(mai_mai_n183_), .Y(mai_mai_n385_));
  NA3        m0357(.A(mai_mai_n385_), .B(mai_mai_n384_), .C(mai_mai_n197_), .Y(mai_mai_n386_));
  NA2        m0358(.A(mai_mai_n386_), .B(mai_mai_n380_), .Y(mai_mai_n387_));
  NO2        m0359(.A(mai_mai_n283_), .B(mai_mai_n183_), .Y(mai_mai_n388_));
  NAi31      m0360(.An(m), .B(f), .C(c), .Y(mai_mai_n389_));
  NOi31      m0361(.An(mai_mai_n376_), .B(mai_mai_n388_), .C(mai_mai_n387_), .Y(mai_mai_n390_));
  NOi32      m0362(.An(c), .Bn(a), .C(b), .Y(mai_mai_n391_));
  NA2        m0363(.A(mai_mai_n391_), .B(mai_mai_n96_), .Y(mai_mai_n392_));
  AN2        m0364(.A(e), .B(d), .Y(mai_mai_n393_));
  NO2        m0365(.A(mai_mai_n112_), .B(mai_mai_n41_), .Y(mai_mai_n394_));
  NO2        m0366(.A(mai_mai_n59_), .B(e), .Y(mai_mai_n395_));
  NOi31      m0367(.An(j), .B(k), .C(i), .Y(mai_mai_n396_));
  NOi21      m0368(.An(mai_mai_n142_), .B(mai_mai_n396_), .Y(mai_mai_n397_));
  NA4        m0369(.A(mai_mai_n271_), .B(mai_mai_n397_), .C(mai_mai_n223_), .D(mai_mai_n101_), .Y(mai_mai_n398_));
  AOI210     m0370(.A0(mai_mai_n398_), .A1(mai_mai_n395_), .B0(mai_mai_n394_), .Y(mai_mai_n399_));
  NO2        m0371(.A(mai_mai_n399_), .B(mai_mai_n392_), .Y(mai_mai_n400_));
  NOi21      m0372(.An(a), .B(b), .Y(mai_mai_n401_));
  NA3        m0373(.A(e), .B(d), .C(c), .Y(mai_mai_n402_));
  NAi21      m0374(.An(mai_mai_n402_), .B(mai_mai_n401_), .Y(mai_mai_n403_));
  AOI210     m0375(.A0(mai_mai_n227_), .A1(mai_mai_n180_), .B0(mai_mai_n403_), .Y(mai_mai_n404_));
  NA2        m0376(.A(mai_mai_n321_), .B(mai_mai_n131_), .Y(mai_mai_n405_));
  OR2        m0377(.A(k), .B(j), .Y(mai_mai_n406_));
  NA2        m0378(.A(l), .B(k), .Y(mai_mai_n407_));
  OR3        m0379(.A(mai_mai_n1278_), .B(mai_mai_n123_), .C(mai_mai_n115_), .Y(mai_mai_n408_));
  INV        m0380(.A(mai_mai_n109_), .Y(mai_mai_n409_));
  NA2        m0381(.A(mai_mai_n333_), .B(mai_mai_n96_), .Y(mai_mai_n410_));
  NO4        m0382(.A(mai_mai_n410_), .B(mai_mai_n77_), .C(mai_mai_n95_), .D(e), .Y(mai_mai_n411_));
  NO3        m0383(.A(mai_mai_n364_), .B(mai_mai_n74_), .C(mai_mai_n112_), .Y(mai_mai_n412_));
  NO2        m0384(.A(mai_mai_n412_), .B(mai_mai_n409_), .Y(mai_mai_n413_));
  NA3        m0385(.A(mai_mai_n413_), .B(mai_mai_n408_), .C(mai_mai_n405_), .Y(mai_mai_n414_));
  NO3        m0386(.A(mai_mai_n414_), .B(mai_mai_n404_), .C(mai_mai_n400_), .Y(mai_mai_n415_));
  NOi21      m0387(.An(d), .B(e), .Y(mai_mai_n416_));
  NAi31      m0388(.An(j), .B(l), .C(i), .Y(mai_mai_n417_));
  INV        m0389(.A(mai_mai_n86_), .Y(mai_mai_n418_));
  NO2        m0390(.A(mai_mai_n334_), .B(mai_mai_n175_), .Y(mai_mai_n419_));
  INV        m0391(.A(mai_mai_n419_), .Y(mai_mai_n420_));
  NA2        m0392(.A(mai_mai_n420_), .B(mai_mai_n209_), .Y(mai_mai_n421_));
  OAI210     m0393(.A0(mai_mai_n108_), .A1(mai_mai_n107_), .B0(n), .Y(mai_mai_n422_));
  NO2        m0394(.A(mai_mai_n422_), .B(mai_mai_n112_), .Y(mai_mai_n423_));
  OA210      m0395(.A0(mai_mai_n210_), .A1(mai_mai_n423_), .B0(mai_mai_n166_), .Y(mai_mai_n424_));
  XO2        m0396(.A(i), .B(h), .Y(mai_mai_n425_));
  BUFFER     m0397(.A(mai_mai_n253_), .Y(mai_mai_n426_));
  NAi31      m0398(.An(c), .B(f), .C(d), .Y(mai_mai_n427_));
  AOI210     m0399(.A0(mai_mai_n236_), .A1(mai_mai_n169_), .B0(mai_mai_n427_), .Y(mai_mai_n428_));
  NA3        m0400(.A(mai_mai_n319_), .B(mai_mai_n80_), .C(mai_mai_n79_), .Y(mai_mai_n429_));
  NA2        m0401(.A(mai_mai_n198_), .B(mai_mai_n91_), .Y(mai_mai_n430_));
  AOI210     m0402(.A0(mai_mai_n430_), .A1(mai_mai_n155_), .B0(mai_mai_n427_), .Y(mai_mai_n431_));
  AOI210     m0403(.A0(mai_mai_n300_), .A1(mai_mai_n35_), .B0(mai_mai_n403_), .Y(mai_mai_n432_));
  NOi31      m0404(.An(mai_mai_n429_), .B(mai_mai_n432_), .C(mai_mai_n431_), .Y(mai_mai_n433_));
  NA3        m0405(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n434_));
  NO2        m0406(.A(mai_mai_n434_), .B(mai_mai_n371_), .Y(mai_mai_n435_));
  INV        m0407(.A(mai_mai_n249_), .Y(mai_mai_n436_));
  NA2        m0408(.A(mai_mai_n436_), .B(mai_mai_n433_), .Y(mai_mai_n437_));
  NO3        m0409(.A(mai_mai_n437_), .B(mai_mai_n424_), .C(mai_mai_n421_), .Y(mai_mai_n438_));
  NA4        m0410(.A(mai_mai_n438_), .B(mai_mai_n415_), .C(mai_mai_n390_), .D(mai_mai_n367_), .Y(mai11));
  NO2        m0411(.A(mai_mai_n62_), .B(f), .Y(mai_mai_n440_));
  NA2        m0412(.A(j), .B(m), .Y(mai_mai_n441_));
  NAi31      m0413(.An(i), .B(m), .C(l), .Y(mai_mai_n442_));
  NA3        m0414(.A(m), .B(k), .C(j), .Y(mai_mai_n443_));
  OAI220     m0415(.A0(mai_mai_n443_), .A1(mai_mai_n112_), .B0(mai_mai_n442_), .B1(mai_mai_n441_), .Y(mai_mai_n444_));
  NA2        m0416(.A(mai_mai_n444_), .B(mai_mai_n440_), .Y(mai_mai_n445_));
  NA2        m0417(.A(mai_mai_n222_), .B(mai_mai_n96_), .Y(mai_mai_n446_));
  NA2        m0418(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n447_));
  NAi31      m0419(.An(d), .B(e), .C(a), .Y(mai_mai_n448_));
  NO2        m0420(.A(mai_mai_n448_), .B(n), .Y(mai_mai_n449_));
  NA2        m0421(.A(mai_mai_n449_), .B(mai_mai_n84_), .Y(mai_mai_n450_));
  NAi41      m0422(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n451_));
  AN2        m0423(.A(mai_mai_n451_), .B(mai_mai_n309_), .Y(mai_mai_n452_));
  AOI210     m0424(.A0(mai_mai_n452_), .A1(mai_mai_n334_), .B0(mai_mai_n229_), .Y(mai_mai_n453_));
  NA2        m0425(.A(j), .B(i), .Y(mai_mai_n454_));
  NAi31      m0426(.An(n), .B(m), .C(k), .Y(mai_mai_n455_));
  NO3        m0427(.A(mai_mai_n455_), .B(mai_mai_n454_), .C(mai_mai_n95_), .Y(mai_mai_n456_));
  NO4        m0428(.A(n), .B(d), .C(mai_mai_n98_), .D(a), .Y(mai_mai_n457_));
  OR2        m0429(.A(n), .B(c), .Y(mai_mai_n458_));
  NO2        m0430(.A(mai_mai_n458_), .B(mai_mai_n128_), .Y(mai_mai_n459_));
  NO2        m0431(.A(mai_mai_n459_), .B(mai_mai_n457_), .Y(mai_mai_n460_));
  NOi32      m0432(.An(m), .Bn(f), .C(i), .Y(mai_mai_n461_));
  AOI220     m0433(.A0(mai_mai_n461_), .A1(mai_mai_n82_), .B0(mai_mai_n444_), .B1(f), .Y(mai_mai_n462_));
  NO2        m0434(.A(mai_mai_n231_), .B(mai_mai_n49_), .Y(mai_mai_n463_));
  NO2        m0435(.A(mai_mai_n462_), .B(mai_mai_n460_), .Y(mai_mai_n464_));
  AOI210     m0436(.A0(mai_mai_n456_), .A1(mai_mai_n453_), .B0(mai_mai_n464_), .Y(mai_mai_n465_));
  NA2        m0437(.A(mai_mai_n120_), .B(mai_mai_n34_), .Y(mai_mai_n466_));
  OAI220     m0438(.A0(mai_mai_n466_), .A1(m), .B0(mai_mai_n447_), .B1(mai_mai_n204_), .Y(mai_mai_n467_));
  NOi41      m0439(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n468_));
  NAi32      m0440(.An(e), .Bn(b), .C(c), .Y(mai_mai_n469_));
  AN2        m0441(.A(mai_mai_n287_), .B(mai_mai_n268_), .Y(mai_mai_n470_));
  OA210      m0442(.A0(n), .A1(mai_mai_n468_), .B0(mai_mai_n467_), .Y(mai_mai_n471_));
  OAI220     m0443(.A0(mai_mai_n336_), .A1(mai_mai_n335_), .B0(mai_mai_n442_), .B1(mai_mai_n441_), .Y(mai_mai_n472_));
  NAi31      m0444(.An(d), .B(c), .C(a), .Y(mai_mai_n473_));
  NO2        m0445(.A(mai_mai_n473_), .B(n), .Y(mai_mai_n474_));
  NA3        m0446(.A(mai_mai_n474_), .B(mai_mai_n472_), .C(e), .Y(mai_mai_n475_));
  NO3        m0447(.A(mai_mai_n56_), .B(mai_mai_n49_), .C(mai_mai_n184_), .Y(mai_mai_n476_));
  NO2        m0448(.A(mai_mai_n201_), .B(mai_mai_n93_), .Y(mai_mai_n477_));
  OAI210     m0449(.A0(mai_mai_n476_), .A1(mai_mai_n337_), .B0(mai_mai_n477_), .Y(mai_mai_n478_));
  NA2        m0450(.A(mai_mai_n478_), .B(mai_mai_n475_), .Y(mai_mai_n479_));
  NO2        m0451(.A(mai_mai_n233_), .B(n), .Y(mai_mai_n480_));
  NO2        m0452(.A(mai_mai_n366_), .B(mai_mai_n480_), .Y(mai_mai_n481_));
  NA2        m0453(.A(mai_mai_n472_), .B(f), .Y(mai_mai_n482_));
  NAi32      m0454(.An(d), .Bn(a), .C(b), .Y(mai_mai_n483_));
  NA2        m0455(.A(h), .B(f), .Y(mai_mai_n484_));
  NO2        m0456(.A(mai_mai_n484_), .B(mai_mai_n77_), .Y(mai_mai_n485_));
  NO2        m0457(.A(mai_mai_n482_), .B(mai_mai_n481_), .Y(mai_mai_n486_));
  NA3        m0458(.A(f), .B(d), .C(b), .Y(mai_mai_n487_));
  NO3        m0459(.A(mai_mai_n486_), .B(mai_mai_n479_), .C(mai_mai_n471_), .Y(mai_mai_n488_));
  AN4        m0460(.A(mai_mai_n488_), .B(mai_mai_n465_), .C(mai_mai_n450_), .D(mai_mai_n445_), .Y(mai_mai_n489_));
  INV        m0461(.A(k), .Y(mai_mai_n490_));
  NA3        m0462(.A(l), .B(mai_mai_n490_), .C(i), .Y(mai_mai_n491_));
  INV        m0463(.A(mai_mai_n491_), .Y(mai_mai_n492_));
  NA3        m0464(.A(mai_mai_n333_), .B(mai_mai_n156_), .C(mai_mai_n96_), .Y(mai_mai_n493_));
  NAi32      m0465(.An(h), .Bn(f), .C(m), .Y(mai_mai_n494_));
  NAi41      m0466(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n495_));
  OAI210     m0467(.A0(mai_mai_n448_), .A1(n), .B0(mai_mai_n495_), .Y(mai_mai_n496_));
  NA2        m0468(.A(mai_mai_n496_), .B(m), .Y(mai_mai_n497_));
  NAi31      m0469(.An(h), .B(m), .C(f), .Y(mai_mai_n498_));
  OR3        m0470(.A(mai_mai_n498_), .B(mai_mai_n233_), .C(mai_mai_n49_), .Y(mai_mai_n499_));
  NA4        m0471(.A(mai_mai_n355_), .B(mai_mai_n103_), .C(mai_mai_n96_), .D(e), .Y(mai_mai_n500_));
  AN2        m0472(.A(mai_mai_n500_), .B(mai_mai_n499_), .Y(mai_mai_n501_));
  OA210      m0473(.A0(mai_mai_n497_), .A1(mai_mai_n494_), .B0(mai_mai_n501_), .Y(mai_mai_n502_));
  NO2        m0474(.A(mai_mai_n494_), .B(mai_mai_n62_), .Y(mai_mai_n503_));
  NO4        m0475(.A(mai_mai_n498_), .B(mai_mai_n458_), .C(mai_mai_n128_), .D(mai_mai_n63_), .Y(mai_mai_n504_));
  OR2        m0476(.A(mai_mai_n504_), .B(mai_mai_n503_), .Y(mai_mai_n505_));
  NAi31      m0477(.An(mai_mai_n505_), .B(mai_mai_n502_), .C(mai_mai_n493_), .Y(mai_mai_n506_));
  NAi31      m0478(.An(f), .B(h), .C(m), .Y(mai_mai_n507_));
  NOi32      m0479(.An(b), .Bn(a), .C(c), .Y(mai_mai_n508_));
  NOi31      m0480(.An(mai_mai_n508_), .B(mai_mai_n295_), .C(mai_mai_n60_), .Y(mai_mai_n509_));
  NOi32      m0481(.An(d), .Bn(a), .C(e), .Y(mai_mai_n510_));
  NA2        m0482(.A(mai_mai_n510_), .B(mai_mai_n96_), .Y(mai_mai_n511_));
  NO2        m0483(.A(n), .B(c), .Y(mai_mai_n512_));
  NA3        m0484(.A(mai_mai_n512_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n513_));
  NOi32      m0485(.An(e), .Bn(a), .C(d), .Y(mai_mai_n514_));
  AOI210     m0486(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n514_), .Y(mai_mai_n515_));
  AOI210     m0487(.A0(mai_mai_n515_), .A1(mai_mai_n183_), .B0(mai_mai_n466_), .Y(mai_mai_n516_));
  AOI210     m0488(.A0(mai_mai_n516_), .A1(mai_mai_n96_), .B0(mai_mai_n509_), .Y(mai_mai_n517_));
  INV        m0489(.A(mai_mai_n517_), .Y(mai_mai_n518_));
  AOI210     m0490(.A0(mai_mai_n506_), .A1(mai_mai_n492_), .B0(mai_mai_n518_), .Y(mai_mai_n519_));
  NO2        m0491(.A(mai_mai_n266_), .B(mai_mai_n55_), .Y(mai_mai_n520_));
  NA3        m0492(.A(mai_mai_n427_), .B(mai_mai_n146_), .C(mai_mai_n145_), .Y(mai_mai_n521_));
  NA2        m0493(.A(mai_mai_n389_), .B(mai_mai_n201_), .Y(mai_mai_n522_));
  OR2        m0494(.A(mai_mai_n522_), .B(mai_mai_n521_), .Y(mai_mai_n523_));
  NA2        m0495(.A(mai_mai_n64_), .B(mai_mai_n96_), .Y(mai_mai_n524_));
  NO2        m0496(.A(mai_mai_n524_), .B(mai_mai_n45_), .Y(mai_mai_n525_));
  AOI220     m0497(.A0(mai_mai_n525_), .A1(mai_mai_n453_), .B0(mai_mai_n523_), .B1(mai_mai_n520_), .Y(mai_mai_n526_));
  NO2        m0498(.A(mai_mai_n526_), .B(mai_mai_n70_), .Y(mai_mai_n527_));
  NOi32      m0499(.An(e), .Bn(c), .C(f), .Y(mai_mai_n528_));
  NOi21      m0500(.An(f), .B(m), .Y(mai_mai_n529_));
  NO2        m0501(.A(mai_mai_n529_), .B(mai_mai_n181_), .Y(mai_mai_n530_));
  AOI220     m0502(.A0(mai_mai_n530_), .A1(mai_mai_n330_), .B0(mai_mai_n528_), .B1(mai_mai_n150_), .Y(mai_mai_n531_));
  NA2        m0503(.A(mai_mai_n531_), .B(mai_mai_n153_), .Y(mai_mai_n532_));
  AOI210     m0504(.A0(mai_mai_n452_), .A1(mai_mai_n334_), .B0(mai_mai_n254_), .Y(mai_mai_n533_));
  NAi21      m0505(.An(k), .B(h), .Y(mai_mai_n534_));
  NO2        m0506(.A(mai_mai_n534_), .B(mai_mai_n224_), .Y(mai_mai_n535_));
  NA2        m0507(.A(mai_mai_n535_), .B(j), .Y(mai_mai_n536_));
  OR2        m0508(.A(mai_mai_n536_), .B(mai_mai_n497_), .Y(mai_mai_n537_));
  NOi31      m0509(.An(m), .B(n), .C(k), .Y(mai_mai_n538_));
  NA2        m0510(.A(j), .B(mai_mai_n538_), .Y(mai_mai_n539_));
  AOI210     m0511(.A0(mai_mai_n334_), .A1(mai_mai_n309_), .B0(mai_mai_n254_), .Y(mai_mai_n540_));
  NAi21      m0512(.An(mai_mai_n539_), .B(mai_mai_n540_), .Y(mai_mai_n541_));
  NO2        m0513(.A(mai_mai_n233_), .B(mai_mai_n49_), .Y(mai_mai_n542_));
  NO2        m0514(.A(mai_mai_n448_), .B(mai_mai_n49_), .Y(mai_mai_n543_));
  NA2        m0515(.A(mai_mai_n542_), .B(mai_mai_n485_), .Y(mai_mai_n544_));
  NA3        m0516(.A(mai_mai_n544_), .B(mai_mai_n541_), .C(mai_mai_n537_), .Y(mai_mai_n545_));
  NA2        m0517(.A(mai_mai_n91_), .B(mai_mai_n36_), .Y(mai_mai_n546_));
  NO2        m0518(.A(k), .B(mai_mai_n184_), .Y(mai_mai_n547_));
  INV        m0519(.A(mai_mai_n302_), .Y(mai_mai_n548_));
  NO2        m0520(.A(mai_mai_n548_), .B(n), .Y(mai_mai_n549_));
  NAi31      m0521(.An(mai_mai_n546_), .B(mai_mai_n549_), .C(mai_mai_n547_), .Y(mai_mai_n550_));
  AN3        m0522(.A(f), .B(d), .C(b), .Y(mai_mai_n551_));
  NO2        m0523(.A(mai_mai_n551_), .B(mai_mai_n111_), .Y(mai_mai_n552_));
  NA3        m0524(.A(mai_mai_n425_), .B(mai_mai_n137_), .C(mai_mai_n184_), .Y(mai_mai_n553_));
  AOI210     m0525(.A0(mai_mai_n552_), .A1(mai_mai_n203_), .B0(mai_mai_n553_), .Y(mai_mai_n554_));
  NAi31      m0526(.An(m), .B(n), .C(k), .Y(mai_mai_n555_));
  NA2        m0527(.A(mai_mai_n554_), .B(j), .Y(mai_mai_n556_));
  NA2        m0528(.A(mai_mai_n556_), .B(mai_mai_n550_), .Y(mai_mai_n557_));
  NO4        m0529(.A(mai_mai_n557_), .B(mai_mai_n545_), .C(mai_mai_n532_), .D(mai_mai_n527_), .Y(mai_mai_n558_));
  NAi31      m0530(.An(m), .B(h), .C(f), .Y(mai_mai_n559_));
  OR3        m0531(.A(mai_mai_n559_), .B(mai_mai_n233_), .C(n), .Y(mai_mai_n560_));
  OA210      m0532(.A0(mai_mai_n448_), .A1(n), .B0(mai_mai_n495_), .Y(mai_mai_n561_));
  NA3        m0533(.A(mai_mai_n353_), .B(mai_mai_n103_), .C(mai_mai_n67_), .Y(mai_mai_n562_));
  OAI210     m0534(.A0(mai_mai_n561_), .A1(mai_mai_n73_), .B0(mai_mai_n562_), .Y(mai_mai_n563_));
  NOi21      m0535(.An(mai_mai_n560_), .B(mai_mai_n563_), .Y(mai_mai_n564_));
  NO2        m0536(.A(mai_mai_n564_), .B(mai_mai_n443_), .Y(mai_mai_n565_));
  NO3        m0537(.A(m), .B(mai_mai_n183_), .C(mai_mai_n51_), .Y(mai_mai_n566_));
  NO2        m0538(.A(mai_mai_n430_), .B(mai_mai_n70_), .Y(mai_mai_n567_));
  OAI210     m0539(.A0(mai_mai_n567_), .A1(mai_mai_n330_), .B0(mai_mai_n566_), .Y(mai_mai_n568_));
  OR2        m0540(.A(mai_mai_n62_), .B(mai_mai_n63_), .Y(mai_mai_n569_));
  NA2        m0541(.A(mai_mai_n508_), .B(mai_mai_n289_), .Y(mai_mai_n570_));
  OA220      m0542(.A0(mai_mai_n539_), .A1(mai_mai_n570_), .B0(mai_mai_n536_), .B1(mai_mai_n569_), .Y(mai_mai_n571_));
  NA3        m0543(.A(mai_mai_n440_), .B(mai_mai_n82_), .C(mai_mai_n81_), .Y(mai_mai_n572_));
  NA2        m0544(.A(h), .B(mai_mai_n37_), .Y(mai_mai_n573_));
  NA2        m0545(.A(mai_mai_n82_), .B(mai_mai_n46_), .Y(mai_mai_n574_));
  OAI220     m0546(.A0(mai_mai_n574_), .A1(mai_mai_n280_), .B0(mai_mai_n573_), .B1(mai_mai_n392_), .Y(mai_mai_n575_));
  AOI210     m0547(.A0(mai_mai_n483_), .A1(mai_mai_n365_), .B0(mai_mai_n49_), .Y(mai_mai_n576_));
  NO2        m0548(.A(mai_mai_n498_), .B(mai_mai_n491_), .Y(mai_mai_n577_));
  AOI210     m0549(.A0(mai_mai_n577_), .A1(mai_mai_n576_), .B0(mai_mai_n575_), .Y(mai_mai_n578_));
  NA4        m0550(.A(mai_mai_n578_), .B(mai_mai_n572_), .C(mai_mai_n571_), .D(mai_mai_n568_), .Y(mai_mai_n579_));
  NO2        m0551(.A(mai_mai_n215_), .B(f), .Y(mai_mai_n580_));
  NA2        m0552(.A(mai_mai_n277_), .B(mai_mai_n120_), .Y(mai_mai_n581_));
  NA2        m0553(.A(mai_mai_n302_), .B(mai_mai_n96_), .Y(mai_mai_n582_));
  OA220      m0554(.A0(mai_mai_n582_), .A1(mai_mai_n466_), .B0(mai_mai_n300_), .B1(mai_mai_n94_), .Y(mai_mai_n583_));
  OAI210     m0555(.A0(mai_mai_n581_), .A1(mai_mai_n529_), .B0(mai_mai_n583_), .Y(mai_mai_n584_));
  NO3        m0556(.A(mai_mai_n341_), .B(mai_mai_n166_), .C(mai_mai_n165_), .Y(mai_mai_n585_));
  NA2        m0557(.A(mai_mai_n585_), .B(mai_mai_n201_), .Y(mai_mai_n586_));
  NA3        m0558(.A(mai_mai_n586_), .B(mai_mai_n217_), .C(j), .Y(mai_mai_n587_));
  NA2        m0559(.A(mai_mai_n391_), .B(mai_mai_n67_), .Y(mai_mai_n588_));
  NA3        m0560(.A(mai_mai_n587_), .B(mai_mai_n429_), .C(mai_mai_n339_), .Y(mai_mai_n589_));
  NO4        m0561(.A(mai_mai_n589_), .B(mai_mai_n584_), .C(mai_mai_n579_), .D(mai_mai_n565_), .Y(mai_mai_n590_));
  NA4        m0562(.A(mai_mai_n590_), .B(mai_mai_n558_), .C(mai_mai_n519_), .D(mai_mai_n489_), .Y(mai08));
  NO2        m0563(.A(k), .B(h), .Y(mai_mai_n592_));
  AO210      m0564(.A0(mai_mai_n215_), .A1(mai_mai_n382_), .B0(mai_mai_n592_), .Y(mai_mai_n593_));
  NO2        m0565(.A(mai_mai_n593_), .B(mai_mai_n252_), .Y(mai_mai_n594_));
  NA2        m0566(.A(mai_mai_n528_), .B(mai_mai_n67_), .Y(mai_mai_n595_));
  NA2        m0567(.A(mai_mai_n595_), .B(mai_mai_n389_), .Y(mai_mai_n596_));
  AOI210     m0568(.A0(mai_mai_n596_), .A1(mai_mai_n594_), .B0(mai_mai_n412_), .Y(mai_mai_n597_));
  NA2        m0569(.A(mai_mai_n67_), .B(mai_mai_n93_), .Y(mai_mai_n598_));
  NO2        m0570(.A(mai_mai_n598_), .B(mai_mai_n52_), .Y(mai_mai_n599_));
  NA2        m0571(.A(mai_mai_n487_), .B(mai_mai_n203_), .Y(mai_mai_n600_));
  NA2        m0572(.A(mai_mai_n600_), .B(mai_mai_n291_), .Y(mai_mai_n601_));
  NA4        m0573(.A(mai_mai_n186_), .B(mai_mai_n120_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n602_));
  AN2        m0574(.A(l), .B(k), .Y(mai_mai_n603_));
  NA2        m0575(.A(mai_mai_n601_), .B(mai_mai_n597_), .Y(mai_mai_n604_));
  AN2        m0576(.A(mai_mai_n449_), .B(mai_mai_n78_), .Y(mai_mai_n605_));
  INV        m0577(.A(mai_mai_n435_), .Y(mai_mai_n606_));
  NO2        m0578(.A(mai_mai_n38_), .B(mai_mai_n183_), .Y(mai_mai_n607_));
  AOI220     m0579(.A0(mai_mai_n530_), .A1(mai_mai_n290_), .B0(mai_mai_n607_), .B1(mai_mai_n480_), .Y(mai_mai_n608_));
  NA2        m0580(.A(mai_mai_n608_), .B(mai_mai_n606_), .Y(mai_mai_n609_));
  NO2        m0581(.A(mai_mai_n452_), .B(mai_mai_n35_), .Y(mai_mai_n610_));
  NA2        m0582(.A(mai_mai_n469_), .B(mai_mai_n115_), .Y(mai_mai_n611_));
  NO2        m0583(.A(mai_mai_n407_), .B(mai_mai_n113_), .Y(mai_mai_n612_));
  AOI210     m0584(.A0(mai_mai_n612_), .A1(mai_mai_n611_), .B0(mai_mai_n610_), .Y(mai_mai_n613_));
  INV        m0585(.A(mai_mai_n613_), .Y(mai_mai_n614_));
  NA2        m0586(.A(mai_mai_n302_), .B(mai_mai_n43_), .Y(mai_mai_n615_));
  NA3        m0587(.A(mai_mai_n586_), .B(mai_mai_n282_), .C(mai_mai_n322_), .Y(mai_mai_n616_));
  NA2        m0588(.A(mai_mai_n603_), .B(mai_mai_n191_), .Y(mai_mai_n617_));
  NO2        m0589(.A(mai_mai_n617_), .B(mai_mai_n276_), .Y(mai_mai_n618_));
  AOI210     m0590(.A0(mai_mai_n618_), .A1(mai_mai_n580_), .B0(mai_mai_n411_), .Y(mai_mai_n619_));
  NA3        m0591(.A(m), .B(l), .C(k), .Y(mai_mai_n620_));
  AOI210     m0592(.A0(mai_mai_n562_), .A1(mai_mai_n560_), .B0(mai_mai_n620_), .Y(mai_mai_n621_));
  NO2        m0593(.A(mai_mai_n451_), .B(mai_mai_n229_), .Y(mai_mai_n622_));
  NOi21      m0594(.An(mai_mai_n622_), .B(mai_mai_n446_), .Y(mai_mai_n623_));
  NA4        m0595(.A(mai_mai_n96_), .B(l), .C(k), .D(mai_mai_n70_), .Y(mai_mai_n624_));
  NA3        m0596(.A(mai_mai_n103_), .B(e), .C(i), .Y(mai_mai_n625_));
  NO2        m0597(.A(mai_mai_n625_), .B(mai_mai_n624_), .Y(mai_mai_n626_));
  NO3        m0598(.A(mai_mai_n626_), .B(mai_mai_n623_), .C(mai_mai_n621_), .Y(mai_mai_n627_));
  NA4        m0599(.A(mai_mai_n627_), .B(mai_mai_n619_), .C(mai_mai_n616_), .D(mai_mai_n615_), .Y(mai_mai_n628_));
  NO4        m0600(.A(mai_mai_n628_), .B(mai_mai_n614_), .C(mai_mai_n609_), .D(mai_mai_n604_), .Y(mai_mai_n629_));
  NA2        m0601(.A(mai_mai_n530_), .B(mai_mai_n330_), .Y(mai_mai_n630_));
  NA2        m0602(.A(mai_mai_n543_), .B(m), .Y(mai_mai_n631_));
  NO3        m0603(.A(mai_mai_n334_), .B(mai_mai_n441_), .C(h), .Y(mai_mai_n632_));
  NA2        m0604(.A(mai_mai_n632_), .B(mai_mai_n96_), .Y(mai_mai_n633_));
  NA3        m0605(.A(mai_mai_n633_), .B(mai_mai_n631_), .C(mai_mai_n630_), .Y(mai_mai_n634_));
  NA2        m0606(.A(mai_mai_n603_), .B(mai_mai_n63_), .Y(mai_mai_n635_));
  NO3        m0607(.A(mai_mai_n585_), .B(mai_mai_n148_), .C(i), .Y(mai_mai_n636_));
  NOi21      m0608(.An(h), .B(j), .Y(mai_mai_n637_));
  NA2        m0609(.A(mai_mai_n637_), .B(f), .Y(mai_mai_n638_));
  INV        m0610(.A(mai_mai_n636_), .Y(mai_mai_n639_));
  OAI220     m0611(.A0(mai_mai_n639_), .A1(mai_mai_n635_), .B0(mai_mai_n501_), .B1(mai_mai_n56_), .Y(mai_mai_n640_));
  AOI210     m0612(.A0(mai_mai_n634_), .A1(l), .B0(mai_mai_n640_), .Y(mai_mai_n641_));
  NO2        m0613(.A(j), .B(i), .Y(mai_mai_n642_));
  NA2        m0614(.A(mai_mai_n65_), .B(l), .Y(mai_mai_n643_));
  NA2        m0615(.A(mai_mai_n642_), .B(mai_mai_n33_), .Y(mai_mai_n644_));
  INV        m0616(.A(mai_mai_n358_), .Y(mai_mai_n645_));
  OA220      m0617(.A0(mai_mai_n645_), .A1(mai_mai_n644_), .B0(mai_mai_n643_), .B1(mai_mai_n497_), .Y(mai_mai_n646_));
  NO3        m0618(.A(mai_mai_n129_), .B(mai_mai_n49_), .C(mai_mai_n93_), .Y(mai_mai_n647_));
  NO3        m0619(.A(mai_mai_n458_), .B(mai_mai_n128_), .C(mai_mai_n63_), .Y(mai_mai_n648_));
  NO2        m0620(.A(mai_mai_n407_), .B(mai_mai_n372_), .Y(mai_mai_n649_));
  OAI210     m0621(.A0(mai_mai_n648_), .A1(mai_mai_n647_), .B0(mai_mai_n649_), .Y(mai_mai_n650_));
  OAI210     m0622(.A0(mai_mai_n631_), .A1(mai_mai_n56_), .B0(mai_mai_n650_), .Y(mai_mai_n651_));
  NA2        m0623(.A(k), .B(j), .Y(mai_mai_n652_));
  NO3        m0624(.A(mai_mai_n252_), .B(mai_mai_n652_), .C(mai_mai_n40_), .Y(mai_mai_n653_));
  AN2        m0625(.A(mai_mai_n653_), .B(mai_mai_n81_), .Y(mai_mai_n654_));
  NO3        m0626(.A(mai_mai_n148_), .B(mai_mai_n329_), .C(mai_mai_n95_), .Y(mai_mai_n655_));
  NA2        m0627(.A(mai_mai_n655_), .B(mai_mai_n212_), .Y(mai_mai_n656_));
  NAi21      m0628(.An(mai_mai_n515_), .B(mai_mai_n75_), .Y(mai_mai_n657_));
  NA2        m0629(.A(mai_mai_n657_), .B(mai_mai_n656_), .Y(mai_mai_n658_));
  NO2        m0630(.A(mai_mai_n252_), .B(mai_mai_n116_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n659_), .B(mai_mai_n530_), .Y(mai_mai_n660_));
  NO2        m0632(.A(mai_mai_n498_), .B(mai_mai_n99_), .Y(mai_mai_n661_));
  OAI210     m0633(.A0(mai_mai_n661_), .A1(mai_mai_n649_), .B0(mai_mai_n576_), .Y(mai_mai_n662_));
  NA2        m0634(.A(mai_mai_n662_), .B(mai_mai_n660_), .Y(mai_mai_n663_));
  OR4        m0635(.A(mai_mai_n663_), .B(mai_mai_n658_), .C(mai_mai_n654_), .D(mai_mai_n651_), .Y(mai_mai_n664_));
  NA3        m0636(.A(f), .B(mai_mai_n470_), .C(mai_mai_n469_), .Y(mai_mai_n665_));
  NA4        m0637(.A(mai_mai_n665_), .B(mai_mai_n186_), .C(mai_mai_n382_), .D(mai_mai_n34_), .Y(mai_mai_n666_));
  OAI220     m0638(.A0(mai_mai_n602_), .A1(mai_mai_n595_), .B0(mai_mai_n280_), .B1(mai_mai_n38_), .Y(mai_mai_n667_));
  INV        m0639(.A(mai_mai_n667_), .Y(mai_mai_n668_));
  NA3        m0640(.A(mai_mai_n461_), .B(mai_mai_n246_), .C(h), .Y(mai_mai_n669_));
  NOi21      m0641(.An(mai_mai_n576_), .B(mai_mai_n669_), .Y(mai_mai_n670_));
  OAI220     m0642(.A0(mai_mai_n669_), .A1(mai_mai_n513_), .B0(mai_mai_n643_), .B1(mai_mai_n569_), .Y(mai_mai_n671_));
  INV        m0643(.A(mai_mai_n671_), .Y(mai_mai_n672_));
  NAi41      m0644(.An(mai_mai_n670_), .B(mai_mai_n672_), .C(mai_mai_n668_), .D(mai_mai_n666_), .Y(mai_mai_n673_));
  NA2        m0645(.A(mai_mai_n649_), .B(mai_mai_n542_), .Y(mai_mai_n674_));
  INV        m0646(.A(mai_mai_n284_), .Y(mai_mai_n675_));
  NA2        m0647(.A(mai_mai_n675_), .B(mai_mai_n674_), .Y(mai_mai_n676_));
  NOi41      m0648(.An(mai_mai_n646_), .B(mai_mai_n676_), .C(mai_mai_n673_), .D(mai_mai_n664_), .Y(mai_mai_n677_));
  OR2        m0649(.A(mai_mai_n602_), .B(mai_mai_n203_), .Y(mai_mai_n678_));
  INV        m0650(.A(mai_mai_n46_), .Y(mai_mai_n679_));
  NO3        m0651(.A(mai_mai_n679_), .B(mai_mai_n644_), .C(mai_mai_n233_), .Y(mai_mai_n680_));
  NO3        m0652(.A(mai_mai_n441_), .B(mai_mai_n76_), .C(h), .Y(mai_mai_n681_));
  AOI210     m0653(.A0(mai_mai_n681_), .A1(mai_mai_n599_), .B0(mai_mai_n680_), .Y(mai_mai_n682_));
  NA3        m0654(.A(mai_mai_n682_), .B(mai_mai_n678_), .C(mai_mai_n342_), .Y(mai_mai_n683_));
  OR2        m0655(.A(mai_mai_n559_), .B(mai_mai_n74_), .Y(mai_mai_n684_));
  NOi31      m0656(.An(b), .B(d), .C(a), .Y(mai_mai_n685_));
  NO2        m0657(.A(mai_mai_n685_), .B(mai_mai_n510_), .Y(mai_mai_n686_));
  NO2        m0658(.A(mai_mai_n686_), .B(n), .Y(mai_mai_n687_));
  NOi21      m0659(.An(mai_mai_n1283_), .B(mai_mai_n687_), .Y(mai_mai_n688_));
  NO2        m0660(.A(mai_mai_n688_), .B(mai_mai_n684_), .Y(mai_mai_n689_));
  NO3        m0661(.A(mai_mai_n529_), .B(mai_mai_n276_), .C(mai_mai_n99_), .Y(mai_mai_n690_));
  NOi21      m0662(.An(mai_mai_n690_), .B(mai_mai_n138_), .Y(mai_mai_n691_));
  INV        m0663(.A(mai_mai_n691_), .Y(mai_mai_n692_));
  OAI210     m0664(.A0(mai_mai_n602_), .A1(mai_mai_n331_), .B0(mai_mai_n692_), .Y(mai_mai_n693_));
  NO2        m0665(.A(mai_mai_n585_), .B(n), .Y(mai_mai_n694_));
  AOI220     m0666(.A0(mai_mai_n659_), .A1(mai_mai_n566_), .B0(mai_mai_n694_), .B1(mai_mai_n594_), .Y(mai_mai_n695_));
  NO2        m0667(.A(mai_mai_n272_), .B(mai_mai_n208_), .Y(mai_mai_n696_));
  OAI210     m0668(.A0(mai_mai_n78_), .A1(mai_mai_n75_), .B0(mai_mai_n696_), .Y(mai_mai_n697_));
  NA2        m0669(.A(mai_mai_n103_), .B(mai_mai_n67_), .Y(mai_mai_n698_));
  AOI210     m0670(.A0(mai_mai_n362_), .A1(mai_mai_n354_), .B0(mai_mai_n698_), .Y(mai_mai_n699_));
  NAi21      m0671(.An(mai_mai_n699_), .B(mai_mai_n697_), .Y(mai_mai_n700_));
  NA2        m0672(.A(mai_mai_n618_), .B(mai_mai_n34_), .Y(mai_mai_n701_));
  NAi21      m0673(.An(mai_mai_n624_), .B(mai_mai_n368_), .Y(mai_mai_n702_));
  NO2        m0674(.A(mai_mai_n229_), .B(i), .Y(mai_mai_n703_));
  OAI210     m0675(.A0(mai_mai_n504_), .A1(mai_mai_n503_), .B0(l), .Y(mai_mai_n704_));
  AN2        m0676(.A(mai_mai_n704_), .B(mai_mai_n702_), .Y(mai_mai_n705_));
  NAi41      m0677(.An(mai_mai_n700_), .B(mai_mai_n705_), .C(mai_mai_n701_), .D(mai_mai_n695_), .Y(mai_mai_n706_));
  NO4        m0678(.A(mai_mai_n706_), .B(mai_mai_n693_), .C(mai_mai_n689_), .D(mai_mai_n683_), .Y(mai_mai_n707_));
  NA4        m0679(.A(mai_mai_n707_), .B(mai_mai_n677_), .C(mai_mai_n641_), .D(mai_mai_n629_), .Y(mai09));
  INV        m0680(.A(mai_mai_n104_), .Y(mai_mai_n709_));
  NA2        m0681(.A(f), .B(e), .Y(mai_mai_n710_));
  NO2        m0682(.A(mai_mai_n196_), .B(mai_mai_n95_), .Y(mai_mai_n711_));
  NA4        m0683(.A(mai_mai_n260_), .B(mai_mai_n397_), .C(mai_mai_n223_), .D(mai_mai_n101_), .Y(mai_mai_n712_));
  AOI210     m0684(.A0(mai_mai_n712_), .A1(m), .B0(mai_mai_n394_), .Y(mai_mai_n713_));
  INV        m0685(.A(mai_mai_n710_), .Y(mai_mai_n714_));
  NA2        m0686(.A(mai_mai_n378_), .B(e), .Y(mai_mai_n715_));
  NO2        m0687(.A(mai_mai_n715_), .B(mai_mai_n427_), .Y(mai_mai_n716_));
  AOI210     m0688(.A0(mai_mai_n714_), .A1(mai_mai_n709_), .B0(mai_mai_n716_), .Y(mai_mai_n717_));
  NO2        m0689(.A(mai_mai_n178_), .B(mai_mai_n183_), .Y(mai_mai_n718_));
  NA3        m0690(.A(m), .B(l), .C(i), .Y(mai_mai_n719_));
  OAI220     m0691(.A0(mai_mai_n498_), .A1(mai_mai_n719_), .B0(mai_mai_n295_), .B1(mai_mai_n442_), .Y(mai_mai_n720_));
  NA4        m0692(.A(mai_mai_n71_), .B(mai_mai_n70_), .C(m), .D(f), .Y(mai_mai_n721_));
  NAi31      m0693(.An(mai_mai_n720_), .B(mai_mai_n721_), .C(mai_mai_n373_), .Y(mai_mai_n722_));
  OR2        m0694(.A(mai_mai_n722_), .B(mai_mai_n718_), .Y(mai_mai_n723_));
  NA3        m0695(.A(mai_mai_n684_), .B(mai_mai_n482_), .C(mai_mai_n434_), .Y(mai_mai_n724_));
  OA210      m0696(.A0(mai_mai_n724_), .A1(mai_mai_n723_), .B0(mai_mai_n687_), .Y(mai_mai_n725_));
  INV        m0697(.A(mai_mai_n108_), .Y(mai_mai_n726_));
  NO2        m0698(.A(mai_mai_n726_), .B(mai_mai_n507_), .Y(mai_mai_n727_));
  INV        m0699(.A(mai_mai_n280_), .Y(mai_mai_n728_));
  NA2        m0700(.A(mai_mai_n289_), .B(j), .Y(mai_mai_n729_));
  NA2        m0701(.A(mai_mai_n727_), .B(d), .Y(mai_mai_n730_));
  NA3        m0702(.A(h), .B(mai_mai_n163_), .C(mai_mai_n31_), .Y(mai_mai_n731_));
  NA3        m0703(.A(mai_mai_n731_), .B(mai_mai_n730_), .C(mai_mai_n531_), .Y(mai_mai_n732_));
  NO2        m0704(.A(mai_mai_n494_), .B(mai_mai_n417_), .Y(mai_mai_n733_));
  NA2        m0705(.A(mai_mai_n733_), .B(mai_mai_n163_), .Y(mai_mai_n734_));
  NOi21      m0706(.An(f), .B(d), .Y(mai_mai_n735_));
  NA2        m0707(.A(mai_mai_n735_), .B(m), .Y(mai_mai_n736_));
  NOi32      m0708(.An(m), .Bn(f), .C(d), .Y(mai_mai_n737_));
  NA4        m0709(.A(mai_mai_n737_), .B(mai_mai_n512_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n738_));
  AN2        m0710(.A(f), .B(d), .Y(mai_mai_n739_));
  NA3        m0711(.A(mai_mai_n401_), .B(mai_mai_n739_), .C(mai_mai_n67_), .Y(mai_mai_n740_));
  NO3        m0712(.A(mai_mai_n740_), .B(mai_mai_n63_), .C(mai_mai_n184_), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n240_), .B(mai_mai_n51_), .Y(mai_mai_n742_));
  NA2        m0714(.A(mai_mai_n100_), .B(mai_mai_n741_), .Y(mai_mai_n743_));
  NA3        m0715(.A(mai_mai_n743_), .B(mai_mai_n738_), .C(mai_mai_n734_), .Y(mai_mai_n744_));
  NO2        m0716(.A(mai_mai_n555_), .B(mai_mai_n276_), .Y(mai_mai_n745_));
  AN2        m0717(.A(mai_mai_n745_), .B(mai_mai_n580_), .Y(mai_mai_n746_));
  INV        m0718(.A(mai_mai_n746_), .Y(mai_mai_n747_));
  NA2        m0719(.A(mai_mai_n510_), .B(mai_mai_n67_), .Y(mai_mai_n748_));
  NO2        m0720(.A(mai_mai_n729_), .B(mai_mai_n748_), .Y(mai_mai_n749_));
  NA3        m0721(.A(mai_mai_n137_), .B(mai_mai_n91_), .C(mai_mai_n90_), .Y(mai_mai_n750_));
  NO2        m0722(.A(mai_mai_n287_), .B(mai_mai_n750_), .Y(mai_mai_n751_));
  NOi31      m0723(.An(mai_mai_n194_), .B(mai_mai_n751_), .C(mai_mai_n749_), .Y(mai_mai_n752_));
  NA2        m0724(.A(c), .B(mai_mai_n98_), .Y(mai_mai_n753_));
  NA3        m0725(.A(mai_mai_n98_), .B(mai_mai_n426_), .C(f), .Y(mai_mai_n754_));
  OR2        m0726(.A(mai_mai_n559_), .B(mai_mai_n455_), .Y(mai_mai_n755_));
  INV        m0727(.A(mai_mai_n755_), .Y(mai_mai_n756_));
  NA2        m0728(.A(mai_mai_n685_), .B(mai_mai_n756_), .Y(mai_mai_n757_));
  NA4        m0729(.A(mai_mai_n757_), .B(mai_mai_n754_), .C(mai_mai_n752_), .D(mai_mai_n747_), .Y(mai_mai_n758_));
  NO4        m0730(.A(mai_mai_n758_), .B(mai_mai_n744_), .C(mai_mai_n732_), .D(mai_mai_n725_), .Y(mai_mai_n759_));
  BUFFER     m0731(.A(mai_mai_n740_), .Y(mai_mai_n760_));
  NA2        m0732(.A(mai_mai_n711_), .B(m), .Y(mai_mai_n761_));
  AOI210     m0733(.A0(mai_mai_n761_), .A1(mai_mai_n247_), .B0(mai_mai_n760_), .Y(mai_mai_n762_));
  NO2        m0734(.A(mai_mai_n280_), .B(mai_mai_n721_), .Y(mai_mai_n763_));
  NA2        m0735(.A(e), .B(d), .Y(mai_mai_n764_));
  OAI220     m0736(.A0(mai_mai_n764_), .A1(c), .B0(mai_mai_n272_), .B1(d), .Y(mai_mai_n765_));
  NA3        m0737(.A(mai_mai_n765_), .B(mai_mai_n385_), .C(mai_mai_n425_), .Y(mai_mai_n766_));
  AOI210     m0738(.A0(mai_mai_n430_), .A1(mai_mai_n155_), .B0(mai_mai_n201_), .Y(mai_mai_n767_));
  AOI210     m0739(.A0(mai_mai_n530_), .A1(mai_mai_n290_), .B0(mai_mai_n767_), .Y(mai_mai_n768_));
  NA2        m0740(.A(mai_mai_n240_), .B(mai_mai_n142_), .Y(mai_mai_n769_));
  NA2        m0741(.A(mai_mai_n741_), .B(mai_mai_n769_), .Y(mai_mai_n770_));
  NA3        m0742(.A(mai_mai_n143_), .B(mai_mai_n68_), .C(mai_mai_n34_), .Y(mai_mai_n771_));
  NA4        m0743(.A(mai_mai_n771_), .B(mai_mai_n770_), .C(mai_mai_n768_), .D(mai_mai_n766_), .Y(mai_mai_n772_));
  NO3        m0744(.A(mai_mai_n772_), .B(mai_mai_n763_), .C(mai_mai_n762_), .Y(mai_mai_n773_));
  NA2        m0745(.A(d), .B(mai_mai_n31_), .Y(mai_mai_n774_));
  OR2        m0746(.A(mai_mai_n774_), .B(mai_mai_n187_), .Y(mai_mai_n775_));
  OAI210     m0747(.A0(mai_mai_n529_), .A1(mai_mai_n55_), .B0(mai_mai_n254_), .Y(mai_mai_n776_));
  AOI220     m0748(.A0(mai_mai_n776_), .A1(mai_mai_n745_), .B0(mai_mai_n520_), .B1(mai_mai_n528_), .Y(mai_mai_n777_));
  OAI210     m0749(.A0(mai_mai_n715_), .A1(mai_mai_n145_), .B0(mai_mai_n777_), .Y(mai_mai_n778_));
  AOI210     m0750(.A0(mai_mai_n100_), .A1(mai_mai_n99_), .B0(mai_mai_n222_), .Y(mai_mai_n779_));
  AN2        m0751(.A(mai_mai_n728_), .B(mai_mai_n720_), .Y(mai_mai_n780_));
  NOi31      m0752(.An(mai_mai_n459_), .B(mai_mai_n736_), .C(mai_mai_n247_), .Y(mai_mai_n781_));
  NO3        m0753(.A(mai_mai_n781_), .B(mai_mai_n780_), .C(mai_mai_n778_), .Y(mai_mai_n782_));
  AO220      m0754(.A0(mai_mai_n385_), .A1(mai_mai_n637_), .B0(mai_mai_n150_), .B1(f), .Y(mai_mai_n783_));
  OAI210     m0755(.A0(mai_mai_n783_), .A1(mai_mai_n388_), .B0(mai_mai_n765_), .Y(mai_mai_n784_));
  NO2        m0756(.A(mai_mai_n372_), .B(mai_mai_n61_), .Y(mai_mai_n785_));
  OAI210     m0757(.A0(mai_mai_n724_), .A1(mai_mai_n785_), .B0(mai_mai_n599_), .Y(mai_mai_n786_));
  AN4        m0758(.A(mai_mai_n786_), .B(mai_mai_n784_), .C(mai_mai_n782_), .D(mai_mai_n775_), .Y(mai_mai_n787_));
  NA4        m0759(.A(mai_mai_n787_), .B(mai_mai_n773_), .C(mai_mai_n759_), .D(mai_mai_n717_), .Y(mai12));
  NO2        m0760(.A(mai_mai_n383_), .B(c), .Y(mai_mai_n789_));
  NO4        m0761(.A(mai_mai_n377_), .B(mai_mai_n215_), .C(mai_mai_n490_), .D(mai_mai_n184_), .Y(mai_mai_n790_));
  NA2        m0762(.A(mai_mai_n790_), .B(mai_mai_n789_), .Y(mai_mai_n791_));
  NO2        m0763(.A(mai_mai_n383_), .B(mai_mai_n98_), .Y(mai_mai_n792_));
  NO2        m0764(.A(mai_mai_n726_), .B(mai_mai_n295_), .Y(mai_mai_n793_));
  NA2        m0765(.A(mai_mai_n793_), .B(mai_mai_n792_), .Y(mai_mai_n794_));
  NA3        m0766(.A(mai_mai_n794_), .B(mai_mai_n791_), .C(mai_mai_n376_), .Y(mai_mai_n795_));
  AOI210     m0767(.A0(mai_mai_n204_), .A1(mai_mai_n286_), .B0(mai_mai_n175_), .Y(mai_mai_n796_));
  BUFFER     m0768(.A(mai_mai_n790_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n327_), .B(mai_mai_n184_), .Y(mai_mai_n798_));
  OAI210     m0770(.A0(mai_mai_n798_), .A1(mai_mai_n797_), .B0(mai_mai_n341_), .Y(mai_mai_n799_));
  NO2        m0771(.A(mai_mai_n546_), .B(mai_mai_n224_), .Y(mai_mai_n800_));
  NO2        m0772(.A(mai_mai_n498_), .B(mai_mai_n719_), .Y(mai_mai_n801_));
  AOI220     m0773(.A0(mai_mai_n801_), .A1(mai_mai_n480_), .B0(mai_mai_n696_), .B1(mai_mai_n800_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n802_), .B(mai_mai_n799_), .Y(mai_mai_n803_));
  NA4        m0775(.A(mai_mai_n378_), .B(mai_mai_n370_), .C(mai_mai_n156_), .D(m), .Y(mai_mai_n804_));
  INV        m0776(.A(mai_mai_n804_), .Y(mai_mai_n805_));
  NO2        m0777(.A(mai_mai_n564_), .B(mai_mai_n74_), .Y(mai_mai_n806_));
  NO4        m0778(.A(mai_mai_n806_), .B(mai_mai_n805_), .C(mai_mai_n803_), .D(mai_mai_n795_), .Y(mai_mai_n807_));
  NO2        m0779(.A(mai_mai_n307_), .B(mai_mai_n306_), .Y(mai_mai_n808_));
  INV        m0780(.A(mai_mai_n495_), .Y(mai_mai_n809_));
  NOi21      m0781(.An(mai_mai_n34_), .B(mai_mai_n555_), .Y(mai_mai_n810_));
  NA2        m0782(.A(mai_mai_n809_), .B(mai_mai_n808_), .Y(mai_mai_n811_));
  INV        m0783(.A(mai_mai_n811_), .Y(mai_mai_n812_));
  NO3        m0784(.A(mai_mai_n698_), .B(mai_mai_n72_), .C(mai_mai_n346_), .Y(mai_mai_n813_));
  NAi21      m0785(.An(mai_mai_n813_), .B(mai_mai_n270_), .Y(mai_mai_n814_));
  NO2        m0786(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n815_));
  NO2        m0787(.A(mai_mai_n422_), .B(mai_mai_n254_), .Y(mai_mai_n816_));
  INV        m0788(.A(mai_mai_n816_), .Y(mai_mai_n817_));
  NO2        m0789(.A(mai_mai_n817_), .B(mai_mai_n124_), .Y(mai_mai_n818_));
  NA2        m0790(.A(mai_mai_n538_), .B(l), .Y(mai_mai_n819_));
  INV        m0791(.A(mai_mai_n304_), .Y(mai_mai_n820_));
  NO4        m0792(.A(mai_mai_n820_), .B(mai_mai_n818_), .C(mai_mai_n814_), .D(mai_mai_n812_), .Y(mai_mai_n821_));
  NA2        m0793(.A(mai_mai_n290_), .B(m), .Y(mai_mai_n822_));
  OAI210     m0794(.A0(mai_mai_n1282_), .A1(mai_mai_n280_), .B0(mai_mai_n822_), .Y(mai_mai_n823_));
  NO2        m0795(.A(mai_mai_n559_), .B(mai_mai_n417_), .Y(mai_mai_n824_));
  NA3        m0796(.A(mai_mai_n289_), .B(j), .C(i), .Y(mai_mai_n825_));
  OAI210     m0797(.A0(mai_mai_n372_), .A1(mai_mai_n260_), .B0(mai_mai_n825_), .Y(mai_mai_n826_));
  OAI220     m0798(.A0(mai_mai_n826_), .A1(mai_mai_n824_), .B0(mai_mai_n576_), .B1(mai_mai_n648_), .Y(mai_mai_n827_));
  NA2        m0799(.A(mai_mai_n514_), .B(mai_mai_n96_), .Y(mai_mai_n828_));
  NA3        m0800(.A(j), .B(mai_mai_n65_), .C(i), .Y(mai_mai_n829_));
  OR2        m0801(.A(mai_mai_n829_), .B(mai_mai_n828_), .Y(mai_mai_n830_));
  NA3        m0802(.A(f), .B(mai_mai_n100_), .C(m), .Y(mai_mai_n831_));
  AOI210     m0803(.A0(mai_mai_n573_), .A1(mai_mai_n831_), .B0(m), .Y(mai_mai_n832_));
  OAI210     m0804(.A0(mai_mai_n832_), .A1(mai_mai_n793_), .B0(mai_mai_n273_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n588_), .B(mai_mai_n748_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n721_), .B(mai_mai_n373_), .Y(mai_mai_n835_));
  NA2        m0807(.A(mai_mai_n192_), .B(h), .Y(mai_mai_n836_));
  NA2        m0808(.A(mai_mai_n836_), .B(mai_mai_n829_), .Y(mai_mai_n837_));
  AOI220     m0809(.A0(mai_mai_n837_), .A1(mai_mai_n221_), .B0(mai_mai_n835_), .B1(mai_mai_n834_), .Y(mai_mai_n838_));
  NA4        m0810(.A(mai_mai_n838_), .B(mai_mai_n833_), .C(mai_mai_n830_), .D(mai_mai_n827_), .Y(mai_mai_n839_));
  NA2        m0811(.A(mai_mai_n563_), .B(mai_mai_n71_), .Y(mai_mai_n840_));
  NA2        m0812(.A(mai_mai_n191_), .B(mai_mai_n321_), .Y(mai_mai_n841_));
  NA2        m0813(.A(mai_mai_n841_), .B(mai_mai_n840_), .Y(mai_mai_n842_));
  OAI210     m0814(.A0(mai_mai_n835_), .A1(mai_mai_n801_), .B0(mai_mai_n457_), .Y(mai_mai_n843_));
  AOI210     m0815(.A0(mai_mai_n357_), .A1(mai_mai_n349_), .B0(mai_mai_n698_), .Y(mai_mai_n844_));
  OAI210     m0816(.A0(mai_mai_n307_), .A1(mai_mai_n306_), .B0(mai_mai_n92_), .Y(mai_mai_n845_));
  AOI210     m0817(.A0(mai_mai_n845_), .A1(mai_mai_n449_), .B0(mai_mai_n844_), .Y(mai_mai_n846_));
  NA2        m0818(.A(mai_mai_n832_), .B(mai_mai_n792_), .Y(mai_mai_n847_));
  NO3        m0819(.A(mai_mai_n1275_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n848_), .B(mai_mai_n533_), .Y(mai_mai_n849_));
  NA4        m0821(.A(mai_mai_n849_), .B(mai_mai_n847_), .C(mai_mai_n846_), .D(mai_mai_n843_), .Y(mai_mai_n850_));
  NO4        m0822(.A(mai_mai_n850_), .B(mai_mai_n842_), .C(mai_mai_n839_), .D(mai_mai_n823_), .Y(mai_mai_n851_));
  NAi21      m0823(.An(mai_mai_n121_), .B(mai_mai_n358_), .Y(mai_mai_n852_));
  NO2        m0824(.A(mai_mai_n229_), .B(mai_mai_n121_), .Y(mai_mai_n853_));
  NA2        m0825(.A(mai_mai_n853_), .B(mai_mai_n418_), .Y(mai_mai_n854_));
  INV        m0826(.A(mai_mai_n412_), .Y(mai_mai_n855_));
  NA2        m0827(.A(mai_mai_n855_), .B(mai_mai_n854_), .Y(mai_mai_n856_));
  NA2        m0828(.A(mai_mai_n201_), .B(mai_mai_n146_), .Y(mai_mai_n857_));
  NO3        m0829(.A(mai_mai_n258_), .B(mai_mai_n378_), .C(mai_mai_n150_), .Y(mai_mai_n858_));
  NOi31      m0830(.An(mai_mai_n857_), .B(mai_mai_n858_), .C(mai_mai_n184_), .Y(mai_mai_n859_));
  OAI220     m0831(.A0(mai_mai_n852_), .A1(mai_mai_n204_), .B0(mai_mai_n825_), .B1(mai_mai_n511_), .Y(mai_mai_n860_));
  NO2        m0832(.A(mai_mai_n560_), .B(mai_mai_n316_), .Y(mai_mai_n861_));
  NA2        m0833(.A(mai_mai_n796_), .B(mai_mai_n789_), .Y(mai_mai_n862_));
  NO3        m0834(.A(mai_mai_n458_), .B(mai_mai_n128_), .C(mai_mai_n183_), .Y(mai_mai_n863_));
  OAI210     m0835(.A0(mai_mai_n863_), .A1(mai_mai_n440_), .B0(mai_mai_n317_), .Y(mai_mai_n864_));
  NA2        m0836(.A(mai_mai_n864_), .B(mai_mai_n862_), .Y(mai_mai_n865_));
  OAI210     m0837(.A0(mai_mai_n796_), .A1(mai_mai_n790_), .B0(mai_mai_n857_), .Y(mai_mai_n866_));
  NA2        m0838(.A(mai_mai_n319_), .B(mai_mai_n317_), .Y(mai_mai_n867_));
  NA3        m0839(.A(mai_mai_n867_), .B(mai_mai_n866_), .C(mai_mai_n230_), .Y(mai_mai_n868_));
  OR4        m0840(.A(mai_mai_n868_), .B(mai_mai_n865_), .C(mai_mai_n861_), .D(mai_mai_n860_), .Y(mai_mai_n869_));
  NO3        m0841(.A(mai_mai_n869_), .B(mai_mai_n859_), .C(mai_mai_n856_), .Y(mai_mai_n870_));
  NA4        m0842(.A(mai_mai_n870_), .B(mai_mai_n851_), .C(mai_mai_n821_), .D(mai_mai_n807_), .Y(mai13));
  NA3        m0843(.A(mai_mai_n214_), .B(b), .C(m), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n416_), .B(f), .Y(mai_mai_n873_));
  NO3        m0845(.A(mai_mai_n873_), .B(mai_mai_n872_), .C(mai_mai_n491_), .Y(mai_mai_n874_));
  NAi32      m0846(.An(d), .Bn(c), .C(e), .Y(mai_mai_n875_));
  NO3        m0847(.A(mai_mai_n875_), .B(mai_mai_n498_), .C(mai_mai_n257_), .Y(mai_mai_n876_));
  NA2        m0848(.A(e), .B(mai_mai_n183_), .Y(mai_mai_n877_));
  NA2        m0849(.A(c), .B(mai_mai_n98_), .Y(mai_mai_n878_));
  NO3        m0850(.A(mai_mai_n878_), .B(mai_mai_n151_), .C(mai_mai_n144_), .Y(mai_mai_n879_));
  NA2        m0851(.A(mai_mai_n416_), .B(c), .Y(mai_mai_n880_));
  NO3        m0852(.A(mai_mai_n494_), .B(mai_mai_n880_), .C(mai_mai_n257_), .Y(mai_mai_n881_));
  OR2        m0853(.A(mai_mai_n879_), .B(mai_mai_n881_), .Y(mai_mai_n882_));
  OR3        m0854(.A(mai_mai_n882_), .B(mai_mai_n876_), .C(mai_mai_n874_), .Y(mai_mai_n883_));
  NAi32      m0855(.An(f), .Bn(e), .C(c), .Y(mai_mai_n884_));
  OR3        m0856(.A(mai_mai_n195_), .B(mai_mai_n151_), .C(mai_mai_n144_), .Y(mai_mai_n885_));
  NO2        m0857(.A(mai_mai_n885_), .B(mai_mai_n884_), .Y(mai_mai_n886_));
  NO2        m0858(.A(mai_mai_n880_), .B(mai_mai_n257_), .Y(mai_mai_n887_));
  NA2        m0859(.A(mai_mai_n535_), .B(mai_mai_n1277_), .Y(mai_mai_n888_));
  NOi21      m0860(.An(mai_mai_n887_), .B(mai_mai_n888_), .Y(mai_mai_n889_));
  NO2        m0861(.A(mai_mai_n652_), .B(mai_mai_n95_), .Y(mai_mai_n890_));
  NOi41      m0862(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n891_));
  NA2        m0863(.A(mai_mai_n891_), .B(mai_mai_n890_), .Y(mai_mai_n892_));
  NO2        m0864(.A(mai_mai_n892_), .B(mai_mai_n884_), .Y(mai_mai_n893_));
  OR3        m0865(.A(e), .B(d), .C(c), .Y(mai_mai_n894_));
  NA3        m0866(.A(k), .B(j), .C(i), .Y(mai_mai_n895_));
  NO3        m0867(.A(mai_mai_n895_), .B(mai_mai_n257_), .C(mai_mai_n73_), .Y(mai_mai_n896_));
  NOi21      m0868(.An(mai_mai_n896_), .B(mai_mai_n894_), .Y(mai_mai_n897_));
  OR4        m0869(.A(mai_mai_n897_), .B(mai_mai_n893_), .C(mai_mai_n889_), .D(mai_mai_n886_), .Y(mai_mai_n898_));
  NA3        m0870(.A(mai_mai_n393_), .B(mai_mai_n282_), .C(mai_mai_n51_), .Y(mai_mai_n899_));
  NO2        m0871(.A(mai_mai_n899_), .B(mai_mai_n888_), .Y(mai_mai_n900_));
  NO2        m0872(.A(mai_mai_n899_), .B(mai_mai_n494_), .Y(mai_mai_n901_));
  NO2        m0873(.A(f), .B(c), .Y(mai_mai_n902_));
  NOi21      m0874(.An(mai_mai_n902_), .B(mai_mai_n377_), .Y(mai_mai_n903_));
  NA2        m0875(.A(mai_mai_n903_), .B(mai_mai_n54_), .Y(mai_mai_n904_));
  OR2        m0876(.A(k), .B(i), .Y(mai_mai_n905_));
  NO3        m0877(.A(mai_mai_n905_), .B(h), .C(l), .Y(mai_mai_n906_));
  NOi31      m0878(.An(mai_mai_n906_), .B(mai_mai_n904_), .C(j), .Y(mai_mai_n907_));
  OR3        m0879(.A(mai_mai_n907_), .B(mai_mai_n901_), .C(mai_mai_n900_), .Y(mai_mai_n908_));
  OR3        m0880(.A(mai_mai_n908_), .B(mai_mai_n898_), .C(mai_mai_n883_), .Y(mai02));
  OR2        m0881(.A(l), .B(k), .Y(mai_mai_n910_));
  OR3        m0882(.A(n), .B(m), .C(i), .Y(mai_mai_n911_));
  NO4        m0883(.A(mai_mai_n911_), .B(h), .C(mai_mai_n910_), .D(mai_mai_n894_), .Y(mai_mai_n912_));
  NOi31      m0884(.An(e), .B(d), .C(c), .Y(mai_mai_n913_));
  AOI210     m0885(.A0(mai_mai_n896_), .A1(mai_mai_n913_), .B0(mai_mai_n876_), .Y(mai_mai_n914_));
  AN3        m0886(.A(m), .B(f), .C(c), .Y(mai_mai_n915_));
  NA2        m0887(.A(mai_mai_n915_), .B(mai_mai_n393_), .Y(mai_mai_n916_));
  OR2        m0888(.A(mai_mai_n895_), .B(mai_mai_n257_), .Y(mai_mai_n917_));
  OR2        m0889(.A(mai_mai_n917_), .B(mai_mai_n916_), .Y(mai_mai_n918_));
  NO2        m0890(.A(mai_mai_n899_), .B(mai_mai_n494_), .Y(mai_mai_n919_));
  NO2        m0891(.A(mai_mai_n919_), .B(mai_mai_n886_), .Y(mai_mai_n920_));
  NA3        m0892(.A(l), .B(k), .C(j), .Y(mai_mai_n921_));
  NA2        m0893(.A(i), .B(h), .Y(mai_mai_n922_));
  NO3        m0894(.A(mai_mai_n922_), .B(mai_mai_n921_), .C(mai_mai_n113_), .Y(mai_mai_n923_));
  NO3        m0895(.A(mai_mai_n122_), .B(mai_mai_n238_), .C(mai_mai_n184_), .Y(mai_mai_n924_));
  AOI210     m0896(.A0(mai_mai_n924_), .A1(mai_mai_n923_), .B0(mai_mai_n889_), .Y(mai_mai_n925_));
  NA3        m0897(.A(c), .B(b), .C(a), .Y(mai_mai_n926_));
  NO3        m0898(.A(mai_mai_n926_), .B(mai_mai_n764_), .C(mai_mai_n183_), .Y(mai_mai_n927_));
  NO2        m0899(.A(mai_mai_n895_), .B(mai_mai_n49_), .Y(mai_mai_n928_));
  AOI210     m0900(.A0(mai_mai_n928_), .A1(mai_mai_n927_), .B0(mai_mai_n900_), .Y(mai_mai_n929_));
  AN4        m0901(.A(mai_mai_n929_), .B(mai_mai_n925_), .C(mai_mai_n920_), .D(mai_mai_n918_), .Y(mai_mai_n930_));
  INV        m0902(.A(mai_mai_n878_), .Y(mai_mai_n931_));
  NA2        m0903(.A(mai_mai_n892_), .B(mai_mai_n885_), .Y(mai_mai_n932_));
  AOI210     m0904(.A0(mai_mai_n932_), .A1(mai_mai_n931_), .B0(mai_mai_n874_), .Y(mai_mai_n933_));
  NAi41      m0905(.An(mai_mai_n912_), .B(mai_mai_n933_), .C(mai_mai_n930_), .D(mai_mai_n914_), .Y(mai03));
  INV        m0906(.A(mai_mai_n845_), .Y(mai_mai_n935_));
  NOi31      m0907(.An(mai_mai_n684_), .B(mai_mai_n722_), .C(mai_mai_n607_), .Y(mai_mai_n936_));
  OAI220     m0908(.A0(mai_mai_n936_), .A1(mai_mai_n588_), .B0(mai_mai_n935_), .B1(mai_mai_n495_), .Y(mai_mai_n937_));
  NOi31      m0909(.An(i), .B(k), .C(j), .Y(mai_mai_n938_));
  NA4        m0910(.A(mai_mai_n938_), .B(mai_mai_n913_), .C(mai_mai_n289_), .D(mai_mai_n282_), .Y(mai_mai_n939_));
  OAI210     m0911(.A0(mai_mai_n698_), .A1(mai_mai_n359_), .B0(mai_mai_n939_), .Y(mai_mai_n940_));
  NOi31      m0912(.An(m), .B(n), .C(f), .Y(mai_mai_n941_));
  NA2        m0913(.A(mai_mai_n425_), .B(l), .Y(mai_mai_n942_));
  NOi31      m0914(.An(mai_mai_n737_), .B(mai_mai_n872_), .C(mai_mai_n942_), .Y(mai_mai_n943_));
  NO3        m0915(.A(mai_mai_n943_), .B(mai_mai_n940_), .C(mai_mai_n844_), .Y(mai_mai_n944_));
  NO2        m0916(.A(mai_mai_n238_), .B(a), .Y(mai_mai_n945_));
  INV        m0917(.A(mai_mai_n876_), .Y(mai_mai_n946_));
  NO2        m0918(.A(mai_mai_n922_), .B(mai_mai_n407_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n70_), .B(m), .Y(mai_mai_n948_));
  AOI210     m0920(.A0(mai_mai_n948_), .A1(mai_mai_n947_), .B0(mai_mai_n906_), .Y(mai_mai_n949_));
  OR2        m0921(.A(mai_mai_n949_), .B(mai_mai_n904_), .Y(mai_mai_n950_));
  NA3        m0922(.A(mai_mai_n950_), .B(mai_mai_n946_), .C(mai_mai_n944_), .Y(mai_mai_n951_));
  NO4        m0923(.A(mai_mai_n951_), .B(mai_mai_n937_), .C(mai_mai_n700_), .D(mai_mai_n479_), .Y(mai_mai_n952_));
  NA2        m0924(.A(c), .B(b), .Y(mai_mai_n953_));
  NO2        m0925(.A(mai_mai_n598_), .B(mai_mai_n953_), .Y(mai_mai_n954_));
  OAI210     m0926(.A0(mai_mai_n736_), .A1(mai_mai_n713_), .B0(mai_mai_n352_), .Y(mai_mai_n955_));
  NA2        m0927(.A(mai_mai_n955_), .B(mai_mai_n954_), .Y(mai_mai_n956_));
  NAi21      m0928(.An(mai_mai_n360_), .B(mai_mai_n954_), .Y(mai_mai_n957_));
  NA2        m0929(.A(mai_mai_n366_), .B(mai_mai_n472_), .Y(mai_mai_n958_));
  OAI210     m0930(.A0(mai_mai_n463_), .A1(mai_mai_n39_), .B0(mai_mai_n945_), .Y(mai_mai_n959_));
  NA3        m0931(.A(mai_mai_n959_), .B(mai_mai_n958_), .C(mai_mai_n957_), .Y(mai_mai_n960_));
  NA2        m0932(.A(mai_mai_n223_), .B(mai_mai_n101_), .Y(mai_mai_n961_));
  OAI210     m0933(.A0(mai_mai_n961_), .A1(mai_mai_n242_), .B0(m), .Y(mai_mai_n962_));
  NAi21      m0934(.An(f), .B(d), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n963_), .B(mai_mai_n926_), .Y(mai_mai_n964_));
  INV        m0936(.A(mai_mai_n964_), .Y(mai_mai_n965_));
  AOI210     m0937(.A0(mai_mai_n962_), .A1(mai_mai_n247_), .B0(mai_mai_n965_), .Y(mai_mai_n966_));
  AOI210     m0938(.A0(mai_mai_n966_), .A1(mai_mai_n96_), .B0(mai_mai_n960_), .Y(mai_mai_n967_));
  INV        m0939(.A(mai_mai_n394_), .Y(mai_mai_n968_));
  NO2        m0940(.A(mai_mai_n157_), .B(mai_mai_n208_), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n969_), .B(m), .Y(mai_mai_n970_));
  NA3        m0942(.A(mai_mai_n779_), .B(mai_mai_n942_), .C(mai_mai_n397_), .Y(mai_mai_n971_));
  OAI210     m0943(.A0(mai_mai_n971_), .A1(mai_mai_n261_), .B0(mai_mai_n395_), .Y(mai_mai_n972_));
  AOI210     m0944(.A0(mai_mai_n972_), .A1(mai_mai_n968_), .B0(mai_mai_n970_), .Y(mai_mai_n973_));
  NA2        m0945(.A(mai_mai_n474_), .B(mai_mai_n348_), .Y(mai_mai_n974_));
  NA2        m0946(.A(mai_mai_n136_), .B(mai_mai_n33_), .Y(mai_mai_n975_));
  AOI210     m0947(.A0(mai_mai_n819_), .A1(mai_mai_n975_), .B0(mai_mai_n184_), .Y(mai_mai_n976_));
  OAI210     m0948(.A0(mai_mai_n976_), .A1(mai_mai_n50_), .B0(mai_mai_n964_), .Y(mai_mai_n977_));
  NO2        m0949(.A(mai_mai_n310_), .B(mai_mai_n309_), .Y(mai_mai_n978_));
  AOI210     m0950(.A0(mai_mai_n969_), .A1(mai_mai_n50_), .B0(mai_mai_n813_), .Y(mai_mai_n979_));
  NAi41      m0951(.An(mai_mai_n978_), .B(mai_mai_n979_), .C(mai_mai_n977_), .D(mai_mai_n974_), .Y(mai_mai_n980_));
  NO2        m0952(.A(mai_mai_n980_), .B(mai_mai_n973_), .Y(mai_mai_n981_));
  NA4        m0953(.A(mai_mai_n981_), .B(mai_mai_n967_), .C(mai_mai_n956_), .D(mai_mai_n952_), .Y(mai00));
  NO2        m0954(.A(mai_mai_n253_), .B(mai_mai_n232_), .Y(mai_mai_n983_));
  NO2        m0955(.A(mai_mai_n983_), .B(mai_mai_n487_), .Y(mai_mai_n984_));
  INV        m0956(.A(mai_mai_n940_), .Y(mai_mai_n985_));
  NO3        m0957(.A(mai_mai_n919_), .B(mai_mai_n813_), .C(mai_mai_n605_), .Y(mai_mai_n986_));
  NA3        m0958(.A(mai_mai_n986_), .B(mai_mai_n985_), .C(mai_mai_n846_), .Y(mai_mai_n987_));
  NA2        m0959(.A(mai_mai_n426_), .B(f), .Y(mai_mai_n988_));
  INV        m0960(.A(mai_mai_n988_), .Y(mai_mai_n989_));
  NO4        m0961(.A(mai_mai_n989_), .B(mai_mai_n987_), .C(mai_mai_n984_), .D(mai_mai_n898_), .Y(mai_mai_n990_));
  NA3        m0962(.A(mai_mai_n143_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n991_));
  NA3        m0963(.A(d), .B(mai_mai_n51_), .C(b), .Y(mai_mai_n992_));
  NOi31      m0964(.An(n), .B(m), .C(i), .Y(mai_mai_n993_));
  NA3        m0965(.A(mai_mai_n993_), .B(mai_mai_n551_), .C(mai_mai_n50_), .Y(mai_mai_n994_));
  OAI210     m0966(.A0(mai_mai_n992_), .A1(mai_mai_n991_), .B0(mai_mai_n994_), .Y(mai_mai_n995_));
  NO3        m0967(.A(mai_mai_n995_), .B(mai_mai_n978_), .C(mai_mai_n781_), .Y(mai_mai_n996_));
  NO3        m0968(.A(mai_mai_n1278_), .B(mai_mai_n296_), .C(mai_mai_n953_), .Y(mai_mai_n997_));
  OR2        m0969(.A(mai_mai_n323_), .B(mai_mai_n115_), .Y(mai_mai_n998_));
  NO2        m0970(.A(h), .B(m), .Y(mai_mai_n999_));
  NO2        m0971(.A(mai_mai_n74_), .B(mai_mai_n73_), .Y(mai_mai_n1000_));
  NA2        m0972(.A(mai_mai_n1000_), .B(mai_mai_n449_), .Y(mai_mai_n1001_));
  NA2        m0973(.A(mai_mai_n152_), .B(mai_mai_n127_), .Y(mai_mai_n1002_));
  NA3        m0974(.A(mai_mai_n1002_), .B(mai_mai_n1001_), .C(mai_mai_n998_), .Y(mai_mai_n1003_));
  NO2        m0975(.A(mai_mai_n1003_), .B(mai_mai_n997_), .Y(mai_mai_n1004_));
  INV        m0976(.A(mai_mai_n132_), .Y(mai_mai_n1005_));
  NA3        m0977(.A(mai_mai_n154_), .B(mai_mai_n95_), .C(m), .Y(mai_mai_n1006_));
  NOi21      m0978(.An(mai_mai_n742_), .B(mai_mai_n1006_), .Y(mai_mai_n1007_));
  NAi21      m0979(.An(mai_mai_n159_), .B(mai_mai_n733_), .Y(mai_mai_n1008_));
  NAi21      m0980(.An(mai_mai_n1007_), .B(mai_mai_n1008_), .Y(mai_mai_n1009_));
  NO2        m0981(.A(mai_mai_n231_), .B(mai_mai_n63_), .Y(mai_mai_n1010_));
  NO3        m0982(.A(mai_mai_n365_), .B(mai_mai_n710_), .C(n), .Y(mai_mai_n1011_));
  AOI210     m0983(.A0(mai_mai_n1011_), .A1(mai_mai_n1010_), .B0(mai_mai_n912_), .Y(mai_mai_n1012_));
  NAi21      m0984(.An(mai_mai_n881_), .B(mai_mai_n1012_), .Y(mai_mai_n1013_));
  NO3        m0985(.A(mai_mai_n1013_), .B(mai_mai_n1009_), .C(mai_mai_n1005_), .Y(mai_mai_n1014_));
  AN3        m0986(.A(mai_mai_n1014_), .B(mai_mai_n1004_), .C(mai_mai_n996_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(mai_mai_n449_), .B(mai_mai_n84_), .Y(mai_mai_n1016_));
  NA2        m0988(.A(mai_mai_n475_), .B(mai_mai_n1016_), .Y(mai_mai_n1017_));
  OAI210     m0989(.A0(mai_mai_n392_), .A1(mai_mai_n102_), .B0(mai_mai_n738_), .Y(mai_mai_n1018_));
  AOI220     m0990(.A0(mai_mai_n1018_), .A1(mai_mai_n971_), .B0(mai_mai_n474_), .B1(mai_mai_n348_), .Y(mai_mai_n1019_));
  OR2        m0991(.A(mai_mai_n229_), .B(mai_mai_n193_), .Y(mai_mai_n1020_));
  NA2        m0992(.A(n), .B(e), .Y(mai_mai_n1021_));
  NO2        m0993(.A(mai_mai_n1021_), .B(mai_mai_n125_), .Y(mai_mai_n1022_));
  NA2        m0994(.A(mai_mai_n297_), .B(mai_mai_n381_), .Y(mai_mai_n1023_));
  NA3        m0995(.A(mai_mai_n1023_), .B(mai_mai_n1020_), .C(mai_mai_n1019_), .Y(mai_mai_n1024_));
  AOI210     m0996(.A0(mai_mai_n1022_), .A1(mai_mai_n727_), .B0(mai_mai_n699_), .Y(mai_mai_n1025_));
  AOI220     m0997(.A0(mai_mai_n810_), .A1(d), .B0(mai_mai_n551_), .B1(mai_mai_n210_), .Y(mai_mai_n1026_));
  NO2        m0998(.A(i), .B(h), .Y(mai_mai_n1027_));
  NO2        m0999(.A(mai_mai_n878_), .B(mai_mai_n617_), .Y(mai_mai_n1028_));
  NO2        m1000(.A(mai_mai_n910_), .B(mai_mai_n113_), .Y(mai_mai_n1029_));
  AN2        m1001(.A(mai_mai_n1029_), .B(mai_mai_n924_), .Y(mai_mai_n1030_));
  OAI210     m1002(.A0(mai_mai_n1030_), .A1(mai_mai_n1028_), .B0(mai_mai_n1027_), .Y(mai_mai_n1031_));
  NA4        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1026_), .C(mai_mai_n1025_), .D(mai_mai_n738_), .Y(mai_mai_n1032_));
  NO4        m1004(.A(mai_mai_n1032_), .B(mai_mai_n1024_), .C(mai_mai_n249_), .D(mai_mai_n1017_), .Y(mai_mai_n1033_));
  NA2        m1005(.A(mai_mai_n714_), .B(mai_mai_n647_), .Y(mai_mai_n1034_));
  NA4        m1006(.A(mai_mai_n1034_), .B(mai_mai_n1033_), .C(mai_mai_n1015_), .D(mai_mai_n990_), .Y(mai01));
  AN2        m1007(.A(mai_mai_n864_), .B(mai_mai_n862_), .Y(mai_mai_n1036_));
  NO2        m1008(.A(mai_mai_n680_), .B(mai_mai_n237_), .Y(mai_mai_n1037_));
  INV        m1009(.A(mai_mai_n332_), .Y(mai_mai_n1038_));
  NA3        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1037_), .C(mai_mai_n1036_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n777_), .B(mai_mai_n281_), .Y(mai_mai_n1040_));
  NA2        m1012(.A(mai_mai_n603_), .B(mai_mai_n79_), .Y(mai_mai_n1041_));
  NO2        m1013(.A(mai_mai_n1041_), .B(mai_mai_n1272_), .Y(mai_mai_n1042_));
  NA2        m1014(.A(mai_mai_n1042_), .B(mai_mai_n542_), .Y(mai_mai_n1043_));
  INV        m1015(.A(mai_mai_n100_), .Y(mai_mai_n1044_));
  NAi21      m1016(.An(mai_mai_n139_), .B(mai_mai_n1043_), .Y(mai_mai_n1045_));
  NO3        m1017(.A(mai_mai_n670_), .B(mai_mai_n575_), .C(mai_mai_n428_), .Y(mai_mai_n1046_));
  NA4        m1018(.A(mai_mai_n603_), .B(mai_mai_n79_), .C(mai_mai_n45_), .D(mai_mai_n183_), .Y(mai_mai_n1047_));
  OA220      m1019(.A0(mai_mai_n1047_), .A1(mai_mai_n569_), .B0(mai_mai_n169_), .B1(mai_mai_n167_), .Y(mai_mai_n1048_));
  NA3        m1020(.A(mai_mai_n1048_), .B(mai_mai_n1046_), .C(mai_mai_n118_), .Y(mai_mai_n1049_));
  NO4        m1021(.A(mai_mai_n1049_), .B(mai_mai_n1045_), .C(mai_mai_n1040_), .D(mai_mai_n1039_), .Y(mai_mai_n1050_));
  NA2        m1022(.A(mai_mai_n452_), .B(mai_mai_n334_), .Y(mai_mai_n1051_));
  BUFFER     m1023(.A(mai_mai_n476_), .Y(mai_mai_n1052_));
  NA2        m1024(.A(mai_mai_n1052_), .B(mai_mai_n1051_), .Y(mai_mai_n1053_));
  AOI210     m1025(.A0(mai_mai_n178_), .A1(mai_mai_n72_), .B0(mai_mai_n183_), .Y(mai_mai_n1054_));
  OAI210     m1026(.A0(mai_mai_n687_), .A1(mai_mai_n366_), .B0(mai_mai_n1054_), .Y(mai_mai_n1055_));
  AN3        m1027(.A(m), .B(l), .C(k), .Y(mai_mai_n1056_));
  OAI210     m1028(.A0(mai_mai_n299_), .A1(mai_mai_n34_), .B0(mai_mai_n1056_), .Y(mai_mai_n1057_));
  NA2        m1029(.A(mai_mai_n177_), .B(mai_mai_n34_), .Y(mai_mai_n1058_));
  AO210      m1030(.A0(mai_mai_n1058_), .A1(mai_mai_n1057_), .B0(mai_mai_n280_), .Y(mai_mai_n1059_));
  NA3        m1031(.A(mai_mai_n1059_), .B(mai_mai_n1055_), .C(mai_mai_n1053_), .Y(mai_mai_n1060_));
  NO2        m1032(.A(mai_mai_n1044_), .B(mai_mai_n502_), .Y(mai_mai_n1061_));
  NA2        m1033(.A(mai_mai_n236_), .B(mai_mai_n169_), .Y(mai_mai_n1062_));
  NA2        m1034(.A(mai_mai_n1062_), .B(mai_mai_n566_), .Y(mai_mai_n1063_));
  NO3        m1035(.A(mai_mai_n698_), .B(mai_mai_n178_), .C(mai_mai_n346_), .Y(mai_mai_n1064_));
  NO2        m1036(.A(mai_mai_n1064_), .B(mai_mai_n813_), .Y(mai_mai_n1065_));
  OAI210     m1037(.A0(mai_mai_n1042_), .A1(mai_mai_n275_), .B0(mai_mai_n576_), .Y(mai_mai_n1066_));
  NA4        m1038(.A(mai_mai_n1066_), .B(mai_mai_n1065_), .C(mai_mai_n1063_), .D(mai_mai_n672_), .Y(mai_mai_n1067_));
  NO3        m1039(.A(mai_mai_n1067_), .B(mai_mai_n1061_), .C(mai_mai_n1060_), .Y(mai_mai_n1068_));
  NA3        m1040(.A(mai_mai_n512_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1069_));
  NO2        m1041(.A(mai_mai_n1069_), .B(mai_mai_n178_), .Y(mai_mai_n1070_));
  AOI210     m1042(.A0(mai_mai_n423_), .A1(mai_mai_n53_), .B0(mai_mai_n1070_), .Y(mai_mai_n1071_));
  OR3        m1043(.A(mai_mai_n1041_), .B(mai_mai_n513_), .C(mai_mai_n1272_), .Y(mai_mai_n1072_));
  NO2        m1044(.A(mai_mai_n1047_), .B(mai_mai_n828_), .Y(mai_mai_n1073_));
  NO2        m1045(.A(mai_mai_n1073_), .B(mai_mai_n995_), .Y(mai_mai_n1074_));
  NA4        m1046(.A(mai_mai_n1074_), .B(mai_mai_n1072_), .C(mai_mai_n1071_), .D(mai_mai_n646_), .Y(mai_mai_n1075_));
  NO2        m1047(.A(m), .B(mai_mai_n203_), .Y(mai_mai_n1076_));
  INV        m1048(.A(mai_mai_n571_), .Y(mai_mai_n1077_));
  NO2        m1049(.A(mai_mai_n308_), .B(mai_mai_n62_), .Y(mai_mai_n1078_));
  INV        m1050(.A(mai_mai_n1078_), .Y(mai_mai_n1079_));
  NA2        m1051(.A(mai_mai_n1079_), .B(mai_mai_n325_), .Y(mai_mai_n1080_));
  NO3        m1052(.A(mai_mai_n1080_), .B(mai_mai_n1077_), .C(mai_mai_n1075_), .Y(mai_mai_n1081_));
  NO2        m1053(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1082_));
  AN2        m1054(.A(mai_mai_n1082_), .B(mai_mai_n530_), .Y(mai_mai_n1083_));
  NA2        m1055(.A(mai_mai_n1083_), .B(mai_mai_n288_), .Y(mai_mai_n1084_));
  INV        m1056(.A(mai_mai_n115_), .Y(mai_mai_n1085_));
  NO3        m1057(.A(mai_mai_n922_), .B(mai_mai_n151_), .C(mai_mai_n70_), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n1085_), .Y(mai_mai_n1087_));
  NA2        m1059(.A(mai_mai_n1087_), .B(mai_mai_n1084_), .Y(mai_mai_n1088_));
  NO2        m1060(.A(mai_mai_n522_), .B(mai_mai_n521_), .Y(mai_mai_n1089_));
  NO4        m1061(.A(mai_mai_n922_), .B(mai_mai_n1089_), .C(mai_mai_n149_), .D(mai_mai_n70_), .Y(mai_mai_n1090_));
  NO3        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1088_), .C(mai_mai_n545_), .Y(mai_mai_n1091_));
  NA4        m1063(.A(mai_mai_n1091_), .B(mai_mai_n1081_), .C(mai_mai_n1068_), .D(mai_mai_n1050_), .Y(mai06));
  NO2        m1064(.A(mai_mai_n347_), .B(mai_mai_n473_), .Y(mai_mai_n1093_));
  OAI210     m1065(.A0(mai_mai_n96_), .A1(mai_mai_n225_), .B0(mai_mai_n1093_), .Y(mai_mai_n1094_));
  NO2        m1066(.A(mai_mai_n195_), .B(mai_mai_n86_), .Y(mai_mai_n1095_));
  OAI210     m1067(.A0(mai_mai_n1095_), .A1(mai_mai_n1086_), .B0(mai_mai_n321_), .Y(mai_mai_n1096_));
  NO3        m1068(.A(mai_mai_n508_), .B(mai_mai_n685_), .C(mai_mai_n510_), .Y(mai_mai_n1097_));
  OR2        m1069(.A(mai_mai_n1097_), .B(mai_mai_n755_), .Y(mai_mai_n1098_));
  NA3        m1070(.A(mai_mai_n1098_), .B(mai_mai_n1096_), .C(mai_mai_n1094_), .Y(mai_mai_n1099_));
  NO3        m1071(.A(mai_mai_n1099_), .B(mai_mai_n1077_), .C(mai_mai_n219_), .Y(mai_mai_n1100_));
  AOI210     m1072(.A0(i), .A1(mai_mai_n468_), .B0(mai_mai_n1076_), .Y(mai_mai_n1101_));
  INV        m1073(.A(mai_mai_n1083_), .Y(mai_mai_n1102_));
  AOI210     m1074(.A0(mai_mai_n1102_), .A1(mai_mai_n1101_), .B0(mai_mai_n286_), .Y(mai_mai_n1103_));
  INV        m1075(.A(mai_mai_n574_), .Y(mai_mai_n1104_));
  NA2        m1076(.A(mai_mai_n1104_), .B(mai_mai_n549_), .Y(mai_mai_n1105_));
  NO2        m1077(.A(mai_mai_n430_), .B(mai_mai_n146_), .Y(mai_mai_n1106_));
  NOi21      m1078(.An(mai_mai_n117_), .B(mai_mai_n45_), .Y(mai_mai_n1107_));
  OAI210     m1079(.A0(mai_mai_n389_), .A1(mai_mai_n213_), .B0(mai_mai_n771_), .Y(mai_mai_n1108_));
  NO3        m1080(.A(mai_mai_n1108_), .B(mai_mai_n1107_), .C(mai_mai_n1106_), .Y(mai_mai_n1109_));
  NA2        m1081(.A(mai_mai_n1109_), .B(mai_mai_n1105_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(mai_mai_n638_), .B(mai_mai_n306_), .Y(mai_mai_n1111_));
  NOi21      m1083(.An(mai_mai_n1111_), .B(mai_mai_n49_), .Y(mai_mai_n1112_));
  NO3        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1110_), .C(mai_mai_n1103_), .Y(mai_mai_n1113_));
  NO2        m1085(.A(mai_mai_n679_), .B(mai_mai_n233_), .Y(mai_mai_n1114_));
  OAI220     m1086(.A0(mai_mai_n624_), .A1(mai_mai_n47_), .B0(mai_mai_n195_), .B1(mai_mai_n524_), .Y(mai_mai_n1115_));
  OAI210     m1087(.A0(mai_mai_n233_), .A1(c), .B0(mai_mai_n548_), .Y(mai_mai_n1116_));
  AOI220     m1088(.A0(mai_mai_n1116_), .A1(mai_mai_n1115_), .B0(mai_mai_n1114_), .B1(mai_mai_n225_), .Y(mai_mai_n1117_));
  OAI220     m1089(.A0(mai_mai_n595_), .A1(mai_mai_n213_), .B0(mai_mai_n427_), .B1(mai_mai_n430_), .Y(mai_mai_n1118_));
  INV        m1090(.A(mai_mai_n507_), .Y(mai_mai_n1119_));
  NOi21      m1091(.An(mai_mai_n1119_), .B(mai_mai_n569_), .Y(mai_mai_n1120_));
  NO2        m1092(.A(mai_mai_n1120_), .B(mai_mai_n1118_), .Y(mai_mai_n1121_));
  NAi31      m1093(.An(mai_mai_n638_), .B(mai_mai_n369_), .C(mai_mai_n177_), .Y(mai_mai_n1122_));
  NA4        m1094(.A(mai_mai_n1122_), .B(mai_mai_n1121_), .C(mai_mai_n1117_), .D(mai_mai_n1026_), .Y(mai_mai_n1123_));
  NOi31      m1095(.An(mai_mai_n1097_), .B(mai_mai_n391_), .C(mai_mai_n333_), .Y(mai_mai_n1124_));
  OR3        m1096(.A(mai_mai_n1124_), .B(mai_mai_n669_), .C(mai_mai_n455_), .Y(mai_mai_n1125_));
  AOI210     m1097(.A0(mai_mai_n485_), .A1(mai_mai_n381_), .B0(mai_mai_n311_), .Y(mai_mai_n1126_));
  NA2        m1098(.A(mai_mai_n1126_), .B(mai_mai_n1125_), .Y(mai_mai_n1127_));
  AN2        m1099(.A(mai_mai_n790_), .B(mai_mai_n789_), .Y(mai_mai_n1128_));
  NO2        m1100(.A(mai_mai_n1128_), .B(mai_mai_n746_), .Y(mai_mai_n1129_));
  INV        m1101(.A(mai_mai_n1129_), .Y(mai_mai_n1130_));
  NAi21      m1102(.An(j), .B(i), .Y(mai_mai_n1131_));
  NO4        m1103(.A(mai_mai_n1089_), .B(mai_mai_n1131_), .C(mai_mai_n377_), .D(mai_mai_n206_), .Y(mai_mai_n1132_));
  NO4        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1130_), .C(mai_mai_n1127_), .D(mai_mai_n1123_), .Y(mai_mai_n1133_));
  NA4        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1113_), .C(mai_mai_n1100_), .D(mai_mai_n1091_), .Y(mai07));
  NOi21      m1106(.An(j), .B(k), .Y(mai_mai_n1135_));
  NA4        m1107(.A(mai_mai_n154_), .B(mai_mai_n91_), .C(mai_mai_n1135_), .D(f), .Y(mai_mai_n1136_));
  NAi21      m1108(.An(f), .B(c), .Y(mai_mai_n1137_));
  OR2        m1109(.A(e), .B(d), .Y(mai_mai_n1138_));
  NO2        m1110(.A(mai_mai_n534_), .B(mai_mai_n272_), .Y(mai_mai_n1139_));
  NA3        m1111(.A(mai_mai_n1139_), .B(mai_mai_n1277_), .C(mai_mai_n154_), .Y(mai_mai_n1140_));
  NOi31      m1112(.An(n), .B(m), .C(b), .Y(mai_mai_n1141_));
  NO3        m1113(.A(mai_mai_n113_), .B(mai_mai_n382_), .C(h), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n1140_), .B(mai_mai_n1136_), .Y(mai_mai_n1143_));
  NOi31      m1115(.An(i), .B(m), .C(h), .Y(mai_mai_n1144_));
  NA2        m1116(.A(mai_mai_n70_), .B(mai_mai_n45_), .Y(mai_mai_n1145_));
  NO2        m1117(.A(mai_mai_n884_), .B(mai_mai_n377_), .Y(mai_mai_n1146_));
  NA3        m1118(.A(mai_mai_n1146_), .B(mai_mai_n1145_), .C(mai_mai_n184_), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n895_), .B(mai_mai_n257_), .Y(mai_mai_n1148_));
  NA2        m1120(.A(mai_mai_n456_), .B(mai_mai_n65_), .Y(mai_mai_n1149_));
  NA2        m1121(.A(mai_mai_n1149_), .B(mai_mai_n1147_), .Y(mai_mai_n1150_));
  NO2        m1122(.A(mai_mai_n1150_), .B(mai_mai_n1143_), .Y(mai_mai_n1151_));
  NO3        m1123(.A(e), .B(d), .C(c), .Y(mai_mai_n1152_));
  NA2        m1124(.A(mai_mai_n1271_), .B(mai_mai_n1152_), .Y(mai_mai_n1153_));
  NO2        m1125(.A(mai_mai_n1153_), .B(mai_mai_n184_), .Y(mai_mai_n1154_));
  NO2        m1126(.A(l), .B(k), .Y(mai_mai_n1155_));
  NOi41      m1127(.An(mai_mai_n461_), .B(mai_mai_n1155_), .C(mai_mai_n402_), .D(mai_mai_n377_), .Y(mai_mai_n1156_));
  NO2        m1128(.A(mai_mai_n1156_), .B(mai_mai_n1154_), .Y(mai_mai_n1157_));
  NO2        m1129(.A(mai_mai_n905_), .B(l), .Y(mai_mai_n1158_));
  NO2        m1130(.A(m), .B(c), .Y(mai_mai_n1159_));
  NA3        m1131(.A(mai_mai_n1159_), .B(mai_mai_n122_), .C(mai_mai_n160_), .Y(mai_mai_n1160_));
  NO2        m1132(.A(mai_mai_n1160_), .B(mai_mai_n1158_), .Y(mai_mai_n1161_));
  NA2        m1133(.A(mai_mai_n1161_), .B(mai_mai_n154_), .Y(mai_mai_n1162_));
  NO2        m1134(.A(mai_mai_n383_), .B(a), .Y(mai_mai_n1163_));
  NA3        m1135(.A(mai_mai_n1163_), .B(mai_mai_n1274_), .C(mai_mai_n96_), .Y(mai_mai_n1164_));
  NA2        m1136(.A(mai_mai_n963_), .B(h), .Y(mai_mai_n1165_));
  NA2        m1137(.A(mai_mai_n119_), .B(mai_mai_n191_), .Y(mai_mai_n1166_));
  NO2        m1138(.A(mai_mai_n1166_), .B(mai_mai_n1165_), .Y(mai_mai_n1167_));
  NOi31      m1139(.An(m), .B(n), .C(b), .Y(mai_mai_n1168_));
  INV        m1140(.A(mai_mai_n1167_), .Y(mai_mai_n1169_));
  NA2        m1141(.A(mai_mai_n915_), .B(mai_mai_n393_), .Y(mai_mai_n1170_));
  NO4        m1142(.A(mai_mai_n1170_), .B(mai_mai_n890_), .C(mai_mai_n377_), .D(mai_mai_n45_), .Y(mai_mai_n1171_));
  OAI210     m1143(.A0(mai_mai_n157_), .A1(mai_mai_n441_), .B0(mai_mai_n891_), .Y(mai_mai_n1172_));
  INV        m1144(.A(mai_mai_n1172_), .Y(mai_mai_n1173_));
  NO2        m1145(.A(mai_mai_n1173_), .B(mai_mai_n1171_), .Y(mai_mai_n1174_));
  AN4        m1146(.A(mai_mai_n1174_), .B(mai_mai_n1169_), .C(mai_mai_n1164_), .D(mai_mai_n1162_), .Y(mai_mai_n1175_));
  NA2        m1147(.A(mai_mai_n1141_), .B(mai_mai_n318_), .Y(mai_mai_n1176_));
  NO2        m1148(.A(mai_mai_n161_), .B(b), .Y(mai_mai_n1177_));
  AOI220     m1149(.A0(mai_mai_n993_), .A1(mai_mai_n1177_), .B0(mai_mai_n923_), .B1(mai_mai_n1170_), .Y(mai_mai_n1178_));
  INV        m1150(.A(mai_mai_n1178_), .Y(mai_mai_n1179_));
  NO4        m1151(.A(mai_mai_n113_), .B(m), .C(f), .D(e), .Y(mai_mai_n1180_));
  NA2        m1152(.A(mai_mai_n246_), .B(h), .Y(mai_mai_n1181_));
  OR2        m1153(.A(e), .B(a), .Y(mai_mai_n1182_));
  NO2        m1154(.A(mai_mai_n1138_), .B(mai_mai_n1137_), .Y(mai_mai_n1183_));
  AOI210     m1155(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1183_), .Y(mai_mai_n1184_));
  NO2        m1156(.A(mai_mai_n1184_), .B(mai_mai_n911_), .Y(mai_mai_n1185_));
  NA2        m1157(.A(mai_mai_n1144_), .B(mai_mai_n1155_), .Y(mai_mai_n1186_));
  INV        m1158(.A(mai_mai_n1186_), .Y(mai_mai_n1187_));
  NA2        m1159(.A(mai_mai_n941_), .B(mai_mai_n346_), .Y(mai_mai_n1188_));
  NO3        m1160(.A(mai_mai_n1187_), .B(mai_mai_n1185_), .C(mai_mai_n1179_), .Y(mai_mai_n1189_));
  NA4        m1161(.A(mai_mai_n1189_), .B(mai_mai_n1175_), .C(mai_mai_n1157_), .D(mai_mai_n1151_), .Y(mai_mai_n1190_));
  NO2        m1162(.A(mai_mai_n329_), .B(j), .Y(mai_mai_n1191_));
  NA3        m1163(.A(m), .B(mai_mai_n1191_), .C(mai_mai_n136_), .Y(mai_mai_n1192_));
  OR2        m1164(.A(n), .B(i), .Y(mai_mai_n1193_));
  OAI210     m1165(.A0(mai_mai_n1193_), .A1(mai_mai_n902_), .B0(mai_mai_n49_), .Y(mai_mai_n1194_));
  AOI220     m1166(.A0(mai_mai_n1194_), .A1(mai_mai_n999_), .B0(mai_mai_n703_), .B1(mai_mai_n168_), .Y(mai_mai_n1195_));
  NO2        m1167(.A(mai_mai_n195_), .B(k), .Y(mai_mai_n1196_));
  NO2        m1168(.A(mai_mai_n911_), .B(h), .Y(mai_mai_n1197_));
  NA3        m1169(.A(mai_mai_n1197_), .B(d), .C(mai_mai_n877_), .Y(mai_mai_n1198_));
  NO2        m1170(.A(mai_mai_n1198_), .B(c), .Y(mai_mai_n1199_));
  NOi21      m1171(.An(d), .B(f), .Y(mai_mai_n1200_));
  NO2        m1172(.A(mai_mai_n1138_), .B(f), .Y(mai_mai_n1201_));
  INV        m1173(.A(mai_mai_n1199_), .Y(mai_mai_n1202_));
  NA3        m1174(.A(mai_mai_n1202_), .B(mai_mai_n1195_), .C(mai_mai_n1192_), .Y(mai_mai_n1203_));
  NO3        m1175(.A(mai_mai_n915_), .B(mai_mai_n902_), .C(mai_mai_n40_), .Y(mai_mai_n1204_));
  NA2        m1176(.A(mai_mai_n1204_), .B(mai_mai_n1148_), .Y(mai_mai_n1205_));
  OAI210     m1177(.A0(mai_mai_n1180_), .A1(mai_mai_n1141_), .B0(mai_mai_n753_), .Y(mai_mai_n1206_));
  NO2        m1178(.A(mai_mai_n875_), .B(mai_mai_n113_), .Y(mai_mai_n1207_));
  NA2        m1179(.A(mai_mai_n1207_), .B(mai_mai_n529_), .Y(mai_mai_n1208_));
  NA3        m1180(.A(mai_mai_n1208_), .B(mai_mai_n1206_), .C(mai_mai_n1205_), .Y(mai_mai_n1209_));
  NA2        m1181(.A(mai_mai_n1159_), .B(mai_mai_n1200_), .Y(mai_mai_n1210_));
  NO2        m1182(.A(mai_mai_n1210_), .B(m), .Y(mai_mai_n1211_));
  NO2        m1183(.A(mai_mai_n129_), .B(mai_mai_n156_), .Y(mai_mai_n1212_));
  OAI210     m1184(.A0(mai_mai_n1212_), .A1(mai_mai_n93_), .B0(mai_mai_n1168_), .Y(mai_mai_n1213_));
  INV        m1185(.A(mai_mai_n1213_), .Y(mai_mai_n1214_));
  NO3        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1211_), .C(mai_mai_n1209_), .Y(mai_mai_n1215_));
  NO2        m1187(.A(mai_mai_n1137_), .B(e), .Y(mai_mai_n1216_));
  NA2        m1188(.A(mai_mai_n1216_), .B(mai_mai_n344_), .Y(mai_mai_n1217_));
  OAI210     m1189(.A0(mai_mai_n1201_), .A1(mai_mai_n948_), .B0(mai_mai_n538_), .Y(mai_mai_n1218_));
  OR3        m1190(.A(mai_mai_n1196_), .B(mai_mai_n1027_), .C(mai_mai_n113_), .Y(mai_mai_n1219_));
  OAI220     m1191(.A0(mai_mai_n1219_), .A1(mai_mai_n1217_), .B0(mai_mai_n1218_), .B1(mai_mai_n379_), .Y(mai_mai_n1220_));
  INV        m1192(.A(mai_mai_n1220_), .Y(mai_mai_n1221_));
  NO2        m1193(.A(mai_mai_n156_), .B(c), .Y(mai_mai_n1222_));
  OAI210     m1194(.A0(mai_mai_n1222_), .A1(mai_mai_n1216_), .B0(mai_mai_n154_), .Y(mai_mai_n1223_));
  AOI220     m1195(.A0(mai_mai_n1223_), .A1(mai_mai_n904_), .B0(mai_mai_n447_), .B1(mai_mai_n306_), .Y(mai_mai_n1224_));
  NO2        m1196(.A(mai_mai_n1182_), .B(f), .Y(mai_mai_n1225_));
  NA2        m1197(.A(mai_mai_n948_), .B(a), .Y(mai_mai_n1226_));
  NO2        m1198(.A(mai_mai_n1226_), .B(mai_mai_n60_), .Y(mai_mai_n1227_));
  NA2        m1199(.A(mai_mai_n1225_), .B(mai_mai_n1145_), .Y(mai_mai_n1228_));
  OAI220     m1200(.A0(mai_mai_n1228_), .A1(mai_mai_n49_), .B0(mai_mai_n1273_), .B1(mai_mai_n149_), .Y(mai_mai_n1229_));
  NA4        m1201(.A(mai_mai_n924_), .B(mai_mai_n921_), .C(mai_mai_n191_), .D(i), .Y(mai_mai_n1230_));
  NA2        m1202(.A(mai_mai_n1142_), .B(mai_mai_n157_), .Y(mai_mai_n1231_));
  NO2        m1203(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1232_));
  OAI210     m1204(.A0(mai_mai_n1182_), .A1(mai_mai_n735_), .B0(mai_mai_n406_), .Y(mai_mai_n1233_));
  OAI210     m1205(.A0(mai_mai_n1233_), .A1(mai_mai_n927_), .B0(mai_mai_n1232_), .Y(mai_mai_n1234_));
  NO2        m1206(.A(mai_mai_n215_), .B(m), .Y(mai_mai_n1235_));
  NO2        m1207(.A(m), .B(i), .Y(mai_mai_n1236_));
  NA2        m1208(.A(mai_mai_n903_), .B(mai_mai_n1235_), .Y(mai_mai_n1237_));
  NA4        m1209(.A(mai_mai_n1237_), .B(mai_mai_n1234_), .C(mai_mai_n1231_), .D(mai_mai_n1230_), .Y(mai_mai_n1238_));
  NO4        m1210(.A(mai_mai_n1238_), .B(mai_mai_n1229_), .C(mai_mai_n1227_), .D(mai_mai_n1224_), .Y(mai_mai_n1239_));
  NA3        m1211(.A(mai_mai_n1239_), .B(mai_mai_n1221_), .C(mai_mai_n1215_), .Y(mai_mai_n1240_));
  NA3        m1212(.A(mai_mai_n815_), .B(mai_mai_n119_), .C(mai_mai_n46_), .Y(mai_mai_n1241_));
  AOI210     m1213(.A0(mai_mai_n127_), .A1(c), .B0(mai_mai_n1241_), .Y(mai_mai_n1242_));
  INV        m1214(.A(mai_mai_n158_), .Y(mai_mai_n1243_));
  NA2        m1215(.A(mai_mai_n1243_), .B(mai_mai_n1197_), .Y(mai_mai_n1244_));
  AO210      m1216(.A0(mai_mai_n114_), .A1(l), .B0(mai_mai_n1176_), .Y(mai_mai_n1245_));
  NA2        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1244_), .Y(mai_mai_n1246_));
  NO2        m1218(.A(mai_mai_n1246_), .B(mai_mai_n1242_), .Y(mai_mai_n1247_));
  NO4        m1219(.A(mai_mai_n195_), .B(mai_mai_n159_), .C(mai_mai_n220_), .D(k), .Y(mai_mai_n1248_));
  NOi21      m1220(.An(mai_mai_n1142_), .B(e), .Y(mai_mai_n1249_));
  NO2        m1221(.A(mai_mai_n1249_), .B(mai_mai_n1248_), .Y(mai_mai_n1250_));
  AN2        m1222(.A(mai_mai_n924_), .B(mai_mai_n910_), .Y(mai_mai_n1251_));
  AOI220     m1223(.A0(mai_mai_n1236_), .A1(mai_mai_n547_), .B0(mai_mai_n1277_), .B1(mai_mai_n137_), .Y(mai_mai_n1252_));
  NOi31      m1224(.An(mai_mai_n30_), .B(mai_mai_n1252_), .C(n), .Y(mai_mai_n1253_));
  AOI210     m1225(.A0(mai_mai_n1251_), .A1(mai_mai_n993_), .B0(mai_mai_n1253_), .Y(mai_mai_n1254_));
  NA2        m1226(.A(mai_mai_n54_), .B(a), .Y(mai_mai_n1255_));
  NO2        m1227(.A(mai_mai_n1188_), .B(mai_mai_n1255_), .Y(mai_mai_n1256_));
  INV        m1228(.A(mai_mai_n1256_), .Y(mai_mai_n1257_));
  NA4        m1229(.A(mai_mai_n1257_), .B(mai_mai_n1254_), .C(mai_mai_n1250_), .D(mai_mai_n1247_), .Y(mai_mai_n1258_));
  OR4        m1230(.A(mai_mai_n1258_), .B(mai_mai_n1240_), .C(mai_mai_n1203_), .D(mai_mai_n1190_), .Y(mai04));
  NOi31      m1231(.An(mai_mai_n1180_), .B(mai_mai_n1181_), .C(mai_mai_n878_), .Y(mai_mai_n1260_));
  NA2        m1232(.A(mai_mai_n1201_), .B(mai_mai_n703_), .Y(mai_mai_n1261_));
  NO2        m1233(.A(mai_mai_n1261_), .B(mai_mai_n872_), .Y(mai_mai_n1262_));
  OR3        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1260_), .C(mai_mai_n893_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n1145_), .B(mai_mai_n73_), .Y(mai_mai_n1264_));
  AOI210     m1236(.A0(mai_mai_n1264_), .A1(mai_mai_n887_), .B0(mai_mai_n1007_), .Y(mai_mai_n1265_));
  NA2        m1237(.A(mai_mai_n1265_), .B(mai_mai_n1031_), .Y(mai_mai_n1266_));
  NO4        m1238(.A(mai_mai_n1266_), .B(mai_mai_n1263_), .C(mai_mai_n901_), .D(mai_mai_n883_), .Y(mai_mai_n1267_));
  NA4        m1239(.A(mai_mai_n1267_), .B(mai_mai_n950_), .C(mai_mai_n939_), .D(mai_mai_n930_), .Y(mai05));
  INV        m1240(.A(m), .Y(mai_mai_n1271_));
  INV        m1241(.A(f), .Y(mai_mai_n1272_));
  INV        m1242(.A(mai_mai_n88_), .Y(mai_mai_n1273_));
  INV        m1243(.A(i), .Y(mai_mai_n1274_));
  INV        m1244(.A(j), .Y(mai_mai_n1275_));
  INV        m1245(.A(mai_mai_n96_), .Y(mai_mai_n1276_));
  INV        m1246(.A(j), .Y(mai_mai_n1277_));
  INV        m1247(.A(mai_mai_n191_), .Y(mai_mai_n1278_));
  INV        m1248(.A(m), .Y(mai_mai_n1279_));
  INV        m1249(.A(m), .Y(mai_mai_n1280_));
  INV        m1250(.A(mai_mai_n260_), .Y(mai_mai_n1281_));
  INV        m1251(.A(mai_mai_n356_), .Y(mai_mai_n1282_));
  INV        m1252(.A(a), .Y(mai_mai_n1283_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA2        u0003(.A(men_men_n31_), .B(men_men_n30_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(u), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(u), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(u), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(u), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(u), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  NO2        u0026(.A(men_men_n54_), .B(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA2        u0031(.A(u), .B(men_men_n59_), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(u), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(u), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(u), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(u), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(u), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(u), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n96_), .C(f), .Y(men_men_n98_));
  AN2        u0070(.A(j), .B(u), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(l), .C(i), .Y(men_men_n100_));
  NOi21      u0072(.An(u), .B(i), .Y(men_men_n101_));
  NOi32      u0073(.An(m), .Bn(j), .C(k), .Y(men_men_n102_));
  AOI220     u0074(.A0(men_men_n102_), .A1(men_men_n101_), .B0(men_men_n100_), .B1(men_men_n99_), .Y(men_men_n103_));
  NO2        u0075(.A(men_men_n103_), .B(f), .Y(men_men_n104_));
  NO4        u0076(.A(men_men_n104_), .B(men_men_n98_), .C(men_men_n95_), .D(men_men_n92_), .Y(men_men_n105_));
  NAi41      u0077(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n106_));
  AN2        u0078(.A(e), .B(b), .Y(men_men_n107_));
  NOi31      u0079(.An(c), .B(h), .C(f), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NOi21      u0081(.An(i), .B(h), .Y(men_men_n110_));
  NA3        u0082(.A(men_men_n110_), .B(u), .C(men_men_n36_), .Y(men_men_n111_));
  INV        u0083(.A(a), .Y(men_men_n112_));
  NA2        u0084(.A(men_men_n107_), .B(men_men_n112_), .Y(men_men_n113_));
  INV        u0085(.A(l), .Y(men_men_n114_));
  NOi21      u0086(.An(m), .B(n), .Y(men_men_n115_));
  NO2        u0087(.A(men_men_n111_), .B(men_men_n88_), .Y(men_men_n116_));
  INV        u0088(.A(b), .Y(men_men_n117_));
  NA2        u0089(.A(l), .B(j), .Y(men_men_n118_));
  AN2        u0090(.A(k), .B(i), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u0092(.A(u), .B(e), .Y(men_men_n121_));
  NOi32      u0093(.An(c), .Bn(a), .C(d), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n115_), .Y(men_men_n123_));
  NO4        u0095(.A(men_men_n123_), .B(men_men_n121_), .C(men_men_n120_), .D(men_men_n117_), .Y(men_men_n124_));
  NO2        u0096(.A(men_men_n124_), .B(men_men_n116_), .Y(men_men_n125_));
  OAI210     u0097(.A0(men_men_n105_), .A1(men_men_n88_), .B0(men_men_n125_), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(j), .Y(men_men_n127_));
  NA3        u0099(.A(men_men_n127_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n128_));
  NOi31      u0100(.An(k), .B(m), .C(i), .Y(men_men_n129_));
  NA3        u0101(.A(men_men_n129_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n130_));
  NA2        u0102(.A(men_men_n130_), .B(men_men_n128_), .Y(men_men_n131_));
  NOi32      u0103(.An(f), .Bn(b), .C(e), .Y(men_men_n132_));
  NAi21      u0104(.An(u), .B(h), .Y(men_men_n133_));
  NAi21      u0105(.An(m), .B(n), .Y(men_men_n134_));
  NAi21      u0106(.An(j), .B(k), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n133_), .Y(men_men_n136_));
  NAi41      u0108(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n137_));
  NAi31      u0109(.An(j), .B(k), .C(h), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n134_), .Y(men_men_n139_));
  AOI210     u0111(.A0(men_men_n136_), .A1(men_men_n132_), .B0(men_men_n139_), .Y(men_men_n140_));
  NO2        u0112(.A(k), .B(j), .Y(men_men_n141_));
  NO2        u0113(.A(men_men_n141_), .B(men_men_n134_), .Y(men_men_n142_));
  AN2        u0114(.A(k), .B(j), .Y(men_men_n143_));
  NAi21      u0115(.An(c), .B(b), .Y(men_men_n144_));
  NA2        u0116(.A(f), .B(d), .Y(men_men_n145_));
  NO4        u0117(.A(men_men_n145_), .B(men_men_n144_), .C(men_men_n143_), .D(men_men_n133_), .Y(men_men_n146_));
  NA2        u0118(.A(h), .B(c), .Y(men_men_n147_));
  NAi31      u0119(.An(f), .B(e), .C(b), .Y(men_men_n148_));
  NA2        u0120(.A(men_men_n146_), .B(men_men_n142_), .Y(men_men_n149_));
  NA2        u0121(.A(d), .B(b), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(f), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n151_), .B(men_men_n150_), .Y(men_men_n152_));
  NA2        u0124(.A(b), .B(a), .Y(men_men_n153_));
  NAi21      u0125(.An(c), .B(d), .Y(men_men_n154_));
  NAi31      u0126(.An(l), .B(k), .C(h), .Y(men_men_n155_));
  NO2        u0127(.A(men_men_n134_), .B(men_men_n155_), .Y(men_men_n156_));
  NA2        u0128(.A(men_men_n156_), .B(men_men_n152_), .Y(men_men_n157_));
  NAi41      u0129(.An(men_men_n131_), .B(men_men_n157_), .C(men_men_n149_), .D(men_men_n140_), .Y(men_men_n158_));
  NAi31      u0130(.An(e), .B(f), .C(b), .Y(men_men_n159_));
  NOi21      u0131(.An(u), .B(d), .Y(men_men_n160_));
  NO2        u0132(.A(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  NOi21      u0133(.An(h), .B(i), .Y(men_men_n162_));
  NOi21      u0134(.An(k), .B(m), .Y(men_men_n163_));
  NA3        u0135(.A(men_men_n163_), .B(men_men_n162_), .C(n), .Y(men_men_n164_));
  NOi21      u0136(.An(men_men_n161_), .B(men_men_n164_), .Y(men_men_n165_));
  NOi21      u0137(.An(h), .B(u), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n145_), .B(men_men_n144_), .Y(men_men_n167_));
  NA2        u0139(.A(men_men_n167_), .B(men_men_n166_), .Y(men_men_n168_));
  NAi31      u0140(.An(l), .B(j), .C(h), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n169_), .B(men_men_n49_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n67_), .Y(men_men_n171_));
  NOi32      u0143(.An(n), .Bn(k), .C(m), .Y(men_men_n172_));
  NA2        u0144(.A(l), .B(i), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  OAI210     u0146(.A0(men_men_n174_), .A1(men_men_n168_), .B0(men_men_n171_), .Y(men_men_n175_));
  NAi31      u0147(.An(d), .B(f), .C(c), .Y(men_men_n176_));
  NAi31      u0148(.An(e), .B(f), .C(c), .Y(men_men_n177_));
  NA2        u0149(.A(j), .B(h), .Y(men_men_n178_));
  OR3        u0150(.A(n), .B(m), .C(k), .Y(men_men_n179_));
  NAi32      u0151(.An(m), .Bn(k), .C(n), .Y(men_men_n180_));
  NO2        u0152(.A(men_men_n180_), .B(men_men_n178_), .Y(men_men_n181_));
  NA2        u0153(.A(men_men_n181_), .B(men_men_n161_), .Y(men_men_n182_));
  NO2        u0154(.A(n), .B(m), .Y(men_men_n183_));
  NA2        u0155(.A(men_men_n183_), .B(men_men_n50_), .Y(men_men_n184_));
  NAi21      u0156(.An(f), .B(e), .Y(men_men_n185_));
  NA2        u0157(.A(d), .B(c), .Y(men_men_n186_));
  NO2        u0158(.A(men_men_n186_), .B(men_men_n185_), .Y(men_men_n187_));
  NOi21      u0159(.An(men_men_n187_), .B(men_men_n184_), .Y(men_men_n188_));
  NAi31      u0160(.An(m), .B(n), .C(b), .Y(men_men_n189_));
  NAi21      u0161(.An(h), .B(f), .Y(men_men_n190_));
  NO2        u0162(.A(men_men_n189_), .B(men_men_n154_), .Y(men_men_n191_));
  NOi32      u0163(.An(f), .Bn(c), .C(d), .Y(men_men_n192_));
  NOi32      u0164(.An(f), .Bn(c), .C(e), .Y(men_men_n193_));
  NO2        u0165(.A(men_men_n193_), .B(men_men_n192_), .Y(men_men_n194_));
  NO3        u0166(.A(n), .B(m), .C(j), .Y(men_men_n195_));
  NA2        u0167(.A(men_men_n195_), .B(k), .Y(men_men_n196_));
  NAi21      u0168(.An(men_men_n188_), .B(men_men_n182_), .Y(men_men_n197_));
  OR4        u0169(.A(men_men_n197_), .B(men_men_n175_), .C(men_men_n165_), .D(men_men_n158_), .Y(men_men_n198_));
  NO4        u0170(.A(men_men_n198_), .B(men_men_n126_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n199_));
  NA3        u0171(.A(m), .B(men_men_n114_), .C(j), .Y(men_men_n200_));
  NAi31      u0172(.An(n), .B(h), .C(u), .Y(men_men_n201_));
  NO2        u0173(.A(men_men_n201_), .B(men_men_n200_), .Y(men_men_n202_));
  NOi32      u0174(.An(m), .Bn(k), .C(l), .Y(men_men_n203_));
  NA3        u0175(.A(men_men_n203_), .B(men_men_n89_), .C(u), .Y(men_men_n204_));
  NO2        u0176(.A(men_men_n204_), .B(n), .Y(men_men_n205_));
  NOi21      u0177(.An(k), .B(j), .Y(men_men_n206_));
  NA4        u0178(.A(men_men_n206_), .B(men_men_n115_), .C(i), .D(u), .Y(men_men_n207_));
  AN2        u0179(.A(i), .B(u), .Y(men_men_n208_));
  NA3        u0180(.A(men_men_n76_), .B(men_men_n208_), .C(men_men_n115_), .Y(men_men_n209_));
  NA2        u0181(.A(men_men_n209_), .B(men_men_n207_), .Y(men_men_n210_));
  NO3        u0182(.A(men_men_n210_), .B(men_men_n205_), .C(men_men_n202_), .Y(men_men_n211_));
  NAi41      u0183(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n212_));
  INV        u0184(.A(men_men_n212_), .Y(men_men_n213_));
  INV        u0185(.A(f), .Y(men_men_n214_));
  INV        u0186(.A(u), .Y(men_men_n215_));
  NOi31      u0187(.An(i), .B(j), .C(h), .Y(men_men_n216_));
  NOi21      u0188(.An(l), .B(m), .Y(men_men_n217_));
  NA2        u0189(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n218_));
  NO3        u0190(.A(men_men_n218_), .B(men_men_n215_), .C(men_men_n214_), .Y(men_men_n219_));
  NA2        u0191(.A(men_men_n219_), .B(men_men_n213_), .Y(men_men_n220_));
  OAI210     u0192(.A0(men_men_n211_), .A1(men_men_n32_), .B0(men_men_n220_), .Y(men_men_n221_));
  NOi21      u0193(.An(n), .B(m), .Y(men_men_n222_));
  NA2        u0194(.A(i), .B(men_men_n222_), .Y(men_men_n223_));
  OA220      u0195(.A0(men_men_n223_), .A1(men_men_n109_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n224_));
  NAi21      u0196(.An(j), .B(h), .Y(men_men_n225_));
  XN2        u0197(.A(i), .B(h), .Y(men_men_n226_));
  NOi31      u0198(.An(k), .B(n), .C(m), .Y(men_men_n227_));
  NAi31      u0199(.An(f), .B(e), .C(c), .Y(men_men_n228_));
  NA4        u0200(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n229_));
  NAi32      u0201(.An(m), .Bn(i), .C(k), .Y(men_men_n230_));
  NO3        u0202(.A(men_men_n230_), .B(men_men_n93_), .C(men_men_n229_), .Y(men_men_n231_));
  INV        u0203(.A(k), .Y(men_men_n232_));
  INV        u0204(.A(men_men_n231_), .Y(men_men_n233_));
  NAi21      u0205(.An(n), .B(a), .Y(men_men_n234_));
  NO2        u0206(.A(men_men_n234_), .B(men_men_n150_), .Y(men_men_n235_));
  NAi41      u0207(.An(u), .B(m), .C(k), .D(h), .Y(men_men_n236_));
  NO2        u0208(.A(men_men_n236_), .B(e), .Y(men_men_n237_));
  NO3        u0209(.A(men_men_n151_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n238_));
  NA2        u0210(.A(men_men_n238_), .B(men_men_n235_), .Y(men_men_n239_));
  AN3        u0211(.A(men_men_n239_), .B(men_men_n233_), .C(men_men_n224_), .Y(men_men_n240_));
  OR2        u0212(.A(h), .B(u), .Y(men_men_n241_));
  NAi41      u0213(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n242_));
  NO2        u0214(.A(men_men_n242_), .B(men_men_n214_), .Y(men_men_n243_));
  NA2        u0215(.A(men_men_n163_), .B(men_men_n110_), .Y(men_men_n244_));
  NAi21      u0216(.An(men_men_n244_), .B(men_men_n243_), .Y(men_men_n245_));
  NO2        u0217(.A(n), .B(a), .Y(men_men_n246_));
  NAi31      u0218(.An(men_men_n236_), .B(men_men_n246_), .C(men_men_n107_), .Y(men_men_n247_));
  AN2        u0219(.A(men_men_n247_), .B(men_men_n245_), .Y(men_men_n248_));
  NAi21      u0220(.An(h), .B(i), .Y(men_men_n249_));
  NA2        u0221(.A(men_men_n183_), .B(k), .Y(men_men_n250_));
  NO2        u0222(.A(men_men_n250_), .B(men_men_n249_), .Y(men_men_n251_));
  NA2        u0223(.A(men_men_n251_), .B(men_men_n192_), .Y(men_men_n252_));
  NA2        u0224(.A(men_men_n252_), .B(men_men_n248_), .Y(men_men_n253_));
  NOi21      u0225(.An(u), .B(e), .Y(men_men_n254_));
  NO2        u0226(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n255_), .B(men_men_n254_), .Y(men_men_n256_));
  NOi32      u0228(.An(l), .Bn(j), .C(i), .Y(men_men_n257_));
  AOI210     u0229(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n257_), .Y(men_men_n258_));
  NO2        u0230(.A(men_men_n249_), .B(men_men_n44_), .Y(men_men_n259_));
  NAi21      u0231(.An(f), .B(u), .Y(men_men_n260_));
  NO2        u0232(.A(men_men_n260_), .B(men_men_n65_), .Y(men_men_n261_));
  NO2        u0233(.A(men_men_n69_), .B(men_men_n118_), .Y(men_men_n262_));
  AOI220     u0234(.A0(men_men_n262_), .A1(men_men_n261_), .B0(men_men_n259_), .B1(men_men_n67_), .Y(men_men_n263_));
  OAI210     u0235(.A0(men_men_n258_), .A1(men_men_n256_), .B0(men_men_n263_), .Y(men_men_n264_));
  NO3        u0236(.A(men_men_n135_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n265_));
  NOi41      u0237(.An(men_men_n240_), .B(men_men_n264_), .C(men_men_n253_), .D(men_men_n221_), .Y(men_men_n266_));
  NO4        u0238(.A(men_men_n202_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n267_));
  NO2        u0239(.A(men_men_n267_), .B(men_men_n113_), .Y(men_men_n268_));
  NA3        u0240(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n269_));
  NAi21      u0241(.An(h), .B(u), .Y(men_men_n270_));
  OR4        u0242(.A(men_men_n270_), .B(men_men_n269_), .C(men_men_n223_), .D(e), .Y(men_men_n271_));
  NO2        u0243(.A(men_men_n244_), .B(men_men_n260_), .Y(men_men_n272_));
  NAi31      u0244(.An(u), .B(k), .C(h), .Y(men_men_n273_));
  NO3        u0245(.A(men_men_n134_), .B(men_men_n273_), .C(l), .Y(men_men_n274_));
  NAi31      u0246(.An(e), .B(d), .C(a), .Y(men_men_n275_));
  NA2        u0247(.A(men_men_n274_), .B(men_men_n132_), .Y(men_men_n276_));
  NA2        u0248(.A(men_men_n276_), .B(men_men_n271_), .Y(men_men_n277_));
  NA4        u0249(.A(men_men_n163_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n118_), .Y(men_men_n278_));
  NA3        u0250(.A(men_men_n163_), .B(men_men_n162_), .C(men_men_n86_), .Y(men_men_n279_));
  NO2        u0251(.A(men_men_n279_), .B(men_men_n194_), .Y(men_men_n280_));
  NOi21      u0252(.An(men_men_n278_), .B(men_men_n280_), .Y(men_men_n281_));
  NA3        u0253(.A(e), .B(c), .C(b), .Y(men_men_n282_));
  NO2        u0254(.A(men_men_n60_), .B(men_men_n282_), .Y(men_men_n283_));
  NAi32      u0255(.An(k), .Bn(i), .C(j), .Y(men_men_n284_));
  NAi31      u0256(.An(h), .B(l), .C(i), .Y(men_men_n285_));
  NA3        u0257(.A(men_men_n285_), .B(men_men_n284_), .C(men_men_n169_), .Y(men_men_n286_));
  NOi21      u0258(.An(men_men_n286_), .B(men_men_n49_), .Y(men_men_n287_));
  OAI210     u0259(.A0(men_men_n261_), .A1(men_men_n283_), .B0(men_men_n287_), .Y(men_men_n288_));
  NAi21      u0260(.An(l), .B(k), .Y(men_men_n289_));
  NO2        u0261(.A(men_men_n289_), .B(men_men_n49_), .Y(men_men_n290_));
  NOi21      u0262(.An(l), .B(j), .Y(men_men_n291_));
  INV        u0263(.A(men_men_n166_), .Y(men_men_n292_));
  NA3        u0264(.A(men_men_n119_), .B(men_men_n118_), .C(u), .Y(men_men_n293_));
  OR3        u0265(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n294_));
  AOI210     u0266(.A0(men_men_n293_), .A1(men_men_n292_), .B0(men_men_n294_), .Y(men_men_n295_));
  INV        u0267(.A(men_men_n295_), .Y(men_men_n296_));
  NAi32      u0268(.An(j), .Bn(h), .C(i), .Y(men_men_n297_));
  NAi21      u0269(.An(m), .B(l), .Y(men_men_n298_));
  NO3        u0270(.A(men_men_n298_), .B(men_men_n297_), .C(men_men_n86_), .Y(men_men_n299_));
  NA2        u0271(.A(h), .B(u), .Y(men_men_n300_));
  NA2        u0272(.A(men_men_n172_), .B(men_men_n45_), .Y(men_men_n301_));
  NO2        u0273(.A(men_men_n301_), .B(men_men_n300_), .Y(men_men_n302_));
  OAI210     u0274(.A0(men_men_n302_), .A1(men_men_n299_), .B0(men_men_n167_), .Y(men_men_n303_));
  NA4        u0275(.A(men_men_n303_), .B(men_men_n296_), .C(men_men_n288_), .D(men_men_n281_), .Y(men_men_n304_));
  NO2        u0276(.A(men_men_n148_), .B(d), .Y(men_men_n305_));
  NA2        u0277(.A(men_men_n305_), .B(men_men_n53_), .Y(men_men_n306_));
  NAi32      u0278(.An(n), .Bn(m), .C(l), .Y(men_men_n307_));
  NO2        u0279(.A(men_men_n307_), .B(men_men_n297_), .Y(men_men_n308_));
  NA2        u0280(.A(men_men_n308_), .B(men_men_n187_), .Y(men_men_n309_));
  NO2        u0281(.A(men_men_n123_), .B(men_men_n117_), .Y(men_men_n310_));
  NAi31      u0282(.An(k), .B(l), .C(j), .Y(men_men_n311_));
  OAI210     u0283(.A0(men_men_n289_), .A1(j), .B0(men_men_n311_), .Y(men_men_n312_));
  NOi21      u0284(.An(men_men_n312_), .B(men_men_n121_), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n313_), .B(men_men_n310_), .Y(men_men_n314_));
  NA3        u0286(.A(men_men_n314_), .B(men_men_n309_), .C(men_men_n306_), .Y(men_men_n315_));
  NO4        u0287(.A(men_men_n315_), .B(men_men_n304_), .C(men_men_n277_), .D(men_men_n268_), .Y(men_men_n316_));
  NAi21      u0288(.An(m), .B(k), .Y(men_men_n317_));
  NO2        u0289(.A(men_men_n226_), .B(men_men_n317_), .Y(men_men_n318_));
  NAi41      u0290(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n319_));
  NAi31      u0291(.An(i), .B(l), .C(h), .Y(men_men_n320_));
  NO4        u0292(.A(men_men_n320_), .B(e), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n321_));
  NA2        u0293(.A(e), .B(c), .Y(men_men_n322_));
  NO3        u0294(.A(men_men_n322_), .B(n), .C(d), .Y(men_men_n323_));
  NOi21      u0295(.An(f), .B(h), .Y(men_men_n324_));
  NAi31      u0296(.An(d), .B(e), .C(b), .Y(men_men_n325_));
  NO2        u0297(.A(men_men_n134_), .B(men_men_n325_), .Y(men_men_n326_));
  NO4        u0298(.A(men_men_n319_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n215_), .Y(men_men_n327_));
  NA2        u0299(.A(men_men_n246_), .B(men_men_n107_), .Y(men_men_n328_));
  NOi31      u0300(.An(l), .B(n), .C(m), .Y(men_men_n329_));
  NAi32      u0301(.An(m), .Bn(j), .C(k), .Y(men_men_n330_));
  NAi41      u0302(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n331_));
  NA2        u0303(.A(men_men_n212_), .B(men_men_n331_), .Y(men_men_n332_));
  NOi31      u0304(.An(j), .B(m), .C(k), .Y(men_men_n333_));
  NO2        u0305(.A(men_men_n127_), .B(men_men_n333_), .Y(men_men_n334_));
  AN3        u0306(.A(h), .B(u), .C(f), .Y(men_men_n335_));
  NAi31      u0307(.An(men_men_n334_), .B(men_men_n335_), .C(men_men_n332_), .Y(men_men_n336_));
  NOi32      u0308(.An(m), .Bn(j), .C(l), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n337_), .B(men_men_n100_), .Y(men_men_n338_));
  NAi32      u0310(.An(men_men_n338_), .Bn(men_men_n201_), .C(men_men_n305_), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n298_), .B(men_men_n297_), .Y(men_men_n340_));
  NO2        u0312(.A(men_men_n218_), .B(u), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n159_), .B(men_men_n86_), .Y(men_men_n342_));
  AOI220     u0314(.A0(men_men_n342_), .A1(men_men_n341_), .B0(men_men_n243_), .B1(men_men_n340_), .Y(men_men_n343_));
  INV        u0315(.A(men_men_n230_), .Y(men_men_n344_));
  NA3        u0316(.A(men_men_n344_), .B(men_men_n335_), .C(men_men_n213_), .Y(men_men_n345_));
  NA4        u0317(.A(men_men_n345_), .B(men_men_n343_), .C(men_men_n339_), .D(men_men_n336_), .Y(men_men_n346_));
  NA3        u0318(.A(h), .B(u), .C(f), .Y(men_men_n347_));
  NO2        u0319(.A(men_men_n347_), .B(men_men_n77_), .Y(men_men_n348_));
  NA2        u0320(.A(men_men_n331_), .B(men_men_n212_), .Y(men_men_n349_));
  NA2        u0321(.A(men_men_n166_), .B(e), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n350_), .B(men_men_n41_), .Y(men_men_n351_));
  AOI220     u0323(.A0(men_men_n351_), .A1(men_men_n310_), .B0(men_men_n349_), .B1(men_men_n348_), .Y(men_men_n352_));
  NOi32      u0324(.An(j), .Bn(u), .C(i), .Y(men_men_n353_));
  NA3        u0325(.A(men_men_n353_), .B(men_men_n289_), .C(men_men_n115_), .Y(men_men_n354_));
  AO210      u0326(.A0(men_men_n113_), .A1(men_men_n32_), .B0(men_men_n354_), .Y(men_men_n355_));
  NOi32      u0327(.An(e), .Bn(b), .C(a), .Y(men_men_n356_));
  AN2        u0328(.A(l), .B(j), .Y(men_men_n357_));
  NO2        u0329(.A(men_men_n317_), .B(men_men_n357_), .Y(men_men_n358_));
  NO3        u0330(.A(men_men_n319_), .B(men_men_n72_), .C(men_men_n215_), .Y(men_men_n359_));
  NA3        u0331(.A(men_men_n209_), .B(men_men_n207_), .C(men_men_n35_), .Y(men_men_n360_));
  AOI220     u0332(.A0(men_men_n360_), .A1(men_men_n356_), .B0(men_men_n359_), .B1(men_men_n358_), .Y(men_men_n361_));
  NO2        u0333(.A(men_men_n325_), .B(n), .Y(men_men_n362_));
  NA2        u0334(.A(men_men_n208_), .B(k), .Y(men_men_n363_));
  NA3        u0335(.A(m), .B(men_men_n114_), .C(men_men_n214_), .Y(men_men_n364_));
  NA4        u0336(.A(men_men_n203_), .B(men_men_n89_), .C(u), .D(men_men_n214_), .Y(men_men_n365_));
  OAI210     u0337(.A0(men_men_n364_), .A1(men_men_n363_), .B0(men_men_n365_), .Y(men_men_n366_));
  NAi41      u0338(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n367_));
  NA2        u0339(.A(men_men_n51_), .B(men_men_n115_), .Y(men_men_n368_));
  NO2        u0340(.A(men_men_n368_), .B(men_men_n367_), .Y(men_men_n369_));
  NA2        u0341(.A(men_men_n366_), .B(men_men_n362_), .Y(men_men_n370_));
  NA4        u0342(.A(men_men_n370_), .B(men_men_n361_), .C(men_men_n355_), .D(men_men_n352_), .Y(men_men_n371_));
  NO4        u0343(.A(men_men_n371_), .B(men_men_n346_), .C(men_men_n327_), .D(men_men_n321_), .Y(men_men_n372_));
  NA4        u0344(.A(men_men_n372_), .B(men_men_n316_), .C(men_men_n266_), .D(men_men_n199_), .Y(men10));
  NA3        u0345(.A(m), .B(k), .C(i), .Y(men_men_n374_));
  NO3        u0346(.A(men_men_n374_), .B(j), .C(men_men_n215_), .Y(men_men_n375_));
  NOi21      u0347(.An(e), .B(f), .Y(men_men_n376_));
  NO4        u0348(.A(men_men_n154_), .B(men_men_n376_), .C(n), .D(men_men_n112_), .Y(men_men_n377_));
  NAi31      u0349(.An(b), .B(f), .C(c), .Y(men_men_n378_));
  INV        u0350(.A(men_men_n378_), .Y(men_men_n379_));
  NOi32      u0351(.An(k), .Bn(h), .C(j), .Y(men_men_n380_));
  NA2        u0352(.A(men_men_n380_), .B(men_men_n222_), .Y(men_men_n381_));
  NA2        u0353(.A(men_men_n164_), .B(men_men_n381_), .Y(men_men_n382_));
  AOI220     u0354(.A0(men_men_n382_), .A1(men_men_n379_), .B0(men_men_n377_), .B1(men_men_n375_), .Y(men_men_n383_));
  AN2        u0355(.A(j), .B(h), .Y(men_men_n384_));
  NA4        u0356(.A(n), .B(f), .C(c), .D(men_men_n117_), .Y(men_men_n385_));
  NOi32      u0357(.An(d), .Bn(a), .C(c), .Y(men_men_n386_));
  NA2        u0358(.A(men_men_n386_), .B(men_men_n185_), .Y(men_men_n387_));
  NAi31      u0359(.An(k), .B(m), .C(j), .Y(men_men_n388_));
  NO3        u0360(.A(men_men_n388_), .B(i), .C(n), .Y(men_men_n389_));
  NOi21      u0361(.An(men_men_n389_), .B(men_men_n387_), .Y(men_men_n390_));
  INV        u0362(.A(men_men_n390_), .Y(men_men_n391_));
  NO2        u0363(.A(men_men_n385_), .B(men_men_n298_), .Y(men_men_n392_));
  NOi32      u0364(.An(f), .Bn(d), .C(c), .Y(men_men_n393_));
  AOI220     u0365(.A0(men_men_n393_), .A1(men_men_n308_), .B0(men_men_n392_), .B1(men_men_n216_), .Y(men_men_n394_));
  NA3        u0366(.A(men_men_n394_), .B(men_men_n391_), .C(men_men_n383_), .Y(men_men_n395_));
  NO2        u0367(.A(men_men_n59_), .B(men_men_n117_), .Y(men_men_n396_));
  NA2        u0368(.A(men_men_n246_), .B(men_men_n396_), .Y(men_men_n397_));
  INV        u0369(.A(e), .Y(men_men_n398_));
  NA2        u0370(.A(men_men_n46_), .B(e), .Y(men_men_n399_));
  OAI220     u0371(.A0(men_men_n399_), .A1(men_men_n200_), .B0(men_men_n204_), .B1(men_men_n398_), .Y(men_men_n400_));
  AN2        u0372(.A(u), .B(e), .Y(men_men_n401_));
  NA3        u0373(.A(men_men_n401_), .B(men_men_n203_), .C(i), .Y(men_men_n402_));
  NA2        u0374(.A(men_men_n91_), .B(men_men_n402_), .Y(men_men_n403_));
  NO2        u0375(.A(men_men_n103_), .B(men_men_n398_), .Y(men_men_n404_));
  NO3        u0376(.A(men_men_n404_), .B(men_men_n403_), .C(men_men_n400_), .Y(men_men_n405_));
  NOi32      u0377(.An(h), .Bn(e), .C(u), .Y(men_men_n406_));
  NA2        u0378(.A(men_men_n406_), .B(m), .Y(men_men_n407_));
  NOi21      u0379(.An(u), .B(h), .Y(men_men_n408_));
  AN3        u0380(.A(m), .B(l), .C(i), .Y(men_men_n409_));
  AN3        u0381(.A(h), .B(u), .C(e), .Y(men_men_n410_));
  NA2        u0382(.A(men_men_n410_), .B(men_men_n100_), .Y(men_men_n411_));
  AOI210     u0383(.A0(men_men_n407_), .A1(men_men_n405_), .B0(men_men_n397_), .Y(men_men_n412_));
  NA3        u0384(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n413_));
  NO2        u0385(.A(men_men_n413_), .B(men_men_n397_), .Y(men_men_n414_));
  NA2        u0386(.A(men_men_n386_), .B(men_men_n86_), .Y(men_men_n415_));
  NAi31      u0387(.An(b), .B(c), .C(a), .Y(men_men_n416_));
  NO2        u0388(.A(men_men_n416_), .B(n), .Y(men_men_n417_));
  OAI210     u0389(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n418_));
  NO2        u0390(.A(men_men_n418_), .B(men_men_n151_), .Y(men_men_n419_));
  NA2        u0391(.A(men_men_n419_), .B(men_men_n417_), .Y(men_men_n420_));
  INV        u0392(.A(men_men_n420_), .Y(men_men_n421_));
  NO4        u0393(.A(men_men_n421_), .B(men_men_n414_), .C(men_men_n412_), .D(men_men_n395_), .Y(men_men_n422_));
  NA2        u0394(.A(i), .B(u), .Y(men_men_n423_));
  NO3        u0395(.A(men_men_n275_), .B(men_men_n423_), .C(c), .Y(men_men_n424_));
  NOi21      u0396(.An(d), .B(c), .Y(men_men_n425_));
  NA2        u0397(.A(men_men_n425_), .B(a), .Y(men_men_n426_));
  NA3        u0398(.A(i), .B(u), .C(f), .Y(men_men_n427_));
  OR2        u0399(.A(men_men_n427_), .B(men_men_n71_), .Y(men_men_n428_));
  NA2        u0400(.A(men_men_n409_), .B(men_men_n408_), .Y(men_men_n429_));
  AOI210     u0401(.A0(men_men_n429_), .A1(men_men_n428_), .B0(men_men_n426_), .Y(men_men_n430_));
  AOI210     u0402(.A0(men_men_n424_), .A1(men_men_n290_), .B0(men_men_n430_), .Y(men_men_n431_));
  OR2        u0403(.A(n), .B(m), .Y(men_men_n432_));
  NO2        u0404(.A(men_men_n416_), .B(men_men_n49_), .Y(men_men_n433_));
  NO3        u0405(.A(men_men_n66_), .B(men_men_n114_), .C(e), .Y(men_men_n434_));
  NAi21      u0406(.An(k), .B(j), .Y(men_men_n435_));
  NA2        u0407(.A(men_men_n434_), .B(men_men_n433_), .Y(men_men_n436_));
  NAi21      u0408(.An(e), .B(d), .Y(men_men_n437_));
  NO2        u0409(.A(men_men_n250_), .B(men_men_n214_), .Y(men_men_n438_));
  NOi31      u0410(.An(n), .B(m), .C(k), .Y(men_men_n439_));
  AOI220     u0411(.A0(men_men_n439_), .A1(men_men_n384_), .B0(men_men_n222_), .B1(men_men_n50_), .Y(men_men_n440_));
  NAi31      u0412(.An(u), .B(f), .C(c), .Y(men_men_n441_));
  OR3        u0413(.A(men_men_n441_), .B(men_men_n440_), .C(e), .Y(men_men_n442_));
  NA2        u0414(.A(men_men_n442_), .B(men_men_n309_), .Y(men_men_n443_));
  NOi41      u0415(.An(men_men_n431_), .B(men_men_n443_), .C(men_men_n1449_), .D(men_men_n264_), .Y(men_men_n444_));
  NOi32      u0416(.An(c), .Bn(a), .C(b), .Y(men_men_n445_));
  NA2        u0417(.A(men_men_n445_), .B(men_men_n115_), .Y(men_men_n446_));
  INV        u0418(.A(men_men_n273_), .Y(men_men_n447_));
  AN2        u0419(.A(e), .B(d), .Y(men_men_n448_));
  NA2        u0420(.A(men_men_n448_), .B(men_men_n447_), .Y(men_men_n449_));
  INV        u0421(.A(men_men_n151_), .Y(men_men_n450_));
  NO2        u0422(.A(men_men_n133_), .B(men_men_n41_), .Y(men_men_n451_));
  NO2        u0423(.A(men_men_n66_), .B(e), .Y(men_men_n452_));
  NOi31      u0424(.An(j), .B(k), .C(i), .Y(men_men_n453_));
  NOi21      u0425(.An(men_men_n169_), .B(men_men_n453_), .Y(men_men_n454_));
  NA2        u0426(.A(men_men_n454_), .B(men_men_n258_), .Y(men_men_n455_));
  AOI220     u0427(.A0(men_men_n455_), .A1(men_men_n452_), .B0(men_men_n451_), .B1(men_men_n450_), .Y(men_men_n456_));
  AOI210     u0428(.A0(men_men_n456_), .A1(men_men_n449_), .B0(men_men_n446_), .Y(men_men_n457_));
  NO2        u0429(.A(men_men_n210_), .B(men_men_n205_), .Y(men_men_n458_));
  NOi21      u0430(.An(a), .B(b), .Y(men_men_n459_));
  NA3        u0431(.A(e), .B(d), .C(c), .Y(men_men_n460_));
  NAi21      u0432(.An(men_men_n460_), .B(men_men_n459_), .Y(men_men_n461_));
  NO2        u0433(.A(men_men_n415_), .B(men_men_n204_), .Y(men_men_n462_));
  NOi21      u0434(.An(men_men_n461_), .B(men_men_n462_), .Y(men_men_n463_));
  AOI210     u0435(.A0(men_men_n267_), .A1(men_men_n458_), .B0(men_men_n463_), .Y(men_men_n464_));
  NO4        u0436(.A(men_men_n190_), .B(men_men_n106_), .C(men_men_n56_), .D(b), .Y(men_men_n465_));
  NA2        u0437(.A(men_men_n379_), .B(men_men_n156_), .Y(men_men_n466_));
  NA2        u0438(.A(l), .B(k), .Y(men_men_n467_));
  NA3        u0439(.A(men_men_n467_), .B(j), .C(men_men_n222_), .Y(men_men_n468_));
  AOI210     u0440(.A0(men_men_n230_), .A1(men_men_n330_), .B0(men_men_n86_), .Y(men_men_n469_));
  NOi21      u0441(.An(men_men_n468_), .B(men_men_n469_), .Y(men_men_n470_));
  OR3        u0442(.A(men_men_n470_), .B(men_men_n147_), .C(men_men_n137_), .Y(men_men_n471_));
  NA3        u0443(.A(men_men_n278_), .B(men_men_n130_), .C(men_men_n128_), .Y(men_men_n472_));
  NA2        u0444(.A(men_men_n386_), .B(men_men_n115_), .Y(men_men_n473_));
  NO4        u0445(.A(men_men_n473_), .B(men_men_n97_), .C(men_men_n114_), .D(e), .Y(men_men_n474_));
  NO3        u0446(.A(men_men_n415_), .B(men_men_n94_), .C(men_men_n133_), .Y(men_men_n475_));
  NO4        u0447(.A(men_men_n475_), .B(men_men_n474_), .C(men_men_n472_), .D(men_men_n321_), .Y(men_men_n476_));
  NA3        u0448(.A(men_men_n476_), .B(men_men_n471_), .C(men_men_n466_), .Y(men_men_n477_));
  NO3        u0449(.A(men_men_n477_), .B(men_men_n464_), .C(men_men_n457_), .Y(men_men_n478_));
  NA2        u0450(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n479_));
  NO2        u0451(.A(men_men_n190_), .B(men_men_n56_), .Y(men_men_n480_));
  NAi31      u0452(.An(j), .B(l), .C(i), .Y(men_men_n481_));
  OAI210     u0453(.A0(men_men_n481_), .A1(men_men_n134_), .B0(men_men_n106_), .Y(men_men_n482_));
  NA2        u0454(.A(men_men_n482_), .B(men_men_n480_), .Y(men_men_n483_));
  NO3        u0455(.A(men_men_n387_), .B(men_men_n338_), .C(men_men_n201_), .Y(men_men_n484_));
  NO2        u0456(.A(men_men_n387_), .B(men_men_n368_), .Y(men_men_n485_));
  NO3        u0457(.A(men_men_n485_), .B(men_men_n484_), .C(men_men_n188_), .Y(men_men_n486_));
  NA4        u0458(.A(men_men_n486_), .B(men_men_n483_), .C(men_men_n479_), .D(men_men_n240_), .Y(men_men_n487_));
  OAI210     u0459(.A0(men_men_n129_), .A1(men_men_n127_), .B0(n), .Y(men_men_n488_));
  NO2        u0460(.A(men_men_n488_), .B(men_men_n133_), .Y(men_men_n489_));
  AN2        u0461(.A(men_men_n489_), .B(men_men_n193_), .Y(men_men_n490_));
  XO2        u0462(.A(i), .B(h), .Y(men_men_n491_));
  NA3        u0463(.A(men_men_n491_), .B(men_men_n163_), .C(n), .Y(men_men_n492_));
  NAi41      u0464(.An(men_men_n299_), .B(men_men_n492_), .C(men_men_n440_), .D(men_men_n381_), .Y(men_men_n493_));
  NOi32      u0465(.An(men_men_n493_), .Bn(men_men_n452_), .C(men_men_n269_), .Y(men_men_n494_));
  NAi31      u0466(.An(c), .B(f), .C(d), .Y(men_men_n495_));
  AOI210     u0467(.A0(men_men_n279_), .A1(men_men_n196_), .B0(men_men_n495_), .Y(men_men_n496_));
  NOi21      u0468(.An(men_men_n84_), .B(men_men_n496_), .Y(men_men_n497_));
  NA3        u0469(.A(men_men_n377_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n498_));
  NA2        u0470(.A(men_men_n227_), .B(men_men_n110_), .Y(men_men_n499_));
  AOI210     u0471(.A0(men_men_n354_), .A1(men_men_n35_), .B0(men_men_n461_), .Y(men_men_n500_));
  NOi21      u0472(.An(men_men_n498_), .B(men_men_n500_), .Y(men_men_n501_));
  AO220      u0473(.A0(men_men_n287_), .A1(men_men_n261_), .B0(men_men_n170_), .B1(men_men_n67_), .Y(men_men_n502_));
  NA3        u0474(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n503_));
  NO2        u0475(.A(men_men_n503_), .B(men_men_n426_), .Y(men_men_n504_));
  NO2        u0476(.A(men_men_n504_), .B(men_men_n295_), .Y(men_men_n505_));
  NAi41      u0477(.An(men_men_n502_), .B(men_men_n505_), .C(men_men_n501_), .D(men_men_n497_), .Y(men_men_n506_));
  NO4        u0478(.A(men_men_n506_), .B(men_men_n494_), .C(men_men_n490_), .D(men_men_n487_), .Y(men_men_n507_));
  NA4        u0479(.A(men_men_n507_), .B(men_men_n478_), .C(men_men_n444_), .D(men_men_n422_), .Y(men11));
  NO2        u0480(.A(men_men_n73_), .B(f), .Y(men_men_n509_));
  NA2        u0481(.A(j), .B(u), .Y(men_men_n510_));
  NAi31      u0482(.An(i), .B(m), .C(l), .Y(men_men_n511_));
  NA3        u0483(.A(m), .B(k), .C(j), .Y(men_men_n512_));
  OAI220     u0484(.A0(men_men_n512_), .A1(men_men_n133_), .B0(men_men_n511_), .B1(men_men_n510_), .Y(men_men_n513_));
  NA2        u0485(.A(men_men_n513_), .B(men_men_n509_), .Y(men_men_n514_));
  NOi32      u0486(.An(e), .Bn(b), .C(f), .Y(men_men_n515_));
  NA2        u0487(.A(men_men_n257_), .B(men_men_n115_), .Y(men_men_n516_));
  NA2        u0488(.A(men_men_n46_), .B(j), .Y(men_men_n517_));
  NO2        u0489(.A(men_men_n517_), .B(men_men_n301_), .Y(men_men_n518_));
  NAi31      u0490(.An(d), .B(e), .C(a), .Y(men_men_n519_));
  NO2        u0491(.A(men_men_n519_), .B(n), .Y(men_men_n520_));
  AOI220     u0492(.A0(men_men_n520_), .A1(men_men_n104_), .B0(men_men_n518_), .B1(men_men_n515_), .Y(men_men_n521_));
  NAi41      u0493(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n522_));
  AN2        u0494(.A(men_men_n522_), .B(men_men_n367_), .Y(men_men_n523_));
  AOI210     u0495(.A0(men_men_n523_), .A1(men_men_n387_), .B0(men_men_n270_), .Y(men_men_n524_));
  NA2        u0496(.A(j), .B(i), .Y(men_men_n525_));
  NAi31      u0497(.An(n), .B(m), .C(k), .Y(men_men_n526_));
  NO3        u0498(.A(men_men_n526_), .B(men_men_n525_), .C(men_men_n114_), .Y(men_men_n527_));
  NO4        u0499(.A(n), .B(d), .C(men_men_n117_), .D(a), .Y(men_men_n528_));
  NO2        u0500(.A(c), .B(men_men_n153_), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n529_), .B(men_men_n528_), .Y(men_men_n530_));
  NOi32      u0502(.An(u), .Bn(f), .C(i), .Y(men_men_n531_));
  AOI220     u0503(.A0(men_men_n531_), .A1(men_men_n102_), .B0(men_men_n513_), .B1(f), .Y(men_men_n532_));
  NO2        u0504(.A(men_men_n532_), .B(men_men_n530_), .Y(men_men_n533_));
  AOI210     u0505(.A0(men_men_n527_), .A1(men_men_n524_), .B0(men_men_n533_), .Y(men_men_n534_));
  NA2        u0506(.A(men_men_n143_), .B(men_men_n34_), .Y(men_men_n535_));
  NOi41      u0507(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n536_));
  NAi32      u0508(.An(e), .Bn(b), .C(c), .Y(men_men_n537_));
  AN2        u0509(.A(men_men_n331_), .B(men_men_n319_), .Y(men_men_n538_));
  NA2        u0510(.A(men_men_n538_), .B(men_men_n537_), .Y(men_men_n539_));
  OAI220     u0511(.A0(men_men_n388_), .A1(i), .B0(men_men_n511_), .B1(men_men_n510_), .Y(men_men_n540_));
  NAi31      u0512(.An(d), .B(c), .C(a), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n541_), .B(n), .Y(men_men_n542_));
  NA3        u0514(.A(men_men_n542_), .B(men_men_n540_), .C(e), .Y(men_men_n543_));
  NO3        u0515(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n215_), .Y(men_men_n544_));
  NO2        u0516(.A(men_men_n228_), .B(men_men_n112_), .Y(men_men_n545_));
  OAI210     u0517(.A0(men_men_n544_), .A1(men_men_n389_), .B0(men_men_n545_), .Y(men_men_n546_));
  NA2        u0518(.A(men_men_n546_), .B(men_men_n543_), .Y(men_men_n547_));
  NO2        u0519(.A(men_men_n275_), .B(n), .Y(men_men_n548_));
  NO2        u0520(.A(men_men_n417_), .B(men_men_n548_), .Y(men_men_n549_));
  NA2        u0521(.A(men_men_n540_), .B(f), .Y(men_men_n550_));
  NAi32      u0522(.An(d), .Bn(a), .C(b), .Y(men_men_n551_));
  NO3        u0523(.A(men_men_n180_), .B(men_men_n178_), .C(u), .Y(men_men_n552_));
  NA2        u0524(.A(men_men_n552_), .B(men_men_n58_), .Y(men_men_n553_));
  OAI210     u0525(.A0(men_men_n550_), .A1(men_men_n549_), .B0(men_men_n553_), .Y(men_men_n554_));
  AN3        u0526(.A(j), .B(h), .C(u), .Y(men_men_n555_));
  NO2        u0527(.A(men_men_n150_), .B(c), .Y(men_men_n556_));
  NA3        u0528(.A(men_men_n556_), .B(men_men_n555_), .C(men_men_n439_), .Y(men_men_n557_));
  NA3        u0529(.A(f), .B(d), .C(b), .Y(men_men_n558_));
  NO4        u0530(.A(men_men_n558_), .B(men_men_n180_), .C(men_men_n178_), .D(u), .Y(men_men_n559_));
  NAi21      u0531(.An(men_men_n559_), .B(men_men_n557_), .Y(men_men_n560_));
  NO3        u0532(.A(men_men_n560_), .B(men_men_n554_), .C(men_men_n547_), .Y(men_men_n561_));
  AN4        u0533(.A(men_men_n561_), .B(men_men_n534_), .C(men_men_n521_), .D(men_men_n514_), .Y(men_men_n562_));
  INV        u0534(.A(k), .Y(men_men_n563_));
  NA3        u0535(.A(l), .B(men_men_n563_), .C(i), .Y(men_men_n564_));
  INV        u0536(.A(men_men_n564_), .Y(men_men_n565_));
  NA3        u0537(.A(men_men_n386_), .B(men_men_n408_), .C(men_men_n115_), .Y(men_men_n566_));
  NAi32      u0538(.An(h), .Bn(f), .C(u), .Y(men_men_n567_));
  NAi41      u0539(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n568_));
  OAI210     u0540(.A0(men_men_n519_), .A1(n), .B0(men_men_n568_), .Y(men_men_n569_));
  NA2        u0541(.A(men_men_n569_), .B(m), .Y(men_men_n570_));
  NAi31      u0542(.An(h), .B(u), .C(f), .Y(men_men_n571_));
  OR3        u0543(.A(men_men_n571_), .B(men_men_n275_), .C(men_men_n49_), .Y(men_men_n572_));
  NA4        u0544(.A(men_men_n408_), .B(men_men_n122_), .C(men_men_n115_), .D(e), .Y(men_men_n573_));
  AN2        u0545(.A(men_men_n573_), .B(men_men_n572_), .Y(men_men_n574_));
  OA210      u0546(.A0(men_men_n570_), .A1(men_men_n567_), .B0(men_men_n574_), .Y(men_men_n575_));
  NO3        u0547(.A(men_men_n567_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n576_));
  NO4        u0548(.A(men_men_n571_), .B(c), .C(men_men_n153_), .D(men_men_n75_), .Y(men_men_n577_));
  OR2        u0549(.A(men_men_n577_), .B(men_men_n576_), .Y(men_men_n578_));
  NAi31      u0550(.An(men_men_n578_), .B(men_men_n575_), .C(men_men_n566_), .Y(men_men_n579_));
  NAi31      u0551(.An(f), .B(h), .C(u), .Y(men_men_n580_));
  NO4        u0552(.A(men_men_n311_), .B(men_men_n580_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n581_));
  NOi21      u0553(.An(b), .B(c), .Y(men_men_n582_));
  NO3        u0554(.A(men_men_n347_), .B(men_men_n69_), .C(men_men_n118_), .Y(men_men_n583_));
  OR2        u0555(.A(men_men_n583_), .B(men_men_n581_), .Y(men_men_n584_));
  NOi32      u0556(.An(d), .Bn(a), .C(e), .Y(men_men_n585_));
  NA2        u0557(.A(men_men_n585_), .B(men_men_n115_), .Y(men_men_n586_));
  NO2        u0558(.A(n), .B(c), .Y(men_men_n587_));
  NA3        u0559(.A(men_men_n587_), .B(men_men_n29_), .C(m), .Y(men_men_n588_));
  NAi32      u0560(.An(n), .Bn(f), .C(m), .Y(men_men_n589_));
  NA3        u0561(.A(men_men_n589_), .B(men_men_n588_), .C(men_men_n586_), .Y(men_men_n590_));
  NOi32      u0562(.An(e), .Bn(a), .C(d), .Y(men_men_n591_));
  AOI210     u0563(.A0(men_men_n29_), .A1(d), .B0(men_men_n591_), .Y(men_men_n592_));
  INV        u0564(.A(men_men_n535_), .Y(men_men_n593_));
  AOI210     u0565(.A0(men_men_n593_), .A1(men_men_n590_), .B0(men_men_n584_), .Y(men_men_n594_));
  OAI210     u0566(.A0(men_men_n245_), .A1(men_men_n89_), .B0(men_men_n594_), .Y(men_men_n595_));
  AOI210     u0567(.A0(men_men_n579_), .A1(men_men_n565_), .B0(men_men_n595_), .Y(men_men_n596_));
  NO3        u0568(.A(men_men_n317_), .B(men_men_n61_), .C(n), .Y(men_men_n597_));
  NA3        u0569(.A(men_men_n495_), .B(men_men_n177_), .C(men_men_n176_), .Y(men_men_n598_));
  NA2        u0570(.A(men_men_n441_), .B(men_men_n228_), .Y(men_men_n599_));
  OR2        u0571(.A(men_men_n599_), .B(men_men_n598_), .Y(men_men_n600_));
  NA2        u0572(.A(men_men_n76_), .B(men_men_n115_), .Y(men_men_n601_));
  NO2        u0573(.A(men_men_n601_), .B(men_men_n45_), .Y(men_men_n602_));
  AOI220     u0574(.A0(men_men_n602_), .A1(men_men_n524_), .B0(men_men_n600_), .B1(men_men_n597_), .Y(men_men_n603_));
  NO2        u0575(.A(men_men_n603_), .B(men_men_n89_), .Y(men_men_n604_));
  NA3        u0576(.A(men_men_n536_), .B(men_men_n333_), .C(men_men_n46_), .Y(men_men_n605_));
  NOi32      u0577(.An(e), .Bn(c), .C(f), .Y(men_men_n606_));
  NOi21      u0578(.An(f), .B(u), .Y(men_men_n607_));
  INV        u0579(.A(men_men_n212_), .Y(men_men_n608_));
  NA2        u0580(.A(men_men_n605_), .B(men_men_n182_), .Y(men_men_n609_));
  AOI210     u0581(.A0(men_men_n523_), .A1(men_men_n387_), .B0(men_men_n300_), .Y(men_men_n610_));
  NA2        u0582(.A(men_men_n610_), .B(men_men_n262_), .Y(men_men_n611_));
  NOi21      u0583(.An(j), .B(l), .Y(men_men_n612_));
  NAi21      u0584(.An(k), .B(h), .Y(men_men_n613_));
  NO2        u0585(.A(men_men_n613_), .B(men_men_n260_), .Y(men_men_n614_));
  NA2        u0586(.A(men_men_n614_), .B(men_men_n612_), .Y(men_men_n615_));
  OR2        u0587(.A(men_men_n615_), .B(men_men_n570_), .Y(men_men_n616_));
  NOi31      u0588(.An(m), .B(n), .C(k), .Y(men_men_n617_));
  NA2        u0589(.A(men_men_n612_), .B(men_men_n617_), .Y(men_men_n618_));
  NAi21      u0590(.An(men_men_n618_), .B(men_men_n386_), .Y(men_men_n619_));
  NO2        u0591(.A(men_men_n275_), .B(men_men_n49_), .Y(men_men_n620_));
  NO2        u0592(.A(men_men_n311_), .B(men_men_n580_), .Y(men_men_n621_));
  NO2        u0593(.A(men_men_n519_), .B(men_men_n49_), .Y(men_men_n622_));
  NA2        u0594(.A(men_men_n622_), .B(men_men_n621_), .Y(men_men_n623_));
  NA4        u0595(.A(men_men_n623_), .B(men_men_n619_), .C(men_men_n616_), .D(men_men_n611_), .Y(men_men_n624_));
  NA2        u0596(.A(men_men_n110_), .B(men_men_n36_), .Y(men_men_n625_));
  NO2        u0597(.A(k), .B(men_men_n215_), .Y(men_men_n626_));
  NO2        u0598(.A(men_men_n517_), .B(men_men_n180_), .Y(men_men_n627_));
  NA3        u0599(.A(men_men_n537_), .B(men_men_n269_), .C(men_men_n148_), .Y(men_men_n628_));
  NA2        u0600(.A(men_men_n491_), .B(men_men_n163_), .Y(men_men_n629_));
  NO3        u0601(.A(men_men_n385_), .B(men_men_n629_), .C(men_men_n89_), .Y(men_men_n630_));
  AOI210     u0602(.A0(men_men_n628_), .A1(men_men_n627_), .B0(men_men_n630_), .Y(men_men_n631_));
  AN3        u0603(.A(f), .B(d), .C(b), .Y(men_men_n632_));
  OAI210     u0604(.A0(men_men_n632_), .A1(men_men_n132_), .B0(n), .Y(men_men_n633_));
  NA3        u0605(.A(men_men_n491_), .B(men_men_n163_), .C(men_men_n215_), .Y(men_men_n634_));
  AOI210     u0606(.A0(men_men_n633_), .A1(men_men_n229_), .B0(men_men_n634_), .Y(men_men_n635_));
  NAi31      u0607(.An(m), .B(n), .C(k), .Y(men_men_n636_));
  OR2        u0608(.A(men_men_n137_), .B(men_men_n61_), .Y(men_men_n637_));
  OAI210     u0609(.A0(men_men_n637_), .A1(men_men_n636_), .B0(men_men_n247_), .Y(men_men_n638_));
  OAI210     u0610(.A0(men_men_n638_), .A1(men_men_n635_), .B0(j), .Y(men_men_n639_));
  NA2        u0611(.A(men_men_n639_), .B(men_men_n631_), .Y(men_men_n640_));
  NO4        u0612(.A(men_men_n640_), .B(men_men_n624_), .C(men_men_n609_), .D(men_men_n604_), .Y(men_men_n641_));
  NA2        u0613(.A(men_men_n377_), .B(men_men_n166_), .Y(men_men_n642_));
  NAi31      u0614(.An(u), .B(h), .C(f), .Y(men_men_n643_));
  OR3        u0615(.A(men_men_n643_), .B(men_men_n275_), .C(n), .Y(men_men_n644_));
  OA210      u0616(.A0(men_men_n519_), .A1(n), .B0(men_men_n568_), .Y(men_men_n645_));
  NA3        u0617(.A(men_men_n406_), .B(men_men_n122_), .C(men_men_n86_), .Y(men_men_n646_));
  OAI210     u0618(.A0(men_men_n645_), .A1(men_men_n93_), .B0(men_men_n646_), .Y(men_men_n647_));
  NOi21      u0619(.An(men_men_n644_), .B(men_men_n647_), .Y(men_men_n648_));
  AOI210     u0620(.A0(men_men_n648_), .A1(men_men_n642_), .B0(men_men_n512_), .Y(men_men_n649_));
  NAi21      u0621(.An(h), .B(j), .Y(men_men_n650_));
  INV        u0622(.A(men_men_n335_), .Y(men_men_n651_));
  OA220      u0623(.A0(men_men_n618_), .A1(men_men_n651_), .B0(men_men_n615_), .B1(men_men_n73_), .Y(men_men_n652_));
  NA3        u0624(.A(men_men_n509_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n653_));
  AN2        u0625(.A(h), .B(f), .Y(men_men_n654_));
  NA2        u0626(.A(men_men_n654_), .B(men_men_n37_), .Y(men_men_n655_));
  NA2        u0627(.A(men_men_n102_), .B(men_men_n46_), .Y(men_men_n656_));
  OAI220     u0628(.A0(men_men_n656_), .A1(men_men_n328_), .B0(men_men_n655_), .B1(men_men_n446_), .Y(men_men_n657_));
  AOI210     u0629(.A0(men_men_n551_), .A1(men_men_n416_), .B0(men_men_n49_), .Y(men_men_n658_));
  INV        u0630(.A(men_men_n657_), .Y(men_men_n659_));
  NA3        u0631(.A(men_men_n659_), .B(men_men_n653_), .C(men_men_n652_), .Y(men_men_n660_));
  NO2        u0632(.A(men_men_n249_), .B(f), .Y(men_men_n661_));
  INV        u0633(.A(men_men_n61_), .Y(men_men_n662_));
  NO2        u0634(.A(men_men_n662_), .B(men_men_n661_), .Y(men_men_n663_));
  NA2        u0635(.A(men_men_n326_), .B(men_men_n143_), .Y(men_men_n664_));
  NA2        u0636(.A(men_men_n134_), .B(men_men_n49_), .Y(men_men_n665_));
  AOI220     u0637(.A0(men_men_n665_), .A1(men_men_n515_), .B0(men_men_n356_), .B1(men_men_n115_), .Y(men_men_n666_));
  OA220      u0638(.A0(men_men_n666_), .A1(men_men_n535_), .B0(men_men_n354_), .B1(men_men_n113_), .Y(men_men_n667_));
  OAI210     u0639(.A0(men_men_n664_), .A1(men_men_n663_), .B0(men_men_n667_), .Y(men_men_n668_));
  NO3        u0640(.A(men_men_n393_), .B(men_men_n193_), .C(men_men_n192_), .Y(men_men_n669_));
  NA2        u0641(.A(men_men_n669_), .B(men_men_n228_), .Y(men_men_n670_));
  NA3        u0642(.A(men_men_n670_), .B(men_men_n251_), .C(j), .Y(men_men_n671_));
  NO3        u0643(.A(men_men_n441_), .B(men_men_n178_), .C(i), .Y(men_men_n672_));
  NA2        u0644(.A(men_men_n445_), .B(men_men_n86_), .Y(men_men_n673_));
  NO4        u0645(.A(men_men_n512_), .B(men_men_n673_), .C(men_men_n133_), .D(men_men_n214_), .Y(men_men_n674_));
  INV        u0646(.A(men_men_n674_), .Y(men_men_n675_));
  NA3        u0647(.A(men_men_n675_), .B(men_men_n671_), .C(men_men_n498_), .Y(men_men_n676_));
  NO4        u0648(.A(men_men_n676_), .B(men_men_n668_), .C(men_men_n660_), .D(men_men_n649_), .Y(men_men_n677_));
  NA4        u0649(.A(men_men_n677_), .B(men_men_n641_), .C(men_men_n596_), .D(men_men_n562_), .Y(men08));
  NO2        u0650(.A(k), .B(h), .Y(men_men_n679_));
  AO210      u0651(.A0(men_men_n249_), .A1(men_men_n435_), .B0(men_men_n679_), .Y(men_men_n680_));
  NO2        u0652(.A(men_men_n680_), .B(men_men_n298_), .Y(men_men_n681_));
  NA2        u0653(.A(men_men_n606_), .B(men_men_n86_), .Y(men_men_n682_));
  INV        u0654(.A(men_men_n475_), .Y(men_men_n683_));
  NA2        u0655(.A(men_men_n86_), .B(men_men_n112_), .Y(men_men_n684_));
  NO2        u0656(.A(men_men_n684_), .B(men_men_n57_), .Y(men_men_n685_));
  NO4        u0657(.A(men_men_n374_), .B(men_men_n114_), .C(j), .D(men_men_n215_), .Y(men_men_n686_));
  NA2        u0658(.A(men_men_n558_), .B(men_men_n229_), .Y(men_men_n687_));
  AOI220     u0659(.A0(men_men_n687_), .A1(men_men_n341_), .B0(men_men_n686_), .B1(men_men_n685_), .Y(men_men_n688_));
  AOI210     u0660(.A0(men_men_n558_), .A1(men_men_n159_), .B0(men_men_n86_), .Y(men_men_n689_));
  NA4        u0661(.A(men_men_n217_), .B(men_men_n143_), .C(men_men_n45_), .D(h), .Y(men_men_n690_));
  AN2        u0662(.A(l), .B(k), .Y(men_men_n691_));
  NA3        u0663(.A(men_men_n691_), .B(men_men_n110_), .C(men_men_n75_), .Y(men_men_n692_));
  OAI210     u0664(.A0(men_men_n690_), .A1(u), .B0(men_men_n692_), .Y(men_men_n693_));
  NA2        u0665(.A(men_men_n693_), .B(men_men_n689_), .Y(men_men_n694_));
  NA4        u0666(.A(men_men_n694_), .B(men_men_n688_), .C(men_men_n683_), .D(men_men_n343_), .Y(men_men_n695_));
  AN2        u0667(.A(men_men_n520_), .B(men_men_n98_), .Y(men_men_n696_));
  NO4        u0668(.A(men_men_n178_), .B(k), .C(men_men_n114_), .D(u), .Y(men_men_n697_));
  AOI210     u0669(.A0(men_men_n697_), .A1(men_men_n687_), .B0(men_men_n504_), .Y(men_men_n698_));
  NO2        u0670(.A(men_men_n38_), .B(men_men_n214_), .Y(men_men_n699_));
  NA2        u0671(.A(men_men_n699_), .B(men_men_n548_), .Y(men_men_n700_));
  NAi31      u0672(.An(men_men_n696_), .B(men_men_n700_), .C(men_men_n698_), .Y(men_men_n701_));
  NO2        u0673(.A(men_men_n523_), .B(men_men_n35_), .Y(men_men_n702_));
  OAI210     u0674(.A0(men_men_n537_), .A1(men_men_n47_), .B0(men_men_n637_), .Y(men_men_n703_));
  NO2        u0675(.A(men_men_n467_), .B(men_men_n134_), .Y(men_men_n704_));
  AOI210     u0676(.A0(men_men_n704_), .A1(men_men_n703_), .B0(men_men_n702_), .Y(men_men_n705_));
  NO3        u0677(.A(men_men_n317_), .B(men_men_n133_), .C(men_men_n41_), .Y(men_men_n706_));
  NAi21      u0678(.An(men_men_n706_), .B(men_men_n692_), .Y(men_men_n707_));
  NA2        u0679(.A(men_men_n680_), .B(men_men_n138_), .Y(men_men_n708_));
  AOI220     u0680(.A0(men_men_n708_), .A1(men_men_n392_), .B0(men_men_n707_), .B1(men_men_n78_), .Y(men_men_n709_));
  OAI210     u0681(.A0(men_men_n705_), .A1(men_men_n89_), .B0(men_men_n709_), .Y(men_men_n710_));
  NA2        u0682(.A(men_men_n356_), .B(men_men_n43_), .Y(men_men_n711_));
  NA3        u0683(.A(men_men_n670_), .B(men_men_n329_), .C(men_men_n380_), .Y(men_men_n712_));
  NA2        u0684(.A(men_men_n691_), .B(men_men_n222_), .Y(men_men_n713_));
  NO2        u0685(.A(men_men_n713_), .B(men_men_n325_), .Y(men_men_n714_));
  AOI210     u0686(.A0(men_men_n714_), .A1(men_men_n661_), .B0(men_men_n474_), .Y(men_men_n715_));
  NA3        u0687(.A(m), .B(l), .C(k), .Y(men_men_n716_));
  AOI210     u0688(.A0(men_men_n646_), .A1(men_men_n644_), .B0(men_men_n716_), .Y(men_men_n717_));
  NO2        u0689(.A(men_men_n522_), .B(men_men_n270_), .Y(men_men_n718_));
  NOi21      u0690(.An(men_men_n718_), .B(men_men_n516_), .Y(men_men_n719_));
  NA4        u0691(.A(men_men_n115_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n720_));
  NA3        u0692(.A(men_men_n122_), .B(men_men_n401_), .C(i), .Y(men_men_n721_));
  NO2        u0693(.A(men_men_n721_), .B(men_men_n720_), .Y(men_men_n722_));
  NO3        u0694(.A(men_men_n722_), .B(men_men_n719_), .C(men_men_n717_), .Y(men_men_n723_));
  NA4        u0695(.A(men_men_n723_), .B(men_men_n715_), .C(men_men_n712_), .D(men_men_n711_), .Y(men_men_n724_));
  NO4        u0696(.A(men_men_n724_), .B(men_men_n710_), .C(men_men_n701_), .D(men_men_n695_), .Y(men_men_n725_));
  NOi31      u0697(.An(u), .B(h), .C(f), .Y(men_men_n726_));
  NA2        u0698(.A(men_men_n622_), .B(men_men_n726_), .Y(men_men_n727_));
  AO210      u0699(.A0(men_men_n727_), .A1(men_men_n572_), .B0(men_men_n525_), .Y(men_men_n728_));
  NO3        u0700(.A(men_men_n387_), .B(men_men_n510_), .C(h), .Y(men_men_n729_));
  AOI210     u0701(.A0(men_men_n729_), .A1(men_men_n115_), .B0(men_men_n485_), .Y(men_men_n730_));
  NA3        u0702(.A(men_men_n730_), .B(men_men_n728_), .C(men_men_n248_), .Y(men_men_n731_));
  NA2        u0703(.A(men_men_n691_), .B(men_men_n75_), .Y(men_men_n732_));
  NO4        u0704(.A(men_men_n669_), .B(men_men_n178_), .C(n), .D(i), .Y(men_men_n733_));
  NOi21      u0705(.An(h), .B(j), .Y(men_men_n734_));
  NA2        u0706(.A(men_men_n734_), .B(f), .Y(men_men_n735_));
  NO2        u0707(.A(men_men_n735_), .B(men_men_n242_), .Y(men_men_n736_));
  NO3        u0708(.A(men_men_n736_), .B(men_men_n733_), .C(men_men_n672_), .Y(men_men_n737_));
  OAI220     u0709(.A0(men_men_n737_), .A1(men_men_n732_), .B0(men_men_n574_), .B1(men_men_n62_), .Y(men_men_n738_));
  AOI210     u0710(.A0(men_men_n731_), .A1(l), .B0(men_men_n738_), .Y(men_men_n739_));
  NO2        u0711(.A(j), .B(i), .Y(men_men_n740_));
  NA3        u0712(.A(men_men_n740_), .B(men_men_n82_), .C(l), .Y(men_men_n741_));
  NA2        u0713(.A(men_men_n740_), .B(men_men_n33_), .Y(men_men_n742_));
  NA2        u0714(.A(men_men_n410_), .B(men_men_n122_), .Y(men_men_n743_));
  OA220      u0715(.A0(men_men_n743_), .A1(men_men_n742_), .B0(men_men_n741_), .B1(men_men_n570_), .Y(men_men_n744_));
  NO3        u0716(.A(men_men_n154_), .B(men_men_n49_), .C(men_men_n112_), .Y(men_men_n745_));
  NO3        u0717(.A(c), .B(men_men_n153_), .C(men_men_n75_), .Y(men_men_n746_));
  NO3        u0718(.A(men_men_n467_), .B(men_men_n427_), .C(j), .Y(men_men_n747_));
  OAI210     u0719(.A0(men_men_n746_), .A1(men_men_n745_), .B0(men_men_n747_), .Y(men_men_n748_));
  OAI210     u0720(.A0(men_men_n727_), .A1(men_men_n62_), .B0(men_men_n748_), .Y(men_men_n749_));
  AOI210     u0721(.A0(men_men_n515_), .A1(n), .B0(men_men_n536_), .Y(men_men_n750_));
  NA2        u0722(.A(men_men_n750_), .B(men_men_n538_), .Y(men_men_n751_));
  NO3        u0723(.A(men_men_n178_), .B(k), .C(men_men_n114_), .Y(men_men_n752_));
  AOI220     u0724(.A0(men_men_n752_), .A1(men_men_n243_), .B0(men_men_n599_), .B1(men_men_n308_), .Y(men_men_n753_));
  NA2        u0725(.A(men_men_n95_), .B(men_men_n86_), .Y(men_men_n754_));
  NA2        u0726(.A(men_men_n754_), .B(men_men_n753_), .Y(men_men_n755_));
  NA2        u0727(.A(men_men_n706_), .B(men_men_n689_), .Y(men_men_n756_));
  NO2        u0728(.A(men_men_n716_), .B(men_men_n93_), .Y(men_men_n757_));
  NA2        u0729(.A(men_men_n757_), .B(men_men_n569_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n758_), .B(men_men_n756_), .Y(men_men_n759_));
  OR3        u0731(.A(men_men_n759_), .B(men_men_n755_), .C(men_men_n749_), .Y(men_men_n760_));
  NO4        u0732(.A(men_men_n467_), .B(men_men_n423_), .C(j), .D(f), .Y(men_men_n761_));
  OAI220     u0733(.A0(men_men_n690_), .A1(men_men_n682_), .B0(men_men_n328_), .B1(men_men_n38_), .Y(men_men_n762_));
  AOI210     u0734(.A0(men_men_n761_), .A1(men_men_n255_), .B0(men_men_n762_), .Y(men_men_n763_));
  NA3        u0735(.A(men_men_n531_), .B(men_men_n291_), .C(h), .Y(men_men_n764_));
  NOi21      u0736(.An(men_men_n658_), .B(men_men_n764_), .Y(men_men_n765_));
  OAI220     u0737(.A0(men_men_n764_), .A1(men_men_n588_), .B0(men_men_n741_), .B1(men_men_n73_), .Y(men_men_n766_));
  INV        u0738(.A(men_men_n766_), .Y(men_men_n767_));
  NAi31      u0739(.An(men_men_n765_), .B(men_men_n767_), .C(men_men_n763_), .Y(men_men_n768_));
  OR2        u0740(.A(men_men_n757_), .B(men_men_n98_), .Y(men_men_n769_));
  AOI220     u0741(.A0(men_men_n769_), .A1(men_men_n235_), .B0(men_men_n747_), .B1(men_men_n620_), .Y(men_men_n770_));
  NO2        u0742(.A(men_men_n645_), .B(men_men_n75_), .Y(men_men_n771_));
  NA2        u0743(.A(men_men_n761_), .B(men_men_n771_), .Y(men_men_n772_));
  OAI210     u0744(.A0(men_men_n716_), .A1(men_men_n643_), .B0(men_men_n503_), .Y(men_men_n773_));
  NA3        u0745(.A(men_men_n246_), .B(men_men_n59_), .C(b), .Y(men_men_n774_));
  AOI220     u0746(.A0(men_men_n587_), .A1(men_men_n29_), .B0(men_men_n445_), .B1(men_men_n86_), .Y(men_men_n775_));
  NA2        u0747(.A(men_men_n775_), .B(men_men_n774_), .Y(men_men_n776_));
  NO2        u0748(.A(men_men_n764_), .B(men_men_n473_), .Y(men_men_n777_));
  AOI210     u0749(.A0(men_men_n776_), .A1(men_men_n773_), .B0(men_men_n777_), .Y(men_men_n778_));
  NA3        u0750(.A(men_men_n778_), .B(men_men_n772_), .C(men_men_n770_), .Y(men_men_n779_));
  NOi41      u0751(.An(men_men_n744_), .B(men_men_n779_), .C(men_men_n768_), .D(men_men_n760_), .Y(men_men_n780_));
  OR3        u0752(.A(men_men_n690_), .B(men_men_n229_), .C(u), .Y(men_men_n781_));
  NO3        u0753(.A(men_men_n334_), .B(men_men_n300_), .C(men_men_n114_), .Y(men_men_n782_));
  NA2        u0754(.A(men_men_n782_), .B(men_men_n751_), .Y(men_men_n783_));
  NA2        u0755(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n784_));
  NO3        u0756(.A(men_men_n784_), .B(men_men_n742_), .C(men_men_n275_), .Y(men_men_n785_));
  INV        u0757(.A(men_men_n785_), .Y(men_men_n786_));
  NA4        u0758(.A(men_men_n786_), .B(men_men_n783_), .C(men_men_n781_), .D(men_men_n394_), .Y(men_men_n787_));
  OR2        u0759(.A(men_men_n643_), .B(men_men_n94_), .Y(men_men_n788_));
  NOi31      u0760(.An(b), .B(d), .C(a), .Y(men_men_n789_));
  NO2        u0761(.A(men_men_n789_), .B(men_men_n585_), .Y(men_men_n790_));
  NO2        u0762(.A(men_men_n790_), .B(n), .Y(men_men_n791_));
  NOi21      u0763(.An(men_men_n775_), .B(men_men_n791_), .Y(men_men_n792_));
  OAI220     u0764(.A0(men_men_n792_), .A1(men_men_n788_), .B0(men_men_n764_), .B1(men_men_n586_), .Y(men_men_n793_));
  INV        u0765(.A(men_men_n537_), .Y(men_men_n794_));
  NO2        u0766(.A(men_men_n325_), .B(men_men_n118_), .Y(men_men_n795_));
  NOi21      u0767(.An(men_men_n795_), .B(men_men_n164_), .Y(men_men_n796_));
  AOI210     u0768(.A0(men_men_n782_), .A1(men_men_n794_), .B0(men_men_n796_), .Y(men_men_n797_));
  INV        u0769(.A(men_men_n797_), .Y(men_men_n798_));
  NA2        u0770(.A(men_men_n192_), .B(men_men_n681_), .Y(men_men_n799_));
  NO2        u0771(.A(men_men_n322_), .B(men_men_n234_), .Y(men_men_n800_));
  OAI210     u0772(.A0(men_men_n98_), .A1(men_men_n95_), .B0(men_men_n800_), .Y(men_men_n801_));
  NA2        u0773(.A(men_men_n122_), .B(men_men_n86_), .Y(men_men_n802_));
  AOI210     u0774(.A0(men_men_n413_), .A1(men_men_n407_), .B0(men_men_n802_), .Y(men_men_n803_));
  NAi21      u0775(.An(men_men_n803_), .B(men_men_n801_), .Y(men_men_n804_));
  NA2        u0776(.A(men_men_n714_), .B(men_men_n34_), .Y(men_men_n805_));
  NAi21      u0777(.An(men_men_n720_), .B(men_men_n424_), .Y(men_men_n806_));
  NA2        u0778(.A(men_men_n697_), .B(men_men_n342_), .Y(men_men_n807_));
  OAI210     u0779(.A0(men_men_n577_), .A1(men_men_n576_), .B0(men_men_n357_), .Y(men_men_n808_));
  AN3        u0780(.A(men_men_n808_), .B(men_men_n807_), .C(men_men_n806_), .Y(men_men_n809_));
  NAi41      u0781(.An(men_men_n804_), .B(men_men_n809_), .C(men_men_n805_), .D(men_men_n799_), .Y(men_men_n810_));
  NO4        u0782(.A(men_men_n810_), .B(men_men_n798_), .C(men_men_n793_), .D(men_men_n787_), .Y(men_men_n811_));
  NA4        u0783(.A(men_men_n811_), .B(men_men_n780_), .C(men_men_n739_), .D(men_men_n725_), .Y(men09));
  INV        u0784(.A(men_men_n123_), .Y(men_men_n813_));
  NA2        u0785(.A(f), .B(e), .Y(men_men_n814_));
  NO2        u0786(.A(men_men_n226_), .B(men_men_n114_), .Y(men_men_n815_));
  NA2        u0787(.A(men_men_n815_), .B(u), .Y(men_men_n816_));
  NA4        u0788(.A(men_men_n311_), .B(men_men_n454_), .C(men_men_n258_), .D(men_men_n120_), .Y(men_men_n817_));
  AOI210     u0789(.A0(men_men_n817_), .A1(u), .B0(men_men_n451_), .Y(men_men_n818_));
  AOI210     u0790(.A0(men_men_n818_), .A1(men_men_n816_), .B0(men_men_n814_), .Y(men_men_n819_));
  NA2        u0791(.A(men_men_n819_), .B(men_men_n813_), .Y(men_men_n820_));
  NO2        u0792(.A(men_men_n204_), .B(men_men_n214_), .Y(men_men_n821_));
  NA3        u0793(.A(m), .B(l), .C(i), .Y(men_men_n822_));
  NA4        u0794(.A(men_men_n90_), .B(men_men_n89_), .C(u), .D(f), .Y(men_men_n823_));
  NA2        u0795(.A(men_men_n823_), .B(men_men_n428_), .Y(men_men_n824_));
  OR2        u0796(.A(men_men_n824_), .B(men_men_n821_), .Y(men_men_n825_));
  NA3        u0797(.A(men_men_n788_), .B(men_men_n550_), .C(men_men_n503_), .Y(men_men_n826_));
  OA210      u0798(.A0(men_men_n826_), .A1(men_men_n825_), .B0(men_men_n791_), .Y(men_men_n827_));
  INV        u0799(.A(men_men_n331_), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n129_), .B(men_men_n127_), .Y(men_men_n829_));
  NO2        u0801(.A(m), .B(men_men_n580_), .Y(men_men_n830_));
  NA2        u0802(.A(men_men_n335_), .B(men_men_n337_), .Y(men_men_n831_));
  OAI210     u0803(.A0(men_men_n204_), .A1(men_men_n214_), .B0(men_men_n831_), .Y(men_men_n832_));
  AOI220     u0804(.A0(men_men_n832_), .A1(men_men_n246_), .B0(men_men_n830_), .B1(men_men_n828_), .Y(men_men_n833_));
  NA2        u0805(.A(men_men_n173_), .B(k), .Y(men_men_n834_));
  NA3        u0806(.A(men_men_n834_), .B(men_men_n680_), .C(men_men_n138_), .Y(men_men_n835_));
  NA3        u0807(.A(men_men_n835_), .B(men_men_n191_), .C(men_men_n31_), .Y(men_men_n836_));
  NA3        u0808(.A(men_men_n836_), .B(men_men_n833_), .C(men_men_n84_), .Y(men_men_n837_));
  NO2        u0809(.A(men_men_n567_), .B(men_men_n481_), .Y(men_men_n838_));
  NA2        u0810(.A(men_men_n838_), .B(men_men_n191_), .Y(men_men_n839_));
  NOi21      u0811(.An(f), .B(d), .Y(men_men_n840_));
  NA2        u0812(.A(men_men_n840_), .B(m), .Y(men_men_n841_));
  NO2        u0813(.A(men_men_n841_), .B(men_men_n52_), .Y(men_men_n842_));
  NOi32      u0814(.An(u), .Bn(f), .C(d), .Y(men_men_n843_));
  NA4        u0815(.A(men_men_n843_), .B(men_men_n587_), .C(men_men_n29_), .D(m), .Y(men_men_n844_));
  NOi21      u0816(.An(men_men_n312_), .B(men_men_n844_), .Y(men_men_n845_));
  INV        u0817(.A(men_men_n845_), .Y(men_men_n846_));
  NA2        u0818(.A(men_men_n311_), .B(men_men_n258_), .Y(men_men_n847_));
  AN2        u0819(.A(f), .B(d), .Y(men_men_n848_));
  NA3        u0820(.A(men_men_n459_), .B(men_men_n848_), .C(men_men_n86_), .Y(men_men_n849_));
  NO3        u0821(.A(men_men_n849_), .B(men_men_n75_), .C(men_men_n215_), .Y(men_men_n850_));
  NA2        u0822(.A(men_men_n847_), .B(men_men_n850_), .Y(men_men_n851_));
  NAi41      u0823(.An(men_men_n472_), .B(men_men_n851_), .C(men_men_n846_), .D(men_men_n839_), .Y(men_men_n852_));
  NO4        u0824(.A(men_men_n607_), .B(men_men_n134_), .C(men_men_n325_), .D(men_men_n155_), .Y(men_men_n853_));
  NO2        u0825(.A(men_men_n636_), .B(men_men_n325_), .Y(men_men_n854_));
  AN2        u0826(.A(men_men_n854_), .B(men_men_n661_), .Y(men_men_n855_));
  NO3        u0827(.A(men_men_n855_), .B(men_men_n853_), .C(men_men_n231_), .Y(men_men_n856_));
  NA2        u0828(.A(men_men_n585_), .B(men_men_n86_), .Y(men_men_n857_));
  NO2        u0829(.A(men_men_n831_), .B(men_men_n857_), .Y(men_men_n858_));
  NOi21      u0830(.An(men_men_n224_), .B(men_men_n858_), .Y(men_men_n859_));
  NA2        u0831(.A(c), .B(men_men_n117_), .Y(men_men_n860_));
  NO2        u0832(.A(men_men_n860_), .B(men_men_n398_), .Y(men_men_n861_));
  NA3        u0833(.A(men_men_n861_), .B(men_men_n493_), .C(f), .Y(men_men_n862_));
  OR2        u0834(.A(men_men_n643_), .B(men_men_n526_), .Y(men_men_n863_));
  INV        u0835(.A(men_men_n863_), .Y(men_men_n864_));
  NA2        u0836(.A(men_men_n790_), .B(men_men_n113_), .Y(men_men_n865_));
  NA2        u0837(.A(men_men_n865_), .B(men_men_n864_), .Y(men_men_n866_));
  NA4        u0838(.A(men_men_n866_), .B(men_men_n862_), .C(men_men_n859_), .D(men_men_n856_), .Y(men_men_n867_));
  NO4        u0839(.A(men_men_n867_), .B(men_men_n852_), .C(men_men_n837_), .D(men_men_n827_), .Y(men_men_n868_));
  OR2        u0840(.A(men_men_n849_), .B(men_men_n75_), .Y(men_men_n869_));
  INV        u0841(.A(men_men_n815_), .Y(men_men_n870_));
  AOI210     u0842(.A0(men_men_n870_), .A1(men_men_n292_), .B0(men_men_n869_), .Y(men_men_n871_));
  NO2        u0843(.A(men_men_n328_), .B(men_men_n823_), .Y(men_men_n872_));
  NO2        u0844(.A(men_men_n138_), .B(men_men_n134_), .Y(men_men_n873_));
  NO2        u0845(.A(men_men_n228_), .B(men_men_n225_), .Y(men_men_n874_));
  AOI220     u0846(.A0(men_men_n874_), .A1(men_men_n227_), .B0(men_men_n305_), .B1(men_men_n873_), .Y(men_men_n875_));
  NO2        u0847(.A(men_men_n418_), .B(men_men_n814_), .Y(men_men_n876_));
  NA2        u0848(.A(men_men_n876_), .B(men_men_n542_), .Y(men_men_n877_));
  NA2        u0849(.A(men_men_n877_), .B(men_men_n875_), .Y(men_men_n878_));
  NA2        u0850(.A(e), .B(d), .Y(men_men_n879_));
  OAI220     u0851(.A0(men_men_n879_), .A1(c), .B0(men_men_n322_), .B1(d), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n608_), .B(men_men_n340_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n284_), .B(men_men_n169_), .Y(men_men_n882_));
  NA2        u0854(.A(men_men_n850_), .B(men_men_n882_), .Y(men_men_n883_));
  NA2        u0855(.A(men_men_n883_), .B(men_men_n881_), .Y(men_men_n884_));
  NO4        u0856(.A(men_men_n884_), .B(men_men_n878_), .C(men_men_n872_), .D(men_men_n871_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n828_), .B(men_men_n31_), .Y(men_men_n886_));
  AO210      u0858(.A0(men_men_n886_), .A1(men_men_n682_), .B0(men_men_n218_), .Y(men_men_n887_));
  OAI220     u0859(.A0(men_men_n607_), .A1(men_men_n61_), .B0(men_men_n300_), .B1(j), .Y(men_men_n888_));
  AOI220     u0860(.A0(men_men_n888_), .A1(men_men_n854_), .B0(men_men_n597_), .B1(men_men_n606_), .Y(men_men_n889_));
  INV        u0861(.A(men_men_n889_), .Y(men_men_n890_));
  OAI210     u0862(.A0(men_men_n815_), .A1(men_men_n882_), .B0(men_men_n843_), .Y(men_men_n891_));
  NO2        u0863(.A(men_men_n891_), .B(men_men_n588_), .Y(men_men_n892_));
  AOI210     u0864(.A0(men_men_n119_), .A1(men_men_n118_), .B0(men_men_n257_), .Y(men_men_n893_));
  NO2        u0865(.A(men_men_n893_), .B(men_men_n844_), .Y(men_men_n894_));
  NOi31      u0866(.An(men_men_n529_), .B(men_men_n841_), .C(men_men_n292_), .Y(men_men_n895_));
  NO4        u0867(.A(men_men_n895_), .B(men_men_n894_), .C(men_men_n892_), .D(men_men_n890_), .Y(men_men_n896_));
  BUFFER     u0868(.A(men_men_n438_), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n897_), .B(men_men_n880_), .Y(men_men_n898_));
  NO2        u0870(.A(men_men_n427_), .B(men_men_n71_), .Y(men_men_n899_));
  OAI210     u0871(.A0(men_men_n826_), .A1(men_men_n899_), .B0(men_men_n685_), .Y(men_men_n900_));
  AN4        u0872(.A(men_men_n900_), .B(men_men_n898_), .C(men_men_n896_), .D(men_men_n887_), .Y(men_men_n901_));
  NA4        u0873(.A(men_men_n901_), .B(men_men_n885_), .C(men_men_n868_), .D(men_men_n820_), .Y(men12));
  NO4        u0874(.A(men_men_n432_), .B(men_men_n249_), .C(men_men_n563_), .D(men_men_n215_), .Y(men_men_n903_));
  NA2        u0875(.A(men_men_n529_), .B(men_men_n899_), .Y(men_men_n904_));
  NO2        u0876(.A(men_men_n437_), .B(men_men_n117_), .Y(men_men_n905_));
  NO2        u0877(.A(men_men_n829_), .B(men_men_n347_), .Y(men_men_n906_));
  NO2        u0878(.A(men_men_n643_), .B(men_men_n374_), .Y(men_men_n907_));
  AOI220     u0879(.A0(men_men_n907_), .A1(men_men_n528_), .B0(men_men_n906_), .B1(men_men_n905_), .Y(men_men_n908_));
  NA3        u0880(.A(men_men_n908_), .B(men_men_n904_), .C(men_men_n431_), .Y(men_men_n909_));
  AOI210     u0881(.A0(men_men_n230_), .A1(men_men_n330_), .B0(men_men_n201_), .Y(men_men_n910_));
  OR2        u0882(.A(men_men_n910_), .B(men_men_n903_), .Y(men_men_n911_));
  NA2        u0883(.A(men_men_n911_), .B(men_men_n393_), .Y(men_men_n912_));
  NO2        u0884(.A(men_men_n625_), .B(men_men_n260_), .Y(men_men_n913_));
  NO2        u0885(.A(men_men_n571_), .B(men_men_n822_), .Y(men_men_n914_));
  AOI220     u0886(.A0(men_men_n914_), .A1(men_men_n548_), .B0(men_men_n800_), .B1(men_men_n913_), .Y(men_men_n915_));
  NO2        u0887(.A(men_men_n154_), .B(men_men_n234_), .Y(men_men_n916_));
  NA3        u0888(.A(men_men_n916_), .B(men_men_n237_), .C(i), .Y(men_men_n917_));
  NA3        u0889(.A(men_men_n917_), .B(men_men_n915_), .C(men_men_n912_), .Y(men_men_n918_));
  OR2        u0890(.A(men_men_n323_), .B(men_men_n905_), .Y(men_men_n919_));
  NA2        u0891(.A(men_men_n919_), .B(men_men_n348_), .Y(men_men_n920_));
  NO3        u0892(.A(men_men_n134_), .B(men_men_n155_), .C(men_men_n215_), .Y(men_men_n921_));
  NA2        u0893(.A(men_men_n921_), .B(men_men_n515_), .Y(men_men_n922_));
  NA2        u0894(.A(men_men_n922_), .B(men_men_n920_), .Y(men_men_n923_));
  NO2        u0895(.A(men_men_n648_), .B(men_men_n45_), .Y(men_men_n924_));
  NO4        u0896(.A(men_men_n924_), .B(men_men_n923_), .C(men_men_n918_), .D(men_men_n909_), .Y(men_men_n925_));
  NO2        u0897(.A(men_men_n364_), .B(men_men_n363_), .Y(men_men_n926_));
  NA2        u0898(.A(men_men_n568_), .B(men_men_n73_), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n537_), .B(men_men_n148_), .Y(men_men_n928_));
  NOi21      u0900(.An(men_men_n34_), .B(men_men_n636_), .Y(men_men_n929_));
  AOI220     u0901(.A0(men_men_n929_), .A1(men_men_n928_), .B0(men_men_n927_), .B1(men_men_n926_), .Y(men_men_n930_));
  OAI210     u0902(.A0(men_men_n247_), .A1(men_men_n45_), .B0(men_men_n930_), .Y(men_men_n931_));
  NA2        u0903(.A(men_men_n424_), .B(men_men_n262_), .Y(men_men_n932_));
  NO3        u0904(.A(men_men_n802_), .B(men_men_n91_), .C(men_men_n398_), .Y(men_men_n933_));
  NAi21      u0905(.An(men_men_n933_), .B(men_men_n932_), .Y(men_men_n934_));
  NO2        u0906(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n935_));
  NO2        u0907(.A(men_men_n488_), .B(men_men_n300_), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n617_), .B(men_men_n357_), .Y(men_men_n937_));
  INV        u0909(.A(men_men_n361_), .Y(men_men_n938_));
  NO3        u0910(.A(men_men_n938_), .B(men_men_n934_), .C(men_men_n931_), .Y(men_men_n939_));
  NA2        u0911(.A(men_men_n340_), .B(u), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n166_), .B(i), .Y(men_men_n941_));
  NA2        u0913(.A(men_men_n46_), .B(i), .Y(men_men_n942_));
  OAI220     u0914(.A0(men_men_n942_), .A1(men_men_n200_), .B0(men_men_n941_), .B1(men_men_n94_), .Y(men_men_n943_));
  INV        u0915(.A(men_men_n943_), .Y(men_men_n944_));
  NO2        u0916(.A(men_men_n148_), .B(men_men_n86_), .Y(men_men_n945_));
  BUFFER     u0917(.A(men_men_n945_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n537_), .B(men_men_n378_), .Y(men_men_n947_));
  AOI210     u0919(.A0(men_men_n947_), .A1(n), .B0(men_men_n946_), .Y(men_men_n948_));
  OAI220     u0920(.A0(men_men_n948_), .A1(men_men_n940_), .B0(men_men_n944_), .B1(men_men_n328_), .Y(men_men_n949_));
  NO2        u0921(.A(men_men_n643_), .B(men_men_n481_), .Y(men_men_n950_));
  NA3        u0922(.A(men_men_n335_), .B(men_men_n612_), .C(i), .Y(men_men_n951_));
  OAI210     u0923(.A0(men_men_n427_), .A1(men_men_n311_), .B0(men_men_n951_), .Y(men_men_n952_));
  OAI220     u0924(.A0(men_men_n952_), .A1(men_men_n950_), .B0(men_men_n658_), .B1(men_men_n746_), .Y(men_men_n953_));
  NA2        u0925(.A(men_men_n591_), .B(men_men_n115_), .Y(men_men_n954_));
  OR3        u0926(.A(men_men_n311_), .B(men_men_n423_), .C(f), .Y(men_men_n955_));
  NA3        u0927(.A(men_men_n612_), .B(men_men_n82_), .C(i), .Y(men_men_n956_));
  OA220      u0928(.A0(men_men_n956_), .A1(men_men_n954_), .B0(men_men_n955_), .B1(men_men_n570_), .Y(men_men_n957_));
  NA3        u0929(.A(men_men_n324_), .B(men_men_n119_), .C(u), .Y(men_men_n958_));
  AOI210     u0930(.A0(men_men_n655_), .A1(men_men_n958_), .B0(m), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n959_), .A1(men_men_n906_), .B0(men_men_n323_), .Y(men_men_n960_));
  NA2        u0932(.A(men_men_n673_), .B(men_men_n857_), .Y(men_men_n961_));
  NA2        u0933(.A(men_men_n823_), .B(men_men_n428_), .Y(men_men_n962_));
  NA2        u0934(.A(i), .B(men_men_n79_), .Y(men_men_n963_));
  NA3        u0935(.A(men_men_n963_), .B(men_men_n956_), .C(men_men_n955_), .Y(men_men_n964_));
  AOI220     u0936(.A0(men_men_n964_), .A1(men_men_n255_), .B0(men_men_n962_), .B1(men_men_n961_), .Y(men_men_n965_));
  NA4        u0937(.A(men_men_n965_), .B(men_men_n960_), .C(men_men_n957_), .D(men_men_n953_), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n913_), .B(men_men_n235_), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n647_), .B(men_men_n90_), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n440_), .B(men_men_n215_), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n919_), .B(men_men_n219_), .Y(men_men_n970_));
  AOI220     u0942(.A0(men_men_n907_), .A1(men_men_n916_), .B0(men_men_n569_), .B1(men_men_n92_), .Y(men_men_n971_));
  NA4        u0943(.A(men_men_n971_), .B(men_men_n970_), .C(men_men_n968_), .D(men_men_n967_), .Y(men_men_n972_));
  OAI210     u0944(.A0(men_men_n962_), .A1(men_men_n914_), .B0(men_men_n528_), .Y(men_men_n973_));
  NO2        u0945(.A(men_men_n402_), .B(men_men_n802_), .Y(men_men_n974_));
  OAI210     u0946(.A0(men_men_n364_), .A1(men_men_n363_), .B0(men_men_n111_), .Y(men_men_n975_));
  AOI210     u0947(.A0(men_men_n975_), .A1(men_men_n520_), .B0(men_men_n974_), .Y(men_men_n976_));
  NA2        u0948(.A(men_men_n959_), .B(men_men_n905_), .Y(men_men_n977_));
  NO3        u0949(.A(l), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n978_));
  AOI220     u0950(.A0(men_men_n978_), .A1(men_men_n610_), .B0(men_men_n627_), .B1(men_men_n515_), .Y(men_men_n979_));
  NA4        u0951(.A(men_men_n979_), .B(men_men_n977_), .C(men_men_n976_), .D(men_men_n973_), .Y(men_men_n980_));
  NO4        u0952(.A(men_men_n980_), .B(men_men_n972_), .C(men_men_n966_), .D(men_men_n949_), .Y(men_men_n981_));
  NAi31      u0953(.An(men_men_n144_), .B(men_men_n410_), .C(n), .Y(men_men_n982_));
  NO3        u0954(.A(men_men_n127_), .B(men_men_n333_), .C(k), .Y(men_men_n983_));
  NA2        u0955(.A(men_men_n475_), .B(i), .Y(men_men_n984_));
  NA2        u0956(.A(men_men_n984_), .B(men_men_n982_), .Y(men_men_n985_));
  NA2        u0957(.A(men_men_n228_), .B(men_men_n177_), .Y(men_men_n986_));
  NAi21      u0958(.An(men_men_n537_), .B(men_men_n969_), .Y(men_men_n987_));
  NO3        u0959(.A(men_men_n427_), .B(men_men_n311_), .C(men_men_n75_), .Y(men_men_n988_));
  AOI220     u0960(.A0(men_men_n988_), .A1(a), .B0(men_men_n465_), .B1(u), .Y(men_men_n989_));
  NA2        u0961(.A(men_men_n989_), .B(men_men_n987_), .Y(men_men_n990_));
  NO2        u0962(.A(men_men_n951_), .B(men_men_n586_), .Y(men_men_n991_));
  NO3        u0963(.A(c), .B(men_men_n153_), .C(men_men_n214_), .Y(men_men_n992_));
  OAI210     u0964(.A0(men_men_n992_), .A1(men_men_n509_), .B0(men_men_n375_), .Y(men_men_n993_));
  OAI220     u0965(.A0(men_men_n907_), .A1(men_men_n914_), .B0(men_men_n529_), .B1(men_men_n417_), .Y(men_men_n994_));
  NA3        u0966(.A(men_men_n994_), .B(men_men_n993_), .C(men_men_n605_), .Y(men_men_n995_));
  OAI210     u0967(.A0(men_men_n910_), .A1(men_men_n903_), .B0(men_men_n986_), .Y(men_men_n996_));
  NA3        u0968(.A(men_men_n947_), .B(men_men_n469_), .C(men_men_n46_), .Y(men_men_n997_));
  AOI210     u0969(.A0(men_men_n377_), .A1(men_men_n375_), .B0(men_men_n327_), .Y(men_men_n998_));
  NA4        u0970(.A(men_men_n998_), .B(men_men_n997_), .C(men_men_n996_), .D(men_men_n271_), .Y(men_men_n999_));
  OR3        u0971(.A(men_men_n999_), .B(men_men_n995_), .C(men_men_n991_), .Y(men_men_n1000_));
  NO3        u0972(.A(men_men_n1000_), .B(men_men_n990_), .C(men_men_n985_), .Y(men_men_n1001_));
  NA4        u0973(.A(men_men_n1001_), .B(men_men_n981_), .C(men_men_n939_), .D(men_men_n925_), .Y(men13));
  NA2        u0974(.A(men_men_n46_), .B(men_men_n89_), .Y(men_men_n1003_));
  NA3        u0975(.A(men_men_n246_), .B(c), .C(m), .Y(men_men_n1004_));
  NO3        u0976(.A(men_men_n1004_), .B(men_men_n1003_), .C(men_men_n564_), .Y(men_men_n1005_));
  NA2        u0977(.A(men_men_n262_), .B(c), .Y(men_men_n1006_));
  NO4        u0978(.A(men_men_n1006_), .B(e), .C(men_men_n941_), .D(a), .Y(men_men_n1007_));
  NA2        u0979(.A(men_men_n143_), .B(men_men_n45_), .Y(men_men_n1008_));
  NO4        u0980(.A(men_men_n1008_), .B(c), .C(men_men_n571_), .D(men_men_n307_), .Y(men_men_n1009_));
  NA2        u0981(.A(men_men_n650_), .B(men_men_n225_), .Y(men_men_n1010_));
  NA2        u0982(.A(men_men_n401_), .B(men_men_n214_), .Y(men_men_n1011_));
  AN2        u0983(.A(d), .B(c), .Y(men_men_n1012_));
  NA2        u0984(.A(men_men_n1012_), .B(men_men_n117_), .Y(men_men_n1013_));
  NO3        u0985(.A(men_men_n1013_), .B(men_men_n1011_), .C(men_men_n180_), .Y(men_men_n1014_));
  NA2        u0986(.A(d), .B(c), .Y(men_men_n1015_));
  NO4        u0987(.A(men_men_n1008_), .B(men_men_n567_), .C(men_men_n1015_), .D(men_men_n307_), .Y(men_men_n1016_));
  AO210      u0988(.A0(men_men_n1014_), .A1(men_men_n1010_), .B0(men_men_n1016_), .Y(men_men_n1017_));
  OR4        u0989(.A(men_men_n1017_), .B(men_men_n1009_), .C(men_men_n1007_), .D(men_men_n1005_), .Y(men_men_n1018_));
  NAi32      u0990(.An(f), .Bn(e), .C(c), .Y(men_men_n1019_));
  NO2        u0991(.A(men_men_n1019_), .B(men_men_n150_), .Y(men_men_n1020_));
  NA2        u0992(.A(men_men_n1020_), .B(u), .Y(men_men_n1021_));
  OR2        u0993(.A(men_men_n225_), .B(men_men_n180_), .Y(men_men_n1022_));
  NO2        u0994(.A(men_men_n1022_), .B(men_men_n1021_), .Y(men_men_n1023_));
  NO2        u0995(.A(men_men_n1015_), .B(men_men_n307_), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n614_), .B(i), .Y(men_men_n1025_));
  NOi21      u0997(.An(men_men_n1024_), .B(men_men_n1025_), .Y(men_men_n1026_));
  NOi41      u0998(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1027_));
  NA2        u0999(.A(men_men_n1027_), .B(l), .Y(men_men_n1028_));
  NO2        u1000(.A(men_men_n1028_), .B(men_men_n1021_), .Y(men_men_n1029_));
  OR3        u1001(.A(e), .B(d), .C(c), .Y(men_men_n1030_));
  NA3        u1002(.A(k), .B(j), .C(i), .Y(men_men_n1031_));
  NO3        u1003(.A(men_men_n1031_), .B(men_men_n307_), .C(men_men_n93_), .Y(men_men_n1032_));
  BUFFER     u1004(.A(men_men_n1032_), .Y(men_men_n1033_));
  OR4        u1005(.A(men_men_n1033_), .B(men_men_n1029_), .C(men_men_n1026_), .D(men_men_n1023_), .Y(men_men_n1034_));
  NA2        u1006(.A(men_men_n448_), .B(men_men_n329_), .Y(men_men_n1035_));
  NO2        u1007(.A(men_men_n1035_), .B(men_men_n1025_), .Y(men_men_n1036_));
  NO4        u1008(.A(men_men_n1035_), .B(men_men_n567_), .C(men_men_n435_), .D(men_men_n45_), .Y(men_men_n1037_));
  NO2        u1009(.A(f), .B(c), .Y(men_men_n1038_));
  NOi21      u1010(.An(men_men_n1038_), .B(men_men_n432_), .Y(men_men_n1039_));
  NA2        u1011(.A(men_men_n1039_), .B(men_men_n59_), .Y(men_men_n1040_));
  NOi21      u1012(.An(men_men_n1450_), .B(men_men_n1040_), .Y(men_men_n1041_));
  OR3        u1013(.A(men_men_n1041_), .B(men_men_n1037_), .C(men_men_n1036_), .Y(men_men_n1042_));
  OR3        u1014(.A(men_men_n1042_), .B(men_men_n1034_), .C(men_men_n1018_), .Y(men02));
  OR3        u1015(.A(h), .B(u), .C(f), .Y(men_men_n1044_));
  NO4        u1016(.A(m), .B(men_men_n1044_), .C(l), .D(men_men_n1030_), .Y(men_men_n1045_));
  NO2        u1017(.A(men_men_n1032_), .B(men_men_n1009_), .Y(men_men_n1046_));
  OR2        u1018(.A(men_men_n1031_), .B(men_men_n307_), .Y(men_men_n1047_));
  OR2        u1019(.A(men_men_n1047_), .B(men_men_n1451_), .Y(men_men_n1048_));
  NO3        u1020(.A(men_men_n1035_), .B(men_men_n1008_), .C(men_men_n567_), .Y(men_men_n1049_));
  NO2        u1021(.A(men_men_n1049_), .B(men_men_n1023_), .Y(men_men_n1050_));
  NA2        u1022(.A(i), .B(h), .Y(men_men_n1051_));
  NO2        u1023(.A(men_men_n1051_), .B(men_men_n134_), .Y(men_men_n1052_));
  NO3        u1024(.A(men_men_n145_), .B(men_men_n282_), .C(men_men_n215_), .Y(men_men_n1053_));
  AOI210     u1025(.A0(men_men_n1053_), .A1(men_men_n1052_), .B0(men_men_n1026_), .Y(men_men_n1054_));
  NA3        u1026(.A(c), .B(b), .C(a), .Y(men_men_n1055_));
  NO3        u1027(.A(men_men_n1055_), .B(men_men_n879_), .C(men_men_n214_), .Y(men_men_n1056_));
  NO3        u1028(.A(men_men_n300_), .B(men_men_n49_), .C(men_men_n114_), .Y(men_men_n1057_));
  AOI210     u1029(.A0(men_men_n1057_), .A1(men_men_n1056_), .B0(men_men_n1036_), .Y(men_men_n1058_));
  AN4        u1030(.A(men_men_n1058_), .B(men_men_n1054_), .C(men_men_n1050_), .D(men_men_n1048_), .Y(men_men_n1059_));
  NO2        u1031(.A(men_men_n1013_), .B(men_men_n1011_), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n1028_), .B(men_men_n1022_), .Y(men_men_n1061_));
  AOI210     u1033(.A0(men_men_n1061_), .A1(men_men_n1060_), .B0(men_men_n1005_), .Y(men_men_n1062_));
  NAi41      u1034(.An(men_men_n1045_), .B(men_men_n1062_), .C(men_men_n1059_), .D(men_men_n1046_), .Y(men03));
  NO2        u1035(.A(men_men_n511_), .B(men_men_n580_), .Y(men_men_n1064_));
  NA4        u1036(.A(men_men_n90_), .B(men_men_n89_), .C(u), .D(men_men_n214_), .Y(men_men_n1065_));
  NA4        u1037(.A(men_men_n555_), .B(m), .C(men_men_n114_), .D(men_men_n214_), .Y(men_men_n1066_));
  NA3        u1038(.A(men_men_n1066_), .B(men_men_n365_), .C(men_men_n1065_), .Y(men_men_n1067_));
  NO3        u1039(.A(men_men_n1067_), .B(men_men_n1064_), .C(men_men_n975_), .Y(men_men_n1068_));
  NOi31      u1040(.An(men_men_n788_), .B(men_men_n832_), .C(men_men_n824_), .Y(men_men_n1069_));
  OAI220     u1041(.A0(men_men_n1069_), .A1(men_men_n673_), .B0(men_men_n1068_), .B1(men_men_n568_), .Y(men_men_n1070_));
  NA4        u1042(.A(i), .B(e), .C(men_men_n335_), .D(men_men_n329_), .Y(men_men_n1071_));
  OAI210     u1043(.A0(men_men_n802_), .A1(men_men_n411_), .B0(men_men_n1071_), .Y(men_men_n1072_));
  NOi31      u1044(.An(m), .B(n), .C(f), .Y(men_men_n1073_));
  NA2        u1045(.A(men_men_n1073_), .B(men_men_n51_), .Y(men_men_n1074_));
  AN2        u1046(.A(e), .B(c), .Y(men_men_n1075_));
  INV        u1047(.A(men_men_n1075_), .Y(men_men_n1076_));
  OAI220     u1048(.A0(men_men_n1076_), .A1(men_men_n1074_), .B0(men_men_n863_), .B1(men_men_n416_), .Y(men_men_n1077_));
  NA2        u1049(.A(men_men_n491_), .B(l), .Y(men_men_n1078_));
  NOi31      u1050(.An(men_men_n843_), .B(men_men_n1004_), .C(men_men_n1078_), .Y(men_men_n1079_));
  NO4        u1051(.A(men_men_n1079_), .B(men_men_n1077_), .C(men_men_n1072_), .D(men_men_n974_), .Y(men_men_n1080_));
  INV        u1052(.A(men_men_n1009_), .Y(men_men_n1081_));
  OR2        u1053(.A(u), .B(men_men_n1040_), .Y(men_men_n1082_));
  NA3        u1054(.A(men_men_n1082_), .B(men_men_n1081_), .C(men_men_n1080_), .Y(men_men_n1083_));
  NO4        u1055(.A(men_men_n1083_), .B(men_men_n1070_), .C(men_men_n804_), .D(men_men_n547_), .Y(men_men_n1084_));
  NA2        u1056(.A(c), .B(b), .Y(men_men_n1085_));
  NO2        u1057(.A(men_men_n684_), .B(men_men_n1085_), .Y(men_men_n1086_));
  OAI210     u1058(.A0(men_men_n841_), .A1(men_men_n818_), .B0(men_men_n405_), .Y(men_men_n1087_));
  OAI210     u1059(.A0(men_men_n1087_), .A1(men_men_n842_), .B0(men_men_n1086_), .Y(men_men_n1088_));
  NAi21      u1060(.An(men_men_n407_), .B(men_men_n1086_), .Y(men_men_n1089_));
  NA3        u1061(.A(men_men_n417_), .B(men_men_n540_), .C(f), .Y(men_men_n1090_));
  NA2        u1062(.A(men_men_n1090_), .B(men_men_n1089_), .Y(men_men_n1091_));
  OAI210     u1063(.A0(k), .A1(men_men_n286_), .B0(u), .Y(men_men_n1092_));
  NO2        u1064(.A(f), .B(men_men_n1055_), .Y(men_men_n1093_));
  INV        u1065(.A(men_men_n1093_), .Y(men_men_n1094_));
  AOI210     u1066(.A0(men_men_n1092_), .A1(men_men_n292_), .B0(men_men_n1094_), .Y(men_men_n1095_));
  AOI210     u1067(.A0(men_men_n1095_), .A1(men_men_n115_), .B0(men_men_n1091_), .Y(men_men_n1096_));
  NA2        u1068(.A(men_men_n451_), .B(men_men_n450_), .Y(men_men_n1097_));
  NO2        u1069(.A(men_men_n186_), .B(men_men_n234_), .Y(men_men_n1098_));
  NA2        u1070(.A(men_men_n1098_), .B(m), .Y(men_men_n1099_));
  NA3        u1071(.A(men_men_n893_), .B(men_men_n1078_), .C(men_men_n454_), .Y(men_men_n1100_));
  OAI210     u1072(.A0(men_men_n1100_), .A1(men_men_n312_), .B0(men_men_n452_), .Y(men_men_n1101_));
  AOI210     u1073(.A0(men_men_n1101_), .A1(men_men_n1097_), .B0(men_men_n1099_), .Y(men_men_n1102_));
  NA2        u1074(.A(men_men_n542_), .B(men_men_n400_), .Y(men_men_n1103_));
  NA2        u1075(.A(men_men_n162_), .B(men_men_n33_), .Y(men_men_n1104_));
  AOI210     u1076(.A0(men_men_n937_), .A1(men_men_n1104_), .B0(men_men_n215_), .Y(men_men_n1105_));
  NA2        u1077(.A(men_men_n1105_), .B(men_men_n1093_), .Y(men_men_n1106_));
  NO2        u1078(.A(men_men_n368_), .B(men_men_n367_), .Y(men_men_n1107_));
  AOI210     u1079(.A0(men_men_n1098_), .A1(men_men_n419_), .B0(men_men_n933_), .Y(men_men_n1108_));
  NAi41      u1080(.An(men_men_n1107_), .B(men_men_n1108_), .C(men_men_n1106_), .D(men_men_n1103_), .Y(men_men_n1109_));
  NO2        u1081(.A(men_men_n1109_), .B(men_men_n1102_), .Y(men_men_n1110_));
  NA4        u1082(.A(men_men_n1110_), .B(men_men_n1096_), .C(men_men_n1088_), .D(men_men_n1084_), .Y(men00));
  AOI210     u1083(.A0(men_men_n299_), .A1(men_men_n215_), .B0(men_men_n274_), .Y(men_men_n1112_));
  NO2        u1084(.A(men_men_n1112_), .B(men_men_n558_), .Y(men_men_n1113_));
  AOI210     u1085(.A0(men_men_n876_), .A1(men_men_n916_), .B0(men_men_n1072_), .Y(men_men_n1114_));
  NO3        u1086(.A(men_men_n1049_), .B(men_men_n933_), .C(men_men_n696_), .Y(men_men_n1115_));
  NA3        u1087(.A(men_men_n1115_), .B(men_men_n1114_), .C(men_men_n976_), .Y(men_men_n1116_));
  NA2        u1088(.A(men_men_n493_), .B(f), .Y(men_men_n1117_));
  OAI210     u1089(.A0(men_men_n983_), .A1(men_men_n40_), .B0(men_men_n629_), .Y(men_men_n1118_));
  NA3        u1090(.A(men_men_n1118_), .B(men_men_n254_), .C(n), .Y(men_men_n1119_));
  AOI210     u1091(.A0(men_men_n1119_), .A1(men_men_n1117_), .B0(men_men_n1013_), .Y(men_men_n1120_));
  NO4        u1092(.A(men_men_n1120_), .B(men_men_n1116_), .C(men_men_n1113_), .D(men_men_n1034_), .Y(men_men_n1121_));
  NA3        u1093(.A(men_men_n172_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1122_));
  NA3        u1094(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1123_));
  NOi31      u1095(.An(n), .B(m), .C(i), .Y(men_men_n1124_));
  NA3        u1096(.A(men_men_n1124_), .B(men_men_n632_), .C(men_men_n51_), .Y(men_men_n1125_));
  OAI210     u1097(.A0(men_men_n1123_), .A1(men_men_n1122_), .B0(men_men_n1125_), .Y(men_men_n1126_));
  INV        u1098(.A(men_men_n557_), .Y(men_men_n1127_));
  NO4        u1099(.A(men_men_n1127_), .B(men_men_n1126_), .C(men_men_n1107_), .D(men_men_n895_), .Y(men_men_n1128_));
  NO4        u1100(.A(men_men_n470_), .B(men_men_n350_), .C(men_men_n1085_), .D(men_men_n59_), .Y(men_men_n1129_));
  NA3        u1101(.A(men_men_n380_), .B(men_men_n222_), .C(u), .Y(men_men_n1130_));
  OA220      u1102(.A0(men_men_n1130_), .A1(men_men_n1123_), .B0(men_men_n381_), .B1(men_men_n137_), .Y(men_men_n1131_));
  NO2        u1103(.A(h), .B(u), .Y(men_men_n1132_));
  NA4        u1104(.A(men_men_n482_), .B(men_men_n448_), .C(men_men_n1132_), .D(c), .Y(men_men_n1133_));
  OAI220     u1105(.A0(men_men_n511_), .A1(men_men_n580_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1134_));
  AOI220     u1106(.A0(men_men_n1134_), .A1(men_men_n520_), .B0(men_men_n921_), .B1(men_men_n556_), .Y(men_men_n1135_));
  AOI220     u1107(.A0(men_men_n318_), .A1(men_men_n243_), .B0(men_men_n181_), .B1(men_men_n152_), .Y(men_men_n1136_));
  NA4        u1108(.A(men_men_n1136_), .B(men_men_n1135_), .C(men_men_n1133_), .D(men_men_n1131_), .Y(men_men_n1137_));
  NO3        u1109(.A(men_men_n1137_), .B(men_men_n1129_), .C(men_men_n264_), .Y(men_men_n1138_));
  INV        u1110(.A(men_men_n321_), .Y(men_men_n1139_));
  AOI210     u1111(.A0(men_men_n243_), .A1(men_men_n340_), .B0(men_men_n559_), .Y(men_men_n1140_));
  NA3        u1112(.A(men_men_n1140_), .B(men_men_n1139_), .C(men_men_n157_), .Y(men_men_n1141_));
  NO2        u1113(.A(men_men_n236_), .B(men_men_n185_), .Y(men_men_n1142_));
  NA2        u1114(.A(men_men_n1142_), .B(men_men_n417_), .Y(men_men_n1143_));
  NA3        u1115(.A(men_men_n183_), .B(men_men_n114_), .C(u), .Y(men_men_n1144_));
  NA3        u1116(.A(men_men_n448_), .B(men_men_n40_), .C(f), .Y(men_men_n1145_));
  NOi31      u1117(.An(j), .B(men_men_n1145_), .C(men_men_n1144_), .Y(men_men_n1146_));
  NAi31      u1118(.An(men_men_n189_), .B(men_men_n838_), .C(men_men_n448_), .Y(men_men_n1147_));
  NAi31      u1119(.An(men_men_n1146_), .B(men_men_n1147_), .C(men_men_n1143_), .Y(men_men_n1148_));
  NO2        u1120(.A(men_men_n273_), .B(men_men_n75_), .Y(men_men_n1149_));
  NO3        u1121(.A(men_men_n416_), .B(men_men_n814_), .C(n), .Y(men_men_n1150_));
  AOI210     u1122(.A0(men_men_n1150_), .A1(men_men_n1149_), .B0(men_men_n1045_), .Y(men_men_n1151_));
  NAi31      u1123(.An(men_men_n1016_), .B(men_men_n1151_), .C(men_men_n74_), .Y(men_men_n1152_));
  NO4        u1124(.A(men_men_n1152_), .B(men_men_n1148_), .C(men_men_n1141_), .D(men_men_n502_), .Y(men_men_n1153_));
  AN3        u1125(.A(men_men_n1153_), .B(men_men_n1138_), .C(men_men_n1128_), .Y(men_men_n1154_));
  NA2        u1126(.A(men_men_n520_), .B(men_men_n104_), .Y(men_men_n1155_));
  NA3        u1127(.A(men_men_n1073_), .B(men_men_n591_), .C(men_men_n447_), .Y(men_men_n1156_));
  NA4        u1128(.A(men_men_n1156_), .B(men_men_n543_), .C(men_men_n1155_), .D(men_men_n239_), .Y(men_men_n1157_));
  NA2        u1129(.A(men_men_n1067_), .B(men_men_n520_), .Y(men_men_n1158_));
  NA4        u1130(.A(men_men_n632_), .B(men_men_n206_), .C(men_men_n222_), .D(men_men_n166_), .Y(men_men_n1159_));
  NA3        u1131(.A(men_men_n1159_), .B(men_men_n1158_), .C(men_men_n296_), .Y(men_men_n1160_));
  OAI210     u1132(.A0(men_men_n446_), .A1(men_men_n121_), .B0(men_men_n844_), .Y(men_men_n1161_));
  AOI220     u1133(.A0(men_men_n1161_), .A1(men_men_n1100_), .B0(men_men_n542_), .B1(men_men_n400_), .Y(men_men_n1162_));
  OR4        u1134(.A(men_men_n1013_), .B(men_men_n270_), .C(men_men_n223_), .D(e), .Y(men_men_n1163_));
  NO2        u1135(.A(men_men_n218_), .B(men_men_n215_), .Y(men_men_n1164_));
  NA2        u1136(.A(n), .B(e), .Y(men_men_n1165_));
  NO2        u1137(.A(men_men_n1165_), .B(men_men_n150_), .Y(men_men_n1166_));
  AOI220     u1138(.A0(men_men_n1166_), .A1(men_men_n272_), .B0(men_men_n828_), .B1(men_men_n1164_), .Y(men_men_n1167_));
  OAI210     u1139(.A0(men_men_n351_), .A1(men_men_n313_), .B0(men_men_n433_), .Y(men_men_n1168_));
  NA4        u1140(.A(men_men_n1168_), .B(men_men_n1167_), .C(men_men_n1163_), .D(men_men_n1162_), .Y(men_men_n1169_));
  AOI210     u1141(.A0(men_men_n1166_), .A1(men_men_n830_), .B0(men_men_n803_), .Y(men_men_n1170_));
  NO2        u1142(.A(men_men_n68_), .B(h), .Y(men_men_n1171_));
  NO3        u1143(.A(men_men_n1013_), .B(men_men_n1011_), .C(men_men_n713_), .Y(men_men_n1172_));
  OAI210     u1144(.A0(men_men_n1053_), .A1(men_men_n1172_), .B0(men_men_n1171_), .Y(men_men_n1173_));
  NA3        u1145(.A(men_men_n1173_), .B(men_men_n1170_), .C(men_men_n846_), .Y(men_men_n1174_));
  NO4        u1146(.A(men_men_n1174_), .B(men_men_n1169_), .C(men_men_n1160_), .D(men_men_n1157_), .Y(men_men_n1175_));
  NA2        u1147(.A(men_men_n819_), .B(men_men_n745_), .Y(men_men_n1176_));
  NA4        u1148(.A(men_men_n1176_), .B(men_men_n1175_), .C(men_men_n1154_), .D(men_men_n1121_), .Y(men01));
  NO4        u1149(.A(men_men_n785_), .B(men_men_n777_), .C(men_men_n462_), .D(men_men_n280_), .Y(men_men_n1178_));
  NA2        u1150(.A(men_men_n1178_), .B(men_men_n993_), .Y(men_men_n1179_));
  NA2        u1151(.A(men_men_n569_), .B(men_men_n92_), .Y(men_men_n1180_));
  NA2        u1152(.A(men_men_n537_), .B(men_men_n269_), .Y(men_men_n1181_));
  NA2        u1153(.A(men_men_n936_), .B(men_men_n1181_), .Y(men_men_n1182_));
  NA3        u1154(.A(men_men_n1182_), .B(men_men_n1180_), .C(men_men_n889_), .Y(men_men_n1183_));
  NA2        u1155(.A(men_men_n691_), .B(men_men_n99_), .Y(men_men_n1184_));
  NO2        u1156(.A(men_men_n1184_), .B(i), .Y(men_men_n1185_));
  OAI210     u1157(.A0(men_men_n764_), .A1(men_men_n586_), .B0(men_men_n1159_), .Y(men_men_n1186_));
  AOI210     u1158(.A0(men_men_n1185_), .A1(men_men_n620_), .B0(men_men_n1186_), .Y(men_men_n1187_));
  INV        u1159(.A(men_men_n119_), .Y(men_men_n1188_));
  OA220      u1160(.A0(men_men_n1188_), .A1(men_men_n566_), .B0(men_men_n645_), .B1(men_men_n365_), .Y(men_men_n1189_));
  NAi41      u1161(.An(men_men_n165_), .B(men_men_n1189_), .C(men_men_n1187_), .D(men_men_n875_), .Y(men_men_n1190_));
  NO3        u1162(.A(men_men_n765_), .B(men_men_n657_), .C(men_men_n496_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n1191_), .B(men_men_n140_), .Y(men_men_n1192_));
  NO4        u1164(.A(men_men_n1192_), .B(men_men_n1190_), .C(men_men_n1183_), .D(men_men_n1179_), .Y(men_men_n1193_));
  NA2        u1165(.A(men_men_n1130_), .B(men_men_n207_), .Y(men_men_n1194_));
  OAI210     u1166(.A0(men_men_n1194_), .A1(men_men_n302_), .B0(men_men_n515_), .Y(men_men_n1195_));
  NOi21      u1167(.An(men_men_n544_), .B(men_men_n563_), .Y(men_men_n1196_));
  NA2        u1168(.A(men_men_n1196_), .B(e), .Y(men_men_n1197_));
  AOI210     u1169(.A0(men_men_n204_), .A1(men_men_n91_), .B0(men_men_n214_), .Y(men_men_n1198_));
  OAI210     u1170(.A0(men_men_n791_), .A1(men_men_n417_), .B0(men_men_n1198_), .Y(men_men_n1199_));
  NA2        u1171(.A(men_men_n203_), .B(men_men_n34_), .Y(men_men_n1200_));
  OR2        u1172(.A(men_men_n1200_), .B(men_men_n328_), .Y(men_men_n1201_));
  NA4        u1173(.A(men_men_n1201_), .B(men_men_n1199_), .C(men_men_n1197_), .D(men_men_n1195_), .Y(men_men_n1202_));
  AOI210     u1174(.A0(men_men_n578_), .A1(men_men_n119_), .B0(men_men_n584_), .Y(men_men_n1203_));
  OAI210     u1175(.A0(men_men_n1188_), .A1(men_men_n575_), .B0(men_men_n1203_), .Y(men_men_n1204_));
  NO3        u1176(.A(men_men_n802_), .B(men_men_n204_), .C(men_men_n398_), .Y(men_men_n1205_));
  NO2        u1177(.A(men_men_n1205_), .B(men_men_n933_), .Y(men_men_n1206_));
  NA2        u1178(.A(men_men_n1206_), .B(men_men_n767_), .Y(men_men_n1207_));
  NO3        u1179(.A(men_men_n1207_), .B(men_men_n1204_), .C(men_men_n1202_), .Y(men_men_n1208_));
  NA3        u1180(.A(men_men_n587_), .B(men_men_n29_), .C(f), .Y(men_men_n1209_));
  NO2        u1181(.A(men_men_n1209_), .B(men_men_n204_), .Y(men_men_n1210_));
  AOI210     u1182(.A0(men_men_n489_), .A1(men_men_n58_), .B0(men_men_n1210_), .Y(men_men_n1211_));
  OR3        u1183(.A(men_men_n1184_), .B(men_men_n588_), .C(i), .Y(men_men_n1212_));
  NO2        u1184(.A(men_men_n207_), .B(men_men_n113_), .Y(men_men_n1213_));
  NO2        u1185(.A(men_men_n1213_), .B(men_men_n1126_), .Y(men_men_n1214_));
  NA4        u1186(.A(men_men_n1214_), .B(men_men_n1212_), .C(men_men_n1211_), .D(men_men_n744_), .Y(men_men_n1215_));
  NO2        u1187(.A(men_men_n941_), .B(men_men_n229_), .Y(men_men_n1216_));
  NO2        u1188(.A(men_men_n942_), .B(men_men_n538_), .Y(men_men_n1217_));
  OAI210     u1189(.A0(men_men_n1217_), .A1(men_men_n1216_), .B0(men_men_n333_), .Y(men_men_n1218_));
  NO3        u1190(.A(men_men_n81_), .B(men_men_n300_), .C(men_men_n45_), .Y(men_men_n1219_));
  NA2        u1191(.A(men_men_n1219_), .B(men_men_n536_), .Y(men_men_n1220_));
  NA2        u1192(.A(men_men_n1220_), .B(men_men_n652_), .Y(men_men_n1221_));
  OR2        u1193(.A(men_men_n1130_), .B(men_men_n1123_), .Y(men_men_n1222_));
  NO2        u1194(.A(men_men_n365_), .B(men_men_n73_), .Y(men_men_n1223_));
  INV        u1195(.A(men_men_n1223_), .Y(men_men_n1224_));
  NA2        u1196(.A(men_men_n1219_), .B(men_men_n794_), .Y(men_men_n1225_));
  NA4        u1197(.A(men_men_n1225_), .B(men_men_n1224_), .C(men_men_n1222_), .D(men_men_n383_), .Y(men_men_n1226_));
  NOi41      u1198(.An(men_men_n1218_), .B(men_men_n1226_), .C(men_men_n1221_), .D(men_men_n1215_), .Y(men_men_n1227_));
  NO2        u1199(.A(men_men_n133_), .B(men_men_n45_), .Y(men_men_n1228_));
  AN2        u1200(.A(men_men_n1228_), .B(men_men_n689_), .Y(men_men_n1229_));
  NA2        u1201(.A(men_men_n1229_), .B(men_men_n333_), .Y(men_men_n1230_));
  INV        u1202(.A(men_men_n137_), .Y(men_men_n1231_));
  NO3        u1203(.A(men_men_n1051_), .B(men_men_n180_), .C(men_men_n89_), .Y(men_men_n1232_));
  AOI220     u1204(.A0(men_men_n1232_), .A1(men_men_n1231_), .B0(men_men_n1219_), .B1(men_men_n945_), .Y(men_men_n1233_));
  NA2        u1205(.A(men_men_n1233_), .B(men_men_n1230_), .Y(men_men_n1234_));
  NO2        u1206(.A(men_men_n599_), .B(men_men_n598_), .Y(men_men_n1235_));
  NO4        u1207(.A(men_men_n1051_), .B(men_men_n1235_), .C(men_men_n179_), .D(men_men_n89_), .Y(men_men_n1236_));
  NO3        u1208(.A(men_men_n1236_), .B(men_men_n1234_), .C(men_men_n624_), .Y(men_men_n1237_));
  NA4        u1209(.A(men_men_n1237_), .B(men_men_n1227_), .C(men_men_n1208_), .D(men_men_n1193_), .Y(men06));
  NO2        u1210(.A(men_men_n399_), .B(men_men_n541_), .Y(men_men_n1239_));
  NA2        u1211(.A(men_men_n265_), .B(men_men_n1239_), .Y(men_men_n1240_));
  NO3        u1212(.A(men_men_n582_), .B(men_men_n789_), .C(men_men_n585_), .Y(men_men_n1241_));
  OR2        u1213(.A(men_men_n1241_), .B(men_men_n863_), .Y(men_men_n1242_));
  NA3        u1214(.A(men_men_n1242_), .B(men_men_n1240_), .C(men_men_n1218_), .Y(men_men_n1243_));
  NO3        u1215(.A(men_men_n1243_), .B(men_men_n1221_), .C(men_men_n253_), .Y(men_men_n1244_));
  NA2        u1216(.A(i), .B(men_men_n946_), .Y(men_men_n1245_));
  AOI210     u1217(.A0(i), .A1(men_men_n539_), .B0(men_men_n1229_), .Y(men_men_n1246_));
  AOI210     u1218(.A0(men_men_n1246_), .A1(men_men_n1245_), .B0(men_men_n330_), .Y(men_men_n1247_));
  OAI210     u1219(.A0(men_men_n91_), .A1(men_men_n40_), .B0(men_men_n656_), .Y(men_men_n1248_));
  NA2        u1220(.A(men_men_n1248_), .B(men_men_n356_), .Y(men_men_n1249_));
  NO2        u1221(.A(men_men_n499_), .B(men_men_n177_), .Y(men_men_n1250_));
  NO2        u1222(.A(men_men_n592_), .B(men_men_n1074_), .Y(men_men_n1251_));
  NO3        u1223(.A(men_men_n1251_), .B(men_men_n139_), .C(men_men_n1250_), .Y(men_men_n1252_));
  OR2        u1224(.A(men_men_n583_), .B(men_men_n581_), .Y(men_men_n1253_));
  NO2        u1225(.A(men_men_n364_), .B(men_men_n138_), .Y(men_men_n1254_));
  AOI210     u1226(.A0(men_men_n1254_), .A1(men_men_n569_), .B0(men_men_n1253_), .Y(men_men_n1255_));
  NA3        u1227(.A(men_men_n1255_), .B(men_men_n1252_), .C(men_men_n1249_), .Y(men_men_n1256_));
  NO2        u1228(.A(men_men_n735_), .B(men_men_n363_), .Y(men_men_n1257_));
  NO3        u1229(.A(men_men_n658_), .B(men_men_n746_), .C(men_men_n620_), .Y(men_men_n1258_));
  NOi21      u1230(.An(men_men_n1257_), .B(men_men_n1258_), .Y(men_men_n1259_));
  AN2        u1231(.A(men_men_n929_), .B(men_men_n628_), .Y(men_men_n1260_));
  NO4        u1232(.A(men_men_n1260_), .B(men_men_n1259_), .C(men_men_n1256_), .D(men_men_n1247_), .Y(men_men_n1261_));
  NO2        u1233(.A(men_men_n784_), .B(men_men_n275_), .Y(men_men_n1262_));
  OAI220     u1234(.A0(men_men_n720_), .A1(men_men_n47_), .B0(men_men_n225_), .B1(men_men_n601_), .Y(men_men_n1263_));
  NO2        u1235(.A(men_men_n275_), .B(c), .Y(men_men_n1264_));
  AOI220     u1236(.A0(men_men_n1264_), .A1(men_men_n1263_), .B0(men_men_n1262_), .B1(men_men_n265_), .Y(men_men_n1265_));
  NO3        u1237(.A(men_men_n241_), .B(men_men_n106_), .C(men_men_n282_), .Y(men_men_n1266_));
  OAI210     u1238(.A0(l), .A1(i), .B0(k), .Y(men_men_n1267_));
  NO3        u1239(.A(men_men_n1267_), .B(men_men_n580_), .C(j), .Y(men_men_n1268_));
  NOi21      u1240(.An(men_men_n1268_), .B(men_men_n73_), .Y(men_men_n1269_));
  NO3        u1241(.A(men_men_n1269_), .B(men_men_n1266_), .C(men_men_n1077_), .Y(men_men_n1270_));
  NA4        u1242(.A(men_men_n775_), .B(men_men_n774_), .C(men_men_n426_), .D(men_men_n857_), .Y(men_men_n1271_));
  NAi31      u1243(.An(men_men_n735_), .B(men_men_n1271_), .C(men_men_n203_), .Y(men_men_n1272_));
  NA3        u1244(.A(men_men_n1272_), .B(men_men_n1270_), .C(men_men_n1265_), .Y(men_men_n1273_));
  OR2        u1245(.A(men_men_n764_), .B(men_men_n526_), .Y(men_men_n1274_));
  OR3        u1246(.A(men_men_n367_), .B(men_men_n225_), .C(men_men_n601_), .Y(men_men_n1275_));
  INV        u1247(.A(men_men_n369_), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n1268_), .B(men_men_n771_), .Y(men_men_n1277_));
  NA4        u1249(.A(men_men_n1277_), .B(men_men_n1276_), .C(men_men_n1275_), .D(men_men_n1274_), .Y(men_men_n1278_));
  AOI220     u1250(.A0(men_men_n1257_), .A1(men_men_n745_), .B0(men_men_n1254_), .B1(men_men_n235_), .Y(men_men_n1279_));
  NO3        u1251(.A(men_men_n855_), .B(men_men_n485_), .C(men_men_n465_), .Y(men_men_n1280_));
  NA3        u1252(.A(men_men_n1280_), .B(men_men_n1279_), .C(men_men_n1225_), .Y(men_men_n1281_));
  NAi21      u1253(.An(j), .B(i), .Y(men_men_n1282_));
  NO4        u1254(.A(men_men_n1235_), .B(men_men_n1282_), .C(men_men_n432_), .D(men_men_n232_), .Y(men_men_n1283_));
  NO4        u1255(.A(men_men_n1283_), .B(men_men_n1281_), .C(men_men_n1278_), .D(men_men_n1273_), .Y(men_men_n1284_));
  NA4        u1256(.A(men_men_n1284_), .B(men_men_n1261_), .C(men_men_n1244_), .D(men_men_n1237_), .Y(men07));
  NOi21      u1257(.An(j), .B(k), .Y(men_men_n1286_));
  NAi32      u1258(.An(m), .Bn(b), .C(n), .Y(men_men_n1287_));
  NO3        u1259(.A(men_men_n1287_), .B(u), .C(f), .Y(men_men_n1288_));
  OAI210     u1260(.A0(men_men_n320_), .A1(j), .B0(men_men_n1288_), .Y(men_men_n1289_));
  NAi21      u1261(.An(f), .B(c), .Y(men_men_n1290_));
  OR2        u1262(.A(e), .B(d), .Y(men_men_n1291_));
  NOi31      u1263(.An(n), .B(m), .C(b), .Y(men_men_n1292_));
  INV        u1264(.A(men_men_n1289_), .Y(men_men_n1293_));
  NOi41      u1265(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1294_));
  NA3        u1266(.A(men_men_n1294_), .B(men_men_n848_), .C(men_men_n401_), .Y(men_men_n1295_));
  INV        u1267(.A(men_men_n1295_), .Y(men_men_n1296_));
  NA2        u1268(.A(men_men_n1053_), .B(men_men_n222_), .Y(men_men_n1297_));
  NO2        u1269(.A(men_men_n1297_), .B(men_men_n61_), .Y(men_men_n1298_));
  NO2        u1270(.A(k), .B(i), .Y(men_men_n1299_));
  NO2        u1271(.A(men_men_n1031_), .B(men_men_n307_), .Y(men_men_n1300_));
  NA2        u1272(.A(men_men_n1171_), .B(men_men_n290_), .Y(men_men_n1301_));
  INV        u1273(.A(men_men_n1301_), .Y(men_men_n1302_));
  NO4        u1274(.A(men_men_n1302_), .B(men_men_n1298_), .C(men_men_n1296_), .D(men_men_n1293_), .Y(men_men_n1303_));
  NO3        u1275(.A(e), .B(d), .C(c), .Y(men_men_n1304_));
  OAI210     u1276(.A0(men_men_n134_), .A1(men_men_n215_), .B0(men_men_n589_), .Y(men_men_n1305_));
  NA2        u1277(.A(men_men_n1305_), .B(men_men_n1304_), .Y(men_men_n1306_));
  INV        u1278(.A(men_men_n1306_), .Y(men_men_n1307_));
  NO3        u1279(.A(n), .B(m), .C(i), .Y(men_men_n1308_));
  OAI210     u1280(.A0(men_men_n1075_), .A1(men_men_n160_), .B0(men_men_n1308_), .Y(men_men_n1309_));
  NO2        u1281(.A(i), .B(u), .Y(men_men_n1310_));
  OR3        u1282(.A(men_men_n1310_), .B(men_men_n1287_), .C(men_men_n72_), .Y(men_men_n1311_));
  OAI220     u1283(.A0(men_men_n1311_), .A1(j), .B0(men_men_n1309_), .B1(f), .Y(men_men_n1312_));
  NA3        u1284(.A(men_men_n679_), .B(men_men_n665_), .C(men_men_n114_), .Y(men_men_n1313_));
  NA3        u1285(.A(men_men_n1292_), .B(l), .C(men_men_n654_), .Y(men_men_n1314_));
  AOI210     u1286(.A0(men_men_n1314_), .A1(men_men_n1313_), .B0(men_men_n45_), .Y(men_men_n1315_));
  NA2        u1287(.A(men_men_n1308_), .B(men_men_n626_), .Y(men_men_n1316_));
  NO3        u1288(.A(men_men_n432_), .B(d), .C(c), .Y(men_men_n1317_));
  NO3        u1289(.A(men_men_n1315_), .B(men_men_n1312_), .C(men_men_n1307_), .Y(men_men_n1318_));
  NO2        u1290(.A(men_men_n151_), .B(h), .Y(men_men_n1319_));
  NO2        u1291(.A(u), .B(c), .Y(men_men_n1320_));
  NO2        u1292(.A(men_men_n437_), .B(a), .Y(men_men_n1321_));
  NA3        u1293(.A(men_men_n1321_), .B(k), .C(men_men_n115_), .Y(men_men_n1322_));
  NO2        u1294(.A(i), .B(h), .Y(men_men_n1323_));
  NA2        u1295(.A(men_men_n1323_), .B(men_men_n222_), .Y(men_men_n1324_));
  AOI210     u1296(.A0(men_men_n254_), .A1(men_men_n117_), .B0(men_men_n515_), .Y(men_men_n1325_));
  NO2        u1297(.A(men_men_n1325_), .B(men_men_n1324_), .Y(men_men_n1326_));
  NO2        u1298(.A(men_men_n742_), .B(men_men_n190_), .Y(men_men_n1327_));
  NOi31      u1299(.An(m), .B(n), .C(b), .Y(men_men_n1328_));
  NOi31      u1300(.An(f), .B(d), .C(c), .Y(men_men_n1329_));
  NA2        u1301(.A(men_men_n1329_), .B(men_men_n1328_), .Y(men_men_n1330_));
  INV        u1302(.A(men_men_n1330_), .Y(men_men_n1331_));
  NO3        u1303(.A(men_men_n1331_), .B(men_men_n1327_), .C(men_men_n1326_), .Y(men_men_n1332_));
  NO3        u1304(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1333_));
  AN2        u1305(.A(men_men_n1332_), .B(men_men_n1322_), .Y(men_men_n1334_));
  NA2        u1306(.A(men_men_n1292_), .B(men_men_n376_), .Y(men_men_n1335_));
  NO2        u1307(.A(men_men_n1335_), .B(men_men_n1010_), .Y(men_men_n1336_));
  NO2        u1308(.A(men_men_n190_), .B(b), .Y(men_men_n1337_));
  NO2        u1309(.A(i), .B(men_men_n214_), .Y(men_men_n1338_));
  NA4        u1310(.A(men_men_n1098_), .B(men_men_n1338_), .C(men_men_n107_), .D(m), .Y(men_men_n1339_));
  NAi21      u1311(.An(men_men_n1336_), .B(men_men_n1339_), .Y(men_men_n1340_));
  NO4        u1312(.A(men_men_n134_), .B(u), .C(f), .D(e), .Y(men_men_n1341_));
  NA2        u1313(.A(men_men_n1299_), .B(h), .Y(men_men_n1342_));
  NA2        u1314(.A(men_men_n195_), .B(men_men_n101_), .Y(men_men_n1343_));
  NOi41      u1315(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1344_));
  NA2        u1316(.A(men_men_n1344_), .B(men_men_n115_), .Y(men_men_n1345_));
  INV        u1317(.A(men_men_n1345_), .Y(men_men_n1346_));
  OR3        u1318(.A(men_men_n526_), .B(men_men_n525_), .C(men_men_n114_), .Y(men_men_n1347_));
  NA2        u1319(.A(men_men_n1073_), .B(men_men_n398_), .Y(men_men_n1348_));
  OAI220     u1320(.A0(men_men_n1348_), .A1(men_men_n425_), .B0(men_men_n1347_), .B1(men_men_n300_), .Y(men_men_n1349_));
  AO210      u1321(.A0(men_men_n1349_), .A1(men_men_n117_), .B0(men_men_n1346_), .Y(men_men_n1350_));
  NO2        u1322(.A(men_men_n1350_), .B(men_men_n1340_), .Y(men_men_n1351_));
  NA4        u1323(.A(men_men_n1351_), .B(men_men_n1334_), .C(men_men_n1318_), .D(men_men_n1303_), .Y(men_men_n1352_));
  NO2        u1324(.A(men_men_n1085_), .B(men_men_n112_), .Y(men_men_n1353_));
  NO2        u1325(.A(c), .B(men_men_n1316_), .Y(men_men_n1354_));
  NA2        u1326(.A(men_men_n216_), .B(men_men_n183_), .Y(men_men_n1355_));
  AOI210     u1327(.A0(men_men_n1355_), .A1(men_men_n1144_), .B0(c), .Y(men_men_n1356_));
  NO2        u1328(.A(men_men_n1356_), .B(men_men_n1354_), .Y(men_men_n1357_));
  NA3        u1329(.A(men_men_n1333_), .B(men_men_n1291_), .C(men_men_n1073_), .Y(men_men_n1358_));
  NAi31      u1330(.An(men_men_n1323_), .B(men_men_n1039_), .C(men_men_n173_), .Y(men_men_n1359_));
  NA2        u1331(.A(men_men_n1359_), .B(men_men_n1358_), .Y(men_men_n1360_));
  INV        u1332(.A(men_men_n1360_), .Y(men_men_n1361_));
  NO3        u1333(.A(m), .B(men_men_n563_), .C(u), .Y(men_men_n1362_));
  NOi21      u1334(.An(men_men_n1355_), .B(men_men_n1362_), .Y(men_men_n1363_));
  AOI210     u1335(.A0(men_men_n1363_), .A1(men_men_n1343_), .B0(men_men_n1019_), .Y(men_men_n1364_));
  INV        u1336(.A(men_men_n49_), .Y(men_men_n1365_));
  NA2        u1337(.A(men_men_n1365_), .B(men_men_n1132_), .Y(men_men_n1366_));
  INV        u1338(.A(men_men_n1366_), .Y(men_men_n1367_));
  OAI220     u1339(.A0(men_men_n650_), .A1(u), .B0(men_men_n225_), .B1(c), .Y(men_men_n1368_));
  AOI210     u1340(.A0(men_men_n1337_), .A1(men_men_n41_), .B0(men_men_n1368_), .Y(men_men_n1369_));
  NO2        u1341(.A(men_men_n134_), .B(l), .Y(men_men_n1370_));
  NO2        u1342(.A(men_men_n225_), .B(k), .Y(men_men_n1371_));
  OAI210     u1343(.A0(men_men_n1371_), .A1(men_men_n1323_), .B0(men_men_n1370_), .Y(men_men_n1372_));
  OAI220     u1344(.A0(men_men_n1372_), .A1(men_men_n31_), .B0(men_men_n1369_), .B1(men_men_n180_), .Y(men_men_n1373_));
  NO3        u1345(.A(men_men_n1347_), .B(men_men_n448_), .C(men_men_n347_), .Y(men_men_n1374_));
  NO4        u1346(.A(men_men_n1374_), .B(men_men_n1373_), .C(men_men_n1367_), .D(men_men_n1364_), .Y(men_men_n1375_));
  NO3        u1347(.A(men_men_n1055_), .B(men_men_n1291_), .C(men_men_n49_), .Y(men_men_n1376_));
  NA2        u1348(.A(men_men_n1056_), .B(men_men_n1448_), .Y(men_men_n1377_));
  NO2        u1349(.A(men_men_n1377_), .B(j), .Y(men_men_n1378_));
  NA3        u1350(.A(men_men_n1353_), .B(men_men_n448_), .C(f), .Y(men_men_n1379_));
  NA2        u1351(.A(men_men_n183_), .B(men_men_n114_), .Y(men_men_n1380_));
  NO2        u1352(.A(men_men_n1286_), .B(men_men_n42_), .Y(men_men_n1381_));
  AOI210     u1353(.A0(men_men_n115_), .A1(men_men_n40_), .B0(men_men_n1381_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n1382_), .B(men_men_n1379_), .Y(men_men_n1383_));
  AOI210     u1355(.A0(men_men_n510_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1384_));
  NA2        u1356(.A(men_men_n1384_), .B(men_men_n1321_), .Y(men_men_n1385_));
  INV        u1357(.A(men_men_n179_), .Y(men_men_n1386_));
  NOi21      u1358(.An(d), .B(f), .Y(men_men_n1387_));
  NO3        u1359(.A(men_men_n1329_), .B(men_men_n1387_), .C(men_men_n40_), .Y(men_men_n1388_));
  NA2        u1360(.A(men_men_n1388_), .B(men_men_n1386_), .Y(men_men_n1389_));
  NA2        u1361(.A(men_men_n1321_), .B(men_men_n1381_), .Y(men_men_n1390_));
  NO2        u1362(.A(men_men_n300_), .B(c), .Y(men_men_n1391_));
  NA2        u1363(.A(men_men_n1391_), .B(men_men_n527_), .Y(men_men_n1392_));
  NA4        u1364(.A(men_men_n1392_), .B(men_men_n1390_), .C(men_men_n1389_), .D(men_men_n1385_), .Y(men_men_n1393_));
  NO3        u1365(.A(men_men_n1393_), .B(men_men_n1383_), .C(men_men_n1378_), .Y(men_men_n1394_));
  NA4        u1366(.A(men_men_n1394_), .B(men_men_n1375_), .C(men_men_n1361_), .D(men_men_n1357_), .Y(men_men_n1395_));
  OAI220     u1367(.A0(men_men_n448_), .A1(men_men_n300_), .B0(men_men_n133_), .B1(men_men_n59_), .Y(men_men_n1396_));
  NA2        u1368(.A(men_men_n1396_), .B(men_men_n1300_), .Y(men_men_n1397_));
  OAI210     u1369(.A0(men_men_n1341_), .A1(men_men_n1292_), .B0(men_men_n860_), .Y(men_men_n1398_));
  OAI210     u1370(.A0(c), .A1(men_men_n134_), .B0(men_men_n179_), .Y(men_men_n1399_));
  NA2        u1371(.A(men_men_n1399_), .B(men_men_n607_), .Y(men_men_n1400_));
  NA3        u1372(.A(men_men_n1400_), .B(men_men_n1398_), .C(men_men_n1397_), .Y(men_men_n1401_));
  NA2        u1373(.A(men_men_n1320_), .B(men_men_n1387_), .Y(men_men_n1402_));
  NO2        u1374(.A(men_men_n1402_), .B(m), .Y(men_men_n1403_));
  NA3        u1375(.A(men_men_n1053_), .B(men_men_n110_), .C(men_men_n222_), .Y(men_men_n1404_));
  NA2        u1376(.A(men_men_n112_), .B(men_men_n1328_), .Y(men_men_n1405_));
  NA2        u1377(.A(men_men_n1405_), .B(men_men_n1404_), .Y(men_men_n1406_));
  NO3        u1378(.A(men_men_n1406_), .B(men_men_n1403_), .C(men_men_n1401_), .Y(men_men_n1407_));
  NO2        u1379(.A(men_men_n1290_), .B(e), .Y(men_men_n1408_));
  NA2        u1380(.A(men_men_n1408_), .B(men_men_n396_), .Y(men_men_n1409_));
  OR3        u1381(.A(men_men_n1371_), .B(men_men_n1171_), .C(men_men_n134_), .Y(men_men_n1410_));
  NO2        u1382(.A(men_men_n1410_), .B(men_men_n1409_), .Y(men_men_n1411_));
  NO3        u1383(.A(men_men_n1347_), .B(men_men_n347_), .C(a), .Y(men_men_n1412_));
  NO2        u1384(.A(men_men_n1412_), .B(men_men_n1411_), .Y(men_men_n1413_));
  NA2        u1385(.A(men_men_n525_), .B(u), .Y(men_men_n1414_));
  AOI210     u1386(.A0(men_men_n1414_), .A1(men_men_n1317_), .B0(men_men_n1376_), .Y(men_men_n1415_));
  NO2        u1387(.A(men_men_n1415_), .B(men_men_n214_), .Y(men_men_n1416_));
  NA2        u1388(.A(men_men_n879_), .B(men_men_n408_), .Y(men_men_n1417_));
  OR2        u1389(.A(men_men_n1417_), .B(men_men_n525_), .Y(men_men_n1418_));
  NO2        u1390(.A(men_men_n1418_), .B(men_men_n179_), .Y(men_men_n1419_));
  NO2        u1391(.A(m), .B(i), .Y(men_men_n1420_));
  NA2        u1392(.A(men_men_n1420_), .B(men_men_n1319_), .Y(men_men_n1421_));
  INV        u1393(.A(men_men_n1421_), .Y(men_men_n1422_));
  NO3        u1394(.A(men_men_n1422_), .B(men_men_n1419_), .C(men_men_n1416_), .Y(men_men_n1423_));
  NA3        u1395(.A(men_men_n1423_), .B(men_men_n1413_), .C(men_men_n1407_), .Y(men_men_n1424_));
  NA3        u1396(.A(men_men_n935_), .B(men_men_n141_), .C(men_men_n46_), .Y(men_men_n1425_));
  NO2        u1397(.A(men_men_n72_), .B(c), .Y(men_men_n1426_));
  NO4        u1398(.A(f), .B(men_men_n189_), .C(men_men_n435_), .D(men_men_n45_), .Y(men_men_n1427_));
  AOI210     u1399(.A0(men_men_n1386_), .A1(men_men_n1426_), .B0(men_men_n1427_), .Y(men_men_n1428_));
  NO2        u1400(.A(men_men_n1290_), .B(men_men_n1380_), .Y(men_men_n1429_));
  NO2        u1401(.A(men_men_n1425_), .B(men_men_n112_), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n1430_), .B(men_men_n1429_), .Y(men_men_n1431_));
  NO2        u1403(.A(men_men_n1379_), .B(men_men_n69_), .Y(men_men_n1432_));
  NO2        u1404(.A(men_men_n1299_), .B(men_men_n119_), .Y(men_men_n1433_));
  NO2        u1405(.A(men_men_n1433_), .B(men_men_n1335_), .Y(men_men_n1434_));
  NO2        u1406(.A(men_men_n1434_), .B(men_men_n1432_), .Y(men_men_n1435_));
  NA3        u1407(.A(men_men_n1435_), .B(men_men_n1431_), .C(men_men_n1428_), .Y(men_men_n1436_));
  OR4        u1408(.A(men_men_n1436_), .B(men_men_n1424_), .C(men_men_n1395_), .D(men_men_n1352_), .Y(men04));
  NOi31      u1409(.An(men_men_n1341_), .B(men_men_n1342_), .C(men_men_n1013_), .Y(men_men_n1438_));
  NO4        u1410(.A(men_men_n1291_), .B(men_men_n1004_), .C(men_men_n467_), .D(j), .Y(men_men_n1439_));
  OR3        u1411(.A(men_men_n1439_), .B(men_men_n1438_), .C(men_men_n1029_), .Y(men_men_n1440_));
  NO2        u1412(.A(men_men_n93_), .B(k), .Y(men_men_n1441_));
  AOI210     u1413(.A0(men_men_n1441_), .A1(men_men_n1024_), .B0(men_men_n1146_), .Y(men_men_n1442_));
  NA2        u1414(.A(men_men_n1442_), .B(men_men_n1173_), .Y(men_men_n1443_));
  NO4        u1415(.A(men_men_n1443_), .B(men_men_n1440_), .C(men_men_n1037_), .D(men_men_n1018_), .Y(men_men_n1444_));
  NA4        u1416(.A(men_men_n1444_), .B(men_men_n1082_), .C(men_men_n1071_), .D(men_men_n1059_), .Y(men05));
  INV        u1417(.A(n), .Y(men_men_n1448_));
  INV        u1418(.A(men_men_n436_), .Y(men_men_n1449_));
  INV        u1419(.A(u), .Y(men_men_n1450_));
  INV        u1420(.A(h), .Y(men_men_n1451_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule