library verilog;
use verilog.vl_types.all;
entity ex3_7_vlg_vec_tst is
end ex3_7_vlg_vec_tst;
