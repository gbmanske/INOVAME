// Benchmark "top" written by ABC on Fri Jun 21 17:49:22 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n140_, new_new_n141_, new_new_n142_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n406_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n542_,
    new_new_n543_, new_new_n544_, new_new_n545_, new_new_n546_,
    new_new_n547_, new_new_n548_, new_new_n549_, new_new_n550_,
    new_new_n551_, new_new_n552_, new_new_n553_, new_new_n554_,
    new_new_n555_, new_new_n556_, new_new_n557_, new_new_n558_,
    new_new_n559_, new_new_n560_, new_new_n561_, new_new_n562_,
    new_new_n563_, new_new_n564_, new_new_n565_, new_new_n566_,
    new_new_n567_, new_new_n568_, new_new_n569_, new_new_n570_,
    new_new_n571_, new_new_n572_, new_new_n573_, new_new_n574_,
    new_new_n575_, new_new_n576_, new_new_n577_, new_new_n578_,
    new_new_n579_, new_new_n580_, new_new_n581_, new_new_n582_,
    new_new_n583_, new_new_n584_, new_new_n585_, new_new_n586_,
    new_new_n587_, new_new_n588_, new_new_n589_, new_new_n591_,
    new_new_n592_, new_new_n593_, new_new_n594_, new_new_n595_,
    new_new_n596_, new_new_n597_, new_new_n598_, new_new_n599_,
    new_new_n600_, new_new_n601_, new_new_n602_, new_new_n603_,
    new_new_n604_, new_new_n605_, new_new_n606_, new_new_n607_,
    new_new_n608_, new_new_n609_, new_new_n610_, new_new_n611_,
    new_new_n612_, new_new_n613_, new_new_n614_, new_new_n615_,
    new_new_n616_, new_new_n617_, new_new_n618_, new_new_n619_,
    new_new_n620_, new_new_n621_, new_new_n622_, new_new_n623_,
    new_new_n624_, new_new_n625_, new_new_n626_, new_new_n627_,
    new_new_n628_, new_new_n629_, new_new_n630_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n653_, new_new_n654_, new_new_n655_, new_new_n656_,
    new_new_n657_, new_new_n658_, new_new_n659_, new_new_n660_,
    new_new_n661_, new_new_n662_, new_new_n663_, new_new_n664_,
    new_new_n665_, new_new_n666_, new_new_n667_, new_new_n668_,
    new_new_n669_, new_new_n670_, new_new_n671_, new_new_n672_,
    new_new_n673_, new_new_n674_, new_new_n675_, new_new_n676_,
    new_new_n677_, new_new_n678_, new_new_n679_, new_new_n680_,
    new_new_n681_, new_new_n682_, new_new_n683_, new_new_n684_,
    new_new_n685_, new_new_n686_, new_new_n687_, new_new_n688_,
    new_new_n689_, new_new_n690_, new_new_n691_, new_new_n692_,
    new_new_n693_, new_new_n694_, new_new_n695_, new_new_n696_,
    new_new_n697_, new_new_n698_, new_new_n699_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n703_, new_new_n704_,
    new_new_n705_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n769_, new_new_n770_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g040(.A(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO2        g062(.A(new_new_n83_), .B(new_new_n63_), .Y(new_new_n85_));
  INV        g063(.A(i_6_), .Y(new_new_n86_));
  NO2        g064(.A(i_2_), .B(i_7_), .Y(new_new_n87_));
  INV        g065(.A(new_new_n87_), .Y(new_new_n88_));
  OAI210     g066(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n88_), .Y(new_new_n89_));
  NAi21      g067(.An(i_6_), .B(i_10_), .Y(new_new_n90_));
  NA2        g068(.A(i_6_), .B(i_9_), .Y(new_new_n91_));
  AOI210     g069(.A0(new_new_n91_), .A1(new_new_n90_), .B0(new_new_n63_), .Y(new_new_n92_));
  NA2        g070(.A(i_2_), .B(i_6_), .Y(new_new_n93_));
  NO3        g071(.A(new_new_n93_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n94_));
  NO2        g072(.A(new_new_n94_), .B(new_new_n92_), .Y(new_new_n95_));
  AOI210     g073(.A0(new_new_n95_), .A1(new_new_n89_), .B0(new_new_n80_), .Y(new_new_n96_));
  AN3        g074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n97_));
  NAi21      g075(.An(i_6_), .B(i_11_), .Y(new_new_n98_));
  NO2        g076(.A(i_5_), .B(i_8_), .Y(new_new_n99_));
  NOi21      g077(.An(new_new_n99_), .B(new_new_n98_), .Y(new_new_n100_));
  AOI220     g078(.A0(new_new_n100_), .A1(new_new_n62_), .B0(new_new_n97_), .B1(new_new_n32_), .Y(new_new_n101_));
  INV        g079(.A(i_7_), .Y(new_new_n102_));
  NA2        g080(.A(new_new_n46_), .B(new_new_n102_), .Y(new_new_n103_));
  NO2        g081(.A(i_0_), .B(i_5_), .Y(new_new_n104_));
  NO2        g082(.A(new_new_n104_), .B(new_new_n86_), .Y(new_new_n105_));
  NA2        g083(.A(i_12_), .B(i_3_), .Y(new_new_n106_));
  INV        g084(.A(new_new_n106_), .Y(new_new_n107_));
  NA3        g085(.A(new_new_n107_), .B(new_new_n105_), .C(new_new_n103_), .Y(new_new_n108_));
  NAi21      g086(.An(i_7_), .B(i_11_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n90_), .C(new_new_n53_), .Y(new_new_n110_));
  AN2        g088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g090(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n113_));
  NO2        g091(.A(i_8_), .B(new_new_n102_), .Y(new_new_n114_));
  NO3        g092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(i_0_), .Y(new_new_n118_));
  NA2        g096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  OAI210     g097(.A0(new_new_n118_), .A1(new_new_n116_), .B0(new_new_n119_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(new_new_n115_), .Y(new_new_n121_));
  NAi41      g099(.An(new_new_n110_), .B(new_new_n121_), .C(new_new_n108_), .D(new_new_n101_), .Y(new_new_n122_));
  NOi21      g100(.An(i_1_), .B(i_5_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(i_11_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n125_));
  NA2        g103(.A(i_7_), .B(new_new_n25_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(new_new_n125_), .Y(new_new_n127_));
  NO2        g105(.A(new_new_n127_), .B(new_new_n46_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n91_), .B(new_new_n90_), .Y(new_new_n129_));
  NAi21      g107(.An(i_3_), .B(i_8_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n62_), .Y(new_new_n131_));
  NOi31      g109(.An(new_new_n131_), .B(new_new_n129_), .C(new_new_n128_), .Y(new_new_n132_));
  NO2        g110(.A(i_1_), .B(new_new_n86_), .Y(new_new_n133_));
  NO2        g111(.A(i_6_), .B(i_5_), .Y(new_new_n134_));
  NA2        g112(.A(new_new_n134_), .B(i_3_), .Y(new_new_n135_));
  AO210      g113(.A0(new_new_n135_), .A1(new_new_n47_), .B0(new_new_n133_), .Y(new_new_n136_));
  OAI220     g114(.A0(new_new_n136_), .A1(new_new_n109_), .B0(new_new_n132_), .B1(new_new_n124_), .Y(new_new_n137_));
  NO3        g115(.A(new_new_n137_), .B(new_new_n122_), .C(new_new_n96_), .Y(new_new_n138_));
  NA3        g116(.A(new_new_n138_), .B(new_new_n79_), .C(new_new_n56_), .Y(ori2));
  NO2        g117(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n140_));
  INV        g118(.A(i_6_), .Y(new_new_n141_));
  NA2        g119(.A(new_new_n141_), .B(new_new_n140_), .Y(new_new_n142_));
  NA4        g120(.A(new_new_n142_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(ori0));
  AN2        g121(.A(i_8_), .B(i_7_), .Y(new_new_n144_));
  NA2        g122(.A(new_new_n144_), .B(i_6_), .Y(new_new_n145_));
  NO2        g123(.A(i_12_), .B(i_13_), .Y(new_new_n146_));
  NAi21      g124(.An(i_5_), .B(i_11_), .Y(new_new_n147_));
  NOi21      g125(.An(new_new_n146_), .B(new_new_n147_), .Y(new_new_n148_));
  NO2        g126(.A(i_0_), .B(i_1_), .Y(new_new_n149_));
  NA2        g127(.A(i_2_), .B(i_3_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n150_), .B(i_4_), .Y(new_new_n151_));
  AN2        g129(.A(new_new_n146_), .B(new_new_n83_), .Y(new_new_n152_));
  NA2        g130(.A(i_1_), .B(i_5_), .Y(new_new_n153_));
  OR2        g131(.A(i_0_), .B(i_1_), .Y(new_new_n154_));
  NO3        g132(.A(new_new_n154_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n155_));
  NAi32      g133(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n156_));
  NAi21      g134(.An(new_new_n156_), .B(new_new_n155_), .Y(new_new_n157_));
  NOi21      g135(.An(i_4_), .B(i_10_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n40_), .Y(new_new_n159_));
  NOi21      g137(.An(i_4_), .B(i_9_), .Y(new_new_n160_));
  NOi21      g138(.An(i_11_), .B(i_13_), .Y(new_new_n161_));
  NA2        g139(.A(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  NAi21      g140(.An(i_12_), .B(i_11_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n163_), .B(i_13_), .Y(new_new_n164_));
  NO2        g142(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n165_));
  NO2        g143(.A(new_new_n73_), .B(i_5_), .Y(new_new_n166_));
  NO2        g144(.A(i_13_), .B(i_10_), .Y(new_new_n167_));
  NA3        g145(.A(new_new_n167_), .B(new_new_n166_), .C(new_new_n44_), .Y(new_new_n168_));
  NO2        g146(.A(i_2_), .B(i_1_), .Y(new_new_n169_));
  NAi21      g147(.An(i_4_), .B(i_12_), .Y(new_new_n170_));
  INV        g148(.A(i_8_), .Y(new_new_n171_));
  NO3        g149(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n172_));
  NO2        g150(.A(i_3_), .B(i_8_), .Y(new_new_n173_));
  NO3        g151(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n174_));
  NA3        g152(.A(new_new_n174_), .B(new_new_n173_), .C(new_new_n40_), .Y(new_new_n175_));
  NO2        g153(.A(new_new_n104_), .B(new_new_n58_), .Y(new_new_n176_));
  INV        g154(.A(new_new_n176_), .Y(new_new_n177_));
  NO2        g155(.A(i_13_), .B(i_9_), .Y(new_new_n178_));
  NAi21      g156(.An(i_12_), .B(i_3_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n44_), .B(i_5_), .Y(new_new_n180_));
  NO2        g158(.A(new_new_n177_), .B(new_new_n175_), .Y(new_new_n181_));
  INV        g159(.A(new_new_n181_), .Y(new_new_n182_));
  NO2        g160(.A(new_new_n182_), .B(i_4_), .Y(new_new_n183_));
  NAi21      g161(.An(i_12_), .B(i_7_), .Y(new_new_n184_));
  NA3        g162(.A(i_13_), .B(new_new_n171_), .C(i_10_), .Y(new_new_n185_));
  NA2        g163(.A(i_0_), .B(i_5_), .Y(new_new_n186_));
  NAi31      g164(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n36_), .B(i_13_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n190_));
  INV        g168(.A(i_13_), .Y(new_new_n191_));
  NO2        g169(.A(i_12_), .B(new_new_n191_), .Y(new_new_n192_));
  NO2        g170(.A(i_12_), .B(new_new_n37_), .Y(new_new_n193_));
  OR2        g171(.A(i_8_), .B(i_7_), .Y(new_new_n194_));
  INV        g172(.A(i_12_), .Y(new_new_n195_));
  NO2        g173(.A(new_new_n44_), .B(new_new_n195_), .Y(new_new_n196_));
  NO3        g174(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n197_));
  NA2        g175(.A(i_2_), .B(i_1_), .Y(new_new_n198_));
  NO3        g176(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n199_));
  NAi21      g177(.An(i_4_), .B(i_3_), .Y(new_new_n200_));
  NO2        g178(.A(i_0_), .B(i_6_), .Y(new_new_n201_));
  NOi41      g179(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n202_));
  NA2        g180(.A(new_new_n202_), .B(new_new_n201_), .Y(new_new_n203_));
  NO2        g181(.A(i_11_), .B(new_new_n191_), .Y(new_new_n204_));
  NOi21      g182(.An(i_1_), .B(i_6_), .Y(new_new_n205_));
  NAi21      g183(.An(i_3_), .B(i_7_), .Y(new_new_n206_));
  NA2        g184(.A(new_new_n195_), .B(i_9_), .Y(new_new_n207_));
  OR4        g185(.A(new_new_n207_), .B(new_new_n206_), .C(new_new_n205_), .D(new_new_n166_), .Y(new_new_n208_));
  NA2        g186(.A(new_new_n73_), .B(i_5_), .Y(new_new_n209_));
  NA2        g187(.A(i_3_), .B(i_9_), .Y(new_new_n210_));
  NAi21      g188(.An(i_7_), .B(i_10_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n211_), .B(new_new_n210_), .Y(new_new_n212_));
  NA3        g190(.A(new_new_n212_), .B(new_new_n209_), .C(new_new_n64_), .Y(new_new_n213_));
  NA2        g191(.A(new_new_n213_), .B(new_new_n208_), .Y(new_new_n214_));
  INV        g192(.A(new_new_n145_), .Y(new_new_n215_));
  NA2        g193(.A(new_new_n195_), .B(i_13_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n216_), .B(new_new_n75_), .Y(new_new_n217_));
  AOI220     g195(.A0(new_new_n217_), .A1(new_new_n215_), .B0(new_new_n214_), .B1(new_new_n204_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n194_), .B(new_new_n37_), .Y(new_new_n219_));
  NA2        g197(.A(i_12_), .B(i_6_), .Y(new_new_n220_));
  OR2        g198(.A(i_13_), .B(i_9_), .Y(new_new_n221_));
  NO3        g199(.A(new_new_n221_), .B(new_new_n220_), .C(new_new_n48_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n200_), .B(i_2_), .Y(new_new_n223_));
  NA3        g201(.A(new_new_n223_), .B(new_new_n222_), .C(new_new_n44_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n204_), .B(i_9_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n209_), .B(new_new_n64_), .Y(new_new_n226_));
  OAI210     g204(.A0(new_new_n226_), .A1(new_new_n225_), .B0(new_new_n224_), .Y(new_new_n227_));
  NO3        g205(.A(i_11_), .B(new_new_n191_), .C(new_new_n25_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n206_), .B(i_8_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n227_), .B(new_new_n219_), .Y(new_new_n230_));
  NA2        g208(.A(new_new_n230_), .B(new_new_n218_), .Y(new_new_n231_));
  NO3        g209(.A(i_12_), .B(new_new_n191_), .C(new_new_n37_), .Y(new_new_n232_));
  NO2        g210(.A(i_2_), .B(new_new_n102_), .Y(new_new_n233_));
  AN2        g211(.A(i_3_), .B(i_10_), .Y(new_new_n234_));
  NO2        g212(.A(i_5_), .B(new_new_n37_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n236_));
  NO2        g214(.A(new_new_n231_), .B(new_new_n183_), .Y(new_new_n237_));
  NO3        g215(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n238_));
  NO2        g216(.A(i_2_), .B(i_3_), .Y(new_new_n239_));
  OR2        g217(.A(i_0_), .B(i_5_), .Y(new_new_n240_));
  NO2        g218(.A(i_12_), .B(i_10_), .Y(new_new_n241_));
  NOi21      g219(.An(i_5_), .B(i_0_), .Y(new_new_n242_));
  NA4        g220(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n243_));
  NO2        g221(.A(i_1_), .B(i_7_), .Y(new_new_n244_));
  NOi21      g222(.An(new_new_n153_), .B(new_new_n105_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n245_), .B(new_new_n126_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n246_), .B(i_3_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n171_), .B(i_9_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n248_), .B(new_new_n176_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n249_), .B(new_new_n46_), .Y(new_new_n250_));
  INV        g228(.A(new_new_n250_), .Y(new_new_n251_));
  AOI210     g229(.A0(new_new_n251_), .A1(new_new_n247_), .B0(new_new_n159_), .Y(new_new_n252_));
  INV        g230(.A(new_new_n252_), .Y(new_new_n253_));
  NOi32      g231(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n254_));
  INV        g232(.A(new_new_n254_), .Y(new_new_n255_));
  INV        g233(.A(new_new_n203_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n187_), .B(new_new_n156_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n156_), .B(new_new_n154_), .Y(new_new_n258_));
  NOi32      g236(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n259_));
  NAi21      g237(.An(i_6_), .B(i_1_), .Y(new_new_n260_));
  NA3        g238(.A(new_new_n260_), .B(new_new_n259_), .C(new_new_n46_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n261_), .B(i_0_), .Y(new_new_n262_));
  OR3        g240(.A(new_new_n262_), .B(new_new_n258_), .C(new_new_n257_), .Y(new_new_n263_));
  NO2        g241(.A(i_1_), .B(new_new_n102_), .Y(new_new_n264_));
  NAi21      g242(.An(i_3_), .B(i_4_), .Y(new_new_n265_));
  NO2        g243(.A(new_new_n265_), .B(i_9_), .Y(new_new_n266_));
  AN2        g244(.A(i_6_), .B(i_7_), .Y(new_new_n267_));
  OAI210     g245(.A0(new_new_n267_), .A1(new_new_n264_), .B0(new_new_n266_), .Y(new_new_n268_));
  NA2        g246(.A(i_2_), .B(i_7_), .Y(new_new_n269_));
  NO2        g247(.A(new_new_n265_), .B(i_10_), .Y(new_new_n270_));
  NA3        g248(.A(new_new_n270_), .B(new_new_n269_), .C(new_new_n201_), .Y(new_new_n271_));
  AOI210     g249(.A0(new_new_n271_), .A1(new_new_n268_), .B0(new_new_n166_), .Y(new_new_n272_));
  AOI210     g250(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n273_));
  OAI210     g251(.A0(new_new_n273_), .A1(new_new_n169_), .B0(new_new_n270_), .Y(new_new_n274_));
  AOI220     g252(.A0(new_new_n270_), .A1(new_new_n244_), .B0(new_new_n197_), .B1(new_new_n169_), .Y(new_new_n275_));
  AOI210     g253(.A0(new_new_n275_), .A1(new_new_n274_), .B0(i_5_), .Y(new_new_n276_));
  NO4        g254(.A(new_new_n276_), .B(new_new_n272_), .C(new_new_n263_), .D(new_new_n256_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n277_), .B(new_new_n255_), .Y(new_new_n278_));
  AN2        g256(.A(i_12_), .B(i_5_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n770_), .B(new_new_n279_), .Y(new_new_n280_));
  NO2        g258(.A(i_11_), .B(i_6_), .Y(new_new_n281_));
  NO2        g259(.A(i_5_), .B(i_10_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n283_));
  NO3        g261(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n284_));
  NO2        g262(.A(i_11_), .B(i_12_), .Y(new_new_n285_));
  NAi21      g263(.An(i_13_), .B(i_0_), .Y(new_new_n286_));
  NO3        g264(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n287_));
  NO2        g265(.A(i_0_), .B(i_11_), .Y(new_new_n288_));
  AN2        g266(.A(i_1_), .B(i_6_), .Y(new_new_n289_));
  NOi21      g267(.An(i_2_), .B(i_12_), .Y(new_new_n290_));
  NAi21      g268(.An(i_9_), .B(i_4_), .Y(new_new_n291_));
  OR2        g269(.A(i_13_), .B(i_10_), .Y(new_new_n292_));
  NO3        g270(.A(new_new_n292_), .B(new_new_n119_), .C(new_new_n291_), .Y(new_new_n293_));
  NO2        g271(.A(new_new_n162_), .B(new_new_n125_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n102_), .B(new_new_n25_), .Y(new_new_n295_));
  NA2        g273(.A(new_new_n232_), .B(new_new_n295_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n296_), .B(new_new_n245_), .Y(new_new_n297_));
  INV        g275(.A(new_new_n297_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n298_), .B(new_new_n26_), .Y(new_new_n299_));
  NA2        g277(.A(new_new_n171_), .B(i_10_), .Y(new_new_n300_));
  NA3        g278(.A(new_new_n209_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n301_), .B(new_new_n300_), .Y(new_new_n302_));
  INV        g280(.A(new_new_n302_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n303_), .B(new_new_n225_), .Y(new_new_n304_));
  NO3        g282(.A(new_new_n304_), .B(new_new_n299_), .C(new_new_n278_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n73_), .B(i_13_), .Y(new_new_n306_));
  NO2        g284(.A(i_10_), .B(i_9_), .Y(new_new_n307_));
  NAi21      g285(.An(i_12_), .B(i_8_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n308_), .B(i_3_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n236_), .B(i_0_), .Y(new_new_n310_));
  NO3        g288(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n311_));
  NA2        g289(.A(new_new_n220_), .B(new_new_n98_), .Y(new_new_n312_));
  NA2        g290(.A(new_new_n312_), .B(new_new_n311_), .Y(new_new_n313_));
  NA2        g291(.A(i_8_), .B(i_9_), .Y(new_new_n314_));
  AOI210     g292(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n315_));
  OR2        g293(.A(new_new_n315_), .B(new_new_n314_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n232_), .B(new_new_n176_), .Y(new_new_n317_));
  OAI220     g295(.A0(new_new_n317_), .A1(new_new_n316_), .B0(new_new_n313_), .B1(new_new_n310_), .Y(new_new_n318_));
  NA2        g296(.A(new_new_n204_), .B(new_new_n235_), .Y(new_new_n319_));
  NO3        g297(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n320_));
  INV        g298(.A(new_new_n320_), .Y(new_new_n321_));
  NA3        g299(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n322_));
  NA4        g300(.A(new_new_n147_), .B(new_new_n117_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n323_));
  OAI220     g301(.A0(new_new_n323_), .A1(new_new_n322_), .B0(new_new_n321_), .B1(new_new_n319_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n324_), .B(new_new_n318_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n97_), .B(i_13_), .Y(new_new_n326_));
  NO2        g304(.A(i_2_), .B(i_13_), .Y(new_new_n327_));
  NO3        g305(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n328_));
  NO2        g306(.A(i_6_), .B(i_7_), .Y(new_new_n329_));
  NO2        g307(.A(i_11_), .B(i_1_), .Y(new_new_n330_));
  NOi21      g308(.An(i_2_), .B(i_7_), .Y(new_new_n331_));
  NO2        g309(.A(i_3_), .B(new_new_n171_), .Y(new_new_n332_));
  NO2        g310(.A(i_6_), .B(i_10_), .Y(new_new_n333_));
  NA3        g311(.A(new_new_n202_), .B(new_new_n161_), .C(new_new_n134_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n154_), .B(i_3_), .Y(new_new_n336_));
  NAi31      g314(.An(new_new_n335_), .B(new_new_n336_), .C(new_new_n192_), .Y(new_new_n337_));
  NA3        g315(.A(new_new_n283_), .B(new_new_n165_), .C(new_new_n151_), .Y(new_new_n338_));
  NA3        g316(.A(new_new_n338_), .B(new_new_n337_), .C(new_new_n334_), .Y(new_new_n339_));
  INV        g317(.A(new_new_n339_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n311_), .B(new_new_n279_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n320_), .B(new_new_n282_), .Y(new_new_n342_));
  NAi21      g320(.An(new_new_n185_), .B(new_new_n285_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n244_), .B(new_new_n186_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n344_), .B(new_new_n343_), .Y(new_new_n345_));
  NA2        g323(.A(new_new_n27_), .B(i_10_), .Y(new_new_n346_));
  NA2        g324(.A(new_new_n238_), .B(new_new_n197_), .Y(new_new_n347_));
  OAI220     g325(.A0(new_new_n347_), .A1(new_new_n301_), .B0(new_new_n346_), .B1(new_new_n326_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(new_new_n345_), .Y(new_new_n349_));
  NA3        g327(.A(new_new_n349_), .B(new_new_n340_), .C(new_new_n325_), .Y(new_new_n350_));
  NA2        g328(.A(new_new_n279_), .B(new_new_n191_), .Y(new_new_n351_));
  NA2        g329(.A(new_new_n267_), .B(new_new_n259_), .Y(new_new_n352_));
  OR2        g330(.A(new_new_n351_), .B(new_new_n352_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n36_), .B(i_8_), .Y(new_new_n354_));
  AOI210     g332(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n293_), .Y(new_new_n355_));
  NA2        g333(.A(new_new_n355_), .B(new_new_n353_), .Y(new_new_n356_));
  INV        g334(.A(new_new_n356_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n209_), .B(new_new_n64_), .Y(new_new_n358_));
  OAI210     g336(.A0(i_8_), .A1(new_new_n358_), .B0(new_new_n136_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n359_), .B(new_new_n294_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n360_), .B(new_new_n357_), .Y(new_new_n361_));
  NO2        g339(.A(i_12_), .B(new_new_n171_), .Y(new_new_n362_));
  NA2        g340(.A(new_new_n44_), .B(i_10_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n363_), .B(i_6_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n154_), .B(i_5_), .Y(new_new_n365_));
  NA3        g343(.A(new_new_n186_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n366_));
  NA2        g344(.A(new_new_n232_), .B(new_new_n84_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n366_), .B(new_new_n367_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n190_), .B(new_new_n189_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n307_), .B(new_new_n188_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n369_), .B(new_new_n370_), .Y(new_new_n371_));
  AOI210     g349(.A0(new_new_n260_), .A1(new_new_n46_), .B0(new_new_n264_), .Y(new_new_n372_));
  NA2        g350(.A(i_0_), .B(new_new_n48_), .Y(new_new_n373_));
  NA3        g351(.A(new_new_n362_), .B(new_new_n228_), .C(new_new_n373_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n372_), .B(new_new_n374_), .Y(new_new_n375_));
  NO3        g353(.A(new_new_n375_), .B(new_new_n371_), .C(new_new_n368_), .Y(new_new_n376_));
  NO4        g354(.A(new_new_n205_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n377_));
  NO3        g355(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n292_), .B(i_1_), .Y(new_new_n379_));
  NOi31      g357(.An(new_new_n379_), .B(new_new_n312_), .C(new_new_n73_), .Y(new_new_n380_));
  NOi21      g358(.An(i_10_), .B(i_6_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n382_));
  AOI220     g360(.A0(new_new_n232_), .A1(new_new_n382_), .B0(new_new_n228_), .B1(new_new_n381_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n310_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n385_));
  NOi31      g363(.An(new_new_n148_), .B(i_10_), .C(new_new_n243_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n386_), .B(new_new_n384_), .Y(new_new_n387_));
  INV        g365(.A(new_new_n239_), .Y(new_new_n388_));
  NO2        g366(.A(i_12_), .B(new_new_n86_), .Y(new_new_n389_));
  NA3        g367(.A(new_new_n389_), .B(new_new_n228_), .C(new_new_n373_), .Y(new_new_n390_));
  NA3        g368(.A(new_new_n281_), .B(new_new_n232_), .C(new_new_n186_), .Y(new_new_n391_));
  AOI210     g369(.A0(new_new_n391_), .A1(new_new_n390_), .B0(new_new_n388_), .Y(new_new_n392_));
  OR2        g370(.A(i_2_), .B(i_5_), .Y(new_new_n393_));
  OR2        g371(.A(new_new_n393_), .B(new_new_n289_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n269_), .B(new_new_n201_), .Y(new_new_n395_));
  AOI210     g373(.A0(new_new_n395_), .A1(new_new_n394_), .B0(new_new_n343_), .Y(new_new_n396_));
  NO2        g374(.A(new_new_n396_), .B(new_new_n392_), .Y(new_new_n397_));
  NA3        g375(.A(new_new_n397_), .B(new_new_n387_), .C(new_new_n376_), .Y(new_new_n398_));
  NO3        g376(.A(new_new_n398_), .B(new_new_n361_), .C(new_new_n350_), .Y(new_new_n399_));
  NA4        g377(.A(new_new_n399_), .B(new_new_n305_), .C(new_new_n253_), .D(new_new_n237_), .Y(ori7));
  NO2        g378(.A(new_new_n93_), .B(new_new_n54_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n109_), .B(new_new_n90_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n770_), .B(new_new_n402_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n333_), .B(new_new_n84_), .Y(new_new_n404_));
  NA2        g382(.A(i_11_), .B(new_new_n171_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n146_), .B(new_new_n405_), .Y(new_new_n406_));
  OAI210     g384(.A0(new_new_n406_), .A1(new_new_n404_), .B0(new_new_n403_), .Y(new_new_n407_));
  NA3        g385(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n195_), .B(i_4_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n409_), .B(i_8_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n106_), .B(new_new_n408_), .Y(new_new_n411_));
  NA2        g389(.A(i_2_), .B(new_new_n86_), .Y(new_new_n412_));
  OAI210     g390(.A0(new_new_n87_), .A1(new_new_n173_), .B0(new_new_n174_), .Y(new_new_n413_));
  NO2        g391(.A(i_7_), .B(new_new_n37_), .Y(new_new_n414_));
  NA2        g392(.A(i_4_), .B(i_8_), .Y(new_new_n415_));
  AOI210     g393(.A0(new_new_n415_), .A1(new_new_n234_), .B0(new_new_n414_), .Y(new_new_n416_));
  OAI220     g394(.A0(new_new_n416_), .A1(new_new_n412_), .B0(new_new_n413_), .B1(i_13_), .Y(new_new_n417_));
  NO4        g395(.A(new_new_n417_), .B(new_new_n411_), .C(new_new_n407_), .D(new_new_n401_), .Y(new_new_n418_));
  AOI210     g396(.A0(new_new_n130_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n419_));
  AOI210     g397(.A0(new_new_n419_), .A1(new_new_n195_), .B0(new_new_n158_), .Y(new_new_n420_));
  OR2        g398(.A(i_6_), .B(i_10_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n421_), .B(new_new_n23_), .Y(new_new_n422_));
  OR3        g400(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n423_));
  INV        g401(.A(new_new_n172_), .Y(new_new_n424_));
  INV        g402(.A(new_new_n422_), .Y(new_new_n425_));
  OA220      g403(.A0(new_new_n425_), .A1(new_new_n388_), .B0(new_new_n420_), .B1(new_new_n221_), .Y(new_new_n426_));
  AOI210     g404(.A0(new_new_n426_), .A1(new_new_n418_), .B0(new_new_n63_), .Y(new_new_n427_));
  NOi21      g405(.An(i_11_), .B(i_7_), .Y(new_new_n428_));
  AO210      g406(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n429_));
  NO2        g407(.A(new_new_n429_), .B(new_new_n428_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n430_), .B(new_new_n178_), .Y(new_new_n431_));
  NA3        g409(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n431_), .B(new_new_n63_), .Y(new_new_n433_));
  OR2        g411(.A(new_new_n275_), .B(new_new_n41_), .Y(new_new_n434_));
  NO3        g412(.A(new_new_n211_), .B(new_new_n179_), .C(new_new_n405_), .Y(new_new_n435_));
  OAI210     g413(.A0(new_new_n435_), .A1(new_new_n192_), .B0(new_new_n63_), .Y(new_new_n436_));
  NA2        g414(.A(new_new_n290_), .B(new_new_n31_), .Y(new_new_n437_));
  OR2        g415(.A(new_new_n179_), .B(new_new_n109_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n438_), .B(new_new_n437_), .Y(new_new_n439_));
  NO2        g417(.A(i_1_), .B(i_4_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n440_), .B(new_new_n439_), .Y(new_new_n441_));
  NO2        g419(.A(i_1_), .B(i_12_), .Y(new_new_n442_));
  NA3        g420(.A(new_new_n442_), .B(new_new_n111_), .C(new_new_n24_), .Y(new_new_n443_));
  BUFFER     g421(.A(new_new_n443_), .Y(new_new_n444_));
  NA4        g422(.A(new_new_n444_), .B(new_new_n441_), .C(new_new_n436_), .D(new_new_n434_), .Y(new_new_n445_));
  OAI210     g423(.A0(new_new_n445_), .A1(new_new_n433_), .B0(i_6_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n432_), .B(new_new_n109_), .Y(new_new_n447_));
  NA2        g425(.A(new_new_n447_), .B(new_new_n389_), .Y(new_new_n448_));
  NO2        g426(.A(i_6_), .B(i_11_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n448_), .B(new_new_n313_), .Y(new_new_n450_));
  NO3        g428(.A(new_new_n421_), .B(new_new_n194_), .C(new_new_n23_), .Y(new_new_n451_));
  AOI210     g429(.A0(i_1_), .A1(new_new_n212_), .B0(new_new_n451_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n452_), .B(new_new_n44_), .Y(new_new_n453_));
  INV        g431(.A(i_2_), .Y(new_new_n454_));
  NA2        g432(.A(new_new_n140_), .B(i_9_), .Y(new_new_n455_));
  NA3        g433(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n46_), .B(i_1_), .Y(new_new_n457_));
  NA3        g435(.A(new_new_n457_), .B(new_new_n220_), .C(new_new_n44_), .Y(new_new_n458_));
  OAI220     g436(.A0(new_new_n458_), .A1(new_new_n456_), .B0(new_new_n455_), .B1(new_new_n454_), .Y(new_new_n459_));
  AOI210     g437(.A0(new_new_n330_), .A1(new_new_n295_), .B0(new_new_n199_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n460_), .B(new_new_n412_), .Y(new_new_n461_));
  NO2        g439(.A(i_11_), .B(new_new_n37_), .Y(new_new_n462_));
  OR2        g440(.A(new_new_n461_), .B(new_new_n459_), .Y(new_new_n463_));
  NO3        g441(.A(new_new_n463_), .B(new_new_n453_), .C(new_new_n450_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n195_), .B(new_new_n102_), .Y(new_new_n465_));
  NO2        g443(.A(new_new_n465_), .B(new_new_n428_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n466_), .B(i_1_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n467_), .B(new_new_n423_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n291_), .B(new_new_n86_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n468_), .B(new_new_n46_), .Y(new_new_n470_));
  NA2        g448(.A(i_3_), .B(new_new_n171_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n471_), .B(new_new_n116_), .Y(new_new_n472_));
  AN2        g450(.A(new_new_n472_), .B(new_new_n364_), .Y(new_new_n473_));
  NO2        g451(.A(new_new_n194_), .B(new_new_n44_), .Y(new_new_n474_));
  NO3        g452(.A(new_new_n474_), .B(new_new_n236_), .C(new_new_n196_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n119_), .B(new_new_n37_), .Y(new_new_n476_));
  NO2        g454(.A(new_new_n476_), .B(i_6_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n86_), .B(i_9_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n478_), .B(new_new_n63_), .Y(new_new_n479_));
  NO2        g457(.A(new_new_n479_), .B(new_new_n442_), .Y(new_new_n480_));
  NO4        g458(.A(new_new_n480_), .B(new_new_n477_), .C(new_new_n475_), .D(i_4_), .Y(new_new_n481_));
  NA2        g459(.A(i_1_), .B(i_3_), .Y(new_new_n482_));
  NO2        g460(.A(new_new_n314_), .B(new_new_n93_), .Y(new_new_n483_));
  AOI210     g461(.A0(new_new_n474_), .A1(new_new_n381_), .B0(new_new_n483_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n484_), .B(new_new_n482_), .Y(new_new_n485_));
  NO3        g463(.A(new_new_n485_), .B(new_new_n481_), .C(new_new_n473_), .Y(new_new_n486_));
  NA4        g464(.A(new_new_n486_), .B(new_new_n470_), .C(new_new_n464_), .D(new_new_n446_), .Y(new_new_n487_));
  AN2        g465(.A(new_new_n202_), .B(new_new_n86_), .Y(new_new_n488_));
  NA2        g466(.A(new_new_n267_), .B(new_new_n266_), .Y(new_new_n489_));
  NO3        g467(.A(new_new_n331_), .B(new_new_n415_), .C(new_new_n86_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n490_), .B(new_new_n25_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n491_), .B(new_new_n489_), .Y(new_new_n492_));
  OAI210     g470(.A0(new_new_n492_), .A1(new_new_n488_), .B0(i_1_), .Y(new_new_n493_));
  AOI210     g471(.A0(new_new_n220_), .A1(new_new_n98_), .B0(i_1_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n265_), .B(i_2_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n495_), .B(new_new_n494_), .Y(new_new_n496_));
  AOI210     g474(.A0(new_new_n496_), .A1(new_new_n493_), .B0(i_13_), .Y(new_new_n497_));
  OR2        g475(.A(i_11_), .B(i_7_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n54_), .B(i_12_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n331_), .B(new_new_n24_), .Y(new_new_n500_));
  AOI220     g478(.A0(new_new_n500_), .A1(new_new_n469_), .B0(new_new_n202_), .B1(new_new_n133_), .Y(new_new_n501_));
  OAI220     g479(.A0(new_new_n501_), .A1(new_new_n41_), .B0(new_new_n769_), .B1(new_new_n93_), .Y(new_new_n502_));
  INV        g480(.A(new_new_n502_), .Y(new_new_n503_));
  INV        g481(.A(new_new_n116_), .Y(new_new_n504_));
  AOI220     g482(.A0(new_new_n504_), .A1(new_new_n72_), .B0(new_new_n281_), .B1(new_new_n457_), .Y(new_new_n505_));
  NO2        g483(.A(new_new_n505_), .B(new_new_n200_), .Y(new_new_n506_));
  AOI210     g484(.A0(new_new_n308_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n507_));
  NOi31      g485(.An(new_new_n507_), .B(new_new_n404_), .C(new_new_n44_), .Y(new_new_n508_));
  NA2        g486(.A(new_new_n129_), .B(i_13_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n456_), .B(new_new_n116_), .Y(new_new_n510_));
  INV        g488(.A(new_new_n510_), .Y(new_new_n511_));
  OAI220     g489(.A0(new_new_n511_), .A1(new_new_n71_), .B0(new_new_n509_), .B1(new_new_n494_), .Y(new_new_n512_));
  NO3        g490(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n102_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n26_), .B(new_new_n171_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n514_), .B(i_7_), .Y(new_new_n515_));
  NO3        g493(.A(new_new_n331_), .B(new_new_n195_), .C(new_new_n86_), .Y(new_new_n516_));
  AOI210     g494(.A0(new_new_n516_), .A1(new_new_n515_), .B0(new_new_n513_), .Y(new_new_n517_));
  AOI220     g495(.A0(new_new_n281_), .A1(new_new_n457_), .B0(new_new_n92_), .B1(new_new_n103_), .Y(new_new_n518_));
  OAI220     g496(.A0(new_new_n518_), .A1(new_new_n410_), .B0(new_new_n517_), .B1(new_new_n424_), .Y(new_new_n519_));
  NO4        g497(.A(new_new_n519_), .B(new_new_n512_), .C(new_new_n508_), .D(new_new_n506_), .Y(new_new_n520_));
  OR2        g498(.A(i_11_), .B(i_6_), .Y(new_new_n521_));
  NA3        g499(.A(new_new_n409_), .B(new_new_n514_), .C(i_7_), .Y(new_new_n522_));
  AOI210     g500(.A0(new_new_n522_), .A1(new_new_n511_), .B0(new_new_n521_), .Y(new_new_n523_));
  NA3        g501(.A(new_new_n290_), .B(new_new_n414_), .C(new_new_n98_), .Y(new_new_n524_));
  NA2        g502(.A(new_new_n449_), .B(i_13_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n103_), .B(new_new_n514_), .Y(new_new_n526_));
  NAi21      g504(.An(i_11_), .B(i_12_), .Y(new_new_n527_));
  NOi41      g505(.An(new_new_n112_), .B(new_new_n527_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n528_));
  NO3        g506(.A(new_new_n331_), .B(new_new_n389_), .C(new_new_n415_), .Y(new_new_n529_));
  AOI220     g507(.A0(new_new_n529_), .A1(new_new_n238_), .B0(new_new_n528_), .B1(new_new_n526_), .Y(new_new_n530_));
  NA3        g508(.A(new_new_n530_), .B(new_new_n525_), .C(new_new_n524_), .Y(new_new_n531_));
  OAI210     g509(.A0(new_new_n531_), .A1(new_new_n523_), .B0(new_new_n63_), .Y(new_new_n532_));
  NO2        g510(.A(i_2_), .B(i_12_), .Y(new_new_n533_));
  NA2        g511(.A(new_new_n264_), .B(new_new_n533_), .Y(new_new_n534_));
  NA2        g512(.A(new_new_n266_), .B(new_new_n264_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n130_), .B(i_2_), .Y(new_new_n536_));
  NA2        g514(.A(new_new_n536_), .B(new_new_n442_), .Y(new_new_n537_));
  NA3        g515(.A(new_new_n537_), .B(new_new_n535_), .C(new_new_n534_), .Y(new_new_n538_));
  NA3        g516(.A(new_new_n538_), .B(new_new_n45_), .C(new_new_n191_), .Y(new_new_n539_));
  NA4        g517(.A(new_new_n539_), .B(new_new_n532_), .C(new_new_n520_), .D(new_new_n503_), .Y(new_new_n540_));
  OR4        g518(.A(new_new_n540_), .B(new_new_n497_), .C(new_new_n487_), .D(new_new_n427_), .Y(ori5));
  NA2        g519(.A(new_new_n466_), .B(new_new_n223_), .Y(new_new_n542_));
  AN2        g520(.A(new_new_n24_), .B(i_10_), .Y(new_new_n543_));
  NA3        g521(.A(new_new_n543_), .B(new_new_n533_), .C(new_new_n109_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n410_), .B(i_11_), .Y(new_new_n545_));
  NA2        g523(.A(new_new_n87_), .B(new_new_n545_), .Y(new_new_n546_));
  NA3        g524(.A(new_new_n546_), .B(new_new_n544_), .C(new_new_n542_), .Y(new_new_n547_));
  NO3        g525(.A(i_11_), .B(new_new_n195_), .C(i_13_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n126_), .B(new_new_n23_), .Y(new_new_n549_));
  NA2        g527(.A(i_12_), .B(i_8_), .Y(new_new_n550_));
  OAI210     g528(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n550_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n307_), .Y(new_new_n552_));
  AOI220     g530(.A0(new_new_n239_), .A1(new_new_n385_), .B0(new_new_n551_), .B1(new_new_n549_), .Y(new_new_n553_));
  INV        g531(.A(new_new_n553_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n554_), .B(new_new_n547_), .Y(new_new_n555_));
  INV        g533(.A(new_new_n161_), .Y(new_new_n556_));
  INV        g534(.A(new_new_n202_), .Y(new_new_n557_));
  OAI210     g535(.A0(new_new_n495_), .A1(new_new_n309_), .B0(new_new_n112_), .Y(new_new_n558_));
  AOI210     g536(.A0(new_new_n558_), .A1(new_new_n557_), .B0(new_new_n556_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n314_), .B(new_new_n26_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n560_), .B(new_new_n295_), .Y(new_new_n561_));
  NA2        g539(.A(new_new_n561_), .B(i_2_), .Y(new_new_n562_));
  INV        g540(.A(new_new_n562_), .Y(new_new_n563_));
  AOI210     g541(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n292_), .Y(new_new_n564_));
  AOI210     g542(.A0(new_new_n564_), .A1(new_new_n563_), .B0(new_new_n559_), .Y(new_new_n565_));
  NO2        g543(.A(new_new_n170_), .B(new_new_n127_), .Y(new_new_n566_));
  OAI210     g544(.A0(new_new_n566_), .A1(new_new_n549_), .B0(i_2_), .Y(new_new_n567_));
  INV        g545(.A(new_new_n162_), .Y(new_new_n568_));
  NO3        g546(.A(new_new_n429_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n569_));
  AOI210     g547(.A0(new_new_n568_), .A1(new_new_n87_), .B0(new_new_n569_), .Y(new_new_n570_));
  AOI210     g548(.A0(new_new_n570_), .A1(new_new_n567_), .B0(new_new_n171_), .Y(new_new_n571_));
  OA210      g549(.A0(new_new_n430_), .A1(new_new_n128_), .B0(i_13_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n172_), .B(new_new_n173_), .Y(new_new_n573_));
  NA2        g551(.A(new_new_n152_), .B(new_new_n405_), .Y(new_new_n574_));
  AOI210     g552(.A0(new_new_n574_), .A1(new_new_n573_), .B0(new_new_n269_), .Y(new_new_n575_));
  AOI210     g553(.A0(new_new_n179_), .A1(new_new_n150_), .B0(new_new_n354_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n576_), .B(new_new_n295_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n103_), .B(new_new_n44_), .Y(new_new_n578_));
  INV        g556(.A(new_new_n233_), .Y(new_new_n579_));
  NA4        g557(.A(new_new_n579_), .B(new_new_n234_), .C(new_new_n126_), .D(new_new_n42_), .Y(new_new_n580_));
  OAI210     g558(.A0(new_new_n580_), .A1(new_new_n578_), .B0(new_new_n577_), .Y(new_new_n581_));
  NO4        g559(.A(new_new_n581_), .B(new_new_n575_), .C(new_new_n572_), .D(new_new_n571_), .Y(new_new_n582_));
  NA2        g560(.A(new_new_n385_), .B(new_new_n28_), .Y(new_new_n583_));
  NA2        g561(.A(new_new_n548_), .B(new_new_n229_), .Y(new_new_n584_));
  NA2        g562(.A(new_new_n584_), .B(new_new_n583_), .Y(new_new_n585_));
  NO2        g563(.A(new_new_n62_), .B(i_12_), .Y(new_new_n586_));
  NO2        g564(.A(new_new_n586_), .B(new_new_n128_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n587_), .B(new_new_n405_), .Y(new_new_n588_));
  AOI220     g566(.A0(new_new_n588_), .A1(new_new_n36_), .B0(new_new_n585_), .B1(new_new_n46_), .Y(new_new_n589_));
  NA4        g567(.A(new_new_n589_), .B(new_new_n582_), .C(new_new_n565_), .D(new_new_n555_), .Y(ori6));
  NA4        g568(.A(new_new_n282_), .B(new_new_n332_), .C(new_new_n71_), .D(new_new_n102_), .Y(new_new_n591_));
  INV        g569(.A(new_new_n591_), .Y(new_new_n592_));
  NO2        g570(.A(new_new_n187_), .B(new_new_n335_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n592_), .B(new_new_n242_), .Y(new_new_n594_));
  OR2        g572(.A(new_new_n594_), .B(i_12_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n389_), .B(new_new_n63_), .Y(new_new_n596_));
  INV        g574(.A(new_new_n596_), .Y(new_new_n597_));
  NA2        g575(.A(new_new_n597_), .B(new_new_n73_), .Y(new_new_n598_));
  INV        g576(.A(new_new_n241_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n75_), .B(new_new_n133_), .Y(new_new_n600_));
  INV        g578(.A(new_new_n126_), .Y(new_new_n601_));
  NA2        g579(.A(new_new_n601_), .B(new_new_n46_), .Y(new_new_n602_));
  AOI210     g580(.A0(new_new_n602_), .A1(new_new_n600_), .B0(new_new_n599_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n205_), .B(i_9_), .Y(new_new_n604_));
  NA2        g582(.A(new_new_n604_), .B(new_new_n586_), .Y(new_new_n605_));
  AOI210     g583(.A0(new_new_n605_), .A1(new_new_n352_), .B0(new_new_n166_), .Y(new_new_n606_));
  NO2        g584(.A(new_new_n32_), .B(i_11_), .Y(new_new_n607_));
  NAi32      g585(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n521_), .B(new_new_n608_), .Y(new_new_n609_));
  OR3        g587(.A(new_new_n609_), .B(new_new_n606_), .C(new_new_n603_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n498_), .B(i_2_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n612_), .B(new_new_n289_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n613_), .B(new_new_n611_), .Y(new_new_n614_));
  OR2        g592(.A(new_new_n430_), .B(new_new_n309_), .Y(new_new_n615_));
  NA3        g593(.A(new_new_n615_), .B(new_new_n149_), .C(new_new_n69_), .Y(new_new_n616_));
  AO210      g594(.A0(new_new_n342_), .A1(new_new_n552_), .B0(new_new_n36_), .Y(new_new_n617_));
  NA3        g595(.A(new_new_n617_), .B(new_new_n616_), .C(new_new_n614_), .Y(new_new_n618_));
  NO2        g596(.A(i_6_), .B(i_11_), .Y(new_new_n619_));
  AOI220     g597(.A0(new_new_n619_), .A1(new_new_n378_), .B0(new_new_n593_), .B1(new_new_n515_), .Y(new_new_n620_));
  NA3        g598(.A(new_new_n269_), .B(new_new_n197_), .C(new_new_n149_), .Y(new_new_n621_));
  NA2        g599(.A(new_new_n284_), .B(new_new_n70_), .Y(new_new_n622_));
  NA4        g600(.A(new_new_n622_), .B(new_new_n621_), .C(new_new_n620_), .D(new_new_n413_), .Y(new_new_n623_));
  AOI210     g601(.A0(new_new_n309_), .A1(new_new_n307_), .B0(new_new_n377_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n421_), .B(new_new_n103_), .Y(new_new_n625_));
  OAI210     g603(.A0(new_new_n625_), .A1(new_new_n113_), .B0(new_new_n288_), .Y(new_new_n626_));
  INV        g604(.A(new_new_n394_), .Y(new_new_n627_));
  NA3        g605(.A(new_new_n627_), .B(new_new_n241_), .C(i_7_), .Y(new_new_n628_));
  NA3        g606(.A(new_new_n628_), .B(new_new_n626_), .C(new_new_n624_), .Y(new_new_n629_));
  NO4        g607(.A(new_new_n629_), .B(new_new_n623_), .C(new_new_n618_), .D(new_new_n610_), .Y(new_new_n630_));
  NA4        g608(.A(new_new_n630_), .B(new_new_n598_), .C(new_new_n595_), .D(new_new_n277_), .Y(ori3));
  NA2        g609(.A(i_12_), .B(i_10_), .Y(new_new_n632_));
  NO2        g610(.A(i_11_), .B(new_new_n195_), .Y(new_new_n633_));
  NA3        g611(.A(new_new_n621_), .B(new_new_n413_), .C(new_new_n268_), .Y(new_new_n634_));
  NA2        g612(.A(new_new_n634_), .B(new_new_n40_), .Y(new_new_n635_));
  NOi21      g613(.An(new_new_n97_), .B(new_new_n561_), .Y(new_new_n636_));
  NO3        g614(.A(new_new_n438_), .B(new_new_n314_), .C(new_new_n133_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n290_), .B(new_new_n45_), .Y(new_new_n638_));
  AN2        g616(.A(new_new_n312_), .B(new_new_n55_), .Y(new_new_n639_));
  NO3        g617(.A(new_new_n639_), .B(new_new_n637_), .C(new_new_n636_), .Y(new_new_n640_));
  AOI210     g618(.A0(new_new_n640_), .A1(new_new_n635_), .B0(new_new_n48_), .Y(new_new_n641_));
  NO4        g619(.A(new_new_n273_), .B(new_new_n279_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n642_));
  NA2        g620(.A(new_new_n166_), .B(new_new_n381_), .Y(new_new_n643_));
  NOi21      g621(.An(new_new_n643_), .B(new_new_n642_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n644_), .B(new_new_n63_), .Y(new_new_n645_));
  NOi21      g623(.An(i_5_), .B(i_9_), .Y(new_new_n646_));
  NA2        g624(.A(new_new_n646_), .B(new_new_n306_), .Y(new_new_n647_));
  BUFFER     g625(.A(new_new_n220_), .Y(new_new_n648_));
  AOI210     g626(.A0(new_new_n648_), .A1(new_new_n330_), .B0(new_new_n490_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n649_), .B(new_new_n647_), .Y(new_new_n650_));
  NO3        g628(.A(new_new_n650_), .B(new_new_n645_), .C(new_new_n641_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n166_), .B(new_new_n24_), .Y(new_new_n652_));
  NO2        g630(.A(new_new_n476_), .B(new_new_n402_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n653_), .B(new_new_n652_), .Y(new_new_n654_));
  INV        g632(.A(new_new_n654_), .Y(new_new_n655_));
  NA2        g633(.A(new_new_n382_), .B(i_0_), .Y(new_new_n656_));
  NO3        g634(.A(new_new_n656_), .B(new_new_n280_), .C(new_new_n87_), .Y(new_new_n657_));
  NO4        g635(.A(new_new_n393_), .B(new_new_n184_), .C(new_new_n292_), .D(new_new_n289_), .Y(new_new_n658_));
  AOI210     g636(.A0(new_new_n658_), .A1(i_11_), .B0(new_new_n657_), .Y(new_new_n659_));
  NA2        g637(.A(new_new_n548_), .B(new_new_n242_), .Y(new_new_n660_));
  AOI210     g638(.A0(new_new_n333_), .A1(new_new_n87_), .B0(new_new_n58_), .Y(new_new_n661_));
  NO2        g639(.A(new_new_n661_), .B(new_new_n660_), .Y(new_new_n662_));
  NO2        g640(.A(new_new_n207_), .B(new_new_n153_), .Y(new_new_n663_));
  NA2        g641(.A(i_0_), .B(i_10_), .Y(new_new_n664_));
  INV        g642(.A(new_new_n363_), .Y(new_new_n665_));
  NO4        g643(.A(new_new_n116_), .B(new_new_n58_), .C(new_new_n471_), .D(i_5_), .Y(new_new_n666_));
  AO220      g644(.A0(new_new_n666_), .A1(new_new_n665_), .B0(new_new_n663_), .B1(i_6_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n667_), .B(new_new_n662_), .Y(new_new_n668_));
  NA3        g646(.A(new_new_n668_), .B(new_new_n659_), .C(new_new_n655_), .Y(new_new_n669_));
  NO2        g647(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n670_));
  NA2        g648(.A(i_11_), .B(i_9_), .Y(new_new_n671_));
  NO3        g649(.A(i_12_), .B(new_new_n671_), .C(new_new_n412_), .Y(new_new_n672_));
  AN2        g650(.A(new_new_n672_), .B(new_new_n670_), .Y(new_new_n673_));
  NA2        g651(.A(new_new_n283_), .B(new_new_n165_), .Y(new_new_n674_));
  NA2        g652(.A(new_new_n674_), .B(new_new_n157_), .Y(new_new_n675_));
  NO2        g653(.A(new_new_n671_), .B(new_new_n73_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n163_), .B(i_0_), .Y(new_new_n677_));
  INV        g655(.A(new_new_n287_), .Y(new_new_n678_));
  NO2        g656(.A(new_new_n678_), .B(new_new_n647_), .Y(new_new_n679_));
  NO3        g657(.A(new_new_n679_), .B(new_new_n675_), .C(new_new_n673_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n462_), .B(new_new_n123_), .Y(new_new_n681_));
  NO2        g659(.A(i_6_), .B(new_new_n681_), .Y(new_new_n682_));
  AOI210     g660(.A0(new_new_n308_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n161_), .B(new_new_n104_), .Y(new_new_n684_));
  NOi32      g662(.An(new_new_n683_), .Bn(new_new_n169_), .C(new_new_n684_), .Y(new_new_n685_));
  NA2        g663(.A(new_new_n414_), .B(new_new_n242_), .Y(new_new_n686_));
  NO2        g664(.A(new_new_n686_), .B(new_new_n638_), .Y(new_new_n687_));
  NO3        g665(.A(new_new_n687_), .B(new_new_n685_), .C(new_new_n682_), .Y(new_new_n688_));
  NOi21      g666(.An(i_7_), .B(i_5_), .Y(new_new_n689_));
  INV        g667(.A(new_new_n240_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n688_), .B(new_new_n680_), .Y(new_new_n691_));
  NO2        g669(.A(new_new_n632_), .B(new_new_n239_), .Y(new_new_n692_));
  OA210      g670(.A0(new_new_n329_), .A1(new_new_n190_), .B0(new_new_n328_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n692_), .B(new_new_n676_), .Y(new_new_n694_));
  NA2        g672(.A(new_new_n676_), .B(new_new_n234_), .Y(new_new_n695_));
  OAI210     g673(.A0(i_2_), .A1(new_new_n168_), .B0(new_new_n695_), .Y(new_new_n696_));
  NA2        g674(.A(new_new_n696_), .B(new_new_n329_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n75_), .B(new_new_n550_), .Y(new_new_n698_));
  NA2        g676(.A(new_new_n698_), .B(i_11_), .Y(new_new_n699_));
  NO2        g677(.A(new_new_n699_), .B(new_new_n47_), .Y(new_new_n700_));
  NA2        g678(.A(new_new_n500_), .B(new_new_n365_), .Y(new_new_n701_));
  NAi21      g679(.An(i_9_), .B(i_5_), .Y(new_new_n702_));
  NO2        g680(.A(new_new_n702_), .B(new_new_n286_), .Y(new_new_n703_));
  NA2        g681(.A(new_new_n703_), .B(new_new_n430_), .Y(new_new_n704_));
  OAI220     g682(.A0(new_new_n704_), .A1(new_new_n86_), .B0(new_new_n701_), .B1(new_new_n162_), .Y(new_new_n705_));
  NO3        g683(.A(new_new_n705_), .B(new_new_n700_), .C(new_new_n356_), .Y(new_new_n706_));
  NA3        g684(.A(new_new_n706_), .B(new_new_n697_), .C(new_new_n694_), .Y(new_new_n707_));
  NO3        g685(.A(new_new_n707_), .B(new_new_n691_), .C(new_new_n669_), .Y(new_new_n708_));
  NO2        g686(.A(i_0_), .B(new_new_n527_), .Y(new_new_n709_));
  AOI210     g687(.A0(new_new_n596_), .A1(new_new_n489_), .B0(new_new_n684_), .Y(new_new_n710_));
  INV        g688(.A(new_new_n710_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n201_), .B(new_new_n193_), .Y(new_new_n712_));
  AOI210     g690(.A0(new_new_n712_), .A1(new_new_n656_), .B0(new_new_n153_), .Y(new_new_n713_));
  INV        g691(.A(new_new_n713_), .Y(new_new_n714_));
  NA2        g692(.A(new_new_n714_), .B(new_new_n711_), .Y(new_new_n715_));
  NO3        g693(.A(new_new_n664_), .B(new_new_n646_), .C(new_new_n170_), .Y(new_new_n716_));
  AOI220     g694(.A0(new_new_n716_), .A1(i_11_), .B0(new_new_n380_), .B1(new_new_n75_), .Y(new_new_n717_));
  NO3        g695(.A(new_new_n180_), .B(new_new_n279_), .C(i_0_), .Y(new_new_n718_));
  OAI210     g696(.A0(new_new_n718_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n719_), .B(new_new_n717_), .Y(new_new_n720_));
  NO2        g698(.A(new_new_n200_), .B(new_new_n93_), .Y(new_new_n721_));
  AOI210     g699(.A0(new_new_n721_), .A1(new_new_n709_), .B0(new_new_n110_), .Y(new_new_n722_));
  OR2        g700(.A(new_new_n722_), .B(i_5_), .Y(new_new_n723_));
  AOI210     g701(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n163_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n724_), .B(new_new_n693_), .Y(new_new_n725_));
  NO3        g703(.A(new_new_n638_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n726_));
  NA2        g704(.A(new_new_n341_), .B(new_new_n334_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n727_), .B(new_new_n726_), .Y(new_new_n728_));
  NA3        g706(.A(new_new_n282_), .B(new_new_n161_), .C(new_new_n160_), .Y(new_new_n729_));
  INV        g707(.A(new_new_n729_), .Y(new_new_n730_));
  NO3        g708(.A(new_new_n671_), .B(new_new_n186_), .C(new_new_n170_), .Y(new_new_n731_));
  NO2        g709(.A(new_new_n731_), .B(new_new_n730_), .Y(new_new_n732_));
  NA4        g710(.A(new_new_n732_), .B(new_new_n728_), .C(new_new_n725_), .D(new_new_n723_), .Y(new_new_n733_));
  NO2        g711(.A(new_new_n86_), .B(i_5_), .Y(new_new_n734_));
  NA3        g712(.A(new_new_n633_), .B(new_new_n111_), .C(new_new_n126_), .Y(new_new_n735_));
  INV        g713(.A(new_new_n735_), .Y(new_new_n736_));
  NA2        g714(.A(new_new_n736_), .B(new_new_n734_), .Y(new_new_n737_));
  NAi21      g715(.An(new_new_n199_), .B(new_new_n200_), .Y(new_new_n738_));
  NO4        g716(.A(new_new_n198_), .B(new_new_n180_), .C(i_0_), .D(i_12_), .Y(new_new_n739_));
  AOI220     g717(.A0(new_new_n739_), .A1(new_new_n738_), .B0(new_new_n592_), .B1(new_new_n164_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n689_), .B(new_new_n327_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n741_), .B(new_new_n479_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n742_), .B(new_new_n677_), .Y(new_new_n743_));
  NA3        g721(.A(new_new_n743_), .B(new_new_n740_), .C(new_new_n737_), .Y(new_new_n744_));
  NO4        g722(.A(new_new_n744_), .B(new_new_n733_), .C(new_new_n720_), .D(new_new_n715_), .Y(new_new_n745_));
  OAI210     g723(.A0(new_new_n611_), .A1(new_new_n607_), .B0(new_new_n37_), .Y(new_new_n746_));
  NA2        g724(.A(new_new_n746_), .B(new_new_n420_), .Y(new_new_n747_));
  NA2        g725(.A(new_new_n747_), .B(new_new_n178_), .Y(new_new_n748_));
  NAi31      g726(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n749_));
  AOI210     g727(.A0(new_new_n119_), .A1(new_new_n70_), .B0(new_new_n749_), .Y(new_new_n750_));
  AOI210     g728(.A0(new_new_n750_), .A1(new_new_n48_), .B0(new_new_n658_), .Y(new_new_n751_));
  AOI210     g729(.A0(new_new_n751_), .A1(new_new_n748_), .B0(new_new_n73_), .Y(new_new_n752_));
  INV        g730(.A(new_new_n276_), .Y(new_new_n753_));
  NO2        g731(.A(new_new_n753_), .B(new_new_n556_), .Y(new_new_n754_));
  OAI210     g732(.A0(new_new_n222_), .A1(new_new_n155_), .B0(new_new_n87_), .Y(new_new_n755_));
  NO2        g733(.A(new_new_n755_), .B(i_11_), .Y(new_new_n756_));
  NO3        g734(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n757_));
  OAI210     g735(.A0(new_new_n690_), .A1(new_new_n235_), .B0(new_new_n757_), .Y(new_new_n758_));
  NO2        g736(.A(new_new_n758_), .B(new_new_n527_), .Y(new_new_n759_));
  INV        g737(.A(new_new_n377_), .Y(new_new_n760_));
  INV        g738(.A(new_new_n257_), .Y(new_new_n761_));
  AOI210     g739(.A0(new_new_n761_), .A1(new_new_n760_), .B0(new_new_n41_), .Y(new_new_n762_));
  NO3        g740(.A(new_new_n762_), .B(new_new_n759_), .C(new_new_n756_), .Y(new_new_n763_));
  INV        g741(.A(new_new_n763_), .Y(new_new_n764_));
  NO3        g742(.A(new_new_n764_), .B(new_new_n754_), .C(new_new_n752_), .Y(new_new_n765_));
  NA4        g743(.A(new_new_n765_), .B(new_new_n745_), .C(new_new_n708_), .D(new_new_n651_), .Y(ori4));
  INV        g744(.A(new_new_n499_), .Y(new_new_n769_));
  INV        g745(.A(i_4_), .Y(new_new_n770_));
endmodule


