//Benchmark atmr_intb_466_0.0156

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n351_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n413_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n388_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n452_, mai_mai_n453_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n389_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n464_, men_men_n465_, men_men_n466_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO3        o027(.A(ori_ori_n49_), .B(x11), .C(x09), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x07), .Y(ori_ori_n54_));
  OAI210     o032(.A0(ori_ori_n54_), .A1(ori_ori_n50_), .B0(ori_ori_n47_), .Y(ori_ori_n55_));
  NOi21      o033(.An(x01), .B(x09), .Y(ori_ori_n56_));
  INV        o034(.A(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n51_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(x09), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o038(.A(x07), .Y(ori_ori_n61_));
  AOI220     o039(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n61_), .Y(ori_ori_n62_));
  INV        o040(.A(ori_ori_n59_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n64_), .B(ori_ori_n24_), .Y(ori_ori_n65_));
  OAI220     o043(.A0(ori_ori_n65_), .A1(ori_ori_n63_), .B0(ori_ori_n62_), .B1(ori_ori_n60_), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n61_), .B(ori_ori_n48_), .Y(ori_ori_n67_));
  OAI210     o045(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n67_), .Y(ori_ori_n68_));
  AOI220     o046(.A0(ori_ori_n68_), .A1(ori_ori_n59_), .B0(ori_ori_n66_), .B1(ori_ori_n31_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(ori_ori_n69_), .A1(ori_ori_n55_), .B0(x05), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n61_), .B(ori_ori_n23_), .Y(ori_ori_n71_));
  NA2        o049(.A(x09), .B(x05), .Y(ori_ori_n72_));
  NA2        o050(.A(x10), .B(x06), .Y(ori_ori_n73_));
  NA3        o051(.A(ori_ori_n73_), .B(ori_ori_n72_), .C(ori_ori_n28_), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n61_), .B(ori_ori_n41_), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n74_), .A1(ori_ori_n71_), .B0(x03), .Y(ori_ori_n76_));
  NOi31      o054(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n77_));
  INV        o055(.A(x07), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n78_), .B(ori_ori_n24_), .Y(ori_ori_n79_));
  NO2        o057(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n80_));
  NO2        o058(.A(ori_ori_n80_), .B(ori_ori_n36_), .Y(ori_ori_n81_));
  OAI210     o059(.A0(ori_ori_n80_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n82_));
  AOI210     o060(.A0(ori_ori_n81_), .A1(ori_ori_n48_), .B0(ori_ori_n82_), .Y(ori_ori_n83_));
  NO2        o061(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n84_));
  NO2        o062(.A(x08), .B(x01), .Y(ori_ori_n85_));
  OAI210     o063(.A0(ori_ori_n85_), .A1(ori_ori_n84_), .B0(ori_ori_n35_), .Y(ori_ori_n86_));
  NA2        o064(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n87_));
  NO3        o065(.A(ori_ori_n86_), .B(ori_ori_n83_), .C(ori_ori_n79_), .Y(ori_ori_n88_));
  AN2        o066(.A(ori_ori_n88_), .B(ori_ori_n76_), .Y(ori_ori_n89_));
  INV        o067(.A(ori_ori_n86_), .Y(ori_ori_n90_));
  NO2        o068(.A(x06), .B(x05), .Y(ori_ori_n91_));
  NA2        o069(.A(x11), .B(x00), .Y(ori_ori_n92_));
  NO2        o070(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n93_));
  NOi21      o071(.An(ori_ori_n92_), .B(ori_ori_n93_), .Y(ori_ori_n94_));
  AOI210     o072(.A0(ori_ori_n91_), .A1(ori_ori_n90_), .B0(ori_ori_n94_), .Y(ori_ori_n95_));
  NOi21      o073(.An(x01), .B(x10), .Y(ori_ori_n96_));
  NO2        o074(.A(ori_ori_n29_), .B(ori_ori_n57_), .Y(ori_ori_n97_));
  NO3        o075(.A(ori_ori_n97_), .B(ori_ori_n96_), .C(x06), .Y(ori_ori_n98_));
  NA2        o076(.A(ori_ori_n98_), .B(ori_ori_n27_), .Y(ori_ori_n99_));
  OAI210     o077(.A0(ori_ori_n95_), .A1(x07), .B0(ori_ori_n99_), .Y(ori_ori_n100_));
  NO3        o078(.A(ori_ori_n100_), .B(ori_ori_n89_), .C(ori_ori_n70_), .Y(ori01));
  INV        o079(.A(x12), .Y(ori_ori_n102_));
  INV        o080(.A(x13), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n96_), .B(ori_ori_n28_), .Y(ori_ori_n104_));
  NO2        o082(.A(x10), .B(x01), .Y(ori_ori_n105_));
  NO2        o083(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(ori_ori_n105_), .Y(ori_ori_n107_));
  NA2        o085(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n109_));
  NOi21      o087(.An(ori_ori_n109_), .B(ori_ori_n58_), .Y(ori_ori_n110_));
  NO2        o088(.A(ori_ori_n35_), .B(x02), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n85_), .B(x13), .Y(ori_ori_n112_));
  NA2        o090(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n113_));
  NA2        o091(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n114_));
  NO2        o092(.A(ori_ori_n114_), .B(x05), .Y(ori_ori_n115_));
  NA2        o093(.A(ori_ori_n35_), .B(ori_ori_n57_), .Y(ori_ori_n116_));
  AOI210     o094(.A0(x13), .A1(ori_ori_n81_), .B0(ori_ori_n110_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n117_), .B(ori_ori_n73_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n119_));
  NA2        o097(.A(x10), .B(ori_ori_n57_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(ori_ori_n119_), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n123_));
  NA3        o101(.A(ori_ori_n123_), .B(ori_ori_n122_), .C(x13), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n125_));
  NOi31      o103(.An(ori_ori_n124_), .B(ori_ori_n125_), .C(ori_ori_n121_), .Y(ori_ori_n126_));
  NO3        o104(.A(ori_ori_n126_), .B(x06), .C(x03), .Y(ori_ori_n127_));
  NO2        o105(.A(ori_ori_n127_), .B(ori_ori_n118_), .Y(ori_ori_n128_));
  NA2        o106(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n129_));
  OAI210     o107(.A0(ori_ori_n85_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n130_), .B(ori_ori_n129_), .Y(ori_ori_n131_));
  NO2        o109(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n133_));
  AOI210     o111(.A0(ori_ori_n133_), .A1(ori_ori_n49_), .B0(ori_ori_n132_), .Y(ori_ori_n134_));
  AN2        o112(.A(ori_ori_n134_), .B(ori_ori_n131_), .Y(ori_ori_n135_));
  NO2        o113(.A(x09), .B(x05), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n136_), .B(ori_ori_n47_), .Y(ori_ori_n137_));
  AOI210     o115(.A0(ori_ori_n137_), .A1(ori_ori_n107_), .B0(ori_ori_n49_), .Y(ori_ori_n138_));
  NA2        o116(.A(x09), .B(x00), .Y(ori_ori_n139_));
  NA2        o117(.A(ori_ori_n109_), .B(ori_ori_n139_), .Y(ori_ori_n140_));
  NO2        o118(.A(ori_ori_n140_), .B(ori_ori_n133_), .Y(ori_ori_n141_));
  NO3        o119(.A(ori_ori_n141_), .B(ori_ori_n138_), .C(ori_ori_n135_), .Y(ori_ori_n142_));
  NO2        o120(.A(x03), .B(x02), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n86_), .B(ori_ori_n103_), .Y(ori_ori_n144_));
  OAI210     o122(.A0(ori_ori_n144_), .A1(ori_ori_n110_), .B0(ori_ori_n143_), .Y(ori_ori_n145_));
  OA210      o123(.A0(ori_ori_n142_), .A1(x11), .B0(ori_ori_n145_), .Y(ori_ori_n146_));
  OAI210     o124(.A0(ori_ori_n128_), .A1(ori_ori_n23_), .B0(ori_ori_n146_), .Y(ori_ori_n147_));
  NA2        o125(.A(ori_ori_n107_), .B(ori_ori_n40_), .Y(ori_ori_n148_));
  NAi21      o126(.An(x06), .B(x10), .Y(ori_ori_n149_));
  NOi21      o127(.An(x01), .B(x13), .Y(ori_ori_n150_));
  NA2        o128(.A(ori_ori_n150_), .B(ori_ori_n149_), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n148_), .B(ori_ori_n41_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n153_));
  NA2        o131(.A(ori_ori_n103_), .B(x01), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n154_), .B(x08), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n153_), .B(ori_ori_n48_), .Y(ori_ori_n156_));
  AOI210     o134(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n157_));
  OAI210     o135(.A0(ori_ori_n156_), .A1(ori_ori_n152_), .B0(ori_ori_n157_), .Y(ori_ori_n158_));
  NA2        o136(.A(x04), .B(x02), .Y(ori_ori_n159_));
  NA2        o137(.A(x10), .B(x05), .Y(ori_ori_n160_));
  NO2        o138(.A(x09), .B(x01), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n109_), .B(x08), .Y(ori_ori_n162_));
  INV        o140(.A(ori_ori_n25_), .Y(ori_ori_n163_));
  NAi21      o141(.An(x13), .B(x00), .Y(ori_ori_n164_));
  AOI210     o142(.A0(ori_ori_n29_), .A1(ori_ori_n48_), .B0(ori_ori_n164_), .Y(ori_ori_n165_));
  AN2        o143(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n97_), .B(x06), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n164_), .B(ori_ori_n36_), .Y(ori_ori_n168_));
  INV        o146(.A(ori_ori_n168_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n167_), .B(ori_ori_n166_), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n170_), .B(ori_ori_n163_), .Y(ori_ori_n171_));
  NOi21      o149(.An(x09), .B(x00), .Y(ori_ori_n172_));
  NO3        o150(.A(ori_ori_n84_), .B(ori_ori_n172_), .C(ori_ori_n47_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n173_), .B(ori_ori_n120_), .Y(ori_ori_n174_));
  NA2        o152(.A(x06), .B(x05), .Y(ori_ori_n175_));
  OAI210     o153(.A0(ori_ori_n175_), .A1(ori_ori_n35_), .B0(ori_ori_n102_), .Y(ori_ori_n176_));
  AOI210     o154(.A0(x10), .A1(ori_ori_n58_), .B0(ori_ori_n176_), .Y(ori_ori_n177_));
  NA2        o155(.A(ori_ori_n177_), .B(ori_ori_n174_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n103_), .B(x12), .Y(ori_ori_n179_));
  AOI210     o157(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n179_), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n181_));
  NA2        o159(.A(ori_ori_n181_), .B(x02), .Y(ori_ori_n182_));
  NA2        o160(.A(ori_ori_n180_), .B(ori_ori_n178_), .Y(ori_ori_n183_));
  NA3        o161(.A(ori_ori_n183_), .B(ori_ori_n171_), .C(ori_ori_n158_), .Y(ori_ori_n184_));
  AOI210     o162(.A0(ori_ori_n147_), .A1(ori_ori_n102_), .B0(ori_ori_n184_), .Y(ori_ori_n185_));
  INV        o163(.A(ori_ori_n74_), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n186_), .B(ori_ori_n131_), .Y(ori_ori_n187_));
  NA2        o165(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n188_));
  NA2        o166(.A(ori_ori_n188_), .B(ori_ori_n130_), .Y(ori_ori_n189_));
  AOI210     o167(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n190_));
  NO2        o168(.A(ori_ori_n119_), .B(x06), .Y(ori_ori_n191_));
  AOI210     o169(.A0(ori_ori_n190_), .A1(ori_ori_n189_), .B0(ori_ori_n191_), .Y(ori_ori_n192_));
  AOI210     o170(.A0(ori_ori_n192_), .A1(ori_ori_n187_), .B0(x12), .Y(ori_ori_n193_));
  INV        o171(.A(ori_ori_n77_), .Y(ori_ori_n194_));
  NO2        o172(.A(x05), .B(ori_ori_n51_), .Y(ori_ori_n195_));
  OAI210     o173(.A0(ori_ori_n195_), .A1(ori_ori_n151_), .B0(ori_ori_n57_), .Y(ori_ori_n196_));
  NA2        o174(.A(ori_ori_n196_), .B(ori_ori_n194_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n96_), .B(x06), .Y(ori_ori_n198_));
  AOI210     o176(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n199_));
  NO3        o177(.A(ori_ori_n199_), .B(ori_ori_n198_), .C(ori_ori_n41_), .Y(ori_ori_n200_));
  INV        o178(.A(ori_ori_n133_), .Y(ori_ori_n201_));
  OAI210     o179(.A0(ori_ori_n201_), .A1(ori_ori_n200_), .B0(x02), .Y(ori_ori_n202_));
  AOI210     o180(.A0(ori_ori_n202_), .A1(ori_ori_n197_), .B0(ori_ori_n23_), .Y(ori_ori_n203_));
  OAI210     o181(.A0(ori_ori_n193_), .A1(ori_ori_n57_), .B0(ori_ori_n203_), .Y(ori_ori_n204_));
  INV        o182(.A(ori_ori_n133_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n206_));
  OAI210     o184(.A0(ori_ori_n80_), .A1(ori_ori_n36_), .B0(ori_ori_n113_), .Y(ori_ori_n207_));
  NO2        o185(.A(ori_ori_n103_), .B(x03), .Y(ori_ori_n208_));
  AOI220     o186(.A0(ori_ori_n208_), .A1(ori_ori_n207_), .B0(ori_ori_n77_), .B1(ori_ori_n206_), .Y(ori_ori_n209_));
  NA2        o187(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n210_));
  INV        o188(.A(ori_ori_n149_), .Y(ori_ori_n211_));
  NOi21      o189(.An(x13), .B(x04), .Y(ori_ori_n212_));
  NO3        o190(.A(ori_ori_n212_), .B(ori_ori_n77_), .C(ori_ori_n172_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n213_), .B(x05), .Y(ori_ori_n214_));
  AOI220     o192(.A0(ori_ori_n214_), .A1(ori_ori_n210_), .B0(ori_ori_n211_), .B1(ori_ori_n57_), .Y(ori_ori_n215_));
  OAI210     o193(.A0(ori_ori_n209_), .A1(ori_ori_n205_), .B0(ori_ori_n215_), .Y(ori_ori_n216_));
  INV        o194(.A(ori_ori_n93_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n217_), .B(x12), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n219_));
  NO2        o197(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n220_));
  NA2        o198(.A(ori_ori_n220_), .B(ori_ori_n165_), .Y(ori_ori_n221_));
  AOI210     o199(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n222_));
  NO2        o200(.A(x06), .B(x00), .Y(ori_ori_n223_));
  NO3        o201(.A(ori_ori_n223_), .B(ori_ori_n222_), .C(ori_ori_n41_), .Y(ori_ori_n224_));
  INV        o202(.A(ori_ori_n73_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n225_), .B(ori_ori_n224_), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n227_));
  NA2        o205(.A(ori_ori_n227_), .B(x03), .Y(ori_ori_n228_));
  OA210      o206(.A0(ori_ori_n228_), .A1(ori_ori_n226_), .B0(ori_ori_n221_), .Y(ori_ori_n229_));
  NA2        o207(.A(x13), .B(ori_ori_n102_), .Y(ori_ori_n230_));
  NA3        o208(.A(ori_ori_n230_), .B(ori_ori_n176_), .C(ori_ori_n94_), .Y(ori_ori_n231_));
  OAI210     o209(.A0(ori_ori_n229_), .A1(ori_ori_n219_), .B0(ori_ori_n231_), .Y(ori_ori_n232_));
  AOI210     o210(.A0(ori_ori_n218_), .A1(ori_ori_n216_), .B0(ori_ori_n232_), .Y(ori_ori_n233_));
  AOI210     o211(.A0(ori_ori_n233_), .A1(ori_ori_n204_), .B0(x07), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n72_), .B(ori_ori_n29_), .Y(ori_ori_n235_));
  NOi31      o213(.An(ori_ori_n129_), .B(ori_ori_n212_), .C(ori_ori_n172_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(ori_ori_n235_), .Y(ori_ori_n237_));
  NO2        o215(.A(x08), .B(x05), .Y(ori_ori_n238_));
  NO2        o216(.A(ori_ori_n238_), .B(ori_ori_n222_), .Y(ori_ori_n239_));
  OAI210     o217(.A0(ori_ori_n77_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n240_));
  INV        o218(.A(ori_ori_n240_), .Y(ori_ori_n241_));
  NO2        o219(.A(x12), .B(x02), .Y(ori_ori_n242_));
  INV        o220(.A(ori_ori_n242_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n243_), .B(ori_ori_n217_), .Y(ori_ori_n244_));
  OA210      o222(.A0(ori_ori_n241_), .A1(ori_ori_n237_), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n246_));
  NO2        o224(.A(ori_ori_n246_), .B(x01), .Y(ori_ori_n247_));
  INV        o225(.A(ori_ori_n247_), .Y(ori_ori_n248_));
  AOI210     o226(.A0(ori_ori_n248_), .A1(ori_ori_n124_), .B0(ori_ori_n29_), .Y(ori_ori_n249_));
  NA2        o227(.A(ori_ori_n103_), .B(x04), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n250_), .B(ori_ori_n28_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n251_), .B(ori_ori_n112_), .Y(ori_ori_n252_));
  NO3        o230(.A(ori_ori_n92_), .B(x12), .C(x03), .Y(ori_ori_n253_));
  OAI210     o231(.A0(ori_ori_n252_), .A1(ori_ori_n249_), .B0(ori_ori_n253_), .Y(ori_ori_n254_));
  NOi21      o232(.An(ori_ori_n235_), .B(ori_ori_n198_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n256_));
  NA2        o234(.A(ori_ori_n255_), .B(ori_ori_n256_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n258_));
  NO3        o236(.A(ori_ori_n258_), .B(ori_ori_n199_), .C(ori_ori_n167_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n219_), .B(ori_ori_n28_), .Y(ori_ori_n260_));
  OAI210     o238(.A0(ori_ori_n259_), .A1(ori_ori_n205_), .B0(ori_ori_n260_), .Y(ori_ori_n261_));
  NA3        o239(.A(ori_ori_n261_), .B(ori_ori_n257_), .C(ori_ori_n254_), .Y(ori_ori_n262_));
  NO3        o240(.A(ori_ori_n262_), .B(ori_ori_n245_), .C(ori_ori_n234_), .Y(ori_ori_n263_));
  OAI210     o241(.A0(ori_ori_n185_), .A1(ori_ori_n61_), .B0(ori_ori_n263_), .Y(ori02));
  AOI210     o242(.A0(ori_ori_n129_), .A1(ori_ori_n86_), .B0(ori_ori_n122_), .Y(ori_ori_n265_));
  NOi21      o243(.An(ori_ori_n213_), .B(ori_ori_n161_), .Y(ori_ori_n266_));
  NO2        o244(.A(ori_ori_n103_), .B(ori_ori_n35_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n266_), .B(ori_ori_n32_), .Y(ori_ori_n268_));
  OAI210     o246(.A0(ori_ori_n268_), .A1(ori_ori_n265_), .B0(ori_ori_n160_), .Y(ori_ori_n269_));
  INV        o247(.A(ori_ori_n160_), .Y(ori_ori_n270_));
  AOI210     o248(.A0(ori_ori_n111_), .A1(ori_ori_n87_), .B0(ori_ori_n199_), .Y(ori_ori_n271_));
  OAI220     o249(.A0(ori_ori_n271_), .A1(ori_ori_n103_), .B0(ori_ori_n86_), .B1(ori_ori_n51_), .Y(ori_ori_n272_));
  AOI220     o250(.A0(ori_ori_n272_), .A1(ori_ori_n270_), .B0(ori_ori_n144_), .B1(ori_ori_n143_), .Y(ori_ori_n273_));
  AOI210     o251(.A0(ori_ori_n273_), .A1(ori_ori_n269_), .B0(ori_ori_n48_), .Y(ori_ori_n274_));
  NO2        o252(.A(x05), .B(x02), .Y(ori_ori_n275_));
  OAI210     o253(.A0(ori_ori_n189_), .A1(ori_ori_n172_), .B0(ori_ori_n275_), .Y(ori_ori_n276_));
  AOI220     o254(.A0(ori_ori_n238_), .A1(ori_ori_n58_), .B0(ori_ori_n56_), .B1(ori_ori_n36_), .Y(ori_ori_n277_));
  NOi21      o255(.An(ori_ori_n267_), .B(ori_ori_n277_), .Y(ori_ori_n278_));
  INV        o256(.A(ori_ori_n278_), .Y(ori_ori_n279_));
  AOI210     o257(.A0(ori_ori_n279_), .A1(ori_ori_n276_), .B0(ori_ori_n133_), .Y(ori_ori_n280_));
  NAi21      o258(.An(ori_ori_n214_), .B(ori_ori_n209_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n227_), .B(ori_ori_n47_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n282_), .B(ori_ori_n281_), .Y(ori_ori_n283_));
  AN2        o261(.A(ori_ori_n208_), .B(ori_ori_n207_), .Y(ori_ori_n284_));
  OAI210     o262(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n285_));
  NA2        o263(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n286_));
  OA210      o264(.A0(ori_ori_n286_), .A1(x08), .B0(ori_ori_n137_), .Y(ori_ori_n287_));
  AOI210     o265(.A0(ori_ori_n287_), .A1(ori_ori_n130_), .B0(ori_ori_n285_), .Y(ori_ori_n288_));
  OAI210     o266(.A0(ori_ori_n288_), .A1(ori_ori_n284_), .B0(ori_ori_n97_), .Y(ori_ori_n289_));
  INV        o267(.A(ori_ori_n143_), .Y(ori_ori_n290_));
  OAI220     o268(.A0(ori_ori_n239_), .A1(ori_ori_n104_), .B0(ori_ori_n290_), .B1(ori_ori_n121_), .Y(ori_ori_n291_));
  NA2        o269(.A(ori_ori_n291_), .B(x13), .Y(ori_ori_n292_));
  NA3        o270(.A(ori_ori_n292_), .B(ori_ori_n289_), .C(ori_ori_n283_), .Y(ori_ori_n293_));
  NO3        o271(.A(ori_ori_n293_), .B(ori_ori_n280_), .C(ori_ori_n274_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n132_), .B(x03), .Y(ori_ori_n295_));
  INV        o273(.A(ori_ori_n164_), .Y(ori_ori_n296_));
  OAI210     o274(.A0(ori_ori_n51_), .A1(ori_ori_n35_), .B0(ori_ori_n36_), .Y(ori_ori_n297_));
  AOI220     o275(.A0(ori_ori_n297_), .A1(ori_ori_n296_), .B0(ori_ori_n181_), .B1(x08), .Y(ori_ori_n298_));
  OAI210     o276(.A0(ori_ori_n298_), .A1(ori_ori_n258_), .B0(ori_ori_n295_), .Y(ori_ori_n299_));
  NA2        o277(.A(ori_ori_n299_), .B(ori_ori_n105_), .Y(ori_ori_n300_));
  NA2        o278(.A(ori_ori_n159_), .B(ori_ori_n154_), .Y(ori_ori_n301_));
  AN2        o279(.A(ori_ori_n301_), .B(ori_ori_n162_), .Y(ori_ori_n302_));
  INV        o280(.A(ori_ori_n56_), .Y(ori_ori_n303_));
  OAI220     o281(.A0(ori_ori_n250_), .A1(ori_ori_n303_), .B0(ori_ori_n122_), .B1(ori_ori_n28_), .Y(ori_ori_n304_));
  OAI210     o282(.A0(ori_ori_n304_), .A1(ori_ori_n302_), .B0(ori_ori_n106_), .Y(ori_ori_n305_));
  NA2        o283(.A(ori_ori_n250_), .B(ori_ori_n102_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n102_), .B(ori_ori_n41_), .Y(ori_ori_n307_));
  NA3        o285(.A(ori_ori_n307_), .B(ori_ori_n306_), .C(ori_ori_n121_), .Y(ori_ori_n308_));
  NA4        o286(.A(ori_ori_n308_), .B(ori_ori_n305_), .C(ori_ori_n300_), .D(ori_ori_n48_), .Y(ori_ori_n309_));
  INV        o287(.A(ori_ori_n181_), .Y(ori_ori_n310_));
  NA2        o288(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n311_));
  OAI220     o289(.A0(ori_ori_n311_), .A1(ori_ori_n413_), .B0(ori_ori_n310_), .B1(ori_ori_n59_), .Y(ori_ori_n312_));
  NA2        o290(.A(ori_ori_n312_), .B(x02), .Y(ori_ori_n313_));
  INV        o291(.A(ori_ori_n220_), .Y(ori_ori_n314_));
  NA2        o292(.A(ori_ori_n179_), .B(x04), .Y(ori_ori_n315_));
  NO3        o293(.A(ori_ori_n179_), .B(ori_ori_n153_), .C(ori_ori_n52_), .Y(ori_ori_n316_));
  OAI210     o294(.A0(ori_ori_n139_), .A1(ori_ori_n36_), .B0(ori_ori_n102_), .Y(ori_ori_n317_));
  OAI210     o295(.A0(ori_ori_n317_), .A1(ori_ori_n173_), .B0(ori_ori_n316_), .Y(ori_ori_n318_));
  NA3        o296(.A(ori_ori_n318_), .B(ori_ori_n313_), .C(x06), .Y(ori_ori_n319_));
  NA2        o297(.A(x09), .B(x03), .Y(ori_ori_n320_));
  OAI220     o298(.A0(ori_ori_n320_), .A1(ori_ori_n120_), .B0(ori_ori_n188_), .B1(ori_ori_n64_), .Y(ori_ori_n321_));
  NO3        o299(.A(ori_ori_n258_), .B(ori_ori_n119_), .C(x08), .Y(ori_ori_n322_));
  INV        o300(.A(ori_ori_n322_), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n324_));
  NO3        o302(.A(ori_ori_n109_), .B(ori_ori_n120_), .C(ori_ori_n38_), .Y(ori_ori_n325_));
  AOI210     o303(.A0(ori_ori_n316_), .A1(ori_ori_n324_), .B0(ori_ori_n325_), .Y(ori_ori_n326_));
  OAI210     o304(.A0(ori_ori_n323_), .A1(ori_ori_n28_), .B0(ori_ori_n326_), .Y(ori_ori_n327_));
  AO220      o305(.A0(ori_ori_n327_), .A1(x04), .B0(ori_ori_n321_), .B1(x05), .Y(ori_ori_n328_));
  AOI210     o306(.A0(ori_ori_n319_), .A1(ori_ori_n309_), .B0(ori_ori_n328_), .Y(ori_ori_n329_));
  OAI210     o307(.A0(ori_ori_n294_), .A1(x12), .B0(ori_ori_n329_), .Y(ori03));
  OR2        o308(.A(ori_ori_n42_), .B(ori_ori_n206_), .Y(ori_ori_n331_));
  AOI210     o309(.A0(ori_ori_n144_), .A1(ori_ori_n102_), .B0(ori_ori_n331_), .Y(ori_ori_n332_));
  AO210      o310(.A0(ori_ori_n314_), .A1(ori_ori_n87_), .B0(ori_ori_n315_), .Y(ori_ori_n333_));
  NA2        o311(.A(ori_ori_n179_), .B(ori_ori_n143_), .Y(ori_ori_n334_));
  NA3        o312(.A(ori_ori_n334_), .B(ori_ori_n333_), .C(ori_ori_n182_), .Y(ori_ori_n335_));
  OAI210     o313(.A0(ori_ori_n335_), .A1(ori_ori_n332_), .B0(x05), .Y(ori_ori_n336_));
  NA2        o314(.A(ori_ori_n331_), .B(x05), .Y(ori_ori_n337_));
  AOI210     o315(.A0(ori_ori_n130_), .A1(ori_ori_n194_), .B0(ori_ori_n337_), .Y(ori_ori_n338_));
  AOI210     o316(.A0(ori_ori_n208_), .A1(ori_ori_n81_), .B0(ori_ori_n115_), .Y(ori_ori_n339_));
  OAI220     o317(.A0(ori_ori_n339_), .A1(ori_ori_n59_), .B0(ori_ori_n286_), .B1(ori_ori_n277_), .Y(ori_ori_n340_));
  OAI210     o318(.A0(ori_ori_n340_), .A1(ori_ori_n338_), .B0(ori_ori_n102_), .Y(ori_ori_n341_));
  AOI210     o319(.A0(ori_ori_n137_), .A1(ori_ori_n60_), .B0(ori_ori_n38_), .Y(ori_ori_n342_));
  NO2        o320(.A(ori_ori_n161_), .B(ori_ori_n125_), .Y(ori_ori_n343_));
  OAI220     o321(.A0(ori_ori_n343_), .A1(ori_ori_n37_), .B0(ori_ori_n140_), .B1(x13), .Y(ori_ori_n344_));
  OAI210     o322(.A0(ori_ori_n344_), .A1(ori_ori_n342_), .B0(x04), .Y(ori_ori_n345_));
  NO3        o323(.A(ori_ori_n307_), .B(ori_ori_n86_), .C(ori_ori_n59_), .Y(ori_ori_n346_));
  AOI210     o324(.A0(ori_ori_n169_), .A1(ori_ori_n102_), .B0(ori_ori_n137_), .Y(ori_ori_n347_));
  OA210      o325(.A0(ori_ori_n155_), .A1(x12), .B0(ori_ori_n125_), .Y(ori_ori_n348_));
  NO3        o326(.A(ori_ori_n348_), .B(ori_ori_n347_), .C(ori_ori_n346_), .Y(ori_ori_n349_));
  NA4        o327(.A(ori_ori_n349_), .B(ori_ori_n345_), .C(ori_ori_n341_), .D(ori_ori_n336_), .Y(ori04));
  NO2        o328(.A(ori_ori_n90_), .B(ori_ori_n39_), .Y(ori_ori_n351_));
  XO2        o329(.A(ori_ori_n351_), .B(ori_ori_n230_), .Y(ori05));
  AOI210     o330(.A0(ori_ori_n72_), .A1(ori_ori_n52_), .B0(ori_ori_n191_), .Y(ori_ori_n353_));
  AOI210     o331(.A0(ori_ori_n353_), .A1(ori_ori_n285_), .B0(ori_ori_n25_), .Y(ori_ori_n354_));
  NA3        o332(.A(ori_ori_n133_), .B(ori_ori_n122_), .C(ori_ori_n31_), .Y(ori_ori_n355_));
  AOI210     o333(.A0(ori_ori_n211_), .A1(ori_ori_n57_), .B0(ori_ori_n91_), .Y(ori_ori_n356_));
  AOI210     o334(.A0(ori_ori_n356_), .A1(ori_ori_n355_), .B0(ori_ori_n24_), .Y(ori_ori_n357_));
  OAI210     o335(.A0(ori_ori_n357_), .A1(ori_ori_n354_), .B0(ori_ori_n102_), .Y(ori_ori_n358_));
  NA2        o336(.A(x11), .B(ori_ori_n31_), .Y(ori_ori_n359_));
  NA2        o337(.A(ori_ori_n23_), .B(ori_ori_n28_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n235_), .B(x03), .Y(ori_ori_n361_));
  OAI220     o339(.A0(ori_ori_n361_), .A1(ori_ori_n360_), .B0(ori_ori_n359_), .B1(ori_ori_n82_), .Y(ori_ori_n362_));
  OAI210     o340(.A0(ori_ori_n26_), .A1(ori_ori_n102_), .B0(x07), .Y(ori_ori_n363_));
  AOI210     o341(.A0(ori_ori_n362_), .A1(x06), .B0(ori_ori_n363_), .Y(ori_ori_n364_));
  AOI210     o342(.A0(ori_ori_n82_), .A1(ori_ori_n31_), .B0(ori_ori_n52_), .Y(ori_ori_n365_));
  NO3        o343(.A(ori_ori_n365_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n366_));
  OR2        o344(.A(x02), .B(ori_ori_n219_), .Y(ori_ori_n367_));
  NA2        o345(.A(ori_ori_n223_), .B(ori_ori_n217_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n368_), .B(ori_ori_n367_), .Y(ori_ori_n369_));
  OAI210     o347(.A0(ori_ori_n369_), .A1(ori_ori_n366_), .B0(ori_ori_n102_), .Y(ori_ori_n370_));
  NA2        o348(.A(ori_ori_n33_), .B(ori_ori_n102_), .Y(ori_ori_n371_));
  AOI210     o349(.A0(ori_ori_n371_), .A1(ori_ori_n93_), .B0(x07), .Y(ori_ori_n372_));
  AOI220     o350(.A0(ori_ori_n372_), .A1(ori_ori_n370_), .B0(ori_ori_n364_), .B1(ori_ori_n358_), .Y(ori_ori_n373_));
  OR2        o351(.A(ori_ori_n246_), .B(ori_ori_n243_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n136_), .B(ori_ori_n28_), .Y(ori_ori_n375_));
  AOI210     o353(.A0(ori_ori_n374_), .A1(ori_ori_n47_), .B0(ori_ori_n375_), .Y(ori_ori_n376_));
  NA2        o354(.A(ori_ori_n376_), .B(ori_ori_n103_), .Y(ori_ori_n377_));
  AOI210     o355(.A0(ori_ori_n315_), .A1(ori_ori_n108_), .B0(ori_ori_n242_), .Y(ori_ori_n378_));
  NOi21      o356(.An(ori_ori_n295_), .B(ori_ori_n125_), .Y(ori_ori_n379_));
  NO2        o357(.A(ori_ori_n379_), .B(ori_ori_n243_), .Y(ori_ori_n380_));
  OAI210     o358(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n381_));
  AOI210     o359(.A0(ori_ori_n230_), .A1(ori_ori_n47_), .B0(ori_ori_n381_), .Y(ori_ori_n382_));
  NO4        o360(.A(ori_ori_n382_), .B(ori_ori_n380_), .C(ori_ori_n378_), .D(x08), .Y(ori_ori_n383_));
  NA2        o361(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n384_));
  NO2        o362(.A(ori_ori_n384_), .B(x03), .Y(ori_ori_n385_));
  NO2        o363(.A(x13), .B(x12), .Y(ori_ori_n386_));
  NO2        o364(.A(ori_ori_n122_), .B(ori_ori_n28_), .Y(ori_ori_n387_));
  NO2        o365(.A(ori_ori_n387_), .B(ori_ori_n247_), .Y(ori_ori_n388_));
  OR3        o366(.A(ori_ori_n388_), .B(x12), .C(x03), .Y(ori_ori_n389_));
  NA3        o367(.A(ori_ori_n310_), .B(ori_ori_n116_), .C(x12), .Y(ori_ori_n390_));
  AO210      o368(.A0(ori_ori_n310_), .A1(ori_ori_n116_), .B0(ori_ori_n230_), .Y(ori_ori_n391_));
  NA4        o369(.A(ori_ori_n391_), .B(ori_ori_n390_), .C(ori_ori_n389_), .D(x08), .Y(ori_ori_n392_));
  AOI210     o370(.A0(ori_ori_n386_), .A1(ori_ori_n385_), .B0(ori_ori_n392_), .Y(ori_ori_n393_));
  AOI210     o371(.A0(ori_ori_n383_), .A1(ori_ori_n377_), .B0(ori_ori_n393_), .Y(ori_ori_n394_));
  INV        o372(.A(x03), .Y(ori_ori_n395_));
  NO2        o373(.A(ori_ori_n136_), .B(ori_ori_n43_), .Y(ori_ori_n396_));
  OAI210     o374(.A0(ori_ori_n396_), .A1(ori_ori_n395_), .B0(ori_ori_n168_), .Y(ori_ori_n397_));
  NA3        o375(.A(ori_ori_n388_), .B(ori_ori_n379_), .C(ori_ori_n306_), .Y(ori_ori_n398_));
  INV        o376(.A(x14), .Y(ori_ori_n399_));
  NO3        o377(.A(ori_ori_n154_), .B(ori_ori_n75_), .C(ori_ori_n57_), .Y(ori_ori_n400_));
  NO2        o378(.A(ori_ori_n400_), .B(ori_ori_n399_), .Y(ori_ori_n401_));
  NA3        o379(.A(ori_ori_n401_), .B(ori_ori_n398_), .C(ori_ori_n397_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n371_), .B(ori_ori_n61_), .Y(ori_ori_n403_));
  NOi21      o381(.An(ori_ori_n250_), .B(ori_ori_n140_), .Y(ori_ori_n404_));
  NO3        o382(.A(ori_ori_n119_), .B(ori_ori_n24_), .C(x06), .Y(ori_ori_n405_));
  INV        o383(.A(ori_ori_n405_), .Y(ori_ori_n406_));
  OAI210     o384(.A0(ori_ori_n44_), .A1(x04), .B0(ori_ori_n406_), .Y(ori_ori_n407_));
  OAI210     o385(.A0(ori_ori_n407_), .A1(ori_ori_n404_), .B0(ori_ori_n102_), .Y(ori_ori_n408_));
  OAI210     o386(.A0(ori_ori_n403_), .A1(ori_ori_n92_), .B0(ori_ori_n408_), .Y(ori_ori_n409_));
  NO4        o387(.A(ori_ori_n409_), .B(ori_ori_n402_), .C(ori_ori_n394_), .D(ori_ori_n373_), .Y(ori06));
  INV        o388(.A(ori_ori_n40_), .Y(ori_ori_n413_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  NOi21      m029(.An(x01), .B(x09), .Y(mai_mai_n52_));
  INV        m030(.A(x00), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  NO2        m032(.A(mai_mai_n54_), .B(mai_mai_n52_), .Y(mai_mai_n55_));
  NA2        m033(.A(x09), .B(mai_mai_n53_), .Y(mai_mai_n56_));
  INV        m034(.A(x07), .Y(mai_mai_n57_));
  INV        m035(.A(mai_mai_n55_), .Y(mai_mai_n58_));
  NA2        m036(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n59_), .B(mai_mai_n24_), .Y(mai_mai_n60_));
  NO2        m038(.A(mai_mai_n60_), .B(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m039(.A(mai_mai_n57_), .B(mai_mai_n48_), .Y(mai_mai_n62_));
  OAI210     m040(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n62_), .Y(mai_mai_n63_));
  AOI220     m041(.A0(mai_mai_n63_), .A1(mai_mai_n55_), .B0(mai_mai_n61_), .B1(mai_mai_n31_), .Y(mai_mai_n64_));
  NO2        m042(.A(mai_mai_n64_), .B(x05), .Y(mai_mai_n65_));
  NO2        m043(.A(mai_mai_n57_), .B(mai_mai_n23_), .Y(mai_mai_n66_));
  NA2        m044(.A(x09), .B(x05), .Y(mai_mai_n67_));
  NA2        m045(.A(x10), .B(x06), .Y(mai_mai_n68_));
  NA3        m046(.A(mai_mai_n68_), .B(mai_mai_n67_), .C(mai_mai_n28_), .Y(mai_mai_n69_));
  OAI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n66_), .B0(x03), .Y(mai_mai_n70_));
  NOi31      m048(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n71_));
  NO2        m049(.A(mai_mai_n452_), .B(mai_mai_n24_), .Y(mai_mai_n72_));
  NO2        m050(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n36_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n73_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n75_));
  AOI210     m053(.A0(mai_mai_n74_), .A1(mai_mai_n48_), .B0(mai_mai_n75_), .Y(mai_mai_n76_));
  NO2        m054(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n77_));
  NO2        m055(.A(x08), .B(x01), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n78_), .A1(mai_mai_n77_), .B0(mai_mai_n35_), .Y(mai_mai_n79_));
  NA2        m057(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n80_));
  NO3        m058(.A(mai_mai_n79_), .B(mai_mai_n76_), .C(mai_mai_n72_), .Y(mai_mai_n81_));
  AN2        m059(.A(mai_mai_n81_), .B(mai_mai_n70_), .Y(mai_mai_n82_));
  INV        m060(.A(mai_mai_n79_), .Y(mai_mai_n83_));
  NO2        m061(.A(x06), .B(x05), .Y(mai_mai_n84_));
  NA2        m062(.A(x11), .B(x00), .Y(mai_mai_n85_));
  NO2        m063(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n86_));
  NOi21      m064(.An(mai_mai_n85_), .B(mai_mai_n86_), .Y(mai_mai_n87_));
  AOI210     m065(.A0(mai_mai_n84_), .A1(mai_mai_n83_), .B0(mai_mai_n87_), .Y(mai_mai_n88_));
  NOi21      m066(.An(x01), .B(x10), .Y(mai_mai_n89_));
  NO2        m067(.A(mai_mai_n29_), .B(mai_mai_n53_), .Y(mai_mai_n90_));
  NO3        m068(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(x06), .Y(mai_mai_n91_));
  NA2        m069(.A(mai_mai_n91_), .B(mai_mai_n27_), .Y(mai_mai_n92_));
  OAI210     m070(.A0(mai_mai_n88_), .A1(x07), .B0(mai_mai_n92_), .Y(mai_mai_n93_));
  NO3        m071(.A(mai_mai_n93_), .B(mai_mai_n82_), .C(mai_mai_n65_), .Y(mai01));
  INV        m072(.A(x12), .Y(mai_mai_n95_));
  INV        m073(.A(x13), .Y(mai_mai_n96_));
  NA2        m074(.A(x08), .B(x04), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n97_), .B(mai_mai_n53_), .Y(mai_mai_n98_));
  NA2        m076(.A(mai_mai_n98_), .B(mai_mai_n84_), .Y(mai_mai_n99_));
  NA2        m077(.A(mai_mai_n89_), .B(mai_mai_n28_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n67_), .Y(mai_mai_n101_));
  NO2        m079(.A(x10), .B(x01), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NA2        m082(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n105_));
  NO3        m083(.A(mai_mai_n105_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n106_));
  AOI210     m084(.A0(mai_mai_n106_), .A1(mai_mai_n104_), .B0(mai_mai_n101_), .Y(mai_mai_n107_));
  AOI210     m085(.A0(mai_mai_n107_), .A1(mai_mai_n99_), .B0(mai_mai_n96_), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n52_), .B(x05), .Y(mai_mai_n109_));
  NOi21      m087(.An(mai_mai_n109_), .B(mai_mai_n54_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n111_));
  NA3        m089(.A(x13), .B(mai_mai_n111_), .C(x06), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n112_), .B(mai_mai_n110_), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n78_), .B(x13), .Y(mai_mai_n114_));
  NA2        m092(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NA2        m094(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n117_), .B(x05), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n118_), .B(mai_mai_n116_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n35_), .B(mai_mai_n53_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n120_), .B(mai_mai_n96_), .Y(mai_mai_n121_));
  AOI210     m099(.A0(mai_mai_n121_), .A1(mai_mai_n74_), .B0(mai_mai_n110_), .Y(mai_mai_n122_));
  AOI210     m100(.A0(mai_mai_n122_), .A1(mai_mai_n119_), .B0(mai_mai_n68_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n124_));
  NA2        m102(.A(x10), .B(mai_mai_n53_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n125_), .B(mai_mai_n124_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n127_));
  NO3        m105(.A(mai_mai_n120_), .B(mai_mai_n73_), .C(mai_mai_n36_), .Y(mai_mai_n128_));
  NO2        m106(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n129_));
  NO3        m107(.A(mai_mai_n129_), .B(mai_mai_n128_), .C(mai_mai_n126_), .Y(mai_mai_n130_));
  NO3        m108(.A(mai_mai_n130_), .B(x06), .C(x03), .Y(mai_mai_n131_));
  NO4        m109(.A(mai_mai_n131_), .B(mai_mai_n123_), .C(mai_mai_n113_), .D(mai_mai_n108_), .Y(mai_mai_n132_));
  NA2        m110(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n133_));
  OAI210     m111(.A0(mai_mai_n78_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n134_), .B(mai_mai_n133_), .Y(mai_mai_n135_));
  NO2        m113(.A(mai_mai_n35_), .B(mai_mai_n47_), .Y(mai_mai_n136_));
  AN2        m114(.A(mai_mai_n84_), .B(mai_mai_n136_), .Y(mai_mai_n137_));
  NO2        m115(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n138_));
  NA2        m116(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n139_));
  AOI210     m117(.A0(mai_mai_n139_), .A1(mai_mai_n49_), .B0(mai_mai_n138_), .Y(mai_mai_n140_));
  OA210      m118(.A0(mai_mai_n140_), .A1(mai_mai_n137_), .B0(mai_mai_n135_), .Y(mai_mai_n141_));
  NO2        m119(.A(x09), .B(x05), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n142_), .B(mai_mai_n47_), .Y(mai_mai_n143_));
  NO2        m121(.A(mai_mai_n104_), .B(mai_mai_n49_), .Y(mai_mai_n144_));
  NA2        m122(.A(x09), .B(x00), .Y(mai_mai_n145_));
  NA2        m123(.A(mai_mai_n109_), .B(mai_mai_n145_), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n71_), .B(mai_mai_n50_), .Y(mai_mai_n147_));
  AOI210     m125(.A0(mai_mai_n147_), .A1(mai_mai_n146_), .B0(mai_mai_n139_), .Y(mai_mai_n148_));
  NO3        m126(.A(mai_mai_n148_), .B(mai_mai_n144_), .C(mai_mai_n141_), .Y(mai_mai_n149_));
  NO2        m127(.A(x03), .B(x02), .Y(mai_mai_n150_));
  NA2        m128(.A(mai_mai_n79_), .B(mai_mai_n96_), .Y(mai_mai_n151_));
  OAI210     m129(.A0(mai_mai_n151_), .A1(mai_mai_n110_), .B0(mai_mai_n150_), .Y(mai_mai_n152_));
  OA210      m130(.A0(mai_mai_n149_), .A1(x11), .B0(mai_mai_n152_), .Y(mai_mai_n153_));
  OAI210     m131(.A0(mai_mai_n132_), .A1(mai_mai_n23_), .B0(mai_mai_n153_), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n104_), .B(mai_mai_n40_), .Y(mai_mai_n155_));
  NAi21      m133(.An(x06), .B(x10), .Y(mai_mai_n156_));
  NOi21      m134(.An(x01), .B(x13), .Y(mai_mai_n157_));
  NA2        m135(.A(mai_mai_n157_), .B(mai_mai_n156_), .Y(mai_mai_n158_));
  BUFFER     m136(.A(mai_mai_n158_), .Y(mai_mai_n159_));
  AOI210     m137(.A0(mai_mai_n159_), .A1(mai_mai_n155_), .B0(mai_mai_n41_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n161_));
  NA2        m139(.A(mai_mai_n96_), .B(x01), .Y(mai_mai_n162_));
  NO2        m140(.A(mai_mai_n162_), .B(x08), .Y(mai_mai_n163_));
  OAI210     m141(.A0(x05), .A1(mai_mai_n163_), .B0(mai_mai_n50_), .Y(mai_mai_n164_));
  AOI210     m142(.A0(mai_mai_n164_), .A1(mai_mai_n161_), .B0(mai_mai_n48_), .Y(mai_mai_n165_));
  AOI210     m143(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n166_));
  OAI210     m144(.A0(mai_mai_n165_), .A1(mai_mai_n160_), .B0(mai_mai_n166_), .Y(mai_mai_n167_));
  NA2        m145(.A(x04), .B(x02), .Y(mai_mai_n168_));
  NA2        m146(.A(x10), .B(x05), .Y(mai_mai_n169_));
  NA2        m147(.A(x09), .B(x06), .Y(mai_mai_n170_));
  AOI210     m148(.A0(mai_mai_n170_), .A1(mai_mai_n169_), .B0(x11), .Y(mai_mai_n171_));
  NO2        m149(.A(x09), .B(x01), .Y(mai_mai_n172_));
  NO3        m150(.A(mai_mai_n172_), .B(mai_mai_n102_), .C(mai_mai_n31_), .Y(mai_mai_n173_));
  OAI210     m151(.A0(mai_mai_n173_), .A1(mai_mai_n171_), .B0(x00), .Y(mai_mai_n174_));
  NO2        m152(.A(mai_mai_n109_), .B(x08), .Y(mai_mai_n175_));
  NA3        m153(.A(mai_mai_n157_), .B(mai_mai_n156_), .C(mai_mai_n50_), .Y(mai_mai_n176_));
  NA2        m154(.A(mai_mai_n89_), .B(x05), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n177_), .B(mai_mai_n176_), .Y(mai_mai_n178_));
  AOI210     m156(.A0(mai_mai_n175_), .A1(x06), .B0(mai_mai_n178_), .Y(mai_mai_n179_));
  OAI210     m157(.A0(mai_mai_n179_), .A1(x11), .B0(mai_mai_n174_), .Y(mai_mai_n180_));
  NAi21      m158(.An(mai_mai_n168_), .B(mai_mai_n180_), .Y(mai_mai_n181_));
  INV        m159(.A(mai_mai_n25_), .Y(mai_mai_n182_));
  NAi21      m160(.An(x13), .B(x00), .Y(mai_mai_n183_));
  AOI210     m161(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n183_), .Y(mai_mai_n184_));
  AOI220     m162(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n185_));
  OAI210     m163(.A0(mai_mai_n169_), .A1(mai_mai_n35_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  AN2        m164(.A(mai_mai_n186_), .B(mai_mai_n184_), .Y(mai_mai_n187_));
  BUFFER     m165(.A(mai_mai_n67_), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n90_), .B(x06), .Y(mai_mai_n189_));
  NO2        m167(.A(mai_mai_n183_), .B(mai_mai_n36_), .Y(mai_mai_n190_));
  INV        m168(.A(mai_mai_n190_), .Y(mai_mai_n191_));
  OAI220     m169(.A0(mai_mai_n191_), .A1(mai_mai_n170_), .B0(mai_mai_n189_), .B1(mai_mai_n188_), .Y(mai_mai_n192_));
  OAI210     m170(.A0(mai_mai_n192_), .A1(mai_mai_n187_), .B0(mai_mai_n182_), .Y(mai_mai_n193_));
  NOi21      m171(.An(x09), .B(x00), .Y(mai_mai_n194_));
  NO3        m172(.A(mai_mai_n77_), .B(mai_mai_n194_), .C(mai_mai_n47_), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n195_), .B(mai_mai_n125_), .Y(mai_mai_n196_));
  NA2        m174(.A(x10), .B(x08), .Y(mai_mai_n197_));
  INV        m175(.A(mai_mai_n197_), .Y(mai_mai_n198_));
  NA2        m176(.A(x06), .B(x05), .Y(mai_mai_n199_));
  OAI210     m177(.A0(mai_mai_n199_), .A1(mai_mai_n35_), .B0(mai_mai_n95_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n95_), .B(mai_mai_n196_), .Y(mai_mai_n201_));
  NO2        m179(.A(mai_mai_n96_), .B(x12), .Y(mai_mai_n202_));
  AOI210     m180(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n202_), .Y(mai_mai_n203_));
  NA2        m181(.A(mai_mai_n89_), .B(mai_mai_n50_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n205_));
  NA2        m183(.A(mai_mai_n205_), .B(x02), .Y(mai_mai_n206_));
  NO2        m184(.A(mai_mai_n206_), .B(mai_mai_n204_), .Y(mai_mai_n207_));
  AOI210     m185(.A0(mai_mai_n203_), .A1(mai_mai_n201_), .B0(mai_mai_n207_), .Y(mai_mai_n208_));
  NA4        m186(.A(mai_mai_n208_), .B(mai_mai_n193_), .C(mai_mai_n181_), .D(mai_mai_n167_), .Y(mai_mai_n209_));
  AOI210     m187(.A0(mai_mai_n154_), .A1(mai_mai_n95_), .B0(mai_mai_n209_), .Y(mai_mai_n210_));
  INV        m188(.A(mai_mai_n69_), .Y(mai_mai_n211_));
  NA2        m189(.A(mai_mai_n211_), .B(mai_mai_n135_), .Y(mai_mai_n212_));
  NA2        m190(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n213_));
  NA2        m191(.A(mai_mai_n213_), .B(mai_mai_n134_), .Y(mai_mai_n214_));
  AOI210     m192(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n124_), .B(x06), .Y(mai_mai_n216_));
  AOI210     m194(.A0(mai_mai_n215_), .A1(mai_mai_n214_), .B0(mai_mai_n216_), .Y(mai_mai_n217_));
  AOI210     m195(.A0(mai_mai_n217_), .A1(mai_mai_n212_), .B0(x12), .Y(mai_mai_n218_));
  INV        m196(.A(mai_mai_n71_), .Y(mai_mai_n219_));
  OAI210     m197(.A0(x09), .A1(mai_mai_n158_), .B0(mai_mai_n53_), .Y(mai_mai_n220_));
  NA2        m198(.A(mai_mai_n220_), .B(mai_mai_n219_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n89_), .B(x06), .Y(mai_mai_n222_));
  AOI210     m200(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n50_), .Y(mai_mai_n223_));
  NO3        m201(.A(mai_mai_n223_), .B(mai_mai_n222_), .C(mai_mai_n41_), .Y(mai_mai_n224_));
  NA4        m202(.A(mai_mai_n156_), .B(mai_mai_n52_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n225_), .B(mai_mai_n139_), .Y(mai_mai_n226_));
  OAI210     m204(.A0(mai_mai_n226_), .A1(mai_mai_n224_), .B0(x02), .Y(mai_mai_n227_));
  AOI210     m205(.A0(mai_mai_n227_), .A1(mai_mai_n221_), .B0(mai_mai_n23_), .Y(mai_mai_n228_));
  OAI210     m206(.A0(mai_mai_n218_), .A1(mai_mai_n53_), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  INV        m207(.A(mai_mai_n139_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n50_), .B(x03), .Y(mai_mai_n231_));
  OAI210     m209(.A0(mai_mai_n73_), .A1(mai_mai_n36_), .B0(mai_mai_n115_), .Y(mai_mai_n232_));
  NO2        m210(.A(mai_mai_n96_), .B(x03), .Y(mai_mai_n233_));
  AOI220     m211(.A0(mai_mai_n233_), .A1(mai_mai_n232_), .B0(mai_mai_n71_), .B1(mai_mai_n231_), .Y(mai_mai_n234_));
  NA2        m212(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n235_));
  INV        m213(.A(mai_mai_n156_), .Y(mai_mai_n236_));
  NOi21      m214(.An(x13), .B(x04), .Y(mai_mai_n237_));
  NO3        m215(.A(mai_mai_n237_), .B(mai_mai_n71_), .C(mai_mai_n194_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n238_), .B(x05), .Y(mai_mai_n239_));
  AOI220     m217(.A0(mai_mai_n239_), .A1(mai_mai_n235_), .B0(mai_mai_n236_), .B1(mai_mai_n53_), .Y(mai_mai_n240_));
  OAI210     m218(.A0(mai_mai_n234_), .A1(mai_mai_n230_), .B0(mai_mai_n240_), .Y(mai_mai_n241_));
  INV        m219(.A(mai_mai_n86_), .Y(mai_mai_n242_));
  NO2        m220(.A(mai_mai_n242_), .B(x12), .Y(mai_mai_n243_));
  NA2        m221(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n244_));
  NO2        m222(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n245_));
  OAI210     m223(.A0(mai_mai_n245_), .A1(mai_mai_n186_), .B0(mai_mai_n184_), .Y(mai_mai_n246_));
  AOI210     m224(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n247_));
  NO2        m225(.A(x06), .B(x00), .Y(mai_mai_n248_));
  NO3        m226(.A(mai_mai_n248_), .B(mai_mai_n247_), .C(mai_mai_n41_), .Y(mai_mai_n249_));
  OAI210     m227(.A0(mai_mai_n97_), .A1(mai_mai_n145_), .B0(mai_mai_n68_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n250_), .B(mai_mai_n249_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n252_), .B(x03), .Y(mai_mai_n253_));
  OA210      m231(.A0(mai_mai_n253_), .A1(mai_mai_n251_), .B0(mai_mai_n246_), .Y(mai_mai_n254_));
  NA2        m232(.A(x13), .B(mai_mai_n95_), .Y(mai_mai_n255_));
  NA3        m233(.A(mai_mai_n255_), .B(mai_mai_n200_), .C(mai_mai_n87_), .Y(mai_mai_n256_));
  OAI210     m234(.A0(mai_mai_n254_), .A1(mai_mai_n244_), .B0(mai_mai_n256_), .Y(mai_mai_n257_));
  AOI210     m235(.A0(mai_mai_n243_), .A1(mai_mai_n241_), .B0(mai_mai_n257_), .Y(mai_mai_n258_));
  AOI210     m236(.A0(mai_mai_n258_), .A1(mai_mai_n229_), .B0(x07), .Y(mai_mai_n259_));
  NA2        m237(.A(mai_mai_n67_), .B(mai_mai_n29_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n237_), .B(mai_mai_n194_), .Y(mai_mai_n261_));
  AOI210     m239(.A0(mai_mai_n261_), .A1(mai_mai_n147_), .B0(mai_mai_n260_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n96_), .B(x06), .Y(mai_mai_n263_));
  INV        m241(.A(mai_mai_n263_), .Y(mai_mai_n264_));
  NO2        m242(.A(x08), .B(x05), .Y(mai_mai_n265_));
  NO2        m243(.A(mai_mai_n265_), .B(mai_mai_n247_), .Y(mai_mai_n266_));
  NA2        m244(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n267_));
  OAI210     m245(.A0(mai_mai_n266_), .A1(mai_mai_n264_), .B0(mai_mai_n267_), .Y(mai_mai_n268_));
  NO2        m246(.A(x12), .B(x02), .Y(mai_mai_n269_));
  INV        m247(.A(mai_mai_n269_), .Y(mai_mai_n270_));
  NO2        m248(.A(mai_mai_n270_), .B(mai_mai_n242_), .Y(mai_mai_n271_));
  OA210      m249(.A0(mai_mai_n268_), .A1(mai_mai_n262_), .B0(mai_mai_n271_), .Y(mai_mai_n272_));
  NA2        m250(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n273_), .B(x01), .Y(mai_mai_n274_));
  NOi21      m252(.An(mai_mai_n78_), .B(mai_mai_n115_), .Y(mai_mai_n275_));
  NO2        m253(.A(mai_mai_n275_), .B(mai_mai_n274_), .Y(mai_mai_n276_));
  NO2        m254(.A(mai_mai_n276_), .B(mai_mai_n29_), .Y(mai_mai_n277_));
  NA2        m255(.A(mai_mai_n263_), .B(mai_mai_n232_), .Y(mai_mai_n278_));
  NA2        m256(.A(mai_mai_n96_), .B(x04), .Y(mai_mai_n279_));
  NA2        m257(.A(mai_mai_n279_), .B(mai_mai_n28_), .Y(mai_mai_n280_));
  OAI210     m258(.A0(mai_mai_n280_), .A1(mai_mai_n114_), .B0(mai_mai_n278_), .Y(mai_mai_n281_));
  NO3        m259(.A(mai_mai_n85_), .B(x12), .C(x03), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n281_), .A1(mai_mai_n277_), .B0(mai_mai_n282_), .Y(mai_mai_n283_));
  AOI210     m261(.A0(mai_mai_n204_), .A1(mai_mai_n199_), .B0(mai_mai_n97_), .Y(mai_mai_n284_));
  NOi21      m262(.An(mai_mai_n260_), .B(mai_mai_n222_), .Y(mai_mai_n285_));
  NO2        m263(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n286_));
  OAI210     m264(.A0(mai_mai_n285_), .A1(mai_mai_n284_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  NO2        m265(.A(mai_mai_n54_), .B(x05), .Y(mai_mai_n288_));
  NO3        m266(.A(mai_mai_n288_), .B(mai_mai_n223_), .C(mai_mai_n189_), .Y(mai_mai_n289_));
  NO2        m267(.A(mai_mai_n244_), .B(mai_mai_n28_), .Y(mai_mai_n290_));
  OAI210     m268(.A0(mai_mai_n289_), .A1(mai_mai_n230_), .B0(mai_mai_n290_), .Y(mai_mai_n291_));
  NA3        m269(.A(mai_mai_n291_), .B(mai_mai_n287_), .C(mai_mai_n283_), .Y(mai_mai_n292_));
  NO3        m270(.A(mai_mai_n292_), .B(mai_mai_n272_), .C(mai_mai_n259_), .Y(mai_mai_n293_));
  OAI210     m271(.A0(mai_mai_n210_), .A1(mai_mai_n57_), .B0(mai_mai_n293_), .Y(mai02));
  AOI210     m272(.A0(mai_mai_n133_), .A1(mai_mai_n79_), .B0(mai_mai_n127_), .Y(mai_mai_n295_));
  NOi21      m273(.An(mai_mai_n238_), .B(mai_mai_n172_), .Y(mai_mai_n296_));
  NO2        m274(.A(mai_mai_n96_), .B(mai_mai_n35_), .Y(mai_mai_n297_));
  NA3        m275(.A(mai_mai_n297_), .B(mai_mai_n198_), .C(mai_mai_n52_), .Y(mai_mai_n298_));
  OAI210     m276(.A0(mai_mai_n296_), .A1(mai_mai_n32_), .B0(mai_mai_n298_), .Y(mai_mai_n299_));
  OAI210     m277(.A0(mai_mai_n299_), .A1(mai_mai_n295_), .B0(mai_mai_n169_), .Y(mai_mai_n300_));
  INV        m278(.A(mai_mai_n169_), .Y(mai_mai_n301_));
  AOI210     m279(.A0(mai_mai_n111_), .A1(mai_mai_n80_), .B0(mai_mai_n223_), .Y(mai_mai_n302_));
  OAI220     m280(.A0(mai_mai_n302_), .A1(mai_mai_n96_), .B0(mai_mai_n79_), .B1(mai_mai_n50_), .Y(mai_mai_n303_));
  AOI220     m281(.A0(mai_mai_n303_), .A1(mai_mai_n301_), .B0(mai_mai_n151_), .B1(mai_mai_n150_), .Y(mai_mai_n304_));
  AOI210     m282(.A0(mai_mai_n304_), .A1(mai_mai_n300_), .B0(mai_mai_n48_), .Y(mai_mai_n305_));
  NO2        m283(.A(x05), .B(x02), .Y(mai_mai_n306_));
  OAI210     m284(.A0(mai_mai_n214_), .A1(mai_mai_n194_), .B0(mai_mai_n306_), .Y(mai_mai_n307_));
  AOI220     m285(.A0(mai_mai_n265_), .A1(mai_mai_n54_), .B0(mai_mai_n52_), .B1(mai_mai_n36_), .Y(mai_mai_n308_));
  NOi21      m286(.An(mai_mai_n297_), .B(mai_mai_n308_), .Y(mai_mai_n309_));
  AOI210     m287(.A0(mai_mai_n237_), .A1(mai_mai_n73_), .B0(mai_mai_n309_), .Y(mai_mai_n310_));
  AOI210     m288(.A0(mai_mai_n310_), .A1(mai_mai_n307_), .B0(mai_mai_n139_), .Y(mai_mai_n311_));
  NAi21      m289(.An(mai_mai_n239_), .B(mai_mai_n234_), .Y(mai_mai_n312_));
  NO2        m290(.A(mai_mai_n252_), .B(mai_mai_n47_), .Y(mai_mai_n313_));
  NA2        m291(.A(mai_mai_n313_), .B(mai_mai_n312_), .Y(mai_mai_n314_));
  AN2        m292(.A(mai_mai_n233_), .B(mai_mai_n232_), .Y(mai_mai_n315_));
  OAI210     m293(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n316_));
  NA2        m294(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n317_));
  OA210      m295(.A0(mai_mai_n317_), .A1(x08), .B0(mai_mai_n143_), .Y(mai_mai_n318_));
  AOI210     m296(.A0(mai_mai_n318_), .A1(mai_mai_n134_), .B0(mai_mai_n316_), .Y(mai_mai_n319_));
  OAI210     m297(.A0(mai_mai_n319_), .A1(mai_mai_n315_), .B0(mai_mai_n90_), .Y(mai_mai_n320_));
  NA3        m298(.A(mai_mai_n90_), .B(mai_mai_n78_), .C(mai_mai_n231_), .Y(mai_mai_n321_));
  NA3        m299(.A(mai_mai_n89_), .B(mai_mai_n77_), .C(mai_mai_n42_), .Y(mai_mai_n322_));
  AOI210     m300(.A0(mai_mai_n322_), .A1(mai_mai_n321_), .B0(x04), .Y(mai_mai_n323_));
  INV        m301(.A(mai_mai_n150_), .Y(mai_mai_n324_));
  OAI220     m302(.A0(mai_mai_n266_), .A1(mai_mai_n100_), .B0(mai_mai_n324_), .B1(mai_mai_n126_), .Y(mai_mai_n325_));
  AOI210     m303(.A0(mai_mai_n325_), .A1(x13), .B0(mai_mai_n323_), .Y(mai_mai_n326_));
  NA3        m304(.A(mai_mai_n326_), .B(mai_mai_n320_), .C(mai_mai_n314_), .Y(mai_mai_n327_));
  NO3        m305(.A(mai_mai_n327_), .B(mai_mai_n311_), .C(mai_mai_n305_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n138_), .B(x03), .Y(mai_mai_n329_));
  INV        m307(.A(mai_mai_n183_), .Y(mai_mai_n330_));
  AOI220     m308(.A0(x08), .A1(mai_mai_n330_), .B0(mai_mai_n205_), .B1(x08), .Y(mai_mai_n331_));
  OAI210     m309(.A0(mai_mai_n331_), .A1(mai_mai_n288_), .B0(mai_mai_n329_), .Y(mai_mai_n332_));
  NA2        m310(.A(mai_mai_n332_), .B(mai_mai_n102_), .Y(mai_mai_n333_));
  NA2        m311(.A(mai_mai_n168_), .B(mai_mai_n162_), .Y(mai_mai_n334_));
  AN2        m312(.A(mai_mai_n334_), .B(mai_mai_n175_), .Y(mai_mai_n335_));
  NO2        m313(.A(mai_mai_n127_), .B(mai_mai_n28_), .Y(mai_mai_n336_));
  OAI210     m314(.A0(mai_mai_n336_), .A1(mai_mai_n335_), .B0(mai_mai_n103_), .Y(mai_mai_n337_));
  NA2        m315(.A(mai_mai_n279_), .B(mai_mai_n95_), .Y(mai_mai_n338_));
  NA2        m316(.A(mai_mai_n95_), .B(mai_mai_n41_), .Y(mai_mai_n339_));
  NA3        m317(.A(mai_mai_n339_), .B(mai_mai_n338_), .C(mai_mai_n126_), .Y(mai_mai_n340_));
  NA4        m318(.A(mai_mai_n340_), .B(mai_mai_n337_), .C(mai_mai_n333_), .D(mai_mai_n48_), .Y(mai_mai_n341_));
  INV        m319(.A(mai_mai_n205_), .Y(mai_mai_n342_));
  NO2        m320(.A(mai_mai_n163_), .B(mai_mai_n40_), .Y(mai_mai_n343_));
  NA2        m321(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n344_));
  OAI220     m322(.A0(mai_mai_n344_), .A1(mai_mai_n343_), .B0(mai_mai_n342_), .B1(mai_mai_n55_), .Y(mai_mai_n345_));
  NA2        m323(.A(mai_mai_n345_), .B(x02), .Y(mai_mai_n346_));
  INV        m324(.A(mai_mai_n245_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n202_), .B(x04), .Y(mai_mai_n348_));
  NO2        m326(.A(mai_mai_n348_), .B(mai_mai_n347_), .Y(mai_mai_n349_));
  NO3        m327(.A(mai_mai_n185_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n350_));
  OAI210     m328(.A0(mai_mai_n350_), .A1(mai_mai_n349_), .B0(mai_mai_n90_), .Y(mai_mai_n351_));
  NO3        m329(.A(mai_mai_n202_), .B(mai_mai_n161_), .C(mai_mai_n51_), .Y(mai_mai_n352_));
  OAI210     m330(.A0(mai_mai_n145_), .A1(mai_mai_n36_), .B0(mai_mai_n95_), .Y(mai_mai_n353_));
  OAI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n195_), .B0(mai_mai_n352_), .Y(mai_mai_n354_));
  NA4        m332(.A(mai_mai_n354_), .B(mai_mai_n351_), .C(mai_mai_n346_), .D(x06), .Y(mai_mai_n355_));
  NA2        m333(.A(x09), .B(x03), .Y(mai_mai_n356_));
  OAI220     m334(.A0(mai_mai_n356_), .A1(mai_mai_n125_), .B0(mai_mai_n213_), .B1(mai_mai_n59_), .Y(mai_mai_n357_));
  OAI220     m335(.A0(mai_mai_n162_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n358_));
  NO3        m336(.A(mai_mai_n288_), .B(mai_mai_n124_), .C(x08), .Y(mai_mai_n359_));
  AOI210     m337(.A0(mai_mai_n358_), .A1(mai_mai_n230_), .B0(mai_mai_n359_), .Y(mai_mai_n360_));
  NO2        m338(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n361_));
  NO3        m339(.A(mai_mai_n109_), .B(mai_mai_n125_), .C(mai_mai_n38_), .Y(mai_mai_n362_));
  AOI210     m340(.A0(mai_mai_n352_), .A1(mai_mai_n361_), .B0(mai_mai_n362_), .Y(mai_mai_n363_));
  OAI210     m341(.A0(mai_mai_n360_), .A1(mai_mai_n28_), .B0(mai_mai_n363_), .Y(mai_mai_n364_));
  AO220      m342(.A0(mai_mai_n364_), .A1(x04), .B0(mai_mai_n357_), .B1(x05), .Y(mai_mai_n365_));
  AOI210     m343(.A0(mai_mai_n355_), .A1(mai_mai_n341_), .B0(mai_mai_n365_), .Y(mai_mai_n366_));
  OAI210     m344(.A0(mai_mai_n328_), .A1(x12), .B0(mai_mai_n366_), .Y(mai03));
  OR2        m345(.A(mai_mai_n42_), .B(mai_mai_n231_), .Y(mai_mai_n368_));
  AOI210     m346(.A0(mai_mai_n151_), .A1(mai_mai_n95_), .B0(mai_mai_n368_), .Y(mai_mai_n369_));
  AO210      m347(.A0(mai_mai_n347_), .A1(mai_mai_n80_), .B0(mai_mai_n348_), .Y(mai_mai_n370_));
  NA2        m348(.A(mai_mai_n202_), .B(mai_mai_n150_), .Y(mai_mai_n371_));
  NA3        m349(.A(mai_mai_n371_), .B(mai_mai_n370_), .C(mai_mai_n206_), .Y(mai_mai_n372_));
  OAI210     m350(.A0(mai_mai_n372_), .A1(mai_mai_n369_), .B0(x05), .Y(mai_mai_n373_));
  NA2        m351(.A(mai_mai_n368_), .B(x05), .Y(mai_mai_n374_));
  AOI210     m352(.A0(mai_mai_n134_), .A1(mai_mai_n219_), .B0(mai_mai_n374_), .Y(mai_mai_n375_));
  AOI210     m353(.A0(mai_mai_n233_), .A1(mai_mai_n74_), .B0(mai_mai_n118_), .Y(mai_mai_n376_));
  OAI220     m354(.A0(mai_mai_n376_), .A1(mai_mai_n55_), .B0(mai_mai_n317_), .B1(mai_mai_n308_), .Y(mai_mai_n377_));
  OAI210     m355(.A0(mai_mai_n377_), .A1(mai_mai_n375_), .B0(mai_mai_n95_), .Y(mai_mai_n378_));
  AOI210     m356(.A0(mai_mai_n143_), .A1(mai_mai_n56_), .B0(mai_mai_n38_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n172_), .B(mai_mai_n129_), .Y(mai_mai_n380_));
  OAI220     m358(.A0(mai_mai_n380_), .A1(mai_mai_n37_), .B0(mai_mai_n146_), .B1(x13), .Y(mai_mai_n381_));
  OAI210     m359(.A0(mai_mai_n381_), .A1(mai_mai_n379_), .B0(x04), .Y(mai_mai_n382_));
  NO3        m360(.A(mai_mai_n339_), .B(mai_mai_n79_), .C(mai_mai_n55_), .Y(mai_mai_n383_));
  AOI210     m361(.A0(mai_mai_n191_), .A1(mai_mai_n95_), .B0(mai_mai_n143_), .Y(mai_mai_n384_));
  OA210      m362(.A0(mai_mai_n163_), .A1(x12), .B0(mai_mai_n129_), .Y(mai_mai_n385_));
  NO3        m363(.A(mai_mai_n385_), .B(mai_mai_n384_), .C(mai_mai_n383_), .Y(mai_mai_n386_));
  NA4        m364(.A(mai_mai_n386_), .B(mai_mai_n382_), .C(mai_mai_n378_), .D(mai_mai_n373_), .Y(mai04));
  NO2        m365(.A(mai_mai_n83_), .B(mai_mai_n39_), .Y(mai_mai_n388_));
  XO2        m366(.A(mai_mai_n388_), .B(mai_mai_n255_), .Y(mai05));
  INV        m367(.A(mai_mai_n51_), .Y(mai_mai_n390_));
  AOI210     m368(.A0(mai_mai_n390_), .A1(mai_mai_n316_), .B0(mai_mai_n25_), .Y(mai_mai_n391_));
  NO2        m369(.A(x06), .B(mai_mai_n24_), .Y(mai_mai_n392_));
  OAI210     m370(.A0(mai_mai_n392_), .A1(mai_mai_n391_), .B0(mai_mai_n95_), .Y(mai_mai_n393_));
  NA2        m371(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n394_));
  NA2        m372(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n395_));
  NA2        m373(.A(mai_mai_n260_), .B(x03), .Y(mai_mai_n396_));
  OAI220     m374(.A0(mai_mai_n396_), .A1(mai_mai_n395_), .B0(mai_mai_n394_), .B1(mai_mai_n75_), .Y(mai_mai_n397_));
  OAI210     m375(.A0(mai_mai_n26_), .A1(mai_mai_n95_), .B0(x07), .Y(mai_mai_n398_));
  AOI210     m376(.A0(mai_mai_n397_), .A1(x06), .B0(mai_mai_n398_), .Y(mai_mai_n399_));
  NA2        m377(.A(mai_mai_n75_), .B(mai_mai_n31_), .Y(mai_mai_n400_));
  NO3        m378(.A(mai_mai_n400_), .B(mai_mai_n23_), .C(x00), .Y(mai_mai_n401_));
  NO2        m379(.A(mai_mai_n396_), .B(mai_mai_n263_), .Y(mai_mai_n402_));
  OR2        m380(.A(mai_mai_n402_), .B(mai_mai_n244_), .Y(mai_mai_n403_));
  NA2        m381(.A(mai_mai_n157_), .B(x05), .Y(mai_mai_n404_));
  NA3        m382(.A(mai_mai_n404_), .B(mai_mai_n248_), .C(mai_mai_n242_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n406_));
  OAI210     m384(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n407_));
  OR3        m385(.A(mai_mai_n407_), .B(mai_mai_n406_), .C(mai_mai_n44_), .Y(mai_mai_n408_));
  NA3        m386(.A(mai_mai_n408_), .B(mai_mai_n405_), .C(mai_mai_n403_), .Y(mai_mai_n409_));
  OAI210     m387(.A0(mai_mai_n409_), .A1(mai_mai_n401_), .B0(mai_mai_n95_), .Y(mai_mai_n410_));
  NA2        m388(.A(mai_mai_n33_), .B(mai_mai_n95_), .Y(mai_mai_n411_));
  AOI210     m389(.A0(mai_mai_n411_), .A1(mai_mai_n86_), .B0(x07), .Y(mai_mai_n412_));
  AOI220     m390(.A0(mai_mai_n412_), .A1(mai_mai_n410_), .B0(mai_mai_n399_), .B1(mai_mai_n393_), .Y(mai_mai_n413_));
  AOI210     m391(.A0(mai_mai_n406_), .A1(x07), .B0(mai_mai_n138_), .Y(mai_mai_n414_));
  OR2        m392(.A(mai_mai_n414_), .B(x03), .Y(mai_mai_n415_));
  NO2        m393(.A(x07), .B(x11), .Y(mai_mai_n416_));
  NO3        m394(.A(mai_mai_n416_), .B(mai_mai_n142_), .C(mai_mai_n28_), .Y(mai_mai_n417_));
  AOI210     m395(.A0(mai_mai_n417_), .A1(mai_mai_n415_), .B0(mai_mai_n47_), .Y(mai_mai_n418_));
  NA2        m396(.A(mai_mai_n418_), .B(mai_mai_n96_), .Y(mai_mai_n419_));
  AOI210     m397(.A0(mai_mai_n348_), .A1(mai_mai_n105_), .B0(mai_mai_n269_), .Y(mai_mai_n420_));
  NOi21      m398(.An(mai_mai_n329_), .B(mai_mai_n129_), .Y(mai_mai_n421_));
  NO2        m399(.A(mai_mai_n421_), .B(mai_mai_n270_), .Y(mai_mai_n422_));
  OAI210     m400(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n423_));
  AOI210     m401(.A0(mai_mai_n255_), .A1(mai_mai_n47_), .B0(mai_mai_n423_), .Y(mai_mai_n424_));
  NO4        m402(.A(mai_mai_n424_), .B(mai_mai_n422_), .C(mai_mai_n420_), .D(x08), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n127_), .B(mai_mai_n28_), .Y(mai_mai_n426_));
  NO2        m404(.A(mai_mai_n426_), .B(mai_mai_n274_), .Y(mai_mai_n427_));
  OR3        m405(.A(mai_mai_n427_), .B(x12), .C(x03), .Y(mai_mai_n428_));
  NA3        m406(.A(mai_mai_n342_), .B(mai_mai_n120_), .C(x12), .Y(mai_mai_n429_));
  AO210      m407(.A0(mai_mai_n342_), .A1(mai_mai_n120_), .B0(mai_mai_n255_), .Y(mai_mai_n430_));
  NA4        m408(.A(mai_mai_n430_), .B(mai_mai_n429_), .C(mai_mai_n428_), .D(x08), .Y(mai_mai_n431_));
  INV        m409(.A(mai_mai_n431_), .Y(mai_mai_n432_));
  AOI210     m410(.A0(mai_mai_n425_), .A1(mai_mai_n419_), .B0(mai_mai_n432_), .Y(mai_mai_n433_));
  OAI210     m411(.A0(x07), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n434_));
  OAI220     m412(.A0(mai_mai_n453_), .A1(mai_mai_n395_), .B0(mai_mai_n142_), .B1(mai_mai_n43_), .Y(mai_mai_n435_));
  OAI210     m413(.A0(mai_mai_n435_), .A1(mai_mai_n434_), .B0(mai_mai_n190_), .Y(mai_mai_n436_));
  NA3        m414(.A(mai_mai_n427_), .B(mai_mai_n421_), .C(mai_mai_n338_), .Y(mai_mai_n437_));
  INV        m415(.A(x14), .Y(mai_mai_n438_));
  NO3        m416(.A(mai_mai_n329_), .B(mai_mai_n100_), .C(x11), .Y(mai_mai_n439_));
  NO3        m417(.A(x06), .B(mai_mai_n339_), .C(mai_mai_n183_), .Y(mai_mai_n440_));
  NO3        m418(.A(mai_mai_n440_), .B(mai_mai_n439_), .C(mai_mai_n438_), .Y(mai_mai_n441_));
  NA3        m419(.A(mai_mai_n441_), .B(mai_mai_n437_), .C(mai_mai_n436_), .Y(mai_mai_n442_));
  AOI220     m420(.A0(mai_mai_n411_), .A1(mai_mai_n57_), .B0(mai_mai_n426_), .B1(mai_mai_n161_), .Y(mai_mai_n443_));
  NOi21      m421(.An(mai_mai_n279_), .B(mai_mai_n146_), .Y(mai_mai_n444_));
  NA2        m422(.A(mai_mai_n286_), .B(mai_mai_n236_), .Y(mai_mai_n445_));
  OAI210     m423(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n445_), .Y(mai_mai_n446_));
  OAI210     m424(.A0(mai_mai_n446_), .A1(mai_mai_n444_), .B0(mai_mai_n95_), .Y(mai_mai_n447_));
  OAI210     m425(.A0(mai_mai_n443_), .A1(mai_mai_n85_), .B0(mai_mai_n447_), .Y(mai_mai_n448_));
  NO4        m426(.A(mai_mai_n448_), .B(mai_mai_n442_), .C(mai_mai_n433_), .D(mai_mai_n413_), .Y(mai06));
  INV        m427(.A(x07), .Y(mai_mai_n452_));
  INV        m428(.A(x07), .Y(mai_mai_n453_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  AOI220     u039(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n61_), .Y(men_men_n62_));
  INV        u040(.A(men_men_n59_), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n29_), .B(x02), .Y(men_men_n64_));
  NA2        u042(.A(men_men_n64_), .B(men_men_n24_), .Y(men_men_n65_));
  OAI220     u043(.A0(men_men_n65_), .A1(men_men_n63_), .B0(men_men_n62_), .B1(men_men_n60_), .Y(men_men_n66_));
  NA2        u044(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n67_));
  OAI210     u045(.A0(men_men_n30_), .A1(x11), .B0(men_men_n67_), .Y(men_men_n68_));
  AOI220     u046(.A0(men_men_n68_), .A1(men_men_n59_), .B0(men_men_n66_), .B1(men_men_n31_), .Y(men_men_n69_));
  AOI210     u047(.A0(men_men_n69_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n70_));
  NA2        u048(.A(x10), .B(x09), .Y(men_men_n71_));
  NO2        u049(.A(men_men_n61_), .B(men_men_n23_), .Y(men_men_n72_));
  NA2        u050(.A(x09), .B(x05), .Y(men_men_n73_));
  NA2        u051(.A(x10), .B(x06), .Y(men_men_n74_));
  NA2        u052(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n76_));
  OAI210     u054(.A0(men_men_n75_), .A1(men_men_n72_), .B0(x03), .Y(men_men_n77_));
  NOi31      u055(.An(x08), .B(x04), .C(x00), .Y(men_men_n78_));
  NO2        u056(.A(x10), .B(x09), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n464_), .B(men_men_n24_), .Y(men_men_n80_));
  NO2        u058(.A(x09), .B(men_men_n41_), .Y(men_men_n81_));
  NO2        u059(.A(men_men_n81_), .B(men_men_n36_), .Y(men_men_n82_));
  OAI210     u060(.A0(men_men_n81_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n83_));
  AOI210     u061(.A0(men_men_n82_), .A1(men_men_n48_), .B0(men_men_n83_), .Y(men_men_n84_));
  NO2        u062(.A(men_men_n36_), .B(x00), .Y(men_men_n85_));
  NO2        u063(.A(x08), .B(x01), .Y(men_men_n86_));
  OAI210     u064(.A0(men_men_n86_), .A1(men_men_n85_), .B0(men_men_n35_), .Y(men_men_n87_));
  NA2        u065(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n88_));
  NO3        u066(.A(men_men_n87_), .B(men_men_n84_), .C(men_men_n80_), .Y(men_men_n89_));
  AN2        u067(.A(men_men_n89_), .B(men_men_n77_), .Y(men_men_n90_));
  INV        u068(.A(men_men_n87_), .Y(men_men_n91_));
  NO2        u069(.A(x06), .B(x05), .Y(men_men_n92_));
  NA2        u070(.A(x11), .B(x00), .Y(men_men_n93_));
  NO2        u071(.A(x11), .B(men_men_n47_), .Y(men_men_n94_));
  NOi21      u072(.An(men_men_n93_), .B(men_men_n94_), .Y(men_men_n95_));
  NOi21      u073(.An(x01), .B(x10), .Y(men_men_n96_));
  NO2        u074(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n97_));
  NO3        u075(.A(men_men_n97_), .B(men_men_n96_), .C(x06), .Y(men_men_n98_));
  NA2        u076(.A(men_men_n98_), .B(men_men_n27_), .Y(men_men_n99_));
  OAI210     u077(.A0(men_men_n465_), .A1(x07), .B0(men_men_n99_), .Y(men_men_n100_));
  NO3        u078(.A(men_men_n100_), .B(men_men_n90_), .C(men_men_n70_), .Y(men01));
  INV        u079(.A(x12), .Y(men_men_n102_));
  INV        u080(.A(x13), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n466_), .B(men_men_n71_), .Y(men_men_n104_));
  NA2        u082(.A(x08), .B(x04), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n105_), .B(men_men_n57_), .Y(men_men_n106_));
  NA2        u084(.A(men_men_n106_), .B(men_men_n104_), .Y(men_men_n107_));
  NA2        u085(.A(men_men_n96_), .B(men_men_n28_), .Y(men_men_n108_));
  NO2        u086(.A(men_men_n108_), .B(men_men_n73_), .Y(men_men_n109_));
  NO2        u087(.A(x10), .B(x01), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n29_), .B(x00), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n111_), .B(men_men_n110_), .Y(men_men_n112_));
  NA2        u090(.A(x04), .B(men_men_n28_), .Y(men_men_n113_));
  NO3        u091(.A(men_men_n113_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n114_));
  AOI210     u092(.A0(men_men_n114_), .A1(men_men_n112_), .B0(men_men_n109_), .Y(men_men_n115_));
  AOI210     u093(.A0(men_men_n115_), .A1(men_men_n107_), .B0(men_men_n103_), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n56_), .B(x05), .Y(men_men_n117_));
  NOi21      u095(.An(men_men_n117_), .B(men_men_n58_), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n35_), .B(x02), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n103_), .B(men_men_n36_), .Y(men_men_n120_));
  NA3        u098(.A(men_men_n120_), .B(men_men_n119_), .C(x06), .Y(men_men_n121_));
  INV        u099(.A(men_men_n121_), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n86_), .B(x13), .Y(men_men_n123_));
  NA2        u101(.A(x09), .B(men_men_n35_), .Y(men_men_n124_));
  NO2        u102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NA2        u103(.A(x13), .B(men_men_n35_), .Y(men_men_n126_));
  NO2        u104(.A(men_men_n126_), .B(x05), .Y(men_men_n127_));
  NO2        u105(.A(men_men_n127_), .B(men_men_n125_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n129_));
  AOI210     u107(.A0(men_men_n57_), .A1(men_men_n82_), .B0(men_men_n118_), .Y(men_men_n130_));
  AOI210     u108(.A0(men_men_n130_), .A1(men_men_n128_), .B0(men_men_n74_), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n132_));
  NA2        u110(.A(x10), .B(men_men_n57_), .Y(men_men_n133_));
  NA2        u111(.A(men_men_n133_), .B(men_men_n132_), .Y(men_men_n134_));
  NA2        u112(.A(men_men_n51_), .B(x05), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n36_), .B(x04), .Y(men_men_n136_));
  NA3        u114(.A(men_men_n136_), .B(men_men_n135_), .C(x13), .Y(men_men_n137_));
  NO3        u115(.A(men_men_n129_), .B(men_men_n81_), .C(men_men_n36_), .Y(men_men_n138_));
  NO2        u116(.A(men_men_n60_), .B(x05), .Y(men_men_n139_));
  NOi41      u117(.An(men_men_n137_), .B(men_men_n139_), .C(men_men_n138_), .D(men_men_n134_), .Y(men_men_n140_));
  NO3        u118(.A(men_men_n140_), .B(x06), .C(x03), .Y(men_men_n141_));
  NO4        u119(.A(men_men_n141_), .B(men_men_n131_), .C(men_men_n122_), .D(men_men_n116_), .Y(men_men_n142_));
  NA2        u120(.A(x13), .B(men_men_n36_), .Y(men_men_n143_));
  OAI210     u121(.A0(men_men_n86_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n144_));
  NA2        u122(.A(men_men_n144_), .B(men_men_n143_), .Y(men_men_n145_));
  NO2        u123(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n146_));
  OA210      u124(.A0(x00), .A1(men_men_n79_), .B0(men_men_n146_), .Y(men_men_n147_));
  NO2        u125(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n29_), .B(x06), .Y(men_men_n149_));
  AN2        u127(.A(men_men_n147_), .B(men_men_n145_), .Y(men_men_n150_));
  NO2        u128(.A(x09), .B(x05), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n151_), .B(men_men_n47_), .Y(men_men_n152_));
  AOI210     u130(.A0(men_men_n152_), .A1(men_men_n112_), .B0(men_men_n49_), .Y(men_men_n153_));
  NA2        u131(.A(x09), .B(x00), .Y(men_men_n154_));
  NA2        u132(.A(men_men_n117_), .B(men_men_n154_), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n78_), .B(men_men_n51_), .Y(men_men_n156_));
  AOI210     u134(.A0(men_men_n156_), .A1(men_men_n155_), .B0(men_men_n149_), .Y(men_men_n157_));
  NO3        u135(.A(men_men_n157_), .B(men_men_n153_), .C(men_men_n150_), .Y(men_men_n158_));
  NO2        u136(.A(x03), .B(x02), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n87_), .B(men_men_n103_), .Y(men_men_n160_));
  OAI210     u138(.A0(men_men_n160_), .A1(men_men_n118_), .B0(men_men_n159_), .Y(men_men_n161_));
  OA210      u139(.A0(men_men_n158_), .A1(x11), .B0(men_men_n161_), .Y(men_men_n162_));
  OAI210     u140(.A0(men_men_n142_), .A1(men_men_n23_), .B0(men_men_n162_), .Y(men_men_n163_));
  NA2        u141(.A(men_men_n112_), .B(men_men_n40_), .Y(men_men_n164_));
  NAi21      u142(.An(x06), .B(x10), .Y(men_men_n165_));
  NOi21      u143(.An(x01), .B(x13), .Y(men_men_n166_));
  NA2        u144(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  OR2        u145(.A(men_men_n167_), .B(x08), .Y(men_men_n168_));
  AOI210     u146(.A0(men_men_n168_), .A1(men_men_n164_), .B0(men_men_n41_), .Y(men_men_n169_));
  NO2        u147(.A(men_men_n29_), .B(x03), .Y(men_men_n170_));
  NA2        u148(.A(men_men_n103_), .B(x01), .Y(men_men_n171_));
  NO2        u149(.A(men_men_n171_), .B(x08), .Y(men_men_n172_));
  OAI210     u150(.A0(x05), .A1(men_men_n172_), .B0(men_men_n51_), .Y(men_men_n173_));
  AOI210     u151(.A0(men_men_n173_), .A1(men_men_n170_), .B0(men_men_n48_), .Y(men_men_n174_));
  AOI210     u152(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n175_));
  OAI210     u153(.A0(men_men_n174_), .A1(men_men_n169_), .B0(men_men_n175_), .Y(men_men_n176_));
  NA2        u154(.A(x04), .B(x02), .Y(men_men_n177_));
  NA2        u155(.A(x10), .B(x05), .Y(men_men_n178_));
  NA2        u156(.A(x09), .B(x06), .Y(men_men_n179_));
  NO2        u157(.A(x09), .B(x01), .Y(men_men_n180_));
  NO3        u158(.A(men_men_n180_), .B(men_men_n110_), .C(men_men_n31_), .Y(men_men_n181_));
  NA2        u159(.A(men_men_n181_), .B(x00), .Y(men_men_n182_));
  NO2        u160(.A(men_men_n117_), .B(x08), .Y(men_men_n183_));
  NA3        u161(.A(men_men_n166_), .B(men_men_n165_), .C(men_men_n51_), .Y(men_men_n184_));
  NA2        u162(.A(men_men_n96_), .B(x05), .Y(men_men_n185_));
  OAI210     u163(.A0(men_men_n185_), .A1(men_men_n120_), .B0(men_men_n184_), .Y(men_men_n186_));
  AOI210     u164(.A0(men_men_n183_), .A1(x06), .B0(men_men_n186_), .Y(men_men_n187_));
  OAI210     u165(.A0(men_men_n187_), .A1(x11), .B0(men_men_n182_), .Y(men_men_n188_));
  NAi21      u166(.An(men_men_n177_), .B(men_men_n188_), .Y(men_men_n189_));
  INV        u167(.A(men_men_n25_), .Y(men_men_n190_));
  NAi21      u168(.An(x13), .B(x00), .Y(men_men_n191_));
  AOI210     u169(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n191_), .Y(men_men_n192_));
  AOI220     u170(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n193_));
  OAI210     u171(.A0(men_men_n178_), .A1(men_men_n35_), .B0(men_men_n193_), .Y(men_men_n194_));
  AN2        u172(.A(men_men_n194_), .B(men_men_n192_), .Y(men_men_n195_));
  NO2        u173(.A(men_men_n97_), .B(x06), .Y(men_men_n196_));
  NO2        u174(.A(men_men_n191_), .B(men_men_n36_), .Y(men_men_n197_));
  INV        u175(.A(men_men_n197_), .Y(men_men_n198_));
  OAI210     u176(.A0(men_men_n198_), .A1(men_men_n179_), .B0(men_men_n74_), .Y(men_men_n199_));
  OAI210     u177(.A0(men_men_n199_), .A1(men_men_n195_), .B0(men_men_n190_), .Y(men_men_n200_));
  NOi21      u178(.An(x09), .B(x00), .Y(men_men_n201_));
  NO3        u179(.A(men_men_n85_), .B(men_men_n201_), .C(men_men_n47_), .Y(men_men_n202_));
  NA2        u180(.A(men_men_n202_), .B(men_men_n133_), .Y(men_men_n203_));
  NA2        u181(.A(x10), .B(x08), .Y(men_men_n204_));
  INV        u182(.A(men_men_n204_), .Y(men_men_n205_));
  NA2        u183(.A(x06), .B(x05), .Y(men_men_n206_));
  OAI210     u184(.A0(men_men_n206_), .A1(men_men_n35_), .B0(men_men_n102_), .Y(men_men_n207_));
  AOI210     u185(.A0(men_men_n205_), .A1(men_men_n58_), .B0(men_men_n207_), .Y(men_men_n208_));
  NA2        u186(.A(men_men_n208_), .B(men_men_n203_), .Y(men_men_n209_));
  NO2        u187(.A(men_men_n103_), .B(x12), .Y(men_men_n210_));
  AOI210     u188(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n210_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n96_), .B(men_men_n51_), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n213_));
  NA2        u191(.A(men_men_n213_), .B(x02), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n214_), .B(men_men_n212_), .Y(men_men_n215_));
  AOI210     u193(.A0(men_men_n211_), .A1(men_men_n209_), .B0(men_men_n215_), .Y(men_men_n216_));
  NA4        u194(.A(men_men_n216_), .B(men_men_n200_), .C(men_men_n189_), .D(men_men_n176_), .Y(men_men_n217_));
  AOI210     u195(.A0(men_men_n163_), .A1(men_men_n102_), .B0(men_men_n217_), .Y(men_men_n218_));
  NA2        u196(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n219_));
  NA2        u197(.A(men_men_n219_), .B(men_men_n144_), .Y(men_men_n220_));
  AOI210     u198(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n221_));
  NO2        u199(.A(men_men_n132_), .B(x06), .Y(men_men_n222_));
  AOI210     u200(.A0(men_men_n221_), .A1(men_men_n220_), .B0(men_men_n222_), .Y(men_men_n223_));
  NO2        u201(.A(men_men_n223_), .B(x12), .Y(men_men_n224_));
  INV        u202(.A(men_men_n78_), .Y(men_men_n225_));
  AOI210     u203(.A0(men_men_n204_), .A1(x05), .B0(men_men_n51_), .Y(men_men_n226_));
  OAI210     u204(.A0(men_men_n226_), .A1(men_men_n167_), .B0(men_men_n57_), .Y(men_men_n227_));
  NA2        u205(.A(men_men_n227_), .B(men_men_n225_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n96_), .B(x06), .Y(men_men_n229_));
  AOI210     u207(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n230_));
  NA4        u208(.A(men_men_n165_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n231_));
  NA2        u209(.A(men_men_n231_), .B(men_men_n149_), .Y(men_men_n232_));
  NA2        u210(.A(men_men_n232_), .B(x02), .Y(men_men_n233_));
  AOI210     u211(.A0(men_men_n233_), .A1(men_men_n228_), .B0(men_men_n23_), .Y(men_men_n234_));
  OAI210     u212(.A0(men_men_n224_), .A1(men_men_n57_), .B0(men_men_n234_), .Y(men_men_n235_));
  INV        u213(.A(men_men_n149_), .Y(men_men_n236_));
  NO2        u214(.A(men_men_n51_), .B(x03), .Y(men_men_n237_));
  OAI210     u215(.A0(men_men_n81_), .A1(men_men_n36_), .B0(men_men_n124_), .Y(men_men_n238_));
  NO2        u216(.A(men_men_n103_), .B(x03), .Y(men_men_n239_));
  AOI220     u217(.A0(men_men_n239_), .A1(men_men_n238_), .B0(men_men_n78_), .B1(men_men_n237_), .Y(men_men_n240_));
  NA2        u218(.A(men_men_n32_), .B(x06), .Y(men_men_n241_));
  INV        u219(.A(men_men_n165_), .Y(men_men_n242_));
  NOi21      u220(.An(x13), .B(x04), .Y(men_men_n243_));
  NO3        u221(.A(men_men_n243_), .B(men_men_n78_), .C(men_men_n201_), .Y(men_men_n244_));
  NO2        u222(.A(men_men_n244_), .B(x05), .Y(men_men_n245_));
  AOI220     u223(.A0(men_men_n245_), .A1(men_men_n241_), .B0(men_men_n242_), .B1(men_men_n57_), .Y(men_men_n246_));
  OAI210     u224(.A0(men_men_n240_), .A1(men_men_n236_), .B0(men_men_n246_), .Y(men_men_n247_));
  INV        u225(.A(men_men_n94_), .Y(men_men_n248_));
  NO2        u226(.A(men_men_n248_), .B(x12), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n250_));
  NO2        u228(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n251_));
  OAI210     u229(.A0(men_men_n251_), .A1(men_men_n194_), .B0(men_men_n192_), .Y(men_men_n252_));
  AOI210     u230(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n253_));
  OAI210     u231(.A0(men_men_n105_), .A1(men_men_n154_), .B0(men_men_n74_), .Y(men_men_n254_));
  INV        u232(.A(men_men_n254_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n256_), .B(x03), .Y(men_men_n257_));
  OA210      u235(.A0(men_men_n257_), .A1(men_men_n255_), .B0(men_men_n252_), .Y(men_men_n258_));
  NA2        u236(.A(x13), .B(men_men_n102_), .Y(men_men_n259_));
  NA3        u237(.A(men_men_n259_), .B(men_men_n207_), .C(men_men_n95_), .Y(men_men_n260_));
  OAI210     u238(.A0(men_men_n258_), .A1(men_men_n250_), .B0(men_men_n260_), .Y(men_men_n261_));
  AOI210     u239(.A0(men_men_n249_), .A1(men_men_n247_), .B0(men_men_n261_), .Y(men_men_n262_));
  AOI210     u240(.A0(men_men_n262_), .A1(men_men_n235_), .B0(x07), .Y(men_men_n263_));
  NA2        u241(.A(men_men_n73_), .B(men_men_n29_), .Y(men_men_n264_));
  BUFFER     u242(.A(men_men_n143_), .Y(men_men_n265_));
  AOI210     u243(.A0(men_men_n265_), .A1(men_men_n156_), .B0(men_men_n264_), .Y(men_men_n266_));
  NO2        u244(.A(men_men_n103_), .B(x06), .Y(men_men_n267_));
  INV        u245(.A(men_men_n267_), .Y(men_men_n268_));
  NO2        u246(.A(x08), .B(x05), .Y(men_men_n269_));
  NO2        u247(.A(men_men_n269_), .B(men_men_n253_), .Y(men_men_n270_));
  OAI210     u248(.A0(men_men_n78_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n271_));
  OAI210     u249(.A0(men_men_n270_), .A1(men_men_n268_), .B0(men_men_n271_), .Y(men_men_n272_));
  NO2        u250(.A(x12), .B(x02), .Y(men_men_n273_));
  INV        u251(.A(men_men_n273_), .Y(men_men_n274_));
  NO2        u252(.A(men_men_n274_), .B(men_men_n248_), .Y(men_men_n275_));
  OA210      u253(.A0(men_men_n272_), .A1(men_men_n266_), .B0(men_men_n275_), .Y(men_men_n276_));
  NA2        u254(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n277_));
  NO2        u255(.A(men_men_n277_), .B(x01), .Y(men_men_n278_));
  NOi21      u256(.An(men_men_n86_), .B(men_men_n124_), .Y(men_men_n279_));
  NO2        u257(.A(men_men_n279_), .B(men_men_n278_), .Y(men_men_n280_));
  AOI210     u258(.A0(men_men_n280_), .A1(men_men_n137_), .B0(men_men_n29_), .Y(men_men_n281_));
  NA2        u259(.A(men_men_n267_), .B(men_men_n238_), .Y(men_men_n282_));
  NA2        u260(.A(men_men_n103_), .B(x04), .Y(men_men_n283_));
  NA2        u261(.A(men_men_n283_), .B(men_men_n28_), .Y(men_men_n284_));
  OAI210     u262(.A0(men_men_n284_), .A1(men_men_n123_), .B0(men_men_n282_), .Y(men_men_n285_));
  NO3        u263(.A(men_men_n93_), .B(x12), .C(x03), .Y(men_men_n286_));
  OAI210     u264(.A0(men_men_n285_), .A1(men_men_n281_), .B0(men_men_n286_), .Y(men_men_n287_));
  AOI210     u265(.A0(men_men_n212_), .A1(men_men_n206_), .B0(men_men_n105_), .Y(men_men_n288_));
  NOi21      u266(.An(men_men_n264_), .B(men_men_n229_), .Y(men_men_n289_));
  NO2        u267(.A(men_men_n25_), .B(x00), .Y(men_men_n290_));
  OAI210     u268(.A0(men_men_n289_), .A1(men_men_n288_), .B0(men_men_n290_), .Y(men_men_n291_));
  NO2        u269(.A(men_men_n58_), .B(x05), .Y(men_men_n292_));
  NO3        u270(.A(men_men_n292_), .B(men_men_n230_), .C(men_men_n196_), .Y(men_men_n293_));
  NO2        u271(.A(men_men_n250_), .B(men_men_n28_), .Y(men_men_n294_));
  OAI210     u272(.A0(men_men_n293_), .A1(men_men_n236_), .B0(men_men_n294_), .Y(men_men_n295_));
  NA3        u273(.A(men_men_n295_), .B(men_men_n291_), .C(men_men_n287_), .Y(men_men_n296_));
  NO3        u274(.A(men_men_n296_), .B(men_men_n276_), .C(men_men_n263_), .Y(men_men_n297_));
  OAI210     u275(.A0(men_men_n218_), .A1(men_men_n61_), .B0(men_men_n297_), .Y(men02));
  NOi21      u276(.An(men_men_n244_), .B(men_men_n180_), .Y(men_men_n299_));
  NA3        u277(.A(x04), .B(men_men_n205_), .C(men_men_n56_), .Y(men_men_n300_));
  OAI210     u278(.A0(men_men_n299_), .A1(men_men_n32_), .B0(men_men_n300_), .Y(men_men_n301_));
  NA2        u279(.A(men_men_n301_), .B(men_men_n178_), .Y(men_men_n302_));
  INV        u280(.A(men_men_n178_), .Y(men_men_n303_));
  AOI210     u281(.A0(men_men_n119_), .A1(men_men_n88_), .B0(men_men_n230_), .Y(men_men_n304_));
  OAI220     u282(.A0(men_men_n304_), .A1(men_men_n103_), .B0(men_men_n87_), .B1(men_men_n51_), .Y(men_men_n305_));
  AOI220     u283(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n160_), .B1(men_men_n159_), .Y(men_men_n306_));
  AOI210     u284(.A0(men_men_n306_), .A1(men_men_n302_), .B0(men_men_n48_), .Y(men_men_n307_));
  NO2        u285(.A(x05), .B(x02), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n220_), .A1(men_men_n201_), .B0(men_men_n308_), .Y(men_men_n309_));
  AOI220     u287(.A0(men_men_n269_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n310_));
  NA2        u288(.A(men_men_n243_), .B(men_men_n81_), .Y(men_men_n311_));
  AOI210     u289(.A0(men_men_n311_), .A1(men_men_n309_), .B0(men_men_n149_), .Y(men_men_n312_));
  NAi21      u290(.An(men_men_n245_), .B(men_men_n240_), .Y(men_men_n313_));
  NO2        u291(.A(men_men_n256_), .B(men_men_n47_), .Y(men_men_n314_));
  NA2        u292(.A(men_men_n314_), .B(men_men_n313_), .Y(men_men_n315_));
  AN2        u293(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n316_));
  OAI210     u294(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n317_));
  NA2        u295(.A(x13), .B(men_men_n28_), .Y(men_men_n318_));
  AOI210     u296(.A0(men_men_n152_), .A1(men_men_n144_), .B0(men_men_n317_), .Y(men_men_n319_));
  OAI210     u297(.A0(men_men_n319_), .A1(men_men_n316_), .B0(men_men_n97_), .Y(men_men_n320_));
  NA3        u298(.A(men_men_n97_), .B(men_men_n86_), .C(men_men_n237_), .Y(men_men_n321_));
  NA3        u299(.A(men_men_n96_), .B(men_men_n85_), .C(men_men_n42_), .Y(men_men_n322_));
  AOI210     u300(.A0(men_men_n322_), .A1(men_men_n321_), .B0(x04), .Y(men_men_n323_));
  INV        u301(.A(men_men_n159_), .Y(men_men_n324_));
  OAI220     u302(.A0(men_men_n270_), .A1(men_men_n108_), .B0(men_men_n324_), .B1(men_men_n134_), .Y(men_men_n325_));
  AOI210     u303(.A0(men_men_n325_), .A1(x13), .B0(men_men_n323_), .Y(men_men_n326_));
  NA3        u304(.A(men_men_n326_), .B(men_men_n320_), .C(men_men_n315_), .Y(men_men_n327_));
  NO3        u305(.A(men_men_n327_), .B(men_men_n312_), .C(men_men_n307_), .Y(men_men_n328_));
  NA2        u306(.A(men_men_n148_), .B(x03), .Y(men_men_n329_));
  INV        u307(.A(men_men_n191_), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n51_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n331_));
  AOI220     u309(.A0(men_men_n331_), .A1(men_men_n330_), .B0(men_men_n213_), .B1(x08), .Y(men_men_n332_));
  OAI210     u310(.A0(men_men_n332_), .A1(men_men_n292_), .B0(men_men_n329_), .Y(men_men_n333_));
  NA2        u311(.A(men_men_n333_), .B(men_men_n110_), .Y(men_men_n334_));
  NA2        u312(.A(men_men_n177_), .B(men_men_n171_), .Y(men_men_n335_));
  AN2        u313(.A(men_men_n335_), .B(men_men_n183_), .Y(men_men_n336_));
  INV        u314(.A(men_men_n56_), .Y(men_men_n337_));
  OAI220     u315(.A0(men_men_n283_), .A1(men_men_n337_), .B0(men_men_n135_), .B1(men_men_n28_), .Y(men_men_n338_));
  OAI210     u316(.A0(men_men_n338_), .A1(men_men_n336_), .B0(men_men_n111_), .Y(men_men_n339_));
  NA2        u317(.A(men_men_n283_), .B(men_men_n102_), .Y(men_men_n340_));
  NA2        u318(.A(men_men_n102_), .B(men_men_n41_), .Y(men_men_n341_));
  NA3        u319(.A(men_men_n341_), .B(men_men_n340_), .C(men_men_n134_), .Y(men_men_n342_));
  NA4        u320(.A(men_men_n342_), .B(men_men_n339_), .C(men_men_n334_), .D(men_men_n48_), .Y(men_men_n343_));
  INV        u321(.A(men_men_n213_), .Y(men_men_n344_));
  NO2        u322(.A(men_men_n172_), .B(men_men_n40_), .Y(men_men_n345_));
  NA2        u323(.A(men_men_n32_), .B(x05), .Y(men_men_n346_));
  OAI220     u324(.A0(men_men_n346_), .A1(men_men_n345_), .B0(men_men_n344_), .B1(men_men_n59_), .Y(men_men_n347_));
  NA2        u325(.A(men_men_n347_), .B(x02), .Y(men_men_n348_));
  INV        u326(.A(men_men_n251_), .Y(men_men_n349_));
  NA2        u327(.A(men_men_n210_), .B(x04), .Y(men_men_n350_));
  NO2        u328(.A(men_men_n350_), .B(men_men_n349_), .Y(men_men_n351_));
  NO3        u329(.A(men_men_n193_), .B(x13), .C(men_men_n31_), .Y(men_men_n352_));
  OAI210     u330(.A0(men_men_n352_), .A1(men_men_n351_), .B0(men_men_n97_), .Y(men_men_n353_));
  NO3        u331(.A(men_men_n210_), .B(men_men_n170_), .C(men_men_n52_), .Y(men_men_n354_));
  OAI210     u332(.A0(men_men_n154_), .A1(men_men_n36_), .B0(men_men_n102_), .Y(men_men_n355_));
  OAI210     u333(.A0(men_men_n355_), .A1(men_men_n202_), .B0(men_men_n354_), .Y(men_men_n356_));
  NA4        u334(.A(men_men_n356_), .B(men_men_n353_), .C(men_men_n348_), .D(x06), .Y(men_men_n357_));
  NA2        u335(.A(x09), .B(x03), .Y(men_men_n358_));
  OAI220     u336(.A0(men_men_n358_), .A1(men_men_n133_), .B0(men_men_n219_), .B1(men_men_n64_), .Y(men_men_n359_));
  OAI220     u337(.A0(men_men_n171_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n360_));
  NO3        u338(.A(men_men_n292_), .B(men_men_n132_), .C(x08), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n360_), .A1(men_men_n236_), .B0(men_men_n361_), .Y(men_men_n362_));
  NO2        u340(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n363_));
  NA2        u341(.A(men_men_n354_), .B(men_men_n363_), .Y(men_men_n364_));
  OAI210     u342(.A0(men_men_n362_), .A1(men_men_n28_), .B0(men_men_n364_), .Y(men_men_n365_));
  AO220      u343(.A0(men_men_n365_), .A1(x04), .B0(men_men_n359_), .B1(x05), .Y(men_men_n366_));
  AOI210     u344(.A0(men_men_n357_), .A1(men_men_n343_), .B0(men_men_n366_), .Y(men_men_n367_));
  OAI210     u345(.A0(men_men_n328_), .A1(x12), .B0(men_men_n367_), .Y(men03));
  OR2        u346(.A(men_men_n42_), .B(men_men_n237_), .Y(men_men_n369_));
  AOI210     u347(.A0(men_men_n160_), .A1(men_men_n102_), .B0(men_men_n369_), .Y(men_men_n370_));
  AO210      u348(.A0(men_men_n349_), .A1(men_men_n88_), .B0(men_men_n350_), .Y(men_men_n371_));
  NA2        u349(.A(men_men_n210_), .B(men_men_n159_), .Y(men_men_n372_));
  NA3        u350(.A(men_men_n372_), .B(men_men_n371_), .C(men_men_n214_), .Y(men_men_n373_));
  OAI210     u351(.A0(men_men_n373_), .A1(men_men_n370_), .B0(x05), .Y(men_men_n374_));
  NA2        u352(.A(men_men_n369_), .B(x05), .Y(men_men_n375_));
  AOI210     u353(.A0(men_men_n144_), .A1(men_men_n225_), .B0(men_men_n375_), .Y(men_men_n376_));
  AOI210     u354(.A0(men_men_n239_), .A1(men_men_n82_), .B0(men_men_n127_), .Y(men_men_n377_));
  OAI220     u355(.A0(men_men_n377_), .A1(men_men_n59_), .B0(men_men_n318_), .B1(men_men_n310_), .Y(men_men_n378_));
  OAI210     u356(.A0(men_men_n378_), .A1(men_men_n376_), .B0(men_men_n102_), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n152_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n380_));
  NO2        u358(.A(men_men_n180_), .B(men_men_n139_), .Y(men_men_n381_));
  OAI220     u359(.A0(men_men_n381_), .A1(men_men_n37_), .B0(men_men_n155_), .B1(x13), .Y(men_men_n382_));
  OAI210     u360(.A0(men_men_n382_), .A1(men_men_n380_), .B0(x04), .Y(men_men_n383_));
  NO3        u361(.A(men_men_n341_), .B(men_men_n87_), .C(men_men_n59_), .Y(men_men_n384_));
  AOI210     u362(.A0(men_men_n198_), .A1(men_men_n102_), .B0(men_men_n152_), .Y(men_men_n385_));
  OA210      u363(.A0(men_men_n172_), .A1(x12), .B0(men_men_n139_), .Y(men_men_n386_));
  NO3        u364(.A(men_men_n386_), .B(men_men_n385_), .C(men_men_n384_), .Y(men_men_n387_));
  NA4        u365(.A(men_men_n387_), .B(men_men_n383_), .C(men_men_n379_), .D(men_men_n374_), .Y(men04));
  NO2        u366(.A(men_men_n91_), .B(men_men_n39_), .Y(men_men_n389_));
  XO2        u367(.A(men_men_n389_), .B(men_men_n259_), .Y(men05));
  INV        u368(.A(men_men_n222_), .Y(men_men_n391_));
  AOI210     u369(.A0(men_men_n391_), .A1(men_men_n317_), .B0(men_men_n25_), .Y(men_men_n392_));
  NAi41      u370(.An(men_men_n79_), .B(men_men_n149_), .C(men_men_n135_), .D(men_men_n31_), .Y(men_men_n393_));
  INV        u371(.A(men_men_n92_), .Y(men_men_n394_));
  AOI210     u372(.A0(men_men_n394_), .A1(men_men_n393_), .B0(men_men_n24_), .Y(men_men_n395_));
  OAI210     u373(.A0(men_men_n395_), .A1(men_men_n392_), .B0(men_men_n102_), .Y(men_men_n396_));
  NA2        u374(.A(x11), .B(men_men_n31_), .Y(men_men_n397_));
  NA2        u375(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n398_));
  NA2        u376(.A(men_men_n264_), .B(x03), .Y(men_men_n399_));
  OAI220     u377(.A0(men_men_n399_), .A1(men_men_n398_), .B0(men_men_n397_), .B1(men_men_n83_), .Y(men_men_n400_));
  OAI210     u378(.A0(men_men_n26_), .A1(men_men_n102_), .B0(x07), .Y(men_men_n401_));
  AOI210     u379(.A0(men_men_n400_), .A1(x06), .B0(men_men_n401_), .Y(men_men_n402_));
  AOI220     u380(.A0(men_men_n83_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n403_));
  NO3        u381(.A(men_men_n403_), .B(men_men_n23_), .C(x00), .Y(men_men_n404_));
  NA2        u382(.A(men_men_n71_), .B(x02), .Y(men_men_n405_));
  AOI210     u383(.A0(men_men_n405_), .A1(men_men_n399_), .B0(men_men_n267_), .Y(men_men_n406_));
  OR2        u384(.A(men_men_n406_), .B(men_men_n250_), .Y(men_men_n407_));
  NO2        u385(.A(men_men_n23_), .B(x10), .Y(men_men_n408_));
  OAI210     u386(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n409_));
  OR3        u387(.A(men_men_n409_), .B(men_men_n408_), .C(men_men_n44_), .Y(men_men_n410_));
  NA2        u388(.A(men_men_n410_), .B(men_men_n407_), .Y(men_men_n411_));
  OAI210     u389(.A0(men_men_n411_), .A1(men_men_n404_), .B0(men_men_n102_), .Y(men_men_n412_));
  NA2        u390(.A(men_men_n33_), .B(men_men_n102_), .Y(men_men_n413_));
  AOI210     u391(.A0(men_men_n413_), .A1(men_men_n94_), .B0(x07), .Y(men_men_n414_));
  AOI220     u392(.A0(men_men_n414_), .A1(men_men_n412_), .B0(men_men_n402_), .B1(men_men_n396_), .Y(men_men_n415_));
  NA3        u393(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n416_));
  AO210      u394(.A0(men_men_n416_), .A1(men_men_n277_), .B0(men_men_n274_), .Y(men_men_n417_));
  AOI210     u395(.A0(men_men_n408_), .A1(men_men_n76_), .B0(men_men_n148_), .Y(men_men_n418_));
  OR2        u396(.A(men_men_n418_), .B(x03), .Y(men_men_n419_));
  NA2        u397(.A(men_men_n363_), .B(men_men_n61_), .Y(men_men_n420_));
  NO2        u398(.A(men_men_n420_), .B(x11), .Y(men_men_n421_));
  NO3        u399(.A(men_men_n421_), .B(men_men_n151_), .C(men_men_n28_), .Y(men_men_n422_));
  AOI220     u400(.A0(men_men_n422_), .A1(men_men_n419_), .B0(men_men_n417_), .B1(men_men_n47_), .Y(men_men_n423_));
  NO4        u401(.A(men_men_n341_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n424_));
  OAI210     u402(.A0(men_men_n424_), .A1(men_men_n423_), .B0(men_men_n103_), .Y(men_men_n425_));
  AOI210     u403(.A0(men_men_n350_), .A1(men_men_n113_), .B0(men_men_n273_), .Y(men_men_n426_));
  NOi21      u404(.An(men_men_n329_), .B(men_men_n139_), .Y(men_men_n427_));
  NO2        u405(.A(men_men_n427_), .B(men_men_n274_), .Y(men_men_n428_));
  OAI210     u406(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n429_));
  AOI210     u407(.A0(men_men_n259_), .A1(men_men_n47_), .B0(men_men_n429_), .Y(men_men_n430_));
  NO4        u408(.A(men_men_n430_), .B(men_men_n428_), .C(men_men_n426_), .D(x08), .Y(men_men_n431_));
  AOI210     u409(.A0(men_men_n408_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n432_));
  NA2        u410(.A(x09), .B(men_men_n41_), .Y(men_men_n433_));
  OAI220     u411(.A0(men_men_n433_), .A1(men_men_n432_), .B0(men_men_n397_), .B1(men_men_n67_), .Y(men_men_n434_));
  NO2        u412(.A(x13), .B(x12), .Y(men_men_n435_));
  NO2        u413(.A(men_men_n135_), .B(men_men_n28_), .Y(men_men_n436_));
  NO2        u414(.A(men_men_n436_), .B(men_men_n278_), .Y(men_men_n437_));
  OR3        u415(.A(men_men_n437_), .B(x12), .C(x03), .Y(men_men_n438_));
  NA3        u416(.A(men_men_n344_), .B(men_men_n129_), .C(x12), .Y(men_men_n439_));
  AO210      u417(.A0(men_men_n344_), .A1(men_men_n129_), .B0(men_men_n259_), .Y(men_men_n440_));
  NA4        u418(.A(men_men_n440_), .B(men_men_n439_), .C(men_men_n438_), .D(x08), .Y(men_men_n441_));
  AOI210     u419(.A0(men_men_n435_), .A1(men_men_n434_), .B0(men_men_n441_), .Y(men_men_n442_));
  AOI210     u420(.A0(men_men_n431_), .A1(men_men_n425_), .B0(men_men_n442_), .Y(men_men_n443_));
  OAI210     u421(.A0(men_men_n420_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n444_));
  NA2        u422(.A(men_men_n303_), .B(x07), .Y(men_men_n445_));
  OAI220     u423(.A0(men_men_n445_), .A1(men_men_n398_), .B0(men_men_n151_), .B1(men_men_n43_), .Y(men_men_n446_));
  OAI210     u424(.A0(men_men_n446_), .A1(men_men_n444_), .B0(men_men_n197_), .Y(men_men_n447_));
  NA3        u425(.A(men_men_n437_), .B(men_men_n427_), .C(men_men_n340_), .Y(men_men_n448_));
  INV        u426(.A(x14), .Y(men_men_n449_));
  NO3        u427(.A(men_men_n329_), .B(men_men_n108_), .C(x11), .Y(men_men_n450_));
  NO3        u428(.A(men_men_n171_), .B(men_men_n76_), .C(men_men_n57_), .Y(men_men_n451_));
  NO3        u429(.A(men_men_n416_), .B(men_men_n341_), .C(men_men_n191_), .Y(men_men_n452_));
  NO4        u430(.A(men_men_n452_), .B(men_men_n451_), .C(men_men_n450_), .D(men_men_n449_), .Y(men_men_n453_));
  NA3        u431(.A(men_men_n453_), .B(men_men_n448_), .C(men_men_n447_), .Y(men_men_n454_));
  AOI220     u432(.A0(men_men_n413_), .A1(men_men_n61_), .B0(men_men_n436_), .B1(men_men_n170_), .Y(men_men_n455_));
  NOi21      u433(.An(men_men_n283_), .B(men_men_n155_), .Y(men_men_n456_));
  NA2        u434(.A(men_men_n290_), .B(men_men_n242_), .Y(men_men_n457_));
  OAI210     u435(.A0(men_men_n44_), .A1(x04), .B0(men_men_n457_), .Y(men_men_n458_));
  OAI210     u436(.A0(men_men_n458_), .A1(men_men_n456_), .B0(men_men_n102_), .Y(men_men_n459_));
  OAI210     u437(.A0(men_men_n455_), .A1(men_men_n93_), .B0(men_men_n459_), .Y(men_men_n460_));
  NO4        u438(.A(men_men_n460_), .B(men_men_n454_), .C(men_men_n443_), .D(men_men_n415_), .Y(men06));
  INV        u439(.A(x07), .Y(men_men_n464_));
  INV        u440(.A(men_men_n95_), .Y(men_men_n465_));
  INV        u441(.A(x01), .Y(men_men_n466_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule