//Benchmark atmr_5xp1_76_0.0156

module atmr_5xp1(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
 wire ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n65_, ori_ori_n69_, ori_ori_n70_, ori_ori_n72_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n65_, mai_mai_n69_, mai_mai_n70_, mai_mai_n72_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n65_, men_men_n69_, men_men_n70_, men_men_n72_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09;
  INV        o00(.A(i_5_), .Y(ori_ori_n18_));
  NO3        o01(.A(i_4_), .B(i_6_), .C(ori_ori_n18_), .Y(ori_ori_n19_));
  INV        o02(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o03(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n21_));
  INV        o04(.A(i_1_), .Y(ori_ori_n22_));
  AOI210     o05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(ori_ori_n23_));
  NA2        o06(.A(ori_ori_n23_), .B(ori_ori_n22_), .Y(ori_ori_n24_));
  NO2        o07(.A(ori_ori_n24_), .B(ori_ori_n21_), .Y(ori_ori_n25_));
  INV        o08(.A(i_6_), .Y(ori_ori_n26_));
  NO2        o09(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n27_));
  INV        o10(.A(i_0_), .Y(ori_ori_n28_));
  NO2        o11(.A(i_2_), .B(i_1_), .Y(ori_ori_n29_));
  OAI210     o12(.A0(ori_ori_n29_), .A1(ori_ori_n28_), .B0(ori_ori_n20_), .Y(ori_ori_n30_));
  NO2        o13(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n31_));
  NO2        o14(.A(i_2_), .B(i_3_), .Y(ori_ori_n32_));
  NO3        o15(.A(ori_ori_n32_), .B(ori_ori_n28_), .C(ori_ori_n22_), .Y(ori_ori_n33_));
  AO220      o16(.A0(ori_ori_n33_), .A1(ori_ori_n31_), .B0(ori_ori_n30_), .B1(ori_ori_n27_), .Y(ori_ori_n34_));
  NA2        o17(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n35_));
  NA2        o18(.A(i_2_), .B(i_3_), .Y(ori_ori_n36_));
  NO2        o19(.A(ori_ori_n36_), .B(ori_ori_n22_), .Y(ori_ori_n37_));
  NO3        o20(.A(ori_ori_n37_), .B(ori_ori_n35_), .C(i_0_), .Y(ori_ori_n38_));
  OR4        o21(.A(ori_ori_n38_), .B(ori_ori_n34_), .C(ori_ori_n25_), .D(ori_ori_n19_), .Y(ori01));
  OR2        o22(.A(i_2_), .B(i_3_), .Y(ori_ori_n40_));
  NA3        o23(.A(ori_ori_n40_), .B(i_0_), .C(i_1_), .Y(ori_ori_n41_));
  NA2        o24(.A(ori_ori_n28_), .B(ori_ori_n18_), .Y(ori_ori_n42_));
  AOI210     o25(.A0(ori_ori_n23_), .A1(ori_ori_n22_), .B0(ori_ori_n26_), .Y(ori_ori_n43_));
  AOI220     o26(.A0(ori_ori_n43_), .A1(ori_ori_n42_), .B0(ori_ori_n41_), .B1(ori_ori_n26_), .Y(ori_ori_n44_));
  NA2        o27(.A(ori_ori_n29_), .B(ori_ori_n18_), .Y(ori_ori_n45_));
  OAI220     o28(.A0(ori_ori_n45_), .A1(ori_ori_n26_), .B0(ori_ori_n35_), .B1(ori_ori_n28_), .Y(ori_ori_n46_));
  NO3        o29(.A(ori_ori_n46_), .B(ori_ori_n44_), .C(i_4_), .Y(ori_ori_n47_));
  NA2        o30(.A(i_0_), .B(i_6_), .Y(ori_ori_n48_));
  OAI210     o31(.A0(i_0_), .A1(i_1_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  NOi31      o32(.An(ori_ori_n49_), .B(ori_ori_n23_), .C(ori_ori_n18_), .Y(ori_ori_n50_));
  NA3        o33(.A(i_1_), .B(i_6_), .C(i_5_), .Y(ori_ori_n51_));
  AOI210     o34(.A0(ori_ori_n51_), .A1(ori_ori_n48_), .B0(ori_ori_n29_), .Y(ori_ori_n52_));
  NO3        o35(.A(ori_ori_n40_), .B(i_6_), .C(i_5_), .Y(ori_ori_n53_));
  NO3        o36(.A(ori_ori_n52_), .B(ori_ori_n50_), .C(ori_ori_n20_), .Y(ori_ori_n54_));
  NA2        o37(.A(ori_ori_n28_), .B(ori_ori_n26_), .Y(ori_ori_n55_));
  NO2        o38(.A(ori_ori_n55_), .B(ori_ori_n20_), .Y(ori_ori_n56_));
  AOI210     o39(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(ori_ori_n57_));
  AO220      o40(.A0(ori_ori_n57_), .A1(ori_ori_n31_), .B0(ori_ori_n37_), .B1(ori_ori_n19_), .Y(ori_ori_n58_));
  AOI210     o41(.A0(ori_ori_n56_), .A1(ori_ori_n36_), .B0(ori_ori_n58_), .Y(ori_ori_n59_));
  OAI210     o42(.A0(ori_ori_n54_), .A1(ori_ori_n47_), .B0(ori_ori_n59_), .Y(ori02));
  NAi21      o43(.An(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n61_));
  NA3        o44(.A(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n62_));
  AOI210     o45(.A0(ori_ori_n56_), .A1(ori_ori_n62_), .B0(ori_ori_n31_), .Y(ori_ori_n63_));
  NA2        o46(.A(ori_ori_n63_), .B(ori_ori_n61_), .Y(ori00));
  OAI210     o47(.A0(ori_ori_n55_), .A1(ori_ori_n37_), .B0(i_5_), .Y(ori_ori_n65_));
  NO2        o48(.A(ori_ori_n65_), .B(ori_ori_n20_), .Y(ori09));
  NOi21      o49(.An(ori_ori_n36_), .B(ori_ori_n32_), .Y(ori07));
  INV        o50(.A(i_3_), .Y(ori08));
  INV        o51(.A(ori_ori_n29_), .Y(ori_ori_n69_));
  NA2        o52(.A(ori07), .B(ori_ori_n69_), .Y(ori_ori_n70_));
  XO2        o53(.A(ori_ori_n70_), .B(ori_ori_n28_), .Y(ori05));
  NO2        o54(.A(i_2_), .B(ori08), .Y(ori_ori_n72_));
  XO2        o55(.A(ori_ori_n72_), .B(i_1_), .Y(ori06));
  NAi21      o56(.An(ori_ori_n53_), .B(ori_ori_n45_), .Y(ori_ori_n74_));
  NA2        o57(.A(ori_ori_n74_), .B(i_0_), .Y(ori_ori_n75_));
  NO2        o58(.A(i_1_), .B(i_6_), .Y(ori_ori_n76_));
  NO3        o59(.A(ori_ori_n76_), .B(ori_ori_n42_), .C(ori_ori_n36_), .Y(ori_ori_n77_));
  NO2        o60(.A(ori_ori_n77_), .B(ori_ori_n38_), .Y(ori_ori_n78_));
  AO210      o61(.A0(ori_ori_n41_), .A1(ori_ori_n24_), .B0(ori_ori_n18_), .Y(ori_ori_n79_));
  NO2        o62(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n80_));
  NO2        o63(.A(ori_ori_n26_), .B(ori_ori_n18_), .Y(ori_ori_n81_));
  OAI210     o64(.A0(ori_ori_n22_), .A1(i_6_), .B0(ori_ori_n18_), .Y(ori_ori_n82_));
  NO2        o65(.A(ori_ori_n82_), .B(ori_ori_n49_), .Y(ori_ori_n83_));
  AOI210     o66(.A0(ori_ori_n81_), .A1(ori_ori_n80_), .B0(ori_ori_n83_), .Y(ori_ori_n84_));
  NA4        o67(.A(ori_ori_n84_), .B(ori_ori_n79_), .C(ori_ori_n78_), .D(ori_ori_n75_), .Y(ori03));
  NA2        o68(.A(ori_ori_n28_), .B(ori08), .Y(ori_ori_n86_));
  OAI210     o69(.A0(ori_ori_n86_), .A1(i_1_), .B0(ori_ori_n62_), .Y(ori_ori_n87_));
  OAI210     o70(.A0(ori_ori_n87_), .A1(ori_ori_n33_), .B0(i_6_), .Y(ori_ori_n88_));
  AOI210     o71(.A0(ori_ori_n32_), .A1(ori_ori_n26_), .B0(ori_ori_n29_), .Y(ori_ori_n89_));
  OR2        o72(.A(ori_ori_n89_), .B(ori_ori_n76_), .Y(ori_ori_n90_));
  NA3        o73(.A(ori_ori_n86_), .B(ori_ori_n76_), .C(i_2_), .Y(ori_ori_n91_));
  NA3        o74(.A(ori_ori_n23_), .B(i_1_), .C(ori_ori_n26_), .Y(ori_ori_n92_));
  NA4        o75(.A(ori_ori_n92_), .B(ori_ori_n91_), .C(ori_ori_n90_), .D(ori_ori_n88_), .Y(ori04));
  INV        m00(.A(i_5_), .Y(mai_mai_n18_));
  NO3        m01(.A(i_4_), .B(i_6_), .C(mai_mai_n18_), .Y(mai_mai_n19_));
  INV        m02(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m03(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n21_));
  INV        m04(.A(i_1_), .Y(mai_mai_n22_));
  AOI210     m05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(mai_mai_n23_));
  NA2        m06(.A(mai_mai_n23_), .B(mai_mai_n22_), .Y(mai_mai_n24_));
  NO2        m07(.A(mai_mai_n24_), .B(mai_mai_n21_), .Y(mai_mai_n25_));
  INV        m08(.A(i_6_), .Y(mai_mai_n26_));
  NO2        m09(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n27_));
  INV        m10(.A(i_0_), .Y(mai_mai_n28_));
  NO2        m11(.A(i_2_), .B(i_1_), .Y(mai_mai_n29_));
  OAI210     m12(.A0(mai_mai_n29_), .A1(mai_mai_n28_), .B0(mai_mai_n20_), .Y(mai_mai_n30_));
  NO2        m13(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n31_));
  NO2        m14(.A(i_2_), .B(i_3_), .Y(mai_mai_n32_));
  NO3        m15(.A(mai_mai_n32_), .B(mai_mai_n28_), .C(mai_mai_n22_), .Y(mai_mai_n33_));
  AO220      m16(.A0(mai_mai_n33_), .A1(mai_mai_n31_), .B0(mai_mai_n30_), .B1(mai_mai_n27_), .Y(mai_mai_n34_));
  NA2        m17(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n35_));
  NA2        m18(.A(i_2_), .B(i_3_), .Y(mai_mai_n36_));
  NO2        m19(.A(mai_mai_n36_), .B(mai_mai_n22_), .Y(mai_mai_n37_));
  NO3        m20(.A(mai_mai_n37_), .B(mai_mai_n35_), .C(i_0_), .Y(mai_mai_n38_));
  OR4        m21(.A(mai_mai_n38_), .B(mai_mai_n34_), .C(mai_mai_n25_), .D(mai_mai_n19_), .Y(mai01));
  OR2        m22(.A(i_2_), .B(i_3_), .Y(mai_mai_n40_));
  NA3        m23(.A(mai_mai_n40_), .B(i_0_), .C(i_1_), .Y(mai_mai_n41_));
  NA2        m24(.A(mai_mai_n28_), .B(mai_mai_n18_), .Y(mai_mai_n42_));
  AOI210     m25(.A0(mai_mai_n23_), .A1(mai_mai_n22_), .B0(mai_mai_n26_), .Y(mai_mai_n43_));
  AOI220     m26(.A0(mai_mai_n43_), .A1(mai_mai_n42_), .B0(mai_mai_n41_), .B1(mai_mai_n26_), .Y(mai_mai_n44_));
  NA2        m27(.A(mai_mai_n29_), .B(mai_mai_n18_), .Y(mai_mai_n45_));
  OAI220     m28(.A0(mai_mai_n45_), .A1(mai_mai_n26_), .B0(mai_mai_n35_), .B1(mai_mai_n28_), .Y(mai_mai_n46_));
  NO3        m29(.A(mai_mai_n46_), .B(mai_mai_n44_), .C(i_4_), .Y(mai_mai_n47_));
  NA2        m30(.A(i_0_), .B(i_6_), .Y(mai_mai_n48_));
  OAI210     m31(.A0(i_0_), .A1(i_1_), .B0(mai_mai_n48_), .Y(mai_mai_n49_));
  NOi31      m32(.An(mai_mai_n49_), .B(mai_mai_n23_), .C(mai_mai_n18_), .Y(mai_mai_n50_));
  NA3        m33(.A(i_1_), .B(i_6_), .C(i_5_), .Y(mai_mai_n51_));
  AOI210     m34(.A0(mai_mai_n51_), .A1(mai_mai_n48_), .B0(mai_mai_n29_), .Y(mai_mai_n52_));
  NO3        m35(.A(mai_mai_n40_), .B(i_6_), .C(i_5_), .Y(mai_mai_n53_));
  NO4        m36(.A(mai_mai_n53_), .B(mai_mai_n52_), .C(mai_mai_n50_), .D(mai_mai_n20_), .Y(mai_mai_n54_));
  NA2        m37(.A(mai_mai_n28_), .B(mai_mai_n26_), .Y(mai_mai_n55_));
  NO2        m38(.A(mai_mai_n55_), .B(mai_mai_n20_), .Y(mai_mai_n56_));
  AOI210     m39(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(mai_mai_n57_));
  AO220      m40(.A0(mai_mai_n57_), .A1(mai_mai_n31_), .B0(mai_mai_n37_), .B1(mai_mai_n19_), .Y(mai_mai_n58_));
  NO2        m41(.A(mai_mai_n56_), .B(mai_mai_n58_), .Y(mai_mai_n59_));
  OAI210     m42(.A0(mai_mai_n54_), .A1(mai_mai_n47_), .B0(mai_mai_n59_), .Y(mai02));
  NAi21      m43(.An(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n61_));
  NA3        m44(.A(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n62_));
  NO2        m45(.A(mai_mai_n56_), .B(mai_mai_n31_), .Y(mai_mai_n63_));
  NA2        m46(.A(mai_mai_n63_), .B(mai_mai_n61_), .Y(mai00));
  NA2        m47(.A(mai_mai_n55_), .B(i_5_), .Y(mai_mai_n65_));
  NO2        m48(.A(mai_mai_n65_), .B(mai_mai_n20_), .Y(mai09));
  NOi21      m49(.An(mai_mai_n36_), .B(mai_mai_n32_), .Y(mai07));
  INV        m50(.A(i_3_), .Y(mai08));
  INV        m51(.A(mai_mai_n29_), .Y(mai_mai_n69_));
  NA2        m52(.A(mai07), .B(mai_mai_n69_), .Y(mai_mai_n70_));
  XO2        m53(.A(mai_mai_n70_), .B(mai_mai_n28_), .Y(mai05));
  NO2        m54(.A(i_2_), .B(mai08), .Y(mai_mai_n72_));
  XO2        m55(.A(mai_mai_n72_), .B(i_1_), .Y(mai06));
  NAi21      m56(.An(mai_mai_n53_), .B(mai_mai_n45_), .Y(mai_mai_n74_));
  NA2        m57(.A(mai_mai_n74_), .B(i_0_), .Y(mai_mai_n75_));
  NO2        m58(.A(i_1_), .B(i_6_), .Y(mai_mai_n76_));
  NO3        m59(.A(mai_mai_n76_), .B(mai_mai_n42_), .C(mai_mai_n36_), .Y(mai_mai_n77_));
  NO2        m60(.A(mai_mai_n77_), .B(mai_mai_n38_), .Y(mai_mai_n78_));
  AO210      m61(.A0(mai_mai_n41_), .A1(mai_mai_n24_), .B0(mai_mai_n18_), .Y(mai_mai_n79_));
  NO2        m62(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n80_));
  NO2        m63(.A(mai_mai_n26_), .B(mai_mai_n18_), .Y(mai_mai_n81_));
  OAI210     m64(.A0(mai_mai_n22_), .A1(i_6_), .B0(mai_mai_n18_), .Y(mai_mai_n82_));
  NO2        m65(.A(mai_mai_n82_), .B(mai_mai_n49_), .Y(mai_mai_n83_));
  AOI210     m66(.A0(mai_mai_n81_), .A1(mai_mai_n80_), .B0(mai_mai_n83_), .Y(mai_mai_n84_));
  NA4        m67(.A(mai_mai_n84_), .B(mai_mai_n79_), .C(mai_mai_n78_), .D(mai_mai_n75_), .Y(mai03));
  NA2        m68(.A(mai_mai_n28_), .B(mai08), .Y(mai_mai_n86_));
  OAI210     m69(.A0(mai_mai_n86_), .A1(i_1_), .B0(mai_mai_n62_), .Y(mai_mai_n87_));
  OAI210     m70(.A0(mai_mai_n87_), .A1(mai_mai_n33_), .B0(i_6_), .Y(mai_mai_n88_));
  AOI210     m71(.A0(mai_mai_n32_), .A1(mai_mai_n26_), .B0(mai_mai_n29_), .Y(mai_mai_n89_));
  OR2        m72(.A(mai_mai_n89_), .B(mai_mai_n76_), .Y(mai_mai_n90_));
  NA3        m73(.A(mai_mai_n86_), .B(mai_mai_n76_), .C(i_2_), .Y(mai_mai_n91_));
  NA3        m74(.A(mai_mai_n23_), .B(i_1_), .C(mai_mai_n26_), .Y(mai_mai_n92_));
  NA4        m75(.A(mai_mai_n92_), .B(mai_mai_n91_), .C(mai_mai_n90_), .D(mai_mai_n88_), .Y(mai04));
  INV        u00(.A(i_5_), .Y(men_men_n18_));
  NO3        u01(.A(i_4_), .B(i_6_), .C(men_men_n18_), .Y(men_men_n19_));
  INV        u02(.A(i_4_), .Y(men_men_n20_));
  NA2        u03(.A(men_men_n20_), .B(i_5_), .Y(men_men_n21_));
  INV        u04(.A(i_1_), .Y(men_men_n22_));
  AOI210     u05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(men_men_n23_));
  NA2        u06(.A(men_men_n23_), .B(men_men_n22_), .Y(men_men_n24_));
  NO2        u07(.A(men_men_n24_), .B(men_men_n21_), .Y(men_men_n25_));
  INV        u08(.A(i_6_), .Y(men_men_n26_));
  NO2        u09(.A(men_men_n26_), .B(i_5_), .Y(men_men_n27_));
  INV        u10(.A(i_0_), .Y(men_men_n28_));
  NO2        u11(.A(i_2_), .B(i_1_), .Y(men_men_n29_));
  OAI210     u12(.A0(men_men_n29_), .A1(men_men_n28_), .B0(men_men_n20_), .Y(men_men_n30_));
  NO2        u13(.A(men_men_n20_), .B(i_5_), .Y(men_men_n31_));
  NO2        u14(.A(i_2_), .B(i_3_), .Y(men_men_n32_));
  NO3        u15(.A(men_men_n32_), .B(men_men_n28_), .C(men_men_n22_), .Y(men_men_n33_));
  AO220      u16(.A0(men_men_n33_), .A1(men_men_n31_), .B0(men_men_n30_), .B1(men_men_n27_), .Y(men_men_n34_));
  NA2        u17(.A(men_men_n26_), .B(i_5_), .Y(men_men_n35_));
  NA2        u18(.A(i_2_), .B(i_3_), .Y(men_men_n36_));
  NO2        u19(.A(men_men_n36_), .B(men_men_n22_), .Y(men_men_n37_));
  NO3        u20(.A(men_men_n37_), .B(men_men_n35_), .C(i_0_), .Y(men_men_n38_));
  OR4        u21(.A(men_men_n38_), .B(men_men_n34_), .C(men_men_n25_), .D(men_men_n19_), .Y(men01));
  OR2        u22(.A(i_2_), .B(i_3_), .Y(men_men_n40_));
  NA3        u23(.A(men_men_n40_), .B(i_0_), .C(i_1_), .Y(men_men_n41_));
  NA2        u24(.A(men_men_n28_), .B(men_men_n18_), .Y(men_men_n42_));
  AOI210     u25(.A0(men_men_n23_), .A1(men_men_n22_), .B0(men_men_n26_), .Y(men_men_n43_));
  AOI220     u26(.A0(men_men_n43_), .A1(men_men_n42_), .B0(men_men_n41_), .B1(men_men_n26_), .Y(men_men_n44_));
  NA2        u27(.A(men_men_n29_), .B(men_men_n18_), .Y(men_men_n45_));
  OAI220     u28(.A0(men_men_n45_), .A1(men_men_n26_), .B0(men_men_n35_), .B1(men_men_n28_), .Y(men_men_n46_));
  NO3        u29(.A(men_men_n46_), .B(men_men_n44_), .C(i_4_), .Y(men_men_n47_));
  NA2        u30(.A(i_0_), .B(i_6_), .Y(men_men_n48_));
  OAI210     u31(.A0(i_0_), .A1(i_1_), .B0(men_men_n48_), .Y(men_men_n49_));
  NOi31      u32(.An(men_men_n49_), .B(men_men_n23_), .C(men_men_n18_), .Y(men_men_n50_));
  NA3        u33(.A(i_1_), .B(i_6_), .C(i_5_), .Y(men_men_n51_));
  AOI210     u34(.A0(men_men_n51_), .A1(men_men_n48_), .B0(men_men_n29_), .Y(men_men_n52_));
  NO3        u35(.A(men_men_n40_), .B(i_6_), .C(i_5_), .Y(men_men_n53_));
  NO4        u36(.A(men_men_n53_), .B(men_men_n52_), .C(men_men_n50_), .D(men_men_n20_), .Y(men_men_n54_));
  NA2        u37(.A(men_men_n28_), .B(men_men_n26_), .Y(men_men_n55_));
  NO2        u38(.A(men_men_n55_), .B(men_men_n20_), .Y(men_men_n56_));
  AOI210     u39(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(men_men_n57_));
  AO220      u40(.A0(men_men_n57_), .A1(men_men_n31_), .B0(men_men_n37_), .B1(men_men_n19_), .Y(men_men_n58_));
  AOI210     u41(.A0(men_men_n56_), .A1(men_men_n36_), .B0(men_men_n58_), .Y(men_men_n59_));
  OAI210     u42(.A0(men_men_n54_), .A1(men_men_n47_), .B0(men_men_n59_), .Y(men02));
  NAi21      u43(.An(men_men_n21_), .B(men_men_n43_), .Y(men_men_n61_));
  NA3        u44(.A(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n62_));
  AOI210     u45(.A0(men_men_n56_), .A1(men_men_n62_), .B0(men_men_n31_), .Y(men_men_n63_));
  NA2        u46(.A(men_men_n63_), .B(men_men_n61_), .Y(men00));
  OAI210     u47(.A0(men_men_n55_), .A1(men_men_n37_), .B0(i_5_), .Y(men_men_n65_));
  NO2        u48(.A(men_men_n65_), .B(men_men_n20_), .Y(men09));
  NOi21      u49(.An(men_men_n36_), .B(men_men_n32_), .Y(men07));
  INV        u50(.A(i_3_), .Y(men08));
  INV        u51(.A(men_men_n29_), .Y(men_men_n69_));
  NA2        u52(.A(men07), .B(men_men_n69_), .Y(men_men_n70_));
  XO2        u53(.A(men_men_n70_), .B(men_men_n28_), .Y(men05));
  NO2        u54(.A(i_2_), .B(men08), .Y(men_men_n72_));
  XO2        u55(.A(men_men_n72_), .B(i_1_), .Y(men06));
  NAi21      u56(.An(men_men_n53_), .B(men_men_n45_), .Y(men_men_n74_));
  NA2        u57(.A(men_men_n74_), .B(i_0_), .Y(men_men_n75_));
  NO2        u58(.A(i_1_), .B(i_6_), .Y(men_men_n76_));
  NO3        u59(.A(men_men_n76_), .B(men_men_n42_), .C(men_men_n36_), .Y(men_men_n77_));
  NO2        u60(.A(men_men_n77_), .B(men_men_n38_), .Y(men_men_n78_));
  AO210      u61(.A0(men_men_n41_), .A1(men_men_n24_), .B0(men_men_n18_), .Y(men_men_n79_));
  NO2        u62(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n80_));
  NO2        u63(.A(men_men_n26_), .B(men_men_n18_), .Y(men_men_n81_));
  OAI210     u64(.A0(men_men_n22_), .A1(i_6_), .B0(men_men_n18_), .Y(men_men_n82_));
  NO2        u65(.A(men_men_n82_), .B(men_men_n49_), .Y(men_men_n83_));
  AOI210     u66(.A0(men_men_n81_), .A1(men_men_n80_), .B0(men_men_n83_), .Y(men_men_n84_));
  NA4        u67(.A(men_men_n84_), .B(men_men_n79_), .C(men_men_n78_), .D(men_men_n75_), .Y(men03));
  NA2        u68(.A(men_men_n28_), .B(men08), .Y(men_men_n86_));
  OAI210     u69(.A0(men_men_n86_), .A1(i_1_), .B0(men_men_n62_), .Y(men_men_n87_));
  OAI210     u70(.A0(men_men_n87_), .A1(men_men_n33_), .B0(i_6_), .Y(men_men_n88_));
  AOI210     u71(.A0(men_men_n32_), .A1(men_men_n26_), .B0(men_men_n29_), .Y(men_men_n89_));
  OR2        u72(.A(men_men_n89_), .B(men_men_n76_), .Y(men_men_n90_));
  NA3        u73(.A(men_men_n86_), .B(men_men_n76_), .C(i_2_), .Y(men_men_n91_));
  NA3        u74(.A(men_men_n23_), .B(i_1_), .C(men_men_n26_), .Y(men_men_n92_));
  NA4        u75(.A(men_men_n92_), .B(men_men_n91_), .C(men_men_n90_), .D(men_men_n88_), .Y(men04));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
endmodule