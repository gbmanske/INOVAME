// Benchmark "top" written by ABC on Fri Jun 21 17:49:24 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n130_, new_new_n131_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n328_, new_new_n329_,
    new_new_n330_, new_new_n331_, new_new_n332_, new_new_n333_,
    new_new_n334_, new_new_n335_, new_new_n336_, new_new_n337_,
    new_new_n338_, new_new_n339_, new_new_n340_, new_new_n341_,
    new_new_n342_, new_new_n343_, new_new_n344_, new_new_n345_,
    new_new_n346_, new_new_n347_, new_new_n348_, new_new_n349_,
    new_new_n350_, new_new_n351_, new_new_n352_, new_new_n353_,
    new_new_n354_, new_new_n355_, new_new_n356_, new_new_n357_,
    new_new_n358_, new_new_n359_, new_new_n360_, new_new_n361_,
    new_new_n362_, new_new_n363_, new_new_n364_, new_new_n365_,
    new_new_n366_, new_new_n367_, new_new_n368_, new_new_n369_,
    new_new_n370_, new_new_n371_, new_new_n372_, new_new_n373_,
    new_new_n374_, new_new_n375_, new_new_n376_, new_new_n377_,
    new_new_n378_, new_new_n379_, new_new_n380_, new_new_n381_,
    new_new_n382_, new_new_n383_, new_new_n384_, new_new_n385_,
    new_new_n386_, new_new_n387_, new_new_n388_, new_new_n389_,
    new_new_n390_, new_new_n391_, new_new_n392_, new_new_n393_,
    new_new_n394_, new_new_n395_, new_new_n396_, new_new_n397_,
    new_new_n398_, new_new_n399_, new_new_n400_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n406_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n448_, new_new_n449_, new_new_n450_,
    new_new_n451_, new_new_n452_, new_new_n453_, new_new_n454_,
    new_new_n455_, new_new_n456_, new_new_n457_, new_new_n458_,
    new_new_n459_, new_new_n460_, new_new_n461_, new_new_n462_,
    new_new_n463_, new_new_n464_, new_new_n465_, new_new_n466_,
    new_new_n467_, new_new_n468_, new_new_n469_, new_new_n470_,
    new_new_n471_, new_new_n472_, new_new_n473_, new_new_n474_,
    new_new_n475_, new_new_n476_, new_new_n477_, new_new_n478_,
    new_new_n479_, new_new_n480_, new_new_n481_, new_new_n482_,
    new_new_n483_, new_new_n484_, new_new_n485_, new_new_n486_,
    new_new_n487_, new_new_n489_, new_new_n490_, new_new_n491_,
    new_new_n492_, new_new_n493_, new_new_n494_, new_new_n495_,
    new_new_n496_, new_new_n497_, new_new_n498_, new_new_n499_,
    new_new_n500_, new_new_n501_, new_new_n502_, new_new_n503_,
    new_new_n504_, new_new_n505_, new_new_n506_, new_new_n507_,
    new_new_n508_, new_new_n509_, new_new_n510_, new_new_n511_,
    new_new_n512_, new_new_n513_, new_new_n514_, new_new_n515_,
    new_new_n516_, new_new_n517_, new_new_n518_, new_new_n519_,
    new_new_n520_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n621_, new_new_n622_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(ori1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  NO2        g027(.A(i_5_), .B(new_new_n45_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA2        g031(.A(new_new_n50_), .B(new_new_n44_), .Y(new_new_n54_));
  NA3        g032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n55_));
  NO2        g033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  OAI210     g035(.A0(new_new_n57_), .A1(new_new_n56_), .B0(new_new_n55_), .Y(new_new_n58_));
  NA2        g036(.A(new_new_n58_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g038(.A(i_1_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA3        g040(.A(new_new_n62_), .B(new_new_n60_), .C(new_new_n31_), .Y(new_new_n63_));
  NA2        g041(.A(i_1_), .B(i_10_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NAi31      g043(.An(new_new_n65_), .B(new_new_n63_), .C(new_new_n59_), .Y(new_new_n66_));
  NA2        g044(.A(new_new_n49_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n75_), .Y(new_new_n76_));
  OAI210     g054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  INV        g056(.A(i_8_), .Y(new_new_n79_));
  NO2        g057(.A(new_new_n79_), .B(new_new_n56_), .Y(new_new_n80_));
  NO2        g058(.A(i_3_), .B(i_9_), .Y(new_new_n81_));
  NO2        g059(.A(i_3_), .B(i_7_), .Y(new_new_n82_));
  NO2        g060(.A(new_new_n81_), .B(new_new_n61_), .Y(new_new_n83_));
  INV        g061(.A(i_6_), .Y(new_new_n84_));
  NO2        g062(.A(i_2_), .B(i_7_), .Y(new_new_n85_));
  INV        g063(.A(new_new_n85_), .Y(new_new_n86_));
  OAI210     g064(.A0(new_new_n83_), .A1(new_new_n80_), .B0(new_new_n86_), .Y(new_new_n87_));
  NAi21      g065(.An(i_6_), .B(i_10_), .Y(new_new_n88_));
  NA2        g066(.A(i_6_), .B(i_9_), .Y(new_new_n89_));
  AOI210     g067(.A0(new_new_n89_), .A1(new_new_n88_), .B0(new_new_n61_), .Y(new_new_n90_));
  NA2        g068(.A(i_2_), .B(i_6_), .Y(new_new_n91_));
  NO3        g069(.A(new_new_n91_), .B(new_new_n48_), .C(new_new_n25_), .Y(new_new_n92_));
  NO2        g070(.A(new_new_n92_), .B(new_new_n90_), .Y(new_new_n93_));
  AOI210     g071(.A0(new_new_n93_), .A1(new_new_n87_), .B0(new_new_n78_), .Y(new_new_n94_));
  AN3        g072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n95_));
  NA2        g073(.A(new_new_n95_), .B(new_new_n32_), .Y(new_new_n96_));
  INV        g074(.A(i_7_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n45_), .B(new_new_n97_), .Y(new_new_n98_));
  NO2        g076(.A(i_0_), .B(i_5_), .Y(new_new_n99_));
  NO2        g077(.A(new_new_n99_), .B(new_new_n84_), .Y(new_new_n100_));
  NA2        g078(.A(i_12_), .B(i_3_), .Y(new_new_n101_));
  INV        g079(.A(new_new_n101_), .Y(new_new_n102_));
  NA3        g080(.A(new_new_n102_), .B(new_new_n100_), .C(new_new_n98_), .Y(new_new_n103_));
  NAi21      g081(.An(i_7_), .B(i_11_), .Y(new_new_n104_));
  NO3        g082(.A(new_new_n104_), .B(new_new_n88_), .C(new_new_n51_), .Y(new_new_n105_));
  AN2        g083(.A(i_2_), .B(i_10_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(i_7_), .Y(new_new_n107_));
  OR2        g085(.A(new_new_n78_), .B(new_new_n56_), .Y(new_new_n108_));
  NA2        g086(.A(i_12_), .B(i_7_), .Y(new_new_n109_));
  NO2        g087(.A(new_new_n61_), .B(new_new_n26_), .Y(new_new_n110_));
  NA2        g088(.A(i_11_), .B(i_12_), .Y(new_new_n111_));
  NAi41      g089(.An(new_new_n105_), .B(new_new_n111_), .C(new_new_n103_), .D(new_new_n96_), .Y(new_new_n112_));
  NOi21      g090(.An(i_1_), .B(i_5_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n113_), .B(i_11_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n115_));
  NA2        g093(.A(i_7_), .B(new_new_n25_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(new_new_n115_), .Y(new_new_n117_));
  NO2        g095(.A(new_new_n117_), .B(new_new_n45_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n89_), .B(new_new_n88_), .Y(new_new_n119_));
  NAi21      g097(.An(i_3_), .B(i_8_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(new_new_n60_), .Y(new_new_n121_));
  NOi31      g099(.An(new_new_n121_), .B(new_new_n119_), .C(new_new_n118_), .Y(new_new_n122_));
  NO2        g100(.A(i_1_), .B(new_new_n84_), .Y(new_new_n123_));
  NO2        g101(.A(i_6_), .B(i_5_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(i_3_), .Y(new_new_n125_));
  AO210      g103(.A0(new_new_n125_), .A1(new_new_n46_), .B0(new_new_n123_), .Y(new_new_n126_));
  OAI220     g104(.A0(new_new_n126_), .A1(new_new_n104_), .B0(new_new_n122_), .B1(new_new_n114_), .Y(new_new_n127_));
  NO3        g105(.A(new_new_n127_), .B(new_new_n112_), .C(new_new_n94_), .Y(new_new_n128_));
  NA3        g106(.A(new_new_n128_), .B(new_new_n77_), .C(new_new_n54_), .Y(ori2));
  NO2        g107(.A(new_new_n61_), .B(new_new_n37_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n621_), .B(new_new_n130_), .Y(new_new_n131_));
  NA4        g109(.A(new_new_n131_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(ori0));
  NO2        g110(.A(i_12_), .B(i_13_), .Y(new_new_n133_));
  NAi21      g111(.An(i_5_), .B(i_11_), .Y(new_new_n134_));
  NO2        g112(.A(i_0_), .B(i_1_), .Y(new_new_n135_));
  NA2        g113(.A(i_2_), .B(i_3_), .Y(new_new_n136_));
  NA2        g114(.A(i_1_), .B(i_5_), .Y(new_new_n137_));
  NOi21      g115(.An(i_4_), .B(i_10_), .Y(new_new_n138_));
  NA2        g116(.A(new_new_n138_), .B(new_new_n40_), .Y(new_new_n139_));
  NOi21      g117(.An(i_4_), .B(i_9_), .Y(new_new_n140_));
  NOi21      g118(.An(i_11_), .B(i_13_), .Y(new_new_n141_));
  NA2        g119(.A(new_new_n141_), .B(new_new_n140_), .Y(new_new_n142_));
  NAi21      g120(.An(i_12_), .B(i_11_), .Y(new_new_n143_));
  NO2        g121(.A(new_new_n71_), .B(new_new_n61_), .Y(new_new_n144_));
  NO2        g122(.A(new_new_n71_), .B(i_5_), .Y(new_new_n145_));
  NO2        g123(.A(i_2_), .B(i_1_), .Y(new_new_n146_));
  NAi21      g124(.An(i_4_), .B(i_12_), .Y(new_new_n147_));
  INV        g125(.A(i_8_), .Y(new_new_n148_));
  NO3        g126(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n149_));
  NO2        g127(.A(i_3_), .B(i_8_), .Y(new_new_n150_));
  NO3        g128(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n151_));
  NO2        g129(.A(new_new_n99_), .B(new_new_n56_), .Y(new_new_n152_));
  NO2        g130(.A(i_13_), .B(i_9_), .Y(new_new_n153_));
  NAi21      g131(.An(i_12_), .B(i_3_), .Y(new_new_n154_));
  NO2        g132(.A(new_new_n43_), .B(i_5_), .Y(new_new_n155_));
  NA3        g133(.A(i_13_), .B(new_new_n148_), .C(i_10_), .Y(new_new_n156_));
  NA2        g134(.A(i_0_), .B(i_5_), .Y(new_new_n157_));
  NAi31      g135(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n158_));
  NO2        g136(.A(new_new_n36_), .B(i_13_), .Y(new_new_n159_));
  NO2        g137(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n45_), .B(new_new_n61_), .Y(new_new_n161_));
  INV        g139(.A(i_13_), .Y(new_new_n162_));
  NO2        g140(.A(i_12_), .B(new_new_n162_), .Y(new_new_n163_));
  NO2        g141(.A(i_12_), .B(new_new_n37_), .Y(new_new_n164_));
  INV        g142(.A(i_12_), .Y(new_new_n165_));
  NO3        g143(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n166_));
  NA2        g144(.A(i_2_), .B(i_1_), .Y(new_new_n167_));
  NO3        g145(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n168_));
  NAi21      g146(.An(i_4_), .B(i_3_), .Y(new_new_n169_));
  NO2        g147(.A(i_0_), .B(i_6_), .Y(new_new_n170_));
  NOi41      g148(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n171_));
  NO2        g149(.A(i_11_), .B(new_new_n162_), .Y(new_new_n172_));
  NOi21      g150(.An(i_1_), .B(i_6_), .Y(new_new_n173_));
  NAi21      g151(.An(i_3_), .B(i_7_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n165_), .B(i_9_), .Y(new_new_n175_));
  OR4        g153(.A(new_new_n175_), .B(new_new_n174_), .C(new_new_n173_), .D(new_new_n145_), .Y(new_new_n176_));
  NA2        g154(.A(new_new_n71_), .B(i_5_), .Y(new_new_n177_));
  NA2        g155(.A(i_3_), .B(i_9_), .Y(new_new_n178_));
  NAi21      g156(.An(i_7_), .B(i_10_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n179_), .B(new_new_n178_), .Y(new_new_n180_));
  NA3        g158(.A(new_new_n180_), .B(new_new_n177_), .C(new_new_n62_), .Y(new_new_n181_));
  NA2        g159(.A(new_new_n181_), .B(new_new_n176_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n182_), .B(new_new_n172_), .Y(new_new_n183_));
  NA2        g161(.A(i_12_), .B(i_6_), .Y(new_new_n184_));
  OR2        g162(.A(i_13_), .B(i_9_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n169_), .B(i_2_), .Y(new_new_n186_));
  NA2        g164(.A(new_new_n172_), .B(i_9_), .Y(new_new_n187_));
  NO3        g165(.A(i_11_), .B(new_new_n162_), .C(new_new_n25_), .Y(new_new_n188_));
  NO3        g166(.A(i_12_), .B(new_new_n162_), .C(new_new_n37_), .Y(new_new_n189_));
  AN2        g167(.A(i_3_), .B(i_10_), .Y(new_new_n190_));
  NO2        g168(.A(i_5_), .B(new_new_n37_), .Y(new_new_n191_));
  NO3        g169(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n192_));
  NO2        g170(.A(i_2_), .B(i_3_), .Y(new_new_n193_));
  OR2        g171(.A(i_0_), .B(i_5_), .Y(new_new_n194_));
  NO2        g172(.A(i_12_), .B(i_10_), .Y(new_new_n195_));
  NOi21      g173(.An(i_5_), .B(i_0_), .Y(new_new_n196_));
  NO2        g174(.A(i_1_), .B(i_7_), .Y(new_new_n197_));
  NOi21      g175(.An(new_new_n137_), .B(new_new_n100_), .Y(new_new_n198_));
  NO2        g176(.A(new_new_n198_), .B(new_new_n116_), .Y(new_new_n199_));
  NA2        g177(.A(new_new_n199_), .B(i_3_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n148_), .B(i_9_), .Y(new_new_n201_));
  NA2        g179(.A(new_new_n201_), .B(new_new_n152_), .Y(new_new_n202_));
  NO2        g180(.A(new_new_n202_), .B(new_new_n45_), .Y(new_new_n203_));
  INV        g181(.A(new_new_n203_), .Y(new_new_n204_));
  AOI210     g182(.A0(new_new_n204_), .A1(new_new_n200_), .B0(new_new_n139_), .Y(new_new_n205_));
  INV        g183(.A(new_new_n205_), .Y(new_new_n206_));
  NOi32      g184(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n207_));
  INV        g185(.A(new_new_n207_), .Y(new_new_n208_));
  NOi32      g186(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n209_));
  NAi21      g187(.An(i_6_), .B(i_1_), .Y(new_new_n210_));
  NA3        g188(.A(new_new_n210_), .B(new_new_n209_), .C(new_new_n45_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n211_), .B(i_0_), .Y(new_new_n212_));
  NO2        g190(.A(i_1_), .B(new_new_n97_), .Y(new_new_n213_));
  NAi21      g191(.An(i_3_), .B(i_4_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n214_), .B(i_9_), .Y(new_new_n215_));
  AN2        g193(.A(i_6_), .B(i_7_), .Y(new_new_n216_));
  OAI210     g194(.A0(new_new_n216_), .A1(new_new_n213_), .B0(new_new_n215_), .Y(new_new_n217_));
  NA2        g195(.A(i_2_), .B(i_7_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n214_), .B(i_10_), .Y(new_new_n219_));
  NA3        g197(.A(new_new_n219_), .B(new_new_n218_), .C(new_new_n170_), .Y(new_new_n220_));
  AOI210     g198(.A0(new_new_n220_), .A1(new_new_n217_), .B0(new_new_n145_), .Y(new_new_n221_));
  AOI210     g199(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n222_));
  OAI210     g200(.A0(new_new_n222_), .A1(new_new_n146_), .B0(new_new_n219_), .Y(new_new_n223_));
  AOI220     g201(.A0(new_new_n219_), .A1(new_new_n197_), .B0(new_new_n166_), .B1(new_new_n146_), .Y(new_new_n224_));
  AOI210     g202(.A0(new_new_n224_), .A1(new_new_n223_), .B0(i_5_), .Y(new_new_n225_));
  NO3        g203(.A(new_new_n225_), .B(new_new_n221_), .C(new_new_n212_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n226_), .B(new_new_n208_), .Y(new_new_n227_));
  AN2        g205(.A(i_12_), .B(i_5_), .Y(new_new_n228_));
  INV        g206(.A(new_new_n228_), .Y(new_new_n229_));
  NO2        g207(.A(i_11_), .B(i_6_), .Y(new_new_n230_));
  NO2        g208(.A(i_5_), .B(i_10_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n232_));
  NO3        g210(.A(new_new_n84_), .B(new_new_n47_), .C(i_9_), .Y(new_new_n233_));
  NO2        g211(.A(i_11_), .B(i_12_), .Y(new_new_n234_));
  NAi21      g212(.An(i_13_), .B(i_0_), .Y(new_new_n235_));
  NO3        g213(.A(i_1_), .B(i_12_), .C(new_new_n84_), .Y(new_new_n236_));
  NO2        g214(.A(i_0_), .B(i_11_), .Y(new_new_n237_));
  AN2        g215(.A(i_1_), .B(i_6_), .Y(new_new_n238_));
  NOi21      g216(.An(i_2_), .B(i_12_), .Y(new_new_n239_));
  NAi21      g217(.An(i_9_), .B(i_4_), .Y(new_new_n240_));
  OR2        g218(.A(i_13_), .B(i_10_), .Y(new_new_n241_));
  NO3        g219(.A(new_new_n241_), .B(new_new_n111_), .C(new_new_n240_), .Y(new_new_n242_));
  NO2        g220(.A(new_new_n142_), .B(new_new_n115_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n97_), .B(new_new_n25_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n189_), .B(new_new_n244_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n245_), .B(new_new_n198_), .Y(new_new_n246_));
  INV        g224(.A(new_new_n246_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n247_), .B(new_new_n26_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n148_), .B(i_10_), .Y(new_new_n249_));
  NA3        g227(.A(new_new_n177_), .B(new_new_n62_), .C(i_2_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n250_), .B(new_new_n249_), .Y(new_new_n251_));
  INV        g229(.A(new_new_n251_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n252_), .B(new_new_n187_), .Y(new_new_n253_));
  NO3        g231(.A(new_new_n253_), .B(new_new_n248_), .C(new_new_n227_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n71_), .B(i_13_), .Y(new_new_n255_));
  NO2        g233(.A(i_10_), .B(i_9_), .Y(new_new_n256_));
  NAi21      g234(.An(i_12_), .B(i_8_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n257_), .B(i_3_), .Y(new_new_n258_));
  NA2        g236(.A(i_8_), .B(i_9_), .Y(new_new_n259_));
  NA2        g237(.A(new_new_n189_), .B(new_new_n152_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n260_), .B(new_new_n259_), .Y(new_new_n261_));
  NA2        g239(.A(new_new_n172_), .B(new_new_n191_), .Y(new_new_n262_));
  NO3        g240(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n263_));
  INV        g241(.A(new_new_n263_), .Y(new_new_n264_));
  NA3        g242(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n265_));
  NA4        g243(.A(new_new_n134_), .B(new_new_n110_), .C(new_new_n78_), .D(new_new_n23_), .Y(new_new_n266_));
  OAI220     g244(.A0(new_new_n266_), .A1(new_new_n265_), .B0(new_new_n264_), .B1(new_new_n262_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n267_), .B(new_new_n261_), .Y(new_new_n268_));
  NA2        g246(.A(new_new_n95_), .B(i_13_), .Y(new_new_n269_));
  NO3        g247(.A(i_4_), .B(new_new_n47_), .C(i_8_), .Y(new_new_n270_));
  NO2        g248(.A(i_6_), .B(i_7_), .Y(new_new_n271_));
  NO2        g249(.A(i_11_), .B(i_1_), .Y(new_new_n272_));
  NOi21      g250(.An(i_2_), .B(i_7_), .Y(new_new_n273_));
  NO2        g251(.A(i_6_), .B(i_10_), .Y(new_new_n274_));
  NA3        g252(.A(new_new_n171_), .B(new_new_n141_), .C(new_new_n124_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n45_), .B(new_new_n43_), .Y(new_new_n276_));
  NA2        g254(.A(new_new_n263_), .B(new_new_n231_), .Y(new_new_n277_));
  NAi21      g255(.An(new_new_n156_), .B(new_new_n234_), .Y(new_new_n278_));
  NA2        g256(.A(new_new_n197_), .B(new_new_n157_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n279_), .B(new_new_n278_), .Y(new_new_n280_));
  NA2        g258(.A(new_new_n27_), .B(i_10_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n192_), .B(new_new_n166_), .Y(new_new_n282_));
  OAI220     g260(.A0(new_new_n282_), .A1(new_new_n250_), .B0(new_new_n281_), .B1(new_new_n269_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n283_), .B(new_new_n280_), .Y(new_new_n284_));
  NA3        g262(.A(new_new_n284_), .B(new_new_n275_), .C(new_new_n268_), .Y(new_new_n285_));
  NA2        g263(.A(new_new_n228_), .B(new_new_n162_), .Y(new_new_n286_));
  NA2        g264(.A(new_new_n216_), .B(new_new_n209_), .Y(new_new_n287_));
  OR2        g265(.A(new_new_n286_), .B(new_new_n287_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n36_), .B(i_8_), .Y(new_new_n289_));
  AOI210     g267(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n242_), .Y(new_new_n290_));
  NA2        g268(.A(new_new_n290_), .B(new_new_n288_), .Y(new_new_n291_));
  INV        g269(.A(new_new_n291_), .Y(new_new_n292_));
  NA2        g270(.A(new_new_n177_), .B(new_new_n62_), .Y(new_new_n293_));
  OAI210     g271(.A0(i_8_), .A1(new_new_n293_), .B0(new_new_n126_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n294_), .B(new_new_n243_), .Y(new_new_n295_));
  NA2        g273(.A(new_new_n295_), .B(new_new_n292_), .Y(new_new_n296_));
  NO2        g274(.A(i_12_), .B(new_new_n148_), .Y(new_new_n297_));
  NA2        g275(.A(new_new_n43_), .B(i_10_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n298_), .B(i_6_), .Y(new_new_n299_));
  NO2        g277(.A(i_0_), .B(i_5_), .Y(new_new_n300_));
  NA3        g278(.A(new_new_n157_), .B(new_new_n69_), .C(new_new_n43_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n189_), .B(new_new_n82_), .Y(new_new_n302_));
  NO2        g280(.A(new_new_n301_), .B(new_new_n302_), .Y(new_new_n303_));
  NA2        g281(.A(new_new_n161_), .B(new_new_n160_), .Y(new_new_n304_));
  NA2        g282(.A(new_new_n256_), .B(new_new_n159_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n304_), .B(new_new_n305_), .Y(new_new_n306_));
  AOI210     g284(.A0(new_new_n210_), .A1(new_new_n45_), .B0(new_new_n213_), .Y(new_new_n307_));
  NA2        g285(.A(i_0_), .B(new_new_n47_), .Y(new_new_n308_));
  NA3        g286(.A(new_new_n297_), .B(new_new_n188_), .C(new_new_n308_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n307_), .B(new_new_n309_), .Y(new_new_n310_));
  NO3        g288(.A(new_new_n310_), .B(new_new_n306_), .C(new_new_n303_), .Y(new_new_n311_));
  NOi21      g289(.An(i_10_), .B(i_6_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n84_), .B(new_new_n25_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n109_), .B(new_new_n23_), .Y(new_new_n314_));
  INV        g292(.A(new_new_n193_), .Y(new_new_n315_));
  NO2        g293(.A(i_12_), .B(new_new_n84_), .Y(new_new_n316_));
  NA3        g294(.A(new_new_n316_), .B(new_new_n188_), .C(new_new_n308_), .Y(new_new_n317_));
  NA3        g295(.A(new_new_n230_), .B(new_new_n189_), .C(new_new_n157_), .Y(new_new_n318_));
  AOI210     g296(.A0(new_new_n318_), .A1(new_new_n317_), .B0(new_new_n315_), .Y(new_new_n319_));
  OR2        g297(.A(i_2_), .B(i_5_), .Y(new_new_n320_));
  OR2        g298(.A(new_new_n320_), .B(new_new_n238_), .Y(new_new_n321_));
  NA2        g299(.A(new_new_n218_), .B(new_new_n170_), .Y(new_new_n322_));
  AOI210     g300(.A0(new_new_n322_), .A1(new_new_n321_), .B0(new_new_n278_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n323_), .B(new_new_n319_), .Y(new_new_n324_));
  NA2        g302(.A(new_new_n324_), .B(new_new_n311_), .Y(new_new_n325_));
  NO3        g303(.A(new_new_n325_), .B(new_new_n296_), .C(new_new_n285_), .Y(new_new_n326_));
  NA4        g304(.A(new_new_n326_), .B(new_new_n254_), .C(new_new_n206_), .D(new_new_n183_), .Y(ori7));
  NO2        g305(.A(new_new_n91_), .B(new_new_n52_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n274_), .B(new_new_n82_), .Y(new_new_n329_));
  NA2        g307(.A(i_11_), .B(new_new_n148_), .Y(new_new_n330_));
  INV        g308(.A(new_new_n133_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n331_), .B(new_new_n329_), .Y(new_new_n332_));
  NA3        g310(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n165_), .B(i_4_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(i_8_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n101_), .B(new_new_n333_), .Y(new_new_n336_));
  NA2        g314(.A(i_2_), .B(new_new_n84_), .Y(new_new_n337_));
  OAI210     g315(.A0(new_new_n85_), .A1(new_new_n150_), .B0(new_new_n151_), .Y(new_new_n338_));
  NO2        g316(.A(i_7_), .B(new_new_n37_), .Y(new_new_n339_));
  NA2        g317(.A(i_4_), .B(i_8_), .Y(new_new_n340_));
  AOI210     g318(.A0(new_new_n340_), .A1(new_new_n190_), .B0(new_new_n339_), .Y(new_new_n341_));
  NO2        g319(.A(new_new_n341_), .B(new_new_n337_), .Y(new_new_n342_));
  NO4        g320(.A(new_new_n342_), .B(new_new_n336_), .C(new_new_n332_), .D(new_new_n328_), .Y(new_new_n343_));
  AOI210     g321(.A0(new_new_n120_), .A1(new_new_n60_), .B0(i_10_), .Y(new_new_n344_));
  AOI210     g322(.A0(new_new_n344_), .A1(new_new_n165_), .B0(new_new_n138_), .Y(new_new_n345_));
  OR2        g323(.A(i_6_), .B(i_10_), .Y(new_new_n346_));
  OR3        g324(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n347_));
  INV        g325(.A(new_new_n149_), .Y(new_new_n348_));
  OR2        g326(.A(new_new_n345_), .B(new_new_n185_), .Y(new_new_n349_));
  AOI210     g327(.A0(new_new_n349_), .A1(new_new_n343_), .B0(new_new_n61_), .Y(new_new_n350_));
  NOi21      g328(.An(i_11_), .B(i_7_), .Y(new_new_n351_));
  AO210      g329(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n352_));
  NO2        g330(.A(new_new_n352_), .B(new_new_n351_), .Y(new_new_n353_));
  NA2        g331(.A(new_new_n353_), .B(new_new_n153_), .Y(new_new_n354_));
  NA3        g332(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n354_), .B(new_new_n61_), .Y(new_new_n356_));
  NO3        g334(.A(new_new_n179_), .B(new_new_n154_), .C(new_new_n330_), .Y(new_new_n357_));
  OAI210     g335(.A0(new_new_n357_), .A1(new_new_n163_), .B0(new_new_n61_), .Y(new_new_n358_));
  NA2        g336(.A(new_new_n239_), .B(new_new_n31_), .Y(new_new_n359_));
  OR2        g337(.A(new_new_n154_), .B(new_new_n104_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n360_), .B(new_new_n359_), .Y(new_new_n361_));
  NO2        g339(.A(i_1_), .B(i_4_), .Y(new_new_n362_));
  NA2        g340(.A(new_new_n362_), .B(new_new_n361_), .Y(new_new_n363_));
  NO2        g341(.A(i_1_), .B(i_12_), .Y(new_new_n364_));
  NA3        g342(.A(new_new_n364_), .B(new_new_n106_), .C(new_new_n24_), .Y(new_new_n365_));
  BUFFER     g343(.A(new_new_n365_), .Y(new_new_n366_));
  NA3        g344(.A(new_new_n366_), .B(new_new_n363_), .C(new_new_n358_), .Y(new_new_n367_));
  OAI210     g345(.A0(new_new_n367_), .A1(new_new_n356_), .B0(i_6_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n355_), .B(new_new_n104_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n369_), .B(new_new_n316_), .Y(new_new_n370_));
  NO2        g348(.A(i_6_), .B(i_11_), .Y(new_new_n371_));
  INV        g349(.A(new_new_n370_), .Y(new_new_n372_));
  NO3        g350(.A(new_new_n346_), .B(i_8_), .C(new_new_n23_), .Y(new_new_n373_));
  AOI210     g351(.A0(i_1_), .A1(new_new_n180_), .B0(new_new_n373_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n374_), .B(new_new_n43_), .Y(new_new_n375_));
  INV        g353(.A(i_2_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n130_), .B(i_9_), .Y(new_new_n377_));
  NA3        g355(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n45_), .B(i_1_), .Y(new_new_n379_));
  NA3        g357(.A(new_new_n379_), .B(new_new_n184_), .C(new_new_n43_), .Y(new_new_n380_));
  OAI220     g358(.A0(new_new_n380_), .A1(new_new_n378_), .B0(new_new_n377_), .B1(new_new_n376_), .Y(new_new_n381_));
  AOI210     g359(.A0(new_new_n272_), .A1(new_new_n244_), .B0(new_new_n168_), .Y(new_new_n382_));
  NO2        g360(.A(new_new_n382_), .B(new_new_n337_), .Y(new_new_n383_));
  OR2        g361(.A(new_new_n383_), .B(new_new_n381_), .Y(new_new_n384_));
  NO3        g362(.A(new_new_n384_), .B(new_new_n375_), .C(new_new_n372_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n165_), .B(new_new_n97_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n386_), .B(new_new_n351_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n387_), .B(i_1_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n388_), .B(new_new_n347_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n240_), .B(new_new_n84_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n389_), .B(new_new_n45_), .Y(new_new_n391_));
  NA2        g369(.A(i_3_), .B(new_new_n148_), .Y(new_new_n392_));
  NO2        g370(.A(new_new_n392_), .B(new_new_n109_), .Y(new_new_n393_));
  AN2        g371(.A(new_new_n393_), .B(new_new_n299_), .Y(new_new_n394_));
  NO2        g372(.A(i_8_), .B(new_new_n43_), .Y(new_new_n395_));
  NA2        g373(.A(i_1_), .B(i_3_), .Y(new_new_n396_));
  NO2        g374(.A(new_new_n259_), .B(new_new_n91_), .Y(new_new_n397_));
  AOI210     g375(.A0(new_new_n395_), .A1(new_new_n312_), .B0(new_new_n397_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n396_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(new_new_n394_), .Y(new_new_n400_));
  NA4        g378(.A(new_new_n400_), .B(new_new_n391_), .C(new_new_n385_), .D(new_new_n368_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n402_));
  NO3        g380(.A(new_new_n273_), .B(new_new_n340_), .C(new_new_n84_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n403_), .B(new_new_n25_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n404_), .B(new_new_n402_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n405_), .B(i_1_), .Y(new_new_n406_));
  INV        g384(.A(i_1_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n214_), .B(i_2_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n406_), .B(i_13_), .Y(new_new_n409_));
  OR2        g387(.A(i_11_), .B(i_7_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n52_), .B(i_12_), .Y(new_new_n411_));
  INV        g389(.A(new_new_n411_), .Y(new_new_n412_));
  NO2        g390(.A(new_new_n273_), .B(new_new_n24_), .Y(new_new_n413_));
  AOI220     g391(.A0(new_new_n413_), .A1(new_new_n390_), .B0(new_new_n171_), .B1(new_new_n123_), .Y(new_new_n414_));
  OAI220     g392(.A0(new_new_n414_), .A1(new_new_n41_), .B0(new_new_n412_), .B1(new_new_n91_), .Y(new_new_n415_));
  INV        g393(.A(new_new_n415_), .Y(new_new_n416_));
  AOI210     g394(.A0(new_new_n257_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n417_));
  NOi31      g395(.An(new_new_n417_), .B(new_new_n329_), .C(new_new_n43_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n119_), .B(i_13_), .Y(new_new_n419_));
  NO2        g397(.A(new_new_n378_), .B(new_new_n109_), .Y(new_new_n420_));
  INV        g398(.A(new_new_n420_), .Y(new_new_n421_));
  OAI220     g399(.A0(new_new_n421_), .A1(new_new_n69_), .B0(new_new_n419_), .B1(new_new_n407_), .Y(new_new_n422_));
  NO3        g400(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n97_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n26_), .B(new_new_n148_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n424_), .B(i_7_), .Y(new_new_n425_));
  NO3        g403(.A(new_new_n273_), .B(new_new_n165_), .C(new_new_n84_), .Y(new_new_n426_));
  AOI210     g404(.A0(new_new_n426_), .A1(new_new_n425_), .B0(new_new_n423_), .Y(new_new_n427_));
  AOI210     g405(.A0(new_new_n230_), .A1(new_new_n379_), .B0(new_new_n90_), .Y(new_new_n428_));
  OAI220     g406(.A0(new_new_n428_), .A1(new_new_n335_), .B0(new_new_n427_), .B1(new_new_n348_), .Y(new_new_n429_));
  NO3        g407(.A(new_new_n429_), .B(new_new_n422_), .C(new_new_n418_), .Y(new_new_n430_));
  OR2        g408(.A(i_11_), .B(i_6_), .Y(new_new_n431_));
  NA3        g409(.A(new_new_n239_), .B(new_new_n339_), .C(i_6_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n371_), .B(i_13_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n98_), .B(new_new_n424_), .Y(new_new_n434_));
  NAi21      g412(.An(i_11_), .B(i_12_), .Y(new_new_n435_));
  NOi41      g413(.An(new_new_n107_), .B(new_new_n435_), .C(i_13_), .D(new_new_n84_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n316_), .B(new_new_n340_), .Y(new_new_n437_));
  AOI220     g415(.A0(new_new_n437_), .A1(new_new_n192_), .B0(new_new_n436_), .B1(new_new_n434_), .Y(new_new_n438_));
  NA3        g416(.A(new_new_n438_), .B(new_new_n433_), .C(new_new_n432_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n439_), .B(new_new_n61_), .Y(new_new_n440_));
  NO2        g418(.A(i_2_), .B(i_12_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n213_), .B(new_new_n441_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n215_), .B(new_new_n213_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n443_), .B(new_new_n442_), .Y(new_new_n444_));
  NA3        g422(.A(new_new_n444_), .B(new_new_n44_), .C(new_new_n162_), .Y(new_new_n445_));
  NA4        g423(.A(new_new_n445_), .B(new_new_n440_), .C(new_new_n430_), .D(new_new_n416_), .Y(new_new_n446_));
  OR4        g424(.A(new_new_n446_), .B(new_new_n409_), .C(new_new_n401_), .D(new_new_n350_), .Y(ori5));
  NA2        g425(.A(new_new_n387_), .B(new_new_n186_), .Y(new_new_n448_));
  AN2        g426(.A(new_new_n24_), .B(i_10_), .Y(new_new_n449_));
  NA3        g427(.A(new_new_n449_), .B(new_new_n441_), .C(new_new_n104_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n335_), .B(i_11_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n85_), .B(new_new_n451_), .Y(new_new_n452_));
  NA3        g430(.A(new_new_n452_), .B(new_new_n450_), .C(new_new_n448_), .Y(new_new_n453_));
  NO3        g431(.A(i_11_), .B(new_new_n165_), .C(i_13_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n455_));
  INV        g433(.A(new_new_n256_), .Y(new_new_n456_));
  AOI220     g434(.A0(new_new_n193_), .A1(new_new_n314_), .B0(i_12_), .B1(new_new_n455_), .Y(new_new_n457_));
  INV        g435(.A(new_new_n457_), .Y(new_new_n458_));
  NO2        g436(.A(new_new_n458_), .B(new_new_n453_), .Y(new_new_n459_));
  INV        g437(.A(new_new_n141_), .Y(new_new_n460_));
  INV        g438(.A(new_new_n171_), .Y(new_new_n461_));
  OAI210     g439(.A0(new_new_n408_), .A1(new_new_n258_), .B0(new_new_n107_), .Y(new_new_n462_));
  AOI210     g440(.A0(new_new_n462_), .A1(new_new_n461_), .B0(new_new_n460_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n259_), .B(new_new_n26_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n464_), .B(new_new_n244_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n465_), .B(i_2_), .Y(new_new_n466_));
  INV        g444(.A(new_new_n466_), .Y(new_new_n467_));
  AOI210     g445(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n241_), .Y(new_new_n468_));
  AOI210     g446(.A0(new_new_n468_), .A1(new_new_n467_), .B0(new_new_n463_), .Y(new_new_n469_));
  NO2        g447(.A(new_new_n147_), .B(new_new_n117_), .Y(new_new_n470_));
  OAI210     g448(.A0(new_new_n470_), .A1(new_new_n455_), .B0(i_2_), .Y(new_new_n471_));
  INV        g449(.A(new_new_n142_), .Y(new_new_n472_));
  NO3        g450(.A(new_new_n352_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n473_));
  AOI210     g451(.A0(new_new_n472_), .A1(new_new_n85_), .B0(new_new_n473_), .Y(new_new_n474_));
  AOI210     g452(.A0(new_new_n474_), .A1(new_new_n471_), .B0(new_new_n148_), .Y(new_new_n475_));
  OA210      g453(.A0(new_new_n353_), .A1(new_new_n118_), .B0(i_13_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n149_), .B(new_new_n150_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n477_), .B(new_new_n218_), .Y(new_new_n478_));
  AOI210     g456(.A0(new_new_n154_), .A1(new_new_n136_), .B0(new_new_n289_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n479_), .B(new_new_n244_), .Y(new_new_n480_));
  NA3        g458(.A(i_2_), .B(new_new_n190_), .C(new_new_n116_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n481_), .B(new_new_n480_), .Y(new_new_n482_));
  NO4        g460(.A(new_new_n482_), .B(new_new_n478_), .C(new_new_n476_), .D(new_new_n475_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n60_), .B(i_12_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n484_), .B(new_new_n118_), .Y(new_new_n485_));
  NO2        g463(.A(new_new_n485_), .B(new_new_n330_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n486_), .B(new_new_n36_), .Y(new_new_n487_));
  NA4        g465(.A(new_new_n487_), .B(new_new_n483_), .C(new_new_n469_), .D(new_new_n459_), .Y(ori6));
  NO2        g466(.A(new_new_n158_), .B(new_new_n276_), .Y(new_new_n489_));
  INV        g467(.A(new_new_n196_), .Y(new_new_n490_));
  OR2        g468(.A(new_new_n490_), .B(i_12_), .Y(new_new_n491_));
  INV        g469(.A(new_new_n195_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n73_), .B(new_new_n123_), .Y(new_new_n493_));
  INV        g471(.A(new_new_n116_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n494_), .B(new_new_n45_), .Y(new_new_n495_));
  AOI210     g473(.A0(new_new_n495_), .A1(new_new_n493_), .B0(new_new_n492_), .Y(new_new_n496_));
  NO2        g474(.A(new_new_n287_), .B(new_new_n145_), .Y(new_new_n497_));
  NO2        g475(.A(new_new_n32_), .B(i_11_), .Y(new_new_n498_));
  NAi32      g476(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n431_), .B(new_new_n499_), .Y(new_new_n500_));
  OR3        g478(.A(new_new_n500_), .B(new_new_n497_), .C(new_new_n496_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n410_), .B(i_2_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n47_), .B(new_new_n37_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(new_new_n238_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n504_), .B(new_new_n502_), .Y(new_new_n505_));
  BUFFER     g483(.A(new_new_n353_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n506_), .B(new_new_n135_), .Y(new_new_n507_));
  AO210      g485(.A0(new_new_n277_), .A1(new_new_n456_), .B0(new_new_n36_), .Y(new_new_n508_));
  NA3        g486(.A(new_new_n508_), .B(new_new_n507_), .C(new_new_n505_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n489_), .B(new_new_n425_), .Y(new_new_n510_));
  NA3        g488(.A(new_new_n218_), .B(new_new_n166_), .C(new_new_n135_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n233_), .B(new_new_n68_), .Y(new_new_n512_));
  NA4        g490(.A(new_new_n512_), .B(new_new_n511_), .C(new_new_n510_), .D(new_new_n338_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n258_), .B(new_new_n256_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n346_), .B(new_new_n98_), .Y(new_new_n515_));
  OAI210     g493(.A0(new_new_n515_), .A1(new_new_n108_), .B0(new_new_n237_), .Y(new_new_n516_));
  INV        g494(.A(new_new_n321_), .Y(new_new_n517_));
  NA3        g495(.A(new_new_n517_), .B(new_new_n195_), .C(i_7_), .Y(new_new_n518_));
  NA3        g496(.A(new_new_n518_), .B(new_new_n516_), .C(new_new_n514_), .Y(new_new_n519_));
  NO4        g497(.A(new_new_n519_), .B(new_new_n513_), .C(new_new_n509_), .D(new_new_n501_), .Y(new_new_n520_));
  NA3        g498(.A(new_new_n520_), .B(new_new_n491_), .C(new_new_n226_), .Y(ori3));
  NA2        g499(.A(i_12_), .B(i_10_), .Y(new_new_n522_));
  NO2        g500(.A(i_11_), .B(new_new_n165_), .Y(new_new_n523_));
  NA3        g501(.A(new_new_n511_), .B(new_new_n338_), .C(new_new_n217_), .Y(new_new_n524_));
  NA2        g502(.A(new_new_n524_), .B(new_new_n40_), .Y(new_new_n525_));
  NOi21      g503(.An(new_new_n95_), .B(new_new_n465_), .Y(new_new_n526_));
  NO3        g504(.A(new_new_n360_), .B(new_new_n259_), .C(new_new_n123_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n239_), .B(new_new_n44_), .Y(new_new_n528_));
  AN2        g506(.A(i_11_), .B(new_new_n53_), .Y(new_new_n529_));
  NO3        g507(.A(new_new_n529_), .B(new_new_n527_), .C(new_new_n526_), .Y(new_new_n530_));
  AOI210     g508(.A0(new_new_n530_), .A1(new_new_n525_), .B0(new_new_n47_), .Y(new_new_n531_));
  NO4        g509(.A(new_new_n222_), .B(new_new_n228_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n145_), .B(new_new_n312_), .Y(new_new_n533_));
  NOi21      g511(.An(new_new_n533_), .B(new_new_n532_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n534_), .B(new_new_n61_), .Y(new_new_n535_));
  NOi21      g513(.An(i_5_), .B(i_9_), .Y(new_new_n536_));
  NA2        g514(.A(new_new_n536_), .B(new_new_n255_), .Y(new_new_n537_));
  BUFFER     g515(.A(new_new_n184_), .Y(new_new_n538_));
  AOI210     g516(.A0(new_new_n538_), .A1(new_new_n272_), .B0(new_new_n403_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n539_), .B(new_new_n537_), .Y(new_new_n540_));
  NO3        g518(.A(new_new_n540_), .B(new_new_n535_), .C(new_new_n531_), .Y(new_new_n541_));
  NA2        g519(.A(new_new_n313_), .B(i_0_), .Y(new_new_n542_));
  NO3        g520(.A(new_new_n542_), .B(new_new_n229_), .C(new_new_n85_), .Y(new_new_n543_));
  NO4        g521(.A(new_new_n320_), .B(i_12_), .C(new_new_n241_), .D(new_new_n238_), .Y(new_new_n544_));
  AOI210     g522(.A0(new_new_n544_), .A1(i_11_), .B0(new_new_n543_), .Y(new_new_n545_));
  NA2        g523(.A(new_new_n454_), .B(new_new_n196_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n85_), .B(new_new_n56_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n547_), .B(new_new_n546_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n175_), .B(new_new_n137_), .Y(new_new_n549_));
  INV        g527(.A(new_new_n298_), .Y(new_new_n550_));
  NO4        g528(.A(new_new_n109_), .B(new_new_n56_), .C(new_new_n392_), .D(i_5_), .Y(new_new_n551_));
  AO220      g529(.A0(new_new_n551_), .A1(new_new_n550_), .B0(new_new_n549_), .B1(i_6_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n552_), .B(new_new_n548_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n553_), .B(new_new_n545_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n555_));
  NA2        g533(.A(i_11_), .B(i_9_), .Y(new_new_n556_));
  NO3        g534(.A(i_12_), .B(new_new_n556_), .C(new_new_n337_), .Y(new_new_n557_));
  AN2        g535(.A(new_new_n557_), .B(new_new_n555_), .Y(new_new_n558_));
  NA2        g536(.A(new_new_n232_), .B(new_new_n144_), .Y(new_new_n559_));
  INV        g537(.A(new_new_n559_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n556_), .B(new_new_n71_), .Y(new_new_n561_));
  INV        g539(.A(new_new_n236_), .Y(new_new_n562_));
  NO2        g540(.A(new_new_n562_), .B(new_new_n537_), .Y(new_new_n563_));
  NO3        g541(.A(new_new_n563_), .B(new_new_n560_), .C(new_new_n558_), .Y(new_new_n564_));
  INV        g542(.A(new_new_n194_), .Y(new_new_n565_));
  INV        g543(.A(new_new_n564_), .Y(new_new_n566_));
  INV        g544(.A(new_new_n522_), .Y(new_new_n567_));
  OA210      g545(.A0(new_new_n271_), .A1(new_new_n161_), .B0(new_new_n270_), .Y(new_new_n568_));
  NA2        g546(.A(new_new_n567_), .B(new_new_n561_), .Y(new_new_n569_));
  NA2        g547(.A(new_new_n413_), .B(new_new_n300_), .Y(new_new_n570_));
  NAi21      g548(.An(i_9_), .B(i_5_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n571_), .B(new_new_n235_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n572_), .B(new_new_n353_), .Y(new_new_n573_));
  OAI220     g551(.A0(new_new_n573_), .A1(new_new_n84_), .B0(new_new_n570_), .B1(new_new_n142_), .Y(new_new_n574_));
  NO2        g552(.A(new_new_n574_), .B(new_new_n291_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n575_), .B(new_new_n569_), .Y(new_new_n576_));
  NO3        g554(.A(new_new_n576_), .B(new_new_n566_), .C(new_new_n554_), .Y(new_new_n577_));
  NO2        g555(.A(i_0_), .B(new_new_n435_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n170_), .B(new_new_n164_), .Y(new_new_n579_));
  AOI210     g557(.A0(new_new_n579_), .A1(new_new_n542_), .B0(new_new_n137_), .Y(new_new_n580_));
  NO3        g558(.A(new_new_n155_), .B(new_new_n228_), .C(i_0_), .Y(new_new_n581_));
  OAI210     g559(.A0(new_new_n581_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n582_));
  INV        g560(.A(new_new_n582_), .Y(new_new_n583_));
  NO2        g561(.A(new_new_n169_), .B(new_new_n91_), .Y(new_new_n584_));
  AOI210     g562(.A0(new_new_n584_), .A1(new_new_n578_), .B0(new_new_n105_), .Y(new_new_n585_));
  OR2        g563(.A(new_new_n585_), .B(i_5_), .Y(new_new_n586_));
  AOI210     g564(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n143_), .Y(new_new_n587_));
  NA2        g565(.A(new_new_n587_), .B(new_new_n568_), .Y(new_new_n588_));
  NO3        g566(.A(new_new_n528_), .B(new_new_n52_), .C(new_new_n47_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n622_), .B(new_new_n589_), .Y(new_new_n590_));
  NA3        g568(.A(new_new_n231_), .B(new_new_n141_), .C(new_new_n140_), .Y(new_new_n591_));
  INV        g569(.A(new_new_n591_), .Y(new_new_n592_));
  NO3        g570(.A(new_new_n556_), .B(new_new_n157_), .C(new_new_n147_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n593_), .B(new_new_n592_), .Y(new_new_n594_));
  NA4        g572(.A(new_new_n594_), .B(new_new_n590_), .C(new_new_n588_), .D(new_new_n586_), .Y(new_new_n595_));
  NO2        g573(.A(new_new_n84_), .B(i_5_), .Y(new_new_n596_));
  NA3        g574(.A(new_new_n523_), .B(new_new_n106_), .C(new_new_n116_), .Y(new_new_n597_));
  INV        g575(.A(new_new_n597_), .Y(new_new_n598_));
  NA2        g576(.A(new_new_n598_), .B(new_new_n596_), .Y(new_new_n599_));
  NAi21      g577(.An(new_new_n168_), .B(new_new_n169_), .Y(new_new_n600_));
  NO4        g578(.A(new_new_n167_), .B(new_new_n155_), .C(i_0_), .D(i_12_), .Y(new_new_n601_));
  NA2        g579(.A(new_new_n601_), .B(new_new_n600_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n602_), .B(new_new_n599_), .Y(new_new_n603_));
  NO4        g581(.A(new_new_n603_), .B(new_new_n595_), .C(new_new_n583_), .D(new_new_n580_), .Y(new_new_n604_));
  OAI210     g582(.A0(new_new_n502_), .A1(new_new_n498_), .B0(new_new_n37_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n605_), .B(new_new_n345_), .Y(new_new_n606_));
  NA2        g584(.A(new_new_n606_), .B(new_new_n153_), .Y(new_new_n607_));
  NAi31      g585(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n68_), .B(new_new_n608_), .Y(new_new_n609_));
  AOI210     g587(.A0(new_new_n609_), .A1(new_new_n47_), .B0(new_new_n544_), .Y(new_new_n610_));
  AOI210     g588(.A0(new_new_n610_), .A1(new_new_n607_), .B0(new_new_n71_), .Y(new_new_n611_));
  INV        g589(.A(new_new_n225_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n612_), .B(new_new_n460_), .Y(new_new_n613_));
  NO3        g591(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n614_));
  OAI210     g592(.A0(new_new_n565_), .A1(new_new_n191_), .B0(new_new_n614_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n615_), .B(new_new_n435_), .Y(new_new_n616_));
  NO3        g594(.A(new_new_n616_), .B(new_new_n613_), .C(new_new_n611_), .Y(new_new_n617_));
  NA4        g595(.A(new_new_n617_), .B(new_new_n604_), .C(new_new_n577_), .D(new_new_n541_), .Y(ori4));
  INV        g596(.A(i_6_), .Y(new_new_n621_));
  INV        g597(.A(new_new_n275_), .Y(new_new_n622_));
endmodule


