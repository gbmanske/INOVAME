//Benchmark atmr_9sym_175_0.0313

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n166_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  NA2        o002(.A(i_4_), .B(ori_ori_n12_), .Y(ori_ori_n13_));
  INV        o003(.A(i_5_), .Y(ori_ori_n14_));
  NOi21      o004(.An(i_3_), .B(i_7_), .Y(ori_ori_n15_));
  INV        o005(.A(i_0_), .Y(ori_ori_n16_));
  NOi21      o006(.An(i_1_), .B(i_3_), .Y(ori_ori_n17_));
  INV        o007(.A(i_4_), .Y(ori_ori_n18_));
  NA2        o008(.A(i_0_), .B(ori_ori_n18_), .Y(ori_ori_n19_));
  INV        o009(.A(i_7_), .Y(ori_ori_n20_));
  NA3        o010(.A(i_6_), .B(i_5_), .C(ori_ori_n20_), .Y(ori_ori_n21_));
  NOi21      o011(.An(i_8_), .B(i_6_), .Y(ori_ori_n22_));
  NOi21      o012(.An(i_1_), .B(i_8_), .Y(ori_ori_n23_));
  AOI220     o013(.A0(ori_ori_n23_), .A1(i_2_), .B0(ori_ori_n22_), .B1(i_5_), .Y(ori_ori_n24_));
  AOI210     o014(.A0(ori_ori_n24_), .A1(ori_ori_n21_), .B0(ori_ori_n19_), .Y(ori_ori_n25_));
  NA2        o015(.A(ori_ori_n25_), .B(ori_ori_n11_), .Y(ori_ori_n26_));
  NA2        o016(.A(i_0_), .B(ori_ori_n14_), .Y(ori_ori_n27_));
  NA2        o017(.A(ori_ori_n16_), .B(i_5_), .Y(ori_ori_n28_));
  NO2        o018(.A(i_2_), .B(i_4_), .Y(ori_ori_n29_));
  NA3        o019(.A(ori_ori_n29_), .B(i_6_), .C(i_8_), .Y(ori_ori_n30_));
  AOI210     o020(.A0(ori_ori_n28_), .A1(ori_ori_n27_), .B0(ori_ori_n30_), .Y(ori_ori_n31_));
  INV        o021(.A(i_2_), .Y(ori_ori_n32_));
  NOi21      o022(.An(i_5_), .B(i_0_), .Y(ori_ori_n33_));
  NOi21      o023(.An(i_6_), .B(i_8_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_7_), .B(i_1_), .Y(ori_ori_n35_));
  NOi21      o025(.An(i_5_), .B(i_6_), .Y(ori_ori_n36_));
  AOI220     o026(.A0(ori_ori_n36_), .A1(ori_ori_n35_), .B0(ori_ori_n34_), .B1(ori_ori_n33_), .Y(ori_ori_n37_));
  NO3        o027(.A(ori_ori_n37_), .B(ori_ori_n32_), .C(i_4_), .Y(ori_ori_n38_));
  NOi21      o028(.An(i_0_), .B(i_4_), .Y(ori_ori_n39_));
  NOi21      o029(.An(i_7_), .B(i_5_), .Y(ori_ori_n40_));
  AN2        o030(.A(ori_ori_n40_), .B(ori_ori_n39_), .Y(ori_ori_n41_));
  INV        o031(.A(i_1_), .Y(ori_ori_n42_));
  NOi21      o032(.An(i_3_), .B(i_0_), .Y(ori_ori_n43_));
  NA2        o033(.A(ori_ori_n43_), .B(ori_ori_n42_), .Y(ori_ori_n44_));
  NA3        o034(.A(i_6_), .B(ori_ori_n14_), .C(i_7_), .Y(ori_ori_n45_));
  AOI210     o035(.A0(ori_ori_n45_), .A1(ori_ori_n21_), .B0(ori_ori_n44_), .Y(ori_ori_n46_));
  NO4        o036(.A(ori_ori_n46_), .B(ori_ori_n41_), .C(ori_ori_n38_), .D(ori_ori_n31_), .Y(ori_ori_n47_));
  NOi21      o037(.An(i_4_), .B(i_0_), .Y(ori_ori_n48_));
  NO2        o038(.A(ori_ori_n22_), .B(ori_ori_n15_), .Y(ori_ori_n49_));
  NA2        o039(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n50_));
  NOi21      o040(.An(i_2_), .B(i_8_), .Y(ori_ori_n51_));
  NO2        o041(.A(ori_ori_n50_), .B(ori_ori_n49_), .Y(ori_ori_n52_));
  INV        o042(.A(ori_ori_n52_), .Y(ori_ori_n53_));
  NOi31      o043(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n54_));
  NA2        o044(.A(ori_ori_n54_), .B(i_0_), .Y(ori_ori_n55_));
  NOi21      o045(.An(i_4_), .B(i_3_), .Y(ori_ori_n56_));
  NOi21      o046(.An(i_1_), .B(i_4_), .Y(ori_ori_n57_));
  OAI210     o047(.A0(ori_ori_n57_), .A1(ori_ori_n56_), .B0(ori_ori_n51_), .Y(ori_ori_n58_));
  NA2        o048(.A(ori_ori_n58_), .B(ori_ori_n55_), .Y(ori_ori_n59_));
  AN2        o049(.A(i_8_), .B(i_7_), .Y(ori_ori_n60_));
  NOi21      o050(.An(i_8_), .B(i_7_), .Y(ori_ori_n61_));
  NA3        o051(.A(ori_ori_n61_), .B(ori_ori_n56_), .C(i_6_), .Y(ori_ori_n62_));
  INV        o052(.A(ori_ori_n62_), .Y(ori_ori_n63_));
  AOI220     o053(.A0(ori_ori_n63_), .A1(ori_ori_n32_), .B0(ori_ori_n59_), .B1(ori_ori_n36_), .Y(ori_ori_n64_));
  NA4        o054(.A(ori_ori_n64_), .B(ori_ori_n53_), .C(ori_ori_n47_), .D(ori_ori_n26_), .Y(ori_ori_n65_));
  NA2        o055(.A(i_8_), .B(i_7_), .Y(ori_ori_n66_));
  NO3        o056(.A(ori_ori_n66_), .B(ori_ori_n13_), .C(i_1_), .Y(ori_ori_n67_));
  NA2        o057(.A(i_8_), .B(ori_ori_n20_), .Y(ori_ori_n68_));
  NOi21      o058(.An(i_1_), .B(i_2_), .Y(ori_ori_n69_));
  NO2        o059(.A(ori_ori_n166_), .B(ori_ori_n68_), .Y(ori_ori_n70_));
  OAI210     o060(.A0(ori_ori_n70_), .A1(ori_ori_n67_), .B0(ori_ori_n14_), .Y(ori_ori_n71_));
  NA3        o061(.A(ori_ori_n61_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n72_));
  NA3        o062(.A(ori_ori_n23_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n73_));
  NA2        o063(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NOi32      o064(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(ori_ori_n75_));
  NA2        o065(.A(ori_ori_n75_), .B(i_3_), .Y(ori_ori_n76_));
  NA2        o066(.A(ori_ori_n17_), .B(i_6_), .Y(ori_ori_n77_));
  NA2        o067(.A(ori_ori_n77_), .B(ori_ori_n76_), .Y(ori_ori_n78_));
  NO2        o068(.A(i_0_), .B(i_4_), .Y(ori_ori_n79_));
  AOI220     o069(.A0(ori_ori_n79_), .A1(ori_ori_n78_), .B0(ori_ori_n74_), .B1(ori_ori_n56_), .Y(ori_ori_n80_));
  NA2        o070(.A(ori_ori_n80_), .B(ori_ori_n71_), .Y(ori_ori_n81_));
  INV        o071(.A(ori_ori_n34_), .Y(ori_ori_n82_));
  NOi21      o072(.An(i_7_), .B(i_8_), .Y(ori_ori_n83_));
  OAI210     o073(.A0(i_8_), .A1(ori_ori_n11_), .B0(ori_ori_n82_), .Y(ori_ori_n84_));
  NA2        o074(.A(ori_ori_n84_), .B(ori_ori_n69_), .Y(ori_ori_n85_));
  AOI220     o075(.A0(ori_ori_n43_), .A1(ori_ori_n42_), .B0(ori_ori_n17_), .B1(ori_ori_n32_), .Y(ori_ori_n86_));
  NA3        o076(.A(ori_ori_n18_), .B(i_5_), .C(i_7_), .Y(ori_ori_n87_));
  NA2        o077(.A(i_4_), .B(i_5_), .Y(ori_ori_n88_));
  NA3        o078(.A(ori_ori_n66_), .B(ori_ori_n17_), .C(ori_ori_n16_), .Y(ori_ori_n89_));
  OAI220     o079(.A0(ori_ori_n89_), .A1(ori_ori_n88_), .B0(ori_ori_n87_), .B1(ori_ori_n86_), .Y(ori_ori_n90_));
  INV        o080(.A(ori_ori_n90_), .Y(ori_ori_n91_));
  NA3        o081(.A(ori_ori_n61_), .B(ori_ori_n32_), .C(i_3_), .Y(ori_ori_n92_));
  NA2        o082(.A(ori_ori_n42_), .B(i_6_), .Y(ori_ori_n93_));
  AOI210     o083(.A0(ori_ori_n93_), .A1(ori_ori_n19_), .B0(ori_ori_n92_), .Y(ori_ori_n94_));
  NOi21      o084(.An(i_2_), .B(i_1_), .Y(ori_ori_n95_));
  AN3        o085(.A(ori_ori_n83_), .B(ori_ori_n95_), .C(ori_ori_n48_), .Y(ori_ori_n96_));
  NAi21      o086(.An(i_6_), .B(i_0_), .Y(ori_ori_n97_));
  NA3        o087(.A(ori_ori_n57_), .B(i_5_), .C(ori_ori_n20_), .Y(ori_ori_n98_));
  NOi21      o088(.An(i_4_), .B(i_6_), .Y(ori_ori_n99_));
  NOi21      o089(.An(i_5_), .B(i_3_), .Y(ori_ori_n100_));
  NA3        o090(.A(ori_ori_n100_), .B(ori_ori_n69_), .C(ori_ori_n99_), .Y(ori_ori_n101_));
  OAI210     o091(.A0(ori_ori_n98_), .A1(ori_ori_n97_), .B0(ori_ori_n101_), .Y(ori_ori_n102_));
  NO3        o092(.A(ori_ori_n102_), .B(ori_ori_n96_), .C(ori_ori_n94_), .Y(ori_ori_n103_));
  AOI220     o093(.A0(i_6_), .A1(i_7_), .B0(ori_ori_n22_), .B1(i_5_), .Y(ori_ori_n104_));
  NOi31      o094(.An(ori_ori_n48_), .B(ori_ori_n104_), .C(i_2_), .Y(ori_ori_n105_));
  NA2        o095(.A(ori_ori_n61_), .B(ori_ori_n12_), .Y(ori_ori_n106_));
  NA2        o096(.A(ori_ori_n34_), .B(ori_ori_n14_), .Y(ori_ori_n107_));
  NOi21      o097(.An(i_3_), .B(i_1_), .Y(ori_ori_n108_));
  NA2        o098(.A(ori_ori_n108_), .B(i_4_), .Y(ori_ori_n109_));
  AOI210     o099(.A0(ori_ori_n107_), .A1(ori_ori_n106_), .B0(ori_ori_n109_), .Y(ori_ori_n110_));
  AOI220     o100(.A0(ori_ori_n83_), .A1(ori_ori_n14_), .B0(ori_ori_n99_), .B1(ori_ori_n20_), .Y(ori_ori_n111_));
  NOi31      o101(.An(ori_ori_n43_), .B(ori_ori_n111_), .C(ori_ori_n32_), .Y(ori_ori_n112_));
  NO3        o102(.A(ori_ori_n112_), .B(ori_ori_n110_), .C(ori_ori_n105_), .Y(ori_ori_n113_));
  NA4        o103(.A(ori_ori_n113_), .B(ori_ori_n103_), .C(ori_ori_n91_), .D(ori_ori_n85_), .Y(ori_ori_n114_));
  NA2        o104(.A(ori_ori_n51_), .B(ori_ori_n15_), .Y(ori_ori_n115_));
  NOi31      o105(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n116_));
  NOi31      o106(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n117_));
  OAI210     o107(.A0(ori_ori_n117_), .A1(ori_ori_n116_), .B0(i_7_), .Y(ori_ori_n118_));
  NA2        o108(.A(ori_ori_n118_), .B(ori_ori_n115_), .Y(ori_ori_n119_));
  NA2        o109(.A(ori_ori_n119_), .B(ori_ori_n39_), .Y(ori_ori_n120_));
  NA2        o110(.A(ori_ori_n56_), .B(ori_ori_n35_), .Y(ori_ori_n121_));
  AOI210     o111(.A0(ori_ori_n121_), .A1(ori_ori_n72_), .B0(ori_ori_n28_), .Y(ori_ori_n122_));
  NA4        o112(.A(ori_ori_n60_), .B(ori_ori_n95_), .C(ori_ori_n16_), .D(ori_ori_n12_), .Y(ori_ori_n123_));
  NAi31      o113(.An(ori_ori_n97_), .B(ori_ori_n83_), .C(ori_ori_n95_), .Y(ori_ori_n124_));
  NA3        o114(.A(ori_ori_n61_), .B(ori_ori_n54_), .C(i_6_), .Y(ori_ori_n125_));
  NA3        o115(.A(ori_ori_n125_), .B(ori_ori_n124_), .C(ori_ori_n123_), .Y(ori_ori_n126_));
  NOi21      o116(.An(i_0_), .B(i_2_), .Y(ori_ori_n127_));
  NA3        o117(.A(ori_ori_n127_), .B(ori_ori_n35_), .C(ori_ori_n99_), .Y(ori_ori_n128_));
  NA3        o118(.A(ori_ori_n48_), .B(ori_ori_n40_), .C(ori_ori_n17_), .Y(ori_ori_n129_));
  NOi32      o119(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n130_));
  NA2        o120(.A(ori_ori_n130_), .B(ori_ori_n116_), .Y(ori_ori_n131_));
  NA3        o121(.A(ori_ori_n127_), .B(ori_ori_n56_), .C(ori_ori_n34_), .Y(ori_ori_n132_));
  NA4        o122(.A(ori_ori_n132_), .B(ori_ori_n131_), .C(ori_ori_n129_), .D(ori_ori_n128_), .Y(ori_ori_n133_));
  NA3        o123(.A(ori_ori_n54_), .B(i_6_), .C(ori_ori_n14_), .Y(ori_ori_n134_));
  NA4        o124(.A(ori_ori_n57_), .B(ori_ori_n36_), .C(ori_ori_n16_), .D(i_8_), .Y(ori_ori_n135_));
  NA4        o125(.A(ori_ori_n57_), .B(ori_ori_n43_), .C(i_5_), .D(ori_ori_n20_), .Y(ori_ori_n136_));
  NA3        o126(.A(ori_ori_n136_), .B(ori_ori_n135_), .C(ori_ori_n134_), .Y(ori_ori_n137_));
  NO4        o127(.A(ori_ori_n137_), .B(ori_ori_n133_), .C(ori_ori_n126_), .D(ori_ori_n122_), .Y(ori_ori_n138_));
  NOi21      o128(.An(i_5_), .B(i_2_), .Y(ori_ori_n139_));
  AOI220     o129(.A0(ori_ori_n139_), .A1(ori_ori_n83_), .B0(ori_ori_n60_), .B1(ori_ori_n29_), .Y(ori_ori_n140_));
  AOI210     o130(.A0(ori_ori_n140_), .A1(ori_ori_n115_), .B0(ori_ori_n93_), .Y(ori_ori_n141_));
  NO4        o131(.A(i_2_), .B(ori_ori_n18_), .C(ori_ori_n11_), .D(ori_ori_n14_), .Y(ori_ori_n142_));
  NA2        o132(.A(i_2_), .B(i_4_), .Y(ori_ori_n143_));
  AOI210     o133(.A0(ori_ori_n97_), .A1(i_3_), .B0(ori_ori_n143_), .Y(ori_ori_n144_));
  NO2        o134(.A(i_8_), .B(i_7_), .Y(ori_ori_n145_));
  OA210      o135(.A0(ori_ori_n144_), .A1(ori_ori_n142_), .B0(ori_ori_n145_), .Y(ori_ori_n146_));
  NA3        o136(.A(ori_ori_n108_), .B(i_0_), .C(ori_ori_n20_), .Y(ori_ori_n147_));
  INV        o137(.A(ori_ori_n147_), .Y(ori_ori_n148_));
  NO3        o138(.A(ori_ori_n148_), .B(ori_ori_n146_), .C(ori_ori_n141_), .Y(ori_ori_n149_));
  NA2        o139(.A(ori_ori_n83_), .B(ori_ori_n12_), .Y(ori_ori_n150_));
  NA3        o140(.A(i_2_), .B(i_1_), .C(ori_ori_n14_), .Y(ori_ori_n151_));
  NA2        o141(.A(ori_ori_n48_), .B(i_3_), .Y(ori_ori_n152_));
  AOI210     o142(.A0(ori_ori_n152_), .A1(ori_ori_n151_), .B0(ori_ori_n150_), .Y(ori_ori_n153_));
  NA3        o143(.A(ori_ori_n127_), .B(ori_ori_n61_), .C(ori_ori_n99_), .Y(ori_ori_n154_));
  OAI210     o144(.A0(ori_ori_n92_), .A1(ori_ori_n28_), .B0(ori_ori_n154_), .Y(ori_ori_n155_));
  NA4        o145(.A(ori_ori_n100_), .B(ori_ori_n60_), .C(ori_ori_n42_), .D(ori_ori_n18_), .Y(ori_ori_n156_));
  NA3        o146(.A(ori_ori_n51_), .B(ori_ori_n33_), .C(ori_ori_n15_), .Y(ori_ori_n157_));
  NOi31      o147(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n158_));
  OAI210     o148(.A0(ori_ori_n130_), .A1(ori_ori_n75_), .B0(ori_ori_n158_), .Y(ori_ori_n159_));
  NA3        o149(.A(ori_ori_n159_), .B(ori_ori_n157_), .C(ori_ori_n156_), .Y(ori_ori_n160_));
  NO3        o150(.A(ori_ori_n160_), .B(ori_ori_n155_), .C(ori_ori_n153_), .Y(ori_ori_n161_));
  NA4        o151(.A(ori_ori_n161_), .B(ori_ori_n149_), .C(ori_ori_n138_), .D(ori_ori_n120_), .Y(ori_ori_n162_));
  OR4        o152(.A(ori_ori_n162_), .B(ori_ori_n114_), .C(ori_ori_n81_), .D(ori_ori_n65_), .Y(ori00));
  INV        o153(.A(i_2_), .Y(ori_ori_n166_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NO2        m008(.A(mai_mai_n16_), .B(mai_mai_n13_), .Y(mai_mai_n19_));
  INV        m009(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m010(.A(i_0_), .B(mai_mai_n20_), .Y(mai_mai_n21_));
  INV        m011(.A(i_7_), .Y(mai_mai_n22_));
  NA3        m012(.A(i_6_), .B(i_5_), .C(mai_mai_n22_), .Y(mai_mai_n23_));
  NOi21      m013(.An(i_8_), .B(i_6_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_1_), .B(i_8_), .Y(mai_mai_n25_));
  AOI220     m015(.A0(mai_mai_n25_), .A1(i_2_), .B0(mai_mai_n24_), .B1(i_5_), .Y(mai_mai_n26_));
  AOI210     m016(.A0(mai_mai_n26_), .A1(mai_mai_n23_), .B0(mai_mai_n21_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n27_), .A1(mai_mai_n11_), .B0(mai_mai_n19_), .Y(mai_mai_n28_));
  NA2        m018(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n29_));
  NA2        m019(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n30_));
  NO2        m020(.A(i_2_), .B(i_4_), .Y(mai_mai_n31_));
  NA3        m021(.A(mai_mai_n31_), .B(i_6_), .C(i_8_), .Y(mai_mai_n32_));
  AOI210     m022(.A0(mai_mai_n30_), .A1(mai_mai_n29_), .B0(mai_mai_n32_), .Y(mai_mai_n33_));
  INV        m023(.A(i_2_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_5_), .B(i_0_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_6_), .B(i_8_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_7_), .B(i_1_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_5_), .B(i_6_), .Y(mai_mai_n38_));
  AOI220     m028(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n36_), .B1(mai_mai_n35_), .Y(mai_mai_n39_));
  NO3        m029(.A(mai_mai_n39_), .B(mai_mai_n34_), .C(i_4_), .Y(mai_mai_n40_));
  NOi21      m030(.An(i_0_), .B(i_4_), .Y(mai_mai_n41_));
  XO2        m031(.A(i_1_), .B(i_3_), .Y(mai_mai_n42_));
  NOi21      m032(.An(i_7_), .B(i_5_), .Y(mai_mai_n43_));
  AN3        m033(.A(mai_mai_n43_), .B(mai_mai_n42_), .C(mai_mai_n41_), .Y(mai_mai_n44_));
  INV        m034(.A(i_1_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_3_), .B(i_0_), .Y(mai_mai_n46_));
  NA2        m036(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NA3        m037(.A(i_6_), .B(mai_mai_n14_), .C(i_7_), .Y(mai_mai_n48_));
  NO2        m038(.A(mai_mai_n48_), .B(mai_mai_n47_), .Y(mai_mai_n49_));
  NO4        m039(.A(mai_mai_n49_), .B(mai_mai_n44_), .C(mai_mai_n40_), .D(mai_mai_n33_), .Y(mai_mai_n50_));
  INV        m040(.A(i_8_), .Y(mai_mai_n51_));
  NA2        m041(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_4_), .B(i_0_), .Y(mai_mai_n53_));
  AOI210     m043(.A0(mai_mai_n53_), .A1(mai_mai_n24_), .B0(mai_mai_n15_), .Y(mai_mai_n54_));
  NA2        m044(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n55_));
  NOi21      m045(.An(i_2_), .B(i_8_), .Y(mai_mai_n56_));
  NO3        m046(.A(mai_mai_n56_), .B(mai_mai_n53_), .C(mai_mai_n41_), .Y(mai_mai_n57_));
  NO3        m047(.A(mai_mai_n57_), .B(mai_mai_n55_), .C(mai_mai_n54_), .Y(mai_mai_n58_));
  INV        m048(.A(mai_mai_n58_), .Y(mai_mai_n59_));
  NOi31      m049(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n60_));
  NA2        m050(.A(mai_mai_n60_), .B(i_0_), .Y(mai_mai_n61_));
  NOi21      m051(.An(i_4_), .B(i_3_), .Y(mai_mai_n62_));
  NOi21      m052(.An(i_1_), .B(i_4_), .Y(mai_mai_n63_));
  OAI210     m053(.A0(mai_mai_n63_), .A1(mai_mai_n62_), .B0(mai_mai_n56_), .Y(mai_mai_n64_));
  NA2        m054(.A(mai_mai_n64_), .B(mai_mai_n61_), .Y(mai_mai_n65_));
  AN2        m055(.A(i_8_), .B(i_7_), .Y(mai_mai_n66_));
  NA2        m056(.A(mai_mai_n66_), .B(mai_mai_n12_), .Y(mai_mai_n67_));
  NOi21      m057(.An(i_8_), .B(i_7_), .Y(mai_mai_n68_));
  NO2        m058(.A(mai_mai_n67_), .B(mai_mai_n55_), .Y(mai_mai_n69_));
  AOI220     m059(.A0(mai_mai_n69_), .A1(mai_mai_n34_), .B0(mai_mai_n65_), .B1(mai_mai_n38_), .Y(mai_mai_n70_));
  NA4        m060(.A(mai_mai_n70_), .B(mai_mai_n59_), .C(mai_mai_n50_), .D(mai_mai_n28_), .Y(mai_mai_n71_));
  NA2        m061(.A(i_8_), .B(i_7_), .Y(mai_mai_n72_));
  NO2        m062(.A(mai_mai_n72_), .B(i_1_), .Y(mai_mai_n73_));
  NA2        m063(.A(i_8_), .B(mai_mai_n22_), .Y(mai_mai_n74_));
  AOI220     m064(.A0(mai_mai_n46_), .A1(i_1_), .B0(mai_mai_n42_), .B1(i_2_), .Y(mai_mai_n75_));
  NOi21      m065(.An(i_1_), .B(i_2_), .Y(mai_mai_n76_));
  NA3        m066(.A(mai_mai_n76_), .B(mai_mai_n53_), .C(i_6_), .Y(mai_mai_n77_));
  OAI210     m067(.A0(mai_mai_n75_), .A1(mai_mai_n74_), .B0(mai_mai_n77_), .Y(mai_mai_n78_));
  OAI210     m068(.A0(mai_mai_n78_), .A1(mai_mai_n73_), .B0(mai_mai_n14_), .Y(mai_mai_n79_));
  NA3        m069(.A(mai_mai_n68_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n80_));
  INV        m070(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NOi32      m071(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n82_), .B(i_3_), .Y(mai_mai_n83_));
  NA3        m073(.A(mai_mai_n18_), .B(i_2_), .C(i_6_), .Y(mai_mai_n84_));
  NA2        m074(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n85_));
  NO2        m075(.A(i_0_), .B(i_4_), .Y(mai_mai_n86_));
  AOI220     m076(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n81_), .B1(mai_mai_n62_), .Y(mai_mai_n87_));
  NA2        m077(.A(mai_mai_n87_), .B(mai_mai_n79_), .Y(mai_mai_n88_));
  NAi21      m078(.An(i_3_), .B(i_6_), .Y(mai_mai_n89_));
  NO2        m079(.A(mai_mai_n89_), .B(mai_mai_n51_), .Y(mai_mai_n90_));
  NA2        m080(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n91_));
  NOi21      m081(.An(i_7_), .B(i_8_), .Y(mai_mai_n92_));
  NOi31      m082(.An(i_6_), .B(i_5_), .C(i_7_), .Y(mai_mai_n93_));
  AOI210     m083(.A0(mai_mai_n92_), .A1(mai_mai_n12_), .B0(mai_mai_n93_), .Y(mai_mai_n94_));
  OAI210     m084(.A0(mai_mai_n94_), .A1(mai_mai_n11_), .B0(mai_mai_n91_), .Y(mai_mai_n95_));
  OAI210     m085(.A0(mai_mai_n95_), .A1(mai_mai_n90_), .B0(mai_mai_n76_), .Y(mai_mai_n96_));
  NA3        m086(.A(mai_mai_n24_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n97_));
  AOI210     m087(.A0(mai_mai_n21_), .A1(mai_mai_n52_), .B0(mai_mai_n97_), .Y(mai_mai_n98_));
  INV        m088(.A(mai_mai_n98_), .Y(mai_mai_n99_));
  NA3        m089(.A(mai_mai_n68_), .B(mai_mai_n34_), .C(i_3_), .Y(mai_mai_n100_));
  NA2        m090(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n101_));
  AOI210     m091(.A0(mai_mai_n101_), .A1(mai_mai_n21_), .B0(mai_mai_n100_), .Y(mai_mai_n102_));
  NOi21      m092(.An(i_2_), .B(i_1_), .Y(mai_mai_n103_));
  AN3        m093(.A(mai_mai_n92_), .B(mai_mai_n103_), .C(mai_mai_n53_), .Y(mai_mai_n104_));
  NAi21      m094(.An(i_6_), .B(i_0_), .Y(mai_mai_n105_));
  NA3        m095(.A(mai_mai_n63_), .B(i_5_), .C(mai_mai_n22_), .Y(mai_mai_n106_));
  NOi21      m096(.An(i_4_), .B(i_6_), .Y(mai_mai_n107_));
  NO2        m097(.A(mai_mai_n106_), .B(mai_mai_n105_), .Y(mai_mai_n108_));
  NA2        m098(.A(mai_mai_n76_), .B(mai_mai_n36_), .Y(mai_mai_n109_));
  NOi21      m099(.An(mai_mai_n43_), .B(mai_mai_n109_), .Y(mai_mai_n110_));
  NO4        m100(.A(mai_mai_n110_), .B(mai_mai_n108_), .C(mai_mai_n104_), .D(mai_mai_n102_), .Y(mai_mai_n111_));
  NOi21      m101(.An(i_6_), .B(i_1_), .Y(mai_mai_n112_));
  AOI220     m102(.A0(mai_mai_n112_), .A1(i_7_), .B0(mai_mai_n24_), .B1(i_5_), .Y(mai_mai_n113_));
  NOi31      m103(.An(mai_mai_n53_), .B(mai_mai_n113_), .C(i_2_), .Y(mai_mai_n114_));
  NA2        m104(.A(mai_mai_n68_), .B(mai_mai_n12_), .Y(mai_mai_n115_));
  NA2        m105(.A(mai_mai_n36_), .B(mai_mai_n14_), .Y(mai_mai_n116_));
  NOi21      m106(.An(i_3_), .B(i_1_), .Y(mai_mai_n117_));
  NA2        m107(.A(mai_mai_n117_), .B(i_4_), .Y(mai_mai_n118_));
  AOI210     m108(.A0(mai_mai_n116_), .A1(mai_mai_n115_), .B0(mai_mai_n118_), .Y(mai_mai_n119_));
  AOI220     m109(.A0(mai_mai_n92_), .A1(mai_mai_n14_), .B0(mai_mai_n107_), .B1(mai_mai_n22_), .Y(mai_mai_n120_));
  NOi31      m110(.An(mai_mai_n46_), .B(mai_mai_n120_), .C(mai_mai_n34_), .Y(mai_mai_n121_));
  NO3        m111(.A(mai_mai_n121_), .B(mai_mai_n119_), .C(mai_mai_n114_), .Y(mai_mai_n122_));
  NA4        m112(.A(mai_mai_n122_), .B(mai_mai_n111_), .C(mai_mai_n99_), .D(mai_mai_n96_), .Y(mai_mai_n123_));
  NA2        m113(.A(mai_mai_n56_), .B(mai_mai_n15_), .Y(mai_mai_n124_));
  NOi31      m114(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n125_));
  NOi31      m115(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n126_));
  OAI210     m116(.A0(mai_mai_n126_), .A1(mai_mai_n125_), .B0(i_7_), .Y(mai_mai_n127_));
  NA3        m117(.A(mai_mai_n36_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n128_));
  NA4        m118(.A(mai_mai_n128_), .B(mai_mai_n127_), .C(mai_mai_n124_), .D(mai_mai_n109_), .Y(mai_mai_n129_));
  NA2        m119(.A(mai_mai_n129_), .B(mai_mai_n41_), .Y(mai_mai_n130_));
  INV        m120(.A(mai_mai_n62_), .Y(mai_mai_n131_));
  AOI210     m121(.A0(mai_mai_n131_), .A1(mai_mai_n80_), .B0(mai_mai_n30_), .Y(mai_mai_n132_));
  NA4        m122(.A(mai_mai_n66_), .B(mai_mai_n103_), .C(mai_mai_n17_), .D(mai_mai_n12_), .Y(mai_mai_n133_));
  NAi31      m123(.An(mai_mai_n105_), .B(mai_mai_n92_), .C(mai_mai_n103_), .Y(mai_mai_n134_));
  NA3        m124(.A(mai_mai_n68_), .B(mai_mai_n60_), .C(i_6_), .Y(mai_mai_n135_));
  NA3        m125(.A(mai_mai_n135_), .B(mai_mai_n134_), .C(mai_mai_n133_), .Y(mai_mai_n136_));
  NOi21      m126(.An(i_0_), .B(i_2_), .Y(mai_mai_n137_));
  NA3        m127(.A(mai_mai_n137_), .B(mai_mai_n37_), .C(mai_mai_n107_), .Y(mai_mai_n138_));
  NA3        m128(.A(mai_mai_n53_), .B(mai_mai_n43_), .C(mai_mai_n18_), .Y(mai_mai_n139_));
  NA2        m129(.A(mai_mai_n137_), .B(mai_mai_n62_), .Y(mai_mai_n140_));
  NA3        m130(.A(mai_mai_n140_), .B(mai_mai_n139_), .C(mai_mai_n138_), .Y(mai_mai_n141_));
  NA4        m131(.A(mai_mai_n60_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n142_));
  NA4        m132(.A(mai_mai_n63_), .B(mai_mai_n38_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n143_));
  NA2        m133(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NO4        m134(.A(mai_mai_n144_), .B(mai_mai_n141_), .C(mai_mai_n136_), .D(mai_mai_n132_), .Y(mai_mai_n145_));
  NOi21      m135(.An(i_5_), .B(i_2_), .Y(mai_mai_n146_));
  NA2        m136(.A(mai_mai_n146_), .B(mai_mai_n92_), .Y(mai_mai_n147_));
  AOI210     m137(.A0(mai_mai_n147_), .A1(mai_mai_n124_), .B0(mai_mai_n101_), .Y(mai_mai_n148_));
  NO3        m138(.A(i_2_), .B(mai_mai_n11_), .C(mai_mai_n14_), .Y(mai_mai_n149_));
  NA2        m139(.A(i_2_), .B(i_4_), .Y(mai_mai_n150_));
  AOI210     m140(.A0(mai_mai_n105_), .A1(mai_mai_n89_), .B0(mai_mai_n150_), .Y(mai_mai_n151_));
  NO2        m141(.A(i_8_), .B(i_7_), .Y(mai_mai_n152_));
  OA210      m142(.A0(mai_mai_n151_), .A1(mai_mai_n149_), .B0(mai_mai_n152_), .Y(mai_mai_n153_));
  NA2        m143(.A(mai_mai_n117_), .B(i_5_), .Y(mai_mai_n154_));
  NO2        m144(.A(mai_mai_n154_), .B(i_4_), .Y(mai_mai_n155_));
  NO3        m145(.A(mai_mai_n155_), .B(mai_mai_n153_), .C(mai_mai_n148_), .Y(mai_mai_n156_));
  NA2        m146(.A(mai_mai_n92_), .B(mai_mai_n12_), .Y(mai_mai_n157_));
  NA3        m147(.A(i_2_), .B(i_1_), .C(mai_mai_n14_), .Y(mai_mai_n158_));
  NA2        m148(.A(mai_mai_n53_), .B(i_3_), .Y(mai_mai_n159_));
  AOI210     m149(.A0(mai_mai_n159_), .A1(mai_mai_n158_), .B0(mai_mai_n157_), .Y(mai_mai_n160_));
  NA3        m150(.A(mai_mai_n66_), .B(mai_mai_n45_), .C(mai_mai_n20_), .Y(mai_mai_n161_));
  NA3        m151(.A(mai_mai_n93_), .B(mai_mai_n117_), .C(i_0_), .Y(mai_mai_n162_));
  NA2        m152(.A(mai_mai_n35_), .B(mai_mai_n15_), .Y(mai_mai_n163_));
  NA3        m153(.A(mai_mai_n163_), .B(mai_mai_n162_), .C(mai_mai_n161_), .Y(mai_mai_n164_));
  NO2        m154(.A(mai_mai_n164_), .B(mai_mai_n160_), .Y(mai_mai_n165_));
  NA4        m155(.A(mai_mai_n165_), .B(mai_mai_n156_), .C(mai_mai_n145_), .D(mai_mai_n130_), .Y(mai_mai_n166_));
  OR4        m156(.A(mai_mai_n166_), .B(mai_mai_n123_), .C(mai_mai_n88_), .D(mai_mai_n71_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  INV        u005(.A(i_0_), .Y(men_men_n16_));
  NOi21      u006(.An(i_1_), .B(i_3_), .Y(men_men_n17_));
  NA3        u007(.A(men_men_n17_), .B(men_men_n16_), .C(i_2_), .Y(men_men_n18_));
  NO2        u008(.A(men_men_n18_), .B(men_men_n13_), .Y(men_men_n19_));
  INV        u009(.A(i_4_), .Y(men_men_n20_));
  NA2        u010(.A(i_0_), .B(men_men_n20_), .Y(men_men_n21_));
  INV        u011(.A(i_7_), .Y(men_men_n22_));
  NA3        u012(.A(i_6_), .B(i_5_), .C(men_men_n22_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  NOi21      u014(.An(i_1_), .B(i_8_), .Y(men_men_n25_));
  AOI220     u015(.A0(men_men_n25_), .A1(i_2_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n26_));
  AOI210     u016(.A0(men_men_n26_), .A1(men_men_n23_), .B0(men_men_n21_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n11_), .B0(men_men_n19_), .Y(men_men_n28_));
  NA2        u018(.A(i_0_), .B(men_men_n14_), .Y(men_men_n29_));
  NA2        u019(.A(men_men_n16_), .B(i_5_), .Y(men_men_n30_));
  NO2        u020(.A(i_2_), .B(i_4_), .Y(men_men_n31_));
  NA3        u021(.A(men_men_n31_), .B(i_6_), .C(i_8_), .Y(men_men_n32_));
  AOI210     u022(.A0(men_men_n30_), .A1(men_men_n29_), .B0(men_men_n32_), .Y(men_men_n33_));
  INV        u023(.A(i_2_), .Y(men_men_n34_));
  NOi21      u024(.An(i_5_), .B(i_0_), .Y(men_men_n35_));
  NOi21      u025(.An(i_6_), .B(i_8_), .Y(men_men_n36_));
  NOi21      u026(.An(i_7_), .B(i_1_), .Y(men_men_n37_));
  NOi21      u027(.An(i_5_), .B(i_6_), .Y(men_men_n38_));
  AOI220     u028(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n36_), .B1(men_men_n35_), .Y(men_men_n39_));
  NO3        u029(.A(men_men_n39_), .B(men_men_n34_), .C(i_4_), .Y(men_men_n40_));
  NOi21      u030(.An(i_0_), .B(i_4_), .Y(men_men_n41_));
  XO2        u031(.A(i_1_), .B(i_3_), .Y(men_men_n42_));
  NOi21      u032(.An(i_7_), .B(i_5_), .Y(men_men_n43_));
  AN3        u033(.A(men_men_n43_), .B(men_men_n42_), .C(men_men_n41_), .Y(men_men_n44_));
  INV        u034(.A(i_1_), .Y(men_men_n45_));
  NOi21      u035(.An(i_3_), .B(i_0_), .Y(men_men_n46_));
  NA2        u036(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u037(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n48_));
  NO4        u038(.A(men_men_n48_), .B(men_men_n44_), .C(men_men_n40_), .D(men_men_n33_), .Y(men_men_n49_));
  INV        u039(.A(i_8_), .Y(men_men_n50_));
  NA2        u040(.A(i_1_), .B(men_men_n11_), .Y(men_men_n51_));
  NO4        u041(.A(men_men_n51_), .B(men_men_n29_), .C(i_2_), .D(men_men_n50_), .Y(men_men_n52_));
  NOi21      u042(.An(i_4_), .B(i_0_), .Y(men_men_n53_));
  INV        u043(.A(men_men_n15_), .Y(men_men_n54_));
  NA2        u044(.A(i_1_), .B(men_men_n14_), .Y(men_men_n55_));
  NOi21      u045(.An(i_2_), .B(i_8_), .Y(men_men_n56_));
  NO2        u046(.A(men_men_n56_), .B(men_men_n41_), .Y(men_men_n57_));
  NO3        u047(.A(men_men_n57_), .B(men_men_n55_), .C(men_men_n54_), .Y(men_men_n58_));
  NO2        u048(.A(men_men_n58_), .B(men_men_n52_), .Y(men_men_n59_));
  NOi31      u049(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n60_));
  NA2        u050(.A(men_men_n60_), .B(i_0_), .Y(men_men_n61_));
  NOi21      u051(.An(i_4_), .B(i_3_), .Y(men_men_n62_));
  NOi21      u052(.An(i_1_), .B(i_4_), .Y(men_men_n63_));
  OAI210     u053(.A0(men_men_n63_), .A1(men_men_n62_), .B0(men_men_n56_), .Y(men_men_n64_));
  NA2        u054(.A(men_men_n64_), .B(men_men_n61_), .Y(men_men_n65_));
  AN2        u055(.A(i_8_), .B(i_7_), .Y(men_men_n66_));
  NA2        u056(.A(men_men_n66_), .B(men_men_n12_), .Y(men_men_n67_));
  NOi21      u057(.An(i_8_), .B(i_7_), .Y(men_men_n68_));
  NA3        u058(.A(men_men_n68_), .B(men_men_n62_), .C(i_6_), .Y(men_men_n69_));
  OAI210     u059(.A0(men_men_n67_), .A1(men_men_n55_), .B0(men_men_n69_), .Y(men_men_n70_));
  AOI220     u060(.A0(men_men_n70_), .A1(men_men_n34_), .B0(men_men_n65_), .B1(men_men_n38_), .Y(men_men_n71_));
  NA4        u061(.A(men_men_n71_), .B(men_men_n59_), .C(men_men_n49_), .D(men_men_n28_), .Y(men_men_n72_));
  NA2        u062(.A(i_8_), .B(men_men_n22_), .Y(men_men_n73_));
  AOI220     u063(.A0(men_men_n46_), .A1(i_1_), .B0(men_men_n42_), .B1(i_2_), .Y(men_men_n74_));
  NOi21      u064(.An(i_1_), .B(i_2_), .Y(men_men_n75_));
  NO2        u065(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n76_));
  NA2        u066(.A(men_men_n76_), .B(men_men_n14_), .Y(men_men_n77_));
  NA3        u067(.A(men_men_n68_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n78_));
  NA3        u068(.A(men_men_n25_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n79_));
  NA2        u069(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NOi32      u070(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n81_));
  NA2        u071(.A(men_men_n81_), .B(i_3_), .Y(men_men_n82_));
  NA3        u072(.A(men_men_n17_), .B(i_2_), .C(i_6_), .Y(men_men_n83_));
  NA2        u073(.A(men_men_n83_), .B(men_men_n82_), .Y(men_men_n84_));
  NO2        u074(.A(i_0_), .B(i_4_), .Y(men_men_n85_));
  AOI220     u075(.A0(men_men_n85_), .A1(men_men_n84_), .B0(men_men_n80_), .B1(men_men_n62_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n86_), .B(men_men_n77_), .Y(men_men_n87_));
  NAi21      u077(.An(i_3_), .B(i_6_), .Y(men_men_n88_));
  NO3        u078(.A(men_men_n88_), .B(i_0_), .C(men_men_n50_), .Y(men_men_n89_));
  NA2        u079(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n90_));
  NOi21      u080(.An(i_7_), .B(i_8_), .Y(men_men_n91_));
  NOi31      u081(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n92_));
  AOI210     u082(.A0(men_men_n91_), .A1(men_men_n12_), .B0(men_men_n92_), .Y(men_men_n93_));
  OAI210     u083(.A0(men_men_n93_), .A1(men_men_n11_), .B0(men_men_n90_), .Y(men_men_n94_));
  OAI210     u084(.A0(men_men_n94_), .A1(men_men_n89_), .B0(men_men_n75_), .Y(men_men_n95_));
  NA3        u085(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n96_));
  AOI210     u086(.A0(men_men_n21_), .A1(men_men_n51_), .B0(men_men_n96_), .Y(men_men_n97_));
  AOI220     u087(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n17_), .B1(men_men_n34_), .Y(men_men_n98_));
  NA3        u088(.A(men_men_n20_), .B(i_5_), .C(i_7_), .Y(men_men_n99_));
  NO2        u089(.A(men_men_n99_), .B(men_men_n98_), .Y(men_men_n100_));
  NO2        u090(.A(men_men_n100_), .B(men_men_n97_), .Y(men_men_n101_));
  NA3        u091(.A(men_men_n68_), .B(men_men_n34_), .C(i_3_), .Y(men_men_n102_));
  NA2        u092(.A(men_men_n45_), .B(i_6_), .Y(men_men_n103_));
  AOI210     u093(.A0(men_men_n103_), .A1(men_men_n21_), .B0(men_men_n102_), .Y(men_men_n104_));
  NAi21      u094(.An(i_6_), .B(i_0_), .Y(men_men_n105_));
  NA3        u095(.A(men_men_n63_), .B(i_5_), .C(men_men_n22_), .Y(men_men_n106_));
  NOi21      u096(.An(i_4_), .B(i_6_), .Y(men_men_n107_));
  NOi21      u097(.An(i_5_), .B(i_3_), .Y(men_men_n108_));
  NA3        u098(.A(men_men_n108_), .B(men_men_n75_), .C(men_men_n107_), .Y(men_men_n109_));
  OAI210     u099(.A0(men_men_n106_), .A1(men_men_n105_), .B0(men_men_n109_), .Y(men_men_n110_));
  NA2        u100(.A(men_men_n75_), .B(men_men_n36_), .Y(men_men_n111_));
  NOi21      u101(.An(men_men_n43_), .B(men_men_n111_), .Y(men_men_n112_));
  NO3        u102(.A(men_men_n112_), .B(men_men_n110_), .C(men_men_n104_), .Y(men_men_n113_));
  NOi21      u103(.An(i_3_), .B(i_1_), .Y(men_men_n114_));
  NA3        u104(.A(men_men_n113_), .B(men_men_n101_), .C(men_men_n95_), .Y(men_men_n115_));
  NA2        u105(.A(men_men_n56_), .B(men_men_n15_), .Y(men_men_n116_));
  NOi31      u106(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n117_));
  NA2        u107(.A(men_men_n117_), .B(i_7_), .Y(men_men_n118_));
  NA3        u108(.A(men_men_n36_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n119_));
  NA4        u109(.A(men_men_n119_), .B(men_men_n118_), .C(men_men_n116_), .D(men_men_n111_), .Y(men_men_n120_));
  NA2        u110(.A(men_men_n120_), .B(men_men_n41_), .Y(men_men_n121_));
  NA2        u111(.A(men_men_n62_), .B(men_men_n37_), .Y(men_men_n122_));
  AOI210     u112(.A0(men_men_n122_), .A1(men_men_n78_), .B0(men_men_n30_), .Y(men_men_n123_));
  NA3        u113(.A(men_men_n68_), .B(men_men_n60_), .C(i_6_), .Y(men_men_n124_));
  INV        u114(.A(men_men_n124_), .Y(men_men_n125_));
  NA2        u115(.A(men_men_n37_), .B(men_men_n107_), .Y(men_men_n126_));
  NA2        u116(.A(men_men_n53_), .B(men_men_n43_), .Y(men_men_n127_));
  NOi32      u117(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n128_));
  NA2        u118(.A(men_men_n62_), .B(men_men_n36_), .Y(men_men_n129_));
  NA3        u119(.A(men_men_n129_), .B(men_men_n127_), .C(men_men_n126_), .Y(men_men_n130_));
  NA3        u120(.A(men_men_n60_), .B(men_men_n14_), .C(i_7_), .Y(men_men_n131_));
  NA4        u121(.A(men_men_n63_), .B(men_men_n38_), .C(men_men_n16_), .D(i_8_), .Y(men_men_n132_));
  NA4        u122(.A(men_men_n63_), .B(men_men_n46_), .C(i_5_), .D(men_men_n22_), .Y(men_men_n133_));
  NA3        u123(.A(men_men_n133_), .B(men_men_n132_), .C(men_men_n131_), .Y(men_men_n134_));
  NO4        u124(.A(men_men_n134_), .B(men_men_n130_), .C(men_men_n125_), .D(men_men_n123_), .Y(men_men_n135_));
  AOI210     u125(.A0(men_men_n66_), .A1(men_men_n31_), .B0(men_men_n91_), .Y(men_men_n136_));
  AOI210     u126(.A0(men_men_n136_), .A1(men_men_n116_), .B0(men_men_n103_), .Y(men_men_n137_));
  NO3        u127(.A(i_2_), .B(men_men_n20_), .C(men_men_n11_), .Y(men_men_n138_));
  NA2        u128(.A(i_2_), .B(i_4_), .Y(men_men_n139_));
  NO2        u129(.A(men_men_n105_), .B(men_men_n139_), .Y(men_men_n140_));
  NO2        u130(.A(i_8_), .B(i_7_), .Y(men_men_n141_));
  OA210      u131(.A0(men_men_n140_), .A1(men_men_n138_), .B0(men_men_n141_), .Y(men_men_n142_));
  NA4        u132(.A(men_men_n114_), .B(i_0_), .C(i_5_), .D(men_men_n22_), .Y(men_men_n143_));
  NO2        u133(.A(men_men_n143_), .B(i_4_), .Y(men_men_n144_));
  NO3        u134(.A(men_men_n144_), .B(men_men_n142_), .C(men_men_n137_), .Y(men_men_n145_));
  NA2        u135(.A(men_men_n91_), .B(men_men_n12_), .Y(men_men_n146_));
  NA2        u136(.A(i_2_), .B(men_men_n14_), .Y(men_men_n147_));
  INV        u137(.A(men_men_n53_), .Y(men_men_n148_));
  AOI210     u138(.A0(men_men_n148_), .A1(men_men_n147_), .B0(men_men_n146_), .Y(men_men_n149_));
  NA2        u139(.A(men_men_n68_), .B(men_men_n107_), .Y(men_men_n150_));
  OAI210     u140(.A0(men_men_n102_), .A1(men_men_n30_), .B0(men_men_n150_), .Y(men_men_n151_));
  NA4        u141(.A(men_men_n108_), .B(men_men_n66_), .C(men_men_n45_), .D(men_men_n20_), .Y(men_men_n152_));
  NA3        u142(.A(men_men_n92_), .B(men_men_n114_), .C(i_0_), .Y(men_men_n153_));
  NA3        u143(.A(men_men_n56_), .B(men_men_n35_), .C(men_men_n15_), .Y(men_men_n154_));
  NOi31      u144(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n155_));
  OAI210     u145(.A0(men_men_n128_), .A1(men_men_n81_), .B0(men_men_n155_), .Y(men_men_n156_));
  NA4        u146(.A(men_men_n156_), .B(men_men_n154_), .C(men_men_n153_), .D(men_men_n152_), .Y(men_men_n157_));
  NO3        u147(.A(men_men_n157_), .B(men_men_n151_), .C(men_men_n149_), .Y(men_men_n158_));
  NA4        u148(.A(men_men_n158_), .B(men_men_n145_), .C(men_men_n135_), .D(men_men_n121_), .Y(men_men_n159_));
  OR4        u149(.A(men_men_n159_), .B(men_men_n115_), .C(men_men_n87_), .D(men_men_n72_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule