// Benchmark "top" written by ABC on Fri Jun 21 17:49:20 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n125_, new_new_n126_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n261_,
    new_new_n262_, new_new_n263_, new_new_n264_, new_new_n265_,
    new_new_n266_, new_new_n267_, new_new_n268_, new_new_n269_,
    new_new_n270_, new_new_n271_, new_new_n272_, new_new_n273_,
    new_new_n274_, new_new_n275_, new_new_n276_, new_new_n277_,
    new_new_n278_, new_new_n279_, new_new_n280_, new_new_n281_,
    new_new_n282_, new_new_n283_, new_new_n284_, new_new_n285_,
    new_new_n286_, new_new_n287_, new_new_n288_, new_new_n289_,
    new_new_n290_, new_new_n291_, new_new_n292_, new_new_n293_,
    new_new_n294_, new_new_n295_, new_new_n296_, new_new_n297_,
    new_new_n298_, new_new_n299_, new_new_n300_, new_new_n301_,
    new_new_n302_, new_new_n303_, new_new_n304_, new_new_n305_,
    new_new_n306_, new_new_n307_, new_new_n308_, new_new_n309_,
    new_new_n310_, new_new_n311_, new_new_n312_, new_new_n313_,
    new_new_n314_, new_new_n315_, new_new_n316_, new_new_n317_,
    new_new_n318_, new_new_n319_, new_new_n320_, new_new_n321_,
    new_new_n322_, new_new_n323_, new_new_n324_, new_new_n325_,
    new_new_n326_, new_new_n327_, new_new_n328_, new_new_n329_,
    new_new_n330_, new_new_n331_, new_new_n332_, new_new_n333_,
    new_new_n334_, new_new_n335_, new_new_n336_, new_new_n337_,
    new_new_n338_, new_new_n339_, new_new_n340_, new_new_n341_,
    new_new_n342_, new_new_n343_, new_new_n344_, new_new_n345_,
    new_new_n346_, new_new_n347_, new_new_n348_, new_new_n349_,
    new_new_n350_, new_new_n351_, new_new_n353_, new_new_n354_,
    new_new_n355_, new_new_n356_, new_new_n357_, new_new_n358_,
    new_new_n359_, new_new_n360_, new_new_n361_, new_new_n362_,
    new_new_n363_, new_new_n364_, new_new_n365_, new_new_n366_,
    new_new_n367_, new_new_n368_, new_new_n369_, new_new_n370_,
    new_new_n371_, new_new_n372_, new_new_n373_, new_new_n374_,
    new_new_n375_, new_new_n376_, new_new_n377_, new_new_n378_,
    new_new_n379_, new_new_n380_, new_new_n381_, new_new_n382_,
    new_new_n383_, new_new_n384_, new_new_n385_, new_new_n386_,
    new_new_n387_, new_new_n388_, new_new_n389_, new_new_n390_,
    new_new_n391_, new_new_n392_, new_new_n393_, new_new_n394_,
    new_new_n395_, new_new_n396_, new_new_n397_, new_new_n399_,
    new_new_n400_, new_new_n401_, new_new_n402_, new_new_n403_,
    new_new_n404_, new_new_n405_, new_new_n406_, new_new_n407_,
    new_new_n408_, new_new_n409_, new_new_n410_, new_new_n411_,
    new_new_n412_, new_new_n413_, new_new_n414_, new_new_n415_,
    new_new_n416_, new_new_n417_, new_new_n418_, new_new_n419_,
    new_new_n420_, new_new_n421_, new_new_n422_, new_new_n423_,
    new_new_n424_, new_new_n425_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n505_, new_new_n506_, new_new_n507_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  OAI210     g027(.A0(new_new_n49_), .A1(i_3_), .B0(new_new_n47_), .Y(new_new_n50_));
  NO2        g028(.A(new_new_n50_), .B(new_new_n46_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NA2        g030(.A(new_new_n51_), .B(new_new_n45_), .Y(new_new_n53_));
  NO2        g031(.A(i_1_), .B(i_6_), .Y(new_new_n54_));
  NAi21      g032(.An(i_2_), .B(i_7_), .Y(new_new_n55_));
  INV        g033(.A(i_1_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n56_), .B(i_6_), .Y(new_new_n57_));
  NA3        g035(.A(new_new_n57_), .B(new_new_n55_), .C(new_new_n31_), .Y(new_new_n58_));
  NA2        g036(.A(i_1_), .B(i_10_), .Y(new_new_n59_));
  NO2        g037(.A(new_new_n59_), .B(i_6_), .Y(new_new_n60_));
  NAi21      g038(.An(new_new_n60_), .B(new_new_n58_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n49_), .B(i_2_), .Y(new_new_n62_));
  AOI210     g040(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(i_1_), .B(i_6_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(new_new_n25_), .Y(new_new_n65_));
  INV        g043(.A(i_0_), .Y(new_new_n66_));
  NAi21      g044(.An(i_5_), .B(i_10_), .Y(new_new_n67_));
  NA2        g045(.A(i_5_), .B(i_9_), .Y(new_new_n68_));
  AOI210     g046(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n66_), .Y(new_new_n69_));
  NO2        g047(.A(new_new_n69_), .B(new_new_n65_), .Y(new_new_n70_));
  OAI210     g048(.A0(new_new_n63_), .A1(new_new_n62_), .B0(new_new_n70_), .Y(new_new_n71_));
  OAI210     g049(.A0(new_new_n71_), .A1(new_new_n61_), .B0(i_0_), .Y(new_new_n72_));
  NA2        g050(.A(i_12_), .B(i_5_), .Y(new_new_n73_));
  NO2        g051(.A(i_3_), .B(i_9_), .Y(new_new_n74_));
  NO2        g052(.A(i_3_), .B(i_7_), .Y(new_new_n75_));
  NO2        g053(.A(new_new_n74_), .B(new_new_n56_), .Y(new_new_n76_));
  INV        g054(.A(i_6_), .Y(new_new_n77_));
  NO2        g055(.A(i_2_), .B(i_7_), .Y(new_new_n78_));
  INV        g056(.A(new_new_n78_), .Y(new_new_n79_));
  NA2        g057(.A(new_new_n76_), .B(new_new_n79_), .Y(new_new_n80_));
  NAi21      g058(.An(i_6_), .B(i_10_), .Y(new_new_n81_));
  NA2        g059(.A(i_6_), .B(i_9_), .Y(new_new_n82_));
  AOI210     g060(.A0(new_new_n82_), .A1(new_new_n81_), .B0(new_new_n56_), .Y(new_new_n83_));
  NA2        g061(.A(i_2_), .B(i_6_), .Y(new_new_n84_));
  INV        g062(.A(new_new_n83_), .Y(new_new_n85_));
  AOI210     g063(.A0(new_new_n85_), .A1(new_new_n80_), .B0(new_new_n73_), .Y(new_new_n86_));
  AN3        g064(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n87_));
  NAi21      g065(.An(i_6_), .B(i_11_), .Y(new_new_n88_));
  NO2        g066(.A(i_5_), .B(i_8_), .Y(new_new_n89_));
  NOi21      g067(.An(new_new_n89_), .B(new_new_n88_), .Y(new_new_n90_));
  AOI220     g068(.A0(new_new_n90_), .A1(new_new_n55_), .B0(new_new_n87_), .B1(new_new_n32_), .Y(new_new_n91_));
  INV        g069(.A(i_7_), .Y(new_new_n92_));
  NA2        g070(.A(new_new_n46_), .B(new_new_n92_), .Y(new_new_n93_));
  NO2        g071(.A(i_0_), .B(i_5_), .Y(new_new_n94_));
  NO2        g072(.A(new_new_n94_), .B(new_new_n77_), .Y(new_new_n95_));
  NA2        g073(.A(i_12_), .B(i_3_), .Y(new_new_n96_));
  INV        g074(.A(new_new_n96_), .Y(new_new_n97_));
  NA3        g075(.A(new_new_n97_), .B(new_new_n95_), .C(new_new_n93_), .Y(new_new_n98_));
  NAi21      g076(.An(i_7_), .B(i_11_), .Y(new_new_n99_));
  AN2        g077(.A(i_2_), .B(i_10_), .Y(new_new_n100_));
  NO2        g078(.A(new_new_n100_), .B(i_7_), .Y(new_new_n101_));
  OR2        g079(.A(new_new_n73_), .B(new_new_n54_), .Y(new_new_n102_));
  NO2        g080(.A(i_8_), .B(new_new_n92_), .Y(new_new_n103_));
  NO3        g081(.A(new_new_n103_), .B(new_new_n102_), .C(new_new_n101_), .Y(new_new_n104_));
  NA2        g082(.A(i_12_), .B(i_7_), .Y(new_new_n105_));
  NA2        g083(.A(i_11_), .B(i_12_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n507_), .B(new_new_n104_), .Y(new_new_n107_));
  NA3        g085(.A(new_new_n107_), .B(new_new_n98_), .C(new_new_n91_), .Y(new_new_n108_));
  NOi21      g086(.An(i_1_), .B(i_5_), .Y(new_new_n109_));
  NA2        g087(.A(new_new_n109_), .B(i_11_), .Y(new_new_n110_));
  NA2        g088(.A(new_new_n92_), .B(new_new_n37_), .Y(new_new_n111_));
  NA2        g089(.A(i_7_), .B(new_new_n25_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n112_), .B(new_new_n111_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n113_), .B(new_new_n46_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n82_), .B(new_new_n81_), .Y(new_new_n115_));
  NAi21      g093(.An(i_3_), .B(i_8_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(new_new_n55_), .Y(new_new_n117_));
  NOi31      g095(.An(new_new_n117_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n118_));
  NO2        g096(.A(i_1_), .B(new_new_n77_), .Y(new_new_n119_));
  NO2        g097(.A(i_6_), .B(i_5_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(i_3_), .Y(new_new_n121_));
  OAI220     g099(.A0(new_new_n121_), .A1(new_new_n99_), .B0(new_new_n118_), .B1(new_new_n110_), .Y(new_new_n122_));
  NO3        g100(.A(new_new_n122_), .B(new_new_n108_), .C(new_new_n86_), .Y(new_new_n123_));
  NA3        g101(.A(new_new_n123_), .B(new_new_n72_), .C(new_new_n53_), .Y(ori2));
  NO2        g102(.A(new_new_n56_), .B(new_new_n37_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n505_), .B(new_new_n125_), .Y(new_new_n126_));
  NA4        g104(.A(new_new_n126_), .B(new_new_n70_), .C(new_new_n62_), .D(new_new_n30_), .Y(ori0));
  NO2        g105(.A(i_0_), .B(i_1_), .Y(new_new_n128_));
  NA2        g106(.A(i_2_), .B(i_3_), .Y(new_new_n129_));
  NO2        g107(.A(new_new_n129_), .B(i_4_), .Y(new_new_n130_));
  NA2        g108(.A(i_1_), .B(i_5_), .Y(new_new_n131_));
  OR2        g109(.A(i_0_), .B(i_1_), .Y(new_new_n132_));
  NO3        g110(.A(new_new_n132_), .B(new_new_n73_), .C(i_13_), .Y(new_new_n133_));
  NAi32      g111(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n134_));
  NAi21      g112(.An(new_new_n134_), .B(new_new_n133_), .Y(new_new_n135_));
  NOi21      g113(.An(i_4_), .B(i_10_), .Y(new_new_n136_));
  NOi21      g114(.An(i_4_), .B(i_9_), .Y(new_new_n137_));
  NOi21      g115(.An(i_11_), .B(i_13_), .Y(new_new_n138_));
  NA2        g116(.A(new_new_n138_), .B(new_new_n137_), .Y(new_new_n139_));
  NO2        g117(.A(new_new_n66_), .B(new_new_n56_), .Y(new_new_n140_));
  NO2        g118(.A(new_new_n66_), .B(i_5_), .Y(new_new_n141_));
  NO2        g119(.A(i_2_), .B(i_1_), .Y(new_new_n142_));
  NAi21      g120(.An(i_4_), .B(i_12_), .Y(new_new_n143_));
  INV        g121(.A(i_8_), .Y(new_new_n144_));
  NO2        g122(.A(i_3_), .B(i_8_), .Y(new_new_n145_));
  NO3        g123(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n146_));
  NO2        g124(.A(new_new_n94_), .B(new_new_n54_), .Y(new_new_n147_));
  NO2        g125(.A(i_13_), .B(i_9_), .Y(new_new_n148_));
  NAi21      g126(.An(i_12_), .B(i_3_), .Y(new_new_n149_));
  NO2        g127(.A(new_new_n44_), .B(i_5_), .Y(new_new_n150_));
  NA2        g128(.A(i_0_), .B(i_5_), .Y(new_new_n151_));
  INV        g129(.A(i_13_), .Y(new_new_n152_));
  NO2        g130(.A(i_12_), .B(new_new_n152_), .Y(new_new_n153_));
  NO2        g131(.A(i_12_), .B(new_new_n37_), .Y(new_new_n154_));
  OR2        g132(.A(i_8_), .B(i_7_), .Y(new_new_n155_));
  INV        g133(.A(i_12_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n44_), .B(new_new_n156_), .Y(new_new_n157_));
  NA2        g135(.A(i_2_), .B(i_1_), .Y(new_new_n158_));
  NO3        g136(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n159_));
  NAi21      g137(.An(i_4_), .B(i_3_), .Y(new_new_n160_));
  NO2        g138(.A(i_0_), .B(i_6_), .Y(new_new_n161_));
  NOi41      g139(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n162_));
  NO2        g140(.A(i_11_), .B(new_new_n152_), .Y(new_new_n163_));
  NOi21      g141(.An(i_1_), .B(i_6_), .Y(new_new_n164_));
  NAi21      g142(.An(i_3_), .B(i_7_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n156_), .B(i_9_), .Y(new_new_n166_));
  OR4        g144(.A(new_new_n166_), .B(new_new_n165_), .C(new_new_n164_), .D(new_new_n141_), .Y(new_new_n167_));
  NA2        g145(.A(new_new_n66_), .B(i_5_), .Y(new_new_n168_));
  NA2        g146(.A(i_3_), .B(i_9_), .Y(new_new_n169_));
  NAi21      g147(.An(i_7_), .B(i_10_), .Y(new_new_n170_));
  NO2        g148(.A(new_new_n170_), .B(new_new_n169_), .Y(new_new_n171_));
  NA3        g149(.A(new_new_n171_), .B(new_new_n168_), .C(new_new_n57_), .Y(new_new_n172_));
  NA2        g150(.A(new_new_n172_), .B(new_new_n167_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(new_new_n163_), .Y(new_new_n174_));
  NA2        g152(.A(i_12_), .B(i_6_), .Y(new_new_n175_));
  OR2        g153(.A(i_13_), .B(i_9_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n160_), .B(i_2_), .Y(new_new_n177_));
  NO2        g155(.A(new_new_n165_), .B(i_8_), .Y(new_new_n178_));
  NO3        g156(.A(i_12_), .B(new_new_n152_), .C(new_new_n37_), .Y(new_new_n179_));
  NO2        g157(.A(i_2_), .B(new_new_n92_), .Y(new_new_n180_));
  AN2        g158(.A(i_3_), .B(i_10_), .Y(new_new_n181_));
  NO2        g159(.A(i_5_), .B(new_new_n37_), .Y(new_new_n182_));
  NO2        g160(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n183_));
  NO2        g161(.A(i_2_), .B(i_3_), .Y(new_new_n184_));
  NO2        g162(.A(i_12_), .B(i_10_), .Y(new_new_n185_));
  NOi21      g163(.An(i_5_), .B(i_0_), .Y(new_new_n186_));
  NOi32      g164(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n187_));
  INV        g165(.A(new_new_n187_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n134_), .B(new_new_n132_), .Y(new_new_n189_));
  NOi32      g167(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n190_));
  NO2        g168(.A(i_1_), .B(new_new_n92_), .Y(new_new_n191_));
  NAi21      g169(.An(i_3_), .B(i_4_), .Y(new_new_n192_));
  NO2        g170(.A(new_new_n192_), .B(i_9_), .Y(new_new_n193_));
  AN2        g171(.A(i_6_), .B(i_7_), .Y(new_new_n194_));
  OAI210     g172(.A0(new_new_n194_), .A1(new_new_n191_), .B0(new_new_n193_), .Y(new_new_n195_));
  NO2        g173(.A(new_new_n192_), .B(i_10_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n195_), .B(new_new_n141_), .Y(new_new_n197_));
  AOI210     g175(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n198_));
  OAI210     g176(.A0(new_new_n198_), .A1(new_new_n142_), .B0(new_new_n196_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n199_), .B(i_5_), .Y(new_new_n200_));
  NO3        g178(.A(new_new_n200_), .B(new_new_n197_), .C(new_new_n189_), .Y(new_new_n201_));
  NO2        g179(.A(new_new_n201_), .B(new_new_n188_), .Y(new_new_n202_));
  AN2        g180(.A(i_12_), .B(i_5_), .Y(new_new_n203_));
  NO2        g181(.A(i_11_), .B(i_6_), .Y(new_new_n204_));
  NO2        g182(.A(i_5_), .B(i_10_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n206_));
  NO3        g184(.A(new_new_n77_), .B(new_new_n47_), .C(i_9_), .Y(new_new_n207_));
  NO2        g185(.A(i_0_), .B(i_11_), .Y(new_new_n208_));
  NOi21      g186(.An(i_2_), .B(i_12_), .Y(new_new_n209_));
  NAi21      g187(.An(i_9_), .B(i_4_), .Y(new_new_n210_));
  OR2        g188(.A(i_13_), .B(i_10_), .Y(new_new_n211_));
  NO3        g189(.A(new_new_n211_), .B(new_new_n106_), .C(new_new_n210_), .Y(new_new_n212_));
  NO2        g190(.A(new_new_n92_), .B(new_new_n25_), .Y(new_new_n213_));
  INV        g191(.A(new_new_n202_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n66_), .B(i_13_), .Y(new_new_n215_));
  NO2        g193(.A(i_10_), .B(i_9_), .Y(new_new_n216_));
  NAi21      g194(.An(i_12_), .B(i_8_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n217_), .B(i_3_), .Y(new_new_n218_));
  NO3        g196(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n219_));
  NA2        g197(.A(new_new_n175_), .B(new_new_n88_), .Y(new_new_n220_));
  NA2        g198(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n221_));
  NA2        g199(.A(i_8_), .B(i_9_), .Y(new_new_n222_));
  NO2        g200(.A(i_7_), .B(i_2_), .Y(new_new_n223_));
  OR2        g201(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n179_), .B(new_new_n147_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  NA2        g204(.A(new_new_n163_), .B(new_new_n182_), .Y(new_new_n227_));
  NO3        g205(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n228_));
  INV        g206(.A(new_new_n228_), .Y(new_new_n229_));
  NO2        g207(.A(new_new_n229_), .B(new_new_n227_), .Y(new_new_n230_));
  NO2        g208(.A(new_new_n230_), .B(new_new_n226_), .Y(new_new_n231_));
  NO2        g209(.A(i_11_), .B(i_1_), .Y(new_new_n232_));
  NOi21      g210(.An(i_2_), .B(i_7_), .Y(new_new_n233_));
  NA3        g211(.A(new_new_n162_), .B(new_new_n138_), .C(new_new_n120_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n132_), .B(i_3_), .Y(new_new_n236_));
  NAi31      g214(.An(new_new_n235_), .B(new_new_n236_), .C(new_new_n153_), .Y(new_new_n237_));
  NA3        g215(.A(new_new_n206_), .B(new_new_n140_), .C(new_new_n130_), .Y(new_new_n238_));
  NA3        g216(.A(new_new_n238_), .B(new_new_n237_), .C(new_new_n234_), .Y(new_new_n239_));
  INV        g217(.A(new_new_n239_), .Y(new_new_n240_));
  NA2        g218(.A(new_new_n219_), .B(new_new_n203_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n228_), .B(new_new_n205_), .Y(new_new_n242_));
  NA2        g220(.A(new_new_n240_), .B(new_new_n231_), .Y(new_new_n243_));
  NA2        g221(.A(new_new_n203_), .B(new_new_n152_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n194_), .B(new_new_n190_), .Y(new_new_n245_));
  OR2        g223(.A(new_new_n244_), .B(new_new_n245_), .Y(new_new_n246_));
  NO2        g224(.A(new_new_n36_), .B(i_8_), .Y(new_new_n247_));
  AOI210     g225(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n212_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n248_), .B(new_new_n246_), .Y(new_new_n249_));
  NA3        g227(.A(new_new_n151_), .B(new_new_n64_), .C(new_new_n44_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n179_), .B(new_new_n75_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n250_), .B(new_new_n251_), .Y(new_new_n252_));
  NO3        g230(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n253_));
  NO2        g231(.A(new_new_n211_), .B(i_1_), .Y(new_new_n254_));
  NOi31      g232(.An(new_new_n254_), .B(new_new_n220_), .C(new_new_n66_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n77_), .B(new_new_n25_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n105_), .B(new_new_n23_), .Y(new_new_n257_));
  NO2        g235(.A(i_12_), .B(new_new_n77_), .Y(new_new_n258_));
  NO3        g236(.A(new_new_n252_), .B(new_new_n249_), .C(new_new_n243_), .Y(new_new_n259_));
  NA3        g237(.A(new_new_n259_), .B(new_new_n214_), .C(new_new_n174_), .Y(ori7));
  NO2        g238(.A(new_new_n84_), .B(new_new_n52_), .Y(new_new_n261_));
  NA2        g239(.A(i_11_), .B(new_new_n144_), .Y(new_new_n262_));
  NA3        g240(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n156_), .B(i_4_), .Y(new_new_n264_));
  NA2        g242(.A(new_new_n264_), .B(i_8_), .Y(new_new_n265_));
  NO2        g243(.A(new_new_n96_), .B(new_new_n263_), .Y(new_new_n266_));
  NA2        g244(.A(i_2_), .B(new_new_n77_), .Y(new_new_n267_));
  OAI210     g245(.A0(new_new_n78_), .A1(new_new_n145_), .B0(new_new_n146_), .Y(new_new_n268_));
  NO2        g246(.A(i_7_), .B(new_new_n37_), .Y(new_new_n269_));
  NA2        g247(.A(i_4_), .B(i_8_), .Y(new_new_n270_));
  AOI210     g248(.A0(new_new_n270_), .A1(new_new_n181_), .B0(new_new_n269_), .Y(new_new_n271_));
  OAI220     g249(.A0(new_new_n271_), .A1(new_new_n267_), .B0(new_new_n268_), .B1(i_13_), .Y(new_new_n272_));
  NO3        g250(.A(new_new_n272_), .B(new_new_n266_), .C(new_new_n261_), .Y(new_new_n273_));
  AOI210     g251(.A0(new_new_n116_), .A1(new_new_n55_), .B0(i_10_), .Y(new_new_n274_));
  AOI210     g252(.A0(new_new_n274_), .A1(new_new_n156_), .B0(new_new_n136_), .Y(new_new_n275_));
  OR2        g253(.A(i_6_), .B(i_10_), .Y(new_new_n276_));
  OR3        g254(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n277_));
  OR2        g255(.A(new_new_n275_), .B(new_new_n176_), .Y(new_new_n278_));
  AOI210     g256(.A0(new_new_n278_), .A1(new_new_n273_), .B0(new_new_n56_), .Y(new_new_n279_));
  NOi21      g257(.An(i_11_), .B(i_7_), .Y(new_new_n280_));
  AO210      g258(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n281_), .B(new_new_n280_), .Y(new_new_n282_));
  NA2        g260(.A(new_new_n282_), .B(new_new_n148_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n283_), .B(new_new_n56_), .Y(new_new_n284_));
  NA2        g262(.A(new_new_n153_), .B(new_new_n56_), .Y(new_new_n285_));
  NO2        g263(.A(i_1_), .B(i_12_), .Y(new_new_n286_));
  INV        g264(.A(new_new_n285_), .Y(new_new_n287_));
  OAI210     g265(.A0(new_new_n287_), .A1(new_new_n284_), .B0(i_6_), .Y(new_new_n288_));
  NO2        g266(.A(i_6_), .B(i_11_), .Y(new_new_n289_));
  INV        g267(.A(new_new_n221_), .Y(new_new_n290_));
  NO3        g268(.A(new_new_n276_), .B(new_new_n155_), .C(new_new_n23_), .Y(new_new_n291_));
  AOI210     g269(.A0(i_1_), .A1(new_new_n171_), .B0(new_new_n291_), .Y(new_new_n292_));
  NO2        g270(.A(new_new_n292_), .B(new_new_n44_), .Y(new_new_n293_));
  INV        g271(.A(i_2_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n125_), .B(i_9_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n46_), .B(i_1_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n295_), .B(new_new_n294_), .Y(new_new_n297_));
  AOI210     g275(.A0(new_new_n232_), .A1(new_new_n213_), .B0(new_new_n159_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n298_), .B(new_new_n267_), .Y(new_new_n299_));
  NO2        g277(.A(i_11_), .B(new_new_n37_), .Y(new_new_n300_));
  OR2        g278(.A(new_new_n299_), .B(new_new_n297_), .Y(new_new_n301_));
  NO3        g279(.A(new_new_n301_), .B(new_new_n293_), .C(new_new_n290_), .Y(new_new_n302_));
  NO2        g280(.A(new_new_n156_), .B(new_new_n92_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n303_), .B(new_new_n280_), .Y(new_new_n304_));
  NA2        g282(.A(new_new_n304_), .B(i_1_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n305_), .B(new_new_n277_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n210_), .B(new_new_n77_), .Y(new_new_n307_));
  NA2        g285(.A(new_new_n306_), .B(new_new_n46_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n155_), .B(new_new_n44_), .Y(new_new_n309_));
  NO3        g287(.A(new_new_n309_), .B(new_new_n183_), .C(new_new_n157_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n106_), .B(new_new_n37_), .Y(new_new_n311_));
  NO2        g289(.A(new_new_n311_), .B(i_6_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n77_), .B(i_9_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n313_), .B(new_new_n56_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n314_), .B(new_new_n286_), .Y(new_new_n315_));
  NO4        g293(.A(new_new_n315_), .B(new_new_n312_), .C(new_new_n310_), .D(i_4_), .Y(new_new_n316_));
  INV        g294(.A(new_new_n316_), .Y(new_new_n317_));
  NA4        g295(.A(new_new_n317_), .B(new_new_n308_), .C(new_new_n302_), .D(new_new_n288_), .Y(new_new_n318_));
  AOI210     g296(.A0(new_new_n175_), .A1(new_new_n88_), .B0(i_1_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n192_), .B(i_2_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n320_), .B(new_new_n319_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n321_), .B(i_13_), .Y(new_new_n322_));
  NO2        g300(.A(new_new_n52_), .B(i_12_), .Y(new_new_n323_));
  INV        g301(.A(new_new_n323_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n233_), .B(new_new_n24_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n325_), .B(new_new_n307_), .Y(new_new_n326_));
  OAI220     g304(.A0(new_new_n326_), .A1(new_new_n41_), .B0(new_new_n324_), .B1(new_new_n84_), .Y(new_new_n327_));
  INV        g305(.A(new_new_n327_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n204_), .B(new_new_n296_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n329_), .B(new_new_n160_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n115_), .B(i_13_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n331_), .B(new_new_n319_), .Y(new_new_n332_));
  NA2        g310(.A(new_new_n26_), .B(new_new_n144_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n83_), .B(new_new_n93_), .Y(new_new_n334_));
  NO2        g312(.A(new_new_n334_), .B(new_new_n265_), .Y(new_new_n335_));
  NO3        g313(.A(new_new_n335_), .B(new_new_n332_), .C(new_new_n330_), .Y(new_new_n336_));
  OR2        g314(.A(i_11_), .B(i_6_), .Y(new_new_n337_));
  NA3        g315(.A(new_new_n264_), .B(new_new_n333_), .C(i_7_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n338_), .B(new_new_n337_), .Y(new_new_n339_));
  NA3        g317(.A(new_new_n209_), .B(new_new_n269_), .C(new_new_n88_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n289_), .B(i_13_), .Y(new_new_n341_));
  NAi21      g319(.An(i_11_), .B(i_12_), .Y(new_new_n342_));
  NOi41      g320(.An(new_new_n101_), .B(new_new_n342_), .C(i_13_), .D(new_new_n77_), .Y(new_new_n343_));
  INV        g321(.A(new_new_n343_), .Y(new_new_n344_));
  NA3        g322(.A(new_new_n344_), .B(new_new_n341_), .C(new_new_n340_), .Y(new_new_n345_));
  OAI210     g323(.A0(new_new_n345_), .A1(new_new_n339_), .B0(new_new_n56_), .Y(new_new_n346_));
  NO2        g324(.A(i_2_), .B(i_12_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n191_), .B(new_new_n347_), .Y(new_new_n348_));
  INV        g326(.A(new_new_n348_), .Y(new_new_n349_));
  NA3        g327(.A(new_new_n349_), .B(new_new_n45_), .C(new_new_n152_), .Y(new_new_n350_));
  NA4        g328(.A(new_new_n350_), .B(new_new_n346_), .C(new_new_n336_), .D(new_new_n328_), .Y(new_new_n351_));
  OR4        g329(.A(new_new_n351_), .B(new_new_n322_), .C(new_new_n318_), .D(new_new_n279_), .Y(ori5));
  NA2        g330(.A(new_new_n304_), .B(new_new_n177_), .Y(new_new_n353_));
  AN2        g331(.A(new_new_n24_), .B(i_10_), .Y(new_new_n354_));
  NA3        g332(.A(new_new_n354_), .B(new_new_n347_), .C(new_new_n99_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n265_), .B(i_11_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n78_), .B(new_new_n356_), .Y(new_new_n357_));
  NA3        g335(.A(new_new_n357_), .B(new_new_n355_), .C(new_new_n353_), .Y(new_new_n358_));
  NO3        g336(.A(i_11_), .B(new_new_n156_), .C(i_13_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n112_), .B(new_new_n23_), .Y(new_new_n360_));
  NA2        g338(.A(i_12_), .B(i_8_), .Y(new_new_n361_));
  OAI210     g339(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n361_), .Y(new_new_n362_));
  INV        g340(.A(new_new_n216_), .Y(new_new_n363_));
  AOI220     g341(.A0(new_new_n184_), .A1(new_new_n257_), .B0(new_new_n362_), .B1(new_new_n360_), .Y(new_new_n364_));
  INV        g342(.A(new_new_n364_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n365_), .B(new_new_n358_), .Y(new_new_n366_));
  INV        g344(.A(new_new_n138_), .Y(new_new_n367_));
  INV        g345(.A(new_new_n162_), .Y(new_new_n368_));
  OAI210     g346(.A0(new_new_n320_), .A1(new_new_n218_), .B0(new_new_n101_), .Y(new_new_n369_));
  AOI210     g347(.A0(new_new_n369_), .A1(new_new_n368_), .B0(new_new_n367_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n222_), .B(new_new_n26_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n371_), .B(new_new_n213_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n372_), .B(i_2_), .Y(new_new_n373_));
  INV        g351(.A(new_new_n373_), .Y(new_new_n374_));
  AOI210     g352(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n211_), .Y(new_new_n375_));
  AOI210     g353(.A0(new_new_n375_), .A1(new_new_n374_), .B0(new_new_n370_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n143_), .B(new_new_n113_), .Y(new_new_n377_));
  OAI210     g355(.A0(new_new_n377_), .A1(new_new_n360_), .B0(i_2_), .Y(new_new_n378_));
  INV        g356(.A(new_new_n139_), .Y(new_new_n379_));
  NO3        g357(.A(new_new_n281_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n380_));
  AOI210     g358(.A0(new_new_n379_), .A1(new_new_n78_), .B0(new_new_n380_), .Y(new_new_n381_));
  AOI210     g359(.A0(new_new_n381_), .A1(new_new_n378_), .B0(new_new_n144_), .Y(new_new_n382_));
  OA210      g360(.A0(new_new_n282_), .A1(new_new_n114_), .B0(i_13_), .Y(new_new_n383_));
  AOI210     g361(.A0(new_new_n149_), .A1(new_new_n129_), .B0(new_new_n247_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n384_), .B(new_new_n213_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n93_), .B(new_new_n44_), .Y(new_new_n386_));
  INV        g364(.A(new_new_n180_), .Y(new_new_n387_));
  NA4        g365(.A(new_new_n387_), .B(new_new_n181_), .C(new_new_n112_), .D(new_new_n42_), .Y(new_new_n388_));
  OAI210     g366(.A0(new_new_n388_), .A1(new_new_n386_), .B0(new_new_n385_), .Y(new_new_n389_));
  NO3        g367(.A(new_new_n389_), .B(new_new_n383_), .C(new_new_n382_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n257_), .B(new_new_n28_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n359_), .B(new_new_n178_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n392_), .B(new_new_n391_), .Y(new_new_n393_));
  NO2        g371(.A(new_new_n55_), .B(i_12_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n394_), .B(new_new_n114_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n395_), .B(new_new_n262_), .Y(new_new_n396_));
  AOI220     g374(.A0(new_new_n396_), .A1(new_new_n36_), .B0(new_new_n393_), .B1(new_new_n46_), .Y(new_new_n397_));
  NA4        g375(.A(new_new_n397_), .B(new_new_n390_), .C(new_new_n376_), .D(new_new_n366_), .Y(ori6));
  OR2        g376(.A(new_new_n506_), .B(i_12_), .Y(new_new_n399_));
  NA2        g377(.A(new_new_n258_), .B(new_new_n56_), .Y(new_new_n400_));
  INV        g378(.A(new_new_n400_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n401_), .B(new_new_n66_), .Y(new_new_n402_));
  INV        g380(.A(new_new_n185_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n68_), .B(new_new_n119_), .Y(new_new_n404_));
  INV        g382(.A(new_new_n112_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n405_), .B(new_new_n46_), .Y(new_new_n406_));
  AOI210     g384(.A0(new_new_n406_), .A1(new_new_n404_), .B0(new_new_n403_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n164_), .B(i_9_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n408_), .B(new_new_n394_), .Y(new_new_n409_));
  AOI210     g387(.A0(new_new_n409_), .A1(new_new_n245_), .B0(new_new_n141_), .Y(new_new_n410_));
  NAi32      g388(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n337_), .B(new_new_n411_), .Y(new_new_n412_));
  OR3        g390(.A(new_new_n412_), .B(new_new_n410_), .C(new_new_n407_), .Y(new_new_n413_));
  BUFFER     g391(.A(new_new_n282_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n414_), .B(new_new_n128_), .Y(new_new_n415_));
  AO210      g393(.A0(new_new_n242_), .A1(new_new_n363_), .B0(new_new_n36_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n416_), .B(new_new_n415_), .Y(new_new_n417_));
  NO2        g395(.A(i_6_), .B(i_11_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n418_), .B(new_new_n253_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n207_), .B(new_new_n63_), .Y(new_new_n420_));
  NA3        g398(.A(new_new_n420_), .B(new_new_n419_), .C(new_new_n268_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n218_), .B(new_new_n216_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n102_), .B(new_new_n208_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n423_), .B(new_new_n422_), .Y(new_new_n424_));
  NO4        g402(.A(new_new_n424_), .B(new_new_n421_), .C(new_new_n417_), .D(new_new_n413_), .Y(new_new_n425_));
  NA4        g403(.A(new_new_n425_), .B(new_new_n402_), .C(new_new_n399_), .D(new_new_n201_), .Y(ori3));
  NA2        g404(.A(i_12_), .B(i_10_), .Y(new_new_n427_));
  NO2        g405(.A(i_11_), .B(new_new_n156_), .Y(new_new_n428_));
  NA2        g406(.A(new_new_n268_), .B(new_new_n195_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n429_), .B(new_new_n40_), .Y(new_new_n430_));
  NOi21      g408(.An(new_new_n87_), .B(new_new_n372_), .Y(new_new_n431_));
  INV        g409(.A(new_new_n431_), .Y(new_new_n432_));
  AOI210     g410(.A0(new_new_n432_), .A1(new_new_n430_), .B0(new_new_n47_), .Y(new_new_n433_));
  NO4        g411(.A(new_new_n198_), .B(new_new_n203_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n141_), .B(i_10_), .Y(new_new_n435_));
  NOi21      g413(.An(new_new_n435_), .B(new_new_n434_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n56_), .Y(new_new_n437_));
  NOi21      g415(.An(i_5_), .B(i_9_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n438_), .B(new_new_n215_), .Y(new_new_n439_));
  BUFFER     g417(.A(new_new_n175_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n440_), .B(new_new_n232_), .Y(new_new_n441_));
  NO2        g419(.A(new_new_n441_), .B(new_new_n439_), .Y(new_new_n442_));
  NO3        g420(.A(new_new_n442_), .B(new_new_n437_), .C(new_new_n433_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n256_), .B(i_0_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n359_), .B(new_new_n186_), .Y(new_new_n445_));
  INV        g423(.A(new_new_n54_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n446_), .B(new_new_n445_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n166_), .B(new_new_n131_), .Y(new_new_n448_));
  NA2        g426(.A(i_0_), .B(i_10_), .Y(new_new_n449_));
  AN2        g427(.A(new_new_n448_), .B(i_6_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n450_), .B(new_new_n447_), .Y(new_new_n451_));
  INV        g429(.A(new_new_n451_), .Y(new_new_n452_));
  NA2        g430(.A(i_11_), .B(i_9_), .Y(new_new_n453_));
  NO3        g431(.A(i_12_), .B(new_new_n453_), .C(new_new_n267_), .Y(new_new_n454_));
  AN2        g432(.A(new_new_n454_), .B(i_5_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n206_), .B(new_new_n140_), .Y(new_new_n456_));
  NA2        g434(.A(new_new_n456_), .B(new_new_n135_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n453_), .B(new_new_n66_), .Y(new_new_n458_));
  NO2        g436(.A(new_new_n457_), .B(new_new_n455_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n300_), .B(new_new_n109_), .Y(new_new_n460_));
  NO2        g438(.A(i_6_), .B(new_new_n460_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n138_), .B(new_new_n94_), .Y(new_new_n462_));
  INV        g440(.A(new_new_n461_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n463_), .B(new_new_n459_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n427_), .B(new_new_n184_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n465_), .B(new_new_n458_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n246_), .B(new_new_n466_), .Y(new_new_n467_));
  NO3        g445(.A(new_new_n467_), .B(new_new_n464_), .C(new_new_n452_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n400_), .B(new_new_n462_), .Y(new_new_n469_));
  INV        g447(.A(new_new_n469_), .Y(new_new_n470_));
  NA2        g448(.A(new_new_n161_), .B(new_new_n154_), .Y(new_new_n471_));
  AOI210     g449(.A0(new_new_n471_), .A1(new_new_n444_), .B0(new_new_n131_), .Y(new_new_n472_));
  INV        g450(.A(new_new_n472_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n473_), .B(new_new_n470_), .Y(new_new_n474_));
  NO3        g452(.A(new_new_n449_), .B(new_new_n438_), .C(new_new_n143_), .Y(new_new_n475_));
  AOI220     g453(.A0(new_new_n475_), .A1(i_11_), .B0(new_new_n255_), .B1(new_new_n68_), .Y(new_new_n476_));
  NO3        g454(.A(new_new_n150_), .B(new_new_n203_), .C(i_0_), .Y(new_new_n477_));
  OAI210     g455(.A0(new_new_n477_), .A1(new_new_n69_), .B0(i_13_), .Y(new_new_n478_));
  NA2        g456(.A(new_new_n478_), .B(new_new_n476_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n241_), .B(new_new_n234_), .Y(new_new_n480_));
  INV        g458(.A(new_new_n480_), .Y(new_new_n481_));
  NA3        g459(.A(new_new_n205_), .B(new_new_n138_), .C(new_new_n137_), .Y(new_new_n482_));
  INV        g460(.A(new_new_n482_), .Y(new_new_n483_));
  NO3        g461(.A(new_new_n453_), .B(new_new_n151_), .C(new_new_n143_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n484_), .B(new_new_n483_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n485_), .B(new_new_n481_), .Y(new_new_n486_));
  NO2        g464(.A(new_new_n77_), .B(i_5_), .Y(new_new_n487_));
  NA3        g465(.A(new_new_n428_), .B(new_new_n100_), .C(new_new_n112_), .Y(new_new_n488_));
  INV        g466(.A(new_new_n488_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n489_), .B(new_new_n487_), .Y(new_new_n490_));
  NAi21      g468(.An(new_new_n159_), .B(new_new_n160_), .Y(new_new_n491_));
  NO4        g469(.A(new_new_n158_), .B(new_new_n150_), .C(i_0_), .D(i_12_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n492_), .B(new_new_n491_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n493_), .B(new_new_n490_), .Y(new_new_n494_));
  NO4        g472(.A(new_new_n494_), .B(new_new_n486_), .C(new_new_n479_), .D(new_new_n474_), .Y(new_new_n495_));
  INV        g473(.A(new_new_n275_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n496_), .B(new_new_n148_), .Y(new_new_n497_));
  NO2        g475(.A(new_new_n497_), .B(new_new_n66_), .Y(new_new_n498_));
  INV        g476(.A(new_new_n200_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n499_), .B(new_new_n367_), .Y(new_new_n500_));
  NO2        g478(.A(new_new_n500_), .B(new_new_n498_), .Y(new_new_n501_));
  NA4        g479(.A(new_new_n501_), .B(new_new_n495_), .C(new_new_n468_), .D(new_new_n443_), .Y(ori4));
  INV        g480(.A(i_6_), .Y(new_new_n505_));
  INV        g481(.A(new_new_n186_), .Y(new_new_n506_));
  INV        g482(.A(new_new_n106_), .Y(new_new_n507_));
endmodule


