//Benchmark atmr_9sym_175_0.0625

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n152_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  INV        o002(.A(i_5_), .Y(ori_ori_n13_));
  NOi21      o003(.An(i_3_), .B(i_7_), .Y(ori_ori_n14_));
  NA3        o004(.A(ori_ori_n14_), .B(i_0_), .C(ori_ori_n13_), .Y(ori_ori_n15_));
  INV        o005(.A(i_0_), .Y(ori_ori_n16_));
  NOi21      o006(.An(i_1_), .B(i_3_), .Y(ori_ori_n17_));
  NA3        o007(.A(ori_ori_n17_), .B(ori_ori_n16_), .C(i_2_), .Y(ori_ori_n18_));
  AOI210     o008(.A0(ori_ori_n18_), .A1(ori_ori_n15_), .B0(ori_ori_n149_), .Y(ori_ori_n19_));
  INV        o009(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o010(.A(i_0_), .B(ori_ori_n20_), .Y(ori_ori_n21_));
  INV        o011(.A(i_7_), .Y(ori_ori_n22_));
  NA2        o012(.A(i_6_), .B(i_5_), .Y(ori_ori_n23_));
  NOi21      o013(.An(i_8_), .B(i_6_), .Y(ori_ori_n24_));
  AOI220     o014(.A0(i_1_), .A1(i_2_), .B0(ori_ori_n24_), .B1(i_5_), .Y(ori_ori_n25_));
  AOI210     o015(.A0(ori_ori_n25_), .A1(ori_ori_n23_), .B0(ori_ori_n21_), .Y(ori_ori_n26_));
  AOI210     o016(.A0(ori_ori_n26_), .A1(ori_ori_n11_), .B0(ori_ori_n19_), .Y(ori_ori_n27_));
  NA2        o017(.A(ori_ori_n16_), .B(i_5_), .Y(ori_ori_n28_));
  NO2        o018(.A(i_2_), .B(i_4_), .Y(ori_ori_n29_));
  NA3        o019(.A(ori_ori_n29_), .B(i_6_), .C(i_8_), .Y(ori_ori_n30_));
  AOI210     o020(.A0(ori_ori_n28_), .A1(ori_ori_n151_), .B0(ori_ori_n30_), .Y(ori_ori_n31_));
  INV        o021(.A(i_2_), .Y(ori_ori_n32_));
  NOi21      o022(.An(i_5_), .B(i_0_), .Y(ori_ori_n33_));
  NOi21      o023(.An(i_6_), .B(i_8_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_5_), .B(i_6_), .Y(ori_ori_n35_));
  AOI220     o025(.A0(ori_ori_n35_), .A1(i_7_), .B0(ori_ori_n34_), .B1(ori_ori_n33_), .Y(ori_ori_n36_));
  NO3        o026(.A(ori_ori_n36_), .B(ori_ori_n32_), .C(i_4_), .Y(ori_ori_n37_));
  NOi21      o027(.An(i_0_), .B(i_4_), .Y(ori_ori_n38_));
  NOi21      o028(.An(i_7_), .B(i_5_), .Y(ori_ori_n39_));
  AN2        o029(.A(ori_ori_n39_), .B(ori_ori_n38_), .Y(ori_ori_n40_));
  INV        o030(.A(i_1_), .Y(ori_ori_n41_));
  NOi21      o031(.An(i_3_), .B(i_0_), .Y(ori_ori_n42_));
  NA2        o032(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NO2        o033(.A(ori_ori_n23_), .B(ori_ori_n43_), .Y(ori_ori_n44_));
  NO4        o034(.A(ori_ori_n44_), .B(ori_ori_n40_), .C(ori_ori_n37_), .D(ori_ori_n31_), .Y(ori_ori_n45_));
  NOi21      o035(.An(i_4_), .B(i_0_), .Y(ori_ori_n46_));
  NO2        o036(.A(ori_ori_n24_), .B(ori_ori_n14_), .Y(ori_ori_n47_));
  NA2        o037(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n48_));
  NOi21      o038(.An(i_2_), .B(i_8_), .Y(ori_ori_n49_));
  NO2        o039(.A(ori_ori_n46_), .B(ori_ori_n38_), .Y(ori_ori_n50_));
  NO3        o040(.A(ori_ori_n50_), .B(ori_ori_n48_), .C(ori_ori_n47_), .Y(ori_ori_n51_));
  INV        o041(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NOi31      o042(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n53_));
  NA2        o043(.A(ori_ori_n53_), .B(i_0_), .Y(ori_ori_n54_));
  NOi21      o044(.An(i_4_), .B(i_3_), .Y(ori_ori_n55_));
  NOi21      o045(.An(i_1_), .B(i_4_), .Y(ori_ori_n56_));
  OAI210     o046(.A0(ori_ori_n56_), .A1(ori_ori_n55_), .B0(ori_ori_n49_), .Y(ori_ori_n57_));
  NA2        o047(.A(ori_ori_n57_), .B(ori_ori_n54_), .Y(ori_ori_n58_));
  AN2        o048(.A(i_8_), .B(i_7_), .Y(ori_ori_n59_));
  INV        o049(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  NOi21      o050(.An(i_8_), .B(i_7_), .Y(ori_ori_n61_));
  NA3        o051(.A(ori_ori_n61_), .B(ori_ori_n55_), .C(i_6_), .Y(ori_ori_n62_));
  OAI210     o052(.A0(ori_ori_n60_), .A1(ori_ori_n48_), .B0(ori_ori_n62_), .Y(ori_ori_n63_));
  AOI220     o053(.A0(ori_ori_n63_), .A1(ori_ori_n32_), .B0(ori_ori_n58_), .B1(ori_ori_n35_), .Y(ori_ori_n64_));
  NA4        o054(.A(ori_ori_n64_), .B(ori_ori_n52_), .C(ori_ori_n45_), .D(ori_ori_n27_), .Y(ori_ori_n65_));
  INV        o055(.A(i_7_), .Y(ori_ori_n66_));
  NO3        o056(.A(ori_ori_n66_), .B(ori_ori_n149_), .C(i_1_), .Y(ori_ori_n67_));
  NOi21      o057(.An(i_1_), .B(i_2_), .Y(ori_ori_n68_));
  NA2        o058(.A(ori_ori_n67_), .B(ori_ori_n13_), .Y(ori_ori_n69_));
  NA3        o059(.A(ori_ori_n61_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n70_));
  NA3        o060(.A(i_1_), .B(i_0_), .C(ori_ori_n13_), .Y(ori_ori_n71_));
  NA2        o061(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n72_));
  NA2        o062(.A(ori_ori_n17_), .B(i_6_), .Y(ori_ori_n73_));
  INV        o063(.A(ori_ori_n73_), .Y(ori_ori_n74_));
  INV        o064(.A(i_0_), .Y(ori_ori_n75_));
  AOI220     o065(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n72_), .B1(ori_ori_n55_), .Y(ori_ori_n76_));
  NA2        o066(.A(ori_ori_n76_), .B(ori_ori_n69_), .Y(ori_ori_n77_));
  NOi21      o067(.An(i_7_), .B(i_8_), .Y(ori_ori_n78_));
  NA2        o068(.A(ori_ori_n78_), .B(ori_ori_n68_), .Y(ori_ori_n79_));
  NA3        o069(.A(ori_ori_n24_), .B(i_2_), .C(ori_ori_n13_), .Y(ori_ori_n80_));
  NO2        o070(.A(i_3_), .B(ori_ori_n80_), .Y(ori_ori_n81_));
  NA2        o071(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n82_));
  NO2        o072(.A(ori_ori_n150_), .B(ori_ori_n82_), .Y(ori_ori_n83_));
  NO2        o073(.A(ori_ori_n83_), .B(ori_ori_n81_), .Y(ori_ori_n84_));
  NA3        o074(.A(ori_ori_n61_), .B(ori_ori_n32_), .C(i_3_), .Y(ori_ori_n85_));
  NA2        o075(.A(ori_ori_n41_), .B(i_6_), .Y(ori_ori_n86_));
  NO2        o076(.A(ori_ori_n86_), .B(ori_ori_n85_), .Y(ori_ori_n87_));
  NAi21      o077(.An(i_6_), .B(i_0_), .Y(ori_ori_n88_));
  NA2        o078(.A(ori_ori_n56_), .B(i_5_), .Y(ori_ori_n89_));
  NOi21      o079(.An(i_4_), .B(i_6_), .Y(ori_ori_n90_));
  NA3        o080(.A(i_5_), .B(ori_ori_n68_), .C(ori_ori_n90_), .Y(ori_ori_n91_));
  OAI210     o081(.A0(ori_ori_n89_), .A1(ori_ori_n88_), .B0(ori_ori_n91_), .Y(ori_ori_n92_));
  NA2        o082(.A(ori_ori_n68_), .B(ori_ori_n34_), .Y(ori_ori_n93_));
  NO2        o083(.A(ori_ori_n92_), .B(ori_ori_n87_), .Y(ori_ori_n94_));
  NOi21      o084(.An(i_6_), .B(i_1_), .Y(ori_ori_n95_));
  AOI220     o085(.A0(ori_ori_n95_), .A1(i_7_), .B0(ori_ori_n24_), .B1(i_5_), .Y(ori_ori_n96_));
  NOi21      o086(.An(ori_ori_n46_), .B(ori_ori_n96_), .Y(ori_ori_n97_));
  NA2        o087(.A(ori_ori_n61_), .B(ori_ori_n12_), .Y(ori_ori_n98_));
  NOi21      o088(.An(i_3_), .B(i_1_), .Y(ori_ori_n99_));
  NA2        o089(.A(ori_ori_n99_), .B(i_4_), .Y(ori_ori_n100_));
  NO2        o090(.A(ori_ori_n98_), .B(ori_ori_n100_), .Y(ori_ori_n101_));
  NOi31      o091(.An(ori_ori_n42_), .B(i_5_), .C(ori_ori_n32_), .Y(ori_ori_n102_));
  NO3        o092(.A(ori_ori_n102_), .B(ori_ori_n101_), .C(ori_ori_n97_), .Y(ori_ori_n103_));
  NA4        o093(.A(ori_ori_n103_), .B(ori_ori_n94_), .C(ori_ori_n84_), .D(ori_ori_n79_), .Y(ori_ori_n104_));
  NA2        o094(.A(ori_ori_n49_), .B(ori_ori_n14_), .Y(ori_ori_n105_));
  NOi31      o095(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n106_));
  NOi31      o096(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n107_));
  OAI210     o097(.A0(ori_ori_n107_), .A1(ori_ori_n106_), .B0(i_7_), .Y(ori_ori_n108_));
  NA3        o098(.A(ori_ori_n108_), .B(ori_ori_n105_), .C(ori_ori_n93_), .Y(ori_ori_n109_));
  NA2        o099(.A(ori_ori_n109_), .B(ori_ori_n38_), .Y(ori_ori_n110_));
  NO2        o100(.A(ori_ori_n70_), .B(ori_ori_n28_), .Y(ori_ori_n111_));
  NA3        o101(.A(ori_ori_n61_), .B(ori_ori_n53_), .C(i_6_), .Y(ori_ori_n112_));
  INV        o102(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  NOi21      o103(.An(i_0_), .B(i_2_), .Y(ori_ori_n114_));
  NA3        o104(.A(ori_ori_n114_), .B(i_7_), .C(ori_ori_n90_), .Y(ori_ori_n115_));
  NOi32      o105(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n116_));
  NA2        o106(.A(ori_ori_n116_), .B(ori_ori_n106_), .Y(ori_ori_n117_));
  NA3        o107(.A(ori_ori_n114_), .B(ori_ori_n55_), .C(ori_ori_n34_), .Y(ori_ori_n118_));
  NA3        o108(.A(ori_ori_n118_), .B(ori_ori_n117_), .C(ori_ori_n115_), .Y(ori_ori_n119_));
  NA3        o109(.A(ori_ori_n53_), .B(i_6_), .C(ori_ori_n13_), .Y(ori_ori_n120_));
  NA3        o110(.A(ori_ori_n56_), .B(ori_ori_n35_), .C(i_8_), .Y(ori_ori_n121_));
  NA3        o111(.A(ori_ori_n56_), .B(ori_ori_n42_), .C(ori_ori_n22_), .Y(ori_ori_n122_));
  NA3        o112(.A(ori_ori_n122_), .B(ori_ori_n121_), .C(ori_ori_n120_), .Y(ori_ori_n123_));
  NO4        o113(.A(ori_ori_n123_), .B(ori_ori_n119_), .C(ori_ori_n113_), .D(ori_ori_n111_), .Y(ori_ori_n124_));
  NA2        o114(.A(ori_ori_n59_), .B(ori_ori_n29_), .Y(ori_ori_n125_));
  AOI210     o115(.A0(ori_ori_n125_), .A1(ori_ori_n105_), .B0(ori_ori_n86_), .Y(ori_ori_n126_));
  NO4        o116(.A(i_2_), .B(ori_ori_n20_), .C(ori_ori_n11_), .D(ori_ori_n13_), .Y(ori_ori_n127_));
  NA2        o117(.A(i_2_), .B(i_4_), .Y(ori_ori_n128_));
  NO2        o118(.A(ori_ori_n88_), .B(ori_ori_n128_), .Y(ori_ori_n129_));
  NO2        o119(.A(i_8_), .B(i_7_), .Y(ori_ori_n130_));
  OA210      o120(.A0(ori_ori_n129_), .A1(ori_ori_n127_), .B0(ori_ori_n130_), .Y(ori_ori_n131_));
  NA3        o121(.A(ori_ori_n99_), .B(i_0_), .C(ori_ori_n22_), .Y(ori_ori_n132_));
  NO2        o122(.A(ori_ori_n132_), .B(i_4_), .Y(ori_ori_n133_));
  NO3        o123(.A(ori_ori_n133_), .B(ori_ori_n131_), .C(ori_ori_n126_), .Y(ori_ori_n134_));
  NA2        o124(.A(ori_ori_n78_), .B(ori_ori_n12_), .Y(ori_ori_n135_));
  NA2        o125(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n136_));
  INV        o126(.A(ori_ori_n46_), .Y(ori_ori_n137_));
  AOI210     o127(.A0(ori_ori_n137_), .A1(ori_ori_n136_), .B0(ori_ori_n135_), .Y(ori_ori_n138_));
  NO2        o128(.A(ori_ori_n85_), .B(ori_ori_n28_), .Y(ori_ori_n139_));
  NA3        o129(.A(ori_ori_n49_), .B(ori_ori_n33_), .C(ori_ori_n14_), .Y(ori_ori_n140_));
  NOi31      o130(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n141_));
  NA2        o131(.A(ori_ori_n116_), .B(ori_ori_n141_), .Y(ori_ori_n142_));
  NA2        o132(.A(ori_ori_n142_), .B(ori_ori_n140_), .Y(ori_ori_n143_));
  NO3        o133(.A(ori_ori_n143_), .B(ori_ori_n139_), .C(ori_ori_n138_), .Y(ori_ori_n144_));
  NA4        o134(.A(ori_ori_n144_), .B(ori_ori_n134_), .C(ori_ori_n124_), .D(ori_ori_n110_), .Y(ori_ori_n145_));
  OR4        o135(.A(ori_ori_n145_), .B(ori_ori_n104_), .C(ori_ori_n77_), .D(ori_ori_n65_), .Y(ori00));
  INV        o136(.A(i_4_), .Y(ori_ori_n149_));
  INV        o137(.A(i_7_), .Y(ori_ori_n150_));
  INV        o138(.A(i_0_), .Y(ori_ori_n151_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NA3        m013(.A(i_6_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_8_), .B(i_6_), .Y(mai_mai_n25_));
  NOi21      m015(.An(i_1_), .B(i_8_), .Y(mai_mai_n26_));
  AOI220     m016(.A0(mai_mai_n26_), .A1(i_2_), .B0(mai_mai_n25_), .B1(i_5_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n22_), .Y(mai_mai_n28_));
  AOI210     m018(.A0(mai_mai_n28_), .A1(mai_mai_n11_), .B0(mai_mai_n20_), .Y(mai_mai_n29_));
  NA2        m019(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n30_));
  NO2        m020(.A(i_2_), .B(i_4_), .Y(mai_mai_n31_));
  NA3        m021(.A(mai_mai_n31_), .B(i_6_), .C(i_8_), .Y(mai_mai_n32_));
  AOI210     m022(.A0(mai_mai_n30_), .A1(i_5_), .B0(mai_mai_n32_), .Y(mai_mai_n33_));
  INV        m023(.A(i_2_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_6_), .B(i_8_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_7_), .B(i_1_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_5_), .B(i_6_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_0_), .B(i_4_), .Y(mai_mai_n38_));
  XO2        m028(.A(i_1_), .B(i_3_), .Y(mai_mai_n39_));
  NOi21      m029(.An(i_7_), .B(i_5_), .Y(mai_mai_n40_));
  AN3        m030(.A(mai_mai_n40_), .B(mai_mai_n39_), .C(mai_mai_n38_), .Y(mai_mai_n41_));
  INV        m031(.A(i_1_), .Y(mai_mai_n42_));
  NOi21      m032(.An(i_3_), .B(i_0_), .Y(mai_mai_n43_));
  NA2        m033(.A(mai_mai_n43_), .B(mai_mai_n42_), .Y(mai_mai_n44_));
  NA3        m034(.A(i_6_), .B(mai_mai_n14_), .C(i_7_), .Y(mai_mai_n45_));
  AOI210     m035(.A0(mai_mai_n45_), .A1(mai_mai_n24_), .B0(mai_mai_n44_), .Y(mai_mai_n46_));
  NO3        m036(.A(mai_mai_n46_), .B(mai_mai_n41_), .C(mai_mai_n33_), .Y(mai_mai_n47_));
  NA2        m037(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n48_));
  NOi21      m038(.An(i_4_), .B(i_0_), .Y(mai_mai_n49_));
  AOI210     m039(.A0(mai_mai_n49_), .A1(mai_mai_n25_), .B0(mai_mai_n15_), .Y(mai_mai_n50_));
  NA2        m040(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n51_));
  NOi21      m041(.An(i_2_), .B(i_8_), .Y(mai_mai_n52_));
  NO3        m042(.A(mai_mai_n52_), .B(mai_mai_n49_), .C(mai_mai_n38_), .Y(mai_mai_n53_));
  NO3        m043(.A(mai_mai_n53_), .B(mai_mai_n51_), .C(mai_mai_n50_), .Y(mai_mai_n54_));
  INV        m044(.A(mai_mai_n54_), .Y(mai_mai_n55_));
  NOi31      m045(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n56_));
  NOi21      m046(.An(i_4_), .B(i_3_), .Y(mai_mai_n57_));
  NOi21      m047(.An(i_1_), .B(i_4_), .Y(mai_mai_n58_));
  AN2        m048(.A(i_8_), .B(i_7_), .Y(mai_mai_n59_));
  NA2        m049(.A(mai_mai_n59_), .B(mai_mai_n12_), .Y(mai_mai_n60_));
  NOi21      m050(.An(i_8_), .B(i_7_), .Y(mai_mai_n61_));
  NA3        m051(.A(mai_mai_n61_), .B(mai_mai_n57_), .C(i_6_), .Y(mai_mai_n62_));
  OAI210     m052(.A0(mai_mai_n60_), .A1(mai_mai_n51_), .B0(mai_mai_n62_), .Y(mai_mai_n63_));
  AOI220     m053(.A0(mai_mai_n63_), .A1(mai_mai_n34_), .B0(mai_mai_n52_), .B1(mai_mai_n37_), .Y(mai_mai_n64_));
  NA4        m054(.A(mai_mai_n64_), .B(mai_mai_n55_), .C(mai_mai_n47_), .D(mai_mai_n29_), .Y(mai_mai_n65_));
  NA2        m055(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n66_));
  AOI220     m056(.A0(mai_mai_n43_), .A1(i_1_), .B0(mai_mai_n39_), .B1(i_2_), .Y(mai_mai_n67_));
  NOi21      m057(.An(i_1_), .B(i_2_), .Y(mai_mai_n68_));
  NO2        m058(.A(mai_mai_n67_), .B(mai_mai_n66_), .Y(mai_mai_n69_));
  NA2        m059(.A(mai_mai_n69_), .B(mai_mai_n14_), .Y(mai_mai_n70_));
  NOi32      m060(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n71_));
  NA2        m061(.A(mai_mai_n71_), .B(i_3_), .Y(mai_mai_n72_));
  NA3        m062(.A(mai_mai_n18_), .B(i_2_), .C(i_6_), .Y(mai_mai_n73_));
  NA2        m063(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  NO2        m064(.A(i_0_), .B(i_4_), .Y(mai_mai_n75_));
  AOI220     m065(.A0(mai_mai_n75_), .A1(mai_mai_n74_), .B0(mai_mai_n26_), .B1(mai_mai_n57_), .Y(mai_mai_n76_));
  NA2        m066(.A(mai_mai_n76_), .B(mai_mai_n70_), .Y(mai_mai_n77_));
  NOi21      m067(.An(i_7_), .B(i_8_), .Y(mai_mai_n78_));
  NOi31      m068(.An(i_6_), .B(i_5_), .C(i_7_), .Y(mai_mai_n79_));
  AOI210     m069(.A0(mai_mai_n78_), .A1(mai_mai_n12_), .B0(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m070(.A(mai_mai_n80_), .B(mai_mai_n11_), .Y(mai_mai_n81_));
  NA2        m071(.A(mai_mai_n81_), .B(mai_mai_n68_), .Y(mai_mai_n82_));
  NA3        m072(.A(mai_mai_n25_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n83_));
  AOI210     m073(.A0(mai_mai_n22_), .A1(mai_mai_n48_), .B0(mai_mai_n83_), .Y(mai_mai_n84_));
  AOI220     m074(.A0(mai_mai_n43_), .A1(mai_mai_n42_), .B0(mai_mai_n18_), .B1(mai_mai_n34_), .Y(mai_mai_n85_));
  NA3        m075(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n86_));
  NO2        m076(.A(mai_mai_n86_), .B(mai_mai_n85_), .Y(mai_mai_n87_));
  NO2        m077(.A(mai_mai_n87_), .B(mai_mai_n84_), .Y(mai_mai_n88_));
  NA3        m078(.A(mai_mai_n61_), .B(mai_mai_n34_), .C(i_3_), .Y(mai_mai_n89_));
  NA2        m079(.A(mai_mai_n42_), .B(i_6_), .Y(mai_mai_n90_));
  AOI210     m080(.A0(mai_mai_n90_), .A1(mai_mai_n22_), .B0(mai_mai_n89_), .Y(mai_mai_n91_));
  NOi21      m081(.An(i_2_), .B(i_1_), .Y(mai_mai_n92_));
  AN3        m082(.A(mai_mai_n78_), .B(mai_mai_n92_), .C(mai_mai_n49_), .Y(mai_mai_n93_));
  NAi21      m083(.An(i_6_), .B(i_0_), .Y(mai_mai_n94_));
  NA3        m084(.A(mai_mai_n58_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n95_));
  NOi21      m085(.An(i_4_), .B(i_6_), .Y(mai_mai_n96_));
  NOi21      m086(.An(i_5_), .B(i_3_), .Y(mai_mai_n97_));
  NO2        m087(.A(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n98_));
  NA2        m088(.A(mai_mai_n68_), .B(mai_mai_n35_), .Y(mai_mai_n99_));
  NOi21      m089(.An(mai_mai_n40_), .B(mai_mai_n99_), .Y(mai_mai_n100_));
  NO4        m090(.A(mai_mai_n100_), .B(mai_mai_n98_), .C(mai_mai_n93_), .D(mai_mai_n91_), .Y(mai_mai_n101_));
  NOi31      m091(.An(mai_mai_n49_), .B(mai_mai_n152_), .C(i_2_), .Y(mai_mai_n102_));
  NA2        m092(.A(mai_mai_n35_), .B(mai_mai_n14_), .Y(mai_mai_n103_));
  NOi21      m093(.An(i_3_), .B(i_1_), .Y(mai_mai_n104_));
  NA2        m094(.A(mai_mai_n104_), .B(i_4_), .Y(mai_mai_n105_));
  NO2        m095(.A(mai_mai_n103_), .B(mai_mai_n105_), .Y(mai_mai_n106_));
  AOI220     m096(.A0(mai_mai_n78_), .A1(mai_mai_n14_), .B0(mai_mai_n96_), .B1(mai_mai_n23_), .Y(mai_mai_n107_));
  NOi31      m097(.An(mai_mai_n43_), .B(mai_mai_n107_), .C(mai_mai_n34_), .Y(mai_mai_n108_));
  NO3        m098(.A(mai_mai_n108_), .B(mai_mai_n106_), .C(mai_mai_n102_), .Y(mai_mai_n109_));
  NA4        m099(.A(mai_mai_n109_), .B(mai_mai_n101_), .C(mai_mai_n88_), .D(mai_mai_n82_), .Y(mai_mai_n110_));
  NA2        m100(.A(mai_mai_n52_), .B(mai_mai_n15_), .Y(mai_mai_n111_));
  INV        m101(.A(mai_mai_n35_), .Y(mai_mai_n112_));
  NA2        m102(.A(mai_mai_n112_), .B(mai_mai_n111_), .Y(mai_mai_n113_));
  NA2        m103(.A(mai_mai_n113_), .B(mai_mai_n38_), .Y(mai_mai_n114_));
  NA4        m104(.A(mai_mai_n59_), .B(mai_mai_n92_), .C(mai_mai_n17_), .D(mai_mai_n12_), .Y(mai_mai_n115_));
  NAi31      m105(.An(mai_mai_n94_), .B(mai_mai_n78_), .C(mai_mai_n92_), .Y(mai_mai_n116_));
  NA3        m106(.A(mai_mai_n61_), .B(mai_mai_n56_), .C(i_6_), .Y(mai_mai_n117_));
  NA3        m107(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(mai_mai_n115_), .Y(mai_mai_n118_));
  NOi21      m108(.An(i_0_), .B(i_2_), .Y(mai_mai_n119_));
  NA3        m109(.A(mai_mai_n119_), .B(mai_mai_n36_), .C(mai_mai_n96_), .Y(mai_mai_n120_));
  NA2        m110(.A(mai_mai_n57_), .B(mai_mai_n35_), .Y(mai_mai_n121_));
  NA2        m111(.A(mai_mai_n121_), .B(mai_mai_n120_), .Y(mai_mai_n122_));
  NA3        m112(.A(mai_mai_n56_), .B(i_6_), .C(i_7_), .Y(mai_mai_n123_));
  NA4        m113(.A(mai_mai_n58_), .B(mai_mai_n37_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n124_));
  NA3        m114(.A(mai_mai_n58_), .B(mai_mai_n43_), .C(i_5_), .Y(mai_mai_n125_));
  NA3        m115(.A(mai_mai_n125_), .B(mai_mai_n124_), .C(mai_mai_n123_), .Y(mai_mai_n126_));
  NO3        m116(.A(mai_mai_n126_), .B(mai_mai_n122_), .C(mai_mai_n118_), .Y(mai_mai_n127_));
  NOi21      m117(.An(i_5_), .B(i_2_), .Y(mai_mai_n128_));
  NA2        m118(.A(mai_mai_n128_), .B(mai_mai_n78_), .Y(mai_mai_n129_));
  AOI210     m119(.A0(mai_mai_n129_), .A1(mai_mai_n111_), .B0(mai_mai_n90_), .Y(mai_mai_n130_));
  NO4        m120(.A(i_2_), .B(mai_mai_n21_), .C(mai_mai_n11_), .D(mai_mai_n14_), .Y(mai_mai_n131_));
  NO2        m121(.A(i_8_), .B(i_7_), .Y(mai_mai_n132_));
  AN2        m122(.A(mai_mai_n131_), .B(mai_mai_n132_), .Y(mai_mai_n133_));
  NA3        m123(.A(mai_mai_n104_), .B(i_0_), .C(i_5_), .Y(mai_mai_n134_));
  NO2        m124(.A(mai_mai_n134_), .B(i_4_), .Y(mai_mai_n135_));
  NO3        m125(.A(mai_mai_n135_), .B(mai_mai_n133_), .C(mai_mai_n130_), .Y(mai_mai_n136_));
  NA2        m126(.A(mai_mai_n78_), .B(mai_mai_n12_), .Y(mai_mai_n137_));
  NA2        m127(.A(i_2_), .B(i_1_), .Y(mai_mai_n138_));
  NA2        m128(.A(mai_mai_n49_), .B(i_3_), .Y(mai_mai_n139_));
  AOI210     m129(.A0(mai_mai_n139_), .A1(mai_mai_n138_), .B0(mai_mai_n137_), .Y(mai_mai_n140_));
  NA2        m130(.A(mai_mai_n61_), .B(mai_mai_n96_), .Y(mai_mai_n141_));
  OAI210     m131(.A0(mai_mai_n89_), .A1(mai_mai_n30_), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  NA3        m132(.A(mai_mai_n97_), .B(mai_mai_n59_), .C(mai_mai_n42_), .Y(mai_mai_n143_));
  NOi31      m133(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n144_));
  NA2        m134(.A(mai_mai_n71_), .B(mai_mai_n144_), .Y(mai_mai_n145_));
  NA2        m135(.A(mai_mai_n145_), .B(mai_mai_n143_), .Y(mai_mai_n146_));
  NO3        m136(.A(mai_mai_n146_), .B(mai_mai_n142_), .C(mai_mai_n140_), .Y(mai_mai_n147_));
  NA4        m137(.A(mai_mai_n147_), .B(mai_mai_n136_), .C(mai_mai_n127_), .D(mai_mai_n114_), .Y(mai_mai_n148_));
  OR4        m138(.A(mai_mai_n148_), .B(mai_mai_n110_), .C(mai_mai_n77_), .D(mai_mai_n65_), .Y(mai00));
  INV        m139(.A(i_8_), .Y(mai_mai_n152_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  INV        u002(.A(i_5_), .Y(men_men_n13_));
  NOi21      u003(.An(i_3_), .B(i_7_), .Y(men_men_n14_));
  INV        u004(.A(i_0_), .Y(men_men_n15_));
  NOi21      u005(.An(i_1_), .B(i_3_), .Y(men_men_n16_));
  INV        u006(.A(i_4_), .Y(men_men_n17_));
  NA2        u007(.A(i_0_), .B(men_men_n17_), .Y(men_men_n18_));
  INV        u008(.A(i_7_), .Y(men_men_n19_));
  NA3        u009(.A(i_6_), .B(i_5_), .C(men_men_n19_), .Y(men_men_n20_));
  NOi21      u010(.An(i_8_), .B(i_6_), .Y(men_men_n21_));
  NOi21      u011(.An(i_1_), .B(i_8_), .Y(men_men_n22_));
  AOI220     u012(.A0(men_men_n22_), .A1(i_2_), .B0(men_men_n21_), .B1(i_5_), .Y(men_men_n23_));
  AOI210     u013(.A0(men_men_n23_), .A1(men_men_n20_), .B0(men_men_n18_), .Y(men_men_n24_));
  NA2        u014(.A(men_men_n24_), .B(men_men_n11_), .Y(men_men_n25_));
  NA2        u015(.A(i_0_), .B(men_men_n13_), .Y(men_men_n26_));
  NA2        u016(.A(men_men_n15_), .B(i_5_), .Y(men_men_n27_));
  NO2        u017(.A(i_2_), .B(i_4_), .Y(men_men_n28_));
  NA3        u018(.A(men_men_n28_), .B(i_6_), .C(i_8_), .Y(men_men_n29_));
  AOI210     u019(.A0(men_men_n27_), .A1(men_men_n26_), .B0(men_men_n29_), .Y(men_men_n30_));
  INV        u020(.A(i_2_), .Y(men_men_n31_));
  NOi21      u021(.An(i_5_), .B(i_0_), .Y(men_men_n32_));
  NOi21      u022(.An(i_6_), .B(i_8_), .Y(men_men_n33_));
  NOi21      u023(.An(i_7_), .B(i_1_), .Y(men_men_n34_));
  NOi21      u024(.An(i_5_), .B(i_6_), .Y(men_men_n35_));
  AOI220     u025(.A0(men_men_n35_), .A1(men_men_n34_), .B0(men_men_n33_), .B1(men_men_n32_), .Y(men_men_n36_));
  NO2        u026(.A(men_men_n36_), .B(i_4_), .Y(men_men_n37_));
  NOi21      u027(.An(i_0_), .B(i_4_), .Y(men_men_n38_));
  XO2        u028(.A(i_1_), .B(i_3_), .Y(men_men_n39_));
  NOi21      u029(.An(i_7_), .B(i_5_), .Y(men_men_n40_));
  AN3        u030(.A(men_men_n40_), .B(men_men_n39_), .C(men_men_n38_), .Y(men_men_n41_));
  INV        u031(.A(i_1_), .Y(men_men_n42_));
  NOi21      u032(.An(i_3_), .B(i_0_), .Y(men_men_n43_));
  NO2        u033(.A(men_men_n20_), .B(i_0_), .Y(men_men_n44_));
  NO4        u034(.A(men_men_n44_), .B(men_men_n41_), .C(men_men_n37_), .D(men_men_n30_), .Y(men_men_n45_));
  INV        u035(.A(i_8_), .Y(men_men_n46_));
  NA2        u036(.A(i_1_), .B(men_men_n11_), .Y(men_men_n47_));
  NO4        u037(.A(men_men_n47_), .B(men_men_n26_), .C(i_2_), .D(men_men_n46_), .Y(men_men_n48_));
  NOi21      u038(.An(i_4_), .B(i_0_), .Y(men_men_n49_));
  AOI210     u039(.A0(men_men_n49_), .A1(men_men_n21_), .B0(men_men_n14_), .Y(men_men_n50_));
  NA2        u040(.A(i_1_), .B(men_men_n13_), .Y(men_men_n51_));
  NOi21      u041(.An(i_2_), .B(i_8_), .Y(men_men_n52_));
  NO3        u042(.A(men_men_n52_), .B(men_men_n49_), .C(men_men_n38_), .Y(men_men_n53_));
  NO3        u043(.A(men_men_n53_), .B(men_men_n51_), .C(men_men_n50_), .Y(men_men_n54_));
  NO2        u044(.A(men_men_n54_), .B(men_men_n48_), .Y(men_men_n55_));
  NOi31      u045(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n56_));
  NA2        u046(.A(men_men_n56_), .B(i_0_), .Y(men_men_n57_));
  NOi21      u047(.An(i_4_), .B(i_3_), .Y(men_men_n58_));
  NOi21      u048(.An(i_1_), .B(i_4_), .Y(men_men_n59_));
  OAI210     u049(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n52_), .Y(men_men_n60_));
  NA2        u050(.A(men_men_n60_), .B(men_men_n57_), .Y(men_men_n61_));
  NOi21      u051(.An(i_8_), .B(i_7_), .Y(men_men_n62_));
  NA2        u052(.A(men_men_n61_), .B(men_men_n35_), .Y(men_men_n63_));
  NA4        u053(.A(men_men_n63_), .B(men_men_n55_), .C(men_men_n45_), .D(men_men_n25_), .Y(men_men_n64_));
  NA2        u054(.A(i_8_), .B(men_men_n19_), .Y(men_men_n65_));
  AOI220     u055(.A0(men_men_n43_), .A1(i_1_), .B0(men_men_n39_), .B1(i_2_), .Y(men_men_n66_));
  NOi21      u056(.An(i_1_), .B(i_2_), .Y(men_men_n67_));
  NA3        u057(.A(men_men_n67_), .B(men_men_n49_), .C(i_6_), .Y(men_men_n68_));
  OAI210     u058(.A0(men_men_n66_), .A1(men_men_n65_), .B0(men_men_n68_), .Y(men_men_n69_));
  NA2        u059(.A(men_men_n69_), .B(men_men_n13_), .Y(men_men_n70_));
  NA3        u060(.A(men_men_n62_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n71_));
  NA3        u061(.A(men_men_n22_), .B(i_0_), .C(men_men_n13_), .Y(men_men_n72_));
  NA2        u062(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n73_));
  NOi32      u063(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n74_));
  NO2        u064(.A(i_0_), .B(i_4_), .Y(men_men_n75_));
  AOI220     u065(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .B1(men_men_n58_), .Y(men_men_n76_));
  NA2        u066(.A(men_men_n76_), .B(men_men_n70_), .Y(men_men_n77_));
  NA2        u067(.A(men_men_n33_), .B(men_men_n32_), .Y(men_men_n78_));
  NOi21      u068(.An(i_7_), .B(i_8_), .Y(men_men_n79_));
  NOi31      u069(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n80_));
  AOI210     u070(.A0(men_men_n79_), .A1(men_men_n12_), .B0(men_men_n80_), .Y(men_men_n81_));
  OAI210     u071(.A0(men_men_n81_), .A1(men_men_n11_), .B0(men_men_n78_), .Y(men_men_n82_));
  NA2        u072(.A(men_men_n82_), .B(men_men_n67_), .Y(men_men_n83_));
  NA3        u073(.A(men_men_n21_), .B(i_2_), .C(men_men_n13_), .Y(men_men_n84_));
  AOI210     u074(.A0(men_men_n18_), .A1(men_men_n47_), .B0(men_men_n84_), .Y(men_men_n85_));
  NA2        u075(.A(men_men_n43_), .B(men_men_n42_), .Y(men_men_n86_));
  NA3        u076(.A(men_men_n17_), .B(i_5_), .C(i_7_), .Y(men_men_n87_));
  NO2        u077(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  NO2        u078(.A(men_men_n88_), .B(men_men_n85_), .Y(men_men_n89_));
  NA3        u079(.A(men_men_n62_), .B(men_men_n31_), .C(i_3_), .Y(men_men_n90_));
  NA2        u080(.A(men_men_n42_), .B(i_6_), .Y(men_men_n91_));
  INV        u081(.A(men_men_n90_), .Y(men_men_n92_));
  NA3        u082(.A(men_men_n59_), .B(i_5_), .C(men_men_n19_), .Y(men_men_n93_));
  NOi21      u083(.An(i_5_), .B(i_3_), .Y(men_men_n94_));
  NA2        u084(.A(men_men_n94_), .B(men_men_n67_), .Y(men_men_n95_));
  OAI210     u085(.A0(men_men_n93_), .A1(i_6_), .B0(men_men_n95_), .Y(men_men_n96_));
  NA2        u086(.A(men_men_n67_), .B(men_men_n33_), .Y(men_men_n97_));
  NOi21      u087(.An(men_men_n40_), .B(men_men_n97_), .Y(men_men_n98_));
  NO3        u088(.A(men_men_n98_), .B(men_men_n96_), .C(men_men_n92_), .Y(men_men_n99_));
  NOi21      u089(.An(i_6_), .B(i_1_), .Y(men_men_n100_));
  AOI220     u090(.A0(men_men_n100_), .A1(i_7_), .B0(men_men_n21_), .B1(i_5_), .Y(men_men_n101_));
  NOi31      u091(.An(men_men_n49_), .B(men_men_n101_), .C(i_2_), .Y(men_men_n102_));
  NOi21      u092(.An(i_3_), .B(i_1_), .Y(men_men_n103_));
  NA2        u093(.A(men_men_n103_), .B(i_4_), .Y(men_men_n104_));
  NO2        u094(.A(i_6_), .B(men_men_n104_), .Y(men_men_n105_));
  NO2        u095(.A(men_men_n105_), .B(men_men_n102_), .Y(men_men_n106_));
  NA4        u096(.A(men_men_n106_), .B(men_men_n99_), .C(men_men_n89_), .D(men_men_n83_), .Y(men_men_n107_));
  NA2        u097(.A(men_men_n52_), .B(men_men_n14_), .Y(men_men_n108_));
  NOi31      u098(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n109_));
  NA2        u099(.A(men_men_n109_), .B(i_7_), .Y(men_men_n110_));
  NA3        u100(.A(men_men_n110_), .B(men_men_n108_), .C(men_men_n97_), .Y(men_men_n111_));
  NA2        u101(.A(men_men_n111_), .B(men_men_n38_), .Y(men_men_n112_));
  NA2        u102(.A(men_men_n58_), .B(men_men_n34_), .Y(men_men_n113_));
  AOI210     u103(.A0(men_men_n113_), .A1(men_men_n71_), .B0(men_men_n27_), .Y(men_men_n114_));
  NA3        u104(.A(men_men_n62_), .B(men_men_n56_), .C(i_6_), .Y(men_men_n115_));
  INV        u105(.A(men_men_n115_), .Y(men_men_n116_));
  NA3        u106(.A(men_men_n49_), .B(men_men_n40_), .C(men_men_n16_), .Y(men_men_n117_));
  INV        u107(.A(men_men_n117_), .Y(men_men_n118_));
  NA3        u108(.A(men_men_n56_), .B(men_men_n13_), .C(i_7_), .Y(men_men_n119_));
  NA4        u109(.A(men_men_n59_), .B(men_men_n35_), .C(men_men_n15_), .D(i_8_), .Y(men_men_n120_));
  NA2        u110(.A(men_men_n120_), .B(men_men_n119_), .Y(men_men_n121_));
  NO4        u111(.A(men_men_n121_), .B(men_men_n118_), .C(men_men_n116_), .D(men_men_n114_), .Y(men_men_n122_));
  AOI210     u112(.A0(i_7_), .A1(men_men_n28_), .B0(men_men_n79_), .Y(men_men_n123_));
  AOI210     u113(.A0(men_men_n123_), .A1(men_men_n108_), .B0(men_men_n91_), .Y(men_men_n124_));
  NO3        u114(.A(i_2_), .B(men_men_n17_), .C(men_men_n11_), .Y(men_men_n125_));
  NA2        u115(.A(i_2_), .B(i_4_), .Y(men_men_n126_));
  AOI210     u116(.A0(i_6_), .A1(i_3_), .B0(men_men_n126_), .Y(men_men_n127_));
  NO2        u117(.A(i_8_), .B(i_7_), .Y(men_men_n128_));
  OA210      u118(.A0(men_men_n127_), .A1(men_men_n125_), .B0(men_men_n128_), .Y(men_men_n129_));
  NA4        u119(.A(men_men_n103_), .B(i_0_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n130_));
  NO2        u120(.A(men_men_n130_), .B(i_4_), .Y(men_men_n131_));
  NO3        u121(.A(men_men_n131_), .B(men_men_n129_), .C(men_men_n124_), .Y(men_men_n132_));
  INV        u122(.A(men_men_n79_), .Y(men_men_n133_));
  NA2        u123(.A(i_2_), .B(men_men_n13_), .Y(men_men_n134_));
  NO2        u124(.A(men_men_n134_), .B(men_men_n133_), .Y(men_men_n135_));
  NA4        u125(.A(men_men_n94_), .B(i_7_), .C(men_men_n42_), .D(men_men_n17_), .Y(men_men_n136_));
  NOi31      u126(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n137_));
  OAI210     u127(.A0(i_4_), .A1(men_men_n74_), .B0(men_men_n137_), .Y(men_men_n138_));
  NA2        u128(.A(men_men_n138_), .B(men_men_n136_), .Y(men_men_n139_));
  NO2        u129(.A(men_men_n139_), .B(men_men_n135_), .Y(men_men_n140_));
  NA4        u130(.A(men_men_n140_), .B(men_men_n132_), .C(men_men_n122_), .D(men_men_n112_), .Y(men_men_n141_));
  OR4        u131(.A(men_men_n141_), .B(men_men_n107_), .C(men_men_n77_), .D(men_men_n64_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule