// Benchmark "top" written by ABC on Thu Jun 20 14:00:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n136_, new_new_n137_, new_new_n138_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n776_, new_new_n777_,
    new_new_n778_, new_new_n779_, new_new_n780_, new_new_n781_,
    new_new_n782_, new_new_n783_, new_new_n784_, new_new_n785_,
    new_new_n786_, new_new_n787_, new_new_n788_, new_new_n789_,
    new_new_n790_, new_new_n791_, new_new_n792_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n825_, new_new_n826_,
    new_new_n827_, new_new_n828_, new_new_n829_, new_new_n830_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n875_,
    new_new_n876_, new_new_n877_, new_new_n878_, new_new_n879_,
    new_new_n880_, new_new_n881_, new_new_n882_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1100_,
    new_new_n1101_, new_new_n1102_, new_new_n1103_, new_new_n1104_,
    new_new_n1105_, new_new_n1106_, new_new_n1107_, new_new_n1108_,
    new_new_n1109_, new_new_n1110_, new_new_n1111_, new_new_n1112_,
    new_new_n1113_, new_new_n1114_, new_new_n1115_, new_new_n1119_,
    new_new_n1120_, new_new_n1121_, new_new_n1122_, new_new_n1123_,
    new_new_n1124_, new_new_n1125_, new_new_n1126_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(zz01));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  OAI210     g0034(.A0(new_new_n56_), .A1(new_new_n53_), .B0(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  NA2        g0038(.A(i_8_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(i_3_), .B(i_9_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_7_), .Y(new_new_n83_));
  NO3        g0061(.A(new_new_n83_), .B(new_new_n82_), .C(new_new_n63_), .Y(new_new_n84_));
  INV        g0062(.A(i_6_), .Y(new_new_n85_));
  OR4        g0063(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n86_));
  INV        g0064(.A(new_new_n86_), .Y(new_new_n87_));
  NO2        g0065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  OAI210     g0066(.A0(new_new_n84_), .A1(i_8_), .B0(new_new_n86_), .Y(new_new_n89_));
  NAi21      g0067(.An(i_6_), .B(i_10_), .Y(new_new_n90_));
  NA2        g0068(.A(i_6_), .B(i_9_), .Y(new_new_n91_));
  AOI210     g0069(.A0(new_new_n91_), .A1(new_new_n90_), .B0(new_new_n63_), .Y(new_new_n92_));
  NA2        g0070(.A(i_2_), .B(i_6_), .Y(new_new_n93_));
  NO3        g0071(.A(new_new_n93_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n94_));
  NO2        g0072(.A(new_new_n94_), .B(new_new_n92_), .Y(new_new_n95_));
  AOI210     g0073(.A0(new_new_n95_), .A1(new_new_n89_), .B0(new_new_n80_), .Y(new_new_n96_));
  AN3        g0074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n97_));
  NAi21      g0075(.An(i_6_), .B(i_11_), .Y(new_new_n98_));
  NO2        g0076(.A(i_5_), .B(i_8_), .Y(new_new_n99_));
  NOi21      g0077(.An(new_new_n99_), .B(new_new_n98_), .Y(new_new_n100_));
  AOI220     g0078(.A0(new_new_n100_), .A1(new_new_n62_), .B0(new_new_n97_), .B1(new_new_n32_), .Y(new_new_n101_));
  INV        g0079(.A(i_7_), .Y(new_new_n102_));
  NA2        g0080(.A(new_new_n47_), .B(new_new_n102_), .Y(new_new_n103_));
  NO2        g0081(.A(i_0_), .B(i_5_), .Y(new_new_n104_));
  NO2        g0082(.A(new_new_n104_), .B(new_new_n85_), .Y(new_new_n105_));
  NA2        g0083(.A(i_12_), .B(i_3_), .Y(new_new_n106_));
  NAi21      g0084(.An(i_7_), .B(i_11_), .Y(new_new_n107_));
  NO3        g0085(.A(new_new_n107_), .B(new_new_n90_), .C(new_new_n54_), .Y(new_new_n108_));
  AN2        g0086(.A(i_2_), .B(i_10_), .Y(new_new_n109_));
  OR2        g0087(.A(new_new_n80_), .B(new_new_n59_), .Y(new_new_n110_));
  NO2        g0088(.A(i_8_), .B(new_new_n102_), .Y(new_new_n111_));
  NA2        g0089(.A(i_12_), .B(i_7_), .Y(new_new_n112_));
  NO2        g0090(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n113_));
  NA2        g0091(.A(new_new_n113_), .B(i_0_), .Y(new_new_n114_));
  NA2        g0092(.A(i_11_), .B(i_12_), .Y(new_new_n115_));
  OAI210     g0093(.A0(new_new_n114_), .A1(new_new_n112_), .B0(new_new_n115_), .Y(new_new_n116_));
  INV        g0094(.A(new_new_n116_), .Y(new_new_n117_));
  NAi31      g0095(.An(new_new_n108_), .B(new_new_n117_), .C(new_new_n101_), .Y(new_new_n118_));
  NOi21      g0096(.An(i_1_), .B(i_5_), .Y(new_new_n119_));
  NA2        g0097(.A(new_new_n119_), .B(i_11_), .Y(new_new_n120_));
  NA2        g0098(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n121_));
  NA2        g0099(.A(i_7_), .B(new_new_n25_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(new_new_n121_), .Y(new_new_n123_));
  NO2        g0101(.A(new_new_n123_), .B(new_new_n47_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n91_), .B(new_new_n90_), .Y(new_new_n125_));
  NAi21      g0103(.An(i_3_), .B(i_8_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(new_new_n62_), .Y(new_new_n127_));
  NOi31      g0105(.An(new_new_n127_), .B(new_new_n125_), .C(new_new_n124_), .Y(new_new_n128_));
  NO2        g0106(.A(i_1_), .B(new_new_n85_), .Y(new_new_n129_));
  NO2        g0107(.A(i_6_), .B(i_5_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n130_), .B(i_3_), .Y(new_new_n131_));
  AO210      g0109(.A0(new_new_n131_), .A1(new_new_n48_), .B0(new_new_n129_), .Y(new_new_n132_));
  OAI220     g0110(.A0(new_new_n132_), .A1(new_new_n107_), .B0(new_new_n128_), .B1(new_new_n120_), .Y(new_new_n133_));
  NO3        g0111(.A(new_new_n133_), .B(new_new_n118_), .C(new_new_n96_), .Y(new_new_n134_));
  NA3        g0112(.A(new_new_n134_), .B(new_new_n79_), .C(new_new_n57_), .Y(zz02));
  NO2        g0113(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n136_));
  NA2        g0114(.A(i_6_), .B(new_new_n25_), .Y(new_new_n137_));
  NA2        g0115(.A(new_new_n137_), .B(new_new_n136_), .Y(new_new_n138_));
  NA4        g0116(.A(new_new_n138_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(zz00));
  AN2        g0117(.A(i_8_), .B(i_7_), .Y(new_new_n140_));
  NA2        g0118(.A(new_new_n140_), .B(i_6_), .Y(new_new_n141_));
  NO2        g0119(.A(i_12_), .B(i_13_), .Y(new_new_n142_));
  NAi21      g0120(.An(i_5_), .B(i_11_), .Y(new_new_n143_));
  NOi21      g0121(.An(new_new_n142_), .B(new_new_n143_), .Y(new_new_n144_));
  NO2        g0122(.A(i_0_), .B(i_1_), .Y(new_new_n145_));
  NA2        g0123(.A(i_2_), .B(i_3_), .Y(new_new_n146_));
  NO2        g0124(.A(new_new_n146_), .B(i_4_), .Y(new_new_n147_));
  NA3        g0125(.A(new_new_n147_), .B(new_new_n145_), .C(new_new_n144_), .Y(new_new_n148_));
  OR2        g0126(.A(new_new_n148_), .B(new_new_n25_), .Y(new_new_n149_));
  AN2        g0127(.A(new_new_n142_), .B(new_new_n82_), .Y(new_new_n150_));
  NO2        g0128(.A(new_new_n150_), .B(new_new_n27_), .Y(new_new_n151_));
  NA2        g0129(.A(i_1_), .B(i_5_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n153_));
  NA2        g0131(.A(new_new_n153_), .B(new_new_n36_), .Y(new_new_n154_));
  NO3        g0132(.A(new_new_n154_), .B(new_new_n152_), .C(new_new_n151_), .Y(new_new_n155_));
  OR2        g0133(.A(i_0_), .B(i_1_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n156_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n157_));
  NAi32      g0135(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n158_));
  NAi21      g0136(.An(new_new_n158_), .B(new_new_n157_), .Y(new_new_n159_));
  NOi21      g0137(.An(i_4_), .B(i_10_), .Y(new_new_n160_));
  NA2        g0138(.A(new_new_n160_), .B(new_new_n40_), .Y(new_new_n161_));
  NO2        g0139(.A(i_3_), .B(i_5_), .Y(new_new_n162_));
  NO3        g0140(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n163_));
  NA2        g0141(.A(new_new_n163_), .B(new_new_n162_), .Y(new_new_n164_));
  OAI210     g0142(.A0(new_new_n164_), .A1(new_new_n161_), .B0(new_new_n159_), .Y(new_new_n165_));
  NO2        g0143(.A(new_new_n165_), .B(new_new_n155_), .Y(new_new_n166_));
  AOI210     g0144(.A0(new_new_n166_), .A1(new_new_n149_), .B0(new_new_n141_), .Y(new_new_n167_));
  NA3        g0145(.A(new_new_n73_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n168_));
  NA2        g0146(.A(i_3_), .B(new_new_n49_), .Y(new_new_n169_));
  NOi21      g0147(.An(i_4_), .B(i_9_), .Y(new_new_n170_));
  NOi21      g0148(.An(i_11_), .B(i_13_), .Y(new_new_n171_));
  NA2        g0149(.A(new_new_n171_), .B(new_new_n170_), .Y(new_new_n172_));
  OR2        g0150(.A(new_new_n172_), .B(new_new_n169_), .Y(new_new_n173_));
  NO2        g0151(.A(i_4_), .B(i_5_), .Y(new_new_n174_));
  NAi21      g0152(.An(i_12_), .B(i_11_), .Y(new_new_n175_));
  NO2        g0153(.A(new_new_n175_), .B(i_13_), .Y(new_new_n176_));
  NA3        g0154(.A(new_new_n176_), .B(new_new_n174_), .C(new_new_n82_), .Y(new_new_n177_));
  AOI210     g0155(.A0(new_new_n177_), .A1(new_new_n173_), .B0(new_new_n168_), .Y(new_new_n178_));
  NO2        g0156(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n179_));
  NA2        g0157(.A(new_new_n179_), .B(new_new_n47_), .Y(new_new_n180_));
  NA2        g0158(.A(new_new_n36_), .B(i_5_), .Y(new_new_n181_));
  NAi31      g0159(.An(new_new_n181_), .B(new_new_n150_), .C(i_11_), .Y(new_new_n182_));
  NA2        g0160(.A(i_3_), .B(i_5_), .Y(new_new_n183_));
  OR2        g0161(.A(new_new_n183_), .B(new_new_n172_), .Y(new_new_n184_));
  AOI210     g0162(.A0(new_new_n184_), .A1(new_new_n182_), .B0(new_new_n180_), .Y(new_new_n185_));
  NO2        g0163(.A(new_new_n73_), .B(i_5_), .Y(new_new_n186_));
  NO2        g0164(.A(i_13_), .B(i_10_), .Y(new_new_n187_));
  NA3        g0165(.A(new_new_n187_), .B(new_new_n186_), .C(new_new_n45_), .Y(new_new_n188_));
  NO2        g0166(.A(i_2_), .B(i_1_), .Y(new_new_n189_));
  NA2        g0167(.A(new_new_n189_), .B(i_3_), .Y(new_new_n190_));
  NAi21      g0168(.An(i_4_), .B(i_12_), .Y(new_new_n191_));
  NO4        g0169(.A(new_new_n191_), .B(new_new_n190_), .C(new_new_n188_), .D(new_new_n25_), .Y(new_new_n192_));
  NO3        g0170(.A(new_new_n192_), .B(new_new_n185_), .C(new_new_n178_), .Y(new_new_n193_));
  INV        g0171(.A(i_8_), .Y(new_new_n194_));
  NO2        g0172(.A(new_new_n194_), .B(i_7_), .Y(new_new_n195_));
  NA2        g0173(.A(new_new_n195_), .B(i_6_), .Y(new_new_n196_));
  NO3        g0174(.A(i_3_), .B(new_new_n85_), .C(new_new_n49_), .Y(new_new_n197_));
  NA2        g0175(.A(new_new_n197_), .B(new_new_n111_), .Y(new_new_n198_));
  NO3        g0176(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n199_));
  NA3        g0177(.A(new_new_n199_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n200_));
  NO3        g0178(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n201_));
  OAI210     g0179(.A0(new_new_n97_), .A1(i_12_), .B0(new_new_n201_), .Y(new_new_n202_));
  AOI210     g0180(.A0(new_new_n202_), .A1(new_new_n200_), .B0(new_new_n198_), .Y(new_new_n203_));
  NO2        g0181(.A(i_3_), .B(i_8_), .Y(new_new_n204_));
  NO3        g0182(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n205_));
  NA3        g0183(.A(new_new_n205_), .B(new_new_n204_), .C(new_new_n40_), .Y(new_new_n206_));
  NO2        g0184(.A(new_new_n104_), .B(new_new_n59_), .Y(new_new_n207_));
  NA2        g0185(.A(new_new_n207_), .B(new_new_n156_), .Y(new_new_n208_));
  NO2        g0186(.A(i_13_), .B(i_9_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(i_6_), .C(new_new_n194_), .Y(new_new_n210_));
  NAi21      g0188(.An(i_12_), .B(i_3_), .Y(new_new_n211_));
  OR2        g0189(.A(new_new_n211_), .B(new_new_n210_), .Y(new_new_n212_));
  NO2        g0190(.A(new_new_n45_), .B(i_5_), .Y(new_new_n213_));
  NO3        g0191(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n214_));
  NA3        g0192(.A(new_new_n214_), .B(new_new_n213_), .C(i_10_), .Y(new_new_n215_));
  OAI220     g0193(.A0(new_new_n215_), .A1(new_new_n212_), .B0(new_new_n208_), .B1(new_new_n206_), .Y(new_new_n216_));
  AOI210     g0194(.A0(new_new_n216_), .A1(i_7_), .B0(new_new_n203_), .Y(new_new_n217_));
  OAI220     g0195(.A0(new_new_n217_), .A1(i_4_), .B0(new_new_n196_), .B1(new_new_n193_), .Y(new_new_n218_));
  NAi21      g0196(.An(i_12_), .B(i_7_), .Y(new_new_n219_));
  NA3        g0197(.A(i_13_), .B(new_new_n194_), .C(i_10_), .Y(new_new_n220_));
  NO2        g0198(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n221_));
  NA2        g0199(.A(i_0_), .B(i_5_), .Y(new_new_n222_));
  NA2        g0200(.A(new_new_n222_), .B(new_new_n105_), .Y(new_new_n223_));
  OAI220     g0201(.A0(new_new_n223_), .A1(new_new_n190_), .B0(new_new_n180_), .B1(new_new_n131_), .Y(new_new_n224_));
  NAi31      g0202(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n36_), .B(i_13_), .Y(new_new_n226_));
  NO2        g0204(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n227_));
  NO2        g0205(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n228_));
  NA3        g0206(.A(new_new_n228_), .B(new_new_n227_), .C(new_new_n226_), .Y(new_new_n229_));
  INV        g0207(.A(i_13_), .Y(new_new_n230_));
  NO2        g0208(.A(i_12_), .B(new_new_n230_), .Y(new_new_n231_));
  NA3        g0209(.A(new_new_n231_), .B(new_new_n199_), .C(new_new_n197_), .Y(new_new_n232_));
  OAI210     g0210(.A0(new_new_n229_), .A1(new_new_n225_), .B0(new_new_n232_), .Y(new_new_n233_));
  AOI220     g0211(.A0(new_new_n233_), .A1(new_new_n140_), .B0(new_new_n224_), .B1(new_new_n221_), .Y(new_new_n234_));
  NO2        g0212(.A(i_12_), .B(new_new_n37_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n183_), .B(i_4_), .Y(new_new_n236_));
  NA2        g0214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  OR2        g0215(.A(i_8_), .B(i_7_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n238_), .B(new_new_n85_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n54_), .B(i_1_), .Y(new_new_n240_));
  NA2        g0218(.A(new_new_n240_), .B(new_new_n239_), .Y(new_new_n241_));
  INV        g0219(.A(i_12_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n45_), .B(new_new_n242_), .Y(new_new_n243_));
  NO3        g0221(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n244_));
  NA2        g0222(.A(i_2_), .B(i_1_), .Y(new_new_n245_));
  NO2        g0223(.A(new_new_n241_), .B(new_new_n237_), .Y(new_new_n246_));
  NO3        g0224(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n247_));
  NAi21      g0225(.An(i_4_), .B(i_3_), .Y(new_new_n248_));
  NO2        g0226(.A(new_new_n248_), .B(new_new_n75_), .Y(new_new_n249_));
  NO2        g0227(.A(i_0_), .B(i_6_), .Y(new_new_n250_));
  NOi41      g0228(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n251_));
  NA2        g0229(.A(new_new_n251_), .B(new_new_n250_), .Y(new_new_n252_));
  NO2        g0230(.A(new_new_n245_), .B(new_new_n183_), .Y(new_new_n253_));
  NAi21      g0231(.An(new_new_n252_), .B(new_new_n253_), .Y(new_new_n254_));
  INV        g0232(.A(new_new_n254_), .Y(new_new_n255_));
  AOI220     g0233(.A0(new_new_n255_), .A1(new_new_n40_), .B0(new_new_n246_), .B1(new_new_n209_), .Y(new_new_n256_));
  NO2        g0234(.A(i_11_), .B(new_new_n230_), .Y(new_new_n257_));
  NOi21      g0235(.An(i_1_), .B(i_6_), .Y(new_new_n258_));
  NAi21      g0236(.An(i_3_), .B(i_7_), .Y(new_new_n259_));
  NA2        g0237(.A(new_new_n242_), .B(i_9_), .Y(new_new_n260_));
  OR4        g0238(.A(new_new_n260_), .B(new_new_n259_), .C(new_new_n258_), .D(new_new_n186_), .Y(new_new_n261_));
  NO2        g0239(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n262_));
  NO2        g0240(.A(i_12_), .B(i_3_), .Y(new_new_n263_));
  NA2        g0241(.A(new_new_n73_), .B(i_5_), .Y(new_new_n264_));
  NA2        g0242(.A(i_3_), .B(i_9_), .Y(new_new_n265_));
  NAi21      g0243(.An(i_7_), .B(i_10_), .Y(new_new_n266_));
  NO2        g0244(.A(new_new_n266_), .B(new_new_n265_), .Y(new_new_n267_));
  NA3        g0245(.A(new_new_n267_), .B(new_new_n264_), .C(new_new_n64_), .Y(new_new_n268_));
  NA2        g0246(.A(new_new_n268_), .B(new_new_n261_), .Y(new_new_n269_));
  NA3        g0247(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n270_));
  INV        g0248(.A(new_new_n141_), .Y(new_new_n271_));
  NA2        g0249(.A(new_new_n242_), .B(i_13_), .Y(new_new_n272_));
  NO2        g0250(.A(new_new_n272_), .B(new_new_n75_), .Y(new_new_n273_));
  AOI220     g0251(.A0(new_new_n273_), .A1(new_new_n271_), .B0(new_new_n269_), .B1(new_new_n257_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n238_), .B(new_new_n37_), .Y(new_new_n275_));
  NA2        g0253(.A(i_12_), .B(i_6_), .Y(new_new_n276_));
  OR2        g0254(.A(i_13_), .B(i_9_), .Y(new_new_n277_));
  NO3        g0255(.A(new_new_n277_), .B(new_new_n276_), .C(new_new_n49_), .Y(new_new_n278_));
  NO2        g0256(.A(new_new_n248_), .B(i_2_), .Y(new_new_n279_));
  NA3        g0257(.A(new_new_n279_), .B(new_new_n278_), .C(new_new_n45_), .Y(new_new_n280_));
  NA2        g0258(.A(new_new_n257_), .B(i_9_), .Y(new_new_n281_));
  OAI210     g0259(.A0(new_new_n73_), .A1(new_new_n281_), .B0(new_new_n280_), .Y(new_new_n282_));
  NA2        g0260(.A(new_new_n153_), .B(new_new_n63_), .Y(new_new_n283_));
  NO3        g0261(.A(i_11_), .B(new_new_n230_), .C(new_new_n25_), .Y(new_new_n284_));
  NO2        g0262(.A(new_new_n259_), .B(i_8_), .Y(new_new_n285_));
  NO2        g0263(.A(i_6_), .B(new_new_n49_), .Y(new_new_n286_));
  NA3        g0264(.A(new_new_n286_), .B(new_new_n285_), .C(new_new_n284_), .Y(new_new_n287_));
  NO3        g0265(.A(new_new_n26_), .B(new_new_n85_), .C(i_5_), .Y(new_new_n288_));
  NA3        g0266(.A(new_new_n288_), .B(new_new_n275_), .C(new_new_n231_), .Y(new_new_n289_));
  AOI210     g0267(.A0(new_new_n289_), .A1(new_new_n287_), .B0(new_new_n283_), .Y(new_new_n290_));
  AOI210     g0268(.A0(new_new_n282_), .A1(new_new_n275_), .B0(new_new_n290_), .Y(new_new_n291_));
  NA4        g0269(.A(new_new_n291_), .B(new_new_n274_), .C(new_new_n256_), .D(new_new_n234_), .Y(new_new_n292_));
  NO3        g0270(.A(i_12_), .B(new_new_n230_), .C(new_new_n37_), .Y(new_new_n293_));
  INV        g0271(.A(new_new_n293_), .Y(new_new_n294_));
  NOi21      g0272(.An(new_new_n162_), .B(new_new_n85_), .Y(new_new_n295_));
  NO3        g0273(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n296_));
  AOI220     g0274(.A0(new_new_n296_), .A1(new_new_n197_), .B0(new_new_n295_), .B1(new_new_n240_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(i_7_), .Y(new_new_n298_));
  NO3        g0276(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n245_), .B(i_0_), .Y(new_new_n300_));
  AOI220     g0278(.A0(new_new_n300_), .A1(new_new_n195_), .B0(new_new_n299_), .B1(new_new_n140_), .Y(new_new_n301_));
  NA2        g0279(.A(new_new_n286_), .B(new_new_n26_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n302_), .B(new_new_n301_), .Y(new_new_n303_));
  NA2        g0281(.A(i_0_), .B(i_1_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n304_), .B(i_2_), .Y(new_new_n305_));
  NO2        g0283(.A(new_new_n60_), .B(i_6_), .Y(new_new_n306_));
  NA3        g0284(.A(new_new_n306_), .B(new_new_n305_), .C(new_new_n162_), .Y(new_new_n307_));
  OAI210     g0285(.A0(new_new_n164_), .A1(new_new_n141_), .B0(new_new_n307_), .Y(new_new_n308_));
  NO3        g0286(.A(new_new_n308_), .B(new_new_n303_), .C(new_new_n298_), .Y(new_new_n309_));
  NO2        g0287(.A(i_3_), .B(i_10_), .Y(new_new_n310_));
  NA3        g0288(.A(new_new_n310_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n311_));
  NO2        g0289(.A(i_2_), .B(new_new_n102_), .Y(new_new_n312_));
  NA2        g0290(.A(i_1_), .B(new_new_n36_), .Y(new_new_n313_));
  NO2        g0291(.A(new_new_n313_), .B(i_8_), .Y(new_new_n314_));
  NOi21      g0292(.An(new_new_n222_), .B(new_new_n104_), .Y(new_new_n315_));
  NA3        g0293(.A(new_new_n315_), .B(new_new_n314_), .C(new_new_n312_), .Y(new_new_n316_));
  AN2        g0294(.A(i_3_), .B(i_10_), .Y(new_new_n317_));
  NA4        g0295(.A(new_new_n317_), .B(new_new_n199_), .C(new_new_n176_), .D(new_new_n174_), .Y(new_new_n318_));
  NO2        g0296(.A(i_5_), .B(new_new_n37_), .Y(new_new_n319_));
  NO2        g0297(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n320_));
  OR2        g0298(.A(new_new_n316_), .B(new_new_n311_), .Y(new_new_n321_));
  OAI220     g0299(.A0(new_new_n321_), .A1(i_6_), .B0(new_new_n309_), .B1(new_new_n294_), .Y(new_new_n322_));
  NO4        g0300(.A(new_new_n322_), .B(new_new_n292_), .C(new_new_n218_), .D(new_new_n167_), .Y(new_new_n323_));
  NO3        g0301(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n324_));
  NO2        g0302(.A(new_new_n60_), .B(new_new_n85_), .Y(new_new_n325_));
  NA2        g0303(.A(new_new_n300_), .B(new_new_n325_), .Y(new_new_n326_));
  NO3        g0304(.A(i_6_), .B(new_new_n194_), .C(i_7_), .Y(new_new_n327_));
  AOI210     g0305(.A0(new_new_n1121_), .A1(new_new_n326_), .B0(new_new_n169_), .Y(new_new_n328_));
  NO2        g0306(.A(i_2_), .B(i_3_), .Y(new_new_n329_));
  OR2        g0307(.A(i_0_), .B(i_5_), .Y(new_new_n330_));
  NA2        g0308(.A(new_new_n222_), .B(new_new_n330_), .Y(new_new_n331_));
  NA4        g0309(.A(new_new_n331_), .B(new_new_n239_), .C(new_new_n329_), .D(i_1_), .Y(new_new_n332_));
  NA3        g0310(.A(new_new_n300_), .B(new_new_n295_), .C(new_new_n111_), .Y(new_new_n333_));
  NAi21      g0311(.An(i_8_), .B(i_7_), .Y(new_new_n334_));
  NO2        g0312(.A(new_new_n334_), .B(i_6_), .Y(new_new_n335_));
  NO2        g0313(.A(new_new_n156_), .B(new_new_n47_), .Y(new_new_n336_));
  NA3        g0314(.A(new_new_n336_), .B(new_new_n335_), .C(new_new_n162_), .Y(new_new_n337_));
  NA3        g0315(.A(new_new_n337_), .B(new_new_n333_), .C(new_new_n332_), .Y(new_new_n338_));
  OAI210     g0316(.A0(new_new_n338_), .A1(new_new_n328_), .B0(i_4_), .Y(new_new_n339_));
  NO2        g0317(.A(i_12_), .B(i_10_), .Y(new_new_n340_));
  NOi21      g0318(.An(i_5_), .B(i_0_), .Y(new_new_n341_));
  AOI210     g0319(.A0(i_2_), .A1(new_new_n49_), .B0(new_new_n102_), .Y(new_new_n342_));
  NO4        g0320(.A(new_new_n342_), .B(new_new_n313_), .C(new_new_n341_), .D(new_new_n126_), .Y(new_new_n343_));
  NA4        g0321(.A(new_new_n83_), .B(new_new_n36_), .C(new_new_n85_), .D(i_8_), .Y(new_new_n344_));
  NA2        g0322(.A(new_new_n343_), .B(new_new_n340_), .Y(new_new_n345_));
  NO2        g0323(.A(i_6_), .B(i_8_), .Y(new_new_n346_));
  NOi21      g0324(.An(i_0_), .B(i_2_), .Y(new_new_n347_));
  AN2        g0325(.A(new_new_n347_), .B(new_new_n346_), .Y(new_new_n348_));
  NO2        g0326(.A(i_1_), .B(i_7_), .Y(new_new_n349_));
  AO220      g0327(.A0(new_new_n349_), .A1(new_new_n348_), .B0(new_new_n335_), .B1(new_new_n240_), .Y(new_new_n350_));
  NA3        g0328(.A(new_new_n350_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n351_));
  NA3        g0329(.A(new_new_n351_), .B(new_new_n345_), .C(new_new_n339_), .Y(new_new_n352_));
  NO3        g0330(.A(new_new_n238_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n353_));
  NO3        g0331(.A(new_new_n334_), .B(i_2_), .C(i_1_), .Y(new_new_n354_));
  OAI210     g0332(.A0(new_new_n354_), .A1(new_new_n353_), .B0(i_6_), .Y(new_new_n355_));
  NA3        g0333(.A(new_new_n258_), .B(new_new_n312_), .C(new_new_n194_), .Y(new_new_n356_));
  AOI210     g0334(.A0(new_new_n356_), .A1(new_new_n355_), .B0(new_new_n331_), .Y(new_new_n357_));
  NOi21      g0335(.An(new_new_n152_), .B(new_new_n105_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n358_), .B(new_new_n122_), .Y(new_new_n359_));
  OAI210     g0337(.A0(new_new_n359_), .A1(new_new_n357_), .B0(i_3_), .Y(new_new_n360_));
  INV        g0338(.A(new_new_n83_), .Y(new_new_n361_));
  NO2        g0339(.A(new_new_n304_), .B(new_new_n81_), .Y(new_new_n362_));
  NA2        g0340(.A(new_new_n362_), .B(new_new_n130_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n93_), .B(new_new_n194_), .Y(new_new_n364_));
  NA3        g0342(.A(new_new_n315_), .B(new_new_n364_), .C(new_new_n63_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n365_), .A1(new_new_n363_), .B0(new_new_n361_), .Y(new_new_n366_));
  NO2        g0344(.A(new_new_n194_), .B(i_9_), .Y(new_new_n367_));
  NA3        g0345(.A(new_new_n367_), .B(new_new_n207_), .C(new_new_n156_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n368_), .B(new_new_n47_), .Y(new_new_n369_));
  NO3        g0347(.A(new_new_n369_), .B(new_new_n366_), .C(new_new_n303_), .Y(new_new_n370_));
  AOI210     g0348(.A0(new_new_n370_), .A1(new_new_n360_), .B0(new_new_n161_), .Y(new_new_n371_));
  AOI210     g0349(.A0(new_new_n352_), .A1(new_new_n324_), .B0(new_new_n371_), .Y(new_new_n372_));
  NOi32      g0350(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n373_));
  INV        g0351(.A(new_new_n373_), .Y(new_new_n374_));
  NAi21      g0352(.An(i_0_), .B(i_6_), .Y(new_new_n375_));
  NAi21      g0353(.An(i_1_), .B(i_5_), .Y(new_new_n376_));
  NA2        g0354(.A(new_new_n376_), .B(new_new_n375_), .Y(new_new_n377_));
  NA2        g0355(.A(new_new_n377_), .B(new_new_n25_), .Y(new_new_n378_));
  OAI210     g0356(.A0(new_new_n378_), .A1(new_new_n158_), .B0(new_new_n252_), .Y(new_new_n379_));
  NAi41      g0357(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n380_));
  OAI220     g0358(.A0(new_new_n380_), .A1(new_new_n376_), .B0(new_new_n225_), .B1(new_new_n158_), .Y(new_new_n381_));
  AOI210     g0359(.A0(new_new_n380_), .A1(new_new_n158_), .B0(new_new_n156_), .Y(new_new_n382_));
  NOi32      g0360(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n383_));
  NAi21      g0361(.An(i_6_), .B(i_1_), .Y(new_new_n384_));
  NA3        g0362(.A(new_new_n384_), .B(new_new_n383_), .C(new_new_n47_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n385_), .B(i_0_), .Y(new_new_n386_));
  OR3        g0364(.A(new_new_n386_), .B(new_new_n382_), .C(new_new_n381_), .Y(new_new_n387_));
  NO2        g0365(.A(i_1_), .B(new_new_n102_), .Y(new_new_n388_));
  NAi21      g0366(.An(i_3_), .B(i_4_), .Y(new_new_n389_));
  NO2        g0367(.A(new_new_n389_), .B(i_9_), .Y(new_new_n390_));
  AN2        g0368(.A(i_6_), .B(i_7_), .Y(new_new_n391_));
  OAI210     g0369(.A0(new_new_n391_), .A1(new_new_n388_), .B0(new_new_n390_), .Y(new_new_n392_));
  NA2        g0370(.A(i_2_), .B(i_7_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n389_), .B(i_10_), .Y(new_new_n394_));
  NA3        g0372(.A(new_new_n394_), .B(new_new_n393_), .C(new_new_n250_), .Y(new_new_n395_));
  AOI210     g0373(.A0(new_new_n395_), .A1(new_new_n392_), .B0(new_new_n186_), .Y(new_new_n396_));
  AOI210     g0374(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n397_));
  OAI210     g0375(.A0(new_new_n397_), .A1(new_new_n189_), .B0(new_new_n394_), .Y(new_new_n398_));
  AOI220     g0376(.A0(new_new_n394_), .A1(new_new_n349_), .B0(new_new_n244_), .B1(new_new_n189_), .Y(new_new_n399_));
  AOI210     g0377(.A0(new_new_n399_), .A1(new_new_n398_), .B0(i_5_), .Y(new_new_n400_));
  NO4        g0378(.A(new_new_n400_), .B(new_new_n396_), .C(new_new_n387_), .D(new_new_n379_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n401_), .B(new_new_n374_), .Y(new_new_n402_));
  NO2        g0380(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n403_));
  AN2        g0381(.A(i_12_), .B(i_5_), .Y(new_new_n404_));
  NO2        g0382(.A(i_4_), .B(new_new_n26_), .Y(new_new_n405_));
  NA2        g0383(.A(new_new_n405_), .B(new_new_n404_), .Y(new_new_n406_));
  NO2        g0384(.A(i_11_), .B(i_6_), .Y(new_new_n407_));
  NA3        g0385(.A(new_new_n407_), .B(new_new_n336_), .C(new_new_n230_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n408_), .B(new_new_n406_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n248_), .B(i_5_), .Y(new_new_n410_));
  NO2        g0388(.A(i_5_), .B(i_10_), .Y(new_new_n411_));
  AOI220     g0389(.A0(new_new_n411_), .A1(new_new_n279_), .B0(new_new_n410_), .B1(new_new_n199_), .Y(new_new_n412_));
  NA2        g0390(.A(new_new_n142_), .B(new_new_n46_), .Y(new_new_n413_));
  NO2        g0391(.A(new_new_n413_), .B(new_new_n412_), .Y(new_new_n414_));
  OAI210     g0392(.A0(new_new_n414_), .A1(new_new_n409_), .B0(new_new_n403_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n148_), .B(new_new_n85_), .Y(new_new_n417_));
  OAI210     g0395(.A0(new_new_n417_), .A1(new_new_n409_), .B0(new_new_n416_), .Y(new_new_n418_));
  NO3        g0396(.A(new_new_n85_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n419_));
  NO2        g0397(.A(i_3_), .B(new_new_n102_), .Y(new_new_n420_));
  NO2        g0398(.A(i_11_), .B(i_12_), .Y(new_new_n421_));
  NA2        g0399(.A(new_new_n411_), .B(new_new_n242_), .Y(new_new_n422_));
  NA3        g0400(.A(new_new_n111_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n423_));
  OAI220     g0401(.A0(new_new_n423_), .A1(new_new_n225_), .B0(new_new_n422_), .B1(new_new_n344_), .Y(new_new_n424_));
  NAi21      g0402(.An(i_13_), .B(i_0_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n425_), .B(new_new_n245_), .Y(new_new_n426_));
  NA2        g0404(.A(new_new_n424_), .B(new_new_n426_), .Y(new_new_n427_));
  NA3        g0405(.A(new_new_n427_), .B(new_new_n418_), .C(new_new_n415_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n45_), .B(new_new_n230_), .Y(new_new_n429_));
  NO3        g0407(.A(i_1_), .B(i_12_), .C(new_new_n85_), .Y(new_new_n430_));
  NO2        g0408(.A(i_0_), .B(i_11_), .Y(new_new_n431_));
  AN2        g0409(.A(i_1_), .B(i_6_), .Y(new_new_n432_));
  NOi21      g0410(.An(i_2_), .B(i_12_), .Y(new_new_n433_));
  NA2        g0411(.A(new_new_n433_), .B(new_new_n432_), .Y(new_new_n434_));
  NO2        g0412(.A(new_new_n434_), .B(new_new_n1119_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n140_), .B(i_9_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n436_), .B(i_4_), .Y(new_new_n437_));
  NA2        g0415(.A(new_new_n435_), .B(new_new_n437_), .Y(new_new_n438_));
  NAi21      g0416(.An(i_9_), .B(i_4_), .Y(new_new_n439_));
  OR2        g0417(.A(i_13_), .B(i_10_), .Y(new_new_n440_));
  NO3        g0418(.A(new_new_n440_), .B(new_new_n115_), .C(new_new_n439_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n172_), .B(new_new_n121_), .Y(new_new_n442_));
  OR2        g0420(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n443_));
  NO2        g0421(.A(new_new_n102_), .B(new_new_n25_), .Y(new_new_n444_));
  NA2        g0422(.A(new_new_n293_), .B(new_new_n444_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n286_), .B(new_new_n214_), .Y(new_new_n446_));
  OAI220     g0424(.A0(new_new_n446_), .A1(new_new_n443_), .B0(new_new_n445_), .B1(new_new_n358_), .Y(new_new_n447_));
  INV        g0425(.A(new_new_n447_), .Y(new_new_n448_));
  AOI210     g0426(.A0(new_new_n448_), .A1(new_new_n438_), .B0(new_new_n26_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n333_), .B(new_new_n332_), .Y(new_new_n450_));
  AOI220     g0428(.A0(new_new_n306_), .A1(new_new_n296_), .B0(new_new_n300_), .B1(new_new_n325_), .Y(new_new_n451_));
  NO2        g0429(.A(new_new_n451_), .B(new_new_n169_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n183_), .B(new_new_n85_), .Y(new_new_n453_));
  AOI220     g0431(.A0(new_new_n453_), .A1(new_new_n305_), .B0(new_new_n288_), .B1(new_new_n214_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n454_), .B(i_7_), .Y(new_new_n455_));
  NO3        g0433(.A(new_new_n455_), .B(new_new_n452_), .C(new_new_n450_), .Y(new_new_n456_));
  NA2        g0434(.A(new_new_n197_), .B(new_new_n97_), .Y(new_new_n457_));
  NA3        g0435(.A(new_new_n336_), .B(new_new_n162_), .C(new_new_n85_), .Y(new_new_n458_));
  AOI210     g0436(.A0(new_new_n458_), .A1(new_new_n457_), .B0(new_new_n334_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n194_), .B(i_10_), .Y(new_new_n460_));
  NA3        g0438(.A(new_new_n264_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n461_));
  NA2        g0439(.A(new_new_n306_), .B(new_new_n240_), .Y(new_new_n462_));
  OAI220     g0440(.A0(new_new_n462_), .A1(new_new_n183_), .B0(new_new_n461_), .B1(new_new_n460_), .Y(new_new_n463_));
  NO2        g0441(.A(i_3_), .B(new_new_n49_), .Y(new_new_n464_));
  NA3        g0442(.A(new_new_n349_), .B(new_new_n348_), .C(new_new_n464_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n327_), .B(new_new_n331_), .Y(new_new_n466_));
  OAI210     g0444(.A0(new_new_n466_), .A1(new_new_n190_), .B0(new_new_n465_), .Y(new_new_n467_));
  NO3        g0445(.A(new_new_n467_), .B(new_new_n463_), .C(new_new_n459_), .Y(new_new_n468_));
  AOI210     g0446(.A0(new_new_n468_), .A1(new_new_n456_), .B0(new_new_n281_), .Y(new_new_n469_));
  NO4        g0447(.A(new_new_n469_), .B(new_new_n449_), .C(new_new_n428_), .D(new_new_n402_), .Y(new_new_n470_));
  NO2        g0448(.A(new_new_n63_), .B(i_4_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n73_), .B(i_13_), .Y(new_new_n472_));
  NA3        g0450(.A(new_new_n472_), .B(new_new_n471_), .C(i_2_), .Y(new_new_n473_));
  NO2        g0451(.A(i_10_), .B(i_9_), .Y(new_new_n474_));
  NAi21      g0452(.An(i_12_), .B(i_8_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n475_), .B(i_3_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n476_), .B(new_new_n474_), .Y(new_new_n477_));
  NO2        g0455(.A(new_new_n47_), .B(i_4_), .Y(new_new_n478_));
  NA2        g0456(.A(new_new_n478_), .B(new_new_n105_), .Y(new_new_n479_));
  OAI220     g0457(.A0(new_new_n479_), .A1(new_new_n206_), .B0(new_new_n477_), .B1(new_new_n473_), .Y(new_new_n480_));
  NA2        g0458(.A(new_new_n320_), .B(i_0_), .Y(new_new_n481_));
  NO3        g0459(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n276_), .B(new_new_n98_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n483_), .B(new_new_n482_), .Y(new_new_n484_));
  NA2        g0462(.A(i_8_), .B(i_9_), .Y(new_new_n485_));
  AOI210     g0463(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n486_));
  OR2        g0464(.A(new_new_n486_), .B(new_new_n485_), .Y(new_new_n487_));
  NA2        g0465(.A(new_new_n293_), .B(new_new_n207_), .Y(new_new_n488_));
  OAI220     g0466(.A0(new_new_n488_), .A1(new_new_n487_), .B0(new_new_n484_), .B1(new_new_n481_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n257_), .B(new_new_n319_), .Y(new_new_n490_));
  NO3        g0468(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n491_));
  AOI210     g0469(.A0(new_new_n263_), .A1(new_new_n189_), .B0(new_new_n491_), .Y(new_new_n492_));
  NA3        g0470(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n493_));
  NA4        g0471(.A(new_new_n143_), .B(new_new_n113_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n494_));
  OAI220     g0472(.A0(new_new_n494_), .A1(new_new_n493_), .B0(new_new_n492_), .B1(new_new_n490_), .Y(new_new_n495_));
  NO3        g0473(.A(new_new_n495_), .B(new_new_n489_), .C(new_new_n480_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n305_), .B(new_new_n107_), .Y(new_new_n497_));
  OR2        g0475(.A(new_new_n497_), .B(new_new_n210_), .Y(new_new_n498_));
  OA210      g0476(.A0(new_new_n368_), .A1(new_new_n102_), .B0(new_new_n307_), .Y(new_new_n499_));
  OA220      g0477(.A0(new_new_n499_), .A1(new_new_n161_), .B0(new_new_n498_), .B1(new_new_n237_), .Y(new_new_n500_));
  NA2        g0478(.A(new_new_n97_), .B(i_13_), .Y(new_new_n501_));
  NA2        g0479(.A(new_new_n453_), .B(new_new_n403_), .Y(new_new_n502_));
  NO2        g0480(.A(i_2_), .B(i_13_), .Y(new_new_n503_));
  NA3        g0481(.A(new_new_n503_), .B(new_new_n160_), .C(new_new_n100_), .Y(new_new_n504_));
  OAI220     g0482(.A0(new_new_n504_), .A1(new_new_n242_), .B0(new_new_n502_), .B1(new_new_n501_), .Y(new_new_n505_));
  NO3        g0483(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n506_));
  NO2        g0484(.A(i_6_), .B(i_7_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n507_), .B(new_new_n506_), .Y(new_new_n508_));
  NO2        g0486(.A(i_11_), .B(i_1_), .Y(new_new_n509_));
  NO2        g0487(.A(new_new_n73_), .B(i_3_), .Y(new_new_n510_));
  OR2        g0488(.A(i_11_), .B(i_8_), .Y(new_new_n511_));
  NOi21      g0489(.An(i_2_), .B(i_7_), .Y(new_new_n512_));
  NAi31      g0490(.An(new_new_n511_), .B(new_new_n512_), .C(new_new_n510_), .Y(new_new_n513_));
  NO2        g0491(.A(new_new_n440_), .B(i_6_), .Y(new_new_n514_));
  NA3        g0492(.A(new_new_n514_), .B(new_new_n471_), .C(new_new_n75_), .Y(new_new_n515_));
  NO2        g0493(.A(new_new_n515_), .B(new_new_n513_), .Y(new_new_n516_));
  NO2        g0494(.A(i_3_), .B(new_new_n194_), .Y(new_new_n517_));
  NO2        g0495(.A(i_6_), .B(i_10_), .Y(new_new_n518_));
  NA4        g0496(.A(new_new_n518_), .B(new_new_n324_), .C(new_new_n517_), .D(new_new_n242_), .Y(new_new_n519_));
  NO2        g0497(.A(new_new_n519_), .B(new_new_n154_), .Y(new_new_n520_));
  NA3        g0498(.A(new_new_n251_), .B(new_new_n171_), .C(new_new_n130_), .Y(new_new_n521_));
  NA2        g0499(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n522_));
  NO2        g0500(.A(new_new_n156_), .B(i_3_), .Y(new_new_n523_));
  NAi31      g0501(.An(new_new_n522_), .B(new_new_n523_), .C(new_new_n231_), .Y(new_new_n524_));
  NA3        g0502(.A(new_new_n416_), .B(new_new_n179_), .C(new_new_n147_), .Y(new_new_n525_));
  NA3        g0503(.A(new_new_n525_), .B(new_new_n524_), .C(new_new_n521_), .Y(new_new_n526_));
  NO4        g0504(.A(new_new_n526_), .B(new_new_n520_), .C(new_new_n516_), .D(new_new_n505_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n491_), .B(new_new_n411_), .Y(new_new_n528_));
  NO2        g0506(.A(new_new_n528_), .B(new_new_n229_), .Y(new_new_n529_));
  NAi21      g0507(.An(new_new_n220_), .B(new_new_n421_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n349_), .B(new_new_n222_), .Y(new_new_n531_));
  NO2        g0509(.A(new_new_n26_), .B(i_5_), .Y(new_new_n532_));
  NO2        g0510(.A(i_0_), .B(new_new_n85_), .Y(new_new_n533_));
  NA3        g0511(.A(new_new_n533_), .B(new_new_n532_), .C(new_new_n140_), .Y(new_new_n534_));
  OR3        g0512(.A(new_new_n313_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n535_));
  OAI220     g0513(.A0(new_new_n535_), .A1(new_new_n534_), .B0(new_new_n531_), .B1(new_new_n530_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n27_), .B(i_10_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n324_), .B(new_new_n244_), .Y(new_new_n538_));
  OAI220     g0516(.A0(new_new_n538_), .A1(new_new_n461_), .B0(new_new_n537_), .B1(new_new_n501_), .Y(new_new_n539_));
  NA4        g0517(.A(new_new_n317_), .B(new_new_n228_), .C(new_new_n73_), .D(new_new_n242_), .Y(new_new_n540_));
  NO2        g0518(.A(new_new_n540_), .B(new_new_n508_), .Y(new_new_n541_));
  NO4        g0519(.A(new_new_n541_), .B(new_new_n539_), .C(new_new_n536_), .D(new_new_n529_), .Y(new_new_n542_));
  NA4        g0520(.A(new_new_n542_), .B(new_new_n527_), .C(new_new_n500_), .D(new_new_n496_), .Y(new_new_n543_));
  NA3        g0521(.A(new_new_n317_), .B(new_new_n176_), .C(new_new_n174_), .Y(new_new_n544_));
  OAI210     g0522(.A0(new_new_n311_), .A1(new_new_n181_), .B0(new_new_n544_), .Y(new_new_n545_));
  AN2        g0523(.A(new_new_n296_), .B(new_new_n239_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n546_), .B(new_new_n545_), .Y(new_new_n547_));
  NA2        g0525(.A(new_new_n120_), .B(new_new_n110_), .Y(new_new_n548_));
  AO220      g0526(.A0(new_new_n548_), .A1(new_new_n482_), .B0(new_new_n441_), .B1(i_6_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n324_), .B(new_new_n163_), .Y(new_new_n550_));
  OAI210     g0528(.A0(new_new_n550_), .A1(new_new_n237_), .B0(new_new_n318_), .Y(new_new_n551_));
  AOI220     g0529(.A0(new_new_n551_), .A1(new_new_n335_), .B0(new_new_n549_), .B1(new_new_n320_), .Y(new_new_n552_));
  NA4        g0530(.A(new_new_n472_), .B(new_new_n471_), .C(new_new_n204_), .D(i_2_), .Y(new_new_n553_));
  INV        g0531(.A(new_new_n553_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n404_), .B(new_new_n230_), .Y(new_new_n555_));
  NA2        g0533(.A(new_new_n373_), .B(new_new_n73_), .Y(new_new_n556_));
  NA2        g0534(.A(new_new_n391_), .B(new_new_n383_), .Y(new_new_n557_));
  AO210      g0535(.A0(new_new_n556_), .A1(new_new_n555_), .B0(new_new_n557_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n36_), .B(i_8_), .Y(new_new_n559_));
  AOI210     g0537(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n441_), .Y(new_new_n560_));
  NA2        g0538(.A(new_new_n560_), .B(new_new_n558_), .Y(new_new_n561_));
  AOI210     g0539(.A0(new_new_n554_), .A1(new_new_n205_), .B0(new_new_n561_), .Y(new_new_n562_));
  NA2        g0540(.A(new_new_n264_), .B(new_new_n64_), .Y(new_new_n563_));
  OAI210     g0541(.A0(i_8_), .A1(new_new_n563_), .B0(new_new_n132_), .Y(new_new_n564_));
  AOI210     g0542(.A0(new_new_n195_), .A1(i_9_), .B0(new_new_n275_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n565_), .B(new_new_n200_), .Y(new_new_n566_));
  OR2        g0544(.A(new_new_n183_), .B(i_4_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n567_), .B(new_new_n85_), .Y(new_new_n568_));
  AOI220     g0546(.A0(new_new_n568_), .A1(new_new_n566_), .B0(new_new_n564_), .B1(new_new_n442_), .Y(new_new_n569_));
  NA4        g0547(.A(new_new_n569_), .B(new_new_n562_), .C(new_new_n552_), .D(new_new_n547_), .Y(new_new_n570_));
  NA2        g0548(.A(new_new_n410_), .B(new_new_n305_), .Y(new_new_n571_));
  OAI210     g0549(.A0(new_new_n406_), .A1(new_new_n168_), .B0(new_new_n571_), .Y(new_new_n572_));
  NO2        g0550(.A(i_12_), .B(new_new_n194_), .Y(new_new_n573_));
  NA2        g0551(.A(new_new_n573_), .B(new_new_n230_), .Y(new_new_n574_));
  NA3        g0552(.A(new_new_n518_), .B(new_new_n174_), .C(new_new_n27_), .Y(new_new_n575_));
  NO3        g0553(.A(new_new_n575_), .B(new_new_n574_), .C(new_new_n497_), .Y(new_new_n576_));
  NOi31      g0554(.An(new_new_n327_), .B(new_new_n440_), .C(new_new_n38_), .Y(new_new_n577_));
  OAI210     g0555(.A0(new_new_n577_), .A1(new_new_n576_), .B0(new_new_n572_), .Y(new_new_n578_));
  NO2        g0556(.A(i_8_), .B(i_7_), .Y(new_new_n579_));
  OAI210     g0557(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n580_));
  NA2        g0558(.A(new_new_n580_), .B(new_new_n228_), .Y(new_new_n581_));
  AOI220     g0559(.A0(new_new_n336_), .A1(new_new_n40_), .B0(new_new_n240_), .B1(new_new_n209_), .Y(new_new_n582_));
  OAI220     g0560(.A0(new_new_n582_), .A1(new_new_n567_), .B0(new_new_n581_), .B1(new_new_n248_), .Y(new_new_n583_));
  NA2        g0561(.A(new_new_n45_), .B(i_10_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n584_), .B(i_6_), .Y(new_new_n585_));
  NA3        g0563(.A(new_new_n585_), .B(new_new_n583_), .C(new_new_n579_), .Y(new_new_n586_));
  AOI220     g0564(.A0(new_new_n453_), .A1(new_new_n336_), .B0(new_new_n253_), .B1(new_new_n250_), .Y(new_new_n587_));
  OAI220     g0565(.A0(new_new_n587_), .A1(new_new_n272_), .B0(new_new_n501_), .B1(new_new_n131_), .Y(new_new_n588_));
  NA2        g0566(.A(new_new_n588_), .B(new_new_n275_), .Y(new_new_n589_));
  NOi31      g0567(.An(new_new_n300_), .B(new_new_n311_), .C(new_new_n181_), .Y(new_new_n590_));
  NA3        g0568(.A(new_new_n317_), .B(new_new_n174_), .C(new_new_n97_), .Y(new_new_n591_));
  NO2        g0569(.A(new_new_n226_), .B(new_new_n45_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n156_), .B(i_5_), .Y(new_new_n593_));
  NA3        g0571(.A(new_new_n593_), .B(new_new_n429_), .C(new_new_n329_), .Y(new_new_n594_));
  OAI210     g0572(.A0(new_new_n594_), .A1(new_new_n592_), .B0(new_new_n591_), .Y(new_new_n595_));
  OAI210     g0573(.A0(new_new_n595_), .A1(new_new_n590_), .B0(new_new_n491_), .Y(new_new_n596_));
  NA4        g0574(.A(new_new_n596_), .B(new_new_n589_), .C(new_new_n586_), .D(new_new_n578_), .Y(new_new_n597_));
  NA3        g0575(.A(new_new_n222_), .B(new_new_n71_), .C(new_new_n45_), .Y(new_new_n598_));
  NA2        g0576(.A(new_new_n293_), .B(new_new_n83_), .Y(new_new_n599_));
  AOI210     g0577(.A0(new_new_n598_), .A1(new_new_n363_), .B0(new_new_n599_), .Y(new_new_n600_));
  NA2        g0578(.A(new_new_n306_), .B(new_new_n296_), .Y(new_new_n601_));
  NO2        g0579(.A(new_new_n601_), .B(new_new_n173_), .Y(new_new_n602_));
  NA2        g0580(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n603_));
  NA2        g0581(.A(new_new_n474_), .B(new_new_n226_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n603_), .B(new_new_n604_), .Y(new_new_n605_));
  AOI210     g0583(.A0(new_new_n384_), .A1(new_new_n47_), .B0(new_new_n388_), .Y(new_new_n606_));
  NA2        g0584(.A(i_0_), .B(new_new_n49_), .Y(new_new_n607_));
  NA3        g0585(.A(new_new_n573_), .B(new_new_n284_), .C(new_new_n607_), .Y(new_new_n608_));
  NO2        g0586(.A(new_new_n606_), .B(new_new_n608_), .Y(new_new_n609_));
  NO4        g0587(.A(new_new_n609_), .B(new_new_n605_), .C(new_new_n602_), .D(new_new_n600_), .Y(new_new_n610_));
  NO4        g0588(.A(new_new_n258_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n611_));
  NO3        g0589(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n612_));
  NO2        g0590(.A(new_new_n238_), .B(new_new_n36_), .Y(new_new_n613_));
  AN2        g0591(.A(new_new_n613_), .B(new_new_n612_), .Y(new_new_n614_));
  OA210      g0592(.A0(new_new_n614_), .A1(new_new_n611_), .B0(new_new_n373_), .Y(new_new_n615_));
  NO2        g0593(.A(new_new_n440_), .B(i_1_), .Y(new_new_n616_));
  NOi31      g0594(.An(new_new_n616_), .B(new_new_n483_), .C(new_new_n73_), .Y(new_new_n617_));
  AN4        g0595(.A(new_new_n617_), .B(new_new_n437_), .C(new_new_n532_), .D(i_2_), .Y(new_new_n618_));
  NO2        g0596(.A(new_new_n451_), .B(new_new_n177_), .Y(new_new_n619_));
  NO3        g0597(.A(new_new_n619_), .B(new_new_n618_), .C(new_new_n615_), .Y(new_new_n620_));
  NOi21      g0598(.An(i_10_), .B(i_6_), .Y(new_new_n621_));
  NO2        g0599(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n622_));
  AOI220     g0600(.A0(new_new_n293_), .A1(new_new_n622_), .B0(new_new_n284_), .B1(new_new_n621_), .Y(new_new_n623_));
  NO2        g0601(.A(new_new_n623_), .B(new_new_n481_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n112_), .B(new_new_n23_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n327_), .B(new_new_n163_), .Y(new_new_n626_));
  AOI220     g0604(.A0(new_new_n626_), .A1(new_new_n462_), .B0(new_new_n184_), .B1(new_new_n182_), .Y(new_new_n627_));
  NO2        g0605(.A(new_new_n199_), .B(new_new_n37_), .Y(new_new_n628_));
  NOi31      g0606(.An(new_new_n144_), .B(new_new_n628_), .C(new_new_n344_), .Y(new_new_n629_));
  NO3        g0607(.A(new_new_n629_), .B(new_new_n627_), .C(new_new_n624_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n556_), .B(new_new_n399_), .Y(new_new_n631_));
  INV        g0609(.A(new_new_n329_), .Y(new_new_n632_));
  NO2        g0610(.A(i_12_), .B(new_new_n85_), .Y(new_new_n633_));
  NA3        g0611(.A(new_new_n633_), .B(new_new_n284_), .C(new_new_n607_), .Y(new_new_n634_));
  NA3        g0612(.A(new_new_n407_), .B(new_new_n293_), .C(new_new_n222_), .Y(new_new_n635_));
  AOI210     g0613(.A0(new_new_n635_), .A1(new_new_n634_), .B0(new_new_n632_), .Y(new_new_n636_));
  NA2        g0614(.A(new_new_n174_), .B(i_0_), .Y(new_new_n637_));
  NO3        g0615(.A(new_new_n637_), .B(new_new_n355_), .C(new_new_n311_), .Y(new_new_n638_));
  OR2        g0616(.A(i_2_), .B(i_5_), .Y(new_new_n639_));
  OR2        g0617(.A(new_new_n639_), .B(new_new_n432_), .Y(new_new_n640_));
  AOI210     g0618(.A0(new_new_n393_), .A1(new_new_n250_), .B0(new_new_n199_), .Y(new_new_n641_));
  AOI210     g0619(.A0(new_new_n641_), .A1(new_new_n640_), .B0(new_new_n530_), .Y(new_new_n642_));
  NO4        g0620(.A(new_new_n642_), .B(new_new_n638_), .C(new_new_n636_), .D(new_new_n631_), .Y(new_new_n643_));
  NA4        g0621(.A(new_new_n643_), .B(new_new_n630_), .C(new_new_n620_), .D(new_new_n610_), .Y(new_new_n644_));
  NO4        g0622(.A(new_new_n644_), .B(new_new_n597_), .C(new_new_n570_), .D(new_new_n543_), .Y(new_new_n645_));
  NA4        g0623(.A(new_new_n645_), .B(new_new_n470_), .C(new_new_n372_), .D(new_new_n323_), .Y(zz07));
  OAI220     g0624(.A0(new_new_n537_), .A1(new_new_n115_), .B0(new_new_n93_), .B1(new_new_n55_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n107_), .B(new_new_n90_), .Y(new_new_n648_));
  NA2        g0626(.A(new_new_n405_), .B(new_new_n648_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n518_), .B(new_new_n83_), .Y(new_new_n650_));
  NA2        g0628(.A(new_new_n142_), .B(i_8_), .Y(new_new_n651_));
  OAI210     g0629(.A0(new_new_n651_), .A1(new_new_n650_), .B0(new_new_n649_), .Y(new_new_n652_));
  NA3        g0630(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n653_));
  NO2        g0631(.A(new_new_n242_), .B(i_4_), .Y(new_new_n654_));
  NA2        g0632(.A(new_new_n654_), .B(i_8_), .Y(new_new_n655_));
  AOI210     g0633(.A0(new_new_n655_), .A1(new_new_n106_), .B0(new_new_n653_), .Y(new_new_n656_));
  NA2        g0634(.A(i_2_), .B(new_new_n85_), .Y(new_new_n657_));
  OAI210     g0635(.A0(new_new_n88_), .A1(new_new_n204_), .B0(new_new_n205_), .Y(new_new_n658_));
  NO2        g0636(.A(i_7_), .B(new_new_n37_), .Y(new_new_n659_));
  NA2        g0637(.A(i_4_), .B(i_8_), .Y(new_new_n660_));
  AOI210     g0638(.A0(new_new_n660_), .A1(new_new_n317_), .B0(new_new_n659_), .Y(new_new_n661_));
  OAI220     g0639(.A0(new_new_n661_), .A1(new_new_n657_), .B0(new_new_n658_), .B1(i_13_), .Y(new_new_n662_));
  NO4        g0640(.A(new_new_n662_), .B(new_new_n656_), .C(new_new_n652_), .D(new_new_n647_), .Y(new_new_n663_));
  AOI210     g0641(.A0(new_new_n126_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n664_));
  AOI210     g0642(.A0(new_new_n664_), .A1(new_new_n242_), .B0(new_new_n160_), .Y(new_new_n665_));
  NO2        g0643(.A(i_10_), .B(new_new_n23_), .Y(new_new_n666_));
  OR3        g0644(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n667_));
  NO3        g0645(.A(new_new_n667_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n668_));
  INV        g0646(.A(new_new_n201_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n668_), .B(new_new_n666_), .Y(new_new_n670_));
  OA220      g0648(.A0(new_new_n670_), .A1(new_new_n632_), .B0(new_new_n665_), .B1(new_new_n277_), .Y(new_new_n671_));
  AOI210     g0649(.A0(new_new_n671_), .A1(new_new_n663_), .B0(new_new_n63_), .Y(new_new_n672_));
  NOi21      g0650(.An(i_11_), .B(i_7_), .Y(new_new_n673_));
  AO210      g0651(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n673_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n675_), .B(new_new_n209_), .Y(new_new_n676_));
  NA3        g0654(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n677_));
  NAi31      g0655(.An(new_new_n677_), .B(new_new_n219_), .C(i_11_), .Y(new_new_n678_));
  AOI210     g0656(.A0(new_new_n678_), .A1(new_new_n676_), .B0(new_new_n63_), .Y(new_new_n679_));
  NA2        g0657(.A(new_new_n87_), .B(new_new_n63_), .Y(new_new_n680_));
  AO210      g0658(.A0(new_new_n680_), .A1(new_new_n399_), .B0(new_new_n41_), .Y(new_new_n681_));
  NO3        g0659(.A(new_new_n266_), .B(new_new_n211_), .C(i_8_), .Y(new_new_n682_));
  OAI210     g0660(.A0(new_new_n682_), .A1(new_new_n231_), .B0(new_new_n63_), .Y(new_new_n683_));
  NA2        g0661(.A(new_new_n433_), .B(new_new_n31_), .Y(new_new_n684_));
  OR2        g0662(.A(new_new_n211_), .B(new_new_n107_), .Y(new_new_n685_));
  INV        g0663(.A(new_new_n684_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n63_), .B(i_9_), .Y(new_new_n687_));
  INV        g0665(.A(i_4_), .Y(new_new_n688_));
  NA2        g0666(.A(new_new_n688_), .B(new_new_n686_), .Y(new_new_n689_));
  NO2        g0667(.A(i_1_), .B(i_12_), .Y(new_new_n690_));
  NA3        g0668(.A(new_new_n690_), .B(new_new_n109_), .C(new_new_n24_), .Y(new_new_n691_));
  NA4        g0669(.A(new_new_n691_), .B(new_new_n689_), .C(new_new_n683_), .D(new_new_n681_), .Y(new_new_n692_));
  OAI210     g0670(.A0(new_new_n692_), .A1(new_new_n679_), .B0(i_6_), .Y(new_new_n693_));
  OAI210     g0671(.A0(new_new_n677_), .A1(new_new_n107_), .B0(new_new_n493_), .Y(new_new_n694_));
  NA2        g0672(.A(new_new_n694_), .B(new_new_n633_), .Y(new_new_n695_));
  NA3        g0673(.A(new_new_n695_), .B(new_new_n560_), .C(new_new_n484_), .Y(new_new_n696_));
  NO4        g0674(.A(new_new_n219_), .B(new_new_n126_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n697_));
  NA2        g0675(.A(new_new_n697_), .B(new_new_n687_), .Y(new_new_n698_));
  NA2        g0676(.A(new_new_n242_), .B(i_6_), .Y(new_new_n699_));
  NO3        g0677(.A(i_10_), .B(new_new_n238_), .C(new_new_n23_), .Y(new_new_n700_));
  AOI210     g0678(.A0(i_1_), .A1(new_new_n267_), .B0(new_new_n700_), .Y(new_new_n701_));
  OAI210     g0679(.A0(new_new_n701_), .A1(new_new_n45_), .B0(new_new_n698_), .Y(new_new_n702_));
  NA3        g0680(.A(new_new_n579_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n703_));
  NA3        g0681(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n704_));
  NA3        g0682(.A(new_new_n1126_), .B(new_new_n276_), .C(new_new_n45_), .Y(new_new_n705_));
  NO2        g0683(.A(new_new_n705_), .B(new_new_n704_), .Y(new_new_n706_));
  NA3        g0684(.A(new_new_n687_), .B(new_new_n329_), .C(i_6_), .Y(new_new_n707_));
  NO2        g0685(.A(new_new_n707_), .B(new_new_n23_), .Y(new_new_n708_));
  AOI210     g0686(.A0(new_new_n509_), .A1(new_new_n444_), .B0(new_new_n247_), .Y(new_new_n709_));
  NO2        g0687(.A(new_new_n709_), .B(new_new_n657_), .Y(new_new_n710_));
  NAi21      g0688(.An(new_new_n703_), .B(new_new_n92_), .Y(new_new_n711_));
  NO2        g0689(.A(i_11_), .B(new_new_n37_), .Y(new_new_n712_));
  NA2        g0690(.A(new_new_n712_), .B(new_new_n24_), .Y(new_new_n713_));
  OAI210     g0691(.A0(new_new_n713_), .A1(i_6_), .B0(new_new_n711_), .Y(new_new_n714_));
  OR4        g0692(.A(new_new_n714_), .B(new_new_n710_), .C(new_new_n708_), .D(new_new_n706_), .Y(new_new_n715_));
  NO3        g0693(.A(new_new_n715_), .B(new_new_n702_), .C(new_new_n696_), .Y(new_new_n716_));
  NO2        g0694(.A(new_new_n242_), .B(new_new_n102_), .Y(new_new_n717_));
  NO2        g0695(.A(new_new_n717_), .B(new_new_n673_), .Y(new_new_n718_));
  NA2        g0696(.A(new_new_n718_), .B(i_1_), .Y(new_new_n719_));
  NO2        g0697(.A(new_new_n719_), .B(new_new_n667_), .Y(new_new_n720_));
  NO2        g0698(.A(new_new_n439_), .B(new_new_n85_), .Y(new_new_n721_));
  NA2        g0699(.A(new_new_n720_), .B(new_new_n47_), .Y(new_new_n722_));
  NA2        g0700(.A(i_3_), .B(new_new_n194_), .Y(new_new_n723_));
  AOI210     g0701(.A0(new_new_n265_), .A1(new_new_n723_), .B0(new_new_n112_), .Y(new_new_n724_));
  AN2        g0702(.A(new_new_n724_), .B(new_new_n585_), .Y(new_new_n725_));
  NO2        g0703(.A(new_new_n238_), .B(new_new_n45_), .Y(new_new_n726_));
  NO3        g0704(.A(new_new_n726_), .B(new_new_n320_), .C(new_new_n243_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n115_), .B(new_new_n37_), .Y(new_new_n728_));
  NO2        g0706(.A(new_new_n728_), .B(i_6_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n85_), .B(i_9_), .Y(new_new_n730_));
  NO2        g0708(.A(new_new_n730_), .B(new_new_n63_), .Y(new_new_n731_));
  NO2        g0709(.A(new_new_n731_), .B(new_new_n690_), .Y(new_new_n732_));
  NO4        g0710(.A(new_new_n732_), .B(new_new_n729_), .C(new_new_n727_), .D(i_4_), .Y(new_new_n733_));
  NA2        g0711(.A(i_1_), .B(i_3_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n485_), .B(new_new_n93_), .Y(new_new_n735_));
  AOI210     g0713(.A0(new_new_n726_), .A1(new_new_n621_), .B0(new_new_n735_), .Y(new_new_n736_));
  NO2        g0714(.A(new_new_n736_), .B(new_new_n734_), .Y(new_new_n737_));
  NO3        g0715(.A(new_new_n737_), .B(new_new_n733_), .C(new_new_n725_), .Y(new_new_n738_));
  NA4        g0716(.A(new_new_n738_), .B(new_new_n722_), .C(new_new_n716_), .D(new_new_n693_), .Y(new_new_n739_));
  NO3        g0717(.A(new_new_n511_), .B(i_3_), .C(i_7_), .Y(new_new_n740_));
  NOi21      g0718(.An(new_new_n740_), .B(i_10_), .Y(new_new_n741_));
  OA210      g0719(.A0(new_new_n741_), .A1(new_new_n251_), .B0(new_new_n85_), .Y(new_new_n742_));
  NA2        g0720(.A(new_new_n391_), .B(new_new_n390_), .Y(new_new_n743_));
  NA3        g0721(.A(new_new_n518_), .B(new_new_n559_), .C(new_new_n47_), .Y(new_new_n744_));
  NO3        g0722(.A(new_new_n512_), .B(new_new_n660_), .C(new_new_n85_), .Y(new_new_n745_));
  NA2        g0723(.A(new_new_n745_), .B(new_new_n25_), .Y(new_new_n746_));
  NA3        g0724(.A(new_new_n160_), .B(new_new_n83_), .C(new_new_n85_), .Y(new_new_n747_));
  NA4        g0725(.A(new_new_n747_), .B(new_new_n746_), .C(new_new_n744_), .D(new_new_n743_), .Y(new_new_n748_));
  OAI210     g0726(.A0(new_new_n748_), .A1(new_new_n742_), .B0(i_1_), .Y(new_new_n749_));
  AOI210     g0727(.A0(new_new_n707_), .A1(new_new_n749_), .B0(i_13_), .Y(new_new_n750_));
  OR2        g0728(.A(i_11_), .B(i_7_), .Y(new_new_n751_));
  NA3        g0729(.A(new_new_n751_), .B(i_3_), .C(new_new_n136_), .Y(new_new_n752_));
  AOI220     g0730(.A0(new_new_n503_), .A1(new_new_n160_), .B0(new_new_n478_), .B1(new_new_n136_), .Y(new_new_n753_));
  OAI210     g0731(.A0(new_new_n753_), .A1(new_new_n45_), .B0(new_new_n752_), .Y(new_new_n754_));
  NO2        g0732(.A(new_new_n512_), .B(new_new_n24_), .Y(new_new_n755_));
  AOI220     g0733(.A0(new_new_n755_), .A1(new_new_n721_), .B0(new_new_n251_), .B1(new_new_n129_), .Y(new_new_n756_));
  OAI220     g0734(.A0(new_new_n756_), .A1(new_new_n41_), .B0(new_new_n55_), .B1(new_new_n93_), .Y(new_new_n757_));
  AOI210     g0735(.A0(new_new_n754_), .A1(new_new_n346_), .B0(new_new_n757_), .Y(new_new_n758_));
  AOI220     g0736(.A0(i_7_), .A1(new_new_n72_), .B0(new_new_n407_), .B1(new_new_n1126_), .Y(new_new_n759_));
  NO2        g0737(.A(new_new_n759_), .B(new_new_n248_), .Y(new_new_n760_));
  AOI210     g0738(.A0(new_new_n475_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n761_));
  NOi31      g0739(.An(new_new_n761_), .B(new_new_n650_), .C(new_new_n45_), .Y(new_new_n762_));
  NA2        g0740(.A(new_new_n125_), .B(i_13_), .Y(new_new_n763_));
  NO2        g0741(.A(new_new_n704_), .B(new_new_n112_), .Y(new_new_n764_));
  INV        g0742(.A(new_new_n764_), .Y(new_new_n765_));
  OAI220     g0743(.A0(new_new_n765_), .A1(new_new_n71_), .B0(new_new_n763_), .B1(new_new_n1122_), .Y(new_new_n766_));
  NO3        g0744(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n102_), .Y(new_new_n767_));
  NA2        g0745(.A(new_new_n26_), .B(new_new_n194_), .Y(new_new_n768_));
  NA2        g0746(.A(new_new_n768_), .B(i_7_), .Y(new_new_n769_));
  NO3        g0747(.A(new_new_n512_), .B(new_new_n242_), .C(new_new_n85_), .Y(new_new_n770_));
  AOI210     g0748(.A0(new_new_n770_), .A1(new_new_n769_), .B0(new_new_n767_), .Y(new_new_n771_));
  OAI220     g0749(.A0(new_new_n1125_), .A1(new_new_n655_), .B0(new_new_n771_), .B1(new_new_n669_), .Y(new_new_n772_));
  NO4        g0750(.A(new_new_n772_), .B(new_new_n766_), .C(new_new_n762_), .D(new_new_n760_), .Y(new_new_n773_));
  OR2        g0751(.A(i_11_), .B(i_6_), .Y(new_new_n774_));
  AOI210     g0752(.A0(new_new_n242_), .A1(new_new_n765_), .B0(new_new_n774_), .Y(new_new_n775_));
  NA2        g0753(.A(new_new_n103_), .B(new_new_n768_), .Y(new_new_n776_));
  NAi21      g0754(.An(i_11_), .B(i_12_), .Y(new_new_n777_));
  NO3        g0755(.A(new_new_n777_), .B(i_13_), .C(new_new_n85_), .Y(new_new_n778_));
  NO3        g0756(.A(new_new_n512_), .B(new_new_n633_), .C(new_new_n660_), .Y(new_new_n779_));
  AOI220     g0757(.A0(new_new_n779_), .A1(new_new_n324_), .B0(new_new_n778_), .B1(new_new_n776_), .Y(new_new_n780_));
  INV        g0758(.A(new_new_n780_), .Y(new_new_n781_));
  OAI210     g0759(.A0(new_new_n781_), .A1(new_new_n775_), .B0(new_new_n63_), .Y(new_new_n782_));
  NO2        g0760(.A(i_2_), .B(i_12_), .Y(new_new_n783_));
  OAI210     g0761(.A0(new_new_n664_), .A1(new_new_n388_), .B0(new_new_n783_), .Y(new_new_n784_));
  NA2        g0762(.A(i_8_), .B(new_new_n25_), .Y(new_new_n785_));
  NO3        g0763(.A(new_new_n785_), .B(new_new_n405_), .C(new_new_n654_), .Y(new_new_n786_));
  OAI210     g0764(.A0(new_new_n786_), .A1(new_new_n390_), .B0(new_new_n388_), .Y(new_new_n787_));
  NO2        g0765(.A(new_new_n126_), .B(i_2_), .Y(new_new_n788_));
  NA2        g0766(.A(new_new_n788_), .B(new_new_n690_), .Y(new_new_n789_));
  NA3        g0767(.A(new_new_n789_), .B(new_new_n787_), .C(new_new_n784_), .Y(new_new_n790_));
  NA3        g0768(.A(new_new_n790_), .B(new_new_n46_), .C(new_new_n230_), .Y(new_new_n791_));
  NA4        g0769(.A(new_new_n791_), .B(new_new_n782_), .C(new_new_n773_), .D(new_new_n758_), .Y(new_new_n792_));
  OR4        g0770(.A(new_new_n792_), .B(new_new_n750_), .C(new_new_n739_), .D(new_new_n672_), .Y(zz05));
  NA3        g0771(.A(new_new_n24_), .B(new_new_n783_), .C(new_new_n107_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n655_), .B(i_11_), .Y(new_new_n795_));
  OAI210     g0773(.A0(new_new_n659_), .A1(new_new_n88_), .B0(new_new_n795_), .Y(new_new_n796_));
  NA3        g0774(.A(new_new_n796_), .B(new_new_n794_), .C(new_new_n560_), .Y(new_new_n797_));
  NO3        g0775(.A(i_11_), .B(new_new_n242_), .C(i_13_), .Y(new_new_n798_));
  NO2        g0776(.A(new_new_n122_), .B(new_new_n23_), .Y(new_new_n799_));
  NA2        g0777(.A(i_12_), .B(i_8_), .Y(new_new_n800_));
  OAI210     g0778(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n800_), .Y(new_new_n801_));
  NA2        g0779(.A(new_new_n801_), .B(new_new_n799_), .Y(new_new_n802_));
  INV        g0780(.A(new_new_n802_), .Y(new_new_n803_));
  NO2        g0781(.A(new_new_n803_), .B(new_new_n797_), .Y(new_new_n804_));
  INV        g0782(.A(new_new_n171_), .Y(new_new_n805_));
  INV        g0783(.A(new_new_n251_), .Y(new_new_n806_));
  INV        g0784(.A(new_new_n476_), .Y(new_new_n807_));
  AOI210     g0785(.A0(new_new_n807_), .A1(new_new_n806_), .B0(new_new_n805_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n485_), .B(new_new_n26_), .Y(new_new_n809_));
  NO2        g0787(.A(new_new_n809_), .B(new_new_n444_), .Y(new_new_n810_));
  INV        g0788(.A(new_new_n808_), .Y(new_new_n811_));
  INV        g0789(.A(new_new_n172_), .Y(new_new_n812_));
  NO3        g0790(.A(new_new_n674_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n813_));
  AOI210     g0791(.A0(new_new_n812_), .A1(new_new_n88_), .B0(new_new_n813_), .Y(new_new_n814_));
  NO2        g0792(.A(new_new_n814_), .B(new_new_n194_), .Y(new_new_n815_));
  OA210      g0793(.A0(new_new_n675_), .A1(new_new_n124_), .B0(i_13_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n201_), .B(new_new_n204_), .Y(new_new_n817_));
  NA2        g0795(.A(new_new_n150_), .B(i_8_), .Y(new_new_n818_));
  AOI210     g0796(.A0(new_new_n818_), .A1(new_new_n817_), .B0(new_new_n393_), .Y(new_new_n819_));
  AOI210     g0797(.A0(new_new_n211_), .A1(new_new_n146_), .B0(new_new_n559_), .Y(new_new_n820_));
  OAI210     g0798(.A0(new_new_n820_), .A1(new_new_n231_), .B0(new_new_n444_), .Y(new_new_n821_));
  NO2        g0799(.A(new_new_n103_), .B(new_new_n45_), .Y(new_new_n822_));
  NA4        g0800(.A(new_new_n102_), .B(new_new_n317_), .C(new_new_n122_), .D(new_new_n43_), .Y(new_new_n823_));
  OAI210     g0801(.A0(new_new_n823_), .A1(new_new_n822_), .B0(new_new_n821_), .Y(new_new_n824_));
  NO4        g0802(.A(new_new_n824_), .B(new_new_n819_), .C(new_new_n816_), .D(new_new_n815_), .Y(new_new_n825_));
  NA2        g0803(.A(new_new_n625_), .B(new_new_n28_), .Y(new_new_n826_));
  NA2        g0804(.A(new_new_n798_), .B(new_new_n285_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n827_), .B(new_new_n826_), .Y(new_new_n828_));
  NO2        g0806(.A(new_new_n62_), .B(i_12_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n828_), .B(new_new_n47_), .Y(new_new_n830_));
  NA4        g0808(.A(new_new_n830_), .B(new_new_n825_), .C(new_new_n811_), .D(new_new_n804_), .Y(zz06));
  NO3        g0809(.A(new_new_n262_), .B(new_new_n319_), .C(i_1_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n186_), .B(new_new_n137_), .Y(new_new_n833_));
  OAI210     g0811(.A0(new_new_n833_), .A1(new_new_n832_), .B0(new_new_n788_), .Y(new_new_n834_));
  NA4        g0812(.A(new_new_n411_), .B(new_new_n517_), .C(new_new_n71_), .D(new_new_n102_), .Y(new_new_n835_));
  INV        g0813(.A(new_new_n835_), .Y(new_new_n836_));
  NO2        g0814(.A(new_new_n225_), .B(new_new_n522_), .Y(new_new_n837_));
  NO2        g0815(.A(i_11_), .B(i_9_), .Y(new_new_n838_));
  NO3        g0816(.A(new_new_n837_), .B(new_new_n836_), .C(new_new_n341_), .Y(new_new_n839_));
  AO210      g0817(.A0(new_new_n839_), .A1(new_new_n834_), .B0(i_12_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n394_), .B(new_new_n349_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n741_), .B(new_new_n71_), .Y(new_new_n842_));
  NA3        g0820(.A(new_new_n680_), .B(new_new_n842_), .C(new_new_n841_), .Y(new_new_n843_));
  INV        g0821(.A(new_new_n198_), .Y(new_new_n844_));
  AOI220     g0822(.A0(new_new_n844_), .A1(new_new_n838_), .B0(new_new_n843_), .B1(new_new_n73_), .Y(new_new_n845_));
  INV        g0823(.A(new_new_n340_), .Y(new_new_n846_));
  NA2        g0824(.A(new_new_n75_), .B(new_new_n129_), .Y(new_new_n847_));
  OAI210     g0825(.A0(new_new_n774_), .A1(i_5_), .B0(new_new_n122_), .Y(new_new_n848_));
  NA2        g0826(.A(new_new_n848_), .B(new_new_n47_), .Y(new_new_n849_));
  AOI210     g0827(.A0(new_new_n849_), .A1(new_new_n847_), .B0(new_new_n846_), .Y(new_new_n850_));
  NO3        g0828(.A(new_new_n258_), .B(new_new_n130_), .C(i_9_), .Y(new_new_n851_));
  NA2        g0829(.A(new_new_n851_), .B(new_new_n829_), .Y(new_new_n852_));
  AOI210     g0830(.A0(new_new_n852_), .A1(new_new_n557_), .B0(new_new_n186_), .Y(new_new_n853_));
  NO2        g0831(.A(new_new_n32_), .B(i_11_), .Y(new_new_n854_));
  NA3        g0832(.A(new_new_n854_), .B(new_new_n507_), .C(new_new_n411_), .Y(new_new_n855_));
  NAi32      g0833(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n856_));
  AOI210     g0834(.A0(new_new_n774_), .A1(new_new_n86_), .B0(new_new_n856_), .Y(new_new_n857_));
  OAI210     g0835(.A0(new_new_n740_), .A1(new_new_n613_), .B0(new_new_n612_), .Y(new_new_n858_));
  NAi31      g0836(.An(new_new_n857_), .B(new_new_n858_), .C(new_new_n855_), .Y(new_new_n859_));
  OR3        g0837(.A(new_new_n859_), .B(new_new_n853_), .C(new_new_n850_), .Y(new_new_n860_));
  NO2        g0838(.A(new_new_n751_), .B(i_2_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n862_));
  NA2        g0840(.A(new_new_n1120_), .B(new_new_n861_), .Y(new_new_n863_));
  AO220      g0841(.A0(new_new_n377_), .A1(new_new_n367_), .B0(new_new_n419_), .B1(i_8_), .Y(new_new_n864_));
  NA3        g0842(.A(new_new_n864_), .B(new_new_n263_), .C(i_7_), .Y(new_new_n865_));
  OR2        g0843(.A(new_new_n675_), .B(new_new_n476_), .Y(new_new_n866_));
  NA3        g0844(.A(new_new_n866_), .B(new_new_n145_), .C(new_new_n69_), .Y(new_new_n867_));
  NA3        g0845(.A(new_new_n867_), .B(new_new_n865_), .C(new_new_n863_), .Y(new_new_n868_));
  AOI220     g0846(.A0(new_new_n1123_), .A1(new_new_n612_), .B0(new_new_n837_), .B1(new_new_n769_), .Y(new_new_n869_));
  NA3        g0847(.A(new_new_n393_), .B(new_new_n244_), .C(new_new_n145_), .Y(new_new_n870_));
  OAI210     g0848(.A0(new_new_n419_), .A1(new_new_n205_), .B0(new_new_n70_), .Y(new_new_n871_));
  NA4        g0849(.A(new_new_n871_), .B(new_new_n870_), .C(new_new_n869_), .D(new_new_n658_), .Y(new_new_n872_));
  AO210      g0850(.A0(new_new_n559_), .A1(new_new_n47_), .B0(new_new_n87_), .Y(new_new_n873_));
  NA3        g0851(.A(new_new_n873_), .B(new_new_n518_), .C(new_new_n222_), .Y(new_new_n874_));
  AOI210     g0852(.A0(new_new_n476_), .A1(new_new_n474_), .B0(new_new_n611_), .Y(new_new_n875_));
  NO2        g0853(.A(i_10_), .B(new_new_n103_), .Y(new_new_n876_));
  OAI210     g0854(.A0(new_new_n876_), .A1(new_new_n110_), .B0(new_new_n431_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n250_), .B(new_new_n47_), .Y(new_new_n878_));
  NA2        g0856(.A(new_new_n878_), .B(new_new_n640_), .Y(new_new_n879_));
  NA3        g0857(.A(new_new_n879_), .B(new_new_n340_), .C(i_7_), .Y(new_new_n880_));
  NA4        g0858(.A(new_new_n880_), .B(new_new_n877_), .C(new_new_n875_), .D(new_new_n874_), .Y(new_new_n881_));
  NO4        g0859(.A(new_new_n881_), .B(new_new_n872_), .C(new_new_n868_), .D(new_new_n860_), .Y(new_new_n882_));
  NA4        g0860(.A(new_new_n882_), .B(new_new_n845_), .C(new_new_n840_), .D(new_new_n401_), .Y(zz03));
  NA2        g0861(.A(i_12_), .B(i_10_), .Y(new_new_n884_));
  NA2        g0862(.A(i_6_), .B(i_7_), .Y(new_new_n885_));
  NO2        g0863(.A(new_new_n885_), .B(i_0_), .Y(new_new_n886_));
  NO2        g0864(.A(i_11_), .B(new_new_n242_), .Y(new_new_n887_));
  OAI210     g0865(.A0(new_new_n886_), .A1(new_new_n300_), .B0(new_new_n887_), .Y(new_new_n888_));
  NO2        g0866(.A(new_new_n888_), .B(new_new_n194_), .Y(new_new_n889_));
  NO3        g0867(.A(new_new_n481_), .B(new_new_n90_), .C(new_new_n45_), .Y(new_new_n890_));
  OA210      g0868(.A0(new_new_n890_), .A1(new_new_n889_), .B0(new_new_n174_), .Y(new_new_n891_));
  NA3        g0869(.A(new_new_n870_), .B(new_new_n658_), .C(new_new_n392_), .Y(new_new_n892_));
  NA2        g0870(.A(new_new_n892_), .B(new_new_n40_), .Y(new_new_n893_));
  NOi21      g0871(.An(new_new_n97_), .B(new_new_n810_), .Y(new_new_n894_));
  NO3        g0872(.A(new_new_n685_), .B(new_new_n485_), .C(new_new_n129_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n433_), .B(new_new_n46_), .Y(new_new_n896_));
  AN2        g0874(.A(new_new_n483_), .B(new_new_n56_), .Y(new_new_n897_));
  NO3        g0875(.A(new_new_n897_), .B(new_new_n895_), .C(new_new_n894_), .Y(new_new_n898_));
  AOI210     g0876(.A0(new_new_n898_), .A1(new_new_n893_), .B0(new_new_n49_), .Y(new_new_n899_));
  NA2        g0877(.A(new_new_n186_), .B(new_new_n621_), .Y(new_new_n900_));
  NA2        g0878(.A(new_new_n761_), .B(new_new_n730_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n347_), .B(new_new_n464_), .Y(new_new_n902_));
  OAI220     g0880(.A0(new_new_n902_), .A1(new_new_n901_), .B0(new_new_n900_), .B1(new_new_n63_), .Y(new_new_n903_));
  NOi21      g0881(.An(i_5_), .B(i_9_), .Y(new_new_n904_));
  NA2        g0882(.A(new_new_n904_), .B(new_new_n472_), .Y(new_new_n905_));
  AOI210     g0883(.A0(new_new_n276_), .A1(new_new_n509_), .B0(new_new_n745_), .Y(new_new_n906_));
  NO3        g0884(.A(new_new_n436_), .B(new_new_n276_), .C(new_new_n73_), .Y(new_new_n907_));
  NO2        g0885(.A(new_new_n175_), .B(new_new_n146_), .Y(new_new_n908_));
  AOI210     g0886(.A0(new_new_n908_), .A1(new_new_n250_), .B0(new_new_n907_), .Y(new_new_n909_));
  OAI220     g0887(.A0(new_new_n909_), .A1(new_new_n181_), .B0(new_new_n906_), .B1(new_new_n905_), .Y(new_new_n910_));
  NO4        g0888(.A(new_new_n910_), .B(new_new_n903_), .C(new_new_n899_), .D(new_new_n891_), .Y(new_new_n911_));
  NOi21      g0889(.An(i_0_), .B(i_10_), .Y(new_new_n912_));
  NA2        g0890(.A(new_new_n186_), .B(new_new_n24_), .Y(new_new_n913_));
  NO2        g0891(.A(new_new_n728_), .B(new_new_n648_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n914_), .B(new_new_n913_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n324_), .B(new_new_n127_), .Y(new_new_n916_));
  NAi21      g0894(.An(new_new_n161_), .B(new_new_n464_), .Y(new_new_n917_));
  OAI220     g0895(.A0(new_new_n917_), .A1(new_new_n878_), .B0(new_new_n916_), .B1(new_new_n422_), .Y(new_new_n918_));
  NO2        g0896(.A(new_new_n918_), .B(new_new_n915_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n411_), .B(new_new_n304_), .Y(new_new_n920_));
  NA2        g0898(.A(new_new_n920_), .B(new_new_n764_), .Y(new_new_n921_));
  NA2        g0899(.A(new_new_n622_), .B(i_0_), .Y(new_new_n922_));
  NO3        g0900(.A(new_new_n922_), .B(new_new_n406_), .C(new_new_n88_), .Y(new_new_n923_));
  NO4        g0901(.A(new_new_n639_), .B(new_new_n219_), .C(new_new_n440_), .D(new_new_n432_), .Y(new_new_n924_));
  AOI210     g0902(.A0(new_new_n924_), .A1(i_11_), .B0(new_new_n923_), .Y(new_new_n925_));
  INV        g0903(.A(new_new_n507_), .Y(new_new_n926_));
  AN2        g0904(.A(new_new_n97_), .B(new_new_n249_), .Y(new_new_n927_));
  NA2        g0905(.A(new_new_n798_), .B(new_new_n341_), .Y(new_new_n928_));
  AOI210     g0906(.A0(new_new_n518_), .A1(new_new_n88_), .B0(new_new_n59_), .Y(new_new_n929_));
  OAI220     g0907(.A0(new_new_n929_), .A1(new_new_n928_), .B0(new_new_n713_), .B1(new_new_n581_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n260_), .B(new_new_n152_), .Y(new_new_n931_));
  NA2        g0909(.A(i_0_), .B(i_10_), .Y(new_new_n932_));
  OAI210     g0910(.A0(new_new_n932_), .A1(new_new_n85_), .B0(new_new_n584_), .Y(new_new_n933_));
  NO4        g0911(.A(new_new_n112_), .B(new_new_n59_), .C(new_new_n723_), .D(i_5_), .Y(new_new_n934_));
  AO220      g0912(.A0(new_new_n934_), .A1(new_new_n933_), .B0(new_new_n931_), .B1(i_6_), .Y(new_new_n935_));
  AOI220     g0913(.A0(new_new_n347_), .A1(new_new_n99_), .B0(new_new_n186_), .B1(new_new_n83_), .Y(new_new_n936_));
  NA2        g0914(.A(new_new_n616_), .B(i_4_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n189_), .B(new_new_n204_), .Y(new_new_n938_));
  OAI220     g0916(.A0(new_new_n938_), .A1(new_new_n928_), .B0(new_new_n937_), .B1(new_new_n936_), .Y(new_new_n939_));
  NO4        g0917(.A(new_new_n939_), .B(new_new_n935_), .C(new_new_n930_), .D(new_new_n927_), .Y(new_new_n940_));
  NA4        g0918(.A(new_new_n940_), .B(new_new_n925_), .C(new_new_n921_), .D(new_new_n919_), .Y(new_new_n941_));
  NA2        g0919(.A(i_11_), .B(i_9_), .Y(new_new_n942_));
  NO3        g0920(.A(i_12_), .B(new_new_n942_), .C(new_new_n657_), .Y(new_new_n943_));
  AO220      g0921(.A0(new_new_n943_), .A1(i_10_), .B0(new_new_n278_), .B1(new_new_n87_), .Y(new_new_n944_));
  NO2        g0922(.A(new_new_n49_), .B(i_7_), .Y(new_new_n945_));
  NAi31      g0923(.An(new_new_n273_), .B(new_new_n490_), .C(new_new_n159_), .Y(new_new_n946_));
  NO2        g0924(.A(new_new_n942_), .B(new_new_n73_), .Y(new_new_n947_));
  NO2        g0925(.A(new_new_n175_), .B(i_0_), .Y(new_new_n948_));
  INV        g0926(.A(new_new_n948_), .Y(new_new_n949_));
  NA2        g0927(.A(new_new_n507_), .B(new_new_n236_), .Y(new_new_n950_));
  AOI210     g0928(.A0(new_new_n391_), .A1(new_new_n42_), .B0(new_new_n430_), .Y(new_new_n951_));
  OAI220     g0929(.A0(new_new_n951_), .A1(new_new_n905_), .B0(new_new_n950_), .B1(new_new_n949_), .Y(new_new_n952_));
  NO3        g0930(.A(new_new_n952_), .B(new_new_n946_), .C(new_new_n944_), .Y(new_new_n953_));
  NA2        g0931(.A(new_new_n712_), .B(new_new_n119_), .Y(new_new_n954_));
  NO2        g0932(.A(i_6_), .B(new_new_n954_), .Y(new_new_n955_));
  AOI210     g0933(.A0(new_new_n475_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n956_));
  NA2        g0934(.A(new_new_n171_), .B(new_new_n104_), .Y(new_new_n957_));
  NOi32      g0935(.An(new_new_n956_), .Bn(new_new_n189_), .C(new_new_n957_), .Y(new_new_n958_));
  AOI210     g0936(.A0(new_new_n659_), .A1(new_new_n341_), .B0(new_new_n249_), .Y(new_new_n959_));
  NO2        g0937(.A(new_new_n959_), .B(new_new_n896_), .Y(new_new_n960_));
  NO3        g0938(.A(new_new_n960_), .B(new_new_n958_), .C(new_new_n955_), .Y(new_new_n961_));
  NOi21      g0939(.An(i_7_), .B(i_5_), .Y(new_new_n962_));
  NOi31      g0940(.An(new_new_n962_), .B(new_new_n912_), .C(new_new_n777_), .Y(new_new_n963_));
  NA3        g0941(.A(new_new_n963_), .B(new_new_n405_), .C(i_6_), .Y(new_new_n964_));
  OA210      g0942(.A0(new_new_n957_), .A1(new_new_n557_), .B0(new_new_n964_), .Y(new_new_n965_));
  NO3        g0943(.A(new_new_n425_), .B(new_new_n380_), .C(new_new_n376_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n270_), .B(new_new_n330_), .Y(new_new_n967_));
  NO2        g0945(.A(new_new_n777_), .B(new_new_n265_), .Y(new_new_n968_));
  AOI210     g0946(.A0(new_new_n968_), .A1(new_new_n967_), .B0(new_new_n966_), .Y(new_new_n969_));
  NA4        g0947(.A(new_new_n969_), .B(new_new_n965_), .C(new_new_n961_), .D(new_new_n953_), .Y(new_new_n970_));
  NO2        g0948(.A(new_new_n913_), .B(new_new_n245_), .Y(new_new_n971_));
  AN2        g0949(.A(new_new_n346_), .B(new_new_n341_), .Y(new_new_n972_));
  AO220      g0950(.A0(new_new_n972_), .A1(new_new_n908_), .B0(new_new_n362_), .B1(new_new_n27_), .Y(new_new_n973_));
  OAI210     g0951(.A0(new_new_n973_), .A1(new_new_n971_), .B0(i_10_), .Y(new_new_n974_));
  NO2        g0952(.A(new_new_n884_), .B(new_new_n329_), .Y(new_new_n975_));
  OA210      g0953(.A0(new_new_n507_), .A1(new_new_n228_), .B0(new_new_n506_), .Y(new_new_n976_));
  OAI210     g0954(.A0(new_new_n976_), .A1(new_new_n975_), .B0(new_new_n947_), .Y(new_new_n977_));
  NA3        g0955(.A(new_new_n506_), .B(new_new_n433_), .C(new_new_n46_), .Y(new_new_n978_));
  OAI210     g0956(.A0(new_new_n917_), .A1(new_new_n926_), .B0(new_new_n978_), .Y(new_new_n979_));
  NO2        g0957(.A(new_new_n263_), .B(new_new_n47_), .Y(new_new_n980_));
  NA2        g0958(.A(new_new_n947_), .B(new_new_n317_), .Y(new_new_n981_));
  OAI210     g0959(.A0(new_new_n980_), .A1(new_new_n188_), .B0(new_new_n981_), .Y(new_new_n982_));
  AOI220     g0960(.A0(new_new_n982_), .A1(new_new_n507_), .B0(new_new_n979_), .B1(new_new_n73_), .Y(new_new_n983_));
  NA3        g0961(.A(new_new_n862_), .B(new_new_n403_), .C(i_12_), .Y(new_new_n984_));
  NA2        g0962(.A(new_new_n93_), .B(new_new_n45_), .Y(new_new_n985_));
  NO2        g0963(.A(new_new_n75_), .B(new_new_n800_), .Y(new_new_n986_));
  AOI220     g0964(.A0(new_new_n986_), .A1(new_new_n985_), .B0(new_new_n174_), .B1(new_new_n648_), .Y(new_new_n987_));
  AOI210     g0965(.A0(new_new_n987_), .A1(new_new_n984_), .B0(new_new_n48_), .Y(new_new_n988_));
  NO3        g0966(.A(new_new_n639_), .B(new_new_n375_), .C(new_new_n24_), .Y(new_new_n989_));
  AOI210     g0967(.A0(new_new_n755_), .A1(new_new_n593_), .B0(new_new_n989_), .Y(new_new_n990_));
  NAi21      g0968(.An(i_9_), .B(i_5_), .Y(new_new_n991_));
  NO2        g0969(.A(new_new_n991_), .B(new_new_n425_), .Y(new_new_n992_));
  NO2        g0970(.A(new_new_n653_), .B(new_new_n106_), .Y(new_new_n993_));
  AOI220     g0971(.A0(new_new_n993_), .A1(i_0_), .B0(new_new_n992_), .B1(new_new_n675_), .Y(new_new_n994_));
  OAI220     g0972(.A0(new_new_n994_), .A1(new_new_n85_), .B0(new_new_n990_), .B1(new_new_n172_), .Y(new_new_n995_));
  NO3        g0973(.A(new_new_n995_), .B(new_new_n988_), .C(new_new_n561_), .Y(new_new_n996_));
  NA4        g0974(.A(new_new_n996_), .B(new_new_n983_), .C(new_new_n977_), .D(new_new_n974_), .Y(new_new_n997_));
  NO3        g0975(.A(new_new_n997_), .B(new_new_n970_), .C(new_new_n941_), .Y(new_new_n998_));
  NO2        g0976(.A(new_new_n912_), .B(new_new_n777_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n1000_));
  NO3        g0978(.A(new_new_n106_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n1001_));
  AO220      g0979(.A0(new_new_n1001_), .A1(new_new_n73_), .B0(new_new_n999_), .B1(new_new_n174_), .Y(new_new_n1002_));
  NO2        g0980(.A(new_new_n743_), .B(new_new_n957_), .Y(new_new_n1003_));
  AOI210     g0981(.A0(new_new_n1002_), .A1(new_new_n364_), .B0(new_new_n1003_), .Y(new_new_n1004_));
  NA2        g0982(.A(new_new_n788_), .B(new_new_n144_), .Y(new_new_n1005_));
  INV        g0983(.A(new_new_n1005_), .Y(new_new_n1006_));
  NA3        g0984(.A(new_new_n1006_), .B(new_new_n730_), .C(new_new_n73_), .Y(new_new_n1007_));
  NO2        g0985(.A(new_new_n858_), .B(new_new_n425_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n886_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n1009_));
  NA2        g0987(.A(new_new_n887_), .B(i_9_), .Y(new_new_n1010_));
  AOI210     g0988(.A0(new_new_n1009_), .A1(new_new_n534_), .B0(new_new_n1010_), .Y(new_new_n1011_));
  OAI210     g0989(.A0(new_new_n250_), .A1(i_9_), .B0(new_new_n235_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n1012_), .A1(new_new_n922_), .B0(new_new_n152_), .Y(new_new_n1013_));
  NO3        g0991(.A(new_new_n1013_), .B(new_new_n1011_), .C(new_new_n1008_), .Y(new_new_n1014_));
  NA3        g0992(.A(new_new_n1014_), .B(new_new_n1007_), .C(new_new_n1004_), .Y(new_new_n1015_));
  NA2        g0993(.A(new_new_n972_), .B(new_new_n393_), .Y(new_new_n1016_));
  AOI210     g0994(.A0(new_new_n311_), .A1(new_new_n161_), .B0(new_new_n1016_), .Y(new_new_n1017_));
  NA3        g0995(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n1018_));
  NA2        g0996(.A(new_new_n945_), .B(new_new_n523_), .Y(new_new_n1019_));
  AOI210     g0997(.A0(new_new_n1018_), .A1(new_new_n161_), .B0(new_new_n1019_), .Y(new_new_n1020_));
  NO2        g0998(.A(new_new_n1020_), .B(new_new_n1017_), .Y(new_new_n1021_));
  NO3        g0999(.A(new_new_n932_), .B(new_new_n904_), .C(new_new_n191_), .Y(new_new_n1022_));
  AOI220     g1000(.A0(new_new_n1022_), .A1(i_11_), .B0(new_new_n617_), .B1(new_new_n75_), .Y(new_new_n1023_));
  NO3        g1001(.A(new_new_n213_), .B(new_new_n404_), .C(i_0_), .Y(new_new_n1024_));
  OAI210     g1002(.A0(new_new_n1024_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n1025_));
  INV        g1003(.A(new_new_n222_), .Y(new_new_n1026_));
  OAI220     g1004(.A0(new_new_n574_), .A1(new_new_n137_), .B0(new_new_n699_), .B1(new_new_n669_), .Y(new_new_n1027_));
  NA3        g1005(.A(new_new_n1027_), .B(new_new_n420_), .C(new_new_n1026_), .Y(new_new_n1028_));
  NA4        g1006(.A(new_new_n1028_), .B(new_new_n1025_), .C(new_new_n1023_), .D(new_new_n1021_), .Y(new_new_n1029_));
  NO2        g1007(.A(new_new_n248_), .B(new_new_n93_), .Y(new_new_n1030_));
  AOI210     g1008(.A0(new_new_n1030_), .A1(new_new_n999_), .B0(new_new_n108_), .Y(new_new_n1031_));
  AOI220     g1009(.A0(new_new_n962_), .A1(new_new_n523_), .B0(new_new_n886_), .B1(new_new_n162_), .Y(new_new_n1032_));
  NA2        g1010(.A(new_new_n367_), .B(new_new_n176_), .Y(new_new_n1033_));
  OA220      g1011(.A0(new_new_n1033_), .A1(new_new_n1032_), .B0(new_new_n1031_), .B1(i_5_), .Y(new_new_n1034_));
  AOI210     g1012(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n175_), .Y(new_new_n1035_));
  NA2        g1013(.A(new_new_n1035_), .B(new_new_n976_), .Y(new_new_n1036_));
  NA3        g1014(.A(new_new_n666_), .B(new_new_n186_), .C(new_new_n83_), .Y(new_new_n1037_));
  NA2        g1015(.A(new_new_n1037_), .B(new_new_n591_), .Y(new_new_n1038_));
  NO3        g1016(.A(new_new_n896_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n1039_));
  NA2        g1017(.A(new_new_n521_), .B(new_new_n504_), .Y(new_new_n1040_));
  NO3        g1018(.A(new_new_n1040_), .B(new_new_n1039_), .C(new_new_n1038_), .Y(new_new_n1041_));
  NA3        g1019(.A(new_new_n945_), .B(new_new_n300_), .C(new_new_n235_), .Y(new_new_n1042_));
  INV        g1020(.A(new_new_n1042_), .Y(new_new_n1043_));
  NA3        g1021(.A(new_new_n411_), .B(new_new_n348_), .C(new_new_n226_), .Y(new_new_n1044_));
  OAI210     g1022(.A0(new_new_n900_), .A1(new_new_n703_), .B0(new_new_n1044_), .Y(new_new_n1045_));
  NOi31      g1023(.An(new_new_n410_), .B(new_new_n1000_), .C(new_new_n245_), .Y(new_new_n1046_));
  NO3        g1024(.A(new_new_n942_), .B(new_new_n222_), .C(new_new_n191_), .Y(new_new_n1047_));
  NO4        g1025(.A(new_new_n1047_), .B(new_new_n1046_), .C(new_new_n1045_), .D(new_new_n1043_), .Y(new_new_n1048_));
  NA4        g1026(.A(new_new_n1048_), .B(new_new_n1041_), .C(new_new_n1036_), .D(new_new_n1034_), .Y(new_new_n1049_));
  AOI210     g1027(.A0(new_new_n616_), .A1(new_new_n573_), .B0(new_new_n668_), .Y(new_new_n1050_));
  NO3        g1028(.A(new_new_n1050_), .B(new_new_n607_), .C(new_new_n361_), .Y(new_new_n1051_));
  NA3        g1029(.A(new_new_n887_), .B(new_new_n109_), .C(new_new_n122_), .Y(new_new_n1052_));
  INV        g1030(.A(new_new_n1052_), .Y(new_new_n1053_));
  AOI210     g1031(.A0(new_new_n1053_), .A1(new_new_n1124_), .B0(new_new_n1051_), .Y(new_new_n1054_));
  NA3        g1032(.A(new_new_n317_), .B(i_5_), .C(new_new_n194_), .Y(new_new_n1055_));
  NAi31      g1033(.An(new_new_n247_), .B(new_new_n1055_), .C(new_new_n248_), .Y(new_new_n1056_));
  NO4        g1034(.A(new_new_n245_), .B(new_new_n213_), .C(i_0_), .D(i_12_), .Y(new_new_n1057_));
  AOI220     g1035(.A0(new_new_n1057_), .A1(new_new_n1056_), .B0(new_new_n836_), .B1(new_new_n176_), .Y(new_new_n1058_));
  AN2        g1036(.A(new_new_n932_), .B(new_new_n152_), .Y(new_new_n1059_));
  NO4        g1037(.A(new_new_n1059_), .B(i_12_), .C(new_new_n703_), .D(new_new_n129_), .Y(new_new_n1060_));
  NA2        g1038(.A(new_new_n1060_), .B(new_new_n222_), .Y(new_new_n1061_));
  NA3        g1039(.A(new_new_n99_), .B(new_new_n621_), .C(i_11_), .Y(new_new_n1062_));
  NO2        g1040(.A(new_new_n1062_), .B(new_new_n154_), .Y(new_new_n1063_));
  NA2        g1041(.A(new_new_n962_), .B(new_new_n503_), .Y(new_new_n1064_));
  OAI220     g1042(.A0(i_7_), .A1(new_new_n1055_), .B0(new_new_n1064_), .B1(new_new_n731_), .Y(new_new_n1065_));
  AOI210     g1043(.A0(new_new_n1065_), .A1(new_new_n948_), .B0(new_new_n1063_), .Y(new_new_n1066_));
  NA4        g1044(.A(new_new_n1066_), .B(new_new_n1061_), .C(new_new_n1058_), .D(new_new_n1054_), .Y(new_new_n1067_));
  NO4        g1045(.A(new_new_n1067_), .B(new_new_n1049_), .C(new_new_n1029_), .D(new_new_n1015_), .Y(new_new_n1068_));
  OAI210     g1046(.A0(new_new_n861_), .A1(new_new_n854_), .B0(new_new_n37_), .Y(new_new_n1069_));
  NA3        g1047(.A(new_new_n956_), .B(new_new_n388_), .C(i_5_), .Y(new_new_n1070_));
  NA3        g1048(.A(new_new_n1070_), .B(new_new_n1069_), .C(new_new_n665_), .Y(new_new_n1071_));
  NA2        g1049(.A(new_new_n1071_), .B(new_new_n209_), .Y(new_new_n1072_));
  AN2        g1050(.A(new_new_n751_), .B(new_new_n389_), .Y(new_new_n1073_));
  NA2        g1051(.A(new_new_n187_), .B(new_new_n189_), .Y(new_new_n1074_));
  AO210      g1052(.A0(new_new_n1073_), .A1(new_new_n33_), .B0(new_new_n1074_), .Y(new_new_n1075_));
  OAI210     g1053(.A0(new_new_n668_), .A1(new_new_n666_), .B0(new_new_n329_), .Y(new_new_n1076_));
  NAi31      g1054(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1077_));
  AOI210     g1055(.A0(new_new_n115_), .A1(new_new_n70_), .B0(new_new_n1077_), .Y(new_new_n1078_));
  NO2        g1056(.A(new_new_n1078_), .B(new_new_n700_), .Y(new_new_n1079_));
  NA3        g1057(.A(new_new_n1079_), .B(new_new_n1076_), .C(new_new_n1075_), .Y(new_new_n1080_));
  NO2        g1058(.A(new_new_n493_), .B(new_new_n276_), .Y(new_new_n1081_));
  NO4        g1059(.A(new_new_n238_), .B(new_new_n143_), .C(new_new_n734_), .D(new_new_n37_), .Y(new_new_n1082_));
  NO3        g1060(.A(new_new_n1082_), .B(new_new_n1081_), .C(new_new_n924_), .Y(new_new_n1083_));
  OAI210     g1061(.A0(new_new_n1062_), .A1(new_new_n146_), .B0(new_new_n1083_), .Y(new_new_n1084_));
  AOI210     g1062(.A0(new_new_n1080_), .A1(new_new_n49_), .B0(new_new_n1084_), .Y(new_new_n1085_));
  AOI210     g1063(.A0(new_new_n1085_), .A1(new_new_n1072_), .B0(new_new_n73_), .Y(new_new_n1086_));
  NO2        g1064(.A(new_new_n614_), .B(new_new_n400_), .Y(new_new_n1087_));
  NO2        g1065(.A(new_new_n1087_), .B(new_new_n805_), .Y(new_new_n1088_));
  OAI210     g1066(.A0(new_new_n80_), .A1(new_new_n55_), .B0(new_new_n107_), .Y(new_new_n1089_));
  NA2        g1067(.A(new_new_n1089_), .B(new_new_n76_), .Y(new_new_n1090_));
  AOI210     g1068(.A0(new_new_n1035_), .A1(new_new_n945_), .B0(new_new_n963_), .Y(new_new_n1091_));
  AOI210     g1069(.A0(new_new_n1091_), .A1(new_new_n1090_), .B0(new_new_n734_), .Y(new_new_n1092_));
  NA2        g1070(.A(new_new_n270_), .B(new_new_n58_), .Y(new_new_n1093_));
  AOI220     g1071(.A0(new_new_n1093_), .A1(new_new_n76_), .B0(new_new_n362_), .B1(new_new_n262_), .Y(new_new_n1094_));
  NO2        g1072(.A(new_new_n1094_), .B(new_new_n242_), .Y(new_new_n1095_));
  NA3        g1073(.A(new_new_n97_), .B(new_new_n319_), .C(new_new_n31_), .Y(new_new_n1096_));
  INV        g1074(.A(new_new_n1096_), .Y(new_new_n1097_));
  NO3        g1075(.A(new_new_n1097_), .B(new_new_n1095_), .C(new_new_n1092_), .Y(new_new_n1098_));
  OAI210     g1076(.A0(new_new_n278_), .A1(new_new_n157_), .B0(new_new_n88_), .Y(new_new_n1099_));
  NA3        g1077(.A(new_new_n809_), .B(new_new_n300_), .C(new_new_n80_), .Y(new_new_n1100_));
  AOI210     g1078(.A0(new_new_n1100_), .A1(new_new_n1099_), .B0(i_11_), .Y(new_new_n1101_));
  NA2        g1079(.A(new_new_n660_), .B(new_new_n219_), .Y(new_new_n1102_));
  OAI210     g1080(.A0(new_new_n1102_), .A1(new_new_n956_), .B0(new_new_n209_), .Y(new_new_n1103_));
  NA2        g1081(.A(new_new_n163_), .B(i_5_), .Y(new_new_n1104_));
  AOI210     g1082(.A0(new_new_n1103_), .A1(new_new_n817_), .B0(new_new_n1104_), .Y(new_new_n1105_));
  NO3        g1083(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n1106_));
  OAI210     g1084(.A0(new_new_n967_), .A1(new_new_n319_), .B0(new_new_n1106_), .Y(new_new_n1107_));
  NO2        g1085(.A(new_new_n1107_), .B(new_new_n777_), .Y(new_new_n1108_));
  NO4        g1086(.A(new_new_n991_), .B(new_new_n511_), .C(new_new_n259_), .D(new_new_n258_), .Y(new_new_n1109_));
  NO2        g1087(.A(new_new_n1109_), .B(new_new_n611_), .Y(new_new_n1110_));
  NO2        g1088(.A(new_new_n857_), .B(new_new_n381_), .Y(new_new_n1111_));
  AOI210     g1089(.A0(new_new_n1111_), .A1(new_new_n1110_), .B0(new_new_n41_), .Y(new_new_n1112_));
  NO4        g1090(.A(new_new_n1112_), .B(new_new_n1108_), .C(new_new_n1105_), .D(new_new_n1101_), .Y(new_new_n1113_));
  OAI210     g1091(.A0(new_new_n1098_), .A1(i_4_), .B0(new_new_n1113_), .Y(new_new_n1114_));
  NO3        g1092(.A(new_new_n1114_), .B(new_new_n1088_), .C(new_new_n1086_), .Y(new_new_n1115_));
  NA4        g1093(.A(new_new_n1115_), .B(new_new_n1068_), .C(new_new_n998_), .D(new_new_n911_), .Y(zz04));
  INV        g1094(.A(i_5_), .Y(new_new_n1119_));
  INV        g1095(.A(new_new_n862_), .Y(new_new_n1120_));
  INV        g1096(.A(new_new_n199_), .Y(new_new_n1121_));
  INV        g1097(.A(i_1_), .Y(new_new_n1122_));
  INV        g1098(.A(new_new_n86_), .Y(new_new_n1123_));
  INV        g1099(.A(i_5_), .Y(new_new_n1124_));
  INV        g1100(.A(new_new_n407_), .Y(new_new_n1125_));
  INV        g1101(.A(i_1_), .Y(new_new_n1126_));
endmodule


