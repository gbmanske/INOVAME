library verilog;
use verilog.vl_types.all;
entity tb_mult is
end tb_mult;
