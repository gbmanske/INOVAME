// Benchmark "top" written by ABC on Fri Jun 21 17:49:26 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n141_, new_new_n143_,
    new_new_n144_, new_new_n145_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1007_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g021(.A(new_new_n35_), .Y(mai1));
  INV        g022(.A(i_11_), .Y(new_new_n45_));
  NO2        g023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g024(.A(i_2_), .Y(new_new_n47_));
  NA2        g025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g026(.A(i_5_), .Y(new_new_n49_));
  NO2        g027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g041(.A(i_1_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g064(.A(i_6_), .Y(new_new_n87_));
  OR4        g065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  NO2        g068(.A(new_new_n89_), .B(new_new_n90_), .Y(new_new_n91_));
  OAI210     g069(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n91_), .Y(new_new_n92_));
  NAi21      g070(.An(i_6_), .B(i_10_), .Y(new_new_n93_));
  NA2        g071(.A(i_6_), .B(i_9_), .Y(new_new_n94_));
  AOI210     g072(.A0(new_new_n94_), .A1(new_new_n93_), .B0(new_new_n64_), .Y(new_new_n95_));
  NA2        g073(.A(i_2_), .B(i_6_), .Y(new_new_n96_));
  NO3        g074(.A(new_new_n96_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n97_));
  NO2        g075(.A(new_new_n97_), .B(new_new_n95_), .Y(new_new_n98_));
  AOI210     g076(.A0(new_new_n98_), .A1(new_new_n92_), .B0(new_new_n81_), .Y(new_new_n99_));
  AN3        g077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n100_));
  NAi21      g078(.An(i_6_), .B(i_11_), .Y(new_new_n101_));
  NO2        g079(.A(i_5_), .B(i_8_), .Y(new_new_n102_));
  NOi21      g080(.An(new_new_n102_), .B(new_new_n101_), .Y(new_new_n103_));
  AOI220     g081(.A0(new_new_n103_), .A1(new_new_n63_), .B0(new_new_n100_), .B1(new_new_n32_), .Y(new_new_n104_));
  INV        g082(.A(i_7_), .Y(new_new_n105_));
  NA2        g083(.A(new_new_n47_), .B(new_new_n105_), .Y(new_new_n106_));
  NO2        g084(.A(i_0_), .B(i_5_), .Y(new_new_n107_));
  NO2        g085(.A(new_new_n107_), .B(new_new_n87_), .Y(new_new_n108_));
  NA2        g086(.A(i_12_), .B(i_3_), .Y(new_new_n109_));
  INV        g087(.A(new_new_n109_), .Y(new_new_n110_));
  NA3        g088(.A(new_new_n110_), .B(new_new_n108_), .C(new_new_n106_), .Y(new_new_n111_));
  NAi21      g089(.An(i_7_), .B(i_11_), .Y(new_new_n112_));
  NO3        g090(.A(new_new_n112_), .B(new_new_n93_), .C(new_new_n54_), .Y(new_new_n113_));
  AN2        g091(.A(i_2_), .B(i_10_), .Y(new_new_n114_));
  NO2        g092(.A(new_new_n114_), .B(i_7_), .Y(new_new_n115_));
  OR2        g093(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n116_));
  NO2        g094(.A(i_8_), .B(new_new_n105_), .Y(new_new_n117_));
  NO3        g095(.A(new_new_n117_), .B(new_new_n116_), .C(new_new_n115_), .Y(new_new_n118_));
  NA2        g096(.A(i_12_), .B(i_7_), .Y(new_new_n119_));
  NO2        g097(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(i_0_), .Y(new_new_n121_));
  NA2        g099(.A(i_11_), .B(i_12_), .Y(new_new_n122_));
  OAI210     g100(.A0(new_new_n121_), .A1(new_new_n119_), .B0(new_new_n122_), .Y(new_new_n123_));
  NO2        g101(.A(new_new_n123_), .B(new_new_n118_), .Y(new_new_n124_));
  NAi41      g102(.An(new_new_n113_), .B(new_new_n124_), .C(new_new_n111_), .D(new_new_n104_), .Y(new_new_n125_));
  NOi21      g103(.An(i_1_), .B(i_5_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(i_11_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n128_));
  NA2        g106(.A(i_7_), .B(new_new_n25_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n129_), .B(new_new_n128_), .Y(new_new_n130_));
  NO2        g108(.A(new_new_n130_), .B(new_new_n47_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n94_), .B(new_new_n93_), .Y(new_new_n132_));
  NAi21      g110(.An(i_3_), .B(i_8_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(new_new_n63_), .Y(new_new_n134_));
  NOi31      g112(.An(new_new_n134_), .B(new_new_n132_), .C(new_new_n131_), .Y(new_new_n135_));
  NO2        g113(.A(i_1_), .B(new_new_n87_), .Y(new_new_n136_));
  NO2        g114(.A(i_6_), .B(i_5_), .Y(new_new_n137_));
  NA2        g115(.A(new_new_n137_), .B(i_3_), .Y(new_new_n138_));
  AO210      g116(.A0(new_new_n138_), .A1(new_new_n48_), .B0(new_new_n136_), .Y(new_new_n139_));
  OAI220     g117(.A0(new_new_n139_), .A1(new_new_n112_), .B0(new_new_n135_), .B1(new_new_n127_), .Y(new_new_n140_));
  NO3        g118(.A(new_new_n140_), .B(new_new_n125_), .C(new_new_n99_), .Y(new_new_n141_));
  NA3        g119(.A(new_new_n141_), .B(new_new_n80_), .C(new_new_n57_), .Y(mai2));
  NO2        g120(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n143_));
  NA2        g121(.A(i_6_), .B(new_new_n25_), .Y(new_new_n144_));
  NA2        g122(.A(new_new_n144_), .B(new_new_n143_), .Y(new_new_n145_));
  NA4        g123(.A(new_new_n145_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(mai0));
  AN2        g124(.A(i_8_), .B(i_7_), .Y(new_new_n147_));
  NA2        g125(.A(new_new_n147_), .B(i_6_), .Y(new_new_n148_));
  NO2        g126(.A(i_12_), .B(i_13_), .Y(new_new_n149_));
  NAi21      g127(.An(i_5_), .B(i_11_), .Y(new_new_n150_));
  NOi21      g128(.An(new_new_n149_), .B(new_new_n150_), .Y(new_new_n151_));
  NO2        g129(.A(i_0_), .B(i_1_), .Y(new_new_n152_));
  NA2        g130(.A(i_2_), .B(i_3_), .Y(new_new_n153_));
  NO2        g131(.A(new_new_n153_), .B(i_4_), .Y(new_new_n154_));
  NA3        g132(.A(new_new_n154_), .B(new_new_n152_), .C(new_new_n151_), .Y(new_new_n155_));
  OR2        g133(.A(new_new_n155_), .B(new_new_n25_), .Y(new_new_n156_));
  AN2        g134(.A(new_new_n149_), .B(new_new_n84_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n157_), .B(new_new_n27_), .Y(new_new_n158_));
  NA2        g136(.A(i_1_), .B(i_5_), .Y(new_new_n159_));
  NO2        g137(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n160_));
  NA2        g138(.A(new_new_n160_), .B(new_new_n36_), .Y(new_new_n161_));
  NO3        g139(.A(new_new_n161_), .B(new_new_n159_), .C(new_new_n158_), .Y(new_new_n162_));
  OR2        g140(.A(i_0_), .B(i_1_), .Y(new_new_n163_));
  NAi32      g141(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n164_));
  NOi21      g142(.An(i_4_), .B(i_10_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n40_), .Y(new_new_n166_));
  NO2        g144(.A(i_3_), .B(i_5_), .Y(new_new_n167_));
  INV        g145(.A(new_new_n162_), .Y(new_new_n168_));
  AOI210     g146(.A0(new_new_n168_), .A1(new_new_n156_), .B0(new_new_n148_), .Y(new_new_n169_));
  NA3        g147(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n170_));
  NA2        g148(.A(i_3_), .B(new_new_n49_), .Y(new_new_n171_));
  NOi21      g149(.An(i_4_), .B(i_9_), .Y(new_new_n172_));
  NOi21      g150(.An(i_11_), .B(i_13_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(new_new_n172_), .Y(new_new_n174_));
  OR2        g152(.A(new_new_n174_), .B(new_new_n171_), .Y(new_new_n175_));
  NO2        g153(.A(i_4_), .B(i_5_), .Y(new_new_n176_));
  NAi21      g154(.An(i_12_), .B(i_11_), .Y(new_new_n177_));
  NO2        g155(.A(new_new_n177_), .B(i_13_), .Y(new_new_n178_));
  NA3        g156(.A(new_new_n178_), .B(new_new_n176_), .C(new_new_n84_), .Y(new_new_n179_));
  AOI210     g157(.A0(new_new_n179_), .A1(new_new_n175_), .B0(new_new_n170_), .Y(new_new_n180_));
  NO2        g158(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n181_));
  NA2        g159(.A(new_new_n181_), .B(new_new_n47_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n36_), .B(i_5_), .Y(new_new_n183_));
  NA2        g161(.A(i_3_), .B(i_5_), .Y(new_new_n184_));
  NO2        g162(.A(new_new_n74_), .B(i_5_), .Y(new_new_n185_));
  NO2        g163(.A(i_13_), .B(i_10_), .Y(new_new_n186_));
  NA3        g164(.A(new_new_n186_), .B(new_new_n185_), .C(new_new_n45_), .Y(new_new_n187_));
  NO2        g165(.A(i_2_), .B(i_1_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n188_), .B(i_3_), .Y(new_new_n189_));
  NAi21      g167(.An(i_4_), .B(i_12_), .Y(new_new_n190_));
  NO4        g168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n187_), .D(new_new_n25_), .Y(new_new_n191_));
  NO2        g169(.A(new_new_n191_), .B(new_new_n180_), .Y(new_new_n192_));
  INV        g170(.A(i_8_), .Y(new_new_n193_));
  NO3        g171(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n194_));
  NA2        g172(.A(new_new_n194_), .B(new_new_n117_), .Y(new_new_n195_));
  NO3        g173(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n196_));
  NA3        g174(.A(new_new_n196_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n197_));
  NO3        g175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n198_));
  OAI210     g176(.A0(new_new_n100_), .A1(i_12_), .B0(new_new_n198_), .Y(new_new_n199_));
  AOI210     g177(.A0(new_new_n199_), .A1(new_new_n197_), .B0(new_new_n195_), .Y(new_new_n200_));
  NO2        g178(.A(i_3_), .B(i_8_), .Y(new_new_n201_));
  NO3        g179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n202_));
  NO2        g180(.A(new_new_n107_), .B(new_new_n59_), .Y(new_new_n203_));
  NO2        g181(.A(i_13_), .B(i_9_), .Y(new_new_n204_));
  NA3        g182(.A(new_new_n204_), .B(i_6_), .C(new_new_n193_), .Y(new_new_n205_));
  NAi21      g183(.An(i_12_), .B(i_3_), .Y(new_new_n206_));
  OR2        g184(.A(new_new_n206_), .B(new_new_n205_), .Y(new_new_n207_));
  NO2        g185(.A(new_new_n45_), .B(i_5_), .Y(new_new_n208_));
  NO3        g186(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n209_));
  NA2        g187(.A(new_new_n209_), .B(new_new_n208_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n210_), .B(new_new_n207_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n211_), .B(new_new_n200_), .Y(new_new_n212_));
  OAI220     g190(.A0(new_new_n212_), .A1(i_4_), .B0(i_7_), .B1(new_new_n192_), .Y(new_new_n213_));
  NAi21      g191(.An(i_12_), .B(i_7_), .Y(new_new_n214_));
  NA3        g192(.A(i_13_), .B(new_new_n193_), .C(i_10_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n216_));
  NA2        g194(.A(i_0_), .B(i_5_), .Y(new_new_n217_));
  OAI220     g195(.A0(new_new_n87_), .A1(new_new_n189_), .B0(new_new_n182_), .B1(new_new_n138_), .Y(new_new_n218_));
  NAi31      g196(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n219_));
  NO2        g197(.A(new_new_n36_), .B(i_13_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n222_));
  INV        g200(.A(i_13_), .Y(new_new_n223_));
  NO2        g201(.A(i_12_), .B(new_new_n223_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n218_), .B(new_new_n216_), .Y(new_new_n225_));
  NO2        g203(.A(i_12_), .B(new_new_n37_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n184_), .B(i_4_), .Y(new_new_n227_));
  NA2        g205(.A(new_new_n227_), .B(new_new_n226_), .Y(new_new_n228_));
  OR2        g206(.A(i_8_), .B(i_7_), .Y(new_new_n229_));
  NO2        g207(.A(new_new_n229_), .B(new_new_n87_), .Y(new_new_n230_));
  NO2        g208(.A(new_new_n54_), .B(i_1_), .Y(new_new_n231_));
  NA2        g209(.A(new_new_n231_), .B(new_new_n230_), .Y(new_new_n232_));
  INV        g210(.A(i_12_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n45_), .B(new_new_n233_), .Y(new_new_n234_));
  NO3        g212(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n235_));
  NA2        g213(.A(i_2_), .B(i_1_), .Y(new_new_n236_));
  NO2        g214(.A(new_new_n232_), .B(new_new_n228_), .Y(new_new_n237_));
  NO3        g215(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n238_));
  NAi21      g216(.An(i_4_), .B(i_3_), .Y(new_new_n239_));
  NO2        g217(.A(i_0_), .B(i_6_), .Y(new_new_n240_));
  NOi41      g218(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n241_), .B(new_new_n240_), .Y(new_new_n242_));
  NO2        g220(.A(new_new_n236_), .B(new_new_n184_), .Y(new_new_n243_));
  NAi21      g221(.An(new_new_n242_), .B(new_new_n243_), .Y(new_new_n244_));
  INV        g222(.A(new_new_n244_), .Y(new_new_n245_));
  AOI220     g223(.A0(new_new_n245_), .A1(new_new_n40_), .B0(new_new_n237_), .B1(new_new_n204_), .Y(new_new_n246_));
  NO2        g224(.A(i_11_), .B(new_new_n223_), .Y(new_new_n247_));
  NOi21      g225(.An(i_1_), .B(i_6_), .Y(new_new_n248_));
  NAi21      g226(.An(i_3_), .B(i_7_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n233_), .B(i_9_), .Y(new_new_n250_));
  OR4        g228(.A(new_new_n250_), .B(new_new_n249_), .C(new_new_n248_), .D(new_new_n185_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n252_));
  NO2        g230(.A(i_12_), .B(i_3_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n74_), .B(i_5_), .Y(new_new_n254_));
  NA2        g232(.A(i_3_), .B(i_9_), .Y(new_new_n255_));
  NAi21      g233(.An(i_7_), .B(i_10_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n256_), .B(new_new_n255_), .Y(new_new_n257_));
  NA3        g235(.A(new_new_n257_), .B(new_new_n254_), .C(new_new_n65_), .Y(new_new_n258_));
  NA2        g236(.A(new_new_n258_), .B(new_new_n251_), .Y(new_new_n259_));
  NA3        g237(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n260_));
  INV        g238(.A(new_new_n148_), .Y(new_new_n261_));
  NA2        g239(.A(new_new_n233_), .B(i_13_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n262_), .B(new_new_n76_), .Y(new_new_n263_));
  AOI220     g241(.A0(new_new_n263_), .A1(new_new_n261_), .B0(new_new_n259_), .B1(new_new_n247_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n229_), .B(new_new_n37_), .Y(new_new_n265_));
  NA2        g243(.A(i_12_), .B(i_6_), .Y(new_new_n266_));
  OR2        g244(.A(i_13_), .B(i_9_), .Y(new_new_n267_));
  NO3        g245(.A(new_new_n267_), .B(new_new_n266_), .C(new_new_n49_), .Y(new_new_n268_));
  NO2        g246(.A(new_new_n239_), .B(i_2_), .Y(new_new_n269_));
  NA3        g247(.A(new_new_n269_), .B(new_new_n268_), .C(new_new_n45_), .Y(new_new_n270_));
  NA2        g248(.A(new_new_n247_), .B(i_9_), .Y(new_new_n271_));
  NA2        g249(.A(new_new_n254_), .B(new_new_n65_), .Y(new_new_n272_));
  OAI210     g250(.A0(new_new_n272_), .A1(new_new_n271_), .B0(new_new_n270_), .Y(new_new_n273_));
  NO3        g251(.A(i_11_), .B(new_new_n223_), .C(new_new_n25_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n249_), .B(i_8_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n273_), .B(new_new_n265_), .Y(new_new_n276_));
  NA4        g254(.A(new_new_n276_), .B(new_new_n264_), .C(new_new_n246_), .D(new_new_n225_), .Y(new_new_n277_));
  NO3        g255(.A(i_12_), .B(new_new_n223_), .C(new_new_n37_), .Y(new_new_n278_));
  INV        g256(.A(new_new_n278_), .Y(new_new_n279_));
  NO3        g257(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n236_), .B(i_0_), .Y(new_new_n281_));
  NA2        g259(.A(i_0_), .B(i_1_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n282_), .B(i_2_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n60_), .B(i_6_), .Y(new_new_n284_));
  NA3        g262(.A(new_new_n284_), .B(new_new_n283_), .C(new_new_n167_), .Y(new_new_n285_));
  NO2        g263(.A(i_3_), .B(i_10_), .Y(new_new_n286_));
  NA3        g264(.A(new_new_n286_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n287_));
  NO2        g265(.A(i_2_), .B(new_new_n105_), .Y(new_new_n288_));
  NA2        g266(.A(i_1_), .B(new_new_n36_), .Y(new_new_n289_));
  NO2        g267(.A(new_new_n289_), .B(i_8_), .Y(new_new_n290_));
  NA2        g268(.A(new_new_n290_), .B(new_new_n288_), .Y(new_new_n291_));
  AN2        g269(.A(i_3_), .B(i_10_), .Y(new_new_n292_));
  NA4        g270(.A(new_new_n292_), .B(new_new_n196_), .C(new_new_n178_), .D(new_new_n176_), .Y(new_new_n293_));
  NO2        g271(.A(i_5_), .B(new_new_n37_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n295_));
  OR2        g273(.A(new_new_n291_), .B(new_new_n287_), .Y(new_new_n296_));
  OAI220     g274(.A0(new_new_n296_), .A1(i_6_), .B0(new_new_n285_), .B1(new_new_n279_), .Y(new_new_n297_));
  NO4        g275(.A(new_new_n297_), .B(new_new_n277_), .C(new_new_n213_), .D(new_new_n169_), .Y(new_new_n298_));
  NO3        g276(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n300_));
  NO3        g278(.A(i_6_), .B(new_new_n193_), .C(i_7_), .Y(new_new_n301_));
  NO2        g279(.A(i_2_), .B(i_3_), .Y(new_new_n302_));
  OR2        g280(.A(i_0_), .B(i_5_), .Y(new_new_n303_));
  NA2        g281(.A(new_new_n217_), .B(new_new_n303_), .Y(new_new_n304_));
  NA4        g282(.A(new_new_n304_), .B(new_new_n230_), .C(new_new_n302_), .D(i_1_), .Y(new_new_n305_));
  NAi21      g283(.An(i_8_), .B(i_7_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n306_), .B(i_6_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n163_), .B(new_new_n47_), .Y(new_new_n308_));
  NA3        g286(.A(new_new_n308_), .B(new_new_n307_), .C(new_new_n167_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n309_), .B(new_new_n305_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n310_), .B(i_4_), .Y(new_new_n311_));
  NO2        g289(.A(i_12_), .B(i_10_), .Y(new_new_n312_));
  NOi21      g290(.An(i_5_), .B(i_0_), .Y(new_new_n313_));
  NA4        g291(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n314_));
  NO2        g292(.A(i_6_), .B(i_8_), .Y(new_new_n315_));
  NOi21      g293(.An(i_0_), .B(i_2_), .Y(new_new_n316_));
  BUFFER     g294(.A(new_new_n316_), .Y(new_new_n317_));
  NO2        g295(.A(i_1_), .B(i_7_), .Y(new_new_n318_));
  AO220      g296(.A0(new_new_n318_), .A1(new_new_n317_), .B0(new_new_n307_), .B1(new_new_n231_), .Y(new_new_n319_));
  NA3        g297(.A(new_new_n319_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n320_), .B(new_new_n311_), .Y(new_new_n321_));
  NO3        g299(.A(new_new_n229_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n322_));
  NO3        g300(.A(new_new_n306_), .B(i_2_), .C(i_1_), .Y(new_new_n323_));
  OAI210     g301(.A0(new_new_n323_), .A1(new_new_n322_), .B0(i_6_), .Y(new_new_n324_));
  NA3        g302(.A(new_new_n248_), .B(new_new_n288_), .C(new_new_n193_), .Y(new_new_n325_));
  AOI210     g303(.A0(new_new_n325_), .A1(new_new_n324_), .B0(new_new_n304_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n326_), .B(i_3_), .Y(new_new_n327_));
  INV        g305(.A(new_new_n85_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n282_), .B(new_new_n82_), .Y(new_new_n329_));
  NA2        g307(.A(new_new_n329_), .B(new_new_n137_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n96_), .B(new_new_n193_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n331_), .B(new_new_n64_), .Y(new_new_n332_));
  AOI210     g310(.A0(new_new_n332_), .A1(new_new_n330_), .B0(new_new_n328_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n193_), .B(i_9_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(new_new_n203_), .Y(new_new_n335_));
  INV        g313(.A(new_new_n333_), .Y(new_new_n336_));
  AOI210     g314(.A0(new_new_n336_), .A1(new_new_n327_), .B0(new_new_n166_), .Y(new_new_n337_));
  AOI210     g315(.A0(new_new_n321_), .A1(new_new_n299_), .B0(new_new_n337_), .Y(new_new_n338_));
  NOi32      g316(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n339_));
  INV        g317(.A(new_new_n339_), .Y(new_new_n340_));
  NAi21      g318(.An(i_0_), .B(i_6_), .Y(new_new_n341_));
  NAi21      g319(.An(i_1_), .B(i_5_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n342_), .B(new_new_n341_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n343_), .B(new_new_n25_), .Y(new_new_n344_));
  OAI210     g322(.A0(new_new_n344_), .A1(new_new_n164_), .B0(new_new_n242_), .Y(new_new_n345_));
  NAi41      g323(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n346_));
  OAI220     g324(.A0(new_new_n346_), .A1(new_new_n342_), .B0(new_new_n219_), .B1(new_new_n164_), .Y(new_new_n347_));
  AOI210     g325(.A0(new_new_n346_), .A1(new_new_n164_), .B0(new_new_n163_), .Y(new_new_n348_));
  OR2        g326(.A(new_new_n348_), .B(new_new_n347_), .Y(new_new_n349_));
  NO2        g327(.A(i_1_), .B(new_new_n105_), .Y(new_new_n350_));
  NAi21      g328(.An(i_3_), .B(i_4_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n351_), .B(i_9_), .Y(new_new_n352_));
  AN2        g330(.A(i_6_), .B(i_7_), .Y(new_new_n353_));
  OAI210     g331(.A0(new_new_n353_), .A1(new_new_n350_), .B0(new_new_n352_), .Y(new_new_n354_));
  NA2        g332(.A(i_2_), .B(i_7_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n351_), .B(i_10_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n354_), .B(new_new_n185_), .Y(new_new_n357_));
  AOI210     g335(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n358_));
  OAI210     g336(.A0(new_new_n358_), .A1(new_new_n188_), .B0(new_new_n356_), .Y(new_new_n359_));
  AOI220     g337(.A0(new_new_n356_), .A1(new_new_n318_), .B0(new_new_n235_), .B1(new_new_n188_), .Y(new_new_n360_));
  AOI210     g338(.A0(new_new_n360_), .A1(new_new_n359_), .B0(i_5_), .Y(new_new_n361_));
  NO4        g339(.A(new_new_n361_), .B(new_new_n357_), .C(new_new_n349_), .D(new_new_n345_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n362_), .B(new_new_n340_), .Y(new_new_n363_));
  AN2        g341(.A(i_12_), .B(i_5_), .Y(new_new_n364_));
  NO2        g342(.A(i_4_), .B(new_new_n26_), .Y(new_new_n365_));
  NA2        g343(.A(new_new_n365_), .B(new_new_n364_), .Y(new_new_n366_));
  NO2        g344(.A(i_11_), .B(i_6_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n239_), .B(i_5_), .Y(new_new_n368_));
  NO2        g346(.A(i_5_), .B(i_10_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n370_));
  NO3        g348(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n371_));
  NO2        g349(.A(i_3_), .B(new_new_n105_), .Y(new_new_n372_));
  NO2        g350(.A(i_11_), .B(i_12_), .Y(new_new_n373_));
  NA3        g351(.A(new_new_n117_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n374_), .B(new_new_n219_), .Y(new_new_n375_));
  NAi21      g353(.An(i_13_), .B(i_0_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n376_), .B(new_new_n236_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n375_), .B(new_new_n377_), .Y(new_new_n378_));
  INV        g356(.A(new_new_n378_), .Y(new_new_n379_));
  NA2        g357(.A(new_new_n45_), .B(new_new_n223_), .Y(new_new_n380_));
  NO3        g358(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n381_));
  NO2        g359(.A(i_0_), .B(i_11_), .Y(new_new_n382_));
  INV        g360(.A(i_5_), .Y(new_new_n383_));
  AN2        g361(.A(i_1_), .B(i_6_), .Y(new_new_n384_));
  NOi21      g362(.An(i_2_), .B(i_12_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n385_), .B(new_new_n384_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n386_), .B(new_new_n383_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n147_), .B(i_9_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n388_), .B(i_4_), .Y(new_new_n389_));
  NA2        g367(.A(new_new_n387_), .B(new_new_n389_), .Y(new_new_n390_));
  NAi21      g368(.An(i_9_), .B(i_4_), .Y(new_new_n391_));
  OR2        g369(.A(i_13_), .B(i_10_), .Y(new_new_n392_));
  NO3        g370(.A(new_new_n392_), .B(new_new_n122_), .C(new_new_n391_), .Y(new_new_n393_));
  OR2        g371(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n105_), .B(new_new_n25_), .Y(new_new_n395_));
  NA2        g373(.A(i_5_), .B(new_new_n209_), .Y(new_new_n396_));
  NO2        g374(.A(new_new_n396_), .B(new_new_n394_), .Y(new_new_n397_));
  INV        g375(.A(new_new_n397_), .Y(new_new_n398_));
  AOI210     g376(.A0(new_new_n398_), .A1(new_new_n390_), .B0(new_new_n26_), .Y(new_new_n399_));
  INV        g377(.A(new_new_n305_), .Y(new_new_n400_));
  AOI220     g378(.A0(new_new_n284_), .A1(new_new_n280_), .B0(new_new_n281_), .B1(new_new_n300_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n401_), .B(new_new_n171_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n402_), .B(new_new_n400_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n193_), .B(i_10_), .Y(new_new_n404_));
  NA3        g382(.A(new_new_n254_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n405_), .B(new_new_n404_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n301_), .B(new_new_n304_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n407_), .B(new_new_n189_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n408_), .B(new_new_n406_), .Y(new_new_n409_));
  AOI210     g387(.A0(new_new_n409_), .A1(new_new_n403_), .B0(new_new_n271_), .Y(new_new_n410_));
  NO4        g388(.A(new_new_n410_), .B(new_new_n399_), .C(new_new_n379_), .D(new_new_n363_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n74_), .B(i_13_), .Y(new_new_n412_));
  NO2        g390(.A(i_10_), .B(i_9_), .Y(new_new_n413_));
  NAi21      g391(.An(i_12_), .B(i_8_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n414_), .B(i_3_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n295_), .B(i_0_), .Y(new_new_n416_));
  NO3        g394(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n417_));
  NA2        g395(.A(new_new_n266_), .B(new_new_n101_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n418_), .B(new_new_n417_), .Y(new_new_n419_));
  NA2        g397(.A(i_8_), .B(i_9_), .Y(new_new_n420_));
  AOI210     g398(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n421_));
  OR2        g399(.A(new_new_n421_), .B(new_new_n420_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n278_), .B(new_new_n203_), .Y(new_new_n423_));
  OAI220     g401(.A0(new_new_n423_), .A1(new_new_n422_), .B0(new_new_n419_), .B1(new_new_n416_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n247_), .B(new_new_n294_), .Y(new_new_n425_));
  NO3        g403(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n426_));
  INV        g404(.A(new_new_n426_), .Y(new_new_n427_));
  NA3        g405(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n428_));
  NA4        g406(.A(new_new_n150_), .B(new_new_n120_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n429_));
  OAI220     g407(.A0(new_new_n429_), .A1(new_new_n428_), .B0(new_new_n427_), .B1(new_new_n425_), .Y(new_new_n430_));
  NO2        g408(.A(new_new_n430_), .B(new_new_n424_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n283_), .B(new_new_n112_), .Y(new_new_n432_));
  OR2        g410(.A(new_new_n432_), .B(new_new_n205_), .Y(new_new_n433_));
  OA210      g411(.A0(new_new_n335_), .A1(new_new_n105_), .B0(new_new_n285_), .Y(new_new_n434_));
  OA220      g412(.A0(new_new_n434_), .A1(new_new_n166_), .B0(new_new_n433_), .B1(new_new_n228_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n100_), .B(i_13_), .Y(new_new_n436_));
  NO2        g414(.A(i_2_), .B(i_13_), .Y(new_new_n437_));
  NO3        g415(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n438_));
  NO2        g416(.A(i_6_), .B(i_7_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n439_), .B(new_new_n438_), .Y(new_new_n440_));
  NO2        g418(.A(i_11_), .B(i_1_), .Y(new_new_n441_));
  OR2        g419(.A(i_11_), .B(i_8_), .Y(new_new_n442_));
  NOi21      g420(.An(i_2_), .B(i_7_), .Y(new_new_n443_));
  NAi31      g421(.An(new_new_n442_), .B(new_new_n443_), .C(i_0_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n392_), .B(i_6_), .Y(new_new_n445_));
  NA3        g423(.A(new_new_n445_), .B(i_1_), .C(new_new_n76_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n446_), .B(new_new_n444_), .Y(new_new_n447_));
  NO2        g425(.A(i_3_), .B(new_new_n193_), .Y(new_new_n448_));
  NO2        g426(.A(i_6_), .B(i_10_), .Y(new_new_n449_));
  NA4        g427(.A(new_new_n449_), .B(new_new_n299_), .C(new_new_n448_), .D(new_new_n233_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n450_), .B(new_new_n161_), .Y(new_new_n451_));
  NA3        g429(.A(new_new_n241_), .B(new_new_n173_), .C(new_new_n137_), .Y(new_new_n452_));
  NA2        g430(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n453_));
  NO2        g431(.A(new_new_n163_), .B(i_3_), .Y(new_new_n454_));
  NAi31      g432(.An(new_new_n453_), .B(new_new_n454_), .C(new_new_n224_), .Y(new_new_n455_));
  NA3        g433(.A(new_new_n370_), .B(new_new_n181_), .C(new_new_n154_), .Y(new_new_n456_));
  NA3        g434(.A(new_new_n456_), .B(new_new_n455_), .C(new_new_n452_), .Y(new_new_n457_));
  NO3        g435(.A(new_new_n457_), .B(new_new_n451_), .C(new_new_n447_), .Y(new_new_n458_));
  NA2        g436(.A(new_new_n417_), .B(new_new_n364_), .Y(new_new_n459_));
  NAi21      g437(.An(new_new_n215_), .B(new_new_n373_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n318_), .B(new_new_n217_), .Y(new_new_n461_));
  NO2        g439(.A(new_new_n26_), .B(i_5_), .Y(new_new_n462_));
  NO2        g440(.A(i_0_), .B(new_new_n87_), .Y(new_new_n463_));
  NA3        g441(.A(new_new_n463_), .B(new_new_n462_), .C(new_new_n147_), .Y(new_new_n464_));
  OR3        g442(.A(new_new_n289_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n465_));
  OAI220     g443(.A0(new_new_n465_), .A1(new_new_n464_), .B0(new_new_n461_), .B1(new_new_n460_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n27_), .B(i_10_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n299_), .B(new_new_n235_), .Y(new_new_n468_));
  OAI220     g446(.A0(new_new_n468_), .A1(new_new_n405_), .B0(new_new_n467_), .B1(new_new_n436_), .Y(new_new_n469_));
  NA4        g447(.A(new_new_n292_), .B(new_new_n222_), .C(new_new_n74_), .D(new_new_n233_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n470_), .B(new_new_n440_), .Y(new_new_n471_));
  NO3        g449(.A(new_new_n471_), .B(new_new_n469_), .C(new_new_n466_), .Y(new_new_n472_));
  NA4        g450(.A(new_new_n472_), .B(new_new_n458_), .C(new_new_n435_), .D(new_new_n431_), .Y(new_new_n473_));
  NA3        g451(.A(new_new_n292_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n474_));
  OAI210     g452(.A0(new_new_n287_), .A1(new_new_n183_), .B0(new_new_n474_), .Y(new_new_n475_));
  AN2        g453(.A(new_new_n280_), .B(new_new_n230_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n476_), .B(new_new_n475_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n127_), .B(new_new_n116_), .Y(new_new_n478_));
  AN2        g456(.A(new_new_n478_), .B(new_new_n417_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n299_), .B(i_0_), .Y(new_new_n480_));
  OAI210     g458(.A0(new_new_n480_), .A1(new_new_n228_), .B0(new_new_n293_), .Y(new_new_n481_));
  AOI220     g459(.A0(new_new_n481_), .A1(new_new_n307_), .B0(new_new_n479_), .B1(new_new_n295_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n339_), .B(new_new_n74_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n36_), .B(i_8_), .Y(new_new_n484_));
  NAi41      g462(.An(new_new_n483_), .B(new_new_n449_), .C(new_new_n484_), .D(new_new_n47_), .Y(new_new_n485_));
  AOI210     g463(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n393_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n486_), .B(new_new_n485_), .Y(new_new_n487_));
  INV        g465(.A(new_new_n487_), .Y(new_new_n488_));
  NO2        g466(.A(i_7_), .B(new_new_n197_), .Y(new_new_n489_));
  OR2        g467(.A(new_new_n184_), .B(i_4_), .Y(new_new_n490_));
  NO2        g468(.A(new_new_n490_), .B(new_new_n87_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n491_), .B(new_new_n489_), .Y(new_new_n492_));
  NA4        g470(.A(new_new_n492_), .B(new_new_n488_), .C(new_new_n482_), .D(new_new_n477_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n368_), .B(new_new_n283_), .Y(new_new_n494_));
  OAI210     g472(.A0(new_new_n366_), .A1(new_new_n170_), .B0(new_new_n494_), .Y(new_new_n495_));
  NO2        g473(.A(i_12_), .B(new_new_n193_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n496_), .B(new_new_n223_), .Y(new_new_n497_));
  NO3        g475(.A(new_new_n1007_), .B(new_new_n497_), .C(new_new_n432_), .Y(new_new_n498_));
  NOi31      g476(.An(new_new_n301_), .B(new_new_n392_), .C(new_new_n38_), .Y(new_new_n499_));
  OAI210     g477(.A0(new_new_n499_), .A1(new_new_n498_), .B0(new_new_n495_), .Y(new_new_n500_));
  AOI220     g478(.A0(new_new_n308_), .A1(new_new_n40_), .B0(new_new_n231_), .B1(new_new_n204_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n501_), .B(new_new_n490_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n45_), .B(i_10_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(i_6_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n504_), .B(new_new_n502_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n243_), .B(new_new_n240_), .Y(new_new_n506_));
  OAI220     g484(.A0(new_new_n506_), .A1(new_new_n262_), .B0(new_new_n436_), .B1(new_new_n138_), .Y(new_new_n507_));
  NA2        g485(.A(new_new_n507_), .B(new_new_n265_), .Y(new_new_n508_));
  NOi31      g486(.An(new_new_n281_), .B(new_new_n287_), .C(new_new_n183_), .Y(new_new_n509_));
  NA3        g487(.A(new_new_n292_), .B(new_new_n176_), .C(new_new_n100_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n220_), .B(new_new_n45_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n163_), .B(i_5_), .Y(new_new_n512_));
  NA3        g490(.A(new_new_n512_), .B(new_new_n380_), .C(new_new_n302_), .Y(new_new_n513_));
  OAI210     g491(.A0(new_new_n513_), .A1(new_new_n511_), .B0(new_new_n510_), .Y(new_new_n514_));
  OAI210     g492(.A0(new_new_n514_), .A1(new_new_n509_), .B0(new_new_n426_), .Y(new_new_n515_));
  NA4        g493(.A(new_new_n515_), .B(new_new_n508_), .C(new_new_n505_), .D(new_new_n500_), .Y(new_new_n516_));
  NA3        g494(.A(new_new_n217_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n517_));
  NA2        g495(.A(new_new_n278_), .B(new_new_n85_), .Y(new_new_n518_));
  AOI210     g496(.A0(new_new_n517_), .A1(new_new_n330_), .B0(new_new_n518_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n284_), .B(new_new_n280_), .Y(new_new_n520_));
  NO2        g498(.A(new_new_n520_), .B(new_new_n175_), .Y(new_new_n521_));
  NA2        g499(.A(new_new_n222_), .B(new_new_n221_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n413_), .B(new_new_n220_), .Y(new_new_n523_));
  NO2        g501(.A(new_new_n522_), .B(new_new_n523_), .Y(new_new_n524_));
  AOI210     g502(.A0(i_6_), .A1(new_new_n47_), .B0(new_new_n350_), .Y(new_new_n525_));
  NA2        g503(.A(i_0_), .B(new_new_n49_), .Y(new_new_n526_));
  NA3        g504(.A(new_new_n496_), .B(new_new_n274_), .C(new_new_n526_), .Y(new_new_n527_));
  NO2        g505(.A(new_new_n525_), .B(new_new_n527_), .Y(new_new_n528_));
  NO4        g506(.A(new_new_n528_), .B(new_new_n524_), .C(new_new_n521_), .D(new_new_n519_), .Y(new_new_n529_));
  NO4        g507(.A(new_new_n248_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n530_));
  NO3        g508(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n229_), .B(new_new_n36_), .Y(new_new_n532_));
  AN2        g510(.A(new_new_n532_), .B(new_new_n531_), .Y(new_new_n533_));
  OA210      g511(.A0(new_new_n533_), .A1(new_new_n530_), .B0(new_new_n339_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n392_), .B(i_1_), .Y(new_new_n535_));
  NOi31      g513(.An(new_new_n535_), .B(new_new_n418_), .C(new_new_n74_), .Y(new_new_n536_));
  AN4        g514(.A(new_new_n536_), .B(new_new_n389_), .C(new_new_n462_), .D(i_2_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n401_), .B(new_new_n179_), .Y(new_new_n538_));
  NO3        g516(.A(new_new_n538_), .B(new_new_n537_), .C(new_new_n534_), .Y(new_new_n539_));
  NOi21      g517(.An(i_10_), .B(i_6_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n541_));
  AOI220     g519(.A0(new_new_n278_), .A1(new_new_n541_), .B0(new_new_n274_), .B1(new_new_n540_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n542_), .B(new_new_n416_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n196_), .B(new_new_n37_), .Y(new_new_n545_));
  NOi31      g523(.An(new_new_n151_), .B(new_new_n545_), .C(new_new_n314_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n546_), .B(new_new_n543_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n483_), .B(new_new_n360_), .Y(new_new_n548_));
  INV        g526(.A(new_new_n302_), .Y(new_new_n549_));
  NO2        g527(.A(i_12_), .B(new_new_n87_), .Y(new_new_n550_));
  NA2        g528(.A(new_new_n176_), .B(i_0_), .Y(new_new_n551_));
  NO3        g529(.A(new_new_n551_), .B(new_new_n324_), .C(new_new_n287_), .Y(new_new_n552_));
  OR2        g530(.A(i_2_), .B(i_5_), .Y(new_new_n553_));
  OR2        g531(.A(new_new_n553_), .B(new_new_n384_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n554_), .B(new_new_n460_), .Y(new_new_n555_));
  NO3        g533(.A(new_new_n555_), .B(new_new_n552_), .C(new_new_n548_), .Y(new_new_n556_));
  NA4        g534(.A(new_new_n556_), .B(new_new_n547_), .C(new_new_n539_), .D(new_new_n529_), .Y(new_new_n557_));
  NO4        g535(.A(new_new_n557_), .B(new_new_n516_), .C(new_new_n493_), .D(new_new_n473_), .Y(new_new_n558_));
  NA4        g536(.A(new_new_n558_), .B(new_new_n411_), .C(new_new_n338_), .D(new_new_n298_), .Y(mai7));
  NO2        g537(.A(new_new_n96_), .B(new_new_n55_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n112_), .B(new_new_n93_), .Y(new_new_n561_));
  NA2        g539(.A(new_new_n365_), .B(new_new_n561_), .Y(new_new_n562_));
  NA2        g540(.A(new_new_n449_), .B(new_new_n85_), .Y(new_new_n563_));
  NA2        g541(.A(i_11_), .B(new_new_n193_), .Y(new_new_n564_));
  INV        g542(.A(new_new_n562_), .Y(new_new_n565_));
  NA3        g543(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n566_));
  NO2        g544(.A(new_new_n233_), .B(i_4_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n567_), .B(i_8_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n109_), .B(new_new_n566_), .Y(new_new_n569_));
  NA2        g547(.A(i_2_), .B(new_new_n87_), .Y(new_new_n570_));
  OAI210     g548(.A0(new_new_n90_), .A1(new_new_n201_), .B0(new_new_n202_), .Y(new_new_n571_));
  NO2        g549(.A(i_7_), .B(new_new_n37_), .Y(new_new_n572_));
  NA2        g550(.A(i_4_), .B(i_8_), .Y(new_new_n573_));
  AOI210     g551(.A0(new_new_n573_), .A1(new_new_n292_), .B0(new_new_n572_), .Y(new_new_n574_));
  OAI220     g552(.A0(new_new_n574_), .A1(new_new_n570_), .B0(new_new_n571_), .B1(i_13_), .Y(new_new_n575_));
  NO4        g553(.A(new_new_n575_), .B(new_new_n569_), .C(new_new_n565_), .D(new_new_n560_), .Y(new_new_n576_));
  AOI210     g554(.A0(new_new_n133_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n577_));
  AOI210     g555(.A0(new_new_n577_), .A1(new_new_n233_), .B0(new_new_n165_), .Y(new_new_n578_));
  OR2        g556(.A(i_6_), .B(i_10_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n579_), .B(new_new_n23_), .Y(new_new_n580_));
  OR3        g558(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n581_));
  NO3        g559(.A(new_new_n581_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n582_));
  INV        g560(.A(new_new_n198_), .Y(new_new_n583_));
  NO2        g561(.A(new_new_n582_), .B(new_new_n580_), .Y(new_new_n584_));
  OA220      g562(.A0(new_new_n584_), .A1(new_new_n549_), .B0(new_new_n578_), .B1(new_new_n267_), .Y(new_new_n585_));
  AOI210     g563(.A0(new_new_n585_), .A1(new_new_n576_), .B0(new_new_n64_), .Y(new_new_n586_));
  NOi21      g564(.An(i_11_), .B(i_7_), .Y(new_new_n587_));
  AO210      g565(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n588_));
  NO2        g566(.A(new_new_n588_), .B(new_new_n587_), .Y(new_new_n589_));
  NA2        g567(.A(new_new_n589_), .B(new_new_n204_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n590_), .B(new_new_n64_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n592_));
  AO210      g570(.A0(new_new_n592_), .A1(new_new_n360_), .B0(new_new_n41_), .Y(new_new_n593_));
  NO3        g571(.A(new_new_n256_), .B(new_new_n206_), .C(new_new_n564_), .Y(new_new_n594_));
  OAI210     g572(.A0(new_new_n594_), .A1(new_new_n224_), .B0(new_new_n64_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n385_), .B(new_new_n31_), .Y(new_new_n596_));
  OR2        g574(.A(new_new_n206_), .B(new_new_n112_), .Y(new_new_n597_));
  NA2        g575(.A(new_new_n597_), .B(new_new_n596_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n64_), .B(i_9_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n599_), .B(i_4_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n600_), .B(new_new_n598_), .Y(new_new_n601_));
  NO2        g579(.A(i_1_), .B(i_12_), .Y(new_new_n602_));
  NA3        g580(.A(new_new_n602_), .B(new_new_n114_), .C(new_new_n24_), .Y(new_new_n603_));
  BUFFER     g581(.A(new_new_n603_), .Y(new_new_n604_));
  NA4        g582(.A(new_new_n604_), .B(new_new_n601_), .C(new_new_n595_), .D(new_new_n593_), .Y(new_new_n605_));
  OAI210     g583(.A0(new_new_n605_), .A1(new_new_n591_), .B0(i_6_), .Y(new_new_n606_));
  NO2        g584(.A(i_6_), .B(i_11_), .Y(new_new_n607_));
  INV        g585(.A(new_new_n419_), .Y(new_new_n608_));
  NO4        g586(.A(new_new_n214_), .B(new_new_n133_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n609_));
  NA2        g587(.A(new_new_n609_), .B(new_new_n599_), .Y(new_new_n610_));
  NA2        g588(.A(new_new_n233_), .B(i_6_), .Y(new_new_n611_));
  NO3        g589(.A(new_new_n579_), .B(new_new_n229_), .C(new_new_n23_), .Y(new_new_n612_));
  AOI210     g590(.A0(i_1_), .A1(new_new_n257_), .B0(new_new_n612_), .Y(new_new_n613_));
  OAI210     g591(.A0(new_new_n613_), .A1(new_new_n45_), .B0(new_new_n610_), .Y(new_new_n614_));
  INV        g592(.A(i_2_), .Y(new_new_n615_));
  NA2        g593(.A(new_new_n143_), .B(i_9_), .Y(new_new_n616_));
  NA3        g594(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n47_), .B(i_1_), .Y(new_new_n618_));
  NA3        g596(.A(new_new_n618_), .B(new_new_n266_), .C(new_new_n45_), .Y(new_new_n619_));
  OAI220     g597(.A0(new_new_n619_), .A1(new_new_n617_), .B0(new_new_n616_), .B1(new_new_n615_), .Y(new_new_n620_));
  NA3        g598(.A(new_new_n599_), .B(new_new_n302_), .C(i_6_), .Y(new_new_n621_));
  NO2        g599(.A(new_new_n621_), .B(new_new_n23_), .Y(new_new_n622_));
  AOI210     g600(.A0(new_new_n441_), .A1(new_new_n395_), .B0(new_new_n238_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n623_), .B(new_new_n570_), .Y(new_new_n624_));
  NO2        g602(.A(i_11_), .B(new_new_n37_), .Y(new_new_n625_));
  OR3        g603(.A(new_new_n624_), .B(new_new_n622_), .C(new_new_n620_), .Y(new_new_n626_));
  NO3        g604(.A(new_new_n626_), .B(new_new_n614_), .C(new_new_n608_), .Y(new_new_n627_));
  NO2        g605(.A(new_new_n233_), .B(new_new_n105_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n628_), .B(new_new_n587_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n629_), .B(i_1_), .Y(new_new_n630_));
  NO2        g608(.A(new_new_n630_), .B(new_new_n581_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n391_), .B(new_new_n87_), .Y(new_new_n632_));
  NA2        g610(.A(new_new_n631_), .B(new_new_n47_), .Y(new_new_n633_));
  NA2        g611(.A(i_3_), .B(new_new_n193_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n634_), .B(new_new_n119_), .Y(new_new_n635_));
  AN2        g613(.A(new_new_n635_), .B(new_new_n504_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n229_), .B(new_new_n45_), .Y(new_new_n637_));
  NO3        g615(.A(new_new_n637_), .B(new_new_n295_), .C(new_new_n234_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n122_), .B(new_new_n37_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n639_), .B(i_6_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n87_), .B(i_9_), .Y(new_new_n641_));
  NO2        g619(.A(new_new_n641_), .B(new_new_n64_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n642_), .B(new_new_n602_), .Y(new_new_n643_));
  NO4        g621(.A(new_new_n643_), .B(new_new_n640_), .C(new_new_n638_), .D(i_4_), .Y(new_new_n644_));
  NA2        g622(.A(i_1_), .B(i_3_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n420_), .B(new_new_n96_), .Y(new_new_n646_));
  AOI210     g624(.A0(new_new_n637_), .A1(new_new_n540_), .B0(new_new_n646_), .Y(new_new_n647_));
  NO2        g625(.A(new_new_n647_), .B(new_new_n645_), .Y(new_new_n648_));
  NO3        g626(.A(new_new_n648_), .B(new_new_n644_), .C(new_new_n636_), .Y(new_new_n649_));
  NA4        g627(.A(new_new_n649_), .B(new_new_n633_), .C(new_new_n627_), .D(new_new_n606_), .Y(new_new_n650_));
  NO3        g628(.A(new_new_n442_), .B(i_3_), .C(i_7_), .Y(new_new_n651_));
  NOi21      g629(.An(new_new_n651_), .B(i_10_), .Y(new_new_n652_));
  OA210      g630(.A0(new_new_n652_), .A1(new_new_n241_), .B0(new_new_n87_), .Y(new_new_n653_));
  NA2        g631(.A(new_new_n353_), .B(new_new_n352_), .Y(new_new_n654_));
  NA3        g632(.A(new_new_n449_), .B(new_new_n484_), .C(new_new_n47_), .Y(new_new_n655_));
  NA3        g633(.A(new_new_n165_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n656_));
  NA3        g634(.A(new_new_n656_), .B(new_new_n655_), .C(new_new_n654_), .Y(new_new_n657_));
  OAI210     g635(.A0(new_new_n657_), .A1(new_new_n653_), .B0(i_1_), .Y(new_new_n658_));
  AOI210     g636(.A0(new_new_n266_), .A1(new_new_n101_), .B0(i_1_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n351_), .B(i_2_), .Y(new_new_n660_));
  NA2        g638(.A(new_new_n660_), .B(new_new_n659_), .Y(new_new_n661_));
  OAI210     g639(.A0(new_new_n621_), .A1(new_new_n414_), .B0(new_new_n661_), .Y(new_new_n662_));
  INV        g640(.A(new_new_n662_), .Y(new_new_n663_));
  AOI210     g641(.A0(new_new_n663_), .A1(new_new_n658_), .B0(i_13_), .Y(new_new_n664_));
  NO2        g642(.A(new_new_n55_), .B(i_12_), .Y(new_new_n665_));
  INV        g643(.A(new_new_n665_), .Y(new_new_n666_));
  NO2        g644(.A(new_new_n443_), .B(new_new_n24_), .Y(new_new_n667_));
  AOI220     g645(.A0(new_new_n667_), .A1(new_new_n632_), .B0(new_new_n241_), .B1(new_new_n136_), .Y(new_new_n668_));
  OAI220     g646(.A0(new_new_n668_), .A1(new_new_n41_), .B0(new_new_n666_), .B1(new_new_n96_), .Y(new_new_n669_));
  INV        g647(.A(new_new_n669_), .Y(new_new_n670_));
  INV        g648(.A(new_new_n119_), .Y(new_new_n671_));
  AOI220     g649(.A0(new_new_n671_), .A1(new_new_n73_), .B0(new_new_n367_), .B1(new_new_n618_), .Y(new_new_n672_));
  NO2        g650(.A(new_new_n672_), .B(new_new_n239_), .Y(new_new_n673_));
  AOI210     g651(.A0(new_new_n414_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n674_));
  NOi31      g652(.An(new_new_n674_), .B(new_new_n563_), .C(new_new_n45_), .Y(new_new_n675_));
  NA2        g653(.A(new_new_n132_), .B(i_13_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n617_), .B(new_new_n119_), .Y(new_new_n677_));
  INV        g655(.A(new_new_n677_), .Y(new_new_n678_));
  OAI220     g656(.A0(new_new_n678_), .A1(new_new_n72_), .B0(new_new_n676_), .B1(new_new_n659_), .Y(new_new_n679_));
  NO3        g657(.A(new_new_n72_), .B(new_new_n32_), .C(new_new_n105_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n26_), .B(new_new_n193_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n681_), .B(i_7_), .Y(new_new_n682_));
  NO3        g660(.A(new_new_n443_), .B(new_new_n233_), .C(new_new_n87_), .Y(new_new_n683_));
  AOI210     g661(.A0(new_new_n683_), .A1(new_new_n682_), .B0(new_new_n680_), .Y(new_new_n684_));
  AOI220     g662(.A0(new_new_n367_), .A1(new_new_n618_), .B0(new_new_n95_), .B1(new_new_n106_), .Y(new_new_n685_));
  OAI220     g663(.A0(new_new_n685_), .A1(new_new_n568_), .B0(new_new_n684_), .B1(new_new_n583_), .Y(new_new_n686_));
  NO4        g664(.A(new_new_n686_), .B(new_new_n679_), .C(new_new_n675_), .D(new_new_n673_), .Y(new_new_n687_));
  OR2        g665(.A(i_11_), .B(i_6_), .Y(new_new_n688_));
  NA3        g666(.A(new_new_n567_), .B(new_new_n681_), .C(i_7_), .Y(new_new_n689_));
  AOI210     g667(.A0(new_new_n689_), .A1(new_new_n678_), .B0(new_new_n688_), .Y(new_new_n690_));
  NA3        g668(.A(new_new_n385_), .B(new_new_n572_), .C(new_new_n101_), .Y(new_new_n691_));
  NA2        g669(.A(new_new_n607_), .B(i_13_), .Y(new_new_n692_));
  NA2        g670(.A(new_new_n106_), .B(new_new_n681_), .Y(new_new_n693_));
  NAi21      g671(.An(i_11_), .B(i_12_), .Y(new_new_n694_));
  NOi41      g672(.An(new_new_n115_), .B(new_new_n694_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n695_));
  NA2        g673(.A(new_new_n695_), .B(new_new_n693_), .Y(new_new_n696_));
  NA3        g674(.A(new_new_n696_), .B(new_new_n692_), .C(new_new_n691_), .Y(new_new_n697_));
  OAI210     g675(.A0(new_new_n697_), .A1(new_new_n690_), .B0(new_new_n64_), .Y(new_new_n698_));
  NO2        g676(.A(i_2_), .B(i_12_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n350_), .B(new_new_n699_), .Y(new_new_n700_));
  NA2        g678(.A(i_8_), .B(new_new_n25_), .Y(new_new_n701_));
  NO3        g679(.A(new_new_n701_), .B(new_new_n365_), .C(new_new_n567_), .Y(new_new_n702_));
  OAI210     g680(.A0(new_new_n702_), .A1(new_new_n352_), .B0(new_new_n350_), .Y(new_new_n703_));
  NO2        g681(.A(new_new_n133_), .B(i_2_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n703_), .B(new_new_n700_), .Y(new_new_n705_));
  NA3        g683(.A(new_new_n705_), .B(new_new_n46_), .C(new_new_n223_), .Y(new_new_n706_));
  NA4        g684(.A(new_new_n706_), .B(new_new_n698_), .C(new_new_n687_), .D(new_new_n670_), .Y(new_new_n707_));
  OR4        g685(.A(new_new_n707_), .B(new_new_n664_), .C(new_new_n650_), .D(new_new_n586_), .Y(mai5));
  NA2        g686(.A(new_new_n629_), .B(new_new_n269_), .Y(new_new_n709_));
  AN2        g687(.A(new_new_n24_), .B(i_10_), .Y(new_new_n710_));
  NA3        g688(.A(new_new_n710_), .B(new_new_n699_), .C(new_new_n112_), .Y(new_new_n711_));
  NO2        g689(.A(new_new_n568_), .B(i_11_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n90_), .B(new_new_n712_), .Y(new_new_n713_));
  NA3        g691(.A(new_new_n713_), .B(new_new_n711_), .C(new_new_n709_), .Y(new_new_n714_));
  NO3        g692(.A(i_11_), .B(new_new_n233_), .C(i_13_), .Y(new_new_n715_));
  NO2        g693(.A(new_new_n129_), .B(new_new_n23_), .Y(new_new_n716_));
  NA2        g694(.A(i_12_), .B(i_8_), .Y(new_new_n717_));
  OAI210     g695(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n717_), .Y(new_new_n718_));
  INV        g696(.A(new_new_n413_), .Y(new_new_n719_));
  AOI220     g697(.A0(new_new_n302_), .A1(new_new_n544_), .B0(new_new_n718_), .B1(new_new_n716_), .Y(new_new_n720_));
  INV        g698(.A(new_new_n720_), .Y(new_new_n721_));
  NO2        g699(.A(new_new_n721_), .B(new_new_n714_), .Y(new_new_n722_));
  INV        g700(.A(new_new_n173_), .Y(new_new_n723_));
  INV        g701(.A(new_new_n241_), .Y(new_new_n724_));
  OAI210     g702(.A0(new_new_n660_), .A1(new_new_n415_), .B0(new_new_n115_), .Y(new_new_n725_));
  AOI210     g703(.A0(new_new_n725_), .A1(new_new_n724_), .B0(new_new_n723_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n420_), .B(new_new_n26_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n727_), .B(new_new_n395_), .Y(new_new_n728_));
  NA2        g706(.A(new_new_n728_), .B(i_2_), .Y(new_new_n729_));
  INV        g707(.A(new_new_n729_), .Y(new_new_n730_));
  AOI210     g708(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n392_), .Y(new_new_n731_));
  AOI210     g709(.A0(new_new_n731_), .A1(new_new_n730_), .B0(new_new_n726_), .Y(new_new_n732_));
  NO2        g710(.A(new_new_n190_), .B(new_new_n130_), .Y(new_new_n733_));
  OAI210     g711(.A0(new_new_n733_), .A1(new_new_n716_), .B0(i_2_), .Y(new_new_n734_));
  INV        g712(.A(new_new_n174_), .Y(new_new_n735_));
  NO3        g713(.A(new_new_n588_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n736_));
  AOI210     g714(.A0(new_new_n735_), .A1(new_new_n90_), .B0(new_new_n736_), .Y(new_new_n737_));
  AOI210     g715(.A0(new_new_n737_), .A1(new_new_n734_), .B0(new_new_n193_), .Y(new_new_n738_));
  OA210      g716(.A0(new_new_n589_), .A1(new_new_n131_), .B0(i_13_), .Y(new_new_n739_));
  NA2        g717(.A(new_new_n198_), .B(new_new_n201_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n157_), .B(new_new_n564_), .Y(new_new_n741_));
  AOI210     g719(.A0(new_new_n741_), .A1(new_new_n740_), .B0(new_new_n355_), .Y(new_new_n742_));
  AOI210     g720(.A0(new_new_n206_), .A1(new_new_n153_), .B0(new_new_n484_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n743_), .B(new_new_n395_), .Y(new_new_n744_));
  NO2        g722(.A(new_new_n106_), .B(new_new_n45_), .Y(new_new_n745_));
  INV        g723(.A(new_new_n288_), .Y(new_new_n746_));
  NA4        g724(.A(new_new_n746_), .B(new_new_n292_), .C(new_new_n129_), .D(new_new_n43_), .Y(new_new_n747_));
  OAI210     g725(.A0(new_new_n747_), .A1(new_new_n745_), .B0(new_new_n744_), .Y(new_new_n748_));
  NO4        g726(.A(new_new_n748_), .B(new_new_n742_), .C(new_new_n739_), .D(new_new_n738_), .Y(new_new_n749_));
  NA2        g727(.A(new_new_n544_), .B(new_new_n28_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n715_), .B(new_new_n275_), .Y(new_new_n751_));
  NA2        g729(.A(new_new_n751_), .B(new_new_n750_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n63_), .B(i_12_), .Y(new_new_n753_));
  NO2        g731(.A(new_new_n753_), .B(new_new_n131_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n754_), .B(new_new_n564_), .Y(new_new_n755_));
  AOI220     g733(.A0(new_new_n755_), .A1(new_new_n36_), .B0(new_new_n752_), .B1(new_new_n47_), .Y(new_new_n756_));
  NA4        g734(.A(new_new_n756_), .B(new_new_n749_), .C(new_new_n732_), .D(new_new_n722_), .Y(mai6));
  NO2        g735(.A(new_new_n185_), .B(new_new_n144_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n758_), .B(new_new_n704_), .Y(new_new_n759_));
  NA4        g737(.A(new_new_n369_), .B(new_new_n448_), .C(new_new_n72_), .D(new_new_n105_), .Y(new_new_n760_));
  INV        g738(.A(new_new_n760_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n219_), .B(new_new_n453_), .Y(new_new_n762_));
  NO2        g740(.A(i_11_), .B(i_9_), .Y(new_new_n763_));
  NO2        g741(.A(new_new_n761_), .B(new_new_n313_), .Y(new_new_n764_));
  AO210      g742(.A0(new_new_n764_), .A1(new_new_n759_), .B0(i_12_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n356_), .B(new_new_n318_), .Y(new_new_n766_));
  NA2        g744(.A(new_new_n550_), .B(new_new_n64_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n652_), .B(new_new_n72_), .Y(new_new_n768_));
  BUFFER     g746(.A(new_new_n592_), .Y(new_new_n769_));
  NA4        g747(.A(new_new_n769_), .B(new_new_n768_), .C(new_new_n767_), .D(new_new_n766_), .Y(new_new_n770_));
  INV        g748(.A(new_new_n195_), .Y(new_new_n771_));
  AOI220     g749(.A0(new_new_n771_), .A1(new_new_n763_), .B0(new_new_n770_), .B1(new_new_n74_), .Y(new_new_n772_));
  INV        g750(.A(new_new_n312_), .Y(new_new_n773_));
  NA2        g751(.A(new_new_n76_), .B(new_new_n136_), .Y(new_new_n774_));
  INV        g752(.A(new_new_n129_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n775_), .B(new_new_n47_), .Y(new_new_n776_));
  AOI210     g754(.A0(new_new_n776_), .A1(new_new_n774_), .B0(new_new_n773_), .Y(new_new_n777_));
  NO2        g755(.A(new_new_n248_), .B(i_9_), .Y(new_new_n778_));
  NA2        g756(.A(new_new_n778_), .B(new_new_n753_), .Y(new_new_n779_));
  NO2        g757(.A(new_new_n779_), .B(new_new_n185_), .Y(new_new_n780_));
  NO2        g758(.A(new_new_n32_), .B(i_11_), .Y(new_new_n781_));
  NA3        g759(.A(new_new_n781_), .B(new_new_n439_), .C(new_new_n369_), .Y(new_new_n782_));
  NAi32      g760(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n783_));
  NO2        g761(.A(new_new_n688_), .B(new_new_n783_), .Y(new_new_n784_));
  OAI210     g762(.A0(new_new_n651_), .A1(new_new_n532_), .B0(new_new_n531_), .Y(new_new_n785_));
  NAi31      g763(.An(new_new_n784_), .B(new_new_n785_), .C(new_new_n782_), .Y(new_new_n786_));
  OR3        g764(.A(new_new_n786_), .B(new_new_n780_), .C(new_new_n777_), .Y(new_new_n787_));
  AO220      g765(.A0(new_new_n343_), .A1(new_new_n334_), .B0(new_new_n371_), .B1(new_new_n564_), .Y(new_new_n788_));
  NA3        g766(.A(new_new_n788_), .B(new_new_n253_), .C(i_7_), .Y(new_new_n789_));
  BUFFER     g767(.A(new_new_n589_), .Y(new_new_n790_));
  NA3        g768(.A(new_new_n790_), .B(new_new_n152_), .C(new_new_n70_), .Y(new_new_n791_));
  OR2        g769(.A(new_new_n719_), .B(new_new_n36_), .Y(new_new_n792_));
  NA3        g770(.A(new_new_n792_), .B(new_new_n791_), .C(new_new_n789_), .Y(new_new_n793_));
  OAI210     g771(.A0(i_6_), .A1(i_11_), .B0(new_new_n88_), .Y(new_new_n794_));
  AOI220     g772(.A0(new_new_n794_), .A1(new_new_n531_), .B0(new_new_n762_), .B1(new_new_n682_), .Y(new_new_n795_));
  NA2        g773(.A(new_new_n371_), .B(new_new_n71_), .Y(new_new_n796_));
  NA3        g774(.A(new_new_n796_), .B(new_new_n795_), .C(new_new_n571_), .Y(new_new_n797_));
  AO210      g775(.A0(new_new_n484_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n798_));
  NA3        g776(.A(new_new_n798_), .B(new_new_n449_), .C(new_new_n217_), .Y(new_new_n799_));
  AOI210     g777(.A0(new_new_n415_), .A1(new_new_n413_), .B0(new_new_n530_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n579_), .B(new_new_n106_), .Y(new_new_n801_));
  OAI210     g779(.A0(new_new_n801_), .A1(new_new_n116_), .B0(new_new_n382_), .Y(new_new_n802_));
  INV        g780(.A(new_new_n554_), .Y(new_new_n803_));
  NA3        g781(.A(new_new_n803_), .B(new_new_n312_), .C(i_7_), .Y(new_new_n804_));
  NA4        g782(.A(new_new_n804_), .B(new_new_n802_), .C(new_new_n800_), .D(new_new_n799_), .Y(new_new_n805_));
  NO4        g783(.A(new_new_n805_), .B(new_new_n797_), .C(new_new_n793_), .D(new_new_n787_), .Y(new_new_n806_));
  NA4        g784(.A(new_new_n806_), .B(new_new_n772_), .C(new_new_n765_), .D(new_new_n362_), .Y(mai3));
  NA2        g785(.A(i_12_), .B(i_10_), .Y(new_new_n808_));
  NA2        g786(.A(i_6_), .B(i_7_), .Y(new_new_n809_));
  NO2        g787(.A(new_new_n809_), .B(i_0_), .Y(new_new_n810_));
  NO2        g788(.A(i_11_), .B(new_new_n233_), .Y(new_new_n811_));
  OAI210     g789(.A0(new_new_n810_), .A1(new_new_n281_), .B0(new_new_n811_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n812_), .B(new_new_n193_), .Y(new_new_n813_));
  NO3        g791(.A(new_new_n416_), .B(new_new_n93_), .C(new_new_n45_), .Y(new_new_n814_));
  OA210      g792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n176_), .Y(new_new_n815_));
  NOi21      g793(.An(new_new_n100_), .B(new_new_n728_), .Y(new_new_n816_));
  NO3        g794(.A(new_new_n597_), .B(new_new_n420_), .C(new_new_n136_), .Y(new_new_n817_));
  AN2        g795(.A(new_new_n418_), .B(new_new_n56_), .Y(new_new_n818_));
  NO3        g796(.A(new_new_n818_), .B(new_new_n817_), .C(new_new_n816_), .Y(new_new_n819_));
  NO2        g797(.A(new_new_n819_), .B(new_new_n49_), .Y(new_new_n820_));
  NO4        g798(.A(new_new_n358_), .B(new_new_n364_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n821_));
  NA2        g799(.A(new_new_n185_), .B(new_new_n540_), .Y(new_new_n822_));
  NOi21      g800(.An(new_new_n822_), .B(new_new_n821_), .Y(new_new_n823_));
  NO2        g801(.A(new_new_n823_), .B(new_new_n64_), .Y(new_new_n824_));
  NOi21      g802(.An(i_5_), .B(i_9_), .Y(new_new_n825_));
  NA2        g803(.A(new_new_n825_), .B(new_new_n412_), .Y(new_new_n826_));
  BUFFER     g804(.A(new_new_n266_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n827_), .B(new_new_n441_), .Y(new_new_n828_));
  NO3        g806(.A(new_new_n388_), .B(new_new_n266_), .C(new_new_n74_), .Y(new_new_n829_));
  NO2        g807(.A(new_new_n177_), .B(new_new_n153_), .Y(new_new_n830_));
  AOI210     g808(.A0(new_new_n830_), .A1(new_new_n240_), .B0(new_new_n829_), .Y(new_new_n831_));
  OAI220     g809(.A0(new_new_n831_), .A1(new_new_n183_), .B0(new_new_n828_), .B1(new_new_n826_), .Y(new_new_n832_));
  NO4        g810(.A(new_new_n832_), .B(new_new_n824_), .C(new_new_n820_), .D(new_new_n815_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n185_), .B(new_new_n24_), .Y(new_new_n834_));
  NO2        g812(.A(new_new_n639_), .B(new_new_n561_), .Y(new_new_n835_));
  NO2        g813(.A(new_new_n835_), .B(new_new_n834_), .Y(new_new_n836_));
  INV        g814(.A(new_new_n836_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n369_), .B(new_new_n282_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n838_), .B(new_new_n677_), .Y(new_new_n839_));
  NA2        g817(.A(new_new_n541_), .B(i_0_), .Y(new_new_n840_));
  NO3        g818(.A(new_new_n840_), .B(new_new_n366_), .C(new_new_n90_), .Y(new_new_n841_));
  NO4        g819(.A(new_new_n553_), .B(new_new_n214_), .C(new_new_n392_), .D(new_new_n384_), .Y(new_new_n842_));
  AOI210     g820(.A0(new_new_n842_), .A1(i_11_), .B0(new_new_n841_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n715_), .B(new_new_n313_), .Y(new_new_n844_));
  AOI210     g822(.A0(new_new_n449_), .A1(new_new_n90_), .B0(new_new_n59_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n845_), .B(new_new_n844_), .Y(new_new_n846_));
  NO2        g824(.A(new_new_n250_), .B(new_new_n159_), .Y(new_new_n847_));
  NA2        g825(.A(i_0_), .B(i_10_), .Y(new_new_n848_));
  INV        g826(.A(new_new_n503_), .Y(new_new_n849_));
  NO4        g827(.A(new_new_n119_), .B(new_new_n59_), .C(new_new_n634_), .D(i_5_), .Y(new_new_n850_));
  AO220      g828(.A0(new_new_n850_), .A1(new_new_n849_), .B0(new_new_n847_), .B1(i_6_), .Y(new_new_n851_));
  AOI220     g829(.A0(new_new_n316_), .A1(new_new_n102_), .B0(new_new_n185_), .B1(new_new_n85_), .Y(new_new_n852_));
  NA2        g830(.A(new_new_n535_), .B(i_4_), .Y(new_new_n853_));
  NA2        g831(.A(new_new_n188_), .B(new_new_n201_), .Y(new_new_n854_));
  OAI220     g832(.A0(new_new_n854_), .A1(new_new_n844_), .B0(new_new_n853_), .B1(new_new_n852_), .Y(new_new_n855_));
  NO3        g833(.A(new_new_n855_), .B(new_new_n851_), .C(new_new_n846_), .Y(new_new_n856_));
  NA4        g834(.A(new_new_n856_), .B(new_new_n843_), .C(new_new_n839_), .D(new_new_n837_), .Y(new_new_n857_));
  NO2        g835(.A(new_new_n107_), .B(new_new_n37_), .Y(new_new_n858_));
  NA2        g836(.A(i_11_), .B(i_9_), .Y(new_new_n859_));
  NO3        g837(.A(i_12_), .B(new_new_n859_), .C(new_new_n570_), .Y(new_new_n860_));
  AN2        g838(.A(new_new_n860_), .B(new_new_n858_), .Y(new_new_n861_));
  NO2        g839(.A(new_new_n49_), .B(i_7_), .Y(new_new_n862_));
  NA2        g840(.A(new_new_n370_), .B(new_new_n181_), .Y(new_new_n863_));
  INV        g841(.A(new_new_n863_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n859_), .B(new_new_n74_), .Y(new_new_n865_));
  NO2        g843(.A(new_new_n177_), .B(i_0_), .Y(new_new_n866_));
  INV        g844(.A(new_new_n866_), .Y(new_new_n867_));
  NA2        g845(.A(new_new_n439_), .B(new_new_n227_), .Y(new_new_n868_));
  AOI210     g846(.A0(new_new_n353_), .A1(new_new_n42_), .B0(new_new_n381_), .Y(new_new_n869_));
  OAI220     g847(.A0(new_new_n869_), .A1(new_new_n826_), .B0(new_new_n868_), .B1(new_new_n867_), .Y(new_new_n870_));
  NO3        g848(.A(new_new_n870_), .B(new_new_n864_), .C(new_new_n861_), .Y(new_new_n871_));
  NA2        g849(.A(new_new_n625_), .B(new_new_n126_), .Y(new_new_n872_));
  NO2        g850(.A(i_6_), .B(new_new_n872_), .Y(new_new_n873_));
  NA2        g851(.A(new_new_n173_), .B(new_new_n107_), .Y(new_new_n874_));
  INV        g852(.A(new_new_n873_), .Y(new_new_n875_));
  NOi21      g853(.An(i_7_), .B(i_5_), .Y(new_new_n876_));
  NOi31      g854(.An(new_new_n876_), .B(i_0_), .C(new_new_n694_), .Y(new_new_n877_));
  NA3        g855(.A(new_new_n877_), .B(new_new_n365_), .C(i_6_), .Y(new_new_n878_));
  BUFFER     g856(.A(new_new_n878_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n376_), .B(new_new_n346_), .C(new_new_n342_), .Y(new_new_n880_));
  NO2        g858(.A(new_new_n260_), .B(new_new_n303_), .Y(new_new_n881_));
  NO2        g859(.A(new_new_n694_), .B(new_new_n255_), .Y(new_new_n882_));
  AOI210     g860(.A0(new_new_n882_), .A1(new_new_n881_), .B0(new_new_n880_), .Y(new_new_n883_));
  NA4        g861(.A(new_new_n883_), .B(new_new_n879_), .C(new_new_n875_), .D(new_new_n871_), .Y(new_new_n884_));
  NO2        g862(.A(new_new_n834_), .B(new_new_n236_), .Y(new_new_n885_));
  AN2        g863(.A(new_new_n315_), .B(new_new_n313_), .Y(new_new_n886_));
  AN2        g864(.A(new_new_n886_), .B(new_new_n830_), .Y(new_new_n887_));
  OAI210     g865(.A0(new_new_n887_), .A1(new_new_n885_), .B0(i_10_), .Y(new_new_n888_));
  NO2        g866(.A(new_new_n808_), .B(new_new_n302_), .Y(new_new_n889_));
  OA210      g867(.A0(new_new_n439_), .A1(new_new_n222_), .B0(new_new_n438_), .Y(new_new_n890_));
  NA2        g868(.A(new_new_n889_), .B(new_new_n865_), .Y(new_new_n891_));
  NA2        g869(.A(new_new_n865_), .B(new_new_n292_), .Y(new_new_n892_));
  OAI210     g870(.A0(i_2_), .A1(new_new_n187_), .B0(new_new_n892_), .Y(new_new_n893_));
  NA2        g871(.A(new_new_n893_), .B(new_new_n439_), .Y(new_new_n894_));
  NA2        g872(.A(new_new_n96_), .B(new_new_n45_), .Y(new_new_n895_));
  NO2        g873(.A(new_new_n76_), .B(new_new_n717_), .Y(new_new_n896_));
  AOI220     g874(.A0(new_new_n896_), .A1(new_new_n895_), .B0(new_new_n176_), .B1(new_new_n561_), .Y(new_new_n897_));
  NO2        g875(.A(new_new_n897_), .B(new_new_n48_), .Y(new_new_n898_));
  NO3        g876(.A(new_new_n553_), .B(new_new_n341_), .C(new_new_n24_), .Y(new_new_n899_));
  AOI210     g877(.A0(new_new_n667_), .A1(new_new_n512_), .B0(new_new_n899_), .Y(new_new_n900_));
  NAi21      g878(.An(i_9_), .B(i_5_), .Y(new_new_n901_));
  NO2        g879(.A(new_new_n901_), .B(new_new_n376_), .Y(new_new_n902_));
  NO2        g880(.A(new_new_n566_), .B(new_new_n109_), .Y(new_new_n903_));
  AOI220     g881(.A0(new_new_n903_), .A1(i_0_), .B0(new_new_n902_), .B1(new_new_n589_), .Y(new_new_n904_));
  OAI220     g882(.A0(new_new_n904_), .A1(new_new_n87_), .B0(new_new_n900_), .B1(new_new_n174_), .Y(new_new_n905_));
  NO3        g883(.A(new_new_n905_), .B(new_new_n898_), .C(new_new_n487_), .Y(new_new_n906_));
  NA4        g884(.A(new_new_n906_), .B(new_new_n894_), .C(new_new_n891_), .D(new_new_n888_), .Y(new_new_n907_));
  NO3        g885(.A(new_new_n907_), .B(new_new_n884_), .C(new_new_n857_), .Y(new_new_n908_));
  NO2        g886(.A(i_0_), .B(new_new_n694_), .Y(new_new_n909_));
  NA2        g887(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n910_));
  INV        g888(.A(new_new_n910_), .Y(new_new_n911_));
  NO3        g889(.A(new_new_n109_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n912_));
  AO220      g890(.A0(new_new_n912_), .A1(new_new_n911_), .B0(new_new_n909_), .B1(new_new_n176_), .Y(new_new_n913_));
  AOI210     g891(.A0(new_new_n767_), .A1(new_new_n654_), .B0(new_new_n874_), .Y(new_new_n914_));
  AOI210     g892(.A0(new_new_n913_), .A1(new_new_n331_), .B0(new_new_n914_), .Y(new_new_n915_));
  NA2        g893(.A(new_new_n704_), .B(new_new_n151_), .Y(new_new_n916_));
  INV        g894(.A(new_new_n916_), .Y(new_new_n917_));
  NA3        g895(.A(new_new_n917_), .B(new_new_n641_), .C(new_new_n74_), .Y(new_new_n918_));
  NO2        g896(.A(new_new_n785_), .B(new_new_n376_), .Y(new_new_n919_));
  NA3        g897(.A(new_new_n810_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n920_));
  NA2        g898(.A(new_new_n811_), .B(i_9_), .Y(new_new_n921_));
  AOI210     g899(.A0(new_new_n920_), .A1(new_new_n464_), .B0(new_new_n921_), .Y(new_new_n922_));
  OAI210     g900(.A0(new_new_n240_), .A1(i_9_), .B0(new_new_n226_), .Y(new_new_n923_));
  AOI210     g901(.A0(new_new_n923_), .A1(new_new_n840_), .B0(new_new_n159_), .Y(new_new_n924_));
  NO3        g902(.A(new_new_n924_), .B(new_new_n922_), .C(new_new_n919_), .Y(new_new_n925_));
  NA3        g903(.A(new_new_n925_), .B(new_new_n918_), .C(new_new_n915_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n886_), .B(new_new_n355_), .Y(new_new_n927_));
  AOI210     g905(.A0(new_new_n287_), .A1(new_new_n166_), .B0(new_new_n927_), .Y(new_new_n928_));
  NA3        g906(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n929_));
  NA2        g907(.A(new_new_n862_), .B(new_new_n454_), .Y(new_new_n930_));
  AOI210     g908(.A0(new_new_n929_), .A1(new_new_n166_), .B0(new_new_n930_), .Y(new_new_n931_));
  NO2        g909(.A(new_new_n931_), .B(new_new_n928_), .Y(new_new_n932_));
  NO3        g910(.A(new_new_n848_), .B(new_new_n825_), .C(new_new_n190_), .Y(new_new_n933_));
  AOI220     g911(.A0(new_new_n933_), .A1(i_11_), .B0(new_new_n536_), .B1(new_new_n76_), .Y(new_new_n934_));
  NO3        g912(.A(new_new_n208_), .B(new_new_n364_), .C(i_0_), .Y(new_new_n935_));
  OAI210     g913(.A0(new_new_n935_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n936_));
  INV        g914(.A(new_new_n217_), .Y(new_new_n937_));
  OAI220     g915(.A0(new_new_n497_), .A1(new_new_n144_), .B0(new_new_n611_), .B1(new_new_n583_), .Y(new_new_n938_));
  NA3        g916(.A(new_new_n938_), .B(new_new_n372_), .C(new_new_n937_), .Y(new_new_n939_));
  NA4        g917(.A(new_new_n939_), .B(new_new_n936_), .C(new_new_n934_), .D(new_new_n932_), .Y(new_new_n940_));
  NO2        g918(.A(new_new_n239_), .B(new_new_n96_), .Y(new_new_n941_));
  AOI210     g919(.A0(new_new_n941_), .A1(new_new_n909_), .B0(new_new_n113_), .Y(new_new_n942_));
  AOI220     g920(.A0(new_new_n876_), .A1(new_new_n454_), .B0(new_new_n810_), .B1(new_new_n167_), .Y(new_new_n943_));
  NA2        g921(.A(new_new_n334_), .B(new_new_n178_), .Y(new_new_n944_));
  OA220      g922(.A0(new_new_n944_), .A1(new_new_n943_), .B0(new_new_n942_), .B1(i_5_), .Y(new_new_n945_));
  AOI210     g923(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n177_), .Y(new_new_n946_));
  NA2        g924(.A(new_new_n946_), .B(new_new_n890_), .Y(new_new_n947_));
  NA3        g925(.A(new_new_n580_), .B(new_new_n185_), .C(new_new_n85_), .Y(new_new_n948_));
  NA2        g926(.A(new_new_n948_), .B(new_new_n510_), .Y(new_new_n949_));
  NA2        g927(.A(new_new_n459_), .B(new_new_n452_), .Y(new_new_n950_));
  NO2        g928(.A(new_new_n950_), .B(new_new_n949_), .Y(new_new_n951_));
  NA3        g929(.A(new_new_n369_), .B(new_new_n173_), .C(new_new_n172_), .Y(new_new_n952_));
  NA3        g930(.A(new_new_n862_), .B(new_new_n281_), .C(new_new_n226_), .Y(new_new_n953_));
  NA2        g931(.A(new_new_n953_), .B(new_new_n952_), .Y(new_new_n954_));
  NO3        g932(.A(new_new_n859_), .B(new_new_n217_), .C(new_new_n190_), .Y(new_new_n955_));
  NO2        g933(.A(new_new_n955_), .B(new_new_n954_), .Y(new_new_n956_));
  NA4        g934(.A(new_new_n956_), .B(new_new_n951_), .C(new_new_n947_), .D(new_new_n945_), .Y(new_new_n957_));
  INV        g935(.A(new_new_n582_), .Y(new_new_n958_));
  NO3        g936(.A(new_new_n958_), .B(new_new_n526_), .C(new_new_n328_), .Y(new_new_n959_));
  NO2        g937(.A(new_new_n87_), .B(i_5_), .Y(new_new_n960_));
  NA3        g938(.A(new_new_n811_), .B(new_new_n114_), .C(new_new_n129_), .Y(new_new_n961_));
  INV        g939(.A(new_new_n961_), .Y(new_new_n962_));
  AOI210     g940(.A0(new_new_n962_), .A1(new_new_n960_), .B0(new_new_n959_), .Y(new_new_n963_));
  NA2        g941(.A(new_new_n292_), .B(i_5_), .Y(new_new_n964_));
  NAi31      g942(.An(new_new_n238_), .B(new_new_n964_), .C(new_new_n239_), .Y(new_new_n965_));
  NO4        g943(.A(new_new_n236_), .B(new_new_n208_), .C(i_0_), .D(i_12_), .Y(new_new_n966_));
  AOI220     g944(.A0(new_new_n966_), .A1(new_new_n965_), .B0(new_new_n761_), .B1(new_new_n178_), .Y(new_new_n967_));
  NA2        g945(.A(new_new_n876_), .B(new_new_n437_), .Y(new_new_n968_));
  NA2        g946(.A(new_new_n65_), .B(new_new_n105_), .Y(new_new_n969_));
  OAI220     g947(.A0(new_new_n969_), .A1(new_new_n964_), .B0(new_new_n968_), .B1(new_new_n642_), .Y(new_new_n970_));
  NA2        g948(.A(new_new_n970_), .B(new_new_n866_), .Y(new_new_n971_));
  NA3        g949(.A(new_new_n971_), .B(new_new_n967_), .C(new_new_n963_), .Y(new_new_n972_));
  NO4        g950(.A(new_new_n972_), .B(new_new_n957_), .C(new_new_n940_), .D(new_new_n926_), .Y(new_new_n973_));
  INV        g951(.A(new_new_n578_), .Y(new_new_n974_));
  NA2        g952(.A(new_new_n974_), .B(new_new_n204_), .Y(new_new_n975_));
  OAI210     g953(.A0(new_new_n582_), .A1(new_new_n580_), .B0(new_new_n302_), .Y(new_new_n976_));
  INV        g954(.A(new_new_n976_), .Y(new_new_n977_));
  NO4        g955(.A(new_new_n229_), .B(new_new_n150_), .C(new_new_n645_), .D(new_new_n37_), .Y(new_new_n978_));
  AOI210     g956(.A0(new_new_n977_), .A1(new_new_n49_), .B0(new_new_n978_), .Y(new_new_n979_));
  AOI210     g957(.A0(new_new_n979_), .A1(new_new_n975_), .B0(new_new_n74_), .Y(new_new_n980_));
  NO2        g958(.A(new_new_n533_), .B(new_new_n361_), .Y(new_new_n981_));
  NO2        g959(.A(new_new_n981_), .B(new_new_n723_), .Y(new_new_n982_));
  AOI210     g960(.A0(new_new_n946_), .A1(new_new_n862_), .B0(new_new_n877_), .Y(new_new_n983_));
  NO2        g961(.A(new_new_n983_), .B(new_new_n645_), .Y(new_new_n984_));
  NA2        g962(.A(new_new_n260_), .B(new_new_n58_), .Y(new_new_n985_));
  AOI220     g963(.A0(new_new_n985_), .A1(new_new_n77_), .B0(new_new_n329_), .B1(new_new_n252_), .Y(new_new_n986_));
  NO2        g964(.A(new_new_n986_), .B(new_new_n233_), .Y(new_new_n987_));
  NA3        g965(.A(new_new_n100_), .B(new_new_n294_), .C(new_new_n31_), .Y(new_new_n988_));
  INV        g966(.A(new_new_n988_), .Y(new_new_n989_));
  NO3        g967(.A(new_new_n989_), .B(new_new_n987_), .C(new_new_n984_), .Y(new_new_n990_));
  NA2        g968(.A(new_new_n268_), .B(new_new_n90_), .Y(new_new_n991_));
  NA3        g969(.A(new_new_n727_), .B(new_new_n281_), .C(new_new_n81_), .Y(new_new_n992_));
  AOI210     g970(.A0(new_new_n992_), .A1(new_new_n991_), .B0(i_11_), .Y(new_new_n993_));
  NO3        g971(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n994_));
  OAI210     g972(.A0(new_new_n881_), .A1(new_new_n294_), .B0(new_new_n994_), .Y(new_new_n995_));
  NO2        g973(.A(new_new_n995_), .B(new_new_n694_), .Y(new_new_n996_));
  NO4        g974(.A(new_new_n901_), .B(new_new_n442_), .C(new_new_n249_), .D(new_new_n248_), .Y(new_new_n997_));
  NO2        g975(.A(new_new_n997_), .B(new_new_n530_), .Y(new_new_n998_));
  INV        g976(.A(new_new_n347_), .Y(new_new_n999_));
  AOI210     g977(.A0(new_new_n999_), .A1(new_new_n998_), .B0(new_new_n41_), .Y(new_new_n1000_));
  NO3        g978(.A(new_new_n1000_), .B(new_new_n996_), .C(new_new_n993_), .Y(new_new_n1001_));
  OAI210     g979(.A0(new_new_n990_), .A1(i_4_), .B0(new_new_n1001_), .Y(new_new_n1002_));
  NO3        g980(.A(new_new_n1002_), .B(new_new_n982_), .C(new_new_n980_), .Y(new_new_n1003_));
  NA4        g981(.A(new_new_n1003_), .B(new_new_n973_), .C(new_new_n908_), .D(new_new_n833_), .Y(mai4));
  INV        g982(.A(new_new_n449_), .Y(new_new_n1007_));
endmodule


