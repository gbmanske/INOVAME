// Benchmark "top" written by ABC on Fri Jun 21 17:49:20 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1029_, new_new_n1030_, new_new_n1031_,
    new_new_n1032_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  NO2        g0029(.A(new_new_n48_), .B(new_new_n47_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g0032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  OAI210     g0033(.A0(new_new_n55_), .A1(new_new_n52_), .B0(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(new_new_n65_), .B(new_new_n61_), .Y(new_new_n66_));
  NA2        g0044(.A(new_new_n51_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g0046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g0047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g0048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g0049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g0050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g0051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g0052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  OAI210     g0053(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n75_), .Y(new_new_n76_));
  OAI210     g0054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g0055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g0056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g0057(.A(new_new_n79_), .B(new_new_n58_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_9_), .Y(new_new_n81_));
  NO2        g0059(.A(i_3_), .B(i_7_), .Y(new_new_n82_));
  INV        g0060(.A(i_6_), .Y(new_new_n83_));
  OR4        g0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n84_));
  INV        g0062(.A(new_new_n84_), .Y(new_new_n85_));
  NO2        g0063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  NA2        g0064(.A(new_new_n80_), .B(i_2_), .Y(new_new_n87_));
  NAi21      g0065(.An(i_6_), .B(i_10_), .Y(new_new_n88_));
  NA2        g0066(.A(i_6_), .B(i_9_), .Y(new_new_n89_));
  AOI210     g0067(.A0(new_new_n89_), .A1(new_new_n88_), .B0(new_new_n63_), .Y(new_new_n90_));
  NA2        g0068(.A(i_2_), .B(i_6_), .Y(new_new_n91_));
  NO3        g0069(.A(new_new_n91_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n92_));
  NO2        g0070(.A(new_new_n92_), .B(new_new_n90_), .Y(new_new_n93_));
  AOI210     g0071(.A0(new_new_n93_), .A1(new_new_n87_), .B0(new_new_n78_), .Y(new_new_n94_));
  AN3        g0072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n95_));
  NAi21      g0073(.An(i_6_), .B(i_11_), .Y(new_new_n96_));
  NO2        g0074(.A(i_5_), .B(i_8_), .Y(new_new_n97_));
  NOi21      g0075(.An(new_new_n97_), .B(new_new_n96_), .Y(new_new_n98_));
  AOI220     g0076(.A0(new_new_n98_), .A1(new_new_n62_), .B0(new_new_n95_), .B1(new_new_n32_), .Y(new_new_n99_));
  INV        g0077(.A(i_7_), .Y(new_new_n100_));
  NA2        g0078(.A(new_new_n47_), .B(new_new_n100_), .Y(new_new_n101_));
  NO2        g0079(.A(i_0_), .B(i_5_), .Y(new_new_n102_));
  NO2        g0080(.A(new_new_n102_), .B(new_new_n83_), .Y(new_new_n103_));
  NA2        g0081(.A(i_12_), .B(i_3_), .Y(new_new_n104_));
  INV        g0082(.A(new_new_n104_), .Y(new_new_n105_));
  NA3        g0083(.A(new_new_n105_), .B(new_new_n103_), .C(new_new_n101_), .Y(new_new_n106_));
  NAi21      g0084(.An(i_7_), .B(i_11_), .Y(new_new_n107_));
  NO3        g0085(.A(new_new_n107_), .B(new_new_n88_), .C(new_new_n53_), .Y(new_new_n108_));
  AN2        g0086(.A(i_2_), .B(i_10_), .Y(new_new_n109_));
  NO2        g0087(.A(new_new_n109_), .B(i_7_), .Y(new_new_n110_));
  OR2        g0088(.A(new_new_n78_), .B(new_new_n58_), .Y(new_new_n111_));
  NO2        g0089(.A(i_8_), .B(new_new_n100_), .Y(new_new_n112_));
  NO3        g0090(.A(new_new_n112_), .B(new_new_n111_), .C(new_new_n110_), .Y(new_new_n113_));
  NA2        g0091(.A(i_12_), .B(i_7_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n115_));
  NA2        g0093(.A(new_new_n115_), .B(i_0_), .Y(new_new_n116_));
  NA2        g0094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  OAI210     g0095(.A0(new_new_n116_), .A1(new_new_n114_), .B0(new_new_n117_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n118_), .B(new_new_n113_), .Y(new_new_n119_));
  NAi41      g0097(.An(new_new_n108_), .B(new_new_n119_), .C(new_new_n106_), .D(new_new_n99_), .Y(new_new_n120_));
  NOi21      g0098(.An(i_1_), .B(i_5_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n121_), .B(i_11_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n100_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g0101(.A(i_7_), .B(new_new_n25_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(new_new_n123_), .Y(new_new_n125_));
  NO2        g0103(.A(new_new_n125_), .B(new_new_n47_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n89_), .B(new_new_n88_), .Y(new_new_n127_));
  NAi21      g0105(.An(i_3_), .B(i_8_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n62_), .Y(new_new_n129_));
  NOi21      g0107(.An(new_new_n129_), .B(new_new_n127_), .Y(new_new_n130_));
  NO2        g0108(.A(i_1_), .B(new_new_n83_), .Y(new_new_n131_));
  NO2        g0109(.A(i_6_), .B(i_5_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(i_3_), .Y(new_new_n133_));
  AO210      g0111(.A0(new_new_n133_), .A1(new_new_n48_), .B0(new_new_n131_), .Y(new_new_n134_));
  OAI220     g0112(.A0(new_new_n134_), .A1(new_new_n107_), .B0(new_new_n130_), .B1(new_new_n122_), .Y(new_new_n135_));
  NO3        g0113(.A(new_new_n135_), .B(new_new_n120_), .C(new_new_n94_), .Y(new_new_n136_));
  NA3        g0114(.A(new_new_n136_), .B(new_new_n77_), .C(new_new_n56_), .Y(mai2));
  NO2        g0115(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n138_));
  NA2        g0116(.A(i_6_), .B(new_new_n25_), .Y(new_new_n139_));
  NA2        g0117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g0118(.A(new_new_n140_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(mai0));
  AN2        g0119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g0121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g0122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g0123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g0124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g0125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NO2        g0126(.A(new_new_n148_), .B(i_4_), .Y(new_new_n149_));
  NA3        g0127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  AN2        g0128(.A(new_new_n144_), .B(new_new_n81_), .Y(new_new_n151_));
  NA2        g0129(.A(i_1_), .B(i_5_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n71_), .B(new_new_n47_), .Y(new_new_n153_));
  NA2        g0131(.A(new_new_n153_), .B(new_new_n36_), .Y(new_new_n154_));
  NO3        g0132(.A(new_new_n154_), .B(new_new_n152_), .C(i_13_), .Y(new_new_n155_));
  OR2        g0133(.A(i_0_), .B(i_1_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n156_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n157_));
  NAi32      g0135(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n158_));
  NAi21      g0136(.An(new_new_n158_), .B(new_new_n157_), .Y(new_new_n159_));
  NOi21      g0137(.An(i_4_), .B(i_10_), .Y(new_new_n160_));
  NA2        g0138(.A(new_new_n160_), .B(new_new_n40_), .Y(new_new_n161_));
  NO2        g0139(.A(i_3_), .B(i_5_), .Y(new_new_n162_));
  NO3        g0140(.A(new_new_n71_), .B(i_2_), .C(i_1_), .Y(new_new_n163_));
  NA2        g0141(.A(new_new_n163_), .B(new_new_n162_), .Y(new_new_n164_));
  OAI210     g0142(.A0(new_new_n164_), .A1(new_new_n161_), .B0(new_new_n159_), .Y(new_new_n165_));
  NO2        g0143(.A(new_new_n165_), .B(new_new_n155_), .Y(new_new_n166_));
  AOI210     g0144(.A0(new_new_n166_), .A1(new_new_n150_), .B0(new_new_n143_), .Y(new_new_n167_));
  NA3        g0145(.A(new_new_n71_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n168_));
  NOi21      g0146(.An(i_4_), .B(i_9_), .Y(new_new_n169_));
  NOi21      g0147(.An(i_11_), .B(i_13_), .Y(new_new_n170_));
  NA2        g0148(.A(new_new_n170_), .B(new_new_n169_), .Y(new_new_n171_));
  BUFFER     g0149(.A(new_new_n171_), .Y(new_new_n172_));
  NO2        g0150(.A(i_4_), .B(i_5_), .Y(new_new_n173_));
  NAi21      g0151(.An(i_12_), .B(i_11_), .Y(new_new_n174_));
  NO2        g0152(.A(new_new_n174_), .B(i_13_), .Y(new_new_n175_));
  NA2        g0153(.A(new_new_n175_), .B(new_new_n173_), .Y(new_new_n176_));
  AOI210     g0154(.A0(new_new_n176_), .A1(new_new_n172_), .B0(new_new_n168_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n71_), .B(new_new_n63_), .Y(new_new_n178_));
  NA2        g0156(.A(new_new_n178_), .B(new_new_n47_), .Y(new_new_n179_));
  NA2        g0157(.A(new_new_n36_), .B(i_5_), .Y(new_new_n180_));
  NAi31      g0158(.An(new_new_n180_), .B(new_new_n151_), .C(i_11_), .Y(new_new_n181_));
  NA2        g0159(.A(i_3_), .B(i_5_), .Y(new_new_n182_));
  AOI210     g0160(.A0(new_new_n171_), .A1(new_new_n181_), .B0(new_new_n179_), .Y(new_new_n183_));
  NO2        g0161(.A(new_new_n71_), .B(i_5_), .Y(new_new_n184_));
  NO2        g0162(.A(i_13_), .B(i_10_), .Y(new_new_n185_));
  NA3        g0163(.A(new_new_n185_), .B(new_new_n184_), .C(new_new_n45_), .Y(new_new_n186_));
  NO2        g0164(.A(i_2_), .B(i_1_), .Y(new_new_n187_));
  NA2        g0165(.A(new_new_n187_), .B(i_3_), .Y(new_new_n188_));
  NAi21      g0166(.An(i_4_), .B(i_12_), .Y(new_new_n189_));
  NO4        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n186_), .D(new_new_n25_), .Y(new_new_n190_));
  NO3        g0168(.A(new_new_n190_), .B(new_new_n183_), .C(new_new_n177_), .Y(new_new_n191_));
  INV        g0169(.A(i_8_), .Y(new_new_n192_));
  NA2        g0170(.A(i_8_), .B(i_6_), .Y(new_new_n193_));
  NO3        g0171(.A(i_3_), .B(new_new_n83_), .C(new_new_n49_), .Y(new_new_n194_));
  NA2        g0172(.A(new_new_n194_), .B(new_new_n112_), .Y(new_new_n195_));
  NO3        g0173(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n196_));
  NA3        g0174(.A(new_new_n196_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n197_));
  NO3        g0175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n198_));
  OAI210     g0176(.A0(new_new_n95_), .A1(i_12_), .B0(new_new_n198_), .Y(new_new_n199_));
  AOI210     g0177(.A0(new_new_n199_), .A1(new_new_n197_), .B0(new_new_n195_), .Y(new_new_n200_));
  NO2        g0178(.A(i_3_), .B(i_8_), .Y(new_new_n201_));
  NO3        g0179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n202_));
  NA3        g0180(.A(new_new_n202_), .B(new_new_n201_), .C(new_new_n40_), .Y(new_new_n203_));
  NO2        g0181(.A(i_13_), .B(i_9_), .Y(new_new_n204_));
  NA3        g0182(.A(new_new_n204_), .B(i_6_), .C(new_new_n192_), .Y(new_new_n205_));
  NAi21      g0183(.An(i_12_), .B(i_3_), .Y(new_new_n206_));
  NO2        g0184(.A(new_new_n45_), .B(i_5_), .Y(new_new_n207_));
  NO3        g0185(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n208_));
  NA3        g0186(.A(new_new_n208_), .B(new_new_n207_), .C(i_10_), .Y(new_new_n209_));
  OAI220     g0187(.A0(new_new_n209_), .A1(new_new_n205_), .B0(new_new_n58_), .B1(new_new_n203_), .Y(new_new_n210_));
  AOI210     g0188(.A0(new_new_n210_), .A1(i_7_), .B0(new_new_n200_), .Y(new_new_n211_));
  OAI220     g0189(.A0(new_new_n211_), .A1(i_4_), .B0(new_new_n193_), .B1(new_new_n191_), .Y(new_new_n212_));
  NAi21      g0190(.An(i_12_), .B(i_7_), .Y(new_new_n213_));
  NA3        g0191(.A(i_13_), .B(new_new_n192_), .C(i_10_), .Y(new_new_n214_));
  NO2        g0192(.A(new_new_n214_), .B(new_new_n213_), .Y(new_new_n215_));
  NA2        g0193(.A(i_0_), .B(i_5_), .Y(new_new_n216_));
  OAI220     g0194(.A0(new_new_n83_), .A1(new_new_n188_), .B0(new_new_n179_), .B1(new_new_n133_), .Y(new_new_n217_));
  NAi31      g0195(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n218_));
  NO2        g0196(.A(new_new_n36_), .B(i_13_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n220_));
  NA3        g0198(.A(new_new_n220_), .B(i_0_), .C(new_new_n219_), .Y(new_new_n221_));
  INV        g0199(.A(i_13_), .Y(new_new_n222_));
  NO2        g0200(.A(i_12_), .B(new_new_n222_), .Y(new_new_n223_));
  NA3        g0201(.A(new_new_n223_), .B(new_new_n196_), .C(new_new_n194_), .Y(new_new_n224_));
  OAI210     g0202(.A0(new_new_n221_), .A1(new_new_n218_), .B0(new_new_n224_), .Y(new_new_n225_));
  AOI220     g0203(.A0(new_new_n225_), .A1(new_new_n142_), .B0(new_new_n217_), .B1(new_new_n215_), .Y(new_new_n226_));
  NO2        g0204(.A(i_12_), .B(new_new_n37_), .Y(new_new_n227_));
  NO2        g0205(.A(new_new_n182_), .B(i_4_), .Y(new_new_n228_));
  NA2        g0206(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n229_));
  OR2        g0207(.A(i_8_), .B(i_7_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n230_), .B(new_new_n83_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n53_), .B(i_1_), .Y(new_new_n232_));
  INV        g0210(.A(i_12_), .Y(new_new_n233_));
  NO3        g0211(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n234_));
  NA2        g0212(.A(i_2_), .B(i_1_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n230_), .B(new_new_n229_), .Y(new_new_n236_));
  NO3        g0214(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n237_));
  NAi21      g0215(.An(i_4_), .B(i_3_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n238_), .B(new_new_n73_), .Y(new_new_n239_));
  NO2        g0217(.A(i_0_), .B(i_6_), .Y(new_new_n240_));
  NOi41      g0218(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n241_));
  NA2        g0219(.A(new_new_n241_), .B(new_new_n240_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n235_), .B(new_new_n182_), .Y(new_new_n243_));
  NAi21      g0221(.An(new_new_n242_), .B(new_new_n243_), .Y(new_new_n244_));
  INV        g0222(.A(new_new_n244_), .Y(new_new_n245_));
  AOI220     g0223(.A0(new_new_n245_), .A1(new_new_n40_), .B0(new_new_n236_), .B1(new_new_n204_), .Y(new_new_n246_));
  NO2        g0224(.A(i_11_), .B(new_new_n222_), .Y(new_new_n247_));
  NOi21      g0225(.An(i_1_), .B(i_6_), .Y(new_new_n248_));
  NAi21      g0226(.An(i_3_), .B(i_7_), .Y(new_new_n249_));
  NO2        g0227(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n250_));
  NO2        g0228(.A(i_12_), .B(i_3_), .Y(new_new_n251_));
  NAi21      g0229(.An(i_7_), .B(i_10_), .Y(new_new_n252_));
  NA3        g0230(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n253_));
  INV        g0231(.A(new_new_n143_), .Y(new_new_n254_));
  NA2        g0232(.A(new_new_n233_), .B(i_13_), .Y(new_new_n255_));
  NO2        g0233(.A(new_new_n255_), .B(new_new_n73_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n256_), .B(new_new_n254_), .Y(new_new_n257_));
  NO2        g0235(.A(new_new_n230_), .B(new_new_n37_), .Y(new_new_n258_));
  NA2        g0236(.A(i_12_), .B(i_6_), .Y(new_new_n259_));
  OR2        g0237(.A(i_13_), .B(i_9_), .Y(new_new_n260_));
  NO3        g0238(.A(new_new_n260_), .B(new_new_n259_), .C(new_new_n49_), .Y(new_new_n261_));
  NO2        g0239(.A(new_new_n238_), .B(i_2_), .Y(new_new_n262_));
  NA3        g0240(.A(new_new_n262_), .B(new_new_n261_), .C(new_new_n45_), .Y(new_new_n263_));
  NA2        g0241(.A(new_new_n247_), .B(i_9_), .Y(new_new_n264_));
  OAI210     g0242(.A0(new_new_n63_), .A1(new_new_n264_), .B0(new_new_n263_), .Y(new_new_n265_));
  NA2        g0243(.A(new_new_n153_), .B(new_new_n63_), .Y(new_new_n266_));
  NO3        g0244(.A(i_11_), .B(new_new_n222_), .C(new_new_n25_), .Y(new_new_n267_));
  NO2        g0245(.A(new_new_n249_), .B(i_8_), .Y(new_new_n268_));
  NO2        g0246(.A(i_6_), .B(new_new_n49_), .Y(new_new_n269_));
  NA3        g0247(.A(new_new_n269_), .B(new_new_n268_), .C(new_new_n267_), .Y(new_new_n270_));
  NO3        g0248(.A(new_new_n26_), .B(new_new_n83_), .C(i_5_), .Y(new_new_n271_));
  NA3        g0249(.A(new_new_n271_), .B(new_new_n258_), .C(new_new_n223_), .Y(new_new_n272_));
  AOI210     g0250(.A0(new_new_n272_), .A1(new_new_n270_), .B0(new_new_n266_), .Y(new_new_n273_));
  AOI210     g0251(.A0(new_new_n265_), .A1(new_new_n258_), .B0(new_new_n273_), .Y(new_new_n274_));
  NA4        g0252(.A(new_new_n274_), .B(new_new_n257_), .C(new_new_n246_), .D(new_new_n226_), .Y(new_new_n275_));
  NO3        g0253(.A(i_12_), .B(new_new_n222_), .C(new_new_n37_), .Y(new_new_n276_));
  INV        g0254(.A(new_new_n276_), .Y(new_new_n277_));
  NA2        g0255(.A(i_8_), .B(new_new_n100_), .Y(new_new_n278_));
  NO3        g0256(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n279_));
  AOI220     g0257(.A0(new_new_n279_), .A1(new_new_n194_), .B0(new_new_n162_), .B1(new_new_n232_), .Y(new_new_n280_));
  NO2        g0258(.A(new_new_n280_), .B(new_new_n278_), .Y(new_new_n281_));
  NO2        g0259(.A(new_new_n235_), .B(i_0_), .Y(new_new_n282_));
  AOI220     g0260(.A0(new_new_n282_), .A1(i_8_), .B0(i_1_), .B1(new_new_n142_), .Y(new_new_n283_));
  NA2        g0261(.A(new_new_n269_), .B(new_new_n26_), .Y(new_new_n284_));
  NO2        g0262(.A(new_new_n284_), .B(new_new_n283_), .Y(new_new_n285_));
  NA2        g0263(.A(i_0_), .B(i_1_), .Y(new_new_n286_));
  NO2        g0264(.A(new_new_n286_), .B(i_2_), .Y(new_new_n287_));
  NO2        g0265(.A(new_new_n59_), .B(i_6_), .Y(new_new_n288_));
  NA2        g0266(.A(new_new_n288_), .B(new_new_n287_), .Y(new_new_n289_));
  OAI210     g0267(.A0(new_new_n164_), .A1(new_new_n143_), .B0(new_new_n289_), .Y(new_new_n290_));
  NO3        g0268(.A(new_new_n290_), .B(new_new_n285_), .C(new_new_n281_), .Y(new_new_n291_));
  NO2        g0269(.A(i_3_), .B(i_10_), .Y(new_new_n292_));
  NA3        g0270(.A(new_new_n292_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n293_));
  NO2        g0271(.A(i_2_), .B(new_new_n100_), .Y(new_new_n294_));
  NA2        g0272(.A(i_1_), .B(new_new_n36_), .Y(new_new_n295_));
  NA3        g0273(.A(new_new_n216_), .B(i_1_), .C(new_new_n294_), .Y(new_new_n296_));
  AN2        g0274(.A(i_3_), .B(i_10_), .Y(new_new_n297_));
  NA4        g0275(.A(new_new_n297_), .B(new_new_n196_), .C(new_new_n175_), .D(new_new_n173_), .Y(new_new_n298_));
  NO2        g0276(.A(i_5_), .B(new_new_n37_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n300_));
  OR2        g0278(.A(new_new_n296_), .B(new_new_n293_), .Y(new_new_n301_));
  OAI220     g0279(.A0(new_new_n301_), .A1(i_6_), .B0(new_new_n291_), .B1(new_new_n277_), .Y(new_new_n302_));
  NO4        g0280(.A(new_new_n302_), .B(new_new_n275_), .C(new_new_n212_), .D(new_new_n167_), .Y(new_new_n303_));
  NO3        g0281(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n59_), .B(new_new_n83_), .Y(new_new_n305_));
  NA2        g0283(.A(new_new_n282_), .B(new_new_n305_), .Y(new_new_n306_));
  NO3        g0284(.A(i_6_), .B(new_new_n192_), .C(i_7_), .Y(new_new_n307_));
  NA2        g0285(.A(new_new_n307_), .B(new_new_n196_), .Y(new_new_n308_));
  AOI210     g0286(.A0(new_new_n308_), .A1(new_new_n306_), .B0(i_5_), .Y(new_new_n309_));
  NO2        g0287(.A(i_2_), .B(i_3_), .Y(new_new_n310_));
  OR2        g0288(.A(i_0_), .B(i_5_), .Y(new_new_n311_));
  NA2        g0289(.A(new_new_n216_), .B(new_new_n311_), .Y(new_new_n312_));
  NA4        g0290(.A(new_new_n312_), .B(new_new_n231_), .C(new_new_n310_), .D(i_1_), .Y(new_new_n313_));
  NA3        g0291(.A(new_new_n282_), .B(new_new_n162_), .C(new_new_n112_), .Y(new_new_n314_));
  NAi21      g0292(.An(i_8_), .B(i_7_), .Y(new_new_n315_));
  NO2        g0293(.A(new_new_n315_), .B(i_6_), .Y(new_new_n316_));
  NO2        g0294(.A(new_new_n156_), .B(new_new_n47_), .Y(new_new_n317_));
  NA2        g0295(.A(new_new_n317_), .B(new_new_n316_), .Y(new_new_n318_));
  NA3        g0296(.A(new_new_n318_), .B(new_new_n314_), .C(new_new_n313_), .Y(new_new_n319_));
  OAI210     g0297(.A0(new_new_n319_), .A1(new_new_n309_), .B0(i_4_), .Y(new_new_n320_));
  NO2        g0298(.A(i_12_), .B(i_10_), .Y(new_new_n321_));
  NOi21      g0299(.An(i_5_), .B(i_0_), .Y(new_new_n322_));
  NO3        g0300(.A(new_new_n295_), .B(new_new_n322_), .C(new_new_n128_), .Y(new_new_n323_));
  NA4        g0301(.A(new_new_n82_), .B(new_new_n36_), .C(new_new_n83_), .D(i_8_), .Y(new_new_n324_));
  NA2        g0302(.A(new_new_n323_), .B(new_new_n321_), .Y(new_new_n325_));
  NO2        g0303(.A(i_6_), .B(i_8_), .Y(new_new_n326_));
  AN2        g0304(.A(i_0_), .B(new_new_n326_), .Y(new_new_n327_));
  NO2        g0305(.A(i_1_), .B(i_7_), .Y(new_new_n328_));
  NA3        g0306(.A(new_new_n326_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n329_));
  NA3        g0307(.A(new_new_n329_), .B(new_new_n325_), .C(new_new_n320_), .Y(new_new_n330_));
  NO3        g0308(.A(new_new_n230_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n331_));
  NO3        g0309(.A(new_new_n315_), .B(i_2_), .C(i_1_), .Y(new_new_n332_));
  OAI210     g0310(.A0(new_new_n332_), .A1(new_new_n331_), .B0(i_6_), .Y(new_new_n333_));
  NA3        g0311(.A(new_new_n248_), .B(new_new_n294_), .C(new_new_n192_), .Y(new_new_n334_));
  AOI210     g0312(.A0(new_new_n334_), .A1(new_new_n333_), .B0(new_new_n312_), .Y(new_new_n335_));
  NOi21      g0313(.An(new_new_n152_), .B(new_new_n103_), .Y(new_new_n336_));
  NO2        g0314(.A(new_new_n336_), .B(new_new_n124_), .Y(new_new_n337_));
  OAI210     g0315(.A0(new_new_n337_), .A1(new_new_n335_), .B0(i_3_), .Y(new_new_n338_));
  NO2        g0316(.A(new_new_n286_), .B(new_new_n79_), .Y(new_new_n339_));
  NA2        g0317(.A(new_new_n339_), .B(new_new_n132_), .Y(new_new_n340_));
  NO2        g0318(.A(new_new_n91_), .B(new_new_n192_), .Y(new_new_n341_));
  NA3        g0319(.A(new_new_n216_), .B(new_new_n341_), .C(new_new_n63_), .Y(new_new_n342_));
  AOI210     g0320(.A0(new_new_n342_), .A1(new_new_n340_), .B0(i_7_), .Y(new_new_n343_));
  NO2        g0321(.A(new_new_n192_), .B(i_9_), .Y(new_new_n344_));
  NA2        g0322(.A(new_new_n344_), .B(new_new_n156_), .Y(new_new_n345_));
  NO2        g0323(.A(new_new_n345_), .B(new_new_n47_), .Y(new_new_n346_));
  NO3        g0324(.A(new_new_n346_), .B(new_new_n343_), .C(new_new_n285_), .Y(new_new_n347_));
  AOI210     g0325(.A0(new_new_n347_), .A1(new_new_n338_), .B0(new_new_n161_), .Y(new_new_n348_));
  AOI210     g0326(.A0(new_new_n330_), .A1(new_new_n304_), .B0(new_new_n348_), .Y(new_new_n349_));
  NOi32      g0327(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n350_));
  INV        g0328(.A(new_new_n350_), .Y(new_new_n351_));
  NAi21      g0329(.An(i_0_), .B(i_6_), .Y(new_new_n352_));
  NAi21      g0330(.An(i_1_), .B(i_5_), .Y(new_new_n353_));
  NA2        g0331(.A(new_new_n353_), .B(new_new_n352_), .Y(new_new_n354_));
  NA2        g0332(.A(new_new_n354_), .B(new_new_n25_), .Y(new_new_n355_));
  OAI210     g0333(.A0(new_new_n355_), .A1(new_new_n158_), .B0(new_new_n242_), .Y(new_new_n356_));
  NAi41      g0334(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n357_));
  OAI220     g0335(.A0(new_new_n357_), .A1(new_new_n353_), .B0(new_new_n218_), .B1(new_new_n158_), .Y(new_new_n358_));
  AOI210     g0336(.A0(new_new_n357_), .A1(new_new_n158_), .B0(new_new_n156_), .Y(new_new_n359_));
  NOi32      g0337(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n360_));
  NAi21      g0338(.An(i_6_), .B(i_1_), .Y(new_new_n361_));
  NA3        g0339(.A(new_new_n361_), .B(new_new_n360_), .C(new_new_n47_), .Y(new_new_n362_));
  NO2        g0340(.A(new_new_n362_), .B(i_0_), .Y(new_new_n363_));
  OR3        g0341(.A(new_new_n363_), .B(new_new_n359_), .C(new_new_n358_), .Y(new_new_n364_));
  NO2        g0342(.A(i_1_), .B(new_new_n100_), .Y(new_new_n365_));
  NAi21      g0343(.An(i_3_), .B(i_4_), .Y(new_new_n366_));
  NO2        g0344(.A(new_new_n366_), .B(i_9_), .Y(new_new_n367_));
  NA2        g0345(.A(i_2_), .B(i_7_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n366_), .B(i_10_), .Y(new_new_n369_));
  NA3        g0347(.A(new_new_n369_), .B(new_new_n368_), .C(new_new_n240_), .Y(new_new_n370_));
  NO2        g0348(.A(new_new_n370_), .B(new_new_n184_), .Y(new_new_n371_));
  AOI210     g0349(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n372_));
  AOI220     g0350(.A0(new_new_n369_), .A1(new_new_n328_), .B0(new_new_n234_), .B1(new_new_n187_), .Y(new_new_n373_));
  NO2        g0351(.A(new_new_n373_), .B(i_5_), .Y(new_new_n374_));
  NO4        g0352(.A(new_new_n374_), .B(new_new_n371_), .C(new_new_n364_), .D(new_new_n356_), .Y(new_new_n375_));
  NO2        g0353(.A(new_new_n375_), .B(new_new_n351_), .Y(new_new_n376_));
  NO2        g0354(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n377_));
  AN2        g0355(.A(i_12_), .B(i_5_), .Y(new_new_n378_));
  NO2        g0356(.A(i_4_), .B(new_new_n26_), .Y(new_new_n379_));
  NA2        g0357(.A(new_new_n379_), .B(new_new_n378_), .Y(new_new_n380_));
  NO2        g0358(.A(i_11_), .B(i_6_), .Y(new_new_n381_));
  NA3        g0359(.A(new_new_n381_), .B(new_new_n317_), .C(new_new_n222_), .Y(new_new_n382_));
  NO2        g0360(.A(new_new_n382_), .B(new_new_n380_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n238_), .B(i_5_), .Y(new_new_n384_));
  NO2        g0362(.A(i_5_), .B(i_10_), .Y(new_new_n385_));
  NA2        g0363(.A(new_new_n144_), .B(new_new_n46_), .Y(new_new_n386_));
  NO2        g0364(.A(new_new_n386_), .B(new_new_n238_), .Y(new_new_n387_));
  OAI210     g0365(.A0(new_new_n387_), .A1(new_new_n383_), .B0(new_new_n377_), .Y(new_new_n388_));
  NO2        g0366(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n389_));
  NO2        g0367(.A(new_new_n150_), .B(new_new_n83_), .Y(new_new_n390_));
  OAI210     g0368(.A0(new_new_n390_), .A1(new_new_n383_), .B0(new_new_n389_), .Y(new_new_n391_));
  NO3        g0369(.A(new_new_n83_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n392_));
  NO2        g0370(.A(i_11_), .B(i_12_), .Y(new_new_n393_));
  NA2        g0371(.A(new_new_n393_), .B(new_new_n36_), .Y(new_new_n394_));
  NO2        g0372(.A(i_9_), .B(new_new_n394_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n385_), .B(new_new_n233_), .Y(new_new_n396_));
  OAI220     g0374(.A0(new_new_n36_), .A1(new_new_n218_), .B0(new_new_n396_), .B1(new_new_n324_), .Y(new_new_n397_));
  NAi21      g0375(.An(i_13_), .B(i_0_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n398_), .B(new_new_n235_), .Y(new_new_n399_));
  OAI210     g0377(.A0(new_new_n397_), .A1(new_new_n395_), .B0(new_new_n399_), .Y(new_new_n400_));
  NA3        g0378(.A(new_new_n400_), .B(new_new_n391_), .C(new_new_n388_), .Y(new_new_n401_));
  NO2        g0379(.A(i_0_), .B(i_11_), .Y(new_new_n402_));
  AN2        g0380(.A(i_1_), .B(i_6_), .Y(new_new_n403_));
  NOi21      g0381(.An(i_2_), .B(i_12_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n404_), .B(new_new_n403_), .Y(new_new_n405_));
  INV        g0383(.A(new_new_n405_), .Y(new_new_n406_));
  NA2        g0384(.A(new_new_n142_), .B(i_9_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(i_4_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n406_), .B(new_new_n408_), .Y(new_new_n409_));
  OR2        g0387(.A(i_13_), .B(i_10_), .Y(new_new_n410_));
  NO2        g0388(.A(new_new_n171_), .B(new_new_n123_), .Y(new_new_n411_));
  BUFFER     g0389(.A(new_new_n214_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n100_), .B(new_new_n25_), .Y(new_new_n413_));
  NA2        g0391(.A(new_new_n276_), .B(new_new_n413_), .Y(new_new_n414_));
  NA2        g0392(.A(new_new_n269_), .B(new_new_n208_), .Y(new_new_n415_));
  OAI220     g0393(.A0(new_new_n415_), .A1(new_new_n412_), .B0(new_new_n414_), .B1(new_new_n336_), .Y(new_new_n416_));
  INV        g0394(.A(new_new_n416_), .Y(new_new_n417_));
  AOI210     g0395(.A0(new_new_n417_), .A1(new_new_n409_), .B0(new_new_n26_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n314_), .B(new_new_n313_), .Y(new_new_n419_));
  AOI220     g0397(.A0(new_new_n288_), .A1(new_new_n279_), .B0(new_new_n282_), .B1(new_new_n305_), .Y(new_new_n420_));
  NO2        g0398(.A(new_new_n420_), .B(i_5_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n182_), .B(new_new_n83_), .Y(new_new_n422_));
  AOI220     g0400(.A0(new_new_n422_), .A1(new_new_n287_), .B0(new_new_n271_), .B1(new_new_n208_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n423_), .B(new_new_n278_), .Y(new_new_n424_));
  NO3        g0402(.A(new_new_n424_), .B(new_new_n421_), .C(new_new_n419_), .Y(new_new_n425_));
  NA2        g0403(.A(new_new_n194_), .B(new_new_n95_), .Y(new_new_n426_));
  NA3        g0404(.A(new_new_n317_), .B(new_new_n162_), .C(new_new_n83_), .Y(new_new_n427_));
  AOI210     g0405(.A0(new_new_n427_), .A1(new_new_n426_), .B0(new_new_n315_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n192_), .B(i_10_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n64_), .B(i_2_), .Y(new_new_n430_));
  NA2        g0408(.A(new_new_n288_), .B(new_new_n232_), .Y(new_new_n431_));
  OAI220     g0409(.A0(new_new_n431_), .A1(new_new_n182_), .B0(new_new_n430_), .B1(new_new_n429_), .Y(new_new_n432_));
  NO2        g0410(.A(i_3_), .B(new_new_n49_), .Y(new_new_n433_));
  NA3        g0411(.A(new_new_n328_), .B(new_new_n327_), .C(new_new_n433_), .Y(new_new_n434_));
  NA2        g0412(.A(new_new_n307_), .B(new_new_n312_), .Y(new_new_n435_));
  OAI210     g0413(.A0(new_new_n435_), .A1(new_new_n188_), .B0(new_new_n434_), .Y(new_new_n436_));
  NO3        g0414(.A(new_new_n436_), .B(new_new_n432_), .C(new_new_n428_), .Y(new_new_n437_));
  AOI210     g0415(.A0(new_new_n437_), .A1(new_new_n425_), .B0(new_new_n264_), .Y(new_new_n438_));
  NO4        g0416(.A(new_new_n438_), .B(new_new_n418_), .C(new_new_n401_), .D(new_new_n376_), .Y(new_new_n439_));
  NO2        g0417(.A(new_new_n71_), .B(i_13_), .Y(new_new_n440_));
  NO2        g0418(.A(i_10_), .B(i_9_), .Y(new_new_n441_));
  NAi21      g0419(.An(i_12_), .B(i_8_), .Y(new_new_n442_));
  NO2        g0420(.A(new_new_n442_), .B(i_3_), .Y(new_new_n443_));
  NA2        g0421(.A(i_2_), .B(new_new_n103_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n444_), .B(new_new_n203_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n300_), .B(i_0_), .Y(new_new_n446_));
  NO3        g0424(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n447_));
  NA2        g0425(.A(new_new_n259_), .B(new_new_n96_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n448_), .B(new_new_n447_), .Y(new_new_n449_));
  NA2        g0427(.A(i_8_), .B(i_9_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n449_), .B(new_new_n446_), .Y(new_new_n451_));
  NO3        g0429(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n452_));
  NA3        g0430(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n453_));
  NA4        g0431(.A(new_new_n145_), .B(new_new_n115_), .C(new_new_n78_), .D(new_new_n23_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n455_));
  NO3        g0433(.A(new_new_n455_), .B(new_new_n451_), .C(new_new_n445_), .Y(new_new_n456_));
  OA210      g0434(.A0(new_new_n345_), .A1(new_new_n100_), .B0(new_new_n289_), .Y(new_new_n457_));
  OA220      g0435(.A0(new_new_n457_), .A1(new_new_n161_), .B0(new_new_n205_), .B1(new_new_n229_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n95_), .B(i_13_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n422_), .B(new_new_n377_), .Y(new_new_n460_));
  NO2        g0438(.A(i_2_), .B(i_13_), .Y(new_new_n461_));
  NA3        g0439(.A(new_new_n461_), .B(new_new_n160_), .C(new_new_n98_), .Y(new_new_n462_));
  OAI220     g0440(.A0(new_new_n462_), .A1(new_new_n233_), .B0(new_new_n460_), .B1(new_new_n459_), .Y(new_new_n463_));
  NO3        g0441(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n464_));
  NO2        g0442(.A(i_6_), .B(i_7_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n465_), .B(new_new_n464_), .Y(new_new_n466_));
  NO2        g0444(.A(i_11_), .B(i_1_), .Y(new_new_n467_));
  OR2        g0445(.A(i_11_), .B(i_8_), .Y(new_new_n468_));
  NOi21      g0446(.An(i_2_), .B(i_7_), .Y(new_new_n469_));
  NAi31      g0447(.An(new_new_n468_), .B(new_new_n469_), .C(i_0_), .Y(new_new_n470_));
  NO2        g0448(.A(new_new_n410_), .B(i_6_), .Y(new_new_n471_));
  NA3        g0449(.A(new_new_n471_), .B(i_1_), .C(new_new_n73_), .Y(new_new_n472_));
  NO2        g0450(.A(new_new_n472_), .B(new_new_n470_), .Y(new_new_n473_));
  NO2        g0451(.A(i_3_), .B(new_new_n192_), .Y(new_new_n474_));
  NO2        g0452(.A(i_6_), .B(i_10_), .Y(new_new_n475_));
  NA4        g0453(.A(new_new_n475_), .B(new_new_n304_), .C(new_new_n474_), .D(new_new_n233_), .Y(new_new_n476_));
  NO2        g0454(.A(new_new_n476_), .B(new_new_n154_), .Y(new_new_n477_));
  NA2        g0455(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n478_));
  NO2        g0456(.A(new_new_n156_), .B(i_3_), .Y(new_new_n479_));
  NO3        g0457(.A(new_new_n477_), .B(new_new_n473_), .C(new_new_n463_), .Y(new_new_n480_));
  NA2        g0458(.A(new_new_n447_), .B(new_new_n378_), .Y(new_new_n481_));
  NA2        g0459(.A(new_new_n452_), .B(new_new_n385_), .Y(new_new_n482_));
  NO2        g0460(.A(new_new_n482_), .B(new_new_n221_), .Y(new_new_n483_));
  NAi21      g0461(.An(new_new_n214_), .B(new_new_n393_), .Y(new_new_n484_));
  NA2        g0462(.A(new_new_n328_), .B(new_new_n216_), .Y(new_new_n485_));
  NO2        g0463(.A(i_0_), .B(new_new_n83_), .Y(new_new_n486_));
  NA3        g0464(.A(new_new_n486_), .B(new_new_n1030_), .C(new_new_n142_), .Y(new_new_n487_));
  OR3        g0465(.A(new_new_n295_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n488_));
  OAI220     g0466(.A0(new_new_n488_), .A1(new_new_n487_), .B0(new_new_n485_), .B1(new_new_n484_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n27_), .B(i_10_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n304_), .B(new_new_n234_), .Y(new_new_n491_));
  OAI220     g0469(.A0(new_new_n491_), .A1(new_new_n430_), .B0(new_new_n490_), .B1(new_new_n459_), .Y(new_new_n492_));
  NA4        g0470(.A(new_new_n297_), .B(new_new_n220_), .C(new_new_n71_), .D(new_new_n233_), .Y(new_new_n493_));
  NO2        g0471(.A(new_new_n493_), .B(new_new_n466_), .Y(new_new_n494_));
  NO4        g0472(.A(new_new_n494_), .B(new_new_n492_), .C(new_new_n489_), .D(new_new_n483_), .Y(new_new_n495_));
  NA4        g0473(.A(new_new_n495_), .B(new_new_n480_), .C(new_new_n458_), .D(new_new_n456_), .Y(new_new_n496_));
  NA3        g0474(.A(new_new_n297_), .B(new_new_n175_), .C(new_new_n173_), .Y(new_new_n497_));
  OAI210     g0475(.A0(new_new_n293_), .A1(new_new_n180_), .B0(new_new_n497_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n231_), .B(new_new_n498_), .Y(new_new_n499_));
  NA2        g0477(.A(new_new_n122_), .B(new_new_n111_), .Y(new_new_n500_));
  AN2        g0478(.A(new_new_n500_), .B(new_new_n447_), .Y(new_new_n501_));
  INV        g0479(.A(new_new_n304_), .Y(new_new_n502_));
  OAI210     g0480(.A0(new_new_n502_), .A1(new_new_n229_), .B0(new_new_n298_), .Y(new_new_n503_));
  AOI220     g0481(.A0(new_new_n503_), .A1(new_new_n316_), .B0(new_new_n501_), .B1(new_new_n300_), .Y(new_new_n504_));
  NA2        g0482(.A(new_new_n350_), .B(new_new_n71_), .Y(new_new_n505_));
  INV        g0483(.A(new_new_n360_), .Y(new_new_n506_));
  NO2        g0484(.A(new_new_n36_), .B(i_8_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n39_), .B(i_13_), .Y(new_new_n508_));
  OAI210     g0486(.A0(i_8_), .A1(new_new_n63_), .B0(new_new_n134_), .Y(new_new_n509_));
  NO2        g0487(.A(i_7_), .B(new_new_n197_), .Y(new_new_n510_));
  OR2        g0488(.A(new_new_n182_), .B(i_4_), .Y(new_new_n511_));
  NO2        g0489(.A(new_new_n511_), .B(new_new_n83_), .Y(new_new_n512_));
  AOI220     g0490(.A0(new_new_n512_), .A1(new_new_n510_), .B0(new_new_n509_), .B1(new_new_n411_), .Y(new_new_n513_));
  NA4        g0491(.A(new_new_n513_), .B(new_new_n508_), .C(new_new_n504_), .D(new_new_n499_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n384_), .B(new_new_n287_), .Y(new_new_n515_));
  NA2        g0493(.A(new_new_n380_), .B(new_new_n515_), .Y(new_new_n516_));
  NO2        g0494(.A(i_12_), .B(new_new_n192_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n517_), .B(new_new_n222_), .Y(new_new_n518_));
  NO2        g0496(.A(i_10_), .B(new_new_n518_), .Y(new_new_n519_));
  NOi31      g0497(.An(new_new_n307_), .B(new_new_n410_), .C(new_new_n38_), .Y(new_new_n520_));
  OAI210     g0498(.A0(new_new_n520_), .A1(new_new_n519_), .B0(new_new_n516_), .Y(new_new_n521_));
  NO2        g0499(.A(i_8_), .B(i_7_), .Y(new_new_n522_));
  OAI210     g0500(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n523_), .B(new_new_n220_), .Y(new_new_n524_));
  OAI220     g0502(.A0(new_new_n47_), .A1(new_new_n511_), .B0(new_new_n524_), .B1(new_new_n238_), .Y(new_new_n525_));
  NA2        g0503(.A(new_new_n45_), .B(i_10_), .Y(new_new_n526_));
  NO2        g0504(.A(new_new_n526_), .B(i_6_), .Y(new_new_n527_));
  NA3        g0505(.A(new_new_n527_), .B(new_new_n525_), .C(new_new_n522_), .Y(new_new_n528_));
  AOI220     g0506(.A0(new_new_n422_), .A1(new_new_n317_), .B0(new_new_n243_), .B1(new_new_n240_), .Y(new_new_n529_));
  OAI220     g0507(.A0(new_new_n529_), .A1(new_new_n255_), .B0(new_new_n459_), .B1(new_new_n133_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n530_), .B(new_new_n258_), .Y(new_new_n531_));
  NOi31      g0509(.An(new_new_n282_), .B(new_new_n293_), .C(new_new_n180_), .Y(new_new_n532_));
  NA3        g0510(.A(new_new_n297_), .B(new_new_n173_), .C(new_new_n95_), .Y(new_new_n533_));
  NO2        g0511(.A(new_new_n156_), .B(i_5_), .Y(new_new_n534_));
  NA2        g0512(.A(new_new_n534_), .B(new_new_n310_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n535_), .B(new_new_n533_), .Y(new_new_n536_));
  OAI210     g0514(.A0(new_new_n536_), .A1(new_new_n532_), .B0(new_new_n452_), .Y(new_new_n537_));
  NA4        g0515(.A(new_new_n537_), .B(new_new_n531_), .C(new_new_n528_), .D(new_new_n521_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n276_), .B(new_new_n82_), .Y(new_new_n539_));
  NO2        g0517(.A(new_new_n340_), .B(new_new_n539_), .Y(new_new_n540_));
  NA2        g0518(.A(new_new_n288_), .B(new_new_n279_), .Y(new_new_n541_));
  NO2        g0519(.A(new_new_n541_), .B(new_new_n172_), .Y(new_new_n542_));
  NA2        g0520(.A(new_new_n220_), .B(i_0_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n441_), .B(new_new_n219_), .Y(new_new_n544_));
  NO2        g0522(.A(new_new_n543_), .B(new_new_n544_), .Y(new_new_n545_));
  AOI210     g0523(.A0(new_new_n361_), .A1(new_new_n47_), .B0(new_new_n365_), .Y(new_new_n546_));
  NA2        g0524(.A(i_0_), .B(new_new_n49_), .Y(new_new_n547_));
  NA3        g0525(.A(new_new_n517_), .B(new_new_n267_), .C(new_new_n547_), .Y(new_new_n548_));
  NO2        g0526(.A(new_new_n546_), .B(new_new_n548_), .Y(new_new_n549_));
  NO4        g0527(.A(new_new_n549_), .B(new_new_n545_), .C(new_new_n542_), .D(new_new_n540_), .Y(new_new_n550_));
  NO4        g0528(.A(new_new_n248_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n551_));
  NO3        g0529(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n552_));
  NO2        g0530(.A(new_new_n230_), .B(new_new_n36_), .Y(new_new_n553_));
  AN2        g0531(.A(new_new_n553_), .B(new_new_n552_), .Y(new_new_n554_));
  OA210      g0532(.A0(new_new_n554_), .A1(new_new_n551_), .B0(new_new_n350_), .Y(new_new_n555_));
  NO2        g0533(.A(new_new_n410_), .B(i_1_), .Y(new_new_n556_));
  NOi31      g0534(.An(new_new_n556_), .B(new_new_n448_), .C(new_new_n71_), .Y(new_new_n557_));
  AN3        g0535(.A(new_new_n557_), .B(new_new_n408_), .C(i_2_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n420_), .B(new_new_n176_), .Y(new_new_n559_));
  NO3        g0537(.A(new_new_n559_), .B(new_new_n558_), .C(new_new_n555_), .Y(new_new_n560_));
  NOi21      g0538(.An(i_10_), .B(i_6_), .Y(new_new_n561_));
  NO2        g0539(.A(new_new_n83_), .B(new_new_n25_), .Y(new_new_n562_));
  AOI220     g0540(.A0(new_new_n276_), .A1(new_new_n562_), .B0(new_new_n267_), .B1(new_new_n561_), .Y(new_new_n563_));
  NO2        g0541(.A(new_new_n563_), .B(new_new_n446_), .Y(new_new_n564_));
  NO2        g0542(.A(new_new_n114_), .B(new_new_n23_), .Y(new_new_n565_));
  NA2        g0543(.A(new_new_n307_), .B(new_new_n163_), .Y(new_new_n566_));
  AOI220     g0544(.A0(new_new_n566_), .A1(new_new_n431_), .B0(new_new_n171_), .B1(new_new_n181_), .Y(new_new_n567_));
  NOi21      g0545(.An(new_new_n146_), .B(new_new_n324_), .Y(new_new_n568_));
  NO3        g0546(.A(new_new_n568_), .B(new_new_n567_), .C(new_new_n564_), .Y(new_new_n569_));
  NO2        g0547(.A(new_new_n505_), .B(new_new_n373_), .Y(new_new_n570_));
  INV        g0548(.A(new_new_n310_), .Y(new_new_n571_));
  NO2        g0549(.A(i_12_), .B(new_new_n83_), .Y(new_new_n572_));
  NA3        g0550(.A(new_new_n572_), .B(new_new_n267_), .C(new_new_n547_), .Y(new_new_n573_));
  NA3        g0551(.A(new_new_n381_), .B(new_new_n276_), .C(new_new_n216_), .Y(new_new_n574_));
  AOI210     g0552(.A0(new_new_n574_), .A1(new_new_n573_), .B0(new_new_n571_), .Y(new_new_n575_));
  NO3        g0553(.A(i_4_), .B(new_new_n333_), .C(new_new_n293_), .Y(new_new_n576_));
  OR2        g0554(.A(i_2_), .B(i_5_), .Y(new_new_n577_));
  OR2        g0555(.A(new_new_n577_), .B(new_new_n403_), .Y(new_new_n578_));
  AOI210     g0556(.A0(new_new_n368_), .A1(new_new_n240_), .B0(new_new_n196_), .Y(new_new_n579_));
  AOI210     g0557(.A0(new_new_n579_), .A1(new_new_n578_), .B0(new_new_n484_), .Y(new_new_n580_));
  NO4        g0558(.A(new_new_n580_), .B(new_new_n576_), .C(new_new_n575_), .D(new_new_n570_), .Y(new_new_n581_));
  NA4        g0559(.A(new_new_n581_), .B(new_new_n569_), .C(new_new_n560_), .D(new_new_n550_), .Y(new_new_n582_));
  NO4        g0560(.A(new_new_n582_), .B(new_new_n538_), .C(new_new_n514_), .D(new_new_n496_), .Y(new_new_n583_));
  NA4        g0561(.A(new_new_n583_), .B(new_new_n439_), .C(new_new_n349_), .D(new_new_n303_), .Y(mai7));
  OAI220     g0562(.A0(new_new_n490_), .A1(new_new_n117_), .B0(new_new_n91_), .B1(new_new_n54_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n107_), .B(new_new_n88_), .Y(new_new_n586_));
  NA2        g0564(.A(new_new_n379_), .B(new_new_n586_), .Y(new_new_n587_));
  NA2        g0565(.A(new_new_n475_), .B(new_new_n82_), .Y(new_new_n588_));
  NA2        g0566(.A(i_11_), .B(new_new_n192_), .Y(new_new_n589_));
  NA2        g0567(.A(new_new_n144_), .B(new_new_n589_), .Y(new_new_n590_));
  OAI210     g0568(.A0(new_new_n590_), .A1(new_new_n588_), .B0(new_new_n587_), .Y(new_new_n591_));
  NA3        g0569(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n233_), .B(i_4_), .Y(new_new_n593_));
  NA2        g0571(.A(new_new_n593_), .B(i_8_), .Y(new_new_n594_));
  NA2        g0572(.A(i_2_), .B(new_new_n83_), .Y(new_new_n595_));
  OAI210     g0573(.A0(new_new_n86_), .A1(new_new_n201_), .B0(new_new_n202_), .Y(new_new_n596_));
  NO2        g0574(.A(i_7_), .B(new_new_n37_), .Y(new_new_n597_));
  NA2        g0575(.A(i_4_), .B(i_8_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n591_), .B(new_new_n585_), .Y(new_new_n599_));
  INV        g0577(.A(new_new_n160_), .Y(new_new_n600_));
  OR2        g0578(.A(i_6_), .B(i_10_), .Y(new_new_n601_));
  NO2        g0579(.A(new_new_n601_), .B(new_new_n23_), .Y(new_new_n602_));
  OR3        g0580(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n603_));
  NO3        g0581(.A(new_new_n603_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n604_));
  INV        g0582(.A(new_new_n198_), .Y(new_new_n605_));
  NO2        g0583(.A(new_new_n604_), .B(new_new_n602_), .Y(new_new_n606_));
  OA220      g0584(.A0(new_new_n606_), .A1(new_new_n571_), .B0(new_new_n600_), .B1(new_new_n260_), .Y(new_new_n607_));
  AOI210     g0585(.A0(new_new_n607_), .A1(new_new_n599_), .B0(new_new_n63_), .Y(new_new_n608_));
  NOi21      g0586(.An(i_11_), .B(i_7_), .Y(new_new_n609_));
  AO210      g0587(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n610_));
  NO2        g0588(.A(new_new_n610_), .B(new_new_n609_), .Y(new_new_n611_));
  NA2        g0589(.A(new_new_n611_), .B(new_new_n204_), .Y(new_new_n612_));
  NA3        g0590(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n613_));
  NAi31      g0591(.An(new_new_n613_), .B(new_new_n213_), .C(i_11_), .Y(new_new_n614_));
  AOI210     g0592(.A0(new_new_n614_), .A1(new_new_n612_), .B0(new_new_n63_), .Y(new_new_n615_));
  NA2        g0593(.A(new_new_n85_), .B(new_new_n63_), .Y(new_new_n616_));
  AO210      g0594(.A0(new_new_n616_), .A1(new_new_n373_), .B0(new_new_n41_), .Y(new_new_n617_));
  NO3        g0595(.A(new_new_n252_), .B(new_new_n206_), .C(new_new_n589_), .Y(new_new_n618_));
  OAI210     g0596(.A0(new_new_n618_), .A1(new_new_n223_), .B0(new_new_n63_), .Y(new_new_n619_));
  NA2        g0597(.A(new_new_n404_), .B(new_new_n31_), .Y(new_new_n620_));
  OR2        g0598(.A(new_new_n206_), .B(new_new_n107_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n621_), .B(new_new_n620_), .Y(new_new_n622_));
  NO2        g0600(.A(new_new_n63_), .B(i_9_), .Y(new_new_n623_));
  NO2        g0601(.A(new_new_n623_), .B(i_4_), .Y(new_new_n624_));
  NA2        g0602(.A(new_new_n624_), .B(new_new_n622_), .Y(new_new_n625_));
  NO2        g0603(.A(i_1_), .B(i_12_), .Y(new_new_n626_));
  NA3        g0604(.A(new_new_n626_), .B(new_new_n109_), .C(new_new_n24_), .Y(new_new_n627_));
  NA4        g0605(.A(new_new_n627_), .B(new_new_n625_), .C(new_new_n619_), .D(new_new_n617_), .Y(new_new_n628_));
  OAI210     g0606(.A0(new_new_n628_), .A1(new_new_n615_), .B0(i_6_), .Y(new_new_n629_));
  OAI210     g0607(.A0(new_new_n613_), .A1(new_new_n107_), .B0(new_new_n453_), .Y(new_new_n630_));
  NA2        g0608(.A(new_new_n630_), .B(new_new_n572_), .Y(new_new_n631_));
  NO2        g0609(.A(new_new_n233_), .B(new_new_n83_), .Y(new_new_n632_));
  NO2        g0610(.A(new_new_n632_), .B(i_11_), .Y(new_new_n633_));
  NA2        g0611(.A(new_new_n631_), .B(new_new_n449_), .Y(new_new_n634_));
  NO4        g0612(.A(new_new_n213_), .B(new_new_n128_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n635_));
  NA2        g0613(.A(new_new_n635_), .B(new_new_n623_), .Y(new_new_n636_));
  NO3        g0614(.A(new_new_n601_), .B(new_new_n230_), .C(new_new_n23_), .Y(new_new_n637_));
  INV        g0615(.A(new_new_n636_), .Y(new_new_n638_));
  NA3        g0616(.A(new_new_n522_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n639_));
  NA2        g0617(.A(new_new_n138_), .B(i_9_), .Y(new_new_n640_));
  NA3        g0618(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n641_));
  NO2        g0619(.A(new_new_n47_), .B(i_1_), .Y(new_new_n642_));
  NA3        g0620(.A(new_new_n642_), .B(new_new_n259_), .C(new_new_n45_), .Y(new_new_n643_));
  OAI220     g0621(.A0(new_new_n643_), .A1(new_new_n641_), .B0(new_new_n640_), .B1(new_new_n1029_), .Y(new_new_n644_));
  NA3        g0622(.A(new_new_n623_), .B(new_new_n310_), .C(i_6_), .Y(new_new_n645_));
  NO2        g0623(.A(new_new_n645_), .B(new_new_n23_), .Y(new_new_n646_));
  AOI210     g0624(.A0(new_new_n467_), .A1(new_new_n413_), .B0(new_new_n237_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n647_), .B(new_new_n595_), .Y(new_new_n648_));
  NAi21      g0626(.An(new_new_n639_), .B(new_new_n90_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n642_), .B(new_new_n259_), .Y(new_new_n650_));
  NO2        g0628(.A(i_11_), .B(new_new_n37_), .Y(new_new_n651_));
  NA2        g0629(.A(new_new_n651_), .B(new_new_n24_), .Y(new_new_n652_));
  OAI210     g0630(.A0(new_new_n652_), .A1(new_new_n650_), .B0(new_new_n649_), .Y(new_new_n653_));
  OR4        g0631(.A(new_new_n653_), .B(new_new_n648_), .C(new_new_n646_), .D(new_new_n644_), .Y(new_new_n654_));
  NO3        g0632(.A(new_new_n654_), .B(new_new_n638_), .C(new_new_n634_), .Y(new_new_n655_));
  NO2        g0633(.A(new_new_n233_), .B(new_new_n100_), .Y(new_new_n656_));
  NO2        g0634(.A(new_new_n656_), .B(new_new_n609_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n657_), .B(i_1_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n658_), .B(new_new_n603_), .Y(new_new_n659_));
  NA2        g0637(.A(new_new_n659_), .B(new_new_n47_), .Y(new_new_n660_));
  NA2        g0638(.A(i_3_), .B(new_new_n192_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n661_), .B(new_new_n114_), .Y(new_new_n662_));
  AN2        g0640(.A(new_new_n662_), .B(new_new_n527_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n83_), .B(i_9_), .Y(new_new_n665_));
  NA2        g0643(.A(i_1_), .B(i_3_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n450_), .B(new_new_n91_), .Y(new_new_n667_));
  AOI210     g0645(.A0(i_11_), .A1(new_new_n561_), .B0(new_new_n667_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n668_), .B(new_new_n666_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n669_), .B(new_new_n663_), .Y(new_new_n670_));
  NA4        g0648(.A(new_new_n670_), .B(new_new_n660_), .C(new_new_n655_), .D(new_new_n629_), .Y(new_new_n671_));
  NO3        g0649(.A(new_new_n468_), .B(i_3_), .C(i_7_), .Y(new_new_n672_));
  NOi21      g0650(.An(new_new_n672_), .B(i_10_), .Y(new_new_n673_));
  OA210      g0651(.A0(new_new_n673_), .A1(new_new_n241_), .B0(new_new_n83_), .Y(new_new_n674_));
  NA2        g0652(.A(i_6_), .B(new_new_n367_), .Y(new_new_n675_));
  NA3        g0653(.A(new_new_n475_), .B(new_new_n507_), .C(new_new_n47_), .Y(new_new_n676_));
  NO3        g0654(.A(new_new_n469_), .B(new_new_n598_), .C(new_new_n83_), .Y(new_new_n677_));
  NA2        g0655(.A(new_new_n677_), .B(new_new_n25_), .Y(new_new_n678_));
  NA3        g0656(.A(new_new_n160_), .B(new_new_n82_), .C(new_new_n83_), .Y(new_new_n679_));
  NA4        g0657(.A(new_new_n679_), .B(new_new_n678_), .C(new_new_n676_), .D(new_new_n675_), .Y(new_new_n680_));
  OAI210     g0658(.A0(new_new_n680_), .A1(new_new_n674_), .B0(i_1_), .Y(new_new_n681_));
  AOI210     g0659(.A0(new_new_n259_), .A1(new_new_n96_), .B0(i_1_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n366_), .B(i_2_), .Y(new_new_n683_));
  NA2        g0661(.A(new_new_n683_), .B(new_new_n682_), .Y(new_new_n684_));
  OAI210     g0662(.A0(new_new_n645_), .A1(new_new_n442_), .B0(new_new_n684_), .Y(new_new_n685_));
  INV        g0663(.A(new_new_n685_), .Y(new_new_n686_));
  AOI210     g0664(.A0(new_new_n686_), .A1(new_new_n681_), .B0(i_13_), .Y(new_new_n687_));
  OR2        g0665(.A(i_11_), .B(i_7_), .Y(new_new_n688_));
  NA3        g0666(.A(new_new_n688_), .B(new_new_n105_), .C(new_new_n138_), .Y(new_new_n689_));
  AOI220     g0667(.A0(new_new_n461_), .A1(new_new_n160_), .B0(i_2_), .B1(new_new_n138_), .Y(new_new_n690_));
  OAI210     g0668(.A0(new_new_n690_), .A1(new_new_n45_), .B0(new_new_n689_), .Y(new_new_n691_));
  NA2        g0669(.A(new_new_n241_), .B(new_new_n131_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n692_), .B(new_new_n41_), .Y(new_new_n693_));
  AOI210     g0671(.A0(new_new_n691_), .A1(new_new_n326_), .B0(new_new_n693_), .Y(new_new_n694_));
  AOI220     g0672(.A0(i_12_), .A1(new_new_n70_), .B0(new_new_n381_), .B1(new_new_n642_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n695_), .B(new_new_n238_), .Y(new_new_n696_));
  AOI210     g0674(.A0(new_new_n442_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n697_));
  NOi31      g0675(.An(new_new_n697_), .B(new_new_n588_), .C(new_new_n45_), .Y(new_new_n698_));
  NA2        g0676(.A(new_new_n127_), .B(i_13_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n641_), .B(new_new_n114_), .Y(new_new_n700_));
  INV        g0678(.A(new_new_n700_), .Y(new_new_n701_));
  OAI220     g0679(.A0(new_new_n701_), .A1(new_new_n69_), .B0(new_new_n699_), .B1(new_new_n682_), .Y(new_new_n702_));
  NO3        g0680(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n100_), .Y(new_new_n703_));
  NA2        g0681(.A(new_new_n26_), .B(new_new_n192_), .Y(new_new_n704_));
  NA2        g0682(.A(new_new_n704_), .B(i_7_), .Y(new_new_n705_));
  NO3        g0683(.A(new_new_n469_), .B(new_new_n233_), .C(new_new_n83_), .Y(new_new_n706_));
  AOI210     g0684(.A0(new_new_n706_), .A1(new_new_n705_), .B0(new_new_n703_), .Y(new_new_n707_));
  AOI220     g0685(.A0(new_new_n381_), .A1(new_new_n642_), .B0(new_new_n90_), .B1(new_new_n101_), .Y(new_new_n708_));
  OAI220     g0686(.A0(new_new_n708_), .A1(new_new_n594_), .B0(new_new_n707_), .B1(new_new_n605_), .Y(new_new_n709_));
  NO4        g0687(.A(new_new_n709_), .B(new_new_n702_), .C(new_new_n698_), .D(new_new_n696_), .Y(new_new_n710_));
  OR2        g0688(.A(i_11_), .B(i_6_), .Y(new_new_n711_));
  NO2        g0689(.A(new_new_n701_), .B(new_new_n711_), .Y(new_new_n712_));
  NA3        g0690(.A(new_new_n404_), .B(new_new_n597_), .C(new_new_n96_), .Y(new_new_n713_));
  NA2        g0691(.A(new_new_n633_), .B(i_13_), .Y(new_new_n714_));
  NAi21      g0692(.An(i_11_), .B(i_12_), .Y(new_new_n715_));
  NO3        g0693(.A(new_new_n469_), .B(new_new_n572_), .C(new_new_n598_), .Y(new_new_n716_));
  NA2        g0694(.A(new_new_n716_), .B(new_new_n304_), .Y(new_new_n717_));
  NA3        g0695(.A(new_new_n717_), .B(new_new_n714_), .C(new_new_n713_), .Y(new_new_n718_));
  OAI210     g0696(.A0(new_new_n718_), .A1(new_new_n712_), .B0(new_new_n63_), .Y(new_new_n719_));
  OAI210     g0697(.A0(new_new_n233_), .A1(new_new_n367_), .B0(new_new_n365_), .Y(new_new_n720_));
  NO2        g0698(.A(new_new_n128_), .B(i_2_), .Y(new_new_n721_));
  NA2        g0699(.A(new_new_n721_), .B(new_new_n626_), .Y(new_new_n722_));
  NA2        g0700(.A(new_new_n722_), .B(new_new_n720_), .Y(new_new_n723_));
  NA3        g0701(.A(new_new_n723_), .B(new_new_n46_), .C(new_new_n222_), .Y(new_new_n724_));
  NA4        g0702(.A(new_new_n724_), .B(new_new_n719_), .C(new_new_n710_), .D(new_new_n694_), .Y(new_new_n725_));
  OR4        g0703(.A(new_new_n725_), .B(new_new_n687_), .C(new_new_n671_), .D(new_new_n608_), .Y(mai5));
  AOI210     g0704(.A0(new_new_n657_), .A1(new_new_n262_), .B0(new_new_n411_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n594_), .B(i_11_), .Y(new_new_n728_));
  OAI210     g0706(.A0(new_new_n597_), .A1(new_new_n86_), .B0(new_new_n728_), .Y(new_new_n729_));
  NA2        g0707(.A(new_new_n729_), .B(new_new_n727_), .Y(new_new_n730_));
  NO3        g0708(.A(i_11_), .B(new_new_n233_), .C(i_13_), .Y(new_new_n731_));
  NO2        g0709(.A(new_new_n124_), .B(new_new_n23_), .Y(new_new_n732_));
  NA2        g0710(.A(i_12_), .B(i_8_), .Y(new_new_n733_));
  OAI210     g0711(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n733_), .Y(new_new_n734_));
  INV        g0712(.A(new_new_n441_), .Y(new_new_n735_));
  AOI220     g0713(.A0(new_new_n310_), .A1(new_new_n565_), .B0(new_new_n734_), .B1(new_new_n732_), .Y(new_new_n736_));
  INV        g0714(.A(new_new_n736_), .Y(new_new_n737_));
  NO2        g0715(.A(new_new_n737_), .B(new_new_n730_), .Y(new_new_n738_));
  INV        g0716(.A(new_new_n170_), .Y(new_new_n739_));
  INV        g0717(.A(new_new_n241_), .Y(new_new_n740_));
  OAI210     g0718(.A0(new_new_n683_), .A1(new_new_n443_), .B0(new_new_n110_), .Y(new_new_n741_));
  AOI210     g0719(.A0(new_new_n741_), .A1(new_new_n740_), .B0(new_new_n739_), .Y(new_new_n742_));
  NO2        g0720(.A(new_new_n450_), .B(new_new_n26_), .Y(new_new_n743_));
  NO2        g0721(.A(new_new_n743_), .B(new_new_n413_), .Y(new_new_n744_));
  NA2        g0722(.A(new_new_n744_), .B(i_2_), .Y(new_new_n745_));
  INV        g0723(.A(new_new_n745_), .Y(new_new_n746_));
  AOI210     g0724(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n410_), .Y(new_new_n747_));
  AOI210     g0725(.A0(new_new_n747_), .A1(new_new_n746_), .B0(new_new_n742_), .Y(new_new_n748_));
  NO2        g0726(.A(new_new_n189_), .B(new_new_n125_), .Y(new_new_n749_));
  OAI210     g0727(.A0(new_new_n749_), .A1(new_new_n732_), .B0(i_2_), .Y(new_new_n750_));
  NO2        g0728(.A(new_new_n750_), .B(new_new_n192_), .Y(new_new_n751_));
  OA210      g0729(.A0(new_new_n611_), .A1(new_new_n126_), .B0(i_13_), .Y(new_new_n752_));
  NA2        g0730(.A(new_new_n198_), .B(new_new_n201_), .Y(new_new_n753_));
  NA2        g0731(.A(new_new_n151_), .B(new_new_n589_), .Y(new_new_n754_));
  AOI210     g0732(.A0(new_new_n754_), .A1(new_new_n753_), .B0(new_new_n368_), .Y(new_new_n755_));
  AOI210     g0733(.A0(new_new_n206_), .A1(new_new_n148_), .B0(new_new_n507_), .Y(new_new_n756_));
  OAI210     g0734(.A0(new_new_n756_), .A1(new_new_n223_), .B0(new_new_n413_), .Y(new_new_n757_));
  NO2        g0735(.A(new_new_n101_), .B(new_new_n45_), .Y(new_new_n758_));
  INV        g0736(.A(new_new_n294_), .Y(new_new_n759_));
  NA4        g0737(.A(new_new_n759_), .B(new_new_n297_), .C(new_new_n124_), .D(new_new_n43_), .Y(new_new_n760_));
  OAI210     g0738(.A0(new_new_n760_), .A1(new_new_n758_), .B0(new_new_n757_), .Y(new_new_n761_));
  NO4        g0739(.A(new_new_n761_), .B(new_new_n755_), .C(new_new_n752_), .D(new_new_n751_), .Y(new_new_n762_));
  NA2        g0740(.A(new_new_n565_), .B(new_new_n28_), .Y(new_new_n763_));
  NA2        g0741(.A(new_new_n731_), .B(new_new_n268_), .Y(new_new_n764_));
  NA2        g0742(.A(new_new_n764_), .B(new_new_n763_), .Y(new_new_n765_));
  NO2        g0743(.A(new_new_n62_), .B(i_12_), .Y(new_new_n766_));
  NO2        g0744(.A(new_new_n766_), .B(new_new_n126_), .Y(new_new_n767_));
  NO2        g0745(.A(new_new_n767_), .B(new_new_n589_), .Y(new_new_n768_));
  AOI220     g0746(.A0(new_new_n768_), .A1(new_new_n36_), .B0(new_new_n765_), .B1(new_new_n47_), .Y(new_new_n769_));
  NA4        g0747(.A(new_new_n769_), .B(new_new_n762_), .C(new_new_n748_), .D(new_new_n738_), .Y(mai6));
  NO3        g0748(.A(new_new_n250_), .B(new_new_n299_), .C(i_1_), .Y(new_new_n771_));
  NO2        g0749(.A(new_new_n184_), .B(new_new_n139_), .Y(new_new_n772_));
  OAI210     g0750(.A0(new_new_n772_), .A1(new_new_n771_), .B0(new_new_n721_), .Y(new_new_n773_));
  NA4        g0751(.A(new_new_n385_), .B(new_new_n474_), .C(new_new_n69_), .D(new_new_n100_), .Y(new_new_n774_));
  INV        g0752(.A(new_new_n774_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n218_), .B(new_new_n478_), .Y(new_new_n776_));
  NO2        g0754(.A(i_11_), .B(i_9_), .Y(new_new_n777_));
  NO3        g0755(.A(new_new_n776_), .B(new_new_n775_), .C(new_new_n322_), .Y(new_new_n778_));
  AO210      g0756(.A0(new_new_n778_), .A1(new_new_n773_), .B0(i_12_), .Y(new_new_n779_));
  NA2        g0757(.A(new_new_n369_), .B(new_new_n328_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n572_), .B(new_new_n63_), .Y(new_new_n781_));
  NA2        g0759(.A(new_new_n673_), .B(new_new_n69_), .Y(new_new_n782_));
  NA4        g0760(.A(new_new_n616_), .B(new_new_n782_), .C(new_new_n781_), .D(new_new_n780_), .Y(new_new_n783_));
  INV        g0761(.A(new_new_n195_), .Y(new_new_n784_));
  AOI220     g0762(.A0(new_new_n784_), .A1(new_new_n777_), .B0(new_new_n783_), .B1(new_new_n71_), .Y(new_new_n785_));
  NO2        g0763(.A(new_new_n32_), .B(i_11_), .Y(new_new_n786_));
  NA3        g0764(.A(new_new_n786_), .B(new_new_n465_), .C(new_new_n385_), .Y(new_new_n787_));
  NAi32      g0765(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n788_));
  AOI210     g0766(.A0(new_new_n711_), .A1(new_new_n84_), .B0(new_new_n788_), .Y(new_new_n789_));
  OAI210     g0767(.A0(new_new_n672_), .A1(new_new_n553_), .B0(new_new_n552_), .Y(new_new_n790_));
  NAi31      g0768(.An(new_new_n789_), .B(new_new_n790_), .C(new_new_n787_), .Y(new_new_n791_));
  NO2        g0769(.A(new_new_n688_), .B(i_2_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n793_));
  OAI210     g0771(.A0(new_new_n793_), .A1(new_new_n403_), .B0(new_new_n355_), .Y(new_new_n794_));
  NA2        g0772(.A(new_new_n794_), .B(new_new_n792_), .Y(new_new_n795_));
  AO220      g0773(.A0(new_new_n354_), .A1(new_new_n344_), .B0(new_new_n392_), .B1(new_new_n589_), .Y(new_new_n796_));
  NA3        g0774(.A(new_new_n796_), .B(new_new_n251_), .C(i_7_), .Y(new_new_n797_));
  NA3        g0775(.A(new_new_n443_), .B(new_new_n147_), .C(new_new_n67_), .Y(new_new_n798_));
  AO210      g0776(.A0(new_new_n482_), .A1(new_new_n735_), .B0(new_new_n36_), .Y(new_new_n799_));
  NA4        g0777(.A(new_new_n799_), .B(new_new_n798_), .C(new_new_n797_), .D(new_new_n795_), .Y(new_new_n800_));
  OAI210     g0778(.A0(new_new_n632_), .A1(i_11_), .B0(new_new_n84_), .Y(new_new_n801_));
  AOI220     g0779(.A0(new_new_n801_), .A1(new_new_n552_), .B0(new_new_n776_), .B1(new_new_n705_), .Y(new_new_n802_));
  NA3        g0780(.A(new_new_n368_), .B(new_new_n234_), .C(new_new_n147_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n392_), .B(new_new_n68_), .Y(new_new_n804_));
  NA4        g0782(.A(new_new_n804_), .B(new_new_n803_), .C(new_new_n802_), .D(new_new_n596_), .Y(new_new_n805_));
  AO210      g0783(.A0(new_new_n507_), .A1(new_new_n47_), .B0(new_new_n85_), .Y(new_new_n806_));
  NA3        g0784(.A(new_new_n806_), .B(new_new_n475_), .C(new_new_n216_), .Y(new_new_n807_));
  AOI210     g0785(.A0(new_new_n443_), .A1(new_new_n441_), .B0(new_new_n551_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n601_), .B(new_new_n101_), .Y(new_new_n809_));
  OAI210     g0787(.A0(new_new_n809_), .A1(new_new_n111_), .B0(new_new_n402_), .Y(new_new_n810_));
  NA2        g0788(.A(new_new_n240_), .B(new_new_n47_), .Y(new_new_n811_));
  NA2        g0789(.A(new_new_n811_), .B(new_new_n578_), .Y(new_new_n812_));
  NA3        g0790(.A(new_new_n812_), .B(new_new_n321_), .C(i_7_), .Y(new_new_n813_));
  NA4        g0791(.A(new_new_n813_), .B(new_new_n810_), .C(new_new_n808_), .D(new_new_n807_), .Y(new_new_n814_));
  NO4        g0792(.A(new_new_n814_), .B(new_new_n805_), .C(new_new_n800_), .D(new_new_n791_), .Y(new_new_n815_));
  NA4        g0793(.A(new_new_n815_), .B(new_new_n785_), .C(new_new_n779_), .D(new_new_n375_), .Y(mai3));
  NA2        g0794(.A(i_6_), .B(i_7_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n817_), .B(i_0_), .Y(new_new_n818_));
  NO2        g0796(.A(i_11_), .B(new_new_n233_), .Y(new_new_n819_));
  OAI210     g0797(.A0(new_new_n818_), .A1(new_new_n282_), .B0(new_new_n819_), .Y(new_new_n820_));
  NO2        g0798(.A(new_new_n820_), .B(new_new_n192_), .Y(new_new_n821_));
  NO3        g0799(.A(new_new_n446_), .B(new_new_n88_), .C(new_new_n45_), .Y(new_new_n822_));
  OA210      g0800(.A0(new_new_n822_), .A1(new_new_n821_), .B0(new_new_n173_), .Y(new_new_n823_));
  INV        g0801(.A(new_new_n803_), .Y(new_new_n824_));
  NA2        g0802(.A(new_new_n824_), .B(new_new_n40_), .Y(new_new_n825_));
  NO3        g0803(.A(new_new_n621_), .B(new_new_n450_), .C(new_new_n131_), .Y(new_new_n826_));
  NA2        g0804(.A(new_new_n404_), .B(new_new_n46_), .Y(new_new_n827_));
  AN2        g0805(.A(new_new_n448_), .B(new_new_n55_), .Y(new_new_n828_));
  NO2        g0806(.A(new_new_n828_), .B(new_new_n826_), .Y(new_new_n829_));
  AOI210     g0807(.A0(new_new_n829_), .A1(new_new_n825_), .B0(new_new_n49_), .Y(new_new_n830_));
  NO4        g0808(.A(new_new_n372_), .B(new_new_n378_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n831_));
  NA2        g0809(.A(new_new_n184_), .B(new_new_n561_), .Y(new_new_n832_));
  NA2        g0810(.A(new_new_n697_), .B(new_new_n665_), .Y(new_new_n833_));
  NA2        g0811(.A(i_0_), .B(new_new_n433_), .Y(new_new_n834_));
  OAI220     g0812(.A0(new_new_n834_), .A1(new_new_n833_), .B0(new_new_n1032_), .B1(new_new_n63_), .Y(new_new_n835_));
  NOi21      g0813(.An(i_5_), .B(i_9_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n836_), .B(new_new_n440_), .Y(new_new_n837_));
  INV        g0815(.A(new_new_n677_), .Y(new_new_n838_));
  NO3        g0816(.A(new_new_n407_), .B(new_new_n259_), .C(new_new_n71_), .Y(new_new_n839_));
  NO2        g0817(.A(new_new_n174_), .B(new_new_n148_), .Y(new_new_n840_));
  AOI210     g0818(.A0(new_new_n840_), .A1(new_new_n240_), .B0(new_new_n839_), .Y(new_new_n841_));
  OAI220     g0819(.A0(new_new_n841_), .A1(new_new_n180_), .B0(new_new_n838_), .B1(new_new_n837_), .Y(new_new_n842_));
  NO4        g0820(.A(new_new_n842_), .B(new_new_n835_), .C(new_new_n830_), .D(new_new_n823_), .Y(new_new_n843_));
  NOi21      g0821(.An(i_0_), .B(i_10_), .Y(new_new_n844_));
  NA2        g0822(.A(new_new_n184_), .B(new_new_n24_), .Y(new_new_n845_));
  NO2        g0823(.A(new_new_n664_), .B(new_new_n586_), .Y(new_new_n846_));
  NO2        g0824(.A(new_new_n846_), .B(new_new_n845_), .Y(new_new_n847_));
  NA2        g0825(.A(new_new_n304_), .B(new_new_n129_), .Y(new_new_n848_));
  NAi21      g0826(.An(new_new_n161_), .B(new_new_n433_), .Y(new_new_n849_));
  OAI220     g0827(.A0(new_new_n849_), .A1(new_new_n811_), .B0(new_new_n848_), .B1(new_new_n396_), .Y(new_new_n850_));
  NO2        g0828(.A(new_new_n850_), .B(new_new_n847_), .Y(new_new_n851_));
  NO2        g0829(.A(new_new_n385_), .B(new_new_n286_), .Y(new_new_n852_));
  NA2        g0830(.A(new_new_n852_), .B(new_new_n700_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n562_), .B(i_0_), .Y(new_new_n854_));
  NO3        g0832(.A(new_new_n854_), .B(new_new_n380_), .C(new_new_n86_), .Y(new_new_n855_));
  NO4        g0833(.A(new_new_n577_), .B(new_new_n213_), .C(new_new_n410_), .D(new_new_n403_), .Y(new_new_n856_));
  AOI210     g0834(.A0(new_new_n856_), .A1(i_11_), .B0(new_new_n855_), .Y(new_new_n857_));
  AN2        g0835(.A(new_new_n95_), .B(new_new_n239_), .Y(new_new_n858_));
  NA2        g0836(.A(new_new_n731_), .B(new_new_n322_), .Y(new_new_n859_));
  AOI210     g0837(.A0(new_new_n475_), .A1(new_new_n86_), .B0(new_new_n58_), .Y(new_new_n860_));
  OAI220     g0838(.A0(new_new_n860_), .A1(new_new_n859_), .B0(new_new_n652_), .B1(new_new_n524_), .Y(new_new_n861_));
  INV        g0839(.A(new_new_n526_), .Y(new_new_n862_));
  NO4        g0840(.A(new_new_n114_), .B(new_new_n58_), .C(new_new_n661_), .D(i_5_), .Y(new_new_n863_));
  AN2        g0841(.A(new_new_n863_), .B(new_new_n862_), .Y(new_new_n864_));
  AOI210     g0842(.A0(i_0_), .A1(new_new_n97_), .B0(new_new_n184_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n556_), .B(i_4_), .Y(new_new_n866_));
  NA2        g0844(.A(new_new_n187_), .B(new_new_n201_), .Y(new_new_n867_));
  OAI220     g0845(.A0(new_new_n867_), .A1(new_new_n859_), .B0(new_new_n866_), .B1(new_new_n865_), .Y(new_new_n868_));
  NO4        g0846(.A(new_new_n868_), .B(new_new_n864_), .C(new_new_n861_), .D(new_new_n858_), .Y(new_new_n869_));
  NA4        g0847(.A(new_new_n869_), .B(new_new_n857_), .C(new_new_n853_), .D(new_new_n851_), .Y(new_new_n870_));
  NO2        g0848(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n871_));
  NA2        g0849(.A(i_11_), .B(i_9_), .Y(new_new_n872_));
  NO3        g0850(.A(i_12_), .B(new_new_n872_), .C(new_new_n595_), .Y(new_new_n873_));
  AO220      g0851(.A0(new_new_n873_), .A1(new_new_n871_), .B0(new_new_n261_), .B1(new_new_n85_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n389_), .B(new_new_n178_), .Y(new_new_n875_));
  NAi31      g0853(.An(new_new_n256_), .B(new_new_n875_), .C(new_new_n159_), .Y(new_new_n876_));
  NO2        g0854(.A(new_new_n872_), .B(new_new_n71_), .Y(new_new_n877_));
  NO2        g0855(.A(new_new_n174_), .B(i_0_), .Y(new_new_n878_));
  INV        g0856(.A(new_new_n878_), .Y(new_new_n879_));
  NA2        g0857(.A(new_new_n465_), .B(new_new_n228_), .Y(new_new_n880_));
  OAI220     g0858(.A0(i_12_), .A1(new_new_n837_), .B0(new_new_n880_), .B1(new_new_n879_), .Y(new_new_n881_));
  NO3        g0859(.A(new_new_n881_), .B(new_new_n876_), .C(new_new_n874_), .Y(new_new_n882_));
  NA2        g0860(.A(new_new_n651_), .B(new_new_n121_), .Y(new_new_n883_));
  NO2        g0861(.A(i_6_), .B(new_new_n883_), .Y(new_new_n884_));
  AOI210     g0862(.A0(new_new_n442_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n170_), .B(new_new_n102_), .Y(new_new_n886_));
  NOi32      g0864(.An(new_new_n885_), .Bn(new_new_n187_), .C(new_new_n886_), .Y(new_new_n887_));
  AOI210     g0865(.A0(new_new_n597_), .A1(new_new_n322_), .B0(new_new_n239_), .Y(new_new_n888_));
  NO2        g0866(.A(new_new_n888_), .B(new_new_n827_), .Y(new_new_n889_));
  NO3        g0867(.A(new_new_n889_), .B(new_new_n887_), .C(new_new_n884_), .Y(new_new_n890_));
  NOi21      g0868(.An(i_7_), .B(i_5_), .Y(new_new_n891_));
  NOi31      g0869(.An(new_new_n891_), .B(new_new_n844_), .C(new_new_n715_), .Y(new_new_n892_));
  NA3        g0870(.A(new_new_n892_), .B(new_new_n379_), .C(i_6_), .Y(new_new_n893_));
  OA210      g0871(.A0(new_new_n886_), .A1(new_new_n506_), .B0(new_new_n893_), .Y(new_new_n894_));
  NO3        g0872(.A(new_new_n398_), .B(new_new_n357_), .C(new_new_n353_), .Y(new_new_n895_));
  NO2        g0873(.A(new_new_n253_), .B(new_new_n311_), .Y(new_new_n896_));
  INV        g0874(.A(new_new_n715_), .Y(new_new_n897_));
  AOI210     g0875(.A0(new_new_n897_), .A1(new_new_n896_), .B0(new_new_n895_), .Y(new_new_n898_));
  NA4        g0876(.A(new_new_n898_), .B(new_new_n894_), .C(new_new_n890_), .D(new_new_n882_), .Y(new_new_n899_));
  AN2        g0877(.A(new_new_n326_), .B(new_new_n322_), .Y(new_new_n900_));
  AO220      g0878(.A0(new_new_n900_), .A1(new_new_n840_), .B0(new_new_n339_), .B1(new_new_n27_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n901_), .B(i_10_), .Y(new_new_n902_));
  OA210      g0880(.A0(new_new_n465_), .A1(new_new_n220_), .B0(new_new_n464_), .Y(new_new_n903_));
  NA3        g0881(.A(new_new_n464_), .B(new_new_n404_), .C(new_new_n46_), .Y(new_new_n904_));
  OAI210     g0882(.A0(new_new_n849_), .A1(i_6_), .B0(new_new_n904_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n877_), .B(new_new_n297_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n186_), .B(new_new_n906_), .Y(new_new_n907_));
  AOI220     g0885(.A0(new_new_n907_), .A1(new_new_n465_), .B0(new_new_n905_), .B1(new_new_n71_), .Y(new_new_n908_));
  NA3        g0886(.A(new_new_n793_), .B(new_new_n377_), .C(new_new_n632_), .Y(new_new_n909_));
  NO2        g0887(.A(new_new_n73_), .B(new_new_n733_), .Y(new_new_n910_));
  AOI210     g0888(.A0(new_new_n173_), .A1(new_new_n586_), .B0(new_new_n910_), .Y(new_new_n911_));
  AOI210     g0889(.A0(new_new_n911_), .A1(new_new_n909_), .B0(new_new_n48_), .Y(new_new_n912_));
  NO3        g0890(.A(new_new_n577_), .B(new_new_n352_), .C(new_new_n24_), .Y(new_new_n913_));
  NO2        g0891(.A(new_new_n534_), .B(new_new_n913_), .Y(new_new_n914_));
  NAi21      g0892(.An(i_9_), .B(i_5_), .Y(new_new_n915_));
  NO2        g0893(.A(new_new_n915_), .B(new_new_n398_), .Y(new_new_n916_));
  NO2        g0894(.A(new_new_n592_), .B(new_new_n104_), .Y(new_new_n917_));
  AOI220     g0895(.A0(new_new_n917_), .A1(i_0_), .B0(new_new_n916_), .B1(new_new_n611_), .Y(new_new_n918_));
  OAI220     g0896(.A0(new_new_n918_), .A1(new_new_n83_), .B0(new_new_n914_), .B1(new_new_n171_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n919_), .B(new_new_n912_), .Y(new_new_n920_));
  NA3        g0898(.A(new_new_n920_), .B(new_new_n908_), .C(new_new_n902_), .Y(new_new_n921_));
  NO3        g0899(.A(new_new_n921_), .B(new_new_n899_), .C(new_new_n870_), .Y(new_new_n922_));
  NO2        g0900(.A(new_new_n844_), .B(new_new_n715_), .Y(new_new_n923_));
  NA2        g0901(.A(new_new_n71_), .B(new_new_n45_), .Y(new_new_n924_));
  INV        g0902(.A(new_new_n924_), .Y(new_new_n925_));
  NO3        g0903(.A(new_new_n104_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n926_));
  AO220      g0904(.A0(new_new_n926_), .A1(new_new_n925_), .B0(new_new_n923_), .B1(new_new_n173_), .Y(new_new_n927_));
  AOI210     g0905(.A0(new_new_n781_), .A1(new_new_n675_), .B0(new_new_n886_), .Y(new_new_n928_));
  AOI210     g0906(.A0(new_new_n927_), .A1(new_new_n341_), .B0(new_new_n928_), .Y(new_new_n929_));
  NA3        g0907(.A(new_new_n146_), .B(new_new_n665_), .C(new_new_n71_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n790_), .B(new_new_n398_), .Y(new_new_n931_));
  NA3        g0909(.A(new_new_n818_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n819_), .B(i_9_), .Y(new_new_n933_));
  AOI210     g0911(.A0(new_new_n932_), .A1(new_new_n487_), .B0(new_new_n933_), .Y(new_new_n934_));
  OAI210     g0912(.A0(new_new_n240_), .A1(i_9_), .B0(new_new_n227_), .Y(new_new_n935_));
  AOI210     g0913(.A0(new_new_n935_), .A1(new_new_n854_), .B0(new_new_n152_), .Y(new_new_n936_));
  NO3        g0914(.A(new_new_n936_), .B(new_new_n934_), .C(new_new_n931_), .Y(new_new_n937_));
  NA3        g0915(.A(new_new_n937_), .B(new_new_n930_), .C(new_new_n929_), .Y(new_new_n938_));
  NA2        g0916(.A(new_new_n900_), .B(new_new_n368_), .Y(new_new_n939_));
  AOI210     g0917(.A0(new_new_n293_), .A1(new_new_n161_), .B0(new_new_n939_), .Y(new_new_n940_));
  NA3        g0918(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n941_));
  NA2        g0919(.A(i_5_), .B(new_new_n479_), .Y(new_new_n942_));
  AOI210     g0920(.A0(new_new_n941_), .A1(new_new_n161_), .B0(new_new_n942_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n943_), .B(new_new_n940_), .Y(new_new_n944_));
  NO3        g0922(.A(new_new_n207_), .B(new_new_n378_), .C(i_0_), .Y(new_new_n945_));
  OAI210     g0923(.A0(new_new_n945_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n946_));
  INV        g0924(.A(new_new_n216_), .Y(new_new_n947_));
  OAI220     g0925(.A0(new_new_n518_), .A1(new_new_n139_), .B0(i_12_), .B1(new_new_n605_), .Y(new_new_n948_));
  NA3        g0926(.A(new_new_n948_), .B(i_7_), .C(new_new_n947_), .Y(new_new_n949_));
  NA3        g0927(.A(new_new_n949_), .B(new_new_n946_), .C(new_new_n944_), .Y(new_new_n950_));
  NO2        g0928(.A(new_new_n238_), .B(new_new_n91_), .Y(new_new_n951_));
  AOI210     g0929(.A0(new_new_n951_), .A1(new_new_n923_), .B0(new_new_n108_), .Y(new_new_n952_));
  AOI220     g0930(.A0(new_new_n891_), .A1(new_new_n479_), .B0(new_new_n818_), .B1(new_new_n162_), .Y(new_new_n953_));
  NA2        g0931(.A(new_new_n344_), .B(new_new_n175_), .Y(new_new_n954_));
  OA220      g0932(.A0(new_new_n954_), .A1(new_new_n953_), .B0(new_new_n952_), .B1(i_5_), .Y(new_new_n955_));
  AOI210     g0933(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n174_), .Y(new_new_n956_));
  NA2        g0934(.A(new_new_n956_), .B(new_new_n903_), .Y(new_new_n957_));
  NA3        g0935(.A(new_new_n602_), .B(new_new_n184_), .C(new_new_n82_), .Y(new_new_n958_));
  NA2        g0936(.A(new_new_n958_), .B(new_new_n533_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n481_), .B(new_new_n462_), .Y(new_new_n960_));
  NO2        g0938(.A(new_new_n960_), .B(new_new_n959_), .Y(new_new_n961_));
  NA3        g0939(.A(i_5_), .B(new_new_n282_), .C(new_new_n227_), .Y(new_new_n962_));
  INV        g0940(.A(new_new_n962_), .Y(new_new_n963_));
  NA3        g0941(.A(new_new_n385_), .B(new_new_n327_), .C(new_new_n219_), .Y(new_new_n964_));
  OAI210     g0942(.A0(new_new_n832_), .A1(new_new_n639_), .B0(new_new_n964_), .Y(new_new_n965_));
  NOi31      g0943(.An(new_new_n384_), .B(new_new_n924_), .C(new_new_n235_), .Y(new_new_n966_));
  NO3        g0944(.A(new_new_n966_), .B(new_new_n965_), .C(new_new_n963_), .Y(new_new_n967_));
  NA4        g0945(.A(new_new_n967_), .B(new_new_n961_), .C(new_new_n957_), .D(new_new_n955_), .Y(new_new_n968_));
  INV        g0946(.A(new_new_n604_), .Y(new_new_n969_));
  NO3        g0947(.A(new_new_n969_), .B(new_new_n547_), .C(i_7_), .Y(new_new_n970_));
  INV        g0948(.A(new_new_n970_), .Y(new_new_n971_));
  NA3        g0949(.A(new_new_n297_), .B(i_5_), .C(new_new_n192_), .Y(new_new_n972_));
  NO4        g0950(.A(new_new_n235_), .B(new_new_n207_), .C(i_0_), .D(i_12_), .Y(new_new_n973_));
  AOI220     g0951(.A0(new_new_n973_), .A1(new_new_n297_), .B0(new_new_n775_), .B1(new_new_n175_), .Y(new_new_n974_));
  BUFFER     g0952(.A(new_new_n152_), .Y(new_new_n975_));
  NO4        g0953(.A(new_new_n975_), .B(i_12_), .C(new_new_n639_), .D(new_new_n131_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n976_), .B(new_new_n216_), .Y(new_new_n977_));
  NA3        g0955(.A(new_new_n97_), .B(new_new_n561_), .C(i_11_), .Y(new_new_n978_));
  NO2        g0956(.A(new_new_n978_), .B(new_new_n154_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n891_), .B(new_new_n461_), .Y(new_new_n980_));
  OAI210     g0958(.A0(i_7_), .A1(new_new_n972_), .B0(new_new_n980_), .Y(new_new_n981_));
  AOI210     g0959(.A0(new_new_n981_), .A1(new_new_n878_), .B0(new_new_n979_), .Y(new_new_n982_));
  NA4        g0960(.A(new_new_n982_), .B(new_new_n977_), .C(new_new_n974_), .D(new_new_n971_), .Y(new_new_n983_));
  NO4        g0961(.A(new_new_n983_), .B(new_new_n968_), .C(new_new_n950_), .D(new_new_n938_), .Y(new_new_n984_));
  OAI210     g0962(.A0(new_new_n792_), .A1(new_new_n786_), .B0(new_new_n37_), .Y(new_new_n985_));
  NA3        g0963(.A(new_new_n885_), .B(new_new_n365_), .C(i_5_), .Y(new_new_n986_));
  NA3        g0964(.A(new_new_n986_), .B(new_new_n985_), .C(new_new_n600_), .Y(new_new_n987_));
  NA2        g0965(.A(new_new_n987_), .B(new_new_n204_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n185_), .B(new_new_n187_), .Y(new_new_n989_));
  AO210      g0967(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n989_), .Y(new_new_n990_));
  OAI210     g0968(.A0(new_new_n604_), .A1(new_new_n602_), .B0(new_new_n310_), .Y(new_new_n991_));
  NAi31      g0969(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n992_));
  AOI210     g0970(.A0(new_new_n117_), .A1(new_new_n68_), .B0(new_new_n992_), .Y(new_new_n993_));
  NO2        g0971(.A(new_new_n993_), .B(new_new_n637_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n994_), .B(new_new_n991_), .C(new_new_n990_), .Y(new_new_n995_));
  NO2        g0973(.A(new_new_n453_), .B(new_new_n259_), .Y(new_new_n996_));
  NO2        g0974(.A(new_new_n996_), .B(new_new_n856_), .Y(new_new_n997_));
  OAI210     g0975(.A0(new_new_n978_), .A1(new_new_n148_), .B0(new_new_n997_), .Y(new_new_n998_));
  AOI210     g0976(.A0(new_new_n995_), .A1(new_new_n49_), .B0(new_new_n998_), .Y(new_new_n999_));
  AOI210     g0977(.A0(new_new_n999_), .A1(new_new_n988_), .B0(new_new_n71_), .Y(new_new_n1000_));
  NO2        g0978(.A(new_new_n554_), .B(new_new_n374_), .Y(new_new_n1001_));
  NO2        g0979(.A(new_new_n1001_), .B(new_new_n739_), .Y(new_new_n1002_));
  NA2        g0980(.A(i_5_), .B(new_new_n74_), .Y(new_new_n1003_));
  AOI210     g0981(.A0(new_new_n956_), .A1(i_5_), .B0(new_new_n892_), .Y(new_new_n1004_));
  AOI210     g0982(.A0(new_new_n1004_), .A1(new_new_n1003_), .B0(new_new_n666_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n253_), .B(new_new_n57_), .Y(new_new_n1006_));
  AOI220     g0984(.A0(new_new_n1006_), .A1(new_new_n74_), .B0(new_new_n339_), .B1(new_new_n250_), .Y(new_new_n1007_));
  NO2        g0985(.A(new_new_n1007_), .B(new_new_n233_), .Y(new_new_n1008_));
  NO2        g0986(.A(new_new_n1008_), .B(new_new_n1005_), .Y(new_new_n1009_));
  OAI210     g0987(.A0(new_new_n261_), .A1(new_new_n157_), .B0(new_new_n86_), .Y(new_new_n1010_));
  NA3        g0988(.A(new_new_n743_), .B(new_new_n282_), .C(new_new_n78_), .Y(new_new_n1011_));
  AOI210     g0989(.A0(new_new_n1011_), .A1(new_new_n1010_), .B0(i_11_), .Y(new_new_n1012_));
  OAI210     g0990(.A0(new_new_n1031_), .A1(new_new_n885_), .B0(new_new_n204_), .Y(new_new_n1013_));
  NA2        g0991(.A(new_new_n163_), .B(i_5_), .Y(new_new_n1014_));
  AOI210     g0992(.A0(new_new_n1013_), .A1(new_new_n753_), .B0(new_new_n1014_), .Y(new_new_n1015_));
  NO3        g0993(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1016_));
  OAI210     g0994(.A0(new_new_n896_), .A1(new_new_n299_), .B0(new_new_n1016_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n1017_), .B(new_new_n715_), .Y(new_new_n1018_));
  NO4        g0996(.A(new_new_n915_), .B(new_new_n468_), .C(new_new_n249_), .D(new_new_n248_), .Y(new_new_n1019_));
  NO2        g0997(.A(new_new_n1019_), .B(new_new_n551_), .Y(new_new_n1020_));
  NO2        g0998(.A(new_new_n789_), .B(new_new_n358_), .Y(new_new_n1021_));
  AOI210     g0999(.A0(new_new_n1021_), .A1(new_new_n1020_), .B0(new_new_n41_), .Y(new_new_n1022_));
  NO4        g1000(.A(new_new_n1022_), .B(new_new_n1018_), .C(new_new_n1015_), .D(new_new_n1012_), .Y(new_new_n1023_));
  OAI210     g1001(.A0(new_new_n1009_), .A1(i_4_), .B0(new_new_n1023_), .Y(new_new_n1024_));
  NO3        g1002(.A(new_new_n1024_), .B(new_new_n1002_), .C(new_new_n1000_), .Y(new_new_n1025_));
  NA4        g1003(.A(new_new_n1025_), .B(new_new_n984_), .C(new_new_n922_), .D(new_new_n843_), .Y(mai4));
  INV        g1004(.A(i_2_), .Y(new_new_n1029_));
  INV        g1005(.A(i_5_), .Y(new_new_n1030_));
  INV        g1006(.A(i_12_), .Y(new_new_n1031_));
  INV        g1007(.A(new_new_n831_), .Y(new_new_n1032_));
endmodule


