library verilog;
use verilog.vl_types.all;
entity divisordefreq2_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        R               : in     vl_logic;
        S               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end divisordefreq2_vlg_sample_tst;
