//Benchmark atmr_9sym_175_0.0625

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n137_, ori_ori_n138_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n164_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  INV        o002(.A(i_5_), .Y(ori_ori_n13_));
  NOi21      o003(.An(i_3_), .B(i_7_), .Y(ori_ori_n14_));
  NA3        o004(.A(ori_ori_n14_), .B(i_0_), .C(ori_ori_n13_), .Y(ori_ori_n15_));
  INV        o005(.A(i_0_), .Y(ori_ori_n16_));
  NOi21      o006(.An(i_1_), .B(i_3_), .Y(ori_ori_n17_));
  NA3        o007(.A(ori_ori_n17_), .B(ori_ori_n16_), .C(i_2_), .Y(ori_ori_n18_));
  AOI210     o008(.A0(ori_ori_n18_), .A1(ori_ori_n15_), .B0(i_6_), .Y(ori_ori_n19_));
  INV        o009(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o010(.A(i_0_), .B(ori_ori_n20_), .Y(ori_ori_n21_));
  INV        o011(.A(i_7_), .Y(ori_ori_n22_));
  NA3        o012(.A(i_6_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n23_));
  NOi21      o013(.An(i_8_), .B(i_6_), .Y(ori_ori_n24_));
  NOi21      o014(.An(i_1_), .B(i_8_), .Y(ori_ori_n25_));
  NO2        o015(.A(ori_ori_n23_), .B(ori_ori_n21_), .Y(ori_ori_n26_));
  AOI210     o016(.A0(ori_ori_n26_), .A1(ori_ori_n11_), .B0(ori_ori_n19_), .Y(ori_ori_n27_));
  NA2        o017(.A(ori_ori_n16_), .B(i_5_), .Y(ori_ori_n28_));
  INV        o018(.A(i_2_), .Y(ori_ori_n29_));
  INV        o019(.A(i_2_), .Y(ori_ori_n30_));
  NOi21      o020(.An(i_5_), .B(i_0_), .Y(ori_ori_n31_));
  NOi21      o021(.An(i_6_), .B(i_8_), .Y(ori_ori_n32_));
  NOi21      o022(.An(i_5_), .B(i_6_), .Y(ori_ori_n33_));
  NOi21      o023(.An(i_0_), .B(i_4_), .Y(ori_ori_n34_));
  INV        o024(.A(i_1_), .Y(ori_ori_n35_));
  NOi21      o025(.An(i_3_), .B(i_0_), .Y(ori_ori_n36_));
  NA2        o026(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n37_));
  NO2        o027(.A(ori_ori_n23_), .B(ori_ori_n37_), .Y(ori_ori_n38_));
  INV        o028(.A(ori_ori_n38_), .Y(ori_ori_n39_));
  NOi21      o029(.An(i_4_), .B(i_0_), .Y(ori_ori_n40_));
  NO2        o030(.A(ori_ori_n24_), .B(ori_ori_n14_), .Y(ori_ori_n41_));
  NA2        o031(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n42_));
  NOi21      o032(.An(i_2_), .B(i_8_), .Y(ori_ori_n43_));
  NO3        o033(.A(ori_ori_n138_), .B(ori_ori_n42_), .C(ori_ori_n41_), .Y(ori_ori_n44_));
  INV        o034(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o035(.A(i_1_), .B(i_3_), .Y(ori_ori_n46_));
  NA2        o036(.A(ori_ori_n46_), .B(i_0_), .Y(ori_ori_n47_));
  NOi21      o037(.An(i_4_), .B(i_3_), .Y(ori_ori_n48_));
  NOi21      o038(.An(i_1_), .B(i_4_), .Y(ori_ori_n49_));
  NA2        o039(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n50_));
  NA2        o040(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n51_));
  BUFFER     o041(.A(i_8_), .Y(ori_ori_n52_));
  NOi21      o042(.An(i_8_), .B(i_7_), .Y(ori_ori_n53_));
  NA2        o043(.A(ori_ori_n51_), .B(ori_ori_n33_), .Y(ori_ori_n54_));
  NA4        o044(.A(ori_ori_n54_), .B(ori_ori_n45_), .C(ori_ori_n39_), .D(ori_ori_n27_), .Y(ori_ori_n55_));
  NA2        o045(.A(i_8_), .B(i_7_), .Y(ori_ori_n56_));
  NO2        o046(.A(ori_ori_n56_), .B(i_6_), .Y(ori_ori_n57_));
  NA2        o047(.A(i_8_), .B(ori_ori_n22_), .Y(ori_ori_n58_));
  NOi21      o048(.An(i_1_), .B(i_2_), .Y(ori_ori_n59_));
  NO2        o049(.A(ori_ori_n137_), .B(ori_ori_n58_), .Y(ori_ori_n60_));
  OAI210     o050(.A0(ori_ori_n60_), .A1(ori_ori_n57_), .B0(ori_ori_n13_), .Y(ori_ori_n61_));
  NA3        o051(.A(ori_ori_n53_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n62_));
  NA3        o052(.A(ori_ori_n25_), .B(i_0_), .C(ori_ori_n13_), .Y(ori_ori_n63_));
  NA2        o053(.A(ori_ori_n63_), .B(ori_ori_n62_), .Y(ori_ori_n64_));
  NA2        o054(.A(ori_ori_n17_), .B(i_6_), .Y(ori_ori_n65_));
  INV        o055(.A(ori_ori_n65_), .Y(ori_ori_n66_));
  INV        o056(.A(i_0_), .Y(ori_ori_n67_));
  AOI220     o057(.A0(ori_ori_n67_), .A1(ori_ori_n66_), .B0(ori_ori_n64_), .B1(ori_ori_n48_), .Y(ori_ori_n68_));
  NA2        o058(.A(ori_ori_n68_), .B(ori_ori_n61_), .Y(ori_ori_n69_));
  NAi21      o059(.An(i_3_), .B(i_6_), .Y(ori_ori_n70_));
  NA2        o060(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n71_));
  NOi21      o061(.An(i_7_), .B(i_8_), .Y(ori_ori_n72_));
  NOi21      o062(.An(i_6_), .B(i_5_), .Y(ori_ori_n73_));
  AOI210     o063(.A0(ori_ori_n72_), .A1(ori_ori_n12_), .B0(ori_ori_n73_), .Y(ori_ori_n74_));
  NA2        o064(.A(ori_ori_n74_), .B(ori_ori_n71_), .Y(ori_ori_n75_));
  NA2        o065(.A(ori_ori_n75_), .B(ori_ori_n59_), .Y(ori_ori_n76_));
  AOI220     o066(.A0(ori_ori_n36_), .A1(ori_ori_n35_), .B0(ori_ori_n17_), .B1(ori_ori_n30_), .Y(ori_ori_n77_));
  NA3        o067(.A(ori_ori_n20_), .B(i_5_), .C(i_7_), .Y(ori_ori_n78_));
  NO2        o068(.A(ori_ori_n78_), .B(ori_ori_n77_), .Y(ori_ori_n79_));
  INV        o069(.A(ori_ori_n79_), .Y(ori_ori_n80_));
  NA2        o070(.A(ori_ori_n53_), .B(ori_ori_n30_), .Y(ori_ori_n81_));
  NA2        o071(.A(ori_ori_n35_), .B(i_6_), .Y(ori_ori_n82_));
  NOi21      o072(.An(i_2_), .B(i_1_), .Y(ori_ori_n83_));
  NAi21      o073(.An(i_6_), .B(i_0_), .Y(ori_ori_n84_));
  NA2        o074(.A(ori_ori_n49_), .B(i_5_), .Y(ori_ori_n85_));
  NOi21      o075(.An(i_4_), .B(i_6_), .Y(ori_ori_n86_));
  NO2        o076(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n87_));
  INV        o077(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  NA2        o078(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n89_));
  NOi21      o079(.An(ori_ori_n40_), .B(ori_ori_n89_), .Y(ori_ori_n90_));
  NA2        o080(.A(ori_ori_n53_), .B(ori_ori_n12_), .Y(ori_ori_n91_));
  INV        o081(.A(ori_ori_n32_), .Y(ori_ori_n92_));
  NOi21      o082(.An(i_3_), .B(i_1_), .Y(ori_ori_n93_));
  NA2        o083(.A(ori_ori_n93_), .B(i_4_), .Y(ori_ori_n94_));
  AOI210     o084(.A0(ori_ori_n92_), .A1(ori_ori_n91_), .B0(ori_ori_n94_), .Y(ori_ori_n95_));
  NOi31      o085(.An(ori_ori_n36_), .B(i_5_), .C(ori_ori_n30_), .Y(ori_ori_n96_));
  NO3        o086(.A(ori_ori_n96_), .B(ori_ori_n95_), .C(ori_ori_n90_), .Y(ori_ori_n97_));
  NA4        o087(.A(ori_ori_n97_), .B(ori_ori_n88_), .C(ori_ori_n80_), .D(ori_ori_n76_), .Y(ori_ori_n98_));
  NA2        o088(.A(ori_ori_n32_), .B(ori_ori_n34_), .Y(ori_ori_n99_));
  INV        o089(.A(ori_ori_n48_), .Y(ori_ori_n100_));
  AOI210     o090(.A0(ori_ori_n100_), .A1(ori_ori_n62_), .B0(ori_ori_n28_), .Y(ori_ori_n101_));
  NA2        o091(.A(ori_ori_n72_), .B(ori_ori_n83_), .Y(ori_ori_n102_));
  NA3        o092(.A(ori_ori_n53_), .B(ori_ori_n46_), .C(i_6_), .Y(ori_ori_n103_));
  NA2        o093(.A(ori_ori_n103_), .B(ori_ori_n102_), .Y(ori_ori_n104_));
  NOi21      o094(.An(i_0_), .B(i_2_), .Y(ori_ori_n105_));
  NA3        o095(.A(ori_ori_n105_), .B(i_7_), .C(ori_ori_n86_), .Y(ori_ori_n106_));
  NA3        o096(.A(ori_ori_n105_), .B(ori_ori_n48_), .C(ori_ori_n32_), .Y(ori_ori_n107_));
  NA2        o097(.A(ori_ori_n107_), .B(ori_ori_n106_), .Y(ori_ori_n108_));
  NA4        o098(.A(ori_ori_n46_), .B(i_6_), .C(ori_ori_n13_), .D(i_7_), .Y(ori_ori_n109_));
  NA3        o099(.A(ori_ori_n49_), .B(ori_ori_n36_), .C(i_5_), .Y(ori_ori_n110_));
  NA2        o100(.A(ori_ori_n110_), .B(ori_ori_n109_), .Y(ori_ori_n111_));
  NO4        o101(.A(ori_ori_n111_), .B(ori_ori_n108_), .C(ori_ori_n104_), .D(ori_ori_n101_), .Y(ori_ori_n112_));
  AOI210     o102(.A0(ori_ori_n52_), .A1(ori_ori_n29_), .B0(ori_ori_n72_), .Y(ori_ori_n113_));
  NO2        o103(.A(ori_ori_n113_), .B(ori_ori_n82_), .Y(ori_ori_n114_));
  NO3        o104(.A(i_2_), .B(ori_ori_n20_), .C(ori_ori_n13_), .Y(ori_ori_n115_));
  NA2        o105(.A(i_2_), .B(i_4_), .Y(ori_ori_n116_));
  AOI210     o106(.A0(ori_ori_n84_), .A1(ori_ori_n70_), .B0(ori_ori_n116_), .Y(ori_ori_n117_));
  NO2        o107(.A(i_8_), .B(i_7_), .Y(ori_ori_n118_));
  OA210      o108(.A0(ori_ori_n117_), .A1(ori_ori_n115_), .B0(ori_ori_n118_), .Y(ori_ori_n119_));
  NA2        o109(.A(ori_ori_n93_), .B(i_0_), .Y(ori_ori_n120_));
  NO2        o110(.A(ori_ori_n120_), .B(i_4_), .Y(ori_ori_n121_));
  NO3        o111(.A(ori_ori_n121_), .B(ori_ori_n119_), .C(ori_ori_n114_), .Y(ori_ori_n122_));
  NA2        o112(.A(ori_ori_n72_), .B(ori_ori_n12_), .Y(ori_ori_n123_));
  NA2        o113(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n124_));
  NA2        o114(.A(ori_ori_n40_), .B(i_3_), .Y(ori_ori_n125_));
  AOI210     o115(.A0(ori_ori_n125_), .A1(ori_ori_n124_), .B0(ori_ori_n123_), .Y(ori_ori_n126_));
  NA2        o116(.A(ori_ori_n105_), .B(ori_ori_n53_), .Y(ori_ori_n127_));
  OAI210     o117(.A0(ori_ori_n81_), .A1(ori_ori_n28_), .B0(ori_ori_n127_), .Y(ori_ori_n128_));
  NA4        o118(.A(i_5_), .B(ori_ori_n52_), .C(ori_ori_n35_), .D(ori_ori_n20_), .Y(ori_ori_n129_));
  NA3        o119(.A(ori_ori_n43_), .B(ori_ori_n31_), .C(ori_ori_n14_), .Y(ori_ori_n130_));
  NA2        o120(.A(ori_ori_n130_), .B(ori_ori_n129_), .Y(ori_ori_n131_));
  NO3        o121(.A(ori_ori_n131_), .B(ori_ori_n128_), .C(ori_ori_n126_), .Y(ori_ori_n132_));
  NA4        o122(.A(ori_ori_n132_), .B(ori_ori_n122_), .C(ori_ori_n112_), .D(ori_ori_n99_), .Y(ori_ori_n133_));
  OR4        o123(.A(ori_ori_n133_), .B(ori_ori_n98_), .C(ori_ori_n69_), .D(ori_ori_n55_), .Y(ori00));
  INV        o124(.A(i_0_), .Y(ori_ori_n137_));
  INV        o125(.A(i_4_), .Y(ori_ori_n138_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NA3        m013(.A(i_6_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_8_), .B(i_6_), .Y(mai_mai_n25_));
  AOI210     m015(.A0(mai_mai_n25_), .A1(i_5_), .B0(i_2_), .Y(mai_mai_n26_));
  AOI210     m016(.A0(mai_mai_n26_), .A1(mai_mai_n24_), .B0(mai_mai_n22_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n27_), .A1(mai_mai_n11_), .B0(mai_mai_n20_), .Y(mai_mai_n28_));
  NA2        m018(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n29_));
  NA2        m019(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n30_));
  NO2        m020(.A(i_2_), .B(i_4_), .Y(mai_mai_n31_));
  NA3        m021(.A(mai_mai_n31_), .B(i_6_), .C(i_8_), .Y(mai_mai_n32_));
  AOI210     m022(.A0(mai_mai_n30_), .A1(mai_mai_n29_), .B0(mai_mai_n32_), .Y(mai_mai_n33_));
  INV        m023(.A(i_2_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_5_), .B(i_0_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_6_), .B(i_8_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_7_), .B(i_1_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_5_), .B(i_6_), .Y(mai_mai_n38_));
  AOI220     m028(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n36_), .B1(mai_mai_n35_), .Y(mai_mai_n39_));
  NO3        m029(.A(mai_mai_n39_), .B(mai_mai_n34_), .C(i_4_), .Y(mai_mai_n40_));
  NOi21      m030(.An(i_0_), .B(i_4_), .Y(mai_mai_n41_));
  XO2        m031(.A(i_1_), .B(i_3_), .Y(mai_mai_n42_));
  NOi21      m032(.An(i_7_), .B(i_5_), .Y(mai_mai_n43_));
  AN3        m033(.A(mai_mai_n43_), .B(mai_mai_n42_), .C(mai_mai_n41_), .Y(mai_mai_n44_));
  INV        m034(.A(i_1_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_3_), .B(i_0_), .Y(mai_mai_n46_));
  NA2        m036(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m037(.A(mai_mai_n24_), .B(mai_mai_n47_), .Y(mai_mai_n48_));
  NO4        m038(.A(mai_mai_n48_), .B(mai_mai_n44_), .C(mai_mai_n40_), .D(mai_mai_n33_), .Y(mai_mai_n49_));
  NOi21      m039(.An(i_4_), .B(i_0_), .Y(mai_mai_n50_));
  AOI210     m040(.A0(mai_mai_n50_), .A1(mai_mai_n25_), .B0(mai_mai_n15_), .Y(mai_mai_n51_));
  NA2        m041(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_2_), .B(i_8_), .Y(mai_mai_n53_));
  NO3        m043(.A(mai_mai_n53_), .B(mai_mai_n50_), .C(mai_mai_n41_), .Y(mai_mai_n54_));
  NO3        m044(.A(mai_mai_n54_), .B(mai_mai_n52_), .C(mai_mai_n51_), .Y(mai_mai_n55_));
  INV        m045(.A(mai_mai_n55_), .Y(mai_mai_n56_));
  NOi31      m046(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n57_));
  NOi21      m047(.An(i_4_), .B(i_3_), .Y(mai_mai_n58_));
  NOi21      m048(.An(i_1_), .B(i_4_), .Y(mai_mai_n59_));
  AN2        m049(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  NA2        m050(.A(mai_mai_n60_), .B(mai_mai_n12_), .Y(mai_mai_n61_));
  NOi21      m051(.An(i_8_), .B(i_7_), .Y(mai_mai_n62_));
  NA3        m052(.A(mai_mai_n62_), .B(mai_mai_n58_), .C(i_6_), .Y(mai_mai_n63_));
  OAI210     m053(.A0(mai_mai_n61_), .A1(mai_mai_n52_), .B0(mai_mai_n63_), .Y(mai_mai_n64_));
  AOI220     m054(.A0(mai_mai_n64_), .A1(mai_mai_n34_), .B0(mai_mai_n53_), .B1(mai_mai_n38_), .Y(mai_mai_n65_));
  NA4        m055(.A(mai_mai_n65_), .B(mai_mai_n56_), .C(mai_mai_n49_), .D(mai_mai_n28_), .Y(mai_mai_n66_));
  NA2        m056(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n67_));
  AOI220     m057(.A0(mai_mai_n46_), .A1(i_1_), .B0(mai_mai_n42_), .B1(i_2_), .Y(mai_mai_n68_));
  NOi21      m058(.An(i_1_), .B(i_2_), .Y(mai_mai_n69_));
  NO2        m059(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n70_));
  NA2        m060(.A(mai_mai_n70_), .B(mai_mai_n14_), .Y(mai_mai_n71_));
  NA3        m061(.A(mai_mai_n62_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n72_));
  NA2        m062(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n73_));
  NA2        m063(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  NOi32      m064(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n75_));
  NA2        m065(.A(mai_mai_n75_), .B(i_3_), .Y(mai_mai_n76_));
  NA3        m066(.A(mai_mai_n18_), .B(i_2_), .C(i_6_), .Y(mai_mai_n77_));
  NA2        m067(.A(mai_mai_n77_), .B(mai_mai_n76_), .Y(mai_mai_n78_));
  NO2        m068(.A(i_0_), .B(i_4_), .Y(mai_mai_n79_));
  AOI220     m069(.A0(mai_mai_n79_), .A1(mai_mai_n78_), .B0(mai_mai_n74_), .B1(mai_mai_n58_), .Y(mai_mai_n80_));
  NA2        m070(.A(mai_mai_n80_), .B(mai_mai_n71_), .Y(mai_mai_n81_));
  NOi21      m071(.An(i_7_), .B(i_8_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n35_), .B(mai_mai_n69_), .Y(mai_mai_n83_));
  AOI220     m073(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n18_), .B1(mai_mai_n34_), .Y(mai_mai_n84_));
  NA3        m074(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n85_));
  NO2        m075(.A(mai_mai_n85_), .B(mai_mai_n84_), .Y(mai_mai_n86_));
  INV        m076(.A(mai_mai_n86_), .Y(mai_mai_n87_));
  NA3        m077(.A(mai_mai_n62_), .B(mai_mai_n34_), .C(i_3_), .Y(mai_mai_n88_));
  NA2        m078(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n89_));
  AOI210     m079(.A0(mai_mai_n89_), .A1(mai_mai_n22_), .B0(mai_mai_n88_), .Y(mai_mai_n90_));
  NOi21      m080(.An(i_2_), .B(i_1_), .Y(mai_mai_n91_));
  AN3        m081(.A(mai_mai_n82_), .B(mai_mai_n91_), .C(mai_mai_n50_), .Y(mai_mai_n92_));
  NAi21      m082(.An(i_6_), .B(i_0_), .Y(mai_mai_n93_));
  NA3        m083(.A(mai_mai_n59_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n94_));
  NOi21      m084(.An(i_4_), .B(i_6_), .Y(mai_mai_n95_));
  NOi21      m085(.An(i_5_), .B(i_3_), .Y(mai_mai_n96_));
  NA3        m086(.A(mai_mai_n96_), .B(mai_mai_n69_), .C(mai_mai_n95_), .Y(mai_mai_n97_));
  OAI210     m087(.A0(mai_mai_n94_), .A1(mai_mai_n93_), .B0(mai_mai_n97_), .Y(mai_mai_n98_));
  NA2        m088(.A(mai_mai_n69_), .B(mai_mai_n36_), .Y(mai_mai_n99_));
  NO3        m089(.A(mai_mai_n98_), .B(mai_mai_n92_), .C(mai_mai_n90_), .Y(mai_mai_n100_));
  NOi31      m090(.An(mai_mai_n50_), .B(mai_mai_n147_), .C(i_2_), .Y(mai_mai_n101_));
  NA2        m091(.A(mai_mai_n36_), .B(mai_mai_n14_), .Y(mai_mai_n102_));
  NOi21      m092(.An(i_3_), .B(i_1_), .Y(mai_mai_n103_));
  NO2        m093(.A(mai_mai_n102_), .B(mai_mai_n148_), .Y(mai_mai_n104_));
  NO2        m094(.A(mai_mai_n104_), .B(mai_mai_n101_), .Y(mai_mai_n105_));
  NA4        m095(.A(mai_mai_n105_), .B(mai_mai_n100_), .C(mai_mai_n87_), .D(mai_mai_n83_), .Y(mai_mai_n106_));
  NA2        m096(.A(mai_mai_n53_), .B(mai_mai_n15_), .Y(mai_mai_n107_));
  NOi31      m097(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n108_));
  NOi31      m098(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n109_));
  OAI210     m099(.A0(mai_mai_n109_), .A1(mai_mai_n108_), .B0(i_7_), .Y(mai_mai_n110_));
  NA3        m100(.A(mai_mai_n110_), .B(mai_mai_n107_), .C(mai_mai_n99_), .Y(mai_mai_n111_));
  NA2        m101(.A(mai_mai_n111_), .B(mai_mai_n41_), .Y(mai_mai_n112_));
  NA2        m102(.A(mai_mai_n58_), .B(mai_mai_n37_), .Y(mai_mai_n113_));
  AOI210     m103(.A0(mai_mai_n113_), .A1(mai_mai_n72_), .B0(mai_mai_n30_), .Y(mai_mai_n114_));
  NA4        m104(.A(mai_mai_n60_), .B(mai_mai_n91_), .C(mai_mai_n17_), .D(mai_mai_n12_), .Y(mai_mai_n115_));
  NA3        m105(.A(mai_mai_n62_), .B(mai_mai_n57_), .C(i_6_), .Y(mai_mai_n116_));
  NA2        m106(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NA3        m107(.A(i_0_), .B(mai_mai_n37_), .C(mai_mai_n95_), .Y(mai_mai_n118_));
  NA3        m108(.A(mai_mai_n50_), .B(mai_mai_n43_), .C(mai_mai_n18_), .Y(mai_mai_n119_));
  NA2        m109(.A(mai_mai_n58_), .B(mai_mai_n36_), .Y(mai_mai_n120_));
  NA3        m110(.A(mai_mai_n120_), .B(mai_mai_n119_), .C(mai_mai_n118_), .Y(mai_mai_n121_));
  NA4        m111(.A(mai_mai_n57_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n122_));
  NA4        m112(.A(mai_mai_n59_), .B(mai_mai_n38_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n123_));
  NA4        m113(.A(mai_mai_n59_), .B(mai_mai_n46_), .C(i_5_), .D(mai_mai_n23_), .Y(mai_mai_n124_));
  NA3        m114(.A(mai_mai_n124_), .B(mai_mai_n123_), .C(mai_mai_n122_), .Y(mai_mai_n125_));
  NO4        m115(.A(mai_mai_n125_), .B(mai_mai_n121_), .C(mai_mai_n117_), .D(mai_mai_n114_), .Y(mai_mai_n126_));
  NOi21      m116(.An(i_5_), .B(i_2_), .Y(mai_mai_n127_));
  AOI220     m117(.A0(mai_mai_n127_), .A1(mai_mai_n82_), .B0(mai_mai_n60_), .B1(mai_mai_n31_), .Y(mai_mai_n128_));
  AOI210     m118(.A0(mai_mai_n128_), .A1(mai_mai_n107_), .B0(mai_mai_n89_), .Y(mai_mai_n129_));
  NO4        m119(.A(i_2_), .B(mai_mai_n21_), .C(mai_mai_n11_), .D(mai_mai_n14_), .Y(mai_mai_n130_));
  NO2        m120(.A(i_8_), .B(i_7_), .Y(mai_mai_n131_));
  AN2        m121(.A(mai_mai_n130_), .B(mai_mai_n131_), .Y(mai_mai_n132_));
  NA4        m122(.A(mai_mai_n103_), .B(i_0_), .C(i_5_), .D(mai_mai_n23_), .Y(mai_mai_n133_));
  NO2        m123(.A(mai_mai_n133_), .B(i_4_), .Y(mai_mai_n134_));
  NO3        m124(.A(mai_mai_n134_), .B(mai_mai_n132_), .C(mai_mai_n129_), .Y(mai_mai_n135_));
  NA2        m125(.A(mai_mai_n82_), .B(mai_mai_n12_), .Y(mai_mai_n136_));
  NO2        m126(.A(mai_mai_n149_), .B(mai_mai_n136_), .Y(mai_mai_n137_));
  NA3        m127(.A(i_0_), .B(mai_mai_n62_), .C(mai_mai_n95_), .Y(mai_mai_n138_));
  OAI210     m128(.A0(mai_mai_n88_), .A1(mai_mai_n30_), .B0(mai_mai_n138_), .Y(mai_mai_n139_));
  NA4        m129(.A(mai_mai_n96_), .B(mai_mai_n60_), .C(mai_mai_n45_), .D(mai_mai_n21_), .Y(mai_mai_n140_));
  INV        m130(.A(mai_mai_n140_), .Y(mai_mai_n141_));
  NO3        m131(.A(mai_mai_n141_), .B(mai_mai_n139_), .C(mai_mai_n137_), .Y(mai_mai_n142_));
  NA4        m132(.A(mai_mai_n142_), .B(mai_mai_n135_), .C(mai_mai_n126_), .D(mai_mai_n112_), .Y(mai_mai_n143_));
  OR4        m133(.A(mai_mai_n143_), .B(mai_mai_n106_), .C(mai_mai_n81_), .D(mai_mai_n66_), .Y(mai00));
  INV        m134(.A(i_8_), .Y(mai_mai_n147_));
  INV        m135(.A(i_3_), .Y(mai_mai_n148_));
  INV        m136(.A(i_3_), .Y(mai_mai_n149_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NO2        u008(.A(men_men_n16_), .B(men_men_n13_), .Y(men_men_n19_));
  INV        u009(.A(i_4_), .Y(men_men_n20_));
  NA2        u010(.A(i_0_), .B(men_men_n20_), .Y(men_men_n21_));
  INV        u011(.A(i_7_), .Y(men_men_n22_));
  NA3        u012(.A(i_6_), .B(i_5_), .C(men_men_n22_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  NOi21      u014(.An(i_1_), .B(i_8_), .Y(men_men_n25_));
  AOI220     u015(.A0(men_men_n25_), .A1(i_2_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n26_));
  AOI210     u016(.A0(men_men_n26_), .A1(men_men_n23_), .B0(men_men_n21_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n11_), .B0(men_men_n19_), .Y(men_men_n28_));
  NA2        u018(.A(men_men_n17_), .B(i_5_), .Y(men_men_n29_));
  INV        u019(.A(i_2_), .Y(men_men_n30_));
  NOi21      u020(.An(i_5_), .B(i_0_), .Y(men_men_n31_));
  NOi21      u021(.An(i_6_), .B(i_8_), .Y(men_men_n32_));
  NOi21      u022(.An(i_7_), .B(i_1_), .Y(men_men_n33_));
  NOi21      u023(.An(i_5_), .B(i_6_), .Y(men_men_n34_));
  AOI220     u024(.A0(men_men_n34_), .A1(men_men_n33_), .B0(men_men_n32_), .B1(men_men_n31_), .Y(men_men_n35_));
  NO3        u025(.A(men_men_n35_), .B(men_men_n30_), .C(i_4_), .Y(men_men_n36_));
  NOi21      u026(.An(i_0_), .B(i_4_), .Y(men_men_n37_));
  XO2        u027(.A(i_1_), .B(i_3_), .Y(men_men_n38_));
  NOi21      u028(.An(i_7_), .B(i_5_), .Y(men_men_n39_));
  AN3        u029(.A(men_men_n39_), .B(men_men_n38_), .C(men_men_n37_), .Y(men_men_n40_));
  INV        u030(.A(i_1_), .Y(men_men_n41_));
  NOi21      u031(.An(i_3_), .B(i_0_), .Y(men_men_n42_));
  NA2        u032(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA3        u033(.A(i_6_), .B(men_men_n14_), .C(i_7_), .Y(men_men_n44_));
  AOI210     u034(.A0(men_men_n44_), .A1(men_men_n23_), .B0(men_men_n43_), .Y(men_men_n45_));
  NO3        u035(.A(men_men_n45_), .B(men_men_n40_), .C(men_men_n36_), .Y(men_men_n46_));
  INV        u036(.A(i_8_), .Y(men_men_n47_));
  NA2        u037(.A(i_1_), .B(men_men_n11_), .Y(men_men_n48_));
  NO4        u038(.A(men_men_n48_), .B(men_men_n164_), .C(i_2_), .D(men_men_n47_), .Y(men_men_n49_));
  NOi21      u039(.An(i_4_), .B(i_0_), .Y(men_men_n50_));
  AOI210     u040(.A0(men_men_n50_), .A1(men_men_n24_), .B0(men_men_n15_), .Y(men_men_n51_));
  NA2        u041(.A(i_1_), .B(men_men_n14_), .Y(men_men_n52_));
  NOi21      u042(.An(i_2_), .B(i_8_), .Y(men_men_n53_));
  NO3        u043(.A(men_men_n53_), .B(men_men_n50_), .C(men_men_n37_), .Y(men_men_n54_));
  NO3        u044(.A(men_men_n54_), .B(men_men_n52_), .C(men_men_n51_), .Y(men_men_n55_));
  NO2        u045(.A(men_men_n55_), .B(men_men_n49_), .Y(men_men_n56_));
  NOi31      u046(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n57_));
  NA2        u047(.A(men_men_n57_), .B(i_0_), .Y(men_men_n58_));
  NOi21      u048(.An(i_4_), .B(i_3_), .Y(men_men_n59_));
  NOi21      u049(.An(i_1_), .B(i_4_), .Y(men_men_n60_));
  OAI210     u050(.A0(men_men_n60_), .A1(men_men_n59_), .B0(men_men_n53_), .Y(men_men_n61_));
  NA2        u051(.A(men_men_n61_), .B(men_men_n58_), .Y(men_men_n62_));
  NOi21      u052(.An(i_8_), .B(i_7_), .Y(men_men_n63_));
  NA3        u053(.A(men_men_n63_), .B(men_men_n59_), .C(i_6_), .Y(men_men_n64_));
  INV        u054(.A(men_men_n64_), .Y(men_men_n65_));
  AOI220     u055(.A0(men_men_n65_), .A1(men_men_n30_), .B0(men_men_n62_), .B1(men_men_n34_), .Y(men_men_n66_));
  NA4        u056(.A(men_men_n66_), .B(men_men_n56_), .C(men_men_n46_), .D(men_men_n28_), .Y(men_men_n67_));
  NA2        u057(.A(i_8_), .B(i_7_), .Y(men_men_n68_));
  NO3        u058(.A(men_men_n68_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n69_));
  NA2        u059(.A(i_8_), .B(men_men_n22_), .Y(men_men_n70_));
  AOI220     u060(.A0(men_men_n42_), .A1(i_1_), .B0(men_men_n38_), .B1(i_2_), .Y(men_men_n71_));
  NOi21      u061(.An(i_1_), .B(i_2_), .Y(men_men_n72_));
  NA3        u062(.A(men_men_n72_), .B(men_men_n50_), .C(i_6_), .Y(men_men_n73_));
  OAI210     u063(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n73_), .Y(men_men_n74_));
  OAI210     u064(.A0(men_men_n74_), .A1(men_men_n69_), .B0(men_men_n14_), .Y(men_men_n75_));
  NA3        u065(.A(men_men_n63_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n76_));
  NA3        u066(.A(men_men_n25_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n77_));
  NA2        u067(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NOi32      u068(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n79_));
  NA2        u069(.A(men_men_n79_), .B(i_3_), .Y(men_men_n80_));
  NA3        u070(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n81_));
  NA2        u071(.A(men_men_n81_), .B(men_men_n80_), .Y(men_men_n82_));
  NO2        u072(.A(i_0_), .B(i_4_), .Y(men_men_n83_));
  AOI220     u073(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n78_), .B1(men_men_n59_), .Y(men_men_n84_));
  NA2        u074(.A(men_men_n84_), .B(men_men_n75_), .Y(men_men_n85_));
  NO3        u075(.A(i_3_), .B(i_0_), .C(men_men_n47_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n87_));
  NOi21      u077(.An(i_7_), .B(i_8_), .Y(men_men_n88_));
  NOi31      u078(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n89_));
  AOI210     u079(.A0(men_men_n88_), .A1(men_men_n12_), .B0(men_men_n89_), .Y(men_men_n90_));
  OAI210     u080(.A0(men_men_n90_), .A1(men_men_n11_), .B0(men_men_n87_), .Y(men_men_n91_));
  OAI210     u081(.A0(men_men_n91_), .A1(men_men_n86_), .B0(men_men_n72_), .Y(men_men_n92_));
  NA3        u082(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n93_));
  AOI210     u083(.A0(men_men_n21_), .A1(men_men_n48_), .B0(men_men_n93_), .Y(men_men_n94_));
  NA3        u084(.A(men_men_n20_), .B(i_5_), .C(i_7_), .Y(men_men_n95_));
  OAI210     u085(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n96_));
  NA3        u086(.A(men_men_n68_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n97_));
  OAI220     u087(.A0(men_men_n97_), .A1(men_men_n96_), .B0(men_men_n95_), .B1(i_2_), .Y(men_men_n98_));
  NO2        u088(.A(men_men_n98_), .B(men_men_n94_), .Y(men_men_n99_));
  NA3        u089(.A(men_men_n63_), .B(men_men_n30_), .C(i_3_), .Y(men_men_n100_));
  NA2        u090(.A(men_men_n41_), .B(i_6_), .Y(men_men_n101_));
  AOI210     u091(.A0(men_men_n101_), .A1(men_men_n21_), .B0(men_men_n100_), .Y(men_men_n102_));
  NOi21      u092(.An(i_2_), .B(i_1_), .Y(men_men_n103_));
  NAi21      u093(.An(i_6_), .B(i_0_), .Y(men_men_n104_));
  NOi21      u094(.An(i_4_), .B(i_6_), .Y(men_men_n105_));
  NA2        u095(.A(men_men_n72_), .B(men_men_n32_), .Y(men_men_n106_));
  NOi21      u096(.An(men_men_n39_), .B(men_men_n106_), .Y(men_men_n107_));
  NO2        u097(.A(men_men_n107_), .B(men_men_n102_), .Y(men_men_n108_));
  NOi21      u098(.An(i_6_), .B(i_1_), .Y(men_men_n109_));
  AOI220     u099(.A0(men_men_n109_), .A1(i_7_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n110_));
  NOi31      u100(.An(men_men_n50_), .B(men_men_n110_), .C(i_2_), .Y(men_men_n111_));
  NA2        u101(.A(men_men_n63_), .B(men_men_n12_), .Y(men_men_n112_));
  NA2        u102(.A(men_men_n32_), .B(men_men_n14_), .Y(men_men_n113_));
  NOi21      u103(.An(i_3_), .B(i_1_), .Y(men_men_n114_));
  NA2        u104(.A(men_men_n114_), .B(i_4_), .Y(men_men_n115_));
  AOI210     u105(.A0(men_men_n113_), .A1(men_men_n112_), .B0(men_men_n115_), .Y(men_men_n116_));
  AOI220     u106(.A0(men_men_n88_), .A1(men_men_n14_), .B0(men_men_n105_), .B1(men_men_n22_), .Y(men_men_n117_));
  NOi31      u107(.An(men_men_n42_), .B(men_men_n117_), .C(men_men_n30_), .Y(men_men_n118_));
  NO3        u108(.A(men_men_n118_), .B(men_men_n116_), .C(men_men_n111_), .Y(men_men_n119_));
  NA4        u109(.A(men_men_n119_), .B(men_men_n108_), .C(men_men_n99_), .D(men_men_n92_), .Y(men_men_n120_));
  NA2        u110(.A(men_men_n53_), .B(men_men_n15_), .Y(men_men_n121_));
  NOi31      u111(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n122_));
  NA2        u112(.A(men_men_n122_), .B(i_7_), .Y(men_men_n123_));
  NA3        u113(.A(men_men_n32_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n124_));
  NA3        u114(.A(men_men_n124_), .B(men_men_n123_), .C(men_men_n121_), .Y(men_men_n125_));
  NA2        u115(.A(men_men_n125_), .B(men_men_n37_), .Y(men_men_n126_));
  NA2        u116(.A(men_men_n59_), .B(men_men_n33_), .Y(men_men_n127_));
  AOI210     u117(.A0(men_men_n127_), .A1(men_men_n76_), .B0(men_men_n29_), .Y(men_men_n128_));
  NAi31      u118(.An(men_men_n104_), .B(men_men_n88_), .C(men_men_n103_), .Y(men_men_n129_));
  NA3        u119(.A(men_men_n63_), .B(men_men_n57_), .C(i_6_), .Y(men_men_n130_));
  NA2        u120(.A(men_men_n130_), .B(men_men_n129_), .Y(men_men_n131_));
  NOi21      u121(.An(i_0_), .B(i_2_), .Y(men_men_n132_));
  NA3        u122(.A(men_men_n132_), .B(men_men_n33_), .C(men_men_n105_), .Y(men_men_n133_));
  NA3        u123(.A(men_men_n50_), .B(men_men_n39_), .C(men_men_n18_), .Y(men_men_n134_));
  NOi32      u124(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n135_));
  NA2        u125(.A(men_men_n135_), .B(men_men_n122_), .Y(men_men_n136_));
  NA3        u126(.A(men_men_n132_), .B(men_men_n59_), .C(men_men_n32_), .Y(men_men_n137_));
  NA4        u127(.A(men_men_n137_), .B(men_men_n136_), .C(men_men_n134_), .D(men_men_n133_), .Y(men_men_n138_));
  NA4        u128(.A(men_men_n57_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n139_));
  INV        u129(.A(men_men_n139_), .Y(men_men_n140_));
  NO4        u130(.A(men_men_n140_), .B(men_men_n138_), .C(men_men_n131_), .D(men_men_n128_), .Y(men_men_n141_));
  NO2        u131(.A(men_men_n121_), .B(men_men_n101_), .Y(men_men_n142_));
  NO3        u132(.A(i_2_), .B(men_men_n11_), .C(men_men_n14_), .Y(men_men_n143_));
  NA2        u133(.A(i_2_), .B(i_4_), .Y(men_men_n144_));
  AOI210     u134(.A0(men_men_n104_), .A1(i_3_), .B0(men_men_n144_), .Y(men_men_n145_));
  NO2        u135(.A(i_8_), .B(i_7_), .Y(men_men_n146_));
  OA210      u136(.A0(men_men_n145_), .A1(men_men_n143_), .B0(men_men_n146_), .Y(men_men_n147_));
  NO2        u137(.A(men_men_n147_), .B(men_men_n142_), .Y(men_men_n148_));
  NA2        u138(.A(men_men_n88_), .B(men_men_n12_), .Y(men_men_n149_));
  NA3        u139(.A(i_2_), .B(i_1_), .C(men_men_n14_), .Y(men_men_n150_));
  NA2        u140(.A(men_men_n50_), .B(i_3_), .Y(men_men_n151_));
  AOI210     u141(.A0(men_men_n151_), .A1(men_men_n150_), .B0(men_men_n149_), .Y(men_men_n152_));
  NA3        u142(.A(men_men_n132_), .B(men_men_n63_), .C(men_men_n105_), .Y(men_men_n153_));
  OAI210     u143(.A0(men_men_n100_), .A1(men_men_n29_), .B0(men_men_n153_), .Y(men_men_n154_));
  NA3        u144(.A(men_men_n53_), .B(men_men_n31_), .C(men_men_n15_), .Y(men_men_n155_));
  NOi31      u145(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n156_));
  OAI210     u146(.A0(men_men_n135_), .A1(men_men_n79_), .B0(men_men_n156_), .Y(men_men_n157_));
  NA2        u147(.A(men_men_n157_), .B(men_men_n155_), .Y(men_men_n158_));
  NO3        u148(.A(men_men_n158_), .B(men_men_n154_), .C(men_men_n152_), .Y(men_men_n159_));
  NA4        u149(.A(men_men_n159_), .B(men_men_n148_), .C(men_men_n141_), .D(men_men_n126_), .Y(men_men_n160_));
  OR4        u150(.A(men_men_n160_), .B(men_men_n120_), .C(men_men_n85_), .D(men_men_n67_), .Y(men00));
  INV        u151(.A(i_0_), .Y(men_men_n164_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule