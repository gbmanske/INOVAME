//Benchmark atmr_max1024_476_0.25

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n426_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  INV        o004(.A(ori_ori_n19_), .Y(ori_ori_n21_));
  NA2        o005(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n22_));
  INV        o006(.A(x5), .Y(ori_ori_n23_));
  NA2        o007(.A(x7), .B(x6), .Y(ori_ori_n24_));
  NA2        o008(.A(x4), .B(x2), .Y(ori_ori_n25_));
  INV        o009(.A(ori_ori_n22_), .Y(ori_ori_n26_));
  NO2        o010(.A(x4), .B(x3), .Y(ori_ori_n27_));
  INV        o011(.A(ori_ori_n27_), .Y(ori_ori_n28_));
  NOi21      o012(.An(ori_ori_n21_), .B(ori_ori_n26_), .Y(ori00));
  NO2        o013(.A(x1), .B(x0), .Y(ori_ori_n30_));
  INV        o014(.A(x6), .Y(ori_ori_n31_));
  NA2        o015(.A(x4), .B(x3), .Y(ori_ori_n32_));
  NO2        o016(.A(ori_ori_n21_), .B(ori_ori_n32_), .Y(ori_ori_n33_));
  NO2        o017(.A(x2), .B(x0), .Y(ori_ori_n34_));
  INV        o018(.A(x3), .Y(ori_ori_n35_));
  NO2        o019(.A(ori_ori_n35_), .B(ori_ori_n18_), .Y(ori_ori_n36_));
  INV        o020(.A(ori_ori_n36_), .Y(ori_ori_n37_));
  INV        o021(.A(x4), .Y(ori_ori_n38_));
  OAI210     o022(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n34_), .Y(ori_ori_n39_));
  INV        o023(.A(x4), .Y(ori_ori_n40_));
  NO2        o024(.A(ori_ori_n40_), .B(ori_ori_n17_), .Y(ori_ori_n41_));
  NA2        o025(.A(ori_ori_n41_), .B(x2), .Y(ori_ori_n42_));
  OAI210     o026(.A0(ori_ori_n42_), .A1(ori_ori_n20_), .B0(ori_ori_n39_), .Y(ori_ori_n43_));
  INV        o027(.A(ori_ori_n30_), .Y(ori_ori_n44_));
  INV        o028(.A(x2), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n45_), .B(ori_ori_n17_), .Y(ori_ori_n46_));
  NA2        o030(.A(ori_ori_n35_), .B(ori_ori_n18_), .Y(ori_ori_n47_));
  NA2        o031(.A(ori_ori_n47_), .B(ori_ori_n46_), .Y(ori_ori_n48_));
  OAI210     o032(.A0(ori_ori_n44_), .A1(ori_ori_n28_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  NO3        o033(.A(ori_ori_n49_), .B(ori_ori_n43_), .C(ori_ori_n33_), .Y(ori01));
  NA2        o034(.A(ori_ori_n35_), .B(x1), .Y(ori_ori_n51_));
  INV        o035(.A(x9), .Y(ori_ori_n52_));
  NO2        o036(.A(ori_ori_n51_), .B(x5), .Y(ori_ori_n53_));
  OAI210     o037(.A0(ori_ori_n36_), .A1(ori_ori_n23_), .B0(ori_ori_n45_), .Y(ori_ori_n54_));
  OAI210     o038(.A0(ori_ori_n47_), .A1(ori_ori_n20_), .B0(ori_ori_n54_), .Y(ori_ori_n55_));
  INV        o039(.A(ori_ori_n55_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(x4), .Y(ori_ori_n57_));
  NA2        o041(.A(ori_ori_n40_), .B(x2), .Y(ori_ori_n58_));
  OAI210     o042(.A0(ori_ori_n58_), .A1(ori_ori_n47_), .B0(x0), .Y(ori_ori_n59_));
  NA2        o043(.A(x5), .B(x3), .Y(ori_ori_n60_));
  NO2        o044(.A(x8), .B(x6), .Y(ori_ori_n61_));
  NO3        o045(.A(ori_ori_n61_), .B(ori_ori_n60_), .C(ori_ori_n45_), .Y(ori_ori_n62_));
  NAi21      o046(.An(x4), .B(x3), .Y(ori_ori_n63_));
  INV        o047(.A(ori_ori_n63_), .Y(ori_ori_n64_));
  NO2        o048(.A(x4), .B(x2), .Y(ori_ori_n65_));
  NO2        o049(.A(ori_ori_n63_), .B(ori_ori_n18_), .Y(ori_ori_n66_));
  NO3        o050(.A(ori_ori_n66_), .B(ori_ori_n62_), .C(ori_ori_n59_), .Y(ori_ori_n67_));
  NA2        o051(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n68_));
  NO2        o052(.A(ori_ori_n68_), .B(ori_ori_n23_), .Y(ori_ori_n69_));
  INV        o053(.A(x8), .Y(ori_ori_n70_));
  NA2        o054(.A(x2), .B(x1), .Y(ori_ori_n71_));
  AOI210     o055(.A0(ori_ori_n47_), .A1(ori_ori_n23_), .B0(ori_ori_n45_), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n37_), .B(ori_ori_n40_), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NA2        o058(.A(x4), .B(ori_ori_n35_), .Y(ori_ori_n75_));
  NO2        o059(.A(ori_ori_n40_), .B(ori_ori_n45_), .Y(ori_ori_n76_));
  NO2        o060(.A(ori_ori_n75_), .B(x1), .Y(ori_ori_n77_));
  NO2        o061(.A(x3), .B(x2), .Y(ori_ori_n78_));
  NA3        o062(.A(ori_ori_n78_), .B(ori_ori_n24_), .C(ori_ori_n23_), .Y(ori_ori_n79_));
  INV        o063(.A(ori_ori_n79_), .Y(ori_ori_n80_));
  NA2        o064(.A(ori_ori_n45_), .B(x1), .Y(ori_ori_n81_));
  OAI210     o065(.A0(ori_ori_n81_), .A1(ori_ori_n32_), .B0(ori_ori_n17_), .Y(ori_ori_n82_));
  NO4        o066(.A(ori_ori_n82_), .B(ori_ori_n80_), .C(ori_ori_n77_), .D(ori_ori_n74_), .Y(ori_ori_n83_));
  AO210      o067(.A0(ori_ori_n67_), .A1(ori_ori_n57_), .B0(ori_ori_n83_), .Y(ori02));
  NA2        o068(.A(ori_ori_n35_), .B(x0), .Y(ori_ori_n85_));
  BUFFER     o069(.A(x0), .Y(ori_ori_n86_));
  NO2        o070(.A(x4), .B(x1), .Y(ori_ori_n87_));
  NA2        o071(.A(ori_ori_n87_), .B(x2), .Y(ori_ori_n88_));
  NOi21      o072(.An(x0), .B(x4), .Y(ori_ori_n89_));
  NO2        o073(.A(ori_ori_n88_), .B(ori_ori_n60_), .Y(ori_ori_n90_));
  NO2        o074(.A(x5), .B(ori_ori_n40_), .Y(ori_ori_n91_));
  NA2        o075(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n92_));
  AOI210     o076(.A0(ori_ori_n92_), .A1(ori_ori_n81_), .B0(ori_ori_n85_), .Y(ori_ori_n93_));
  OAI210     o077(.A0(ori_ori_n93_), .A1(ori_ori_n30_), .B0(ori_ori_n91_), .Y(ori_ori_n94_));
  NAi21      o078(.An(x0), .B(x4), .Y(ori_ori_n95_));
  NO2        o079(.A(ori_ori_n95_), .B(x1), .Y(ori_ori_n96_));
  NO2        o080(.A(x7), .B(x0), .Y(ori_ori_n97_));
  NO2        o081(.A(ori_ori_n65_), .B(ori_ori_n76_), .Y(ori_ori_n98_));
  NO2        o082(.A(ori_ori_n98_), .B(x3), .Y(ori_ori_n99_));
  OAI210     o083(.A0(ori_ori_n97_), .A1(ori_ori_n96_), .B0(ori_ori_n99_), .Y(ori_ori_n100_));
  NA2        o084(.A(x5), .B(x0), .Y(ori_ori_n101_));
  NO2        o085(.A(ori_ori_n40_), .B(x2), .Y(ori_ori_n102_));
  NA3        o086(.A(ori_ori_n100_), .B(ori_ori_n94_), .C(ori_ori_n31_), .Y(ori_ori_n103_));
  NO2        o087(.A(ori_ori_n103_), .B(ori_ori_n90_), .Y(ori_ori_n104_));
  NO3        o088(.A(ori_ori_n60_), .B(ori_ori_n58_), .C(ori_ori_n22_), .Y(ori_ori_n105_));
  NO2        o089(.A(ori_ori_n25_), .B(ori_ori_n23_), .Y(ori_ori_n106_));
  NA2        o090(.A(x7), .B(x3), .Y(ori_ori_n107_));
  NO2        o091(.A(ori_ori_n75_), .B(x5), .Y(ori_ori_n108_));
  NO2        o092(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n109_));
  INV        o093(.A(x7), .Y(ori_ori_n110_));
  NA2        o094(.A(ori_ori_n110_), .B(ori_ori_n18_), .Y(ori_ori_n111_));
  NA2        o095(.A(ori_ori_n111_), .B(ori_ori_n109_), .Y(ori_ori_n112_));
  NO2        o096(.A(ori_ori_n23_), .B(x4), .Y(ori_ori_n113_));
  NO2        o097(.A(ori_ori_n113_), .B(ori_ori_n89_), .Y(ori_ori_n114_));
  NO2        o098(.A(ori_ori_n114_), .B(ori_ori_n112_), .Y(ori_ori_n115_));
  NA2        o099(.A(x5), .B(x1), .Y(ori_ori_n116_));
  INV        o100(.A(ori_ori_n116_), .Y(ori_ori_n117_));
  NAi21      o101(.An(x2), .B(x7), .Y(ori_ori_n118_));
  NO2        o102(.A(ori_ori_n118_), .B(ori_ori_n40_), .Y(ori_ori_n119_));
  NA2        o103(.A(ori_ori_n119_), .B(ori_ori_n53_), .Y(ori_ori_n120_));
  NA2        o104(.A(ori_ori_n120_), .B(x6), .Y(ori_ori_n121_));
  NO3        o105(.A(ori_ori_n121_), .B(ori_ori_n115_), .C(ori_ori_n105_), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n122_), .B(ori_ori_n104_), .Y(ori_ori_n123_));
  NO2        o107(.A(ori_ori_n101_), .B(ori_ori_n98_), .Y(ori_ori_n124_));
  NA2        o108(.A(ori_ori_n23_), .B(ori_ori_n18_), .Y(ori_ori_n125_));
  NA2        o109(.A(ori_ori_n23_), .B(ori_ori_n17_), .Y(ori_ori_n126_));
  NA3        o110(.A(ori_ori_n126_), .B(ori_ori_n125_), .C(ori_ori_n22_), .Y(ori_ori_n127_));
  AN2        o111(.A(ori_ori_n127_), .B(ori_ori_n102_), .Y(ori_ori_n128_));
  NA2        o112(.A(x8), .B(x0), .Y(ori_ori_n129_));
  NO2        o113(.A(ori_ori_n110_), .B(ori_ori_n23_), .Y(ori_ori_n130_));
  INV        o114(.A(x4), .Y(ori_ori_n131_));
  NA2        o115(.A(ori_ori_n131_), .B(ori_ori_n130_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n129_), .B(ori_ori_n132_), .Y(ori_ori_n133_));
  NA2        o117(.A(x2), .B(x0), .Y(ori_ori_n134_));
  NA2        o118(.A(x4), .B(x1), .Y(ori_ori_n135_));
  NAi21      o119(.An(ori_ori_n87_), .B(ori_ori_n135_), .Y(ori_ori_n136_));
  NOi31      o120(.An(ori_ori_n136_), .B(ori_ori_n113_), .C(ori_ori_n134_), .Y(ori_ori_n137_));
  NO4        o121(.A(ori_ori_n137_), .B(ori_ori_n133_), .C(ori_ori_n128_), .D(ori_ori_n124_), .Y(ori_ori_n138_));
  NO2        o122(.A(ori_ori_n138_), .B(ori_ori_n35_), .Y(ori_ori_n139_));
  NO2        o123(.A(ori_ori_n127_), .B(ori_ori_n58_), .Y(ori_ori_n140_));
  INV        o124(.A(ori_ori_n91_), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n81_), .B(ori_ori_n17_), .Y(ori_ori_n142_));
  AOI210     o126(.A0(ori_ori_n30_), .A1(ori_ori_n70_), .B0(ori_ori_n142_), .Y(ori_ori_n143_));
  NO3        o127(.A(ori_ori_n143_), .B(ori_ori_n141_), .C(x7), .Y(ori_ori_n144_));
  NA3        o128(.A(ori_ori_n136_), .B(ori_ori_n141_), .C(ori_ori_n34_), .Y(ori_ori_n145_));
  OAI210     o129(.A0(ori_ori_n126_), .A1(ori_ori_n98_), .B0(ori_ori_n145_), .Y(ori_ori_n146_));
  NO3        o130(.A(ori_ori_n146_), .B(ori_ori_n144_), .C(ori_ori_n140_), .Y(ori_ori_n147_));
  NO2        o131(.A(ori_ori_n147_), .B(x3), .Y(ori_ori_n148_));
  NO3        o132(.A(ori_ori_n148_), .B(ori_ori_n139_), .C(ori_ori_n123_), .Y(ori03));
  NO2        o133(.A(ori_ori_n40_), .B(x3), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n60_), .B(x6), .Y(ori_ori_n151_));
  NA2        o135(.A(x6), .B(ori_ori_n23_), .Y(ori_ori_n152_));
  NO2        o136(.A(ori_ori_n152_), .B(x4), .Y(ori_ori_n153_));
  AN2        o137(.A(ori_ori_n151_), .B(ori_ori_n46_), .Y(ori_ori_n154_));
  INV        o138(.A(ori_ori_n154_), .Y(ori_ori_n155_));
  NA2        o139(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n156_));
  NA2        o140(.A(x9), .B(ori_ori_n45_), .Y(ori_ori_n157_));
  NO3        o141(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n158_));
  NO2        o142(.A(x5), .B(x1), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n156_), .B(ori_ori_n125_), .Y(ori_ori_n160_));
  NO3        o144(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n161_));
  NO2        o145(.A(ori_ori_n161_), .B(ori_ori_n160_), .Y(ori_ori_n162_));
  INV        o146(.A(ori_ori_n162_), .Y(ori_ori_n163_));
  AOI220     o147(.A0(ori_ori_n163_), .A1(ori_ori_n40_), .B0(ori_ori_n158_), .B1(ori_ori_n91_), .Y(ori_ori_n164_));
  NA2        o148(.A(ori_ori_n164_), .B(ori_ori_n155_), .Y(ori_ori_n165_));
  NO2        o149(.A(ori_ori_n40_), .B(ori_ori_n35_), .Y(ori_ori_n166_));
  NA2        o150(.A(ori_ori_n166_), .B(ori_ori_n19_), .Y(ori_ori_n167_));
  NO2        o151(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n168_));
  NO2        o152(.A(ori_ori_n168_), .B(x6), .Y(ori_ori_n169_));
  NOi21      o153(.An(ori_ori_n65_), .B(ori_ori_n169_), .Y(ori_ori_n170_));
  NA2        o154(.A(ori_ori_n52_), .B(ori_ori_n70_), .Y(ori_ori_n171_));
  NA3        o155(.A(ori_ori_n171_), .B(ori_ori_n168_), .C(x6), .Y(ori_ori_n172_));
  AOI210     o156(.A0(ori_ori_n172_), .A1(ori_ori_n170_), .B0(ori_ori_n110_), .Y(ori_ori_n173_));
  OR2        o157(.A(ori_ori_n173_), .B(ori_ori_n130_), .Y(ori_ori_n174_));
  NA2        o158(.A(ori_ori_n35_), .B(ori_ori_n45_), .Y(ori_ori_n175_));
  NA2        o159(.A(ori_ori_n102_), .B(ori_ori_n69_), .Y(ori_ori_n176_));
  NA2        o160(.A(x6), .B(ori_ori_n40_), .Y(ori_ori_n177_));
  NA2        o161(.A(ori_ori_n61_), .B(x4), .Y(ori_ori_n178_));
  AOI210     o162(.A0(ori_ori_n178_), .A1(ori_ori_n177_), .B0(ori_ori_n60_), .Y(ori_ori_n179_));
  NA2        o163(.A(x5), .B(ori_ori_n96_), .Y(ori_ori_n180_));
  INV        o164(.A(ori_ori_n53_), .Y(ori_ori_n181_));
  NA2        o165(.A(ori_ori_n181_), .B(ori_ori_n180_), .Y(ori_ori_n182_));
  OAI210     o166(.A0(ori_ori_n182_), .A1(ori_ori_n179_), .B0(x2), .Y(ori_ori_n183_));
  NA3        o167(.A(ori_ori_n183_), .B(ori_ori_n176_), .C(ori_ori_n174_), .Y(ori_ori_n184_));
  AOI210     o168(.A0(ori_ori_n165_), .A1(x8), .B0(ori_ori_n184_), .Y(ori_ori_n185_));
  NO2        o169(.A(ori_ori_n70_), .B(x3), .Y(ori_ori_n186_));
  NA2        o170(.A(ori_ori_n186_), .B(ori_ori_n153_), .Y(ori_ori_n187_));
  NO2        o171(.A(ori_ori_n68_), .B(ori_ori_n23_), .Y(ori_ori_n188_));
  AOI210     o172(.A0(ori_ori_n169_), .A1(ori_ori_n113_), .B0(ori_ori_n188_), .Y(ori_ori_n189_));
  AOI210     o173(.A0(ori_ori_n189_), .A1(ori_ori_n187_), .B0(x2), .Y(ori_ori_n190_));
  AOI220     o174(.A0(ori_ori_n153_), .A1(ori_ori_n142_), .B0(x2), .B1(ori_ori_n53_), .Y(ori_ori_n191_));
  NA2        o175(.A(ori_ori_n156_), .B(x6), .Y(ori_ori_n192_));
  NO2        o176(.A(ori_ori_n156_), .B(x6), .Y(ori_ori_n193_));
  INV        o177(.A(ori_ori_n193_), .Y(ori_ori_n194_));
  NA3        o178(.A(ori_ori_n194_), .B(ori_ori_n192_), .C(ori_ori_n106_), .Y(ori_ori_n195_));
  NA3        o179(.A(ori_ori_n195_), .B(ori_ori_n191_), .C(ori_ori_n110_), .Y(ori_ori_n196_));
  NO2        o180(.A(ori_ori_n101_), .B(x3), .Y(ori_ori_n197_));
  NA2        o181(.A(x6), .B(x2), .Y(ori_ori_n198_));
  NA2        o182(.A(x4), .B(ori_ori_n197_), .Y(ori_ori_n199_));
  NO2        o183(.A(x3), .B(ori_ori_n152_), .Y(ori_ori_n200_));
  BUFFER     o184(.A(ori_ori_n200_), .Y(ori_ori_n201_));
  NA2        o185(.A(ori_ori_n201_), .B(ori_ori_n34_), .Y(ori_ori_n202_));
  AOI210     o186(.A0(ori_ori_n202_), .A1(ori_ori_n199_), .B0(x8), .Y(ori_ori_n203_));
  NA2        o187(.A(x0), .B(ori_ori_n20_), .Y(ori_ori_n204_));
  NO2        o188(.A(ori_ori_n204_), .B(ori_ori_n175_), .Y(ori_ori_n205_));
  NO4        o189(.A(ori_ori_n205_), .B(ori_ori_n203_), .C(ori_ori_n196_), .D(ori_ori_n190_), .Y(ori_ori_n206_));
  NA2        o190(.A(ori_ori_n193_), .B(x2), .Y(ori_ori_n207_));
  OAI210     o191(.A0(x0), .A1(x6), .B0(ori_ori_n36_), .Y(ori_ori_n208_));
  AOI210     o192(.A0(ori_ori_n208_), .A1(ori_ori_n207_), .B0(ori_ori_n141_), .Y(ori_ori_n209_));
  NOi21      o193(.An(ori_ori_n198_), .B(ori_ori_n17_), .Y(ori_ori_n210_));
  NA3        o194(.A(ori_ori_n210_), .B(ori_ori_n159_), .C(ori_ori_n32_), .Y(ori_ori_n211_));
  AOI210     o195(.A0(ori_ori_n31_), .A1(ori_ori_n45_), .B0(x0), .Y(ori_ori_n212_));
  NA3        o196(.A(ori_ori_n212_), .B(ori_ori_n117_), .C(ori_ori_n28_), .Y(ori_ori_n213_));
  NA2        o197(.A(x3), .B(x2), .Y(ori_ori_n214_));
  AOI220     o198(.A0(ori_ori_n214_), .A1(ori_ori_n175_), .B0(ori_ori_n213_), .B1(ori_ori_n211_), .Y(ori_ori_n215_));
  NO2        o199(.A(ori_ori_n212_), .B(ori_ori_n210_), .Y(ori_ori_n216_));
  AOI220     o200(.A0(ori_ori_n216_), .A1(ori_ori_n64_), .B0(ori_ori_n18_), .B1(ori_ori_n27_), .Y(ori_ori_n217_));
  NO2        o201(.A(ori_ori_n217_), .B(ori_ori_n23_), .Y(ori_ori_n218_));
  NA3        o202(.A(ori_ori_n31_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n219_));
  NO2        o203(.A(ori_ori_n212_), .B(ori_ori_n210_), .Y(ori_ori_n220_));
  INV        o204(.A(ori_ori_n160_), .Y(ori_ori_n221_));
  NA2        o205(.A(ori_ori_n31_), .B(ori_ori_n35_), .Y(ori_ori_n222_));
  NO2        o206(.A(ori_ori_n177_), .B(ori_ori_n221_), .Y(ori_ori_n223_));
  AO210      o207(.A0(ori_ori_n220_), .A1(ori_ori_n108_), .B0(ori_ori_n223_), .Y(ori_ori_n224_));
  NO4        o208(.A(ori_ori_n224_), .B(ori_ori_n218_), .C(ori_ori_n215_), .D(ori_ori_n209_), .Y(ori_ori_n225_));
  OAI210     o209(.A0(ori_ori_n206_), .A1(ori_ori_n185_), .B0(ori_ori_n225_), .Y(ori04));
  NA2        o210(.A(ori_ori_n45_), .B(ori_ori_n186_), .Y(ori_ori_n227_));
  NA2        o211(.A(x6), .B(ori_ori_n227_), .Y(ori_ori_n228_));
  NA2        o212(.A(ori_ori_n228_), .B(x6), .Y(ori_ori_n229_));
  OAI210     o213(.A0(ori_ori_n86_), .A1(ori_ori_n81_), .B0(ori_ori_n129_), .Y(ori_ori_n230_));
  NA3        o214(.A(ori_ori_n230_), .B(x6), .C(x3), .Y(ori_ori_n231_));
  AOI210     o215(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n232_));
  OAI220     o216(.A0(ori_ori_n232_), .A1(ori_ori_n222_), .B0(ori_ori_n312_), .B1(ori_ori_n219_), .Y(ori_ori_n233_));
  INV        o217(.A(ori_ori_n233_), .Y(ori_ori_n234_));
  NA2        o218(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n235_));
  INV        o219(.A(ori_ori_n235_), .Y(ori_ori_n236_));
  NA2        o220(.A(ori_ori_n236_), .B(ori_ori_n61_), .Y(ori_ori_n237_));
  NA3        o221(.A(ori_ori_n237_), .B(ori_ori_n234_), .C(ori_ori_n231_), .Y(ori_ori_n238_));
  NA2        o222(.A(ori_ori_n158_), .B(ori_ori_n65_), .Y(ori_ori_n239_));
  NA2        o223(.A(ori_ori_n239_), .B(ori_ori_n110_), .Y(ori_ori_n240_));
  AOI210     o224(.A0(ori_ori_n238_), .A1(x4), .B0(ori_ori_n240_), .Y(ori_ori_n241_));
  NA3        o225(.A(x0), .B(ori_ori_n157_), .C(ori_ori_n70_), .Y(ori_ori_n242_));
  XO2        o226(.A(x4), .B(x0), .Y(ori_ori_n243_));
  NA2        o227(.A(x4), .B(ori_ori_n71_), .Y(ori_ori_n244_));
  AOI210     o228(.A0(ori_ori_n244_), .A1(ori_ori_n242_), .B0(x3), .Y(ori_ori_n245_));
  NO2        o229(.A(ori_ori_n243_), .B(x2), .Y(ori_ori_n246_));
  INV        o230(.A(ori_ori_n246_), .Y(ori_ori_n247_));
  NA3        o231(.A(ori_ori_n247_), .B(ori_ori_n167_), .C(x6), .Y(ori_ori_n248_));
  NO2        o232(.A(ori_ori_n30_), .B(x2), .Y(ori_ori_n249_));
  OAI220     o233(.A0(ori_ori_n313_), .A1(x6), .B0(ori_ori_n248_), .B1(ori_ori_n245_), .Y(ori_ori_n250_));
  AO220      o234(.A0(x7), .A1(ori_ori_n250_), .B0(ori_ori_n241_), .B1(ori_ori_n229_), .Y(ori_ori_n251_));
  NA2        o235(.A(ori_ori_n249_), .B(x6), .Y(ori_ori_n252_));
  AOI210     o236(.A0(x6), .A1(x1), .B0(ori_ori_n109_), .Y(ori_ori_n253_));
  NA2        o237(.A(ori_ori_n311_), .B(x0), .Y(ori_ori_n254_));
  NA2        o238(.A(ori_ori_n65_), .B(x6), .Y(ori_ori_n255_));
  OAI210     o239(.A0(ori_ori_n254_), .A1(ori_ori_n253_), .B0(ori_ori_n255_), .Y(ori_ori_n256_));
  AOI220     o240(.A0(ori_ori_n256_), .A1(ori_ori_n252_), .B0(ori_ori_n161_), .B1(ori_ori_n41_), .Y(ori_ori_n257_));
  NA2        o241(.A(ori_ori_n257_), .B(ori_ori_n251_), .Y(ori_ori_n258_));
  NA2        o242(.A(ori_ori_n150_), .B(ori_ori_n110_), .Y(ori_ori_n259_));
  NA3        o243(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n260_));
  NA2        o244(.A(ori_ori_n166_), .B(x0), .Y(ori_ori_n261_));
  OAI220     o245(.A0(ori_ori_n261_), .A1(ori_ori_n157_), .B0(ori_ori_n260_), .B1(x2), .Y(ori_ori_n262_));
  INV        o246(.A(ori_ori_n262_), .Y(ori_ori_n263_));
  AOI210     o247(.A0(ori_ori_n263_), .A1(ori_ori_n259_), .B0(ori_ori_n23_), .Y(ori_ori_n264_));
  NAi21      o248(.An(ori_ori_n42_), .B(ori_ori_n130_), .Y(ori_ori_n265_));
  INV        o249(.A(ori_ori_n265_), .Y(ori_ori_n266_));
  OAI210     o250(.A0(ori_ori_n266_), .A1(ori_ori_n264_), .B0(x6), .Y(ori_ori_n267_));
  AOI220     o251(.A0(x7), .A1(ori_ori_n166_), .B0(ori_ori_n150_), .B1(ori_ori_n110_), .Y(ori_ori_n268_));
  INV        o252(.A(x1), .Y(ori_ori_n269_));
  OAI210     o253(.A0(ori_ori_n268_), .A1(x8), .B0(ori_ori_n269_), .Y(ori_ori_n270_));
  NAi31      o254(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n271_));
  OAI210     o255(.A0(ori_ori_n271_), .A1(x4), .B0(ori_ori_n118_), .Y(ori_ori_n272_));
  NA2        o256(.A(ori_ori_n272_), .B(ori_ori_n107_), .Y(ori_ori_n273_));
  NO2        o257(.A(ori_ori_n110_), .B(x0), .Y(ori_ori_n274_));
  NA2        o258(.A(ori_ori_n274_), .B(ori_ori_n186_), .Y(ori_ori_n275_));
  NA3        o259(.A(ori_ori_n275_), .B(x1), .C(ori_ori_n273_), .Y(ori_ori_n276_));
  NA2        o260(.A(ori_ori_n270_), .B(ori_ori_n276_), .Y(ori_ori_n277_));
  INV        o261(.A(ori_ori_n95_), .Y(ori_ori_n278_));
  NO2        o262(.A(ori_ori_n278_), .B(ori_ori_n35_), .Y(ori_ori_n279_));
  NO2        o263(.A(x1), .B(x0), .Y(ori_ori_n280_));
  NO2        o264(.A(ori_ori_n280_), .B(x3), .Y(ori_ori_n281_));
  NO3        o265(.A(ori_ori_n281_), .B(ori_ori_n279_), .C(x2), .Y(ori_ori_n282_));
  OAI210     o266(.A0(x4), .A1(ori_ori_n35_), .B0(ori_ori_n243_), .Y(ori_ori_n283_));
  INV        o267(.A(ori_ori_n260_), .Y(ori_ori_n284_));
  AOI220     o268(.A0(ori_ori_n284_), .A1(ori_ori_n70_), .B0(ori_ori_n283_), .B1(ori_ori_n110_), .Y(ori_ori_n285_));
  NO2        o269(.A(ori_ori_n285_), .B(ori_ori_n45_), .Y(ori_ori_n286_));
  NO2        o270(.A(ori_ori_n286_), .B(ori_ori_n282_), .Y(ori_ori_n287_));
  AOI210     o271(.A0(ori_ori_n287_), .A1(ori_ori_n277_), .B0(ori_ori_n23_), .Y(ori_ori_n288_));
  NA4        o272(.A(ori_ori_n27_), .B(ori_ori_n70_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n289_));
  NO3        o273(.A(ori_ori_n312_), .B(ori_ori_n129_), .C(ori_ori_n32_), .Y(ori_ori_n290_));
  NA2        o274(.A(ori_ori_n290_), .B(x7), .Y(ori_ori_n291_));
  NA2        o275(.A(ori_ori_n109_), .B(ori_ori_n96_), .Y(ori_ori_n292_));
  NA3        o276(.A(ori_ori_n292_), .B(ori_ori_n291_), .C(ori_ori_n289_), .Y(ori_ori_n293_));
  OAI210     o277(.A0(ori_ori_n293_), .A1(ori_ori_n288_), .B0(ori_ori_n31_), .Y(ori_ori_n294_));
  INV        o278(.A(ori_ori_n274_), .Y(ori_ori_n295_));
  NO4        o279(.A(ori_ori_n295_), .B(ori_ori_n60_), .C(x4), .D(ori_ori_n45_), .Y(ori_ori_n296_));
  NA2        o280(.A(x3), .B(x7), .Y(ori_ori_n297_));
  NO2        o281(.A(ori_ori_n116_), .B(ori_ori_n97_), .Y(ori_ori_n298_));
  NA2        o282(.A(ori_ori_n298_), .B(ori_ori_n297_), .Y(ori_ori_n299_));
  NO2        o283(.A(ori_ori_n299_), .B(ori_ori_n25_), .Y(ori_ori_n300_));
  OAI220     o284(.A0(x3), .A1(x2), .B0(ori_ori_n116_), .B1(ori_ori_n35_), .Y(ori_ori_n301_));
  NA2        o285(.A(x3), .B(ori_ori_n45_), .Y(ori_ori_n302_));
  NO2        o286(.A(ori_ori_n111_), .B(ori_ori_n302_), .Y(ori_ori_n303_));
  AOI220     o287(.A0(ori_ori_n303_), .A1(x0), .B0(ori_ori_n301_), .B1(ori_ori_n97_), .Y(ori_ori_n304_));
  NO2        o288(.A(ori_ori_n304_), .B(ori_ori_n177_), .Y(ori_ori_n305_));
  NO3        o289(.A(ori_ori_n305_), .B(ori_ori_n300_), .C(ori_ori_n296_), .Y(ori_ori_n306_));
  NA3        o290(.A(ori_ori_n306_), .B(ori_ori_n294_), .C(ori_ori_n267_), .Y(ori_ori_n307_));
  AOI210     o291(.A0(ori_ori_n258_), .A1(ori_ori_n23_), .B0(ori_ori_n307_), .Y(ori05));
  INV        o292(.A(x4), .Y(ori_ori_n311_));
  INV        o293(.A(x2), .Y(ori_ori_n312_));
  INV        o294(.A(ori_ori_n63_), .Y(ori_ori_n313_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  NOi21      m004(.An(mai_mai_n20_), .B(x7), .Y(mai_mai_n21_));
  NAi21      m005(.An(mai_mai_n21_), .B(mai_mai_n19_), .Y(mai_mai_n22_));
  NA2        m006(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n23_));
  INV        m007(.A(x5), .Y(mai_mai_n24_));
  NA2        m008(.A(x7), .B(x6), .Y(mai_mai_n25_));
  NA2        m009(.A(x8), .B(x3), .Y(mai_mai_n26_));
  NA2        m010(.A(x4), .B(x2), .Y(mai_mai_n27_));
  NO4        m011(.A(mai_mai_n27_), .B(mai_mai_n26_), .C(mai_mai_n25_), .D(mai_mai_n24_), .Y(mai_mai_n28_));
  NO2        m012(.A(mai_mai_n28_), .B(mai_mai_n23_), .Y(mai_mai_n29_));
  NO2        m013(.A(x4), .B(x3), .Y(mai_mai_n30_));
  INV        m014(.A(mai_mai_n30_), .Y(mai_mai_n31_));
  AN2        m015(.A(x2), .B(mai_mai_n19_), .Y(mai_mai_n32_));
  NOi31      m016(.An(mai_mai_n22_), .B(mai_mai_n32_), .C(mai_mai_n29_), .Y(mai00));
  NO2        m017(.A(x1), .B(x0), .Y(mai_mai_n34_));
  INV        m018(.A(x6), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n35_), .B(mai_mai_n24_), .Y(mai_mai_n36_));
  AN2        m020(.A(x8), .B(x7), .Y(mai_mai_n37_));
  NA3        m021(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(mai_mai_n34_), .Y(mai_mai_n38_));
  NA2        m022(.A(x4), .B(x3), .Y(mai_mai_n39_));
  AOI210     m023(.A0(mai_mai_n38_), .A1(mai_mai_n22_), .B0(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m024(.A(x2), .B(x0), .Y(mai_mai_n41_));
  INV        m025(.A(x3), .Y(mai_mai_n42_));
  NO2        m026(.A(mai_mai_n42_), .B(mai_mai_n18_), .Y(mai_mai_n43_));
  INV        m027(.A(mai_mai_n43_), .Y(mai_mai_n44_));
  NO2        m028(.A(mai_mai_n36_), .B(x4), .Y(mai_mai_n45_));
  OAI210     m029(.A0(mai_mai_n45_), .A1(mai_mai_n44_), .B0(mai_mai_n41_), .Y(mai_mai_n46_));
  INV        m030(.A(x4), .Y(mai_mai_n47_));
  NO2        m031(.A(mai_mai_n47_), .B(mai_mai_n17_), .Y(mai_mai_n48_));
  NA2        m032(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n49_));
  OAI210     m033(.A0(mai_mai_n49_), .A1(mai_mai_n20_), .B0(mai_mai_n46_), .Y(mai_mai_n50_));
  NA2        m034(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n51_));
  AOI220     m035(.A0(mai_mai_n51_), .A1(mai_mai_n34_), .B0(mai_mai_n21_), .B1(mai_mai_n19_), .Y(mai_mai_n52_));
  INV        m036(.A(x2), .Y(mai_mai_n53_));
  NO2        m037(.A(mai_mai_n53_), .B(mai_mai_n17_), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n42_), .B(mai_mai_n18_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  OAI210     m040(.A0(mai_mai_n52_), .A1(mai_mai_n31_), .B0(mai_mai_n56_), .Y(mai_mai_n57_));
  NO3        m041(.A(mai_mai_n57_), .B(mai_mai_n50_), .C(mai_mai_n40_), .Y(mai01));
  NA2        m042(.A(x8), .B(x7), .Y(mai_mai_n59_));
  NA2        m043(.A(mai_mai_n42_), .B(x1), .Y(mai_mai_n60_));
  INV        m044(.A(x9), .Y(mai_mai_n61_));
  NO2        m045(.A(mai_mai_n61_), .B(mai_mai_n35_), .Y(mai_mai_n62_));
  INV        m046(.A(mai_mai_n62_), .Y(mai_mai_n63_));
  NO2        m047(.A(mai_mai_n63_), .B(mai_mai_n60_), .Y(mai_mai_n64_));
  NO2        m048(.A(x7), .B(x6), .Y(mai_mai_n65_));
  NO2        m049(.A(mai_mai_n60_), .B(x5), .Y(mai_mai_n66_));
  NO2        m050(.A(x8), .B(x2), .Y(mai_mai_n67_));
  OA210      m051(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n65_), .Y(mai_mai_n68_));
  OAI210     m052(.A0(mai_mai_n43_), .A1(mai_mai_n24_), .B0(mai_mai_n53_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n55_), .A1(mai_mai_n20_), .B0(mai_mai_n69_), .Y(mai_mai_n70_));
  NAi21      m054(.An(x1), .B(x5), .Y(mai_mai_n71_));
  NO2        m055(.A(mai_mai_n70_), .B(mai_mai_n68_), .Y(mai_mai_n72_));
  OAI210     m056(.A0(mai_mai_n72_), .A1(mai_mai_n64_), .B0(x4), .Y(mai_mai_n73_));
  NA2        m057(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n74_));
  OAI210     m058(.A0(mai_mai_n74_), .A1(mai_mai_n55_), .B0(x0), .Y(mai_mai_n75_));
  NA2        m059(.A(x5), .B(x3), .Y(mai_mai_n76_));
  NO2        m060(.A(x8), .B(x6), .Y(mai_mai_n77_));
  NO4        m061(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(mai_mai_n65_), .D(mai_mai_n53_), .Y(mai_mai_n78_));
  NAi21      m062(.An(x4), .B(x3), .Y(mai_mai_n79_));
  INV        m063(.A(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m064(.A(mai_mai_n80_), .B(mai_mai_n21_), .Y(mai_mai_n81_));
  NO2        m065(.A(x4), .B(x2), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(x3), .Y(mai_mai_n83_));
  NO3        m067(.A(mai_mai_n83_), .B(mai_mai_n81_), .C(mai_mai_n18_), .Y(mai_mai_n84_));
  NO3        m068(.A(mai_mai_n84_), .B(mai_mai_n78_), .C(mai_mai_n75_), .Y(mai_mai_n85_));
  NO3        m069(.A(x6), .B(mai_mai_n42_), .C(x1), .Y(mai_mai_n86_));
  INV        m070(.A(x4), .Y(mai_mai_n87_));
  NA2        m071(.A(mai_mai_n86_), .B(mai_mai_n87_), .Y(mai_mai_n88_));
  NA2        m072(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n89_), .B(mai_mai_n24_), .Y(mai_mai_n90_));
  INV        m074(.A(x8), .Y(mai_mai_n91_));
  NA2        m075(.A(x2), .B(x1), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n91_), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n90_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n25_), .Y(mai_mai_n95_));
  AOI210     m079(.A0(mai_mai_n55_), .A1(mai_mai_n24_), .B0(mai_mai_n53_), .Y(mai_mai_n96_));
  OAI210     m080(.A0(mai_mai_n44_), .A1(mai_mai_n36_), .B0(mai_mai_n47_), .Y(mai_mai_n97_));
  NO3        m081(.A(mai_mai_n97_), .B(mai_mai_n96_), .C(mai_mai_n95_), .Y(mai_mai_n98_));
  NA2        m082(.A(x4), .B(mai_mai_n42_), .Y(mai_mai_n99_));
  NO2        m083(.A(mai_mai_n47_), .B(mai_mai_n53_), .Y(mai_mai_n100_));
  OAI210     m084(.A0(mai_mai_n100_), .A1(mai_mai_n42_), .B0(mai_mai_n18_), .Y(mai_mai_n101_));
  AOI210     m085(.A0(mai_mai_n99_), .A1(mai_mai_n51_), .B0(mai_mai_n101_), .Y(mai_mai_n102_));
  NO2        m086(.A(x3), .B(x2), .Y(mai_mai_n103_));
  NA2        m087(.A(mai_mai_n53_), .B(x1), .Y(mai_mai_n104_));
  OAI210     m088(.A0(mai_mai_n104_), .A1(mai_mai_n39_), .B0(mai_mai_n17_), .Y(mai_mai_n105_));
  NO3        m089(.A(mai_mai_n105_), .B(mai_mai_n102_), .C(mai_mai_n98_), .Y(mai_mai_n106_));
  AO220      m090(.A0(mai_mai_n106_), .A1(mai_mai_n88_), .B0(mai_mai_n85_), .B1(mai_mai_n73_), .Y(mai02));
  NO2        m091(.A(x3), .B(mai_mai_n53_), .Y(mai_mai_n108_));
  NO2        m092(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n109_));
  AOI220     m093(.A0(mai_mai_n53_), .A1(mai_mai_n109_), .B0(mai_mai_n108_), .B1(x4), .Y(mai_mai_n110_));
  NO3        m094(.A(mai_mai_n110_), .B(x7), .C(x5), .Y(mai_mai_n111_));
  OR2        m095(.A(x8), .B(x0), .Y(mai_mai_n112_));
  INV        m096(.A(mai_mai_n112_), .Y(mai_mai_n113_));
  NAi21      m097(.An(x2), .B(x8), .Y(mai_mai_n114_));
  INV        m098(.A(mai_mai_n114_), .Y(mai_mai_n115_));
  NO2        m099(.A(x4), .B(x1), .Y(mai_mai_n116_));
  NO3        m100(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n117_));
  NOi21      m101(.An(x0), .B(x4), .Y(mai_mai_n118_));
  NAi21      m102(.An(x8), .B(x7), .Y(mai_mai_n119_));
  NO2        m103(.A(mai_mai_n119_), .B(mai_mai_n61_), .Y(mai_mai_n120_));
  AOI220     m104(.A0(mai_mai_n120_), .A1(mai_mai_n118_), .B0(mai_mai_n117_), .B1(x0), .Y(mai_mai_n121_));
  NO2        m105(.A(mai_mai_n121_), .B(mai_mai_n76_), .Y(mai_mai_n122_));
  NO2        m106(.A(x5), .B(mai_mai_n47_), .Y(mai_mai_n123_));
  NA2        m107(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n124_));
  AOI210     m108(.A0(mai_mai_n124_), .A1(mai_mai_n104_), .B0(x3), .Y(mai_mai_n125_));
  OAI210     m109(.A0(mai_mai_n125_), .A1(mai_mai_n34_), .B0(mai_mai_n123_), .Y(mai_mai_n126_));
  NAi21      m110(.An(x0), .B(x4), .Y(mai_mai_n127_));
  NO2        m111(.A(mai_mai_n127_), .B(x1), .Y(mai_mai_n128_));
  NO2        m112(.A(x7), .B(x0), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n82_), .B(mai_mai_n100_), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n130_), .B(x3), .Y(mai_mai_n131_));
  OAI210     m115(.A0(mai_mai_n129_), .A1(mai_mai_n128_), .B0(mai_mai_n131_), .Y(mai_mai_n132_));
  NO2        m116(.A(x7), .B(mai_mai_n42_), .Y(mai_mai_n133_));
  NA2        m117(.A(x5), .B(x0), .Y(mai_mai_n134_));
  NO2        m118(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n135_));
  NA3        m119(.A(mai_mai_n135_), .B(mai_mai_n134_), .C(mai_mai_n133_), .Y(mai_mai_n136_));
  NA4        m120(.A(mai_mai_n136_), .B(mai_mai_n132_), .C(mai_mai_n126_), .D(mai_mai_n35_), .Y(mai_mai_n137_));
  NO3        m121(.A(mai_mai_n137_), .B(mai_mai_n122_), .C(mai_mai_n111_), .Y(mai_mai_n138_));
  NO3        m122(.A(mai_mai_n76_), .B(mai_mai_n74_), .C(mai_mai_n23_), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n27_), .B(mai_mai_n24_), .Y(mai_mai_n140_));
  AOI220     m124(.A0(x0), .A1(mai_mai_n140_), .B0(mai_mai_n66_), .B1(mai_mai_n17_), .Y(mai_mai_n141_));
  NO2        m125(.A(mai_mai_n141_), .B(mai_mai_n59_), .Y(mai_mai_n142_));
  NA2        m126(.A(x7), .B(x3), .Y(mai_mai_n143_));
  NO2        m127(.A(mai_mai_n99_), .B(x5), .Y(mai_mai_n144_));
  NO2        m128(.A(x9), .B(x7), .Y(mai_mai_n145_));
  NOi21      m129(.An(x8), .B(x0), .Y(mai_mai_n146_));
  NO2        m130(.A(mai_mai_n42_), .B(x2), .Y(mai_mai_n147_));
  INV        m131(.A(x7), .Y(mai_mai_n148_));
  AOI220     m132(.A0(x7), .A1(mai_mai_n147_), .B0(mai_mai_n108_), .B1(mai_mai_n37_), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n24_), .B(x4), .Y(mai_mai_n150_));
  NO2        m134(.A(mai_mai_n150_), .B(mai_mai_n118_), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n151_), .B(mai_mai_n149_), .Y(mai_mai_n152_));
  AOI210     m136(.A0(mai_mai_n146_), .A1(mai_mai_n144_), .B0(mai_mai_n152_), .Y(mai_mai_n153_));
  OAI210     m137(.A0(mai_mai_n143_), .A1(mai_mai_n49_), .B0(mai_mai_n153_), .Y(mai_mai_n154_));
  NA2        m138(.A(x5), .B(x1), .Y(mai_mai_n155_));
  INV        m139(.A(mai_mai_n155_), .Y(mai_mai_n156_));
  AOI210     m140(.A0(mai_mai_n156_), .A1(mai_mai_n118_), .B0(mai_mai_n35_), .Y(mai_mai_n157_));
  NO2        m141(.A(mai_mai_n61_), .B(mai_mai_n91_), .Y(mai_mai_n158_));
  NO3        m142(.A(x2), .B(mai_mai_n158_), .C(mai_mai_n47_), .Y(mai_mai_n159_));
  NA2        m143(.A(mai_mai_n159_), .B(mai_mai_n66_), .Y(mai_mai_n160_));
  NAi31      m144(.An(mai_mai_n76_), .B(mai_mai_n37_), .C(mai_mai_n34_), .Y(mai_mai_n161_));
  NA3        m145(.A(mai_mai_n161_), .B(mai_mai_n160_), .C(mai_mai_n157_), .Y(mai_mai_n162_));
  NO4        m146(.A(mai_mai_n162_), .B(mai_mai_n154_), .C(mai_mai_n142_), .D(mai_mai_n139_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n163_), .B(mai_mai_n138_), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n134_), .B(mai_mai_n130_), .Y(mai_mai_n165_));
  NA2        m149(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n166_));
  NA2        m150(.A(mai_mai_n24_), .B(mai_mai_n17_), .Y(mai_mai_n167_));
  NA3        m151(.A(mai_mai_n167_), .B(mai_mai_n166_), .C(mai_mai_n23_), .Y(mai_mai_n168_));
  AN2        m152(.A(mai_mai_n168_), .B(mai_mai_n135_), .Y(mai_mai_n169_));
  NO2        m153(.A(mai_mai_n148_), .B(mai_mai_n24_), .Y(mai_mai_n170_));
  NA2        m154(.A(x2), .B(x0), .Y(mai_mai_n171_));
  NA2        m155(.A(x4), .B(x1), .Y(mai_mai_n172_));
  NAi21      m156(.An(mai_mai_n116_), .B(mai_mai_n172_), .Y(mai_mai_n173_));
  NOi31      m157(.An(mai_mai_n173_), .B(mai_mai_n150_), .C(mai_mai_n171_), .Y(mai_mai_n174_));
  NO3        m158(.A(mai_mai_n174_), .B(mai_mai_n169_), .C(mai_mai_n165_), .Y(mai_mai_n175_));
  NO2        m159(.A(mai_mai_n175_), .B(mai_mai_n42_), .Y(mai_mai_n176_));
  NO2        m160(.A(mai_mai_n168_), .B(mai_mai_n74_), .Y(mai_mai_n177_));
  INV        m161(.A(mai_mai_n123_), .Y(mai_mai_n178_));
  NA2        m162(.A(mai_mai_n173_), .B(mai_mai_n41_), .Y(mai_mai_n179_));
  OAI210     m163(.A0(mai_mai_n167_), .A1(mai_mai_n130_), .B0(mai_mai_n179_), .Y(mai_mai_n180_));
  NO2        m164(.A(mai_mai_n180_), .B(mai_mai_n177_), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n181_), .B(x3), .Y(mai_mai_n182_));
  NO3        m166(.A(mai_mai_n182_), .B(mai_mai_n176_), .C(mai_mai_n164_), .Y(mai03));
  NO2        m167(.A(mai_mai_n47_), .B(x3), .Y(mai_mai_n184_));
  NO2        m168(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n185_));
  NO2        m169(.A(mai_mai_n53_), .B(x1), .Y(mai_mai_n186_));
  INV        m170(.A(mai_mai_n62_), .Y(mai_mai_n187_));
  NO2        m171(.A(mai_mai_n187_), .B(mai_mai_n17_), .Y(mai_mai_n188_));
  NA2        m172(.A(mai_mai_n188_), .B(mai_mai_n184_), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n76_), .B(x6), .Y(mai_mai_n190_));
  NA2        m174(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n192_));
  NA2        m176(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n193_), .B(mai_mai_n191_), .Y(mai_mai_n194_));
  NA2        m178(.A(x9), .B(mai_mai_n53_), .Y(mai_mai_n195_));
  NA2        m179(.A(mai_mai_n195_), .B(x4), .Y(mai_mai_n196_));
  NA2        m180(.A(mai_mai_n191_), .B(mai_mai_n79_), .Y(mai_mai_n197_));
  AOI210     m181(.A0(mai_mai_n24_), .A1(x3), .B0(mai_mai_n171_), .Y(mai_mai_n198_));
  AOI220     m182(.A0(mai_mai_n198_), .A1(mai_mai_n197_), .B0(mai_mai_n196_), .B1(mai_mai_n194_), .Y(mai_mai_n199_));
  NO2        m183(.A(x5), .B(x1), .Y(mai_mai_n200_));
  AOI220     m184(.A0(mai_mai_n200_), .A1(mai_mai_n17_), .B0(mai_mai_n103_), .B1(x5), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n193_), .B(mai_mai_n166_), .Y(mai_mai_n202_));
  NO3        m186(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n203_));
  NO2        m187(.A(mai_mai_n203_), .B(mai_mai_n202_), .Y(mai_mai_n204_));
  OAI210     m188(.A0(mai_mai_n201_), .A1(mai_mai_n63_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  NA2        m189(.A(mai_mai_n205_), .B(mai_mai_n47_), .Y(mai_mai_n206_));
  NA3        m190(.A(mai_mai_n206_), .B(mai_mai_n199_), .C(mai_mai_n189_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n47_), .B(mai_mai_n42_), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n208_), .B(mai_mai_n19_), .Y(mai_mai_n209_));
  NO2        m193(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n210_));
  INV        m194(.A(x6), .Y(mai_mai_n211_));
  NA2        m195(.A(mai_mai_n61_), .B(mai_mai_n91_), .Y(mai_mai_n212_));
  AO210      m196(.A0(x7), .A1(mai_mai_n209_), .B0(mai_mai_n170_), .Y(mai_mai_n213_));
  NA2        m197(.A(mai_mai_n42_), .B(mai_mai_n53_), .Y(mai_mai_n214_));
  OAI210     m198(.A0(mai_mai_n214_), .A1(mai_mai_n24_), .B0(mai_mai_n167_), .Y(mai_mai_n215_));
  NO2        m199(.A(mai_mai_n172_), .B(x6), .Y(mai_mai_n216_));
  AOI220     m200(.A0(mai_mai_n216_), .A1(mai_mai_n215_), .B0(mai_mai_n135_), .B1(mai_mai_n90_), .Y(mai_mai_n217_));
  NA2        m201(.A(x6), .B(mai_mai_n47_), .Y(mai_mai_n218_));
  OAI210     m202(.A0(mai_mai_n113_), .A1(mai_mai_n77_), .B0(x4), .Y(mai_mai_n219_));
  AOI210     m203(.A0(mai_mai_n219_), .A1(mai_mai_n218_), .B0(mai_mai_n76_), .Y(mai_mai_n220_));
  NO2        m204(.A(mai_mai_n61_), .B(x6), .Y(mai_mai_n221_));
  NO2        m205(.A(mai_mai_n155_), .B(mai_mai_n42_), .Y(mai_mai_n222_));
  OAI210     m206(.A0(mai_mai_n222_), .A1(mai_mai_n202_), .B0(mai_mai_n221_), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n185_), .B(mai_mai_n128_), .Y(mai_mai_n224_));
  NA3        m208(.A(mai_mai_n193_), .B(mai_mai_n123_), .C(x6), .Y(mai_mai_n225_));
  OAI210     m209(.A0(mai_mai_n91_), .A1(mai_mai_n35_), .B0(mai_mai_n66_), .Y(mai_mai_n226_));
  NA4        m210(.A(mai_mai_n226_), .B(mai_mai_n225_), .C(mai_mai_n224_), .D(mai_mai_n223_), .Y(mai_mai_n227_));
  OAI210     m211(.A0(mai_mai_n227_), .A1(mai_mai_n220_), .B0(x2), .Y(mai_mai_n228_));
  NA3        m212(.A(mai_mai_n228_), .B(mai_mai_n217_), .C(mai_mai_n213_), .Y(mai_mai_n229_));
  AOI210     m213(.A0(mai_mai_n207_), .A1(x8), .B0(mai_mai_n229_), .Y(mai_mai_n230_));
  NO3        m214(.A(mai_mai_n89_), .B(mai_mai_n77_), .C(mai_mai_n24_), .Y(mai_mai_n231_));
  AOI210     m215(.A0(mai_mai_n211_), .A1(mai_mai_n150_), .B0(mai_mai_n231_), .Y(mai_mai_n232_));
  NO2        m216(.A(mai_mai_n232_), .B(x2), .Y(mai_mai_n233_));
  NO2        m217(.A(x4), .B(mai_mai_n53_), .Y(mai_mai_n234_));
  NA2        m218(.A(mai_mai_n234_), .B(mai_mai_n66_), .Y(mai_mai_n235_));
  NO2        m219(.A(mai_mai_n134_), .B(x9), .Y(mai_mai_n236_));
  NA2        m220(.A(mai_mai_n42_), .B(mai_mai_n17_), .Y(mai_mai_n237_));
  NO2        m221(.A(mai_mai_n237_), .B(mai_mai_n24_), .Y(mai_mai_n238_));
  OAI210     m222(.A0(mai_mai_n238_), .A1(mai_mai_n236_), .B0(mai_mai_n116_), .Y(mai_mai_n239_));
  NA2        m223(.A(mai_mai_n193_), .B(x6), .Y(mai_mai_n240_));
  NA2        m224(.A(mai_mai_n240_), .B(mai_mai_n140_), .Y(mai_mai_n241_));
  NA4        m225(.A(mai_mai_n241_), .B(mai_mai_n239_), .C(mai_mai_n235_), .D(mai_mai_n148_), .Y(mai_mai_n242_));
  NA2        m226(.A(mai_mai_n185_), .B(mai_mai_n210_), .Y(mai_mai_n243_));
  NO2        m227(.A(mai_mai_n134_), .B(mai_mai_n18_), .Y(mai_mai_n244_));
  AOI210     m228(.A0(x3), .A1(x2), .B0(mai_mai_n47_), .Y(mai_mai_n245_));
  INV        m229(.A(mai_mai_n245_), .Y(mai_mai_n246_));
  NO2        m230(.A(mai_mai_n244_), .B(mai_mai_n246_), .Y(mai_mai_n247_));
  NA2        m231(.A(mai_mai_n247_), .B(mai_mai_n243_), .Y(mai_mai_n248_));
  INV        m232(.A(mai_mai_n243_), .Y(mai_mai_n249_));
  NO3        m233(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n250_));
  NA2        m234(.A(mai_mai_n104_), .B(mai_mai_n24_), .Y(mai_mai_n251_));
  NA2        m235(.A(mai_mai_n251_), .B(mai_mai_n250_), .Y(mai_mai_n252_));
  OAI210     m236(.A0(mai_mai_n252_), .A1(mai_mai_n42_), .B0(mai_mai_n397_), .Y(mai_mai_n253_));
  OAI210     m237(.A0(mai_mai_n253_), .A1(mai_mai_n249_), .B0(mai_mai_n248_), .Y(mai_mai_n254_));
  NA2        m238(.A(x4), .B(x0), .Y(mai_mai_n255_));
  NA2        m239(.A(mai_mai_n190_), .B(mai_mai_n41_), .Y(mai_mai_n256_));
  AOI210     m240(.A0(mai_mai_n256_), .A1(mai_mai_n254_), .B0(x8), .Y(mai_mai_n257_));
  OAI210     m241(.A0(mai_mai_n244_), .A1(mai_mai_n200_), .B0(x6), .Y(mai_mai_n258_));
  NO2        m242(.A(mai_mai_n258_), .B(mai_mai_n214_), .Y(mai_mai_n259_));
  NO4        m243(.A(mai_mai_n259_), .B(mai_mai_n257_), .C(mai_mai_n242_), .D(mai_mai_n233_), .Y(mai_mai_n260_));
  NO2        m244(.A(x3), .B(mai_mai_n35_), .Y(mai_mai_n261_));
  NA2        m245(.A(mai_mai_n261_), .B(x2), .Y(mai_mai_n262_));
  NA2        m246(.A(x6), .B(mai_mai_n43_), .Y(mai_mai_n263_));
  AOI210     m247(.A0(mai_mai_n263_), .A1(mai_mai_n262_), .B0(mai_mai_n178_), .Y(mai_mai_n264_));
  NA3        m248(.A(x0), .B(mai_mai_n200_), .C(mai_mai_n39_), .Y(mai_mai_n265_));
  AOI210     m249(.A0(mai_mai_n35_), .A1(mai_mai_n53_), .B0(x0), .Y(mai_mai_n266_));
  NA3        m250(.A(mai_mai_n266_), .B(mai_mai_n156_), .C(mai_mai_n31_), .Y(mai_mai_n267_));
  NA2        m251(.A(x3), .B(x2), .Y(mai_mai_n268_));
  AOI220     m252(.A0(mai_mai_n268_), .A1(mai_mai_n214_), .B0(mai_mai_n267_), .B1(mai_mai_n265_), .Y(mai_mai_n269_));
  NAi21      m253(.An(x4), .B(x0), .Y(mai_mai_n270_));
  NO3        m254(.A(mai_mai_n270_), .B(mai_mai_n43_), .C(x2), .Y(mai_mai_n271_));
  OAI210     m255(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n271_), .Y(mai_mai_n272_));
  OAI220     m256(.A0(mai_mai_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n273_));
  NO2        m257(.A(x9), .B(x8), .Y(mai_mai_n274_));
  NA3        m258(.A(mai_mai_n274_), .B(mai_mai_n35_), .C(mai_mai_n53_), .Y(mai_mai_n275_));
  OAI210     m259(.A0(mai_mai_n266_), .A1(x0), .B0(mai_mai_n275_), .Y(mai_mai_n276_));
  AOI220     m260(.A0(mai_mai_n276_), .A1(mai_mai_n80_), .B0(mai_mai_n273_), .B1(mai_mai_n30_), .Y(mai_mai_n277_));
  AOI210     m261(.A0(mai_mai_n277_), .A1(mai_mai_n272_), .B0(mai_mai_n24_), .Y(mai_mai_n278_));
  INV        m262(.A(mai_mai_n202_), .Y(mai_mai_n279_));
  NA2        m263(.A(mai_mai_n35_), .B(mai_mai_n42_), .Y(mai_mai_n280_));
  OR2        m264(.A(mai_mai_n280_), .B(mai_mai_n255_), .Y(mai_mai_n281_));
  OAI220     m265(.A0(mai_mai_n281_), .A1(mai_mai_n155_), .B0(mai_mai_n218_), .B1(mai_mai_n279_), .Y(mai_mai_n282_));
  NO4        m266(.A(mai_mai_n282_), .B(mai_mai_n278_), .C(mai_mai_n269_), .D(mai_mai_n264_), .Y(mai_mai_n283_));
  OAI210     m267(.A0(mai_mai_n260_), .A1(mai_mai_n230_), .B0(mai_mai_n283_), .Y(mai04));
  NA2        m268(.A(mai_mai_n250_), .B(mai_mai_n83_), .Y(mai_mai_n285_));
  NA2        m269(.A(mai_mai_n237_), .B(mai_mai_n35_), .Y(mai_mai_n286_));
  INV        m270(.A(mai_mai_n89_), .Y(mai_mai_n287_));
  NO2        m271(.A(mai_mai_n287_), .B(mai_mai_n35_), .Y(mai_mai_n288_));
  NO2        m272(.A(mai_mai_n268_), .B(mai_mai_n192_), .Y(mai_mai_n289_));
  NA2        m273(.A(x9), .B(x0), .Y(mai_mai_n290_));
  NO2        m274(.A(mai_mai_n74_), .B(mai_mai_n290_), .Y(mai_mai_n291_));
  OAI210     m275(.A0(mai_mai_n291_), .A1(mai_mai_n289_), .B0(mai_mai_n91_), .Y(mai_mai_n292_));
  NA2        m276(.A(mai_mai_n292_), .B(mai_mai_n288_), .Y(mai_mai_n293_));
  NA2        m277(.A(mai_mai_n293_), .B(mai_mai_n286_), .Y(mai_mai_n294_));
  NO2        m278(.A(mai_mai_n195_), .B(x3), .Y(mai_mai_n295_));
  INV        m279(.A(mai_mai_n295_), .Y(mai_mai_n296_));
  NA2        m280(.A(mai_mai_n18_), .B(mai_mai_n62_), .Y(mai_mai_n297_));
  NA2        m281(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n298_));
  NA3        m282(.A(mai_mai_n399_), .B(mai_mai_n297_), .C(mai_mai_n296_), .Y(mai_mai_n299_));
  OAI210     m283(.A0(mai_mai_n109_), .A1(x3), .B0(mai_mai_n271_), .Y(mai_mai_n300_));
  NA2        m284(.A(mai_mai_n300_), .B(mai_mai_n148_), .Y(mai_mai_n301_));
  AOI210     m285(.A0(mai_mai_n299_), .A1(x4), .B0(mai_mai_n301_), .Y(mai_mai_n302_));
  NOi21      m286(.An(x4), .B(x0), .Y(mai_mai_n303_));
  AOI220     m287(.A0(x2), .A1(x8), .B0(mai_mai_n303_), .B1(mai_mai_n92_), .Y(mai_mai_n304_));
  NO2        m288(.A(mai_mai_n304_), .B(x3), .Y(mai_mai_n305_));
  INV        m289(.A(mai_mai_n92_), .Y(mai_mai_n306_));
  NO2        m290(.A(mai_mai_n91_), .B(x4), .Y(mai_mai_n307_));
  AOI220     m291(.A0(mai_mai_n307_), .A1(mai_mai_n43_), .B0(mai_mai_n118_), .B1(mai_mai_n306_), .Y(mai_mai_n308_));
  NO3        m292(.A(mai_mai_n212_), .B(mai_mai_n27_), .C(mai_mai_n23_), .Y(mai_mai_n309_));
  INV        m293(.A(mai_mai_n309_), .Y(mai_mai_n310_));
  NA4        m294(.A(mai_mai_n310_), .B(mai_mai_n308_), .C(mai_mai_n209_), .D(x6), .Y(mai_mai_n311_));
  NO2        m295(.A(mai_mai_n171_), .B(mai_mai_n91_), .Y(mai_mai_n312_));
  NO2        m296(.A(mai_mai_n42_), .B(x0), .Y(mai_mai_n313_));
  OR2        m297(.A(mai_mai_n307_), .B(mai_mai_n313_), .Y(mai_mai_n314_));
  NO2        m298(.A(mai_mai_n146_), .B(mai_mai_n104_), .Y(mai_mai_n315_));
  AOI220     m299(.A0(mai_mai_n315_), .A1(mai_mai_n314_), .B0(mai_mai_n312_), .B1(mai_mai_n60_), .Y(mai_mai_n316_));
  NO2        m300(.A(mai_mai_n146_), .B(mai_mai_n79_), .Y(mai_mai_n317_));
  NO2        m301(.A(mai_mai_n34_), .B(x2), .Y(mai_mai_n318_));
  NOi21      m302(.An(mai_mai_n116_), .B(mai_mai_n26_), .Y(mai_mai_n319_));
  AOI210     m303(.A0(mai_mai_n318_), .A1(mai_mai_n317_), .B0(mai_mai_n319_), .Y(mai_mai_n320_));
  OAI210     m304(.A0(mai_mai_n316_), .A1(mai_mai_n61_), .B0(mai_mai_n320_), .Y(mai_mai_n321_));
  OAI220     m305(.A0(mai_mai_n321_), .A1(x6), .B0(mai_mai_n311_), .B1(mai_mai_n305_), .Y(mai_mai_n322_));
  OAI210     m306(.A0(mai_mai_n62_), .A1(mai_mai_n47_), .B0(mai_mai_n41_), .Y(mai_mai_n323_));
  OAI210     m307(.A0(mai_mai_n323_), .A1(mai_mai_n91_), .B0(mai_mai_n281_), .Y(mai_mai_n324_));
  AOI210     m308(.A0(mai_mai_n324_), .A1(mai_mai_n18_), .B0(mai_mai_n148_), .Y(mai_mai_n325_));
  AO220      m309(.A0(mai_mai_n325_), .A1(mai_mai_n322_), .B0(mai_mai_n302_), .B1(mai_mai_n294_), .Y(mai_mai_n326_));
  NA2        m310(.A(mai_mai_n82_), .B(x6), .Y(mai_mai_n327_));
  AOI220     m311(.A0(mai_mai_n396_), .A1(mai_mai_n34_), .B0(mai_mai_n203_), .B1(mai_mai_n48_), .Y(mai_mai_n328_));
  NA3        m312(.A(mai_mai_n328_), .B(mai_mai_n326_), .C(mai_mai_n285_), .Y(mai_mai_n329_));
  AOI210     m313(.A0(mai_mai_n186_), .A1(x8), .B0(mai_mai_n109_), .Y(mai_mai_n330_));
  NA2        m314(.A(mai_mai_n330_), .B(mai_mai_n298_), .Y(mai_mai_n331_));
  NA3        m315(.A(mai_mai_n331_), .B(mai_mai_n184_), .C(mai_mai_n148_), .Y(mai_mai_n332_));
  OAI210     m316(.A0(mai_mai_n27_), .A1(x1), .B0(mai_mai_n214_), .Y(mai_mai_n333_));
  AO220      m317(.A0(mai_mai_n333_), .A1(mai_mai_n145_), .B0(mai_mai_n108_), .B1(x4), .Y(mai_mai_n334_));
  NA3        m318(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n335_));
  NO2        m319(.A(mai_mai_n335_), .B(mai_mai_n306_), .Y(mai_mai_n336_));
  AOI210     m320(.A0(mai_mai_n334_), .A1(mai_mai_n113_), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  AOI210     m321(.A0(mai_mai_n337_), .A1(mai_mai_n332_), .B0(mai_mai_n24_), .Y(mai_mai_n338_));
  NA3        m322(.A(mai_mai_n115_), .B(mai_mai_n208_), .C(x0), .Y(mai_mai_n339_));
  OAI210     m323(.A0(mai_mai_n184_), .A1(mai_mai_n67_), .B0(mai_mai_n192_), .Y(mai_mai_n340_));
  NO2        m324(.A(mai_mai_n340_), .B(mai_mai_n24_), .Y(mai_mai_n341_));
  AOI210     m325(.A0(mai_mai_n114_), .A1(mai_mai_n112_), .B0(mai_mai_n41_), .Y(mai_mai_n342_));
  NOi31      m326(.An(mai_mai_n342_), .B(mai_mai_n313_), .C(mai_mai_n172_), .Y(mai_mai_n343_));
  OAI210     m327(.A0(mai_mai_n343_), .A1(mai_mai_n341_), .B0(mai_mai_n145_), .Y(mai_mai_n344_));
  NA2        m328(.A(mai_mai_n344_), .B(mai_mai_n339_), .Y(mai_mai_n345_));
  OAI210     m329(.A0(mai_mai_n345_), .A1(mai_mai_n338_), .B0(x6), .Y(mai_mai_n346_));
  AOI210     m330(.A0(mai_mai_n400_), .A1(x0), .B0(mai_mai_n31_), .Y(mai_mai_n347_));
  AOI220     m331(.A0(mai_mai_n398_), .A1(mai_mai_n208_), .B0(mai_mai_n184_), .B1(mai_mai_n148_), .Y(mai_mai_n348_));
  AOI210     m332(.A0(mai_mai_n120_), .A1(mai_mai_n234_), .B0(x1), .Y(mai_mai_n349_));
  OAI210     m333(.A0(mai_mai_n348_), .A1(x8), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  NO4        m334(.A(mai_mai_n119_), .B(mai_mai_n270_), .C(x9), .D(x2), .Y(mai_mai_n351_));
  NOi21      m335(.An(mai_mai_n117_), .B(mai_mai_n171_), .Y(mai_mai_n352_));
  NO3        m336(.A(mai_mai_n352_), .B(mai_mai_n351_), .C(mai_mai_n18_), .Y(mai_mai_n353_));
  NA2        m337(.A(mai_mai_n317_), .B(mai_mai_n148_), .Y(mai_mai_n354_));
  NA3        m338(.A(mai_mai_n354_), .B(mai_mai_n353_), .C(mai_mai_n49_), .Y(mai_mai_n355_));
  OAI210     m339(.A0(mai_mai_n350_), .A1(mai_mai_n347_), .B0(mai_mai_n355_), .Y(mai_mai_n356_));
  NOi31      m340(.An(mai_mai_n398_), .B(mai_mai_n31_), .C(x8), .Y(mai_mai_n357_));
  NO2        m341(.A(mai_mai_n117_), .B(mai_mai_n42_), .Y(mai_mai_n358_));
  NOi31      m342(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n359_));
  AOI210     m343(.A0(mai_mai_n118_), .A1(x3), .B0(mai_mai_n303_), .Y(mai_mai_n360_));
  NA2        m344(.A(x3), .B(mai_mai_n360_), .Y(mai_mai_n361_));
  NO3        m345(.A(mai_mai_n361_), .B(mai_mai_n358_), .C(x2), .Y(mai_mai_n362_));
  AOI210     m346(.A0(x9), .A1(mai_mai_n47_), .B0(mai_mai_n335_), .Y(mai_mai_n363_));
  NA2        m347(.A(mai_mai_n363_), .B(mai_mai_n91_), .Y(mai_mai_n364_));
  NO2        m348(.A(mai_mai_n364_), .B(mai_mai_n53_), .Y(mai_mai_n365_));
  NO3        m349(.A(mai_mai_n365_), .B(mai_mai_n362_), .C(mai_mai_n357_), .Y(mai_mai_n366_));
  AOI210     m350(.A0(mai_mai_n366_), .A1(mai_mai_n356_), .B0(mai_mai_n24_), .Y(mai_mai_n367_));
  NO3        m351(.A(mai_mai_n61_), .B(x4), .C(x1), .Y(mai_mai_n368_));
  NO3        m352(.A(mai_mai_n67_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n369_));
  AOI220     m353(.A0(mai_mai_n369_), .A1(mai_mai_n245_), .B0(mai_mai_n368_), .B1(mai_mai_n342_), .Y(mai_mai_n370_));
  NO2        m354(.A(mai_mai_n370_), .B(mai_mai_n103_), .Y(mai_mai_n371_));
  NA2        m355(.A(mai_mai_n371_), .B(x7), .Y(mai_mai_n372_));
  NA2        m356(.A(mai_mai_n212_), .B(x7), .Y(mai_mai_n373_));
  NA2        m357(.A(mai_mai_n373_), .B(mai_mai_n128_), .Y(mai_mai_n374_));
  NA2        m358(.A(mai_mai_n374_), .B(mai_mai_n372_), .Y(mai_mai_n375_));
  OAI210     m359(.A0(mai_mai_n375_), .A1(mai_mai_n367_), .B0(mai_mai_n35_), .Y(mai_mai_n376_));
  INV        m360(.A(mai_mai_n192_), .Y(mai_mai_n377_));
  NO4        m361(.A(mai_mai_n377_), .B(mai_mai_n76_), .C(x4), .D(mai_mai_n53_), .Y(mai_mai_n378_));
  NO2        m362(.A(mai_mai_n161_), .B(mai_mai_n27_), .Y(mai_mai_n379_));
  AOI220     m363(.A0(mai_mai_n313_), .A1(mai_mai_n91_), .B0(mai_mai_n146_), .B1(mai_mai_n186_), .Y(mai_mai_n380_));
  NA2        m364(.A(mai_mai_n380_), .B(mai_mai_n89_), .Y(mai_mai_n381_));
  NA2        m365(.A(mai_mai_n381_), .B(mai_mai_n170_), .Y(mai_mai_n382_));
  AOI210     m366(.A0(x2), .A1(mai_mai_n26_), .B0(mai_mai_n71_), .Y(mai_mai_n383_));
  NO3        m367(.A(mai_mai_n359_), .B(x3), .C(mai_mai_n53_), .Y(mai_mai_n384_));
  NO2        m368(.A(mai_mai_n384_), .B(mai_mai_n383_), .Y(mai_mai_n385_));
  INV        m369(.A(mai_mai_n385_), .Y(mai_mai_n386_));
  NA2        m370(.A(mai_mai_n386_), .B(x0), .Y(mai_mai_n387_));
  AOI210     m371(.A0(mai_mai_n387_), .A1(mai_mai_n382_), .B0(mai_mai_n218_), .Y(mai_mai_n388_));
  INV        m372(.A(x5), .Y(mai_mai_n389_));
  NO4        m373(.A(mai_mai_n104_), .B(mai_mai_n389_), .C(mai_mai_n59_), .D(mai_mai_n31_), .Y(mai_mai_n390_));
  NO4        m374(.A(mai_mai_n390_), .B(mai_mai_n388_), .C(mai_mai_n379_), .D(mai_mai_n378_), .Y(mai_mai_n391_));
  NA3        m375(.A(mai_mai_n391_), .B(mai_mai_n376_), .C(mai_mai_n346_), .Y(mai_mai_n392_));
  AOI210     m376(.A0(mai_mai_n329_), .A1(mai_mai_n24_), .B0(mai_mai_n392_), .Y(mai05));
  INV        m377(.A(mai_mai_n327_), .Y(mai_mai_n396_));
  INV        m378(.A(x4), .Y(mai_mai_n397_));
  INV        m379(.A(x0), .Y(mai_mai_n398_));
  INV        m380(.A(mai_mai_n77_), .Y(mai_mai_n399_));
  INV        m381(.A(mai_mai_n37_), .Y(mai_mai_n400_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  AN2        u016(.A(men_men_n32_), .B(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  AN2        u021(.A(x8), .B(x7), .Y(men_men_n38_));
  NA2        u022(.A(men_men_n38_), .B(men_men_n35_), .Y(men_men_n39_));
  NA2        u023(.A(x4), .B(x3), .Y(men_men_n40_));
  AOI210     u024(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n40_), .Y(men_men_n41_));
  NO2        u025(.A(x2), .B(x0), .Y(men_men_n42_));
  INV        u026(.A(x3), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n44_));
  INV        u028(.A(men_men_n44_), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n37_), .B(x4), .Y(men_men_n46_));
  OAI210     u030(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n42_), .Y(men_men_n47_));
  INV        u031(.A(x4), .Y(men_men_n48_));
  NO2        u032(.A(men_men_n48_), .B(men_men_n17_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(x2), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n50_), .B(men_men_n47_), .Y(men_men_n51_));
  NA2        u035(.A(men_men_n38_), .B(men_men_n37_), .Y(men_men_n52_));
  AOI220     u036(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n53_));
  INV        u037(.A(x2), .Y(men_men_n54_));
  NO2        u038(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n56_));
  NA2        u040(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  OAI210     u041(.A0(men_men_n53_), .A1(men_men_n32_), .B0(men_men_n57_), .Y(men_men_n58_));
  NO3        u042(.A(men_men_n58_), .B(men_men_n51_), .C(men_men_n41_), .Y(men01));
  NA2        u043(.A(x8), .B(x7), .Y(men_men_n60_));
  NA2        u044(.A(men_men_n43_), .B(x1), .Y(men_men_n61_));
  INV        u045(.A(x9), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n61_), .B(men_men_n60_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n61_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  NO2        u051(.A(men_men_n67_), .B(x1), .Y(men_men_n68_));
  OA210      u052(.A0(men_men_n68_), .A1(men_men_n65_), .B0(men_men_n64_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n56_), .A1(men_men_n20_), .B0(men_men_n70_), .Y(men_men_n71_));
  NAi31      u055(.An(x1), .B(x9), .C(x5), .Y(men_men_n72_));
  OAI220     u056(.A0(men_men_n72_), .A1(men_men_n43_), .B0(men_men_n71_), .B1(men_men_n69_), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n48_), .B(x2), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n56_), .B0(x0), .Y(men_men_n76_));
  NA2        u060(.A(x5), .B(x3), .Y(men_men_n77_));
  NAi21      u061(.An(x4), .B(x3), .Y(men_men_n78_));
  INV        u062(.A(men_men_n78_), .Y(men_men_n79_));
  NO2        u063(.A(men_men_n79_), .B(men_men_n22_), .Y(men_men_n80_));
  NO2        u064(.A(x4), .B(x2), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n81_), .B(x3), .Y(men_men_n82_));
  NO3        u066(.A(men_men_n82_), .B(men_men_n80_), .C(men_men_n18_), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n83_), .B(men_men_n76_), .Y(men_men_n84_));
  NO4        u068(.A(men_men_n21_), .B(x6), .C(men_men_n43_), .D(x1), .Y(men_men_n85_));
  NA2        u069(.A(men_men_n62_), .B(men_men_n48_), .Y(men_men_n86_));
  INV        u070(.A(men_men_n86_), .Y(men_men_n87_));
  OAI210     u071(.A0(men_men_n85_), .A1(men_men_n65_), .B0(men_men_n87_), .Y(men_men_n88_));
  NA2        u072(.A(x3), .B(men_men_n18_), .Y(men_men_n89_));
  NO2        u073(.A(men_men_n89_), .B(men_men_n25_), .Y(men_men_n90_));
  INV        u074(.A(x8), .Y(men_men_n91_));
  NO2        u075(.A(x2), .B(men_men_n90_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n26_), .Y(men_men_n93_));
  AOI210     u077(.A0(men_men_n56_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n94_));
  OAI210     u078(.A0(men_men_n45_), .A1(men_men_n37_), .B0(men_men_n48_), .Y(men_men_n95_));
  NO3        u079(.A(men_men_n95_), .B(men_men_n94_), .C(men_men_n93_), .Y(men_men_n96_));
  NA2        u080(.A(x4), .B(men_men_n43_), .Y(men_men_n97_));
  NO2        u081(.A(men_men_n48_), .B(men_men_n54_), .Y(men_men_n98_));
  OAI210     u082(.A0(men_men_n98_), .A1(men_men_n43_), .B0(men_men_n18_), .Y(men_men_n99_));
  AOI210     u083(.A0(men_men_n97_), .A1(men_men_n52_), .B0(men_men_n99_), .Y(men_men_n100_));
  NO2        u084(.A(x3), .B(x2), .Y(men_men_n101_));
  NA2        u085(.A(men_men_n101_), .B(men_men_n25_), .Y(men_men_n102_));
  AOI210     u086(.A0(x8), .A1(x6), .B0(men_men_n102_), .Y(men_men_n103_));
  NA2        u087(.A(men_men_n54_), .B(x1), .Y(men_men_n104_));
  OAI210     u088(.A0(men_men_n104_), .A1(men_men_n40_), .B0(men_men_n17_), .Y(men_men_n105_));
  NO4        u089(.A(men_men_n105_), .B(men_men_n103_), .C(men_men_n100_), .D(men_men_n96_), .Y(men_men_n106_));
  AO220      u090(.A0(men_men_n106_), .A1(men_men_n88_), .B0(men_men_n84_), .B1(men_men_n74_), .Y(men02));
  NO2        u091(.A(x3), .B(men_men_n54_), .Y(men_men_n108_));
  NA2        u092(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n109_));
  NA2        u093(.A(men_men_n43_), .B(x0), .Y(men_men_n110_));
  OAI210     u094(.A0(men_men_n86_), .A1(men_men_n109_), .B0(men_men_n110_), .Y(men_men_n111_));
  NA2        u095(.A(men_men_n111_), .B(x1), .Y(men_men_n112_));
  NO3        u096(.A(men_men_n112_), .B(x7), .C(x5), .Y(men_men_n113_));
  NA2        u097(.A(x9), .B(x2), .Y(men_men_n114_));
  OR2        u098(.A(x8), .B(x0), .Y(men_men_n115_));
  INV        u099(.A(men_men_n115_), .Y(men_men_n116_));
  OAI210     u100(.A0(men_men_n114_), .A1(x7), .B0(men_men_n116_), .Y(men_men_n117_));
  NO2        u101(.A(x4), .B(x1), .Y(men_men_n118_));
  NA3        u102(.A(men_men_n118_), .B(men_men_n117_), .C(men_men_n60_), .Y(men_men_n119_));
  NOi21      u103(.An(x0), .B(x1), .Y(men_men_n120_));
  NO3        u104(.A(x9), .B(x8), .C(x7), .Y(men_men_n121_));
  NOi21      u105(.An(x0), .B(x4), .Y(men_men_n122_));
  NO2        u106(.A(x8), .B(men_men_n62_), .Y(men_men_n123_));
  AOI220     u107(.A0(men_men_n123_), .A1(men_men_n122_), .B0(men_men_n121_), .B1(men_men_n120_), .Y(men_men_n124_));
  AOI210     u108(.A0(men_men_n124_), .A1(men_men_n119_), .B0(men_men_n77_), .Y(men_men_n125_));
  NO2        u109(.A(x5), .B(men_men_n48_), .Y(men_men_n126_));
  NA2        u110(.A(x2), .B(men_men_n18_), .Y(men_men_n127_));
  NA2        u111(.A(men_men_n35_), .B(men_men_n126_), .Y(men_men_n128_));
  NAi21      u112(.An(x0), .B(x4), .Y(men_men_n129_));
  NO2        u113(.A(x7), .B(x0), .Y(men_men_n130_));
  NO2        u114(.A(men_men_n81_), .B(men_men_n98_), .Y(men_men_n131_));
  NO2        u115(.A(men_men_n21_), .B(men_men_n43_), .Y(men_men_n132_));
  NA2        u116(.A(x5), .B(x0), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n48_), .B(x2), .Y(men_men_n134_));
  NA3        u118(.A(men_men_n134_), .B(men_men_n133_), .C(men_men_n132_), .Y(men_men_n135_));
  NA3        u119(.A(men_men_n135_), .B(men_men_n128_), .C(men_men_n36_), .Y(men_men_n136_));
  NO3        u120(.A(men_men_n136_), .B(men_men_n125_), .C(men_men_n113_), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n138_));
  AOI220     u122(.A0(men_men_n120_), .A1(men_men_n138_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n139_));
  NO3        u123(.A(men_men_n139_), .B(men_men_n60_), .C(men_men_n62_), .Y(men_men_n140_));
  NA2        u124(.A(x7), .B(x3), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n97_), .B(x5), .Y(men_men_n142_));
  NO2        u126(.A(x9), .B(x7), .Y(men_men_n143_));
  NOi21      u127(.An(x8), .B(x0), .Y(men_men_n144_));
  OA210      u128(.A0(men_men_n143_), .A1(x1), .B0(men_men_n144_), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n43_), .B(x2), .Y(men_men_n146_));
  INV        u130(.A(x7), .Y(men_men_n147_));
  AOI220     u131(.A0(x1), .A1(men_men_n146_), .B0(men_men_n108_), .B1(men_men_n38_), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n25_), .B(x4), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n149_), .B(men_men_n122_), .Y(men_men_n150_));
  NO2        u134(.A(men_men_n150_), .B(men_men_n148_), .Y(men_men_n151_));
  AOI210     u135(.A0(men_men_n145_), .A1(men_men_n142_), .B0(men_men_n151_), .Y(men_men_n152_));
  OAI210     u136(.A0(men_men_n141_), .A1(men_men_n50_), .B0(men_men_n152_), .Y(men_men_n153_));
  NA2        u137(.A(x5), .B(x1), .Y(men_men_n154_));
  INV        u138(.A(men_men_n154_), .Y(men_men_n155_));
  AOI210     u139(.A0(men_men_n155_), .A1(men_men_n122_), .B0(men_men_n36_), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n62_), .B(men_men_n91_), .Y(men_men_n157_));
  NAi21      u141(.An(x2), .B(x7), .Y(men_men_n158_));
  NAi31      u142(.An(men_men_n77_), .B(men_men_n38_), .C(men_men_n35_), .Y(men_men_n159_));
  NA2        u143(.A(men_men_n159_), .B(men_men_n156_), .Y(men_men_n160_));
  NO3        u144(.A(men_men_n160_), .B(men_men_n153_), .C(men_men_n140_), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n161_), .B(men_men_n137_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n163_));
  NA2        u147(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n164_));
  NA2        u148(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n165_));
  NA3        u149(.A(men_men_n165_), .B(men_men_n164_), .C(men_men_n24_), .Y(men_men_n166_));
  AN2        u150(.A(men_men_n166_), .B(men_men_n134_), .Y(men_men_n167_));
  NA2        u151(.A(x8), .B(x0), .Y(men_men_n168_));
  NO2        u152(.A(men_men_n147_), .B(men_men_n25_), .Y(men_men_n169_));
  NO2        u153(.A(men_men_n120_), .B(x4), .Y(men_men_n170_));
  NA2        u154(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  AOI210     u155(.A0(men_men_n168_), .A1(men_men_n127_), .B0(men_men_n171_), .Y(men_men_n172_));
  NA2        u156(.A(x2), .B(x0), .Y(men_men_n173_));
  NA2        u157(.A(x4), .B(x1), .Y(men_men_n174_));
  NAi21      u158(.An(men_men_n118_), .B(men_men_n174_), .Y(men_men_n175_));
  NOi31      u159(.An(men_men_n175_), .B(men_men_n149_), .C(men_men_n173_), .Y(men_men_n176_));
  NO4        u160(.A(men_men_n176_), .B(men_men_n172_), .C(men_men_n167_), .D(men_men_n163_), .Y(men_men_n177_));
  NO2        u161(.A(men_men_n177_), .B(men_men_n43_), .Y(men_men_n178_));
  NO2        u162(.A(men_men_n166_), .B(men_men_n75_), .Y(men_men_n179_));
  INV        u163(.A(men_men_n126_), .Y(men_men_n180_));
  NO2        u164(.A(men_men_n104_), .B(men_men_n17_), .Y(men_men_n181_));
  AOI210     u165(.A0(men_men_n35_), .A1(men_men_n91_), .B0(men_men_n181_), .Y(men_men_n182_));
  NO3        u166(.A(men_men_n182_), .B(men_men_n180_), .C(x7), .Y(men_men_n183_));
  NA3        u167(.A(men_men_n175_), .B(men_men_n180_), .C(men_men_n42_), .Y(men_men_n184_));
  OAI210     u168(.A0(men_men_n165_), .A1(men_men_n131_), .B0(men_men_n184_), .Y(men_men_n185_));
  NO3        u169(.A(men_men_n185_), .B(men_men_n183_), .C(men_men_n179_), .Y(men_men_n186_));
  NO2        u170(.A(men_men_n186_), .B(x3), .Y(men_men_n187_));
  NO3        u171(.A(men_men_n187_), .B(men_men_n178_), .C(men_men_n162_), .Y(men03));
  NO2        u172(.A(men_men_n54_), .B(x1), .Y(men_men_n189_));
  OAI210     u173(.A0(men_men_n189_), .A1(men_men_n25_), .B0(x6), .Y(men_men_n190_));
  OAI220     u174(.A0(men_men_n190_), .A1(men_men_n17_), .B0(x6), .B1(men_men_n104_), .Y(men_men_n191_));
  NA2        u175(.A(men_men_n191_), .B(x4), .Y(men_men_n192_));
  NO2        u176(.A(men_men_n77_), .B(x6), .Y(men_men_n193_));
  NA2        u177(.A(x6), .B(men_men_n25_), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n194_), .B(x4), .Y(men_men_n195_));
  NO2        u179(.A(men_men_n18_), .B(x0), .Y(men_men_n196_));
  AO220      u180(.A0(men_men_n196_), .A1(men_men_n195_), .B0(men_men_n193_), .B1(men_men_n55_), .Y(men_men_n197_));
  NA2        u181(.A(men_men_n197_), .B(men_men_n62_), .Y(men_men_n198_));
  NA2        u182(.A(x3), .B(men_men_n17_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n199_), .B(men_men_n194_), .Y(men_men_n200_));
  AOI210     u184(.A0(men_men_n25_), .A1(x3), .B0(men_men_n173_), .Y(men_men_n201_));
  AOI220     u185(.A0(men_men_n201_), .A1(men_men_n25_), .B0(x9), .B1(men_men_n200_), .Y(men_men_n202_));
  NO3        u186(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n203_));
  NO2        u187(.A(x5), .B(x1), .Y(men_men_n204_));
  AOI220     u188(.A0(men_men_n204_), .A1(men_men_n17_), .B0(men_men_n101_), .B1(x5), .Y(men_men_n205_));
  NO2        u189(.A(men_men_n199_), .B(men_men_n164_), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n205_), .B(men_men_n36_), .Y(men_men_n207_));
  NA2        u191(.A(men_men_n207_), .B(men_men_n48_), .Y(men_men_n208_));
  NA4        u192(.A(men_men_n208_), .B(men_men_n202_), .C(men_men_n198_), .D(men_men_n192_), .Y(men_men_n209_));
  NO2        u193(.A(x3), .B(men_men_n17_), .Y(men_men_n210_));
  NO2        u194(.A(men_men_n210_), .B(x6), .Y(men_men_n211_));
  NOi21      u195(.An(men_men_n81_), .B(men_men_n211_), .Y(men_men_n212_));
  NA2        u196(.A(men_men_n62_), .B(men_men_n91_), .Y(men_men_n213_));
  NO2        u197(.A(men_men_n212_), .B(men_men_n147_), .Y(men_men_n214_));
  OR2        u198(.A(men_men_n214_), .B(men_men_n169_), .Y(men_men_n215_));
  NA2        u199(.A(men_men_n43_), .B(men_men_n54_), .Y(men_men_n216_));
  NO3        u200(.A(men_men_n174_), .B(men_men_n62_), .C(x6), .Y(men_men_n217_));
  AOI220     u201(.A0(men_men_n217_), .A1(men_men_n54_), .B0(men_men_n134_), .B1(men_men_n90_), .Y(men_men_n218_));
  NA2        u202(.A(x6), .B(men_men_n48_), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n154_), .B(men_men_n43_), .Y(men_men_n220_));
  NO2        u204(.A(men_men_n220_), .B(men_men_n206_), .Y(men_men_n221_));
  NA2        u205(.A(men_men_n126_), .B(x6), .Y(men_men_n222_));
  NA2        u206(.A(men_men_n222_), .B(men_men_n221_), .Y(men_men_n223_));
  NA2        u207(.A(men_men_n223_), .B(x2), .Y(men_men_n224_));
  NA3        u208(.A(men_men_n224_), .B(men_men_n218_), .C(men_men_n215_), .Y(men_men_n225_));
  AOI210     u209(.A0(men_men_n209_), .A1(x8), .B0(men_men_n225_), .Y(men_men_n226_));
  NO2        u210(.A(men_men_n91_), .B(x3), .Y(men_men_n227_));
  NA2        u211(.A(men_men_n227_), .B(men_men_n195_), .Y(men_men_n228_));
  INV        u212(.A(men_men_n228_), .Y(men_men_n229_));
  NO2        u213(.A(x4), .B(men_men_n54_), .Y(men_men_n230_));
  AOI220     u214(.A0(men_men_n195_), .A1(men_men_n181_), .B0(men_men_n230_), .B1(men_men_n65_), .Y(men_men_n231_));
  NA2        u215(.A(men_men_n62_), .B(x6), .Y(men_men_n232_));
  NA3        u216(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n233_));
  INV        u217(.A(men_men_n232_), .Y(men_men_n234_));
  NA2        u218(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n235_));
  NA2        u219(.A(men_men_n234_), .B(men_men_n118_), .Y(men_men_n236_));
  NO2        u220(.A(men_men_n199_), .B(x6), .Y(men_men_n237_));
  NA2        u221(.A(men_men_n157_), .B(men_men_n138_), .Y(men_men_n238_));
  NA4        u222(.A(men_men_n238_), .B(men_men_n236_), .C(men_men_n231_), .D(men_men_n147_), .Y(men_men_n239_));
  NO2        u223(.A(x9), .B(x6), .Y(men_men_n240_));
  NO2        u224(.A(men_men_n133_), .B(men_men_n18_), .Y(men_men_n241_));
  NAi21      u225(.An(men_men_n241_), .B(men_men_n233_), .Y(men_men_n242_));
  NAi21      u226(.An(x1), .B(x4), .Y(men_men_n243_));
  AOI210     u227(.A0(x3), .A1(x2), .B0(men_men_n48_), .Y(men_men_n244_));
  OAI210     u228(.A0(men_men_n133_), .A1(x3), .B0(men_men_n244_), .Y(men_men_n245_));
  AOI220     u229(.A0(men_men_n245_), .A1(men_men_n243_), .B0(men_men_n242_), .B1(men_men_n240_), .Y(men_men_n246_));
  INV        u230(.A(men_men_n246_), .Y(men_men_n247_));
  NA2        u231(.A(men_men_n62_), .B(x2), .Y(men_men_n248_));
  NO2        u232(.A(men_men_n248_), .B(x3), .Y(men_men_n249_));
  NO3        u233(.A(x9), .B(x6), .C(x0), .Y(men_men_n250_));
  NA2        u234(.A(x6), .B(x2), .Y(men_men_n251_));
  NO2        u235(.A(men_men_n251_), .B(men_men_n164_), .Y(men_men_n252_));
  NO2        u236(.A(men_men_n250_), .B(men_men_n252_), .Y(men_men_n253_));
  OAI220     u237(.A0(men_men_n253_), .A1(men_men_n43_), .B0(men_men_n170_), .B1(men_men_n46_), .Y(men_men_n254_));
  OAI210     u238(.A0(men_men_n254_), .A1(men_men_n249_), .B0(men_men_n247_), .Y(men_men_n255_));
  NO2        u239(.A(men_men_n426_), .B(men_men_n194_), .Y(men_men_n256_));
  OR3        u240(.A(men_men_n256_), .B(men_men_n193_), .C(men_men_n142_), .Y(men_men_n257_));
  NA2        u241(.A(x4), .B(x0), .Y(men_men_n258_));
  NO3        u242(.A(men_men_n72_), .B(men_men_n258_), .C(x6), .Y(men_men_n259_));
  AOI210     u243(.A0(men_men_n257_), .A1(men_men_n42_), .B0(men_men_n259_), .Y(men_men_n260_));
  AOI210     u244(.A0(men_men_n260_), .A1(men_men_n255_), .B0(x8), .Y(men_men_n261_));
  INV        u245(.A(men_men_n232_), .Y(men_men_n262_));
  OAI210     u246(.A0(men_men_n241_), .A1(men_men_n204_), .B0(men_men_n262_), .Y(men_men_n263_));
  INV        u247(.A(men_men_n168_), .Y(men_men_n264_));
  OAI210     u248(.A0(men_men_n264_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n265_));
  AOI210     u249(.A0(men_men_n265_), .A1(men_men_n263_), .B0(men_men_n216_), .Y(men_men_n266_));
  NO4        u250(.A(men_men_n266_), .B(men_men_n261_), .C(men_men_n239_), .D(men_men_n229_), .Y(men_men_n267_));
  NO2        u251(.A(men_men_n157_), .B(x1), .Y(men_men_n268_));
  NO3        u252(.A(men_men_n268_), .B(x3), .C(men_men_n36_), .Y(men_men_n269_));
  OAI210     u253(.A0(men_men_n269_), .A1(men_men_n237_), .B0(x2), .Y(men_men_n270_));
  OAI210     u254(.A0(men_men_n264_), .A1(x6), .B0(men_men_n44_), .Y(men_men_n271_));
  AOI210     u255(.A0(men_men_n271_), .A1(men_men_n270_), .B0(men_men_n180_), .Y(men_men_n272_));
  NOi21      u256(.An(men_men_n251_), .B(men_men_n17_), .Y(men_men_n273_));
  NA3        u257(.A(men_men_n273_), .B(men_men_n204_), .C(men_men_n40_), .Y(men_men_n274_));
  AOI210     u258(.A0(men_men_n36_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n275_));
  NA3        u259(.A(men_men_n275_), .B(men_men_n155_), .C(men_men_n32_), .Y(men_men_n276_));
  NA2        u260(.A(x3), .B(x2), .Y(men_men_n277_));
  AOI220     u261(.A0(men_men_n277_), .A1(men_men_n216_), .B0(men_men_n276_), .B1(men_men_n274_), .Y(men_men_n278_));
  NAi21      u262(.An(x4), .B(x0), .Y(men_men_n279_));
  NO3        u263(.A(men_men_n279_), .B(men_men_n44_), .C(x2), .Y(men_men_n280_));
  OAI210     u264(.A0(x6), .A1(men_men_n18_), .B0(men_men_n280_), .Y(men_men_n281_));
  OAI220     u265(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n282_));
  NO2        u266(.A(x9), .B(x8), .Y(men_men_n283_));
  NA2        u267(.A(men_men_n36_), .B(men_men_n54_), .Y(men_men_n284_));
  OAI210     u268(.A0(men_men_n275_), .A1(men_men_n273_), .B0(men_men_n284_), .Y(men_men_n285_));
  AOI220     u269(.A0(men_men_n285_), .A1(men_men_n79_), .B0(men_men_n282_), .B1(men_men_n31_), .Y(men_men_n286_));
  AOI210     u270(.A0(men_men_n286_), .A1(men_men_n281_), .B0(men_men_n25_), .Y(men_men_n287_));
  NA3        u271(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n288_));
  OAI210     u272(.A0(men_men_n275_), .A1(men_men_n273_), .B0(men_men_n288_), .Y(men_men_n289_));
  NA2        u273(.A(men_men_n36_), .B(men_men_n43_), .Y(men_men_n290_));
  OR2        u274(.A(men_men_n290_), .B(men_men_n258_), .Y(men_men_n291_));
  NO2        u275(.A(men_men_n291_), .B(men_men_n154_), .Y(men_men_n292_));
  AO210      u276(.A0(men_men_n289_), .A1(men_men_n142_), .B0(men_men_n292_), .Y(men_men_n293_));
  NO4        u277(.A(men_men_n293_), .B(men_men_n287_), .C(men_men_n278_), .D(men_men_n272_), .Y(men_men_n294_));
  OAI210     u278(.A0(men_men_n267_), .A1(men_men_n226_), .B0(men_men_n294_), .Y(men04));
  OAI210     u279(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n296_));
  NA3        u280(.A(men_men_n296_), .B(men_men_n250_), .C(men_men_n82_), .Y(men_men_n297_));
  NO2        u281(.A(x2), .B(x1), .Y(men_men_n298_));
  OAI210     u282(.A0(men_men_n235_), .A1(men_men_n298_), .B0(men_men_n36_), .Y(men_men_n299_));
  NO2        u283(.A(men_men_n298_), .B(men_men_n279_), .Y(men_men_n300_));
  AOI210     u284(.A0(men_men_n62_), .A1(x4), .B0(men_men_n109_), .Y(men_men_n301_));
  OAI210     u285(.A0(men_men_n301_), .A1(men_men_n300_), .B0(men_men_n227_), .Y(men_men_n302_));
  NO2        u286(.A(men_men_n248_), .B(men_men_n89_), .Y(men_men_n303_));
  NO2        u287(.A(men_men_n303_), .B(men_men_n36_), .Y(men_men_n304_));
  NO2        u288(.A(men_men_n277_), .B(men_men_n196_), .Y(men_men_n305_));
  NA2        u289(.A(x9), .B(x0), .Y(men_men_n306_));
  AOI210     u290(.A0(men_men_n89_), .A1(men_men_n75_), .B0(men_men_n306_), .Y(men_men_n307_));
  OAI210     u291(.A0(men_men_n307_), .A1(men_men_n305_), .B0(men_men_n91_), .Y(men_men_n308_));
  NA3        u292(.A(men_men_n308_), .B(men_men_n304_), .C(men_men_n302_), .Y(men_men_n309_));
  NA2        u293(.A(men_men_n309_), .B(men_men_n299_), .Y(men_men_n310_));
  NO3        u294(.A(men_men_n232_), .B(x2), .C(men_men_n18_), .Y(men_men_n311_));
  INV        u295(.A(men_men_n311_), .Y(men_men_n312_));
  OAI210     u296(.A0(men_men_n115_), .A1(men_men_n104_), .B0(men_men_n168_), .Y(men_men_n313_));
  NA3        u297(.A(men_men_n313_), .B(x6), .C(x3), .Y(men_men_n314_));
  NOi21      u298(.An(men_men_n144_), .B(men_men_n127_), .Y(men_men_n315_));
  AOI210     u299(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n316_));
  OAI220     u300(.A0(men_men_n316_), .A1(men_men_n290_), .B0(men_men_n248_), .B1(men_men_n288_), .Y(men_men_n317_));
  AOI210     u301(.A0(men_men_n315_), .A1(x6), .B0(men_men_n317_), .Y(men_men_n318_));
  NO2        u302(.A(men_men_n104_), .B(men_men_n17_), .Y(men_men_n319_));
  AOI210     u303(.A0(men_men_n303_), .A1(men_men_n91_), .B0(men_men_n319_), .Y(men_men_n320_));
  NA4        u304(.A(men_men_n320_), .B(men_men_n318_), .C(men_men_n314_), .D(men_men_n312_), .Y(men_men_n321_));
  OAI210     u305(.A0(x1), .A1(x3), .B0(men_men_n280_), .Y(men_men_n322_));
  NA3        u306(.A(men_men_n213_), .B(men_men_n203_), .C(men_men_n81_), .Y(men_men_n323_));
  NA3        u307(.A(men_men_n323_), .B(men_men_n322_), .C(men_men_n147_), .Y(men_men_n324_));
  AOI210     u308(.A0(men_men_n321_), .A1(x4), .B0(men_men_n324_), .Y(men_men_n325_));
  NA2        u309(.A(men_men_n300_), .B(men_men_n91_), .Y(men_men_n326_));
  NOi21      u310(.An(x4), .B(x0), .Y(men_men_n327_));
  XO2        u311(.A(x4), .B(x0), .Y(men_men_n328_));
  OAI210     u312(.A0(men_men_n328_), .A1(men_men_n114_), .B0(men_men_n243_), .Y(men_men_n329_));
  NA2        u313(.A(men_men_n329_), .B(x8), .Y(men_men_n330_));
  AOI210     u314(.A0(men_men_n330_), .A1(men_men_n326_), .B0(x3), .Y(men_men_n331_));
  NO2        u315(.A(men_men_n91_), .B(x4), .Y(men_men_n332_));
  NA2        u316(.A(men_men_n332_), .B(men_men_n44_), .Y(men_men_n333_));
  NO3        u317(.A(men_men_n328_), .B(men_men_n157_), .C(x2), .Y(men_men_n334_));
  NO2        u318(.A(men_men_n28_), .B(men_men_n24_), .Y(men_men_n335_));
  NO2        u319(.A(men_men_n335_), .B(men_men_n334_), .Y(men_men_n336_));
  NA3        u320(.A(men_men_n336_), .B(men_men_n333_), .C(x6), .Y(men_men_n337_));
  OAI220     u321(.A0(men_men_n279_), .A1(men_men_n89_), .B0(men_men_n173_), .B1(men_men_n91_), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n144_), .B(men_men_n104_), .Y(men_men_n339_));
  NO2        u323(.A(men_men_n338_), .B(men_men_n339_), .Y(men_men_n340_));
  NO2        u324(.A(men_men_n144_), .B(men_men_n78_), .Y(men_men_n341_));
  NO2        u325(.A(men_men_n340_), .B(men_men_n62_), .Y(men_men_n342_));
  OAI220     u326(.A0(men_men_n342_), .A1(x6), .B0(men_men_n337_), .B1(men_men_n331_), .Y(men_men_n343_));
  OAI210     u327(.A0(x6), .A1(men_men_n48_), .B0(men_men_n42_), .Y(men_men_n344_));
  OAI210     u328(.A0(men_men_n344_), .A1(men_men_n91_), .B0(men_men_n291_), .Y(men_men_n345_));
  AOI210     u329(.A0(men_men_n345_), .A1(men_men_n18_), .B0(men_men_n147_), .Y(men_men_n346_));
  AO220      u330(.A0(men_men_n346_), .A1(men_men_n343_), .B0(men_men_n325_), .B1(men_men_n310_), .Y(men_men_n347_));
  AOI210     u331(.A0(x6), .A1(x1), .B0(men_men_n146_), .Y(men_men_n348_));
  NA2        u332(.A(men_men_n332_), .B(x0), .Y(men_men_n349_));
  NO2        u333(.A(men_men_n349_), .B(men_men_n348_), .Y(men_men_n350_));
  INV        u334(.A(men_men_n350_), .Y(men_men_n351_));
  NA3        u335(.A(men_men_n351_), .B(men_men_n347_), .C(men_men_n297_), .Y(men_men_n352_));
  AO220      u336(.A0(x4), .A1(men_men_n143_), .B0(men_men_n108_), .B1(x4), .Y(men_men_n353_));
  NA2        u337(.A(x3), .B(x0), .Y(men_men_n354_));
  NO2        u338(.A(men_men_n354_), .B(x2), .Y(men_men_n355_));
  AOI210     u339(.A0(men_men_n353_), .A1(men_men_n116_), .B0(men_men_n355_), .Y(men_men_n356_));
  NO2        u340(.A(men_men_n356_), .B(men_men_n25_), .Y(men_men_n357_));
  OAI210     u341(.A0(x4), .A1(men_men_n66_), .B0(men_men_n196_), .Y(men_men_n358_));
  NA3        u342(.A(men_men_n189_), .B(men_men_n210_), .C(x8), .Y(men_men_n359_));
  AOI210     u343(.A0(men_men_n359_), .A1(men_men_n358_), .B0(men_men_n25_), .Y(men_men_n360_));
  AOI210     u344(.A0(x2), .A1(men_men_n115_), .B0(men_men_n42_), .Y(men_men_n361_));
  NOi31      u345(.An(men_men_n361_), .B(x3), .C(men_men_n174_), .Y(men_men_n362_));
  OAI210     u346(.A0(men_men_n362_), .A1(men_men_n360_), .B0(men_men_n143_), .Y(men_men_n363_));
  NAi31      u347(.An(men_men_n50_), .B(men_men_n268_), .C(men_men_n169_), .Y(men_men_n364_));
  NA2        u348(.A(men_men_n364_), .B(men_men_n363_), .Y(men_men_n365_));
  OAI210     u349(.A0(men_men_n365_), .A1(men_men_n357_), .B0(x6), .Y(men_men_n366_));
  OAI210     u350(.A0(men_men_n157_), .A1(men_men_n48_), .B0(men_men_n130_), .Y(men_men_n367_));
  NA3        u351(.A(men_men_n55_), .B(men_men_n38_), .C(men_men_n31_), .Y(men_men_n368_));
  AOI220     u352(.A0(men_men_n368_), .A1(men_men_n367_), .B0(men_men_n40_), .B1(men_men_n32_), .Y(men_men_n369_));
  AOI210     u353(.A0(men_men_n123_), .A1(men_men_n230_), .B0(x1), .Y(men_men_n370_));
  INV        u354(.A(men_men_n370_), .Y(men_men_n371_));
  NAi31      u355(.An(x2), .B(x8), .C(x0), .Y(men_men_n372_));
  OAI210     u356(.A0(men_men_n372_), .A1(x4), .B0(men_men_n158_), .Y(men_men_n373_));
  NA3        u357(.A(men_men_n373_), .B(men_men_n141_), .C(x9), .Y(men_men_n374_));
  NO4        u358(.A(x8), .B(men_men_n279_), .C(x9), .D(x2), .Y(men_men_n375_));
  NOi21      u359(.An(men_men_n121_), .B(men_men_n173_), .Y(men_men_n376_));
  NO3        u360(.A(men_men_n376_), .B(men_men_n375_), .C(men_men_n18_), .Y(men_men_n377_));
  NO3        u361(.A(x9), .B(men_men_n147_), .C(x0), .Y(men_men_n378_));
  AOI220     u362(.A0(men_men_n378_), .A1(men_men_n227_), .B0(men_men_n341_), .B1(men_men_n147_), .Y(men_men_n379_));
  NA4        u363(.A(men_men_n379_), .B(men_men_n377_), .C(men_men_n374_), .D(men_men_n50_), .Y(men_men_n380_));
  OAI210     u364(.A0(men_men_n371_), .A1(men_men_n369_), .B0(men_men_n380_), .Y(men_men_n381_));
  AOI210     u365(.A0(men_men_n38_), .A1(x9), .B0(men_men_n129_), .Y(men_men_n382_));
  NO3        u366(.A(men_men_n382_), .B(men_men_n121_), .C(men_men_n43_), .Y(men_men_n383_));
  NOi31      u367(.An(x1), .B(x8), .C(x7), .Y(men_men_n384_));
  AOI220     u368(.A0(men_men_n384_), .A1(men_men_n327_), .B0(men_men_n122_), .B1(x3), .Y(men_men_n385_));
  AOI210     u369(.A0(men_men_n243_), .A1(men_men_n60_), .B0(men_men_n120_), .Y(men_men_n386_));
  OAI210     u370(.A0(men_men_n386_), .A1(x3), .B0(men_men_n385_), .Y(men_men_n387_));
  NO3        u371(.A(men_men_n387_), .B(men_men_n383_), .C(x2), .Y(men_men_n388_));
  OAI220     u372(.A0(men_men_n328_), .A1(men_men_n283_), .B0(men_men_n279_), .B1(men_men_n43_), .Y(men_men_n389_));
  NA2        u373(.A(men_men_n389_), .B(men_men_n147_), .Y(men_men_n390_));
  NO2        u374(.A(men_men_n390_), .B(men_men_n54_), .Y(men_men_n391_));
  NO2        u375(.A(men_men_n391_), .B(men_men_n388_), .Y(men_men_n392_));
  AOI210     u376(.A0(men_men_n392_), .A1(men_men_n381_), .B0(men_men_n25_), .Y(men_men_n393_));
  NA4        u377(.A(men_men_n31_), .B(men_men_n91_), .C(x2), .D(men_men_n17_), .Y(men_men_n394_));
  NO3        u378(.A(men_men_n62_), .B(x4), .C(x1), .Y(men_men_n395_));
  AOI220     u379(.A0(x1), .A1(men_men_n244_), .B0(men_men_n395_), .B1(men_men_n361_), .Y(men_men_n396_));
  NO2        u380(.A(men_men_n396_), .B(men_men_n101_), .Y(men_men_n397_));
  NO3        u381(.A(men_men_n248_), .B(men_men_n168_), .C(men_men_n40_), .Y(men_men_n398_));
  OAI210     u382(.A0(men_men_n398_), .A1(men_men_n397_), .B0(x7), .Y(men_men_n399_));
  NA2        u383(.A(men_men_n399_), .B(men_men_n394_), .Y(men_men_n400_));
  OAI210     u384(.A0(men_men_n400_), .A1(men_men_n393_), .B0(men_men_n36_), .Y(men_men_n401_));
  NO2        u385(.A(men_men_n378_), .B(men_men_n196_), .Y(men_men_n402_));
  NO4        u386(.A(men_men_n402_), .B(men_men_n77_), .C(x4), .D(men_men_n54_), .Y(men_men_n403_));
  NA2        u387(.A(men_men_n235_), .B(men_men_n21_), .Y(men_men_n404_));
  NO2        u388(.A(men_men_n154_), .B(men_men_n130_), .Y(men_men_n405_));
  NA2        u389(.A(men_men_n405_), .B(men_men_n404_), .Y(men_men_n406_));
  AOI210     u390(.A0(men_men_n406_), .A1(men_men_n159_), .B0(men_men_n28_), .Y(men_men_n407_));
  AOI220     u391(.A0(x3), .A1(men_men_n91_), .B0(men_men_n144_), .B1(men_men_n189_), .Y(men_men_n408_));
  NA3        u392(.A(men_men_n408_), .B(men_men_n372_), .C(men_men_n89_), .Y(men_men_n409_));
  NA2        u393(.A(men_men_n409_), .B(men_men_n169_), .Y(men_men_n410_));
  OAI220     u394(.A0(men_men_n426_), .A1(men_men_n67_), .B0(men_men_n154_), .B1(men_men_n43_), .Y(men_men_n411_));
  AOI210     u395(.A0(men_men_n158_), .A1(men_men_n27_), .B0(men_men_n72_), .Y(men_men_n412_));
  OAI210     u396(.A0(men_men_n143_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n413_));
  NO3        u397(.A(men_men_n384_), .B(x3), .C(men_men_n54_), .Y(men_men_n414_));
  AOI210     u398(.A0(men_men_n414_), .A1(men_men_n413_), .B0(men_men_n412_), .Y(men_men_n415_));
  INV        u399(.A(men_men_n415_), .Y(men_men_n416_));
  AOI220     u400(.A0(men_men_n416_), .A1(x0), .B0(men_men_n411_), .B1(men_men_n130_), .Y(men_men_n417_));
  AOI210     u401(.A0(men_men_n417_), .A1(men_men_n410_), .B0(men_men_n219_), .Y(men_men_n418_));
  NA2        u402(.A(x9), .B(x5), .Y(men_men_n419_));
  NO4        u403(.A(men_men_n104_), .B(men_men_n419_), .C(men_men_n60_), .D(men_men_n32_), .Y(men_men_n420_));
  NO4        u404(.A(men_men_n420_), .B(men_men_n418_), .C(men_men_n407_), .D(men_men_n403_), .Y(men_men_n421_));
  NA3        u405(.A(men_men_n421_), .B(men_men_n401_), .C(men_men_n366_), .Y(men_men_n422_));
  AOI210     u406(.A0(men_men_n352_), .A1(men_men_n25_), .B0(men_men_n422_), .Y(men05));
  INV        u407(.A(x9), .Y(men_men_n426_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule