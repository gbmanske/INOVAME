//Benchmark atmr_max1024_476_0.125

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n354_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n462_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  INV        o005(.A(ori_ori_n19_), .Y(ori_ori_n22_));
  NA2        o006(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n23_));
  INV        o007(.A(x5), .Y(ori_ori_n24_));
  NA2        o008(.A(x7), .B(x6), .Y(ori_ori_n25_));
  NA2        o009(.A(x4), .B(x2), .Y(ori_ori_n26_));
  INV        o010(.A(ori_ori_n23_), .Y(ori_ori_n27_));
  NO2        o011(.A(x4), .B(x3), .Y(ori_ori_n28_));
  INV        o012(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  NOi21      o013(.An(ori_ori_n22_), .B(ori_ori_n27_), .Y(ori00));
  NO2        o014(.A(x1), .B(x0), .Y(ori_ori_n31_));
  INV        o015(.A(x6), .Y(ori_ori_n32_));
  NO2        o016(.A(ori_ori_n32_), .B(ori_ori_n24_), .Y(ori_ori_n33_));
  NA2        o017(.A(x4), .B(x3), .Y(ori_ori_n34_));
  NO2        o018(.A(ori_ori_n22_), .B(ori_ori_n34_), .Y(ori_ori_n35_));
  NO2        o019(.A(x2), .B(x0), .Y(ori_ori_n36_));
  INV        o020(.A(x3), .Y(ori_ori_n37_));
  NO2        o021(.A(ori_ori_n37_), .B(ori_ori_n18_), .Y(ori_ori_n38_));
  INV        o022(.A(ori_ori_n38_), .Y(ori_ori_n39_));
  NO2        o023(.A(ori_ori_n33_), .B(x4), .Y(ori_ori_n40_));
  OAI210     o024(.A0(ori_ori_n40_), .A1(ori_ori_n39_), .B0(ori_ori_n36_), .Y(ori_ori_n41_));
  INV        o025(.A(x4), .Y(ori_ori_n42_));
  NO2        o026(.A(ori_ori_n42_), .B(ori_ori_n17_), .Y(ori_ori_n43_));
  NA2        o027(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n44_));
  OAI210     o028(.A0(ori_ori_n44_), .A1(ori_ori_n20_), .B0(ori_ori_n41_), .Y(ori_ori_n45_));
  INV        o029(.A(ori_ori_n31_), .Y(ori_ori_n46_));
  INV        o030(.A(x2), .Y(ori_ori_n47_));
  NO2        o031(.A(ori_ori_n47_), .B(ori_ori_n17_), .Y(ori_ori_n48_));
  NA2        o032(.A(ori_ori_n37_), .B(ori_ori_n18_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(ori_ori_n48_), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n46_), .A1(ori_ori_n29_), .B0(ori_ori_n50_), .Y(ori_ori_n51_));
  NO3        o035(.A(ori_ori_n51_), .B(ori_ori_n45_), .C(ori_ori_n35_), .Y(ori01));
  NA2        o036(.A(x8), .B(x7), .Y(ori_ori_n53_));
  NA2        o037(.A(ori_ori_n37_), .B(x1), .Y(ori_ori_n54_));
  NO2        o038(.A(x7), .B(x6), .Y(ori_ori_n55_));
  NO2        o039(.A(ori_ori_n54_), .B(x5), .Y(ori_ori_n56_));
  NO2        o040(.A(x8), .B(x2), .Y(ori_ori_n57_));
  INV        o041(.A(ori_ori_n57_), .Y(ori_ori_n58_));
  OAI210     o042(.A0(ori_ori_n38_), .A1(ori_ori_n24_), .B0(ori_ori_n47_), .Y(ori_ori_n59_));
  OAI210     o043(.A0(ori_ori_n49_), .A1(ori_ori_n20_), .B0(ori_ori_n59_), .Y(ori_ori_n60_));
  INV        o044(.A(ori_ori_n60_), .Y(ori_ori_n61_));
  NA2        o045(.A(ori_ori_n61_), .B(x4), .Y(ori_ori_n62_));
  NA2        o046(.A(ori_ori_n42_), .B(x2), .Y(ori_ori_n63_));
  OAI210     o047(.A0(ori_ori_n63_), .A1(ori_ori_n49_), .B0(x0), .Y(ori_ori_n64_));
  NA2        o048(.A(x5), .B(x3), .Y(ori_ori_n65_));
  NO2        o049(.A(x8), .B(x6), .Y(ori_ori_n66_));
  NO4        o050(.A(ori_ori_n66_), .B(ori_ori_n65_), .C(ori_ori_n55_), .D(ori_ori_n47_), .Y(ori_ori_n67_));
  NAi21      o051(.An(x4), .B(x3), .Y(ori_ori_n68_));
  INV        o052(.A(ori_ori_n68_), .Y(ori_ori_n69_));
  NO2        o053(.A(x4), .B(x2), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n68_), .B(ori_ori_n18_), .Y(ori_ori_n71_));
  NO3        o055(.A(ori_ori_n71_), .B(ori_ori_n67_), .C(ori_ori_n64_), .Y(ori_ori_n72_));
  NA2        o056(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n73_), .B(ori_ori_n24_), .Y(ori_ori_n74_));
  INV        o058(.A(x8), .Y(ori_ori_n75_));
  NA2        o059(.A(x2), .B(x1), .Y(ori_ori_n76_));
  INV        o060(.A(ori_ori_n74_), .Y(ori_ori_n77_));
  NO2        o061(.A(ori_ori_n77_), .B(ori_ori_n25_), .Y(ori_ori_n78_));
  AOI210     o062(.A0(ori_ori_n49_), .A1(ori_ori_n24_), .B0(ori_ori_n47_), .Y(ori_ori_n79_));
  OAI210     o063(.A0(ori_ori_n39_), .A1(ori_ori_n33_), .B0(ori_ori_n42_), .Y(ori_ori_n80_));
  NO3        o064(.A(ori_ori_n80_), .B(ori_ori_n79_), .C(ori_ori_n78_), .Y(ori_ori_n81_));
  NA2        o065(.A(x4), .B(ori_ori_n37_), .Y(ori_ori_n82_));
  NO2        o066(.A(ori_ori_n42_), .B(ori_ori_n47_), .Y(ori_ori_n83_));
  NO2        o067(.A(ori_ori_n82_), .B(x1), .Y(ori_ori_n84_));
  NO2        o068(.A(x3), .B(x2), .Y(ori_ori_n85_));
  NA3        o069(.A(ori_ori_n85_), .B(ori_ori_n25_), .C(ori_ori_n24_), .Y(ori_ori_n86_));
  INV        o070(.A(ori_ori_n86_), .Y(ori_ori_n87_));
  NA2        o071(.A(ori_ori_n47_), .B(x1), .Y(ori_ori_n88_));
  OAI210     o072(.A0(ori_ori_n88_), .A1(ori_ori_n34_), .B0(ori_ori_n17_), .Y(ori_ori_n89_));
  NO4        o073(.A(ori_ori_n89_), .B(ori_ori_n87_), .C(ori_ori_n84_), .D(ori_ori_n81_), .Y(ori_ori_n90_));
  AO210      o074(.A0(ori_ori_n72_), .A1(ori_ori_n62_), .B0(ori_ori_n90_), .Y(ori02));
  NO2        o075(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n92_));
  NA2        o076(.A(ori_ori_n37_), .B(x0), .Y(ori_ori_n93_));
  BUFFER     o077(.A(x0), .Y(ori_ori_n94_));
  INV        o078(.A(ori_ori_n94_), .Y(ori_ori_n95_));
  NO2        o079(.A(x4), .B(x1), .Y(ori_ori_n96_));
  NA2        o080(.A(ori_ori_n96_), .B(x2), .Y(ori_ori_n97_));
  NOi21      o081(.An(x0), .B(x1), .Y(ori_ori_n98_));
  NOi21      o082(.An(x0), .B(x4), .Y(ori_ori_n99_));
  NO2        o083(.A(ori_ori_n97_), .B(ori_ori_n65_), .Y(ori_ori_n100_));
  NO2        o084(.A(x5), .B(ori_ori_n42_), .Y(ori_ori_n101_));
  NA2        o085(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n102_));
  AOI210     o086(.A0(ori_ori_n102_), .A1(ori_ori_n88_), .B0(ori_ori_n93_), .Y(ori_ori_n103_));
  OAI210     o087(.A0(ori_ori_n103_), .A1(ori_ori_n31_), .B0(ori_ori_n101_), .Y(ori_ori_n104_));
  NAi21      o088(.An(x0), .B(x4), .Y(ori_ori_n105_));
  NO2        o089(.A(ori_ori_n105_), .B(x1), .Y(ori_ori_n106_));
  NO2        o090(.A(x7), .B(x0), .Y(ori_ori_n107_));
  NO2        o091(.A(ori_ori_n70_), .B(ori_ori_n83_), .Y(ori_ori_n108_));
  NO2        o092(.A(ori_ori_n108_), .B(x3), .Y(ori_ori_n109_));
  OAI210     o093(.A0(ori_ori_n107_), .A1(ori_ori_n106_), .B0(ori_ori_n109_), .Y(ori_ori_n110_));
  NA2        o094(.A(x5), .B(x0), .Y(ori_ori_n111_));
  NO2        o095(.A(ori_ori_n42_), .B(x2), .Y(ori_ori_n112_));
  NA3        o096(.A(ori_ori_n110_), .B(ori_ori_n104_), .C(ori_ori_n32_), .Y(ori_ori_n113_));
  NO2        o097(.A(ori_ori_n113_), .B(ori_ori_n100_), .Y(ori_ori_n114_));
  NO3        o098(.A(ori_ori_n65_), .B(ori_ori_n63_), .C(ori_ori_n23_), .Y(ori_ori_n115_));
  NO2        o099(.A(ori_ori_n26_), .B(ori_ori_n24_), .Y(ori_ori_n116_));
  NA2        o100(.A(x7), .B(x3), .Y(ori_ori_n117_));
  NO2        o101(.A(ori_ori_n82_), .B(x5), .Y(ori_ori_n118_));
  NO2        o102(.A(ori_ori_n37_), .B(x2), .Y(ori_ori_n119_));
  INV        o103(.A(x7), .Y(ori_ori_n120_));
  NA2        o104(.A(ori_ori_n120_), .B(ori_ori_n18_), .Y(ori_ori_n121_));
  NA2        o105(.A(ori_ori_n121_), .B(ori_ori_n119_), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n24_), .B(x4), .Y(ori_ori_n123_));
  NO2        o107(.A(ori_ori_n123_), .B(ori_ori_n99_), .Y(ori_ori_n124_));
  NO2        o108(.A(ori_ori_n124_), .B(ori_ori_n122_), .Y(ori_ori_n125_));
  INV        o109(.A(ori_ori_n125_), .Y(ori_ori_n126_));
  OAI210     o110(.A0(ori_ori_n117_), .A1(ori_ori_n44_), .B0(ori_ori_n126_), .Y(ori_ori_n127_));
  NA2        o111(.A(x5), .B(x1), .Y(ori_ori_n128_));
  INV        o112(.A(ori_ori_n128_), .Y(ori_ori_n129_));
  AOI210     o113(.A0(ori_ori_n129_), .A1(ori_ori_n99_), .B0(ori_ori_n32_), .Y(ori_ori_n130_));
  NAi21      o114(.An(x2), .B(x7), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n131_), .B(ori_ori_n42_), .Y(ori_ori_n132_));
  NA2        o116(.A(ori_ori_n132_), .B(ori_ori_n56_), .Y(ori_ori_n133_));
  NA2        o117(.A(ori_ori_n133_), .B(ori_ori_n130_), .Y(ori_ori_n134_));
  NO3        o118(.A(ori_ori_n134_), .B(ori_ori_n127_), .C(ori_ori_n115_), .Y(ori_ori_n135_));
  NO2        o119(.A(ori_ori_n135_), .B(ori_ori_n114_), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n111_), .B(ori_ori_n108_), .Y(ori_ori_n137_));
  NA2        o121(.A(ori_ori_n24_), .B(ori_ori_n18_), .Y(ori_ori_n138_));
  NA2        o122(.A(ori_ori_n24_), .B(ori_ori_n17_), .Y(ori_ori_n139_));
  NA3        o123(.A(ori_ori_n139_), .B(ori_ori_n138_), .C(ori_ori_n23_), .Y(ori_ori_n140_));
  AN2        o124(.A(ori_ori_n140_), .B(ori_ori_n112_), .Y(ori_ori_n141_));
  NA2        o125(.A(x8), .B(x0), .Y(ori_ori_n142_));
  NO2        o126(.A(ori_ori_n120_), .B(ori_ori_n24_), .Y(ori_ori_n143_));
  NA2        o127(.A(x2), .B(x0), .Y(ori_ori_n144_));
  NA2        o128(.A(x4), .B(x1), .Y(ori_ori_n145_));
  NAi21      o129(.An(ori_ori_n96_), .B(ori_ori_n145_), .Y(ori_ori_n146_));
  NOi31      o130(.An(ori_ori_n146_), .B(ori_ori_n123_), .C(ori_ori_n144_), .Y(ori_ori_n147_));
  NO3        o131(.A(ori_ori_n147_), .B(ori_ori_n141_), .C(ori_ori_n137_), .Y(ori_ori_n148_));
  NO2        o132(.A(ori_ori_n148_), .B(ori_ori_n37_), .Y(ori_ori_n149_));
  NO2        o133(.A(ori_ori_n140_), .B(ori_ori_n63_), .Y(ori_ori_n150_));
  INV        o134(.A(ori_ori_n101_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n88_), .B(ori_ori_n17_), .Y(ori_ori_n152_));
  AOI210     o136(.A0(ori_ori_n31_), .A1(ori_ori_n75_), .B0(ori_ori_n152_), .Y(ori_ori_n153_));
  NO3        o137(.A(ori_ori_n153_), .B(ori_ori_n151_), .C(x7), .Y(ori_ori_n154_));
  NA3        o138(.A(ori_ori_n146_), .B(ori_ori_n151_), .C(ori_ori_n36_), .Y(ori_ori_n155_));
  OAI210     o139(.A0(ori_ori_n139_), .A1(ori_ori_n108_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NO3        o140(.A(ori_ori_n156_), .B(ori_ori_n154_), .C(ori_ori_n150_), .Y(ori_ori_n157_));
  NO2        o141(.A(ori_ori_n157_), .B(x3), .Y(ori_ori_n158_));
  NO3        o142(.A(ori_ori_n158_), .B(ori_ori_n149_), .C(ori_ori_n136_), .Y(ori03));
  NO2        o143(.A(ori_ori_n42_), .B(x3), .Y(ori_ori_n160_));
  NO2        o144(.A(x6), .B(ori_ori_n24_), .Y(ori_ori_n161_));
  NA2        o145(.A(x6), .B(ori_ori_n24_), .Y(ori_ori_n162_));
  NO2        o146(.A(ori_ori_n162_), .B(x4), .Y(ori_ori_n163_));
  NO2        o147(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n164_));
  NA2        o148(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n165_));
  NO3        o149(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n166_));
  NO2        o150(.A(x5), .B(x1), .Y(ori_ori_n167_));
  NO2        o151(.A(ori_ori_n165_), .B(ori_ori_n138_), .Y(ori_ori_n168_));
  NO3        o152(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n169_));
  NO2        o153(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  INV        o154(.A(ori_ori_n170_), .Y(ori_ori_n171_));
  AOI220     o155(.A0(ori_ori_n171_), .A1(ori_ori_n42_), .B0(ori_ori_n166_), .B1(ori_ori_n101_), .Y(ori_ori_n172_));
  INV        o156(.A(ori_ori_n172_), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n42_), .B(ori_ori_n37_), .Y(ori_ori_n174_));
  NA2        o158(.A(ori_ori_n174_), .B(ori_ori_n19_), .Y(ori_ori_n175_));
  NO2        o159(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n176_));
  NO2        o160(.A(ori_ori_n176_), .B(x6), .Y(ori_ori_n177_));
  NOi21      o161(.An(ori_ori_n70_), .B(ori_ori_n177_), .Y(ori_ori_n178_));
  NA2        o162(.A(ori_ori_n176_), .B(x6), .Y(ori_ori_n179_));
  AOI210     o163(.A0(ori_ori_n179_), .A1(ori_ori_n178_), .B0(ori_ori_n120_), .Y(ori_ori_n180_));
  OR2        o164(.A(ori_ori_n180_), .B(ori_ori_n143_), .Y(ori_ori_n181_));
  NA2        o165(.A(ori_ori_n37_), .B(ori_ori_n47_), .Y(ori_ori_n182_));
  NA2        o166(.A(ori_ori_n112_), .B(ori_ori_n74_), .Y(ori_ori_n183_));
  NA2        o167(.A(x6), .B(ori_ori_n42_), .Y(ori_ori_n184_));
  OAI210     o168(.A0(ori_ori_n95_), .A1(ori_ori_n66_), .B0(x4), .Y(ori_ori_n185_));
  AOI210     o169(.A0(ori_ori_n185_), .A1(ori_ori_n184_), .B0(ori_ori_n65_), .Y(ori_ori_n186_));
  NA2        o170(.A(ori_ori_n161_), .B(ori_ori_n106_), .Y(ori_ori_n187_));
  NA3        o171(.A(ori_ori_n165_), .B(ori_ori_n101_), .C(x6), .Y(ori_ori_n188_));
  INV        o172(.A(ori_ori_n56_), .Y(ori_ori_n189_));
  NA3        o173(.A(ori_ori_n189_), .B(ori_ori_n188_), .C(ori_ori_n187_), .Y(ori_ori_n190_));
  OAI210     o174(.A0(ori_ori_n190_), .A1(ori_ori_n186_), .B0(x2), .Y(ori_ori_n191_));
  NA3        o175(.A(ori_ori_n191_), .B(ori_ori_n183_), .C(ori_ori_n181_), .Y(ori_ori_n192_));
  AOI210     o176(.A0(ori_ori_n173_), .A1(x8), .B0(ori_ori_n192_), .Y(ori_ori_n193_));
  NO2        o177(.A(ori_ori_n75_), .B(x3), .Y(ori_ori_n194_));
  NA2        o178(.A(ori_ori_n194_), .B(ori_ori_n163_), .Y(ori_ori_n195_));
  NO2        o179(.A(ori_ori_n73_), .B(ori_ori_n24_), .Y(ori_ori_n196_));
  AOI210     o180(.A0(ori_ori_n177_), .A1(ori_ori_n123_), .B0(ori_ori_n196_), .Y(ori_ori_n197_));
  AOI210     o181(.A0(ori_ori_n197_), .A1(ori_ori_n195_), .B0(x2), .Y(ori_ori_n198_));
  AOI220     o182(.A0(ori_ori_n163_), .A1(ori_ori_n152_), .B0(x2), .B1(ori_ori_n56_), .Y(ori_ori_n199_));
  NA2        o183(.A(ori_ori_n37_), .B(ori_ori_n17_), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n200_), .B(ori_ori_n24_), .Y(ori_ori_n201_));
  NA2        o185(.A(ori_ori_n201_), .B(ori_ori_n96_), .Y(ori_ori_n202_));
  NA2        o186(.A(ori_ori_n165_), .B(x6), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n165_), .B(x6), .Y(ori_ori_n204_));
  INV        o188(.A(ori_ori_n204_), .Y(ori_ori_n205_));
  NA3        o189(.A(ori_ori_n205_), .B(ori_ori_n203_), .C(ori_ori_n116_), .Y(ori_ori_n206_));
  NA4        o190(.A(ori_ori_n206_), .B(ori_ori_n202_), .C(ori_ori_n199_), .D(ori_ori_n120_), .Y(ori_ori_n207_));
  NA2        o191(.A(ori_ori_n161_), .B(ori_ori_n176_), .Y(ori_ori_n208_));
  NAi21      o192(.An(x1), .B(x4), .Y(ori_ori_n209_));
  AOI210     o193(.A0(x3), .A1(x2), .B0(ori_ori_n42_), .Y(ori_ori_n210_));
  OAI210     o194(.A0(ori_ori_n111_), .A1(x3), .B0(ori_ori_n210_), .Y(ori_ori_n211_));
  NA2        o195(.A(ori_ori_n211_), .B(ori_ori_n209_), .Y(ori_ori_n212_));
  NA2        o196(.A(ori_ori_n212_), .B(ori_ori_n208_), .Y(ori_ori_n213_));
  NA2        o197(.A(x6), .B(x2), .Y(ori_ori_n214_));
  NA2        o198(.A(x4), .B(ori_ori_n213_), .Y(ori_ori_n215_));
  NO2        o199(.A(x3), .B(ori_ori_n162_), .Y(ori_ori_n216_));
  BUFFER     o200(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  NA2        o201(.A(x4), .B(x0), .Y(ori_ori_n218_));
  NA2        o202(.A(ori_ori_n217_), .B(ori_ori_n36_), .Y(ori_ori_n219_));
  AOI210     o203(.A0(ori_ori_n219_), .A1(ori_ori_n215_), .B0(x8), .Y(ori_ori_n220_));
  OAI210     o204(.A0(x0), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n221_));
  NO2        o205(.A(ori_ori_n221_), .B(ori_ori_n182_), .Y(ori_ori_n222_));
  NO4        o206(.A(ori_ori_n222_), .B(ori_ori_n220_), .C(ori_ori_n207_), .D(ori_ori_n198_), .Y(ori_ori_n223_));
  OAI210     o207(.A0(x1), .A1(ori_ori_n204_), .B0(x2), .Y(ori_ori_n224_));
  OAI210     o208(.A0(x0), .A1(x6), .B0(ori_ori_n38_), .Y(ori_ori_n225_));
  AOI210     o209(.A0(ori_ori_n225_), .A1(ori_ori_n224_), .B0(ori_ori_n151_), .Y(ori_ori_n226_));
  NOi21      o210(.An(ori_ori_n214_), .B(ori_ori_n17_), .Y(ori_ori_n227_));
  NA3        o211(.A(ori_ori_n227_), .B(ori_ori_n167_), .C(ori_ori_n34_), .Y(ori_ori_n228_));
  AOI210     o212(.A0(ori_ori_n32_), .A1(ori_ori_n47_), .B0(x0), .Y(ori_ori_n229_));
  NA3        o213(.A(ori_ori_n229_), .B(ori_ori_n129_), .C(ori_ori_n29_), .Y(ori_ori_n230_));
  NA2        o214(.A(x3), .B(x2), .Y(ori_ori_n231_));
  AOI220     o215(.A0(ori_ori_n231_), .A1(ori_ori_n182_), .B0(ori_ori_n230_), .B1(ori_ori_n228_), .Y(ori_ori_n232_));
  NAi21      o216(.An(x4), .B(x0), .Y(ori_ori_n233_));
  NO3        o217(.A(ori_ori_n233_), .B(ori_ori_n38_), .C(x2), .Y(ori_ori_n234_));
  OAI210     o218(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n234_), .Y(ori_ori_n235_));
  OAI220     o219(.A0(ori_ori_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n236_));
  NO2        o220(.A(ori_ori_n229_), .B(ori_ori_n227_), .Y(ori_ori_n237_));
  AOI220     o221(.A0(ori_ori_n237_), .A1(ori_ori_n69_), .B0(ori_ori_n236_), .B1(ori_ori_n28_), .Y(ori_ori_n238_));
  AOI210     o222(.A0(ori_ori_n238_), .A1(ori_ori_n235_), .B0(ori_ori_n24_), .Y(ori_ori_n239_));
  NO2        o223(.A(ori_ori_n229_), .B(ori_ori_n227_), .Y(ori_ori_n240_));
  INV        o224(.A(ori_ori_n168_), .Y(ori_ori_n241_));
  NA2        o225(.A(ori_ori_n32_), .B(ori_ori_n37_), .Y(ori_ori_n242_));
  OR2        o226(.A(ori_ori_n242_), .B(ori_ori_n218_), .Y(ori_ori_n243_));
  OAI220     o227(.A0(ori_ori_n243_), .A1(ori_ori_n128_), .B0(ori_ori_n184_), .B1(ori_ori_n241_), .Y(ori_ori_n244_));
  AO210      o228(.A0(ori_ori_n240_), .A1(ori_ori_n118_), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  NO4        o229(.A(ori_ori_n245_), .B(ori_ori_n239_), .C(ori_ori_n232_), .D(ori_ori_n226_), .Y(ori_ori_n246_));
  OAI210     o230(.A0(ori_ori_n223_), .A1(ori_ori_n193_), .B0(ori_ori_n246_), .Y(ori04));
  NO2        o231(.A(x2), .B(x1), .Y(ori_ori_n248_));
  OAI210     o232(.A0(ori_ori_n200_), .A1(ori_ori_n248_), .B0(ori_ori_n32_), .Y(ori_ori_n249_));
  INV        o233(.A(ori_ori_n233_), .Y(ori_ori_n250_));
  OAI210     o234(.A0(ori_ori_n47_), .A1(ori_ori_n250_), .B0(ori_ori_n194_), .Y(ori_ori_n251_));
  NO2        o235(.A(ori_ori_n231_), .B(ori_ori_n164_), .Y(ori_ori_n252_));
  NA2        o236(.A(ori_ori_n252_), .B(ori_ori_n75_), .Y(ori_ori_n253_));
  NA3        o237(.A(ori_ori_n253_), .B(x6), .C(ori_ori_n251_), .Y(ori_ori_n254_));
  NA2        o238(.A(ori_ori_n254_), .B(ori_ori_n249_), .Y(ori_ori_n255_));
  OAI210     o239(.A0(ori_ori_n94_), .A1(ori_ori_n88_), .B0(ori_ori_n142_), .Y(ori_ori_n256_));
  NA3        o240(.A(ori_ori_n256_), .B(x6), .C(x3), .Y(ori_ori_n257_));
  AOI210     o241(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n258_));
  NO2        o242(.A(ori_ori_n258_), .B(ori_ori_n242_), .Y(ori_ori_n259_));
  INV        o243(.A(ori_ori_n259_), .Y(ori_ori_n260_));
  NA2        o244(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n261_));
  INV        o245(.A(ori_ori_n261_), .Y(ori_ori_n262_));
  NA2        o246(.A(ori_ori_n262_), .B(ori_ori_n66_), .Y(ori_ori_n263_));
  NA3        o247(.A(ori_ori_n263_), .B(ori_ori_n260_), .C(ori_ori_n257_), .Y(ori_ori_n264_));
  OAI210     o248(.A0(ori_ori_n92_), .A1(x3), .B0(ori_ori_n234_), .Y(ori_ori_n265_));
  NA2        o249(.A(ori_ori_n166_), .B(ori_ori_n70_), .Y(ori_ori_n266_));
  NA3        o250(.A(ori_ori_n266_), .B(ori_ori_n265_), .C(ori_ori_n120_), .Y(ori_ori_n267_));
  AOI210     o251(.A0(ori_ori_n264_), .A1(x4), .B0(ori_ori_n267_), .Y(ori_ori_n268_));
  NOi21      o252(.An(x4), .B(x0), .Y(ori_ori_n269_));
  XO2        o253(.A(x4), .B(x0), .Y(ori_ori_n270_));
  INV        o254(.A(ori_ori_n209_), .Y(ori_ori_n271_));
  AOI220     o255(.A0(ori_ori_n271_), .A1(x8), .B0(ori_ori_n269_), .B1(ori_ori_n76_), .Y(ori_ori_n272_));
  NO2        o256(.A(ori_ori_n272_), .B(x3), .Y(ori_ori_n273_));
  INV        o257(.A(ori_ori_n76_), .Y(ori_ori_n274_));
  NO2        o258(.A(ori_ori_n75_), .B(x4), .Y(ori_ori_n275_));
  AOI220     o259(.A0(ori_ori_n275_), .A1(ori_ori_n38_), .B0(ori_ori_n99_), .B1(ori_ori_n274_), .Y(ori_ori_n276_));
  NO2        o260(.A(ori_ori_n270_), .B(x2), .Y(ori_ori_n277_));
  INV        o261(.A(ori_ori_n277_), .Y(ori_ori_n278_));
  NA4        o262(.A(ori_ori_n278_), .B(ori_ori_n276_), .C(ori_ori_n175_), .D(x6), .Y(ori_ori_n279_));
  NO2        o263(.A(ori_ori_n144_), .B(ori_ori_n75_), .Y(ori_ori_n280_));
  NA2        o264(.A(ori_ori_n280_), .B(ori_ori_n54_), .Y(ori_ori_n281_));
  NO2        o265(.A(x8), .B(ori_ori_n68_), .Y(ori_ori_n282_));
  NO2        o266(.A(ori_ori_n31_), .B(x2), .Y(ori_ori_n283_));
  NA2        o267(.A(ori_ori_n283_), .B(ori_ori_n282_), .Y(ori_ori_n284_));
  NA2        o268(.A(ori_ori_n281_), .B(ori_ori_n284_), .Y(ori_ori_n285_));
  OAI220     o269(.A0(ori_ori_n285_), .A1(x6), .B0(ori_ori_n279_), .B1(ori_ori_n273_), .Y(ori_ori_n286_));
  NA2        o270(.A(ori_ori_n42_), .B(ori_ori_n36_), .Y(ori_ori_n287_));
  OAI210     o271(.A0(ori_ori_n287_), .A1(ori_ori_n75_), .B0(ori_ori_n243_), .Y(ori_ori_n288_));
  AOI210     o272(.A0(ori_ori_n288_), .A1(ori_ori_n18_), .B0(ori_ori_n120_), .Y(ori_ori_n289_));
  AO220      o273(.A0(ori_ori_n289_), .A1(ori_ori_n286_), .B0(ori_ori_n268_), .B1(ori_ori_n255_), .Y(ori_ori_n290_));
  NA2        o274(.A(ori_ori_n283_), .B(x6), .Y(ori_ori_n291_));
  AOI210     o275(.A0(x6), .A1(x1), .B0(ori_ori_n119_), .Y(ori_ori_n292_));
  NA2        o276(.A(ori_ori_n275_), .B(x0), .Y(ori_ori_n293_));
  NA2        o277(.A(ori_ori_n70_), .B(x6), .Y(ori_ori_n294_));
  OAI210     o278(.A0(ori_ori_n293_), .A1(ori_ori_n292_), .B0(ori_ori_n294_), .Y(ori_ori_n295_));
  AOI220     o279(.A0(ori_ori_n295_), .A1(ori_ori_n291_), .B0(ori_ori_n169_), .B1(ori_ori_n43_), .Y(ori_ori_n296_));
  NA2        o280(.A(ori_ori_n296_), .B(ori_ori_n290_), .Y(ori_ori_n297_));
  INV        o281(.A(ori_ori_n92_), .Y(ori_ori_n298_));
  NA2        o282(.A(ori_ori_n298_), .B(ori_ori_n261_), .Y(ori_ori_n299_));
  NA3        o283(.A(ori_ori_n299_), .B(ori_ori_n160_), .C(ori_ori_n120_), .Y(ori_ori_n300_));
  NA3        o284(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n301_));
  NA2        o285(.A(ori_ori_n174_), .B(x0), .Y(ori_ori_n302_));
  OAI220     o286(.A0(ori_ori_n302_), .A1(x2), .B0(ori_ori_n301_), .B1(ori_ori_n274_), .Y(ori_ori_n303_));
  INV        o287(.A(ori_ori_n303_), .Y(ori_ori_n304_));
  AOI210     o288(.A0(ori_ori_n304_), .A1(ori_ori_n300_), .B0(ori_ori_n24_), .Y(ori_ori_n305_));
  NA2        o289(.A(ori_ori_n305_), .B(x6), .Y(ori_ori_n306_));
  NO2        o290(.A(ori_ori_n29_), .B(x0), .Y(ori_ori_n307_));
  NA2        o291(.A(ori_ori_n160_), .B(ori_ori_n120_), .Y(ori_ori_n308_));
  OAI210     o292(.A0(ori_ori_n308_), .A1(x8), .B0(ori_ori_n354_), .Y(ori_ori_n309_));
  NAi31      o293(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n310_));
  OAI210     o294(.A0(ori_ori_n310_), .A1(x4), .B0(ori_ori_n131_), .Y(ori_ori_n311_));
  NA3        o295(.A(ori_ori_n311_), .B(ori_ori_n117_), .C(x9), .Y(ori_ori_n312_));
  NA2        o296(.A(ori_ori_n282_), .B(ori_ori_n120_), .Y(ori_ori_n313_));
  NA4        o297(.A(ori_ori_n313_), .B(x1), .C(ori_ori_n312_), .D(ori_ori_n44_), .Y(ori_ori_n314_));
  OAI210     o298(.A0(ori_ori_n309_), .A1(ori_ori_n307_), .B0(ori_ori_n314_), .Y(ori_ori_n315_));
  INV        o299(.A(ori_ori_n105_), .Y(ori_ori_n316_));
  NO2        o300(.A(ori_ori_n316_), .B(ori_ori_n37_), .Y(ori_ori_n317_));
  AOI210     o301(.A0(ori_ori_n209_), .A1(ori_ori_n53_), .B0(ori_ori_n98_), .Y(ori_ori_n318_));
  NO2        o302(.A(ori_ori_n318_), .B(x3), .Y(ori_ori_n319_));
  NO3        o303(.A(ori_ori_n319_), .B(ori_ori_n317_), .C(x2), .Y(ori_ori_n320_));
  OAI210     o304(.A0(ori_ori_n233_), .A1(ori_ori_n37_), .B0(ori_ori_n270_), .Y(ori_ori_n321_));
  INV        o305(.A(ori_ori_n301_), .Y(ori_ori_n322_));
  AOI220     o306(.A0(ori_ori_n322_), .A1(ori_ori_n75_), .B0(ori_ori_n321_), .B1(ori_ori_n120_), .Y(ori_ori_n323_));
  NO2        o307(.A(ori_ori_n323_), .B(ori_ori_n47_), .Y(ori_ori_n324_));
  NO2        o308(.A(ori_ori_n324_), .B(ori_ori_n320_), .Y(ori_ori_n325_));
  AOI210     o309(.A0(ori_ori_n325_), .A1(ori_ori_n315_), .B0(ori_ori_n24_), .Y(ori_ori_n326_));
  NA4        o310(.A(ori_ori_n28_), .B(ori_ori_n75_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n327_));
  NO3        o311(.A(ori_ori_n57_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n328_));
  NA2        o312(.A(ori_ori_n328_), .B(ori_ori_n210_), .Y(ori_ori_n329_));
  NO2        o313(.A(ori_ori_n329_), .B(ori_ori_n85_), .Y(ori_ori_n330_));
  NA2        o314(.A(ori_ori_n330_), .B(x7), .Y(ori_ori_n331_));
  INV        o315(.A(x7), .Y(ori_ori_n332_));
  NA3        o316(.A(ori_ori_n332_), .B(ori_ori_n119_), .C(ori_ori_n106_), .Y(ori_ori_n333_));
  NA3        o317(.A(ori_ori_n333_), .B(ori_ori_n331_), .C(ori_ori_n327_), .Y(ori_ori_n334_));
  OAI210     o318(.A0(ori_ori_n334_), .A1(ori_ori_n326_), .B0(ori_ori_n32_), .Y(ori_ori_n335_));
  INV        o319(.A(ori_ori_n164_), .Y(ori_ori_n336_));
  NO4        o320(.A(ori_ori_n336_), .B(ori_ori_n65_), .C(x4), .D(ori_ori_n47_), .Y(ori_ori_n337_));
  NA2        o321(.A(ori_ori_n200_), .B(ori_ori_n21_), .Y(ori_ori_n338_));
  NO2        o322(.A(ori_ori_n128_), .B(ori_ori_n107_), .Y(ori_ori_n339_));
  NA2        o323(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n340_));
  NO2        o324(.A(ori_ori_n340_), .B(ori_ori_n26_), .Y(ori_ori_n341_));
  NA2        o325(.A(ori_ori_n310_), .B(ori_ori_n73_), .Y(ori_ori_n342_));
  NA2        o326(.A(ori_ori_n342_), .B(ori_ori_n143_), .Y(ori_ori_n343_));
  OAI220     o327(.A0(x3), .A1(ori_ori_n58_), .B0(ori_ori_n128_), .B1(ori_ori_n37_), .Y(ori_ori_n344_));
  NA2        o328(.A(x3), .B(ori_ori_n47_), .Y(ori_ori_n345_));
  NO2        o329(.A(ori_ori_n121_), .B(ori_ori_n345_), .Y(ori_ori_n346_));
  AOI220     o330(.A0(ori_ori_n346_), .A1(x0), .B0(ori_ori_n344_), .B1(ori_ori_n107_), .Y(ori_ori_n347_));
  AOI210     o331(.A0(ori_ori_n347_), .A1(ori_ori_n343_), .B0(ori_ori_n184_), .Y(ori_ori_n348_));
  NO3        o332(.A(ori_ori_n348_), .B(ori_ori_n341_), .C(ori_ori_n337_), .Y(ori_ori_n349_));
  NA3        o333(.A(ori_ori_n349_), .B(ori_ori_n335_), .C(ori_ori_n306_), .Y(ori_ori_n350_));
  AOI210     o334(.A0(ori_ori_n297_), .A1(ori_ori_n24_), .B0(ori_ori_n350_), .Y(ori05));
  INV        o335(.A(x1), .Y(ori_ori_n354_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  AN2        m021(.A(x8), .B(x7), .Y(mai_mai_n38_));
  NA3        m022(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m023(.A(x4), .B(x3), .Y(mai_mai_n40_));
  AOI210     m024(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(x2), .B(x0), .Y(mai_mai_n42_));
  INV        m026(.A(x3), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n44_));
  INV        m028(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n42_), .Y(mai_mai_n47_));
  INV        m031(.A(x4), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(x2), .Y(mai_mai_n50_));
  OAI210     m034(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n47_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n38_), .B(mai_mai_n37_), .Y(mai_mai_n52_));
  AOI220     m036(.A0(mai_mai_n52_), .A1(mai_mai_n35_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n53_));
  INV        m037(.A(x2), .Y(mai_mai_n54_));
  NO2        m038(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  OAI210     m041(.A0(mai_mai_n53_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai01));
  NA2        m043(.A(x8), .B(x7), .Y(mai_mai_n60_));
  NA2        m044(.A(mai_mai_n43_), .B(x1), .Y(mai_mai_n61_));
  INV        m045(.A(x9), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n62_), .B(mai_mai_n36_), .Y(mai_mai_n63_));
  NO3        m047(.A(mai_mai_n36_), .B(mai_mai_n61_), .C(mai_mai_n60_), .Y(mai_mai_n64_));
  NO2        m048(.A(x7), .B(x6), .Y(mai_mai_n65_));
  NO2        m049(.A(mai_mai_n61_), .B(x5), .Y(mai_mai_n66_));
  NO2        m050(.A(x8), .B(x2), .Y(mai_mai_n67_));
  OA210      m051(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n65_), .Y(mai_mai_n68_));
  OAI210     m052(.A0(mai_mai_n44_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n56_), .A1(mai_mai_n20_), .B0(mai_mai_n69_), .Y(mai_mai_n70_));
  NAi31      m054(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n71_));
  NO2        m055(.A(mai_mai_n70_), .B(mai_mai_n68_), .Y(mai_mai_n72_));
  OAI210     m056(.A0(mai_mai_n72_), .A1(mai_mai_n64_), .B0(x4), .Y(mai_mai_n73_));
  NA2        m057(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n74_));
  OAI210     m058(.A0(mai_mai_n74_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n75_));
  NA2        m059(.A(x5), .B(x3), .Y(mai_mai_n76_));
  NO2        m060(.A(x8), .B(x6), .Y(mai_mai_n77_));
  NO4        m061(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(mai_mai_n65_), .D(mai_mai_n54_), .Y(mai_mai_n78_));
  NAi21      m062(.An(x4), .B(x3), .Y(mai_mai_n79_));
  INV        m063(.A(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m064(.A(mai_mai_n80_), .B(mai_mai_n22_), .Y(mai_mai_n81_));
  NO2        m065(.A(x4), .B(x2), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(x3), .Y(mai_mai_n83_));
  NO3        m067(.A(mai_mai_n83_), .B(mai_mai_n81_), .C(mai_mai_n18_), .Y(mai_mai_n84_));
  NO3        m068(.A(mai_mai_n84_), .B(mai_mai_n78_), .C(mai_mai_n75_), .Y(mai_mai_n85_));
  NO4        m069(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n43_), .D(x1), .Y(mai_mai_n86_));
  NA2        m070(.A(mai_mai_n62_), .B(mai_mai_n48_), .Y(mai_mai_n87_));
  INV        m071(.A(mai_mai_n87_), .Y(mai_mai_n88_));
  OAI210     m072(.A0(mai_mai_n86_), .A1(mai_mai_n66_), .B0(mai_mai_n88_), .Y(mai_mai_n89_));
  NA2        m073(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n90_), .B(mai_mai_n25_), .Y(mai_mai_n91_));
  INV        m075(.A(x8), .Y(mai_mai_n92_));
  NA2        m076(.A(x2), .B(x1), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n92_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n91_), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n95_), .B(mai_mai_n26_), .Y(mai_mai_n96_));
  AOI210     m080(.A0(mai_mai_n56_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n97_));
  OAI210     m081(.A0(mai_mai_n45_), .A1(mai_mai_n37_), .B0(mai_mai_n48_), .Y(mai_mai_n98_));
  NO3        m082(.A(mai_mai_n98_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n99_));
  NA2        m083(.A(x4), .B(mai_mai_n43_), .Y(mai_mai_n100_));
  NO2        m084(.A(mai_mai_n48_), .B(mai_mai_n54_), .Y(mai_mai_n101_));
  OAI210     m085(.A0(mai_mai_n101_), .A1(mai_mai_n43_), .B0(mai_mai_n18_), .Y(mai_mai_n102_));
  AOI210     m086(.A0(mai_mai_n100_), .A1(mai_mai_n52_), .B0(mai_mai_n102_), .Y(mai_mai_n103_));
  NO2        m087(.A(x3), .B(x2), .Y(mai_mai_n104_));
  NA2        m088(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n105_));
  OAI210     m089(.A0(mai_mai_n105_), .A1(mai_mai_n40_), .B0(mai_mai_n17_), .Y(mai_mai_n106_));
  NO3        m090(.A(mai_mai_n106_), .B(mai_mai_n103_), .C(mai_mai_n99_), .Y(mai_mai_n107_));
  AO220      m091(.A0(mai_mai_n107_), .A1(mai_mai_n89_), .B0(mai_mai_n85_), .B1(mai_mai_n73_), .Y(mai02));
  NO2        m092(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n109_));
  NO2        m093(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n110_));
  AOI220     m094(.A0(mai_mai_n54_), .A1(mai_mai_n110_), .B0(mai_mai_n109_), .B1(x4), .Y(mai_mai_n111_));
  NO3        m095(.A(mai_mai_n111_), .B(x7), .C(x5), .Y(mai_mai_n112_));
  NA2        m096(.A(x9), .B(x2), .Y(mai_mai_n113_));
  OR2        m097(.A(x8), .B(x0), .Y(mai_mai_n114_));
  INV        m098(.A(mai_mai_n114_), .Y(mai_mai_n115_));
  NAi21      m099(.An(x2), .B(x8), .Y(mai_mai_n116_));
  INV        m100(.A(mai_mai_n116_), .Y(mai_mai_n117_));
  NO2        m101(.A(x4), .B(x1), .Y(mai_mai_n118_));
  NOi21      m102(.An(x0), .B(x1), .Y(mai_mai_n119_));
  NO3        m103(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n120_));
  NOi21      m104(.An(x0), .B(x4), .Y(mai_mai_n121_));
  NO2        m105(.A(x8), .B(mai_mai_n62_), .Y(mai_mai_n122_));
  AOI220     m106(.A0(mai_mai_n122_), .A1(mai_mai_n121_), .B0(mai_mai_n120_), .B1(mai_mai_n119_), .Y(mai_mai_n123_));
  NO2        m107(.A(mai_mai_n123_), .B(mai_mai_n76_), .Y(mai_mai_n124_));
  NO2        m108(.A(x5), .B(mai_mai_n48_), .Y(mai_mai_n125_));
  NA2        m109(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n126_));
  AOI210     m110(.A0(mai_mai_n126_), .A1(mai_mai_n105_), .B0(x3), .Y(mai_mai_n127_));
  OAI210     m111(.A0(mai_mai_n127_), .A1(mai_mai_n35_), .B0(mai_mai_n125_), .Y(mai_mai_n128_));
  NAi21      m112(.An(x0), .B(x4), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n129_), .B(x1), .Y(mai_mai_n130_));
  NO2        m114(.A(x7), .B(x0), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n82_), .B(mai_mai_n101_), .Y(mai_mai_n132_));
  NO2        m116(.A(mai_mai_n132_), .B(x3), .Y(mai_mai_n133_));
  OAI210     m117(.A0(mai_mai_n131_), .A1(mai_mai_n130_), .B0(mai_mai_n133_), .Y(mai_mai_n134_));
  NO2        m118(.A(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n135_));
  NA2        m119(.A(x5), .B(x0), .Y(mai_mai_n136_));
  NO2        m120(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n137_));
  NA3        m121(.A(mai_mai_n137_), .B(mai_mai_n136_), .C(mai_mai_n135_), .Y(mai_mai_n138_));
  NA4        m122(.A(mai_mai_n138_), .B(mai_mai_n134_), .C(mai_mai_n128_), .D(mai_mai_n36_), .Y(mai_mai_n139_));
  NO3        m123(.A(mai_mai_n139_), .B(mai_mai_n124_), .C(mai_mai_n112_), .Y(mai_mai_n140_));
  NO3        m124(.A(mai_mai_n76_), .B(mai_mai_n74_), .C(mai_mai_n24_), .Y(mai_mai_n141_));
  NO2        m125(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n142_));
  AOI220     m126(.A0(mai_mai_n119_), .A1(mai_mai_n142_), .B0(mai_mai_n66_), .B1(mai_mai_n17_), .Y(mai_mai_n143_));
  NO3        m127(.A(mai_mai_n143_), .B(mai_mai_n60_), .C(mai_mai_n62_), .Y(mai_mai_n144_));
  NA2        m128(.A(x7), .B(x3), .Y(mai_mai_n145_));
  NO2        m129(.A(mai_mai_n100_), .B(x5), .Y(mai_mai_n146_));
  NO2        m130(.A(x9), .B(x7), .Y(mai_mai_n147_));
  NOi21      m131(.An(x8), .B(x0), .Y(mai_mai_n148_));
  NO2        m132(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n149_));
  INV        m133(.A(x7), .Y(mai_mai_n150_));
  NA2        m134(.A(mai_mai_n150_), .B(mai_mai_n18_), .Y(mai_mai_n151_));
  AOI220     m135(.A0(mai_mai_n151_), .A1(mai_mai_n149_), .B0(mai_mai_n109_), .B1(mai_mai_n38_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n153_), .B(mai_mai_n121_), .Y(mai_mai_n154_));
  NO2        m138(.A(mai_mai_n154_), .B(mai_mai_n152_), .Y(mai_mai_n155_));
  AOI210     m139(.A0(mai_mai_n148_), .A1(mai_mai_n146_), .B0(mai_mai_n155_), .Y(mai_mai_n156_));
  OAI210     m140(.A0(mai_mai_n145_), .A1(mai_mai_n50_), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  NA2        m141(.A(x5), .B(x1), .Y(mai_mai_n158_));
  INV        m142(.A(mai_mai_n158_), .Y(mai_mai_n159_));
  AOI210     m143(.A0(mai_mai_n159_), .A1(mai_mai_n121_), .B0(mai_mai_n36_), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n62_), .B(mai_mai_n92_), .Y(mai_mai_n161_));
  NAi21      m145(.An(x2), .B(x7), .Y(mai_mai_n162_));
  NAi31      m146(.An(mai_mai_n76_), .B(mai_mai_n38_), .C(mai_mai_n35_), .Y(mai_mai_n163_));
  NA2        m147(.A(mai_mai_n163_), .B(mai_mai_n160_), .Y(mai_mai_n164_));
  NO4        m148(.A(mai_mai_n164_), .B(mai_mai_n157_), .C(mai_mai_n144_), .D(mai_mai_n141_), .Y(mai_mai_n165_));
  NO2        m149(.A(mai_mai_n165_), .B(mai_mai_n140_), .Y(mai_mai_n166_));
  NO2        m150(.A(mai_mai_n136_), .B(mai_mai_n132_), .Y(mai_mai_n167_));
  NA2        m151(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n168_));
  NA2        m152(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n169_));
  NA3        m153(.A(mai_mai_n169_), .B(mai_mai_n168_), .C(mai_mai_n24_), .Y(mai_mai_n170_));
  AN2        m154(.A(mai_mai_n170_), .B(mai_mai_n137_), .Y(mai_mai_n171_));
  NA2        m155(.A(x8), .B(x0), .Y(mai_mai_n172_));
  NO2        m156(.A(mai_mai_n150_), .B(mai_mai_n25_), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n119_), .B(x4), .Y(mai_mai_n174_));
  NA2        m158(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  AOI210     m159(.A0(mai_mai_n172_), .A1(mai_mai_n126_), .B0(mai_mai_n175_), .Y(mai_mai_n176_));
  NA2        m160(.A(x2), .B(x0), .Y(mai_mai_n177_));
  NA2        m161(.A(x4), .B(x1), .Y(mai_mai_n178_));
  NAi21      m162(.An(mai_mai_n118_), .B(mai_mai_n178_), .Y(mai_mai_n179_));
  NOi31      m163(.An(mai_mai_n179_), .B(mai_mai_n153_), .C(mai_mai_n177_), .Y(mai_mai_n180_));
  NO4        m164(.A(mai_mai_n180_), .B(mai_mai_n176_), .C(mai_mai_n171_), .D(mai_mai_n167_), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n181_), .B(mai_mai_n43_), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n170_), .B(mai_mai_n74_), .Y(mai_mai_n183_));
  INV        m167(.A(mai_mai_n125_), .Y(mai_mai_n184_));
  NO2        m168(.A(mai_mai_n105_), .B(mai_mai_n17_), .Y(mai_mai_n185_));
  NO3        m169(.A(mai_mai_n105_), .B(mai_mai_n184_), .C(x7), .Y(mai_mai_n186_));
  NA3        m170(.A(mai_mai_n179_), .B(mai_mai_n184_), .C(mai_mai_n42_), .Y(mai_mai_n187_));
  OAI210     m171(.A0(mai_mai_n169_), .A1(mai_mai_n132_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  NO3        m172(.A(mai_mai_n188_), .B(mai_mai_n186_), .C(mai_mai_n183_), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n189_), .B(x3), .Y(mai_mai_n190_));
  NO3        m174(.A(mai_mai_n190_), .B(mai_mai_n182_), .C(mai_mai_n166_), .Y(mai03));
  NO2        m175(.A(mai_mai_n48_), .B(x3), .Y(mai_mai_n192_));
  NO2        m176(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n193_));
  INV        m177(.A(mai_mai_n193_), .Y(mai_mai_n194_));
  NO2        m178(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n195_));
  OAI210     m179(.A0(mai_mai_n195_), .A1(mai_mai_n25_), .B0(mai_mai_n63_), .Y(mai_mai_n196_));
  OAI220     m180(.A0(mai_mai_n196_), .A1(mai_mai_n17_), .B0(mai_mai_n194_), .B1(mai_mai_n105_), .Y(mai_mai_n197_));
  NA2        m181(.A(mai_mai_n197_), .B(mai_mai_n192_), .Y(mai_mai_n198_));
  NO2        m182(.A(mai_mai_n76_), .B(x6), .Y(mai_mai_n199_));
  NA2        m183(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n200_));
  NO2        m184(.A(mai_mai_n200_), .B(x4), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n202_));
  AO220      m186(.A0(mai_mai_n202_), .A1(mai_mai_n201_), .B0(mai_mai_n199_), .B1(mai_mai_n55_), .Y(mai_mai_n203_));
  NA2        m187(.A(mai_mai_n203_), .B(mai_mai_n62_), .Y(mai_mai_n204_));
  NA2        m188(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n205_));
  NO2        m189(.A(mai_mai_n205_), .B(mai_mai_n200_), .Y(mai_mai_n206_));
  NA2        m190(.A(x9), .B(mai_mai_n54_), .Y(mai_mai_n207_));
  NA2        m191(.A(mai_mai_n200_), .B(mai_mai_n79_), .Y(mai_mai_n208_));
  AOI210     m192(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n177_), .Y(mai_mai_n209_));
  AOI220     m193(.A0(mai_mai_n209_), .A1(mai_mai_n208_), .B0(x9), .B1(mai_mai_n206_), .Y(mai_mai_n210_));
  NO2        m194(.A(x5), .B(x1), .Y(mai_mai_n211_));
  AOI220     m195(.A0(mai_mai_n211_), .A1(mai_mai_n17_), .B0(mai_mai_n104_), .B1(x5), .Y(mai_mai_n212_));
  NO2        m196(.A(mai_mai_n205_), .B(mai_mai_n168_), .Y(mai_mai_n213_));
  INV        m197(.A(mai_mai_n213_), .Y(mai_mai_n214_));
  OAI210     m198(.A0(mai_mai_n212_), .A1(mai_mai_n36_), .B0(mai_mai_n214_), .Y(mai_mai_n215_));
  NA2        m199(.A(mai_mai_n215_), .B(mai_mai_n48_), .Y(mai_mai_n216_));
  NA4        m200(.A(mai_mai_n216_), .B(mai_mai_n210_), .C(mai_mai_n204_), .D(mai_mai_n198_), .Y(mai_mai_n217_));
  NO2        m201(.A(mai_mai_n48_), .B(mai_mai_n43_), .Y(mai_mai_n218_));
  NA2        m202(.A(mai_mai_n218_), .B(mai_mai_n19_), .Y(mai_mai_n219_));
  NO2        m203(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n220_));
  NO2        m204(.A(mai_mai_n220_), .B(x6), .Y(mai_mai_n221_));
  NOi21      m205(.An(mai_mai_n82_), .B(mai_mai_n221_), .Y(mai_mai_n222_));
  NA2        m206(.A(mai_mai_n62_), .B(mai_mai_n92_), .Y(mai_mai_n223_));
  NO2        m207(.A(mai_mai_n222_), .B(mai_mai_n150_), .Y(mai_mai_n224_));
  AO210      m208(.A0(mai_mai_n224_), .A1(mai_mai_n219_), .B0(mai_mai_n173_), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n43_), .B(mai_mai_n54_), .Y(mai_mai_n226_));
  NO3        m210(.A(mai_mai_n178_), .B(mai_mai_n62_), .C(x6), .Y(mai_mai_n227_));
  AOI220     m211(.A0(mai_mai_n227_), .A1(mai_mai_n17_), .B0(mai_mai_n137_), .B1(mai_mai_n91_), .Y(mai_mai_n228_));
  NA2        m212(.A(x6), .B(mai_mai_n48_), .Y(mai_mai_n229_));
  NO2        m213(.A(mai_mai_n229_), .B(mai_mai_n76_), .Y(mai_mai_n230_));
  NO2        m214(.A(mai_mai_n158_), .B(mai_mai_n43_), .Y(mai_mai_n231_));
  OAI210     m215(.A0(mai_mai_n231_), .A1(mai_mai_n213_), .B0(mai_mai_n435_), .Y(mai_mai_n232_));
  NA2        m216(.A(mai_mai_n193_), .B(mai_mai_n130_), .Y(mai_mai_n233_));
  NA3        m217(.A(mai_mai_n205_), .B(mai_mai_n125_), .C(x6), .Y(mai_mai_n234_));
  OAI210     m218(.A0(mai_mai_n92_), .A1(mai_mai_n36_), .B0(mai_mai_n66_), .Y(mai_mai_n235_));
  NA4        m219(.A(mai_mai_n235_), .B(mai_mai_n234_), .C(mai_mai_n233_), .D(mai_mai_n232_), .Y(mai_mai_n236_));
  OAI210     m220(.A0(mai_mai_n236_), .A1(mai_mai_n230_), .B0(x2), .Y(mai_mai_n237_));
  NA3        m221(.A(mai_mai_n237_), .B(mai_mai_n228_), .C(mai_mai_n225_), .Y(mai_mai_n238_));
  AOI210     m222(.A0(mai_mai_n217_), .A1(x8), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  NO2        m223(.A(mai_mai_n92_), .B(x3), .Y(mai_mai_n240_));
  NO3        m224(.A(mai_mai_n90_), .B(mai_mai_n77_), .C(mai_mai_n25_), .Y(mai_mai_n241_));
  AOI210     m225(.A0(mai_mai_n221_), .A1(mai_mai_n153_), .B0(mai_mai_n241_), .Y(mai_mai_n242_));
  NO2        m226(.A(mai_mai_n242_), .B(x2), .Y(mai_mai_n243_));
  NO2        m227(.A(x4), .B(mai_mai_n54_), .Y(mai_mai_n244_));
  AOI220     m228(.A0(mai_mai_n201_), .A1(mai_mai_n185_), .B0(mai_mai_n244_), .B1(mai_mai_n66_), .Y(mai_mai_n245_));
  NA2        m229(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n246_));
  NA3        m230(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n247_));
  AOI210     m231(.A0(mai_mai_n247_), .A1(mai_mai_n136_), .B0(mai_mai_n246_), .Y(mai_mai_n248_));
  NA2        m232(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n249_));
  NO2        m233(.A(mai_mai_n249_), .B(mai_mai_n25_), .Y(mai_mai_n250_));
  OAI210     m234(.A0(mai_mai_n250_), .A1(mai_mai_n248_), .B0(mai_mai_n118_), .Y(mai_mai_n251_));
  NA2        m235(.A(mai_mai_n205_), .B(x6), .Y(mai_mai_n252_));
  NO2        m236(.A(mai_mai_n205_), .B(x6), .Y(mai_mai_n253_));
  NA2        m237(.A(mai_mai_n252_), .B(mai_mai_n142_), .Y(mai_mai_n254_));
  NA4        m238(.A(mai_mai_n254_), .B(mai_mai_n251_), .C(mai_mai_n245_), .D(mai_mai_n150_), .Y(mai_mai_n255_));
  NA2        m239(.A(mai_mai_n193_), .B(mai_mai_n220_), .Y(mai_mai_n256_));
  NO2        m240(.A(x9), .B(x6), .Y(mai_mai_n257_));
  NO2        m241(.A(mai_mai_n136_), .B(mai_mai_n18_), .Y(mai_mai_n258_));
  NAi21      m242(.An(mai_mai_n258_), .B(mai_mai_n247_), .Y(mai_mai_n259_));
  NAi21      m243(.An(x1), .B(x4), .Y(mai_mai_n260_));
  AOI220     m244(.A0(mai_mai_n48_), .A1(mai_mai_n260_), .B0(mai_mai_n259_), .B1(mai_mai_n257_), .Y(mai_mai_n261_));
  NA2        m245(.A(mai_mai_n261_), .B(mai_mai_n256_), .Y(mai_mai_n262_));
  NA2        m246(.A(mai_mai_n62_), .B(x2), .Y(mai_mai_n263_));
  NO2        m247(.A(mai_mai_n263_), .B(mai_mai_n256_), .Y(mai_mai_n264_));
  NO3        m248(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n265_));
  NA2        m249(.A(mai_mai_n105_), .B(mai_mai_n25_), .Y(mai_mai_n266_));
  NA2        m250(.A(x6), .B(x2), .Y(mai_mai_n267_));
  NO2        m251(.A(mai_mai_n267_), .B(mai_mai_n168_), .Y(mai_mai_n268_));
  AOI210     m252(.A0(mai_mai_n266_), .A1(mai_mai_n265_), .B0(mai_mai_n268_), .Y(mai_mai_n269_));
  OAI220     m253(.A0(mai_mai_n269_), .A1(mai_mai_n43_), .B0(mai_mai_n174_), .B1(mai_mai_n46_), .Y(mai_mai_n270_));
  OAI210     m254(.A0(mai_mai_n270_), .A1(mai_mai_n264_), .B0(mai_mai_n262_), .Y(mai_mai_n271_));
  NA2        m255(.A(x4), .B(x0), .Y(mai_mai_n272_));
  NA2        m256(.A(mai_mai_n199_), .B(mai_mai_n42_), .Y(mai_mai_n273_));
  AOI210     m257(.A0(mai_mai_n273_), .A1(mai_mai_n271_), .B0(x8), .Y(mai_mai_n274_));
  OAI210     m258(.A0(mai_mai_n258_), .A1(mai_mai_n211_), .B0(x6), .Y(mai_mai_n275_));
  INV        m259(.A(mai_mai_n172_), .Y(mai_mai_n276_));
  OAI210     m260(.A0(mai_mai_n276_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n277_));
  AOI210     m261(.A0(mai_mai_n277_), .A1(mai_mai_n275_), .B0(mai_mai_n226_), .Y(mai_mai_n278_));
  NO4        m262(.A(mai_mai_n278_), .B(mai_mai_n274_), .C(mai_mai_n255_), .D(mai_mai_n243_), .Y(mai_mai_n279_));
  NO2        m263(.A(mai_mai_n161_), .B(x1), .Y(mai_mai_n280_));
  NO3        m264(.A(mai_mai_n280_), .B(x3), .C(mai_mai_n36_), .Y(mai_mai_n281_));
  OAI210     m265(.A0(mai_mai_n281_), .A1(mai_mai_n253_), .B0(x2), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n276_), .A1(x6), .B0(mai_mai_n44_), .Y(mai_mai_n283_));
  AOI210     m267(.A0(mai_mai_n283_), .A1(mai_mai_n282_), .B0(mai_mai_n184_), .Y(mai_mai_n284_));
  NOi21      m268(.An(mai_mai_n267_), .B(mai_mai_n17_), .Y(mai_mai_n285_));
  NA3        m269(.A(mai_mai_n285_), .B(mai_mai_n211_), .C(mai_mai_n40_), .Y(mai_mai_n286_));
  AOI210     m270(.A0(mai_mai_n36_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n287_));
  NA3        m271(.A(mai_mai_n287_), .B(mai_mai_n159_), .C(mai_mai_n32_), .Y(mai_mai_n288_));
  NA2        m272(.A(x3), .B(x2), .Y(mai_mai_n289_));
  AOI220     m273(.A0(mai_mai_n289_), .A1(mai_mai_n226_), .B0(mai_mai_n288_), .B1(mai_mai_n286_), .Y(mai_mai_n290_));
  NAi21      m274(.An(x4), .B(x0), .Y(mai_mai_n291_));
  NO3        m275(.A(mai_mai_n291_), .B(mai_mai_n44_), .C(x2), .Y(mai_mai_n292_));
  OAI210     m276(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n292_), .Y(mai_mai_n293_));
  OAI220     m277(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n294_));
  NO2        m278(.A(x9), .B(x8), .Y(mai_mai_n295_));
  NA3        m279(.A(mai_mai_n295_), .B(mai_mai_n36_), .C(mai_mai_n54_), .Y(mai_mai_n296_));
  OAI210     m280(.A0(mai_mai_n287_), .A1(mai_mai_n285_), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  AOI220     m281(.A0(mai_mai_n297_), .A1(mai_mai_n80_), .B0(mai_mai_n294_), .B1(mai_mai_n31_), .Y(mai_mai_n298_));
  AOI210     m282(.A0(mai_mai_n298_), .A1(mai_mai_n293_), .B0(mai_mai_n25_), .Y(mai_mai_n299_));
  NA3        m283(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n300_));
  OAI210     m284(.A0(mai_mai_n287_), .A1(mai_mai_n285_), .B0(mai_mai_n300_), .Y(mai_mai_n301_));
  INV        m285(.A(mai_mai_n213_), .Y(mai_mai_n302_));
  NA2        m286(.A(mai_mai_n36_), .B(mai_mai_n43_), .Y(mai_mai_n303_));
  OR2        m287(.A(mai_mai_n303_), .B(mai_mai_n272_), .Y(mai_mai_n304_));
  OAI220     m288(.A0(mai_mai_n304_), .A1(mai_mai_n158_), .B0(mai_mai_n229_), .B1(mai_mai_n302_), .Y(mai_mai_n305_));
  AO210      m289(.A0(mai_mai_n301_), .A1(mai_mai_n146_), .B0(mai_mai_n305_), .Y(mai_mai_n306_));
  NO4        m290(.A(mai_mai_n306_), .B(mai_mai_n299_), .C(mai_mai_n290_), .D(mai_mai_n284_), .Y(mai_mai_n307_));
  OAI210     m291(.A0(mai_mai_n279_), .A1(mai_mai_n239_), .B0(mai_mai_n307_), .Y(mai04));
  OAI210     m292(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n309_));
  NA3        m293(.A(mai_mai_n309_), .B(mai_mai_n265_), .C(mai_mai_n83_), .Y(mai_mai_n310_));
  NO2        m294(.A(x2), .B(x1), .Y(mai_mai_n311_));
  OAI210     m295(.A0(mai_mai_n249_), .A1(mai_mai_n311_), .B0(mai_mai_n36_), .Y(mai_mai_n312_));
  NO2        m296(.A(mai_mai_n311_), .B(mai_mai_n291_), .Y(mai_mai_n313_));
  NA2        m297(.A(mai_mai_n313_), .B(mai_mai_n240_), .Y(mai_mai_n314_));
  NO2        m298(.A(mai_mai_n263_), .B(mai_mai_n90_), .Y(mai_mai_n315_));
  NO2        m299(.A(mai_mai_n315_), .B(mai_mai_n36_), .Y(mai_mai_n316_));
  NO2        m300(.A(mai_mai_n289_), .B(mai_mai_n202_), .Y(mai_mai_n317_));
  NA2        m301(.A(x9), .B(x0), .Y(mai_mai_n318_));
  AOI210     m302(.A0(mai_mai_n90_), .A1(mai_mai_n74_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  OAI210     m303(.A0(mai_mai_n319_), .A1(mai_mai_n317_), .B0(mai_mai_n92_), .Y(mai_mai_n320_));
  NA3        m304(.A(mai_mai_n320_), .B(mai_mai_n316_), .C(mai_mai_n314_), .Y(mai_mai_n321_));
  NA2        m305(.A(mai_mai_n321_), .B(mai_mai_n312_), .Y(mai_mai_n322_));
  NO2        m306(.A(mai_mai_n207_), .B(x3), .Y(mai_mai_n323_));
  INV        m307(.A(mai_mai_n323_), .Y(mai_mai_n324_));
  NOi21      m308(.An(mai_mai_n148_), .B(mai_mai_n126_), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n263_), .A1(mai_mai_n300_), .B0(mai_mai_n303_), .Y(mai_mai_n326_));
  AOI210     m310(.A0(mai_mai_n325_), .A1(mai_mai_n63_), .B0(mai_mai_n326_), .Y(mai_mai_n327_));
  NA3        m311(.A(mai_mai_n437_), .B(mai_mai_n327_), .C(mai_mai_n324_), .Y(mai_mai_n328_));
  OAI210     m312(.A0(mai_mai_n110_), .A1(x3), .B0(mai_mai_n292_), .Y(mai_mai_n329_));
  NA2        m313(.A(mai_mai_n329_), .B(mai_mai_n150_), .Y(mai_mai_n330_));
  AOI210     m314(.A0(mai_mai_n328_), .A1(x4), .B0(mai_mai_n330_), .Y(mai_mai_n331_));
  NA3        m315(.A(mai_mai_n313_), .B(mai_mai_n207_), .C(mai_mai_n92_), .Y(mai_mai_n332_));
  NOi21      m316(.An(x4), .B(x0), .Y(mai_mai_n333_));
  XO2        m317(.A(x4), .B(x0), .Y(mai_mai_n334_));
  OAI210     m318(.A0(mai_mai_n334_), .A1(mai_mai_n113_), .B0(mai_mai_n260_), .Y(mai_mai_n335_));
  AOI220     m319(.A0(mai_mai_n335_), .A1(x8), .B0(mai_mai_n333_), .B1(mai_mai_n93_), .Y(mai_mai_n336_));
  AOI210     m320(.A0(mai_mai_n336_), .A1(mai_mai_n332_), .B0(x3), .Y(mai_mai_n337_));
  INV        m321(.A(mai_mai_n93_), .Y(mai_mai_n338_));
  NO2        m322(.A(mai_mai_n92_), .B(x4), .Y(mai_mai_n339_));
  AOI220     m323(.A0(mai_mai_n339_), .A1(mai_mai_n44_), .B0(mai_mai_n121_), .B1(mai_mai_n338_), .Y(mai_mai_n340_));
  NO3        m324(.A(mai_mai_n334_), .B(mai_mai_n161_), .C(x2), .Y(mai_mai_n341_));
  NO3        m325(.A(mai_mai_n223_), .B(mai_mai_n28_), .C(mai_mai_n24_), .Y(mai_mai_n342_));
  NO2        m326(.A(mai_mai_n342_), .B(mai_mai_n341_), .Y(mai_mai_n343_));
  NA4        m327(.A(mai_mai_n343_), .B(mai_mai_n340_), .C(mai_mai_n219_), .D(x6), .Y(mai_mai_n344_));
  OAI220     m328(.A0(mai_mai_n291_), .A1(mai_mai_n90_), .B0(mai_mai_n177_), .B1(mai_mai_n92_), .Y(mai_mai_n345_));
  NO2        m329(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n346_));
  OR2        m330(.A(mai_mai_n339_), .B(mai_mai_n346_), .Y(mai_mai_n347_));
  NO2        m331(.A(mai_mai_n148_), .B(mai_mai_n105_), .Y(mai_mai_n348_));
  AOI220     m332(.A0(mai_mai_n348_), .A1(mai_mai_n347_), .B0(mai_mai_n345_), .B1(mai_mai_n61_), .Y(mai_mai_n349_));
  NO2        m333(.A(mai_mai_n148_), .B(mai_mai_n79_), .Y(mai_mai_n350_));
  NO2        m334(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n351_));
  NOi21      m335(.An(mai_mai_n118_), .B(mai_mai_n27_), .Y(mai_mai_n352_));
  AOI210     m336(.A0(mai_mai_n351_), .A1(mai_mai_n350_), .B0(mai_mai_n352_), .Y(mai_mai_n353_));
  OAI210     m337(.A0(mai_mai_n349_), .A1(mai_mai_n62_), .B0(mai_mai_n353_), .Y(mai_mai_n354_));
  OAI220     m338(.A0(mai_mai_n354_), .A1(x6), .B0(mai_mai_n344_), .B1(mai_mai_n337_), .Y(mai_mai_n355_));
  OAI210     m339(.A0(mai_mai_n63_), .A1(mai_mai_n48_), .B0(mai_mai_n42_), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n356_), .A1(mai_mai_n92_), .B0(mai_mai_n304_), .Y(mai_mai_n357_));
  AOI210     m341(.A0(mai_mai_n357_), .A1(mai_mai_n18_), .B0(mai_mai_n150_), .Y(mai_mai_n358_));
  AO220      m342(.A0(mai_mai_n358_), .A1(mai_mai_n355_), .B0(mai_mai_n331_), .B1(mai_mai_n322_), .Y(mai_mai_n359_));
  NA2        m343(.A(mai_mai_n82_), .B(x6), .Y(mai_mai_n360_));
  INV        m344(.A(mai_mai_n360_), .Y(mai_mai_n361_));
  NA2        m345(.A(mai_mai_n361_), .B(mai_mai_n35_), .Y(mai_mai_n362_));
  NA3        m346(.A(mai_mai_n362_), .B(mai_mai_n359_), .C(mai_mai_n310_), .Y(mai_mai_n363_));
  AOI210     m347(.A0(mai_mai_n195_), .A1(x8), .B0(mai_mai_n110_), .Y(mai_mai_n364_));
  INV        m348(.A(mai_mai_n364_), .Y(mai_mai_n365_));
  NA3        m349(.A(mai_mai_n365_), .B(mai_mai_n192_), .C(mai_mai_n150_), .Y(mai_mai_n366_));
  OAI210     m350(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n226_), .Y(mai_mai_n367_));
  AO220      m351(.A0(mai_mai_n367_), .A1(mai_mai_n147_), .B0(mai_mai_n109_), .B1(x4), .Y(mai_mai_n368_));
  NA3        m352(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n369_));
  NO2        m353(.A(mai_mai_n369_), .B(mai_mai_n338_), .Y(mai_mai_n370_));
  AOI210     m354(.A0(mai_mai_n368_), .A1(mai_mai_n115_), .B0(mai_mai_n370_), .Y(mai_mai_n371_));
  AOI210     m355(.A0(mai_mai_n371_), .A1(mai_mai_n366_), .B0(mai_mai_n25_), .Y(mai_mai_n372_));
  NA3        m356(.A(mai_mai_n117_), .B(mai_mai_n218_), .C(x0), .Y(mai_mai_n373_));
  OAI210     m357(.A0(mai_mai_n192_), .A1(mai_mai_n67_), .B0(mai_mai_n202_), .Y(mai_mai_n374_));
  NA3        m358(.A(mai_mai_n195_), .B(mai_mai_n220_), .C(x8), .Y(mai_mai_n375_));
  AOI210     m359(.A0(mai_mai_n375_), .A1(mai_mai_n374_), .B0(mai_mai_n25_), .Y(mai_mai_n376_));
  AOI210     m360(.A0(mai_mai_n116_), .A1(mai_mai_n114_), .B0(mai_mai_n42_), .Y(mai_mai_n377_));
  NOi31      m361(.An(mai_mai_n377_), .B(mai_mai_n346_), .C(mai_mai_n178_), .Y(mai_mai_n378_));
  OAI210     m362(.A0(mai_mai_n378_), .A1(mai_mai_n376_), .B0(mai_mai_n147_), .Y(mai_mai_n379_));
  NAi31      m363(.An(mai_mai_n50_), .B(mai_mai_n280_), .C(mai_mai_n173_), .Y(mai_mai_n380_));
  NA3        m364(.A(mai_mai_n380_), .B(mai_mai_n379_), .C(mai_mai_n373_), .Y(mai_mai_n381_));
  OAI210     m365(.A0(mai_mai_n381_), .A1(mai_mai_n372_), .B0(x6), .Y(mai_mai_n382_));
  INV        m366(.A(mai_mai_n131_), .Y(mai_mai_n383_));
  NA3        m367(.A(mai_mai_n55_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n384_));
  AOI220     m368(.A0(mai_mai_n384_), .A1(mai_mai_n383_), .B0(mai_mai_n40_), .B1(mai_mai_n32_), .Y(mai_mai_n385_));
  AOI220     m369(.A0(mai_mai_n436_), .A1(mai_mai_n218_), .B0(mai_mai_n192_), .B1(mai_mai_n150_), .Y(mai_mai_n386_));
  AOI210     m370(.A0(mai_mai_n122_), .A1(mai_mai_n244_), .B0(x1), .Y(mai_mai_n387_));
  OAI210     m371(.A0(mai_mai_n386_), .A1(x8), .B0(mai_mai_n387_), .Y(mai_mai_n388_));
  NO4        m372(.A(x8), .B(mai_mai_n291_), .C(x9), .D(x2), .Y(mai_mai_n389_));
  NOi21      m373(.An(mai_mai_n120_), .B(mai_mai_n177_), .Y(mai_mai_n390_));
  NO3        m374(.A(mai_mai_n390_), .B(mai_mai_n389_), .C(mai_mai_n18_), .Y(mai_mai_n391_));
  NO3        m375(.A(x9), .B(mai_mai_n150_), .C(x0), .Y(mai_mai_n392_));
  AOI220     m376(.A0(mai_mai_n392_), .A1(mai_mai_n240_), .B0(mai_mai_n350_), .B1(mai_mai_n150_), .Y(mai_mai_n393_));
  NA3        m377(.A(mai_mai_n393_), .B(mai_mai_n391_), .C(mai_mai_n50_), .Y(mai_mai_n394_));
  OAI210     m378(.A0(mai_mai_n388_), .A1(mai_mai_n385_), .B0(mai_mai_n394_), .Y(mai_mai_n395_));
  NOi31      m379(.An(mai_mai_n436_), .B(mai_mai_n32_), .C(x8), .Y(mai_mai_n396_));
  AOI210     m380(.A0(mai_mai_n38_), .A1(x9), .B0(mai_mai_n129_), .Y(mai_mai_n397_));
  NO3        m381(.A(mai_mai_n397_), .B(mai_mai_n120_), .C(mai_mai_n43_), .Y(mai_mai_n398_));
  NOi31      m382(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n399_));
  AOI220     m383(.A0(mai_mai_n399_), .A1(mai_mai_n333_), .B0(mai_mai_n121_), .B1(x3), .Y(mai_mai_n400_));
  AOI210     m384(.A0(mai_mai_n260_), .A1(mai_mai_n60_), .B0(mai_mai_n119_), .Y(mai_mai_n401_));
  OAI210     m385(.A0(mai_mai_n401_), .A1(x3), .B0(mai_mai_n400_), .Y(mai_mai_n402_));
  NO3        m386(.A(mai_mai_n402_), .B(mai_mai_n398_), .C(x2), .Y(mai_mai_n403_));
  NO2        m387(.A(mai_mai_n403_), .B(mai_mai_n396_), .Y(mai_mai_n404_));
  AOI210     m388(.A0(mai_mai_n404_), .A1(mai_mai_n395_), .B0(mai_mai_n25_), .Y(mai_mai_n405_));
  NO3        m389(.A(mai_mai_n62_), .B(x4), .C(x1), .Y(mai_mai_n406_));
  NA2        m390(.A(mai_mai_n406_), .B(mai_mai_n377_), .Y(mai_mai_n407_));
  NO2        m391(.A(mai_mai_n407_), .B(mai_mai_n104_), .Y(mai_mai_n408_));
  NO3        m392(.A(mai_mai_n263_), .B(mai_mai_n172_), .C(mai_mai_n40_), .Y(mai_mai_n409_));
  OAI210     m393(.A0(mai_mai_n409_), .A1(mai_mai_n408_), .B0(x7), .Y(mai_mai_n410_));
  NA2        m394(.A(mai_mai_n223_), .B(x7), .Y(mai_mai_n411_));
  NA3        m395(.A(mai_mai_n411_), .B(mai_mai_n149_), .C(mai_mai_n130_), .Y(mai_mai_n412_));
  NA2        m396(.A(mai_mai_n412_), .B(mai_mai_n410_), .Y(mai_mai_n413_));
  OAI210     m397(.A0(mai_mai_n413_), .A1(mai_mai_n405_), .B0(mai_mai_n36_), .Y(mai_mai_n414_));
  NO2        m398(.A(mai_mai_n392_), .B(mai_mai_n202_), .Y(mai_mai_n415_));
  NO4        m399(.A(mai_mai_n415_), .B(mai_mai_n76_), .C(x4), .D(mai_mai_n54_), .Y(mai_mai_n416_));
  NO2        m400(.A(mai_mai_n163_), .B(mai_mai_n28_), .Y(mai_mai_n417_));
  AOI220     m401(.A0(mai_mai_n346_), .A1(mai_mai_n92_), .B0(mai_mai_n148_), .B1(mai_mai_n195_), .Y(mai_mai_n418_));
  NA2        m402(.A(mai_mai_n418_), .B(mai_mai_n90_), .Y(mai_mai_n419_));
  NA2        m403(.A(mai_mai_n419_), .B(mai_mai_n173_), .Y(mai_mai_n420_));
  AOI210     m404(.A0(mai_mai_n162_), .A1(mai_mai_n27_), .B0(mai_mai_n71_), .Y(mai_mai_n421_));
  OAI210     m405(.A0(mai_mai_n147_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n422_));
  NO3        m406(.A(mai_mai_n399_), .B(x3), .C(mai_mai_n54_), .Y(mai_mai_n423_));
  AOI210     m407(.A0(mai_mai_n423_), .A1(mai_mai_n422_), .B0(mai_mai_n421_), .Y(mai_mai_n424_));
  INV        m408(.A(mai_mai_n424_), .Y(mai_mai_n425_));
  NA2        m409(.A(mai_mai_n425_), .B(x0), .Y(mai_mai_n426_));
  AOI210     m410(.A0(mai_mai_n426_), .A1(mai_mai_n420_), .B0(mai_mai_n229_), .Y(mai_mai_n427_));
  NA2        m411(.A(x9), .B(x5), .Y(mai_mai_n428_));
  NO4        m412(.A(mai_mai_n105_), .B(mai_mai_n428_), .C(mai_mai_n60_), .D(mai_mai_n32_), .Y(mai_mai_n429_));
  NO4        m413(.A(mai_mai_n429_), .B(mai_mai_n427_), .C(mai_mai_n417_), .D(mai_mai_n416_), .Y(mai_mai_n430_));
  NA3        m414(.A(mai_mai_n430_), .B(mai_mai_n414_), .C(mai_mai_n382_), .Y(mai_mai_n431_));
  AOI210     m415(.A0(mai_mai_n363_), .A1(mai_mai_n25_), .B0(mai_mai_n431_), .Y(mai05));
  INV        m416(.A(x6), .Y(mai_mai_n435_));
  INV        m417(.A(x0), .Y(mai_mai_n436_));
  INV        m418(.A(mai_mai_n77_), .Y(mai_mai_n437_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  AN2        u021(.A(x8), .B(x7), .Y(men_men_n38_));
  NA3        u022(.A(men_men_n38_), .B(men_men_n37_), .C(men_men_n35_), .Y(men_men_n39_));
  NA2        u023(.A(x4), .B(x3), .Y(men_men_n40_));
  AOI210     u024(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n40_), .Y(men_men_n41_));
  NO2        u025(.A(x2), .B(x0), .Y(men_men_n42_));
  INV        u026(.A(x3), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n44_));
  INV        u028(.A(men_men_n44_), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n37_), .B(x4), .Y(men_men_n46_));
  OAI210     u030(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n42_), .Y(men_men_n47_));
  INV        u031(.A(x4), .Y(men_men_n48_));
  NO2        u032(.A(men_men_n48_), .B(men_men_n17_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(x2), .Y(men_men_n50_));
  OAI210     u034(.A0(men_men_n50_), .A1(men_men_n20_), .B0(men_men_n47_), .Y(men_men_n51_));
  NA2        u035(.A(men_men_n38_), .B(men_men_n37_), .Y(men_men_n52_));
  AOI220     u036(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n53_));
  INV        u037(.A(x2), .Y(men_men_n54_));
  NO2        u038(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n56_));
  NA2        u040(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  OAI210     u041(.A0(men_men_n53_), .A1(men_men_n32_), .B0(men_men_n57_), .Y(men_men_n58_));
  NO3        u042(.A(men_men_n58_), .B(men_men_n51_), .C(men_men_n41_), .Y(men01));
  NA2        u043(.A(x8), .B(x7), .Y(men_men_n60_));
  NA2        u044(.A(men_men_n43_), .B(x1), .Y(men_men_n61_));
  INV        u045(.A(x9), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n62_), .B(men_men_n36_), .Y(men_men_n63_));
  INV        u047(.A(men_men_n63_), .Y(men_men_n64_));
  NO3        u048(.A(men_men_n64_), .B(men_men_n61_), .C(men_men_n60_), .Y(men_men_n65_));
  NO2        u049(.A(x7), .B(x6), .Y(men_men_n66_));
  NO2        u050(.A(men_men_n61_), .B(x5), .Y(men_men_n67_));
  NO2        u051(.A(x8), .B(x2), .Y(men_men_n68_));
  INV        u052(.A(men_men_n68_), .Y(men_men_n69_));
  NO2        u053(.A(men_men_n69_), .B(x1), .Y(men_men_n70_));
  OA210      u054(.A0(men_men_n70_), .A1(men_men_n67_), .B0(men_men_n66_), .Y(men_men_n71_));
  OAI210     u055(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n72_));
  OAI210     u056(.A0(men_men_n56_), .A1(men_men_n20_), .B0(men_men_n72_), .Y(men_men_n73_));
  NAi31      u057(.An(x1), .B(x9), .C(x5), .Y(men_men_n74_));
  OAI220     u058(.A0(men_men_n74_), .A1(men_men_n43_), .B0(men_men_n73_), .B1(men_men_n71_), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n65_), .B0(x4), .Y(men_men_n76_));
  NA2        u060(.A(men_men_n48_), .B(x2), .Y(men_men_n77_));
  OAI210     u061(.A0(men_men_n77_), .A1(men_men_n56_), .B0(x0), .Y(men_men_n78_));
  NA2        u062(.A(x5), .B(x3), .Y(men_men_n79_));
  NO2        u063(.A(x8), .B(x6), .Y(men_men_n80_));
  NO4        u064(.A(men_men_n80_), .B(men_men_n79_), .C(men_men_n66_), .D(men_men_n54_), .Y(men_men_n81_));
  NAi21      u065(.An(x4), .B(x3), .Y(men_men_n82_));
  INV        u066(.A(men_men_n82_), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n83_), .B(men_men_n22_), .Y(men_men_n84_));
  NO2        u068(.A(x4), .B(x2), .Y(men_men_n85_));
  NO2        u069(.A(men_men_n85_), .B(x3), .Y(men_men_n86_));
  NO3        u070(.A(men_men_n86_), .B(men_men_n84_), .C(men_men_n18_), .Y(men_men_n87_));
  NO3        u071(.A(men_men_n87_), .B(men_men_n81_), .C(men_men_n78_), .Y(men_men_n88_));
  NO4        u072(.A(men_men_n21_), .B(x6), .C(men_men_n43_), .D(x1), .Y(men_men_n89_));
  NA2        u073(.A(men_men_n62_), .B(men_men_n48_), .Y(men_men_n90_));
  INV        u074(.A(men_men_n90_), .Y(men_men_n91_));
  OAI210     u075(.A0(men_men_n89_), .A1(men_men_n67_), .B0(men_men_n91_), .Y(men_men_n92_));
  NA2        u076(.A(x3), .B(men_men_n18_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n25_), .Y(men_men_n94_));
  INV        u078(.A(x8), .Y(men_men_n95_));
  NA2        u079(.A(x2), .B(x1), .Y(men_men_n96_));
  NO2        u080(.A(men_men_n96_), .B(men_men_n26_), .Y(men_men_n97_));
  AOI210     u081(.A0(men_men_n56_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n98_));
  OAI210     u082(.A0(men_men_n45_), .A1(men_men_n37_), .B0(men_men_n48_), .Y(men_men_n99_));
  NO3        u083(.A(men_men_n99_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n100_));
  NA2        u084(.A(x4), .B(men_men_n43_), .Y(men_men_n101_));
  NO2        u085(.A(men_men_n48_), .B(men_men_n54_), .Y(men_men_n102_));
  AOI210     u086(.A0(men_men_n101_), .A1(men_men_n52_), .B0(x1), .Y(men_men_n103_));
  NO2        u087(.A(x3), .B(x2), .Y(men_men_n104_));
  NA3        u088(.A(men_men_n104_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n105_));
  AOI210     u089(.A0(x8), .A1(x6), .B0(men_men_n105_), .Y(men_men_n106_));
  NA2        u090(.A(men_men_n54_), .B(x1), .Y(men_men_n107_));
  OAI210     u091(.A0(men_men_n107_), .A1(men_men_n40_), .B0(men_men_n17_), .Y(men_men_n108_));
  NO4        u092(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n103_), .D(men_men_n100_), .Y(men_men_n109_));
  AO220      u093(.A0(men_men_n109_), .A1(men_men_n92_), .B0(men_men_n88_), .B1(men_men_n76_), .Y(men02));
  NO2        u094(.A(x3), .B(men_men_n54_), .Y(men_men_n111_));
  NA2        u095(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n43_), .B(x0), .Y(men_men_n113_));
  OAI210     u097(.A0(men_men_n90_), .A1(men_men_n112_), .B0(men_men_n113_), .Y(men_men_n114_));
  AOI220     u098(.A0(men_men_n114_), .A1(x1), .B0(men_men_n111_), .B1(x4), .Y(men_men_n115_));
  NO3        u099(.A(men_men_n115_), .B(x7), .C(x5), .Y(men_men_n116_));
  NA2        u100(.A(x9), .B(x2), .Y(men_men_n117_));
  OR2        u101(.A(x8), .B(x0), .Y(men_men_n118_));
  INV        u102(.A(men_men_n118_), .Y(men_men_n119_));
  NAi21      u103(.An(x2), .B(x8), .Y(men_men_n120_));
  OAI210     u104(.A0(men_men_n117_), .A1(x7), .B0(men_men_n119_), .Y(men_men_n121_));
  NO2        u105(.A(x4), .B(x1), .Y(men_men_n122_));
  NA3        u106(.A(men_men_n122_), .B(men_men_n121_), .C(men_men_n60_), .Y(men_men_n123_));
  NOi21      u107(.An(x0), .B(x1), .Y(men_men_n124_));
  NO3        u108(.A(x9), .B(x8), .C(x7), .Y(men_men_n125_));
  NOi21      u109(.An(x0), .B(x4), .Y(men_men_n126_));
  NAi21      u110(.An(x8), .B(x7), .Y(men_men_n127_));
  NO2        u111(.A(men_men_n127_), .B(men_men_n62_), .Y(men_men_n128_));
  AOI220     u112(.A0(men_men_n128_), .A1(men_men_n126_), .B0(men_men_n125_), .B1(men_men_n124_), .Y(men_men_n129_));
  AOI210     u113(.A0(men_men_n129_), .A1(men_men_n123_), .B0(men_men_n79_), .Y(men_men_n130_));
  NO2        u114(.A(x5), .B(men_men_n48_), .Y(men_men_n131_));
  NA2        u115(.A(x2), .B(men_men_n18_), .Y(men_men_n132_));
  NA2        u116(.A(men_men_n35_), .B(men_men_n131_), .Y(men_men_n133_));
  NAi21      u117(.An(x0), .B(x4), .Y(men_men_n134_));
  NO2        u118(.A(men_men_n134_), .B(x1), .Y(men_men_n135_));
  NO2        u119(.A(x7), .B(x0), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n85_), .B(men_men_n102_), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n137_), .B(x3), .Y(men_men_n138_));
  OAI210     u122(.A0(men_men_n136_), .A1(men_men_n135_), .B0(men_men_n138_), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n21_), .B(men_men_n43_), .Y(men_men_n140_));
  NA2        u124(.A(x5), .B(x0), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n48_), .B(x2), .Y(men_men_n142_));
  NA3        u126(.A(men_men_n142_), .B(men_men_n141_), .C(men_men_n140_), .Y(men_men_n143_));
  NA4        u127(.A(men_men_n143_), .B(men_men_n139_), .C(men_men_n133_), .D(men_men_n36_), .Y(men_men_n144_));
  NO3        u128(.A(men_men_n144_), .B(men_men_n130_), .C(men_men_n116_), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n146_));
  AOI220     u130(.A0(men_men_n124_), .A1(men_men_n146_), .B0(men_men_n67_), .B1(men_men_n17_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n147_), .B(men_men_n60_), .C(men_men_n62_), .Y(men_men_n148_));
  NA2        u132(.A(x7), .B(x3), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n101_), .B(x5), .Y(men_men_n150_));
  NO2        u134(.A(x9), .B(x7), .Y(men_men_n151_));
  NOi21      u135(.An(x8), .B(x0), .Y(men_men_n152_));
  OA210      u136(.A0(men_men_n151_), .A1(x1), .B0(men_men_n152_), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n43_), .B(x2), .Y(men_men_n154_));
  INV        u138(.A(x7), .Y(men_men_n155_));
  NA2        u139(.A(men_men_n155_), .B(men_men_n18_), .Y(men_men_n156_));
  AOI220     u140(.A0(men_men_n156_), .A1(men_men_n154_), .B0(men_men_n111_), .B1(men_men_n38_), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n25_), .B(x4), .Y(men_men_n158_));
  NO2        u142(.A(men_men_n158_), .B(men_men_n126_), .Y(men_men_n159_));
  NO2        u143(.A(men_men_n159_), .B(men_men_n157_), .Y(men_men_n160_));
  AOI210     u144(.A0(men_men_n153_), .A1(men_men_n150_), .B0(men_men_n160_), .Y(men_men_n161_));
  OAI210     u145(.A0(men_men_n149_), .A1(men_men_n50_), .B0(men_men_n161_), .Y(men_men_n162_));
  NA2        u146(.A(x5), .B(x1), .Y(men_men_n163_));
  INV        u147(.A(men_men_n163_), .Y(men_men_n164_));
  AOI210     u148(.A0(men_men_n164_), .A1(men_men_n126_), .B0(men_men_n36_), .Y(men_men_n165_));
  NO2        u149(.A(men_men_n62_), .B(men_men_n95_), .Y(men_men_n166_));
  NAi21      u150(.An(x2), .B(x7), .Y(men_men_n167_));
  NO3        u151(.A(men_men_n167_), .B(men_men_n166_), .C(men_men_n48_), .Y(men_men_n168_));
  NA2        u152(.A(men_men_n168_), .B(men_men_n67_), .Y(men_men_n169_));
  NAi31      u153(.An(men_men_n79_), .B(men_men_n38_), .C(men_men_n35_), .Y(men_men_n170_));
  NA3        u154(.A(men_men_n170_), .B(men_men_n169_), .C(men_men_n165_), .Y(men_men_n171_));
  NO3        u155(.A(men_men_n171_), .B(men_men_n162_), .C(men_men_n148_), .Y(men_men_n172_));
  NO2        u156(.A(men_men_n172_), .B(men_men_n145_), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n141_), .B(men_men_n137_), .Y(men_men_n174_));
  NA2        u158(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n175_));
  NA2        u159(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n176_));
  NA3        u160(.A(men_men_n176_), .B(men_men_n175_), .C(men_men_n24_), .Y(men_men_n177_));
  AN2        u161(.A(men_men_n177_), .B(men_men_n142_), .Y(men_men_n178_));
  NA2        u162(.A(x8), .B(x0), .Y(men_men_n179_));
  NO2        u163(.A(men_men_n155_), .B(men_men_n25_), .Y(men_men_n180_));
  NO2        u164(.A(men_men_n124_), .B(x4), .Y(men_men_n181_));
  NA2        u165(.A(men_men_n181_), .B(men_men_n180_), .Y(men_men_n182_));
  AOI210     u166(.A0(men_men_n179_), .A1(men_men_n132_), .B0(men_men_n182_), .Y(men_men_n183_));
  NA2        u167(.A(x2), .B(x0), .Y(men_men_n184_));
  NA2        u168(.A(x4), .B(x1), .Y(men_men_n185_));
  NAi21      u169(.An(men_men_n122_), .B(men_men_n185_), .Y(men_men_n186_));
  NOi31      u170(.An(men_men_n186_), .B(men_men_n158_), .C(men_men_n184_), .Y(men_men_n187_));
  NO4        u171(.A(men_men_n187_), .B(men_men_n183_), .C(men_men_n178_), .D(men_men_n174_), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n188_), .B(men_men_n43_), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n177_), .B(men_men_n77_), .Y(men_men_n190_));
  INV        u174(.A(men_men_n131_), .Y(men_men_n191_));
  NO2        u175(.A(men_men_n107_), .B(men_men_n17_), .Y(men_men_n192_));
  AOI210     u176(.A0(men_men_n35_), .A1(men_men_n95_), .B0(men_men_n192_), .Y(men_men_n193_));
  NO3        u177(.A(men_men_n193_), .B(men_men_n191_), .C(x7), .Y(men_men_n194_));
  NA3        u178(.A(men_men_n186_), .B(men_men_n191_), .C(men_men_n42_), .Y(men_men_n195_));
  OAI210     u179(.A0(men_men_n176_), .A1(men_men_n137_), .B0(men_men_n195_), .Y(men_men_n196_));
  NO3        u180(.A(men_men_n196_), .B(men_men_n194_), .C(men_men_n190_), .Y(men_men_n197_));
  NO2        u181(.A(men_men_n197_), .B(x3), .Y(men_men_n198_));
  NO3        u182(.A(men_men_n198_), .B(men_men_n189_), .C(men_men_n173_), .Y(men03));
  NO2        u183(.A(men_men_n48_), .B(x3), .Y(men_men_n200_));
  NO2        u184(.A(x6), .B(men_men_n25_), .Y(men_men_n201_));
  INV        u185(.A(men_men_n63_), .Y(men_men_n202_));
  OAI220     u186(.A0(men_men_n202_), .A1(men_men_n17_), .B0(x6), .B1(men_men_n107_), .Y(men_men_n203_));
  NA2        u187(.A(men_men_n203_), .B(men_men_n200_), .Y(men_men_n204_));
  NO2        u188(.A(men_men_n79_), .B(x6), .Y(men_men_n205_));
  NA2        u189(.A(x6), .B(men_men_n25_), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n206_), .B(x4), .Y(men_men_n207_));
  NO2        u191(.A(men_men_n18_), .B(x0), .Y(men_men_n208_));
  NA2        u192(.A(men_men_n205_), .B(men_men_n62_), .Y(men_men_n209_));
  NA2        u193(.A(x3), .B(men_men_n17_), .Y(men_men_n210_));
  NO2        u194(.A(men_men_n210_), .B(men_men_n206_), .Y(men_men_n211_));
  NA2        u195(.A(x9), .B(men_men_n54_), .Y(men_men_n212_));
  NA2        u196(.A(men_men_n212_), .B(x4), .Y(men_men_n213_));
  NA2        u197(.A(men_men_n206_), .B(men_men_n82_), .Y(men_men_n214_));
  AOI210     u198(.A0(men_men_n25_), .A1(x3), .B0(men_men_n184_), .Y(men_men_n215_));
  AOI220     u199(.A0(men_men_n215_), .A1(men_men_n214_), .B0(men_men_n213_), .B1(men_men_n211_), .Y(men_men_n216_));
  NO3        u200(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n217_));
  NO2        u201(.A(x5), .B(x1), .Y(men_men_n218_));
  AOI220     u202(.A0(men_men_n218_), .A1(men_men_n17_), .B0(men_men_n104_), .B1(x5), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n210_), .B(men_men_n175_), .Y(men_men_n220_));
  NO3        u204(.A(x3), .B(x2), .C(x1), .Y(men_men_n221_));
  NO2        u205(.A(men_men_n221_), .B(men_men_n220_), .Y(men_men_n222_));
  OAI210     u206(.A0(men_men_n219_), .A1(men_men_n64_), .B0(men_men_n222_), .Y(men_men_n223_));
  AOI220     u207(.A0(men_men_n223_), .A1(men_men_n48_), .B0(men_men_n217_), .B1(men_men_n131_), .Y(men_men_n224_));
  NA4        u208(.A(men_men_n224_), .B(men_men_n216_), .C(men_men_n209_), .D(men_men_n204_), .Y(men_men_n225_));
  NO2        u209(.A(men_men_n48_), .B(men_men_n43_), .Y(men_men_n226_));
  NA2        u210(.A(men_men_n226_), .B(men_men_n19_), .Y(men_men_n227_));
  NO2        u211(.A(x3), .B(men_men_n17_), .Y(men_men_n228_));
  NO2        u212(.A(men_men_n228_), .B(x6), .Y(men_men_n229_));
  NOi21      u213(.An(men_men_n85_), .B(men_men_n229_), .Y(men_men_n230_));
  NA2        u214(.A(men_men_n62_), .B(men_men_n95_), .Y(men_men_n231_));
  NA3        u215(.A(men_men_n231_), .B(men_men_n228_), .C(x6), .Y(men_men_n232_));
  AOI210     u216(.A0(men_men_n232_), .A1(men_men_n230_), .B0(men_men_n155_), .Y(men_men_n233_));
  AO210      u217(.A0(men_men_n233_), .A1(men_men_n227_), .B0(men_men_n180_), .Y(men_men_n234_));
  NA2        u218(.A(men_men_n43_), .B(men_men_n54_), .Y(men_men_n235_));
  OAI210     u219(.A0(men_men_n235_), .A1(men_men_n25_), .B0(men_men_n176_), .Y(men_men_n236_));
  NO3        u220(.A(men_men_n185_), .B(men_men_n62_), .C(x6), .Y(men_men_n237_));
  AOI220     u221(.A0(men_men_n237_), .A1(men_men_n236_), .B0(men_men_n142_), .B1(men_men_n94_), .Y(men_men_n238_));
  NA2        u222(.A(x6), .B(men_men_n48_), .Y(men_men_n239_));
  OAI210     u223(.A0(men_men_n119_), .A1(men_men_n80_), .B0(x4), .Y(men_men_n240_));
  AOI210     u224(.A0(men_men_n240_), .A1(men_men_n239_), .B0(men_men_n79_), .Y(men_men_n241_));
  NO2        u225(.A(men_men_n62_), .B(x6), .Y(men_men_n242_));
  NO2        u226(.A(men_men_n163_), .B(men_men_n43_), .Y(men_men_n243_));
  OAI210     u227(.A0(men_men_n243_), .A1(men_men_n220_), .B0(men_men_n242_), .Y(men_men_n244_));
  NA2        u228(.A(men_men_n201_), .B(men_men_n135_), .Y(men_men_n245_));
  NA3        u229(.A(men_men_n210_), .B(men_men_n131_), .C(x6), .Y(men_men_n246_));
  OAI210     u230(.A0(men_men_n95_), .A1(men_men_n36_), .B0(men_men_n67_), .Y(men_men_n247_));
  NA4        u231(.A(men_men_n247_), .B(men_men_n246_), .C(men_men_n245_), .D(men_men_n244_), .Y(men_men_n248_));
  OAI210     u232(.A0(men_men_n248_), .A1(men_men_n241_), .B0(x2), .Y(men_men_n249_));
  NA3        u233(.A(men_men_n249_), .B(men_men_n238_), .C(men_men_n234_), .Y(men_men_n250_));
  AOI210     u234(.A0(men_men_n225_), .A1(x8), .B0(men_men_n250_), .Y(men_men_n251_));
  NO2        u235(.A(men_men_n95_), .B(x3), .Y(men_men_n252_));
  NA2        u236(.A(men_men_n252_), .B(men_men_n207_), .Y(men_men_n253_));
  NO3        u237(.A(men_men_n93_), .B(men_men_n80_), .C(men_men_n25_), .Y(men_men_n254_));
  AOI210     u238(.A0(men_men_n229_), .A1(men_men_n158_), .B0(men_men_n254_), .Y(men_men_n255_));
  AOI210     u239(.A0(men_men_n255_), .A1(men_men_n253_), .B0(x2), .Y(men_men_n256_));
  NO2        u240(.A(x4), .B(men_men_n54_), .Y(men_men_n257_));
  AOI220     u241(.A0(men_men_n207_), .A1(men_men_n192_), .B0(men_men_n257_), .B1(men_men_n67_), .Y(men_men_n258_));
  NA2        u242(.A(men_men_n62_), .B(x6), .Y(men_men_n259_));
  NA3        u243(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n260_));
  AOI210     u244(.A0(men_men_n260_), .A1(men_men_n141_), .B0(men_men_n259_), .Y(men_men_n261_));
  NA2        u245(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n262_));
  NA2        u246(.A(men_men_n261_), .B(men_men_n122_), .Y(men_men_n263_));
  NA2        u247(.A(men_men_n210_), .B(x6), .Y(men_men_n264_));
  NO2        u248(.A(men_men_n210_), .B(x6), .Y(men_men_n265_));
  NAi21      u249(.An(men_men_n166_), .B(men_men_n265_), .Y(men_men_n266_));
  NA3        u250(.A(men_men_n266_), .B(men_men_n264_), .C(men_men_n146_), .Y(men_men_n267_));
  NA4        u251(.A(men_men_n267_), .B(men_men_n263_), .C(men_men_n258_), .D(men_men_n155_), .Y(men_men_n268_));
  NA2        u252(.A(men_men_n201_), .B(men_men_n228_), .Y(men_men_n269_));
  NO2        u253(.A(x9), .B(x6), .Y(men_men_n270_));
  NO2        u254(.A(men_men_n141_), .B(men_men_n18_), .Y(men_men_n271_));
  NAi21      u255(.An(men_men_n271_), .B(men_men_n260_), .Y(men_men_n272_));
  NAi21      u256(.An(x1), .B(x4), .Y(men_men_n273_));
  AOI210     u257(.A0(x3), .A1(x2), .B0(men_men_n48_), .Y(men_men_n274_));
  OAI210     u258(.A0(men_men_n141_), .A1(x3), .B0(men_men_n274_), .Y(men_men_n275_));
  AOI220     u259(.A0(men_men_n275_), .A1(men_men_n273_), .B0(men_men_n272_), .B1(men_men_n270_), .Y(men_men_n276_));
  INV        u260(.A(men_men_n276_), .Y(men_men_n277_));
  NA2        u261(.A(men_men_n62_), .B(x2), .Y(men_men_n278_));
  NO2        u262(.A(men_men_n278_), .B(men_men_n269_), .Y(men_men_n279_));
  NO3        u263(.A(x9), .B(x6), .C(x0), .Y(men_men_n280_));
  NA2        u264(.A(x6), .B(x2), .Y(men_men_n281_));
  NO2        u265(.A(men_men_n281_), .B(men_men_n175_), .Y(men_men_n282_));
  NO2        u266(.A(men_men_n280_), .B(men_men_n282_), .Y(men_men_n283_));
  OAI220     u267(.A0(men_men_n283_), .A1(men_men_n43_), .B0(men_men_n181_), .B1(men_men_n46_), .Y(men_men_n284_));
  OAI210     u268(.A0(men_men_n284_), .A1(men_men_n279_), .B0(men_men_n277_), .Y(men_men_n285_));
  NA2        u269(.A(x9), .B(men_men_n43_), .Y(men_men_n286_));
  NO2        u270(.A(men_men_n286_), .B(men_men_n206_), .Y(men_men_n287_));
  OR3        u271(.A(men_men_n287_), .B(men_men_n205_), .C(men_men_n150_), .Y(men_men_n288_));
  NA2        u272(.A(x4), .B(x0), .Y(men_men_n289_));
  NO3        u273(.A(men_men_n74_), .B(men_men_n289_), .C(x6), .Y(men_men_n290_));
  AOI210     u274(.A0(men_men_n288_), .A1(men_men_n42_), .B0(men_men_n290_), .Y(men_men_n291_));
  AOI210     u275(.A0(men_men_n291_), .A1(men_men_n285_), .B0(x8), .Y(men_men_n292_));
  INV        u276(.A(men_men_n259_), .Y(men_men_n293_));
  OAI210     u277(.A0(men_men_n271_), .A1(men_men_n218_), .B0(men_men_n293_), .Y(men_men_n294_));
  INV        u278(.A(men_men_n179_), .Y(men_men_n295_));
  NO2        u279(.A(men_men_n294_), .B(men_men_n235_), .Y(men_men_n296_));
  NO4        u280(.A(men_men_n296_), .B(men_men_n292_), .C(men_men_n268_), .D(men_men_n256_), .Y(men_men_n297_));
  NO2        u281(.A(men_men_n166_), .B(x1), .Y(men_men_n298_));
  NO3        u282(.A(men_men_n298_), .B(x3), .C(men_men_n36_), .Y(men_men_n299_));
  OAI210     u283(.A0(men_men_n299_), .A1(men_men_n265_), .B0(x2), .Y(men_men_n300_));
  OAI210     u284(.A0(men_men_n295_), .A1(x6), .B0(men_men_n44_), .Y(men_men_n301_));
  AOI210     u285(.A0(men_men_n301_), .A1(men_men_n300_), .B0(men_men_n191_), .Y(men_men_n302_));
  NOi21      u286(.An(men_men_n281_), .B(men_men_n17_), .Y(men_men_n303_));
  NA3        u287(.A(men_men_n303_), .B(men_men_n218_), .C(men_men_n40_), .Y(men_men_n304_));
  AOI210     u288(.A0(men_men_n36_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n305_));
  NA3        u289(.A(men_men_n305_), .B(men_men_n164_), .C(men_men_n32_), .Y(men_men_n306_));
  NA2        u290(.A(x3), .B(x2), .Y(men_men_n307_));
  AOI220     u291(.A0(men_men_n307_), .A1(men_men_n235_), .B0(men_men_n306_), .B1(men_men_n304_), .Y(men_men_n308_));
  NAi21      u292(.An(x4), .B(x0), .Y(men_men_n309_));
  NO3        u293(.A(men_men_n309_), .B(men_men_n44_), .C(x2), .Y(men_men_n310_));
  OAI210     u294(.A0(x6), .A1(men_men_n18_), .B0(men_men_n310_), .Y(men_men_n311_));
  NO2        u295(.A(x9), .B(x8), .Y(men_men_n312_));
  NA3        u296(.A(men_men_n312_), .B(men_men_n36_), .C(men_men_n54_), .Y(men_men_n313_));
  OAI210     u297(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n313_), .Y(men_men_n314_));
  AOI220     u298(.A0(men_men_n314_), .A1(men_men_n83_), .B0(men_men_n18_), .B1(men_men_n31_), .Y(men_men_n315_));
  AOI210     u299(.A0(men_men_n315_), .A1(men_men_n311_), .B0(men_men_n25_), .Y(men_men_n316_));
  NA3        u300(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n317_));
  OAI210     u301(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n317_), .Y(men_men_n318_));
  INV        u302(.A(men_men_n220_), .Y(men_men_n319_));
  NO2        u303(.A(men_men_n239_), .B(men_men_n319_), .Y(men_men_n320_));
  AO210      u304(.A0(men_men_n318_), .A1(men_men_n150_), .B0(men_men_n320_), .Y(men_men_n321_));
  NO4        u305(.A(men_men_n321_), .B(men_men_n316_), .C(men_men_n308_), .D(men_men_n302_), .Y(men_men_n322_));
  OAI210     u306(.A0(men_men_n297_), .A1(men_men_n251_), .B0(men_men_n322_), .Y(men04));
  OAI210     u307(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n324_));
  NA3        u308(.A(men_men_n324_), .B(men_men_n280_), .C(men_men_n86_), .Y(men_men_n325_));
  NO2        u309(.A(x2), .B(x1), .Y(men_men_n326_));
  OAI210     u310(.A0(men_men_n262_), .A1(men_men_n326_), .B0(men_men_n36_), .Y(men_men_n327_));
  AOI210     u311(.A0(men_men_n62_), .A1(x4), .B0(men_men_n112_), .Y(men_men_n328_));
  NA2        u312(.A(men_men_n328_), .B(men_men_n252_), .Y(men_men_n329_));
  NO2        u313(.A(men_men_n278_), .B(men_men_n93_), .Y(men_men_n330_));
  NO2        u314(.A(men_men_n330_), .B(men_men_n36_), .Y(men_men_n331_));
  NO2        u315(.A(men_men_n307_), .B(men_men_n208_), .Y(men_men_n332_));
  NA2        u316(.A(x9), .B(x0), .Y(men_men_n333_));
  AOI210     u317(.A0(men_men_n93_), .A1(men_men_n77_), .B0(men_men_n333_), .Y(men_men_n334_));
  OAI210     u318(.A0(men_men_n334_), .A1(men_men_n332_), .B0(men_men_n95_), .Y(men_men_n335_));
  NA3        u319(.A(men_men_n335_), .B(men_men_n331_), .C(men_men_n329_), .Y(men_men_n336_));
  NA2        u320(.A(men_men_n336_), .B(men_men_n327_), .Y(men_men_n337_));
  NO2        u321(.A(men_men_n212_), .B(men_men_n113_), .Y(men_men_n338_));
  NO3        u322(.A(men_men_n259_), .B(men_men_n120_), .C(men_men_n18_), .Y(men_men_n339_));
  NO2        u323(.A(men_men_n339_), .B(men_men_n338_), .Y(men_men_n340_));
  OAI210     u324(.A0(men_men_n118_), .A1(men_men_n107_), .B0(men_men_n179_), .Y(men_men_n341_));
  NA3        u325(.A(men_men_n341_), .B(x6), .C(x3), .Y(men_men_n342_));
  NOi21      u326(.An(men_men_n152_), .B(men_men_n132_), .Y(men_men_n343_));
  NO2        u327(.A(men_men_n278_), .B(men_men_n317_), .Y(men_men_n344_));
  AOI210     u328(.A0(men_men_n343_), .A1(men_men_n63_), .B0(men_men_n344_), .Y(men_men_n345_));
  NA2        u329(.A(x2), .B(men_men_n17_), .Y(men_men_n346_));
  OAI210     u330(.A0(men_men_n107_), .A1(men_men_n17_), .B0(men_men_n346_), .Y(men_men_n347_));
  AOI220     u331(.A0(men_men_n347_), .A1(men_men_n80_), .B0(men_men_n330_), .B1(men_men_n95_), .Y(men_men_n348_));
  NA4        u332(.A(men_men_n348_), .B(men_men_n345_), .C(men_men_n342_), .D(men_men_n340_), .Y(men_men_n349_));
  OAI210     u333(.A0(x1), .A1(x3), .B0(men_men_n310_), .Y(men_men_n350_));
  NA3        u334(.A(men_men_n231_), .B(men_men_n217_), .C(men_men_n85_), .Y(men_men_n351_));
  NA3        u335(.A(men_men_n351_), .B(men_men_n350_), .C(men_men_n155_), .Y(men_men_n352_));
  AOI210     u336(.A0(men_men_n349_), .A1(x4), .B0(men_men_n352_), .Y(men_men_n353_));
  NOi21      u337(.An(x4), .B(x0), .Y(men_men_n354_));
  XO2        u338(.A(x4), .B(x0), .Y(men_men_n355_));
  AOI220     u339(.A0(x2), .A1(x8), .B0(men_men_n354_), .B1(men_men_n96_), .Y(men_men_n356_));
  AOI210     u340(.A0(men_men_n356_), .A1(men_men_n309_), .B0(x3), .Y(men_men_n357_));
  NO2        u341(.A(men_men_n95_), .B(x4), .Y(men_men_n358_));
  NA2        u342(.A(men_men_n358_), .B(men_men_n44_), .Y(men_men_n359_));
  NO3        u343(.A(men_men_n355_), .B(men_men_n166_), .C(x2), .Y(men_men_n360_));
  NO3        u344(.A(men_men_n231_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n361_));
  NO2        u345(.A(men_men_n361_), .B(men_men_n360_), .Y(men_men_n362_));
  NA4        u346(.A(men_men_n362_), .B(men_men_n359_), .C(men_men_n227_), .D(x6), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n152_), .B(men_men_n107_), .Y(men_men_n364_));
  AOI210     u348(.A0(men_men_n462_), .A1(men_men_n61_), .B0(men_men_n364_), .Y(men_men_n365_));
  NO2        u349(.A(men_men_n152_), .B(men_men_n82_), .Y(men_men_n366_));
  NO2        u350(.A(men_men_n35_), .B(x2), .Y(men_men_n367_));
  NOi21      u351(.An(men_men_n122_), .B(men_men_n27_), .Y(men_men_n368_));
  AOI210     u352(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n368_), .Y(men_men_n369_));
  OAI210     u353(.A0(men_men_n365_), .A1(men_men_n62_), .B0(men_men_n369_), .Y(men_men_n370_));
  OAI220     u354(.A0(men_men_n370_), .A1(x6), .B0(men_men_n363_), .B1(men_men_n357_), .Y(men_men_n371_));
  OAI210     u355(.A0(men_men_n63_), .A1(men_men_n48_), .B0(men_men_n42_), .Y(men_men_n372_));
  NO2        u356(.A(men_men_n372_), .B(men_men_n95_), .Y(men_men_n373_));
  AOI210     u357(.A0(men_men_n373_), .A1(men_men_n18_), .B0(men_men_n155_), .Y(men_men_n374_));
  AO220      u358(.A0(men_men_n374_), .A1(men_men_n371_), .B0(men_men_n353_), .B1(men_men_n337_), .Y(men_men_n375_));
  NA2        u359(.A(men_men_n367_), .B(x6), .Y(men_men_n376_));
  AOI210     u360(.A0(x6), .A1(x1), .B0(men_men_n154_), .Y(men_men_n377_));
  NA2        u361(.A(men_men_n358_), .B(x0), .Y(men_men_n378_));
  NA2        u362(.A(men_men_n85_), .B(x6), .Y(men_men_n379_));
  OAI210     u363(.A0(men_men_n378_), .A1(men_men_n377_), .B0(men_men_n379_), .Y(men_men_n380_));
  AOI220     u364(.A0(men_men_n380_), .A1(men_men_n376_), .B0(men_men_n221_), .B1(men_men_n49_), .Y(men_men_n381_));
  NA3        u365(.A(men_men_n381_), .B(men_men_n375_), .C(men_men_n325_), .Y(men_men_n382_));
  NA3        u366(.A(x2), .B(men_men_n200_), .C(men_men_n155_), .Y(men_men_n383_));
  AO220      u367(.A0(x4), .A1(men_men_n151_), .B0(men_men_n111_), .B1(x4), .Y(men_men_n384_));
  NA3        u368(.A(x7), .B(x3), .C(x0), .Y(men_men_n385_));
  NA2        u369(.A(men_men_n226_), .B(x0), .Y(men_men_n386_));
  NO2        u370(.A(men_men_n386_), .B(men_men_n212_), .Y(men_men_n387_));
  AOI210     u371(.A0(men_men_n384_), .A1(men_men_n119_), .B0(men_men_n387_), .Y(men_men_n388_));
  AOI210     u372(.A0(men_men_n388_), .A1(men_men_n383_), .B0(men_men_n25_), .Y(men_men_n389_));
  OAI210     u373(.A0(men_men_n200_), .A1(men_men_n68_), .B0(men_men_n208_), .Y(men_men_n390_));
  NA3        u374(.A(x2), .B(men_men_n228_), .C(x8), .Y(men_men_n391_));
  AOI210     u375(.A0(men_men_n391_), .A1(men_men_n390_), .B0(men_men_n25_), .Y(men_men_n392_));
  AOI210     u376(.A0(men_men_n120_), .A1(men_men_n118_), .B0(men_men_n42_), .Y(men_men_n393_));
  NOi31      u377(.An(men_men_n393_), .B(x3), .C(men_men_n185_), .Y(men_men_n394_));
  OAI210     u378(.A0(men_men_n394_), .A1(men_men_n392_), .B0(men_men_n151_), .Y(men_men_n395_));
  NAi31      u379(.An(men_men_n50_), .B(men_men_n298_), .C(men_men_n180_), .Y(men_men_n396_));
  NA2        u380(.A(men_men_n396_), .B(men_men_n395_), .Y(men_men_n397_));
  OAI210     u381(.A0(men_men_n397_), .A1(men_men_n389_), .B0(x6), .Y(men_men_n398_));
  OAI210     u382(.A0(men_men_n166_), .A1(men_men_n48_), .B0(men_men_n136_), .Y(men_men_n399_));
  NA3        u383(.A(men_men_n55_), .B(men_men_n38_), .C(men_men_n31_), .Y(men_men_n400_));
  AOI220     u384(.A0(men_men_n400_), .A1(men_men_n399_), .B0(men_men_n40_), .B1(men_men_n32_), .Y(men_men_n401_));
  NO2        u385(.A(men_men_n155_), .B(x0), .Y(men_men_n402_));
  AOI220     u386(.A0(men_men_n402_), .A1(men_men_n226_), .B0(men_men_n200_), .B1(men_men_n155_), .Y(men_men_n403_));
  AOI210     u387(.A0(men_men_n128_), .A1(men_men_n257_), .B0(x1), .Y(men_men_n404_));
  OAI210     u388(.A0(men_men_n403_), .A1(x8), .B0(men_men_n404_), .Y(men_men_n405_));
  NAi31      u389(.An(x2), .B(x8), .C(x0), .Y(men_men_n406_));
  OAI210     u390(.A0(men_men_n406_), .A1(x4), .B0(men_men_n167_), .Y(men_men_n407_));
  NA3        u391(.A(men_men_n407_), .B(men_men_n149_), .C(x9), .Y(men_men_n408_));
  NO4        u392(.A(men_men_n127_), .B(men_men_n309_), .C(x9), .D(x2), .Y(men_men_n409_));
  NOi21      u393(.An(men_men_n125_), .B(men_men_n184_), .Y(men_men_n410_));
  NO3        u394(.A(men_men_n410_), .B(men_men_n409_), .C(men_men_n18_), .Y(men_men_n411_));
  NO3        u395(.A(x9), .B(men_men_n155_), .C(x0), .Y(men_men_n412_));
  AOI220     u396(.A0(men_men_n412_), .A1(men_men_n252_), .B0(men_men_n366_), .B1(men_men_n155_), .Y(men_men_n413_));
  NA3        u397(.A(men_men_n413_), .B(men_men_n411_), .C(men_men_n408_), .Y(men_men_n414_));
  OAI210     u398(.A0(men_men_n405_), .A1(men_men_n401_), .B0(men_men_n414_), .Y(men_men_n415_));
  NOi31      u399(.An(men_men_n402_), .B(men_men_n32_), .C(x8), .Y(men_men_n416_));
  NO2        u400(.A(men_men_n125_), .B(men_men_n43_), .Y(men_men_n417_));
  NOi31      u401(.An(x1), .B(x8), .C(x7), .Y(men_men_n418_));
  AOI210     u402(.A0(men_men_n126_), .A1(x3), .B0(men_men_n354_), .Y(men_men_n419_));
  NA2        u403(.A(x3), .B(men_men_n419_), .Y(men_men_n420_));
  NO3        u404(.A(men_men_n420_), .B(men_men_n417_), .C(x2), .Y(men_men_n421_));
  OAI220     u405(.A0(men_men_n355_), .A1(men_men_n312_), .B0(men_men_n309_), .B1(men_men_n43_), .Y(men_men_n422_));
  AOI210     u406(.A0(x9), .A1(men_men_n48_), .B0(men_men_n385_), .Y(men_men_n423_));
  AOI220     u407(.A0(men_men_n423_), .A1(men_men_n95_), .B0(men_men_n422_), .B1(men_men_n155_), .Y(men_men_n424_));
  NO2        u408(.A(men_men_n424_), .B(men_men_n54_), .Y(men_men_n425_));
  NO3        u409(.A(men_men_n425_), .B(men_men_n421_), .C(men_men_n416_), .Y(men_men_n426_));
  AOI210     u410(.A0(men_men_n426_), .A1(men_men_n415_), .B0(men_men_n25_), .Y(men_men_n427_));
  NA4        u411(.A(men_men_n31_), .B(men_men_n95_), .C(x2), .D(men_men_n17_), .Y(men_men_n428_));
  NO3        u412(.A(men_men_n62_), .B(x4), .C(x1), .Y(men_men_n429_));
  NO3        u413(.A(men_men_n68_), .B(men_men_n18_), .C(x0), .Y(men_men_n430_));
  AOI220     u414(.A0(men_men_n430_), .A1(men_men_n274_), .B0(men_men_n429_), .B1(men_men_n393_), .Y(men_men_n431_));
  NO2        u415(.A(men_men_n431_), .B(men_men_n104_), .Y(men_men_n432_));
  NO3        u416(.A(men_men_n278_), .B(men_men_n179_), .C(men_men_n40_), .Y(men_men_n433_));
  OAI210     u417(.A0(men_men_n433_), .A1(men_men_n432_), .B0(x7), .Y(men_men_n434_));
  NA3        u418(.A(men_men_n62_), .B(men_men_n154_), .C(men_men_n135_), .Y(men_men_n435_));
  NA3        u419(.A(men_men_n435_), .B(men_men_n434_), .C(men_men_n428_), .Y(men_men_n436_));
  OAI210     u420(.A0(men_men_n436_), .A1(men_men_n427_), .B0(men_men_n36_), .Y(men_men_n437_));
  NO2        u421(.A(men_men_n412_), .B(men_men_n208_), .Y(men_men_n438_));
  NO4        u422(.A(men_men_n438_), .B(men_men_n79_), .C(x4), .D(men_men_n54_), .Y(men_men_n439_));
  NA2        u423(.A(men_men_n262_), .B(men_men_n21_), .Y(men_men_n440_));
  NO2        u424(.A(men_men_n163_), .B(men_men_n136_), .Y(men_men_n441_));
  NA2        u425(.A(men_men_n441_), .B(men_men_n440_), .Y(men_men_n442_));
  AOI210     u426(.A0(men_men_n442_), .A1(men_men_n170_), .B0(men_men_n28_), .Y(men_men_n443_));
  AOI220     u427(.A0(x3), .A1(men_men_n95_), .B0(men_men_n152_), .B1(x2), .Y(men_men_n444_));
  NA3        u428(.A(men_men_n444_), .B(men_men_n406_), .C(men_men_n93_), .Y(men_men_n445_));
  NA2        u429(.A(men_men_n445_), .B(men_men_n180_), .Y(men_men_n446_));
  OAI220     u430(.A0(men_men_n286_), .A1(men_men_n69_), .B0(men_men_n163_), .B1(men_men_n43_), .Y(men_men_n447_));
  NA2        u431(.A(x3), .B(men_men_n54_), .Y(men_men_n448_));
  AOI210     u432(.A0(men_men_n167_), .A1(men_men_n27_), .B0(men_men_n74_), .Y(men_men_n449_));
  NO3        u433(.A(men_men_n418_), .B(x3), .C(men_men_n54_), .Y(men_men_n450_));
  NO2        u434(.A(men_men_n450_), .B(men_men_n449_), .Y(men_men_n451_));
  OAI210     u435(.A0(men_men_n156_), .A1(men_men_n448_), .B0(men_men_n451_), .Y(men_men_n452_));
  AOI220     u436(.A0(men_men_n452_), .A1(x0), .B0(men_men_n447_), .B1(men_men_n136_), .Y(men_men_n453_));
  AOI210     u437(.A0(men_men_n453_), .A1(men_men_n446_), .B0(men_men_n239_), .Y(men_men_n454_));
  NA2        u438(.A(x9), .B(x5), .Y(men_men_n455_));
  NO4        u439(.A(men_men_n107_), .B(men_men_n455_), .C(men_men_n60_), .D(men_men_n32_), .Y(men_men_n456_));
  NO4        u440(.A(men_men_n456_), .B(men_men_n454_), .C(men_men_n443_), .D(men_men_n439_), .Y(men_men_n457_));
  NA3        u441(.A(men_men_n457_), .B(men_men_n437_), .C(men_men_n398_), .Y(men_men_n458_));
  AOI210     u442(.A0(men_men_n382_), .A1(men_men_n25_), .B0(men_men_n458_), .Y(men05));
  INV        u443(.A(men_men_n184_), .Y(men_men_n462_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule