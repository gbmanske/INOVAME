// Benchmark "top" written by ABC on Thu Jun 20 14:00:11 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n142_, new_new_n143_,
    new_new_n144_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1045_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  OR4        g0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g0067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  NO2        g0068(.A(new_new_n89_), .B(new_new_n90_), .Y(new_new_n91_));
  OAI210     g0069(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n91_), .Y(new_new_n92_));
  NAi21      g0070(.An(i_6_), .B(i_10_), .Y(new_new_n93_));
  NA2        g0071(.A(i_6_), .B(i_9_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n93_), .B0(new_new_n64_), .Y(new_new_n95_));
  NA2        g0073(.A(i_2_), .B(i_6_), .Y(new_new_n96_));
  NO3        g0074(.A(new_new_n96_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n97_));
  NO2        g0075(.A(new_new_n97_), .B(new_new_n95_), .Y(new_new_n98_));
  AOI210     g0076(.A0(new_new_n98_), .A1(new_new_n92_), .B0(new_new_n81_), .Y(new_new_n99_));
  AN3        g0077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n100_));
  NAi21      g0078(.An(i_6_), .B(i_11_), .Y(new_new_n101_));
  NO2        g0079(.A(i_5_), .B(i_8_), .Y(new_new_n102_));
  NOi21      g0080(.An(new_new_n102_), .B(new_new_n101_), .Y(new_new_n103_));
  AOI220     g0081(.A0(new_new_n103_), .A1(new_new_n63_), .B0(new_new_n100_), .B1(new_new_n32_), .Y(new_new_n104_));
  INV        g0082(.A(i_7_), .Y(new_new_n105_));
  NA2        g0083(.A(new_new_n47_), .B(new_new_n105_), .Y(new_new_n106_));
  NO2        g0084(.A(i_0_), .B(i_5_), .Y(new_new_n107_));
  NO2        g0085(.A(new_new_n107_), .B(new_new_n87_), .Y(new_new_n108_));
  NA2        g0086(.A(i_12_), .B(i_3_), .Y(new_new_n109_));
  INV        g0087(.A(new_new_n109_), .Y(new_new_n110_));
  NA3        g0088(.A(new_new_n110_), .B(new_new_n108_), .C(new_new_n106_), .Y(new_new_n111_));
  NAi21      g0089(.An(i_7_), .B(i_11_), .Y(new_new_n112_));
  NO3        g0090(.A(new_new_n112_), .B(new_new_n93_), .C(new_new_n54_), .Y(new_new_n113_));
  AN2        g0091(.A(i_2_), .B(i_10_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n114_), .B(i_7_), .Y(new_new_n115_));
  OR2        g0093(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n116_));
  NO2        g0094(.A(i_8_), .B(new_new_n105_), .Y(new_new_n117_));
  NO3        g0095(.A(new_new_n117_), .B(new_new_n116_), .C(new_new_n115_), .Y(new_new_n118_));
  NA2        g0096(.A(i_12_), .B(i_7_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n120_));
  NA2        g0098(.A(i_11_), .B(i_12_), .Y(new_new_n121_));
  INV        g0099(.A(new_new_n121_), .Y(new_new_n122_));
  NO2        g0100(.A(new_new_n122_), .B(new_new_n118_), .Y(new_new_n123_));
  NAi41      g0101(.An(new_new_n113_), .B(new_new_n123_), .C(new_new_n111_), .D(new_new_n104_), .Y(new_new_n124_));
  NOi21      g0102(.An(i_1_), .B(i_5_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(i_11_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n127_));
  NA2        g0105(.A(i_7_), .B(new_new_n25_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n127_), .Y(new_new_n129_));
  NO2        g0107(.A(new_new_n129_), .B(new_new_n47_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n94_), .B(new_new_n93_), .Y(new_new_n131_));
  NAi21      g0109(.An(i_3_), .B(i_8_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(new_new_n63_), .Y(new_new_n133_));
  NOi31      g0111(.An(new_new_n133_), .B(new_new_n131_), .C(new_new_n130_), .Y(new_new_n134_));
  NO2        g0112(.A(i_1_), .B(new_new_n87_), .Y(new_new_n135_));
  NO2        g0113(.A(i_6_), .B(i_5_), .Y(new_new_n136_));
  NA2        g0114(.A(new_new_n136_), .B(i_3_), .Y(new_new_n137_));
  AO210      g0115(.A0(new_new_n137_), .A1(new_new_n48_), .B0(new_new_n135_), .Y(new_new_n138_));
  OAI220     g0116(.A0(new_new_n138_), .A1(new_new_n112_), .B0(new_new_n134_), .B1(new_new_n126_), .Y(new_new_n139_));
  NO3        g0117(.A(new_new_n139_), .B(new_new_n124_), .C(new_new_n99_), .Y(new_new_n140_));
  NA3        g0118(.A(new_new_n140_), .B(new_new_n80_), .C(new_new_n57_), .Y(mai2));
  NO2        g0119(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n142_));
  NA2        g0120(.A(i_6_), .B(new_new_n25_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(new_new_n142_), .Y(new_new_n144_));
  NA4        g0122(.A(new_new_n144_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(mai0));
  AN2        g0123(.A(i_8_), .B(i_7_), .Y(new_new_n146_));
  NA2        g0124(.A(new_new_n146_), .B(i_6_), .Y(new_new_n147_));
  NO2        g0125(.A(i_12_), .B(i_13_), .Y(new_new_n148_));
  NAi21      g0126(.An(i_5_), .B(i_11_), .Y(new_new_n149_));
  NOi21      g0127(.An(new_new_n148_), .B(new_new_n149_), .Y(new_new_n150_));
  NO2        g0128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NA2        g0129(.A(i_2_), .B(i_3_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(i_4_), .Y(new_new_n153_));
  AN2        g0131(.A(new_new_n148_), .B(new_new_n84_), .Y(new_new_n154_));
  NA2        g0132(.A(i_1_), .B(i_5_), .Y(new_new_n155_));
  NO2        g0133(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n156_));
  OR2        g0134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g0137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g0138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g0139(.A(new_new_n161_), .B(new_new_n40_), .Y(new_new_n162_));
  NO2        g0140(.A(i_3_), .B(i_5_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n164_));
  NA3        g0142(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n165_));
  NA2        g0143(.A(i_3_), .B(new_new_n49_), .Y(new_new_n166_));
  NOi21      g0144(.An(i_4_), .B(i_9_), .Y(new_new_n167_));
  NOi21      g0145(.An(i_11_), .B(i_13_), .Y(new_new_n168_));
  NA2        g0146(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n169_));
  OR2        g0147(.A(new_new_n169_), .B(new_new_n166_), .Y(new_new_n170_));
  NO2        g0148(.A(i_4_), .B(i_5_), .Y(new_new_n171_));
  NAi21      g0149(.An(i_12_), .B(i_11_), .Y(new_new_n172_));
  NO2        g0150(.A(new_new_n172_), .B(i_13_), .Y(new_new_n173_));
  NA3        g0151(.A(new_new_n173_), .B(new_new_n171_), .C(new_new_n84_), .Y(new_new_n174_));
  AOI210     g0152(.A0(new_new_n174_), .A1(new_new_n170_), .B0(new_new_n165_), .Y(new_new_n175_));
  NO2        g0153(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n176_));
  NA2        g0154(.A(new_new_n176_), .B(new_new_n47_), .Y(new_new_n177_));
  NAi31      g0155(.An(i_4_), .B(new_new_n154_), .C(i_11_), .Y(new_new_n178_));
  NA2        g0156(.A(i_3_), .B(i_5_), .Y(new_new_n179_));
  OR2        g0157(.A(new_new_n179_), .B(new_new_n169_), .Y(new_new_n180_));
  AOI210     g0158(.A0(new_new_n180_), .A1(new_new_n178_), .B0(new_new_n177_), .Y(new_new_n181_));
  NO2        g0159(.A(new_new_n74_), .B(i_5_), .Y(new_new_n182_));
  NO2        g0160(.A(i_13_), .B(i_10_), .Y(new_new_n183_));
  NA3        g0161(.A(new_new_n183_), .B(new_new_n182_), .C(new_new_n45_), .Y(new_new_n184_));
  NO2        g0162(.A(i_2_), .B(i_1_), .Y(new_new_n185_));
  NA2        g0163(.A(new_new_n185_), .B(i_3_), .Y(new_new_n186_));
  NAi21      g0164(.An(i_4_), .B(i_12_), .Y(new_new_n187_));
  NO4        g0165(.A(new_new_n187_), .B(new_new_n186_), .C(new_new_n184_), .D(new_new_n25_), .Y(new_new_n188_));
  NO3        g0166(.A(new_new_n188_), .B(new_new_n181_), .C(new_new_n175_), .Y(new_new_n189_));
  INV        g0167(.A(i_8_), .Y(new_new_n190_));
  NO2        g0168(.A(new_new_n190_), .B(i_7_), .Y(new_new_n191_));
  NA2        g0169(.A(new_new_n191_), .B(i_6_), .Y(new_new_n192_));
  NO3        g0170(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(new_new_n117_), .Y(new_new_n194_));
  NO3        g0172(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n195_));
  NO3        g0173(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n196_));
  NA2        g0174(.A(i_12_), .B(new_new_n196_), .Y(new_new_n197_));
  NO2        g0175(.A(new_new_n197_), .B(new_new_n194_), .Y(new_new_n198_));
  NO2        g0176(.A(i_3_), .B(i_8_), .Y(new_new_n199_));
  NO3        g0177(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n200_));
  NO2        g0178(.A(new_new_n107_), .B(new_new_n59_), .Y(new_new_n201_));
  NO2        g0179(.A(i_13_), .B(i_9_), .Y(new_new_n202_));
  NA3        g0180(.A(new_new_n202_), .B(i_6_), .C(new_new_n190_), .Y(new_new_n203_));
  NAi21      g0181(.An(i_12_), .B(i_3_), .Y(new_new_n204_));
  OR2        g0182(.A(new_new_n204_), .B(new_new_n203_), .Y(new_new_n205_));
  NO2        g0183(.A(new_new_n45_), .B(i_5_), .Y(new_new_n206_));
  NO3        g0184(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n207_));
  NA3        g0185(.A(new_new_n207_), .B(new_new_n206_), .C(i_10_), .Y(new_new_n208_));
  NO2        g0186(.A(new_new_n208_), .B(new_new_n205_), .Y(new_new_n209_));
  NO2        g0187(.A(new_new_n209_), .B(new_new_n198_), .Y(new_new_n210_));
  OAI220     g0188(.A0(new_new_n210_), .A1(i_4_), .B0(new_new_n192_), .B1(new_new_n189_), .Y(new_new_n211_));
  NAi21      g0189(.An(i_12_), .B(i_7_), .Y(new_new_n212_));
  NA3        g0190(.A(i_13_), .B(new_new_n190_), .C(i_10_), .Y(new_new_n213_));
  NO2        g0191(.A(new_new_n213_), .B(new_new_n212_), .Y(new_new_n214_));
  NA2        g0192(.A(i_0_), .B(i_5_), .Y(new_new_n215_));
  NA2        g0193(.A(new_new_n215_), .B(new_new_n108_), .Y(new_new_n216_));
  OAI220     g0194(.A0(new_new_n216_), .A1(new_new_n186_), .B0(new_new_n177_), .B1(new_new_n137_), .Y(new_new_n217_));
  NAi31      g0195(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n218_));
  NO2        g0196(.A(new_new_n36_), .B(i_13_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n220_));
  NO2        g0198(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n221_));
  INV        g0199(.A(i_13_), .Y(new_new_n222_));
  NO2        g0200(.A(i_12_), .B(new_new_n222_), .Y(new_new_n223_));
  NA2        g0201(.A(new_new_n217_), .B(new_new_n214_), .Y(new_new_n224_));
  NO2        g0202(.A(i_12_), .B(new_new_n37_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n179_), .B(i_4_), .Y(new_new_n226_));
  NA2        g0204(.A(new_new_n226_), .B(new_new_n225_), .Y(new_new_n227_));
  OR2        g0205(.A(i_8_), .B(i_7_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n228_), .B(new_new_n87_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n54_), .B(i_1_), .Y(new_new_n230_));
  NA2        g0208(.A(new_new_n230_), .B(new_new_n229_), .Y(new_new_n231_));
  INV        g0209(.A(i_12_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n45_), .B(new_new_n232_), .Y(new_new_n233_));
  NO3        g0211(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n234_));
  NA2        g0212(.A(i_2_), .B(i_1_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n231_), .B(new_new_n227_), .Y(new_new_n236_));
  NO3        g0214(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n237_));
  NAi21      g0215(.An(i_4_), .B(i_3_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n238_), .B(new_new_n76_), .Y(new_new_n239_));
  NO2        g0217(.A(i_0_), .B(i_6_), .Y(new_new_n240_));
  NOi41      g0218(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n241_));
  NA2        g0219(.A(new_new_n241_), .B(new_new_n240_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n235_), .B(new_new_n179_), .Y(new_new_n243_));
  NAi21      g0221(.An(new_new_n242_), .B(new_new_n243_), .Y(new_new_n244_));
  INV        g0222(.A(new_new_n244_), .Y(new_new_n245_));
  AOI220     g0223(.A0(new_new_n245_), .A1(new_new_n40_), .B0(new_new_n236_), .B1(new_new_n202_), .Y(new_new_n246_));
  NO2        g0224(.A(i_11_), .B(new_new_n222_), .Y(new_new_n247_));
  NOi21      g0225(.An(i_1_), .B(i_6_), .Y(new_new_n248_));
  NAi21      g0226(.An(i_3_), .B(i_7_), .Y(new_new_n249_));
  NA2        g0227(.A(new_new_n232_), .B(i_9_), .Y(new_new_n250_));
  OR4        g0228(.A(new_new_n250_), .B(new_new_n249_), .C(new_new_n248_), .D(new_new_n182_), .Y(new_new_n251_));
  NO2        g0229(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n252_));
  NO2        g0230(.A(i_12_), .B(i_3_), .Y(new_new_n253_));
  NA2        g0231(.A(new_new_n74_), .B(i_5_), .Y(new_new_n254_));
  NA2        g0232(.A(i_3_), .B(i_9_), .Y(new_new_n255_));
  NAi21      g0233(.An(i_7_), .B(i_10_), .Y(new_new_n256_));
  NO2        g0234(.A(new_new_n256_), .B(new_new_n255_), .Y(new_new_n257_));
  NA3        g0235(.A(new_new_n257_), .B(new_new_n254_), .C(new_new_n65_), .Y(new_new_n258_));
  NA2        g0236(.A(new_new_n258_), .B(new_new_n251_), .Y(new_new_n259_));
  NA3        g0237(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n260_));
  INV        g0238(.A(new_new_n147_), .Y(new_new_n261_));
  NA2        g0239(.A(new_new_n232_), .B(i_13_), .Y(new_new_n262_));
  NO2        g0240(.A(new_new_n262_), .B(new_new_n76_), .Y(new_new_n263_));
  AOI220     g0241(.A0(new_new_n263_), .A1(new_new_n261_), .B0(new_new_n259_), .B1(new_new_n247_), .Y(new_new_n264_));
  NO2        g0242(.A(new_new_n228_), .B(new_new_n37_), .Y(new_new_n265_));
  NA2        g0243(.A(i_12_), .B(i_6_), .Y(new_new_n266_));
  OR2        g0244(.A(i_13_), .B(i_9_), .Y(new_new_n267_));
  NO3        g0245(.A(new_new_n267_), .B(new_new_n266_), .C(new_new_n49_), .Y(new_new_n268_));
  NO2        g0246(.A(new_new_n238_), .B(i_2_), .Y(new_new_n269_));
  NA3        g0247(.A(new_new_n269_), .B(new_new_n268_), .C(new_new_n45_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n247_), .B(i_9_), .Y(new_new_n271_));
  NA2        g0249(.A(new_new_n254_), .B(new_new_n65_), .Y(new_new_n272_));
  OAI210     g0250(.A0(new_new_n272_), .A1(new_new_n271_), .B0(new_new_n270_), .Y(new_new_n273_));
  NA2        g0251(.A(new_new_n156_), .B(new_new_n64_), .Y(new_new_n274_));
  NO3        g0252(.A(i_11_), .B(new_new_n222_), .C(new_new_n25_), .Y(new_new_n275_));
  NO2        g0253(.A(new_new_n249_), .B(i_8_), .Y(new_new_n276_));
  NO2        g0254(.A(i_6_), .B(new_new_n49_), .Y(new_new_n277_));
  NA3        g0255(.A(new_new_n277_), .B(new_new_n276_), .C(new_new_n275_), .Y(new_new_n278_));
  NO3        g0256(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n279_));
  NA3        g0257(.A(new_new_n279_), .B(new_new_n265_), .C(new_new_n223_), .Y(new_new_n280_));
  AOI210     g0258(.A0(new_new_n280_), .A1(new_new_n278_), .B0(new_new_n274_), .Y(new_new_n281_));
  AOI210     g0259(.A0(new_new_n273_), .A1(new_new_n265_), .B0(new_new_n281_), .Y(new_new_n282_));
  NA4        g0260(.A(new_new_n282_), .B(new_new_n264_), .C(new_new_n246_), .D(new_new_n224_), .Y(new_new_n283_));
  NO3        g0261(.A(i_12_), .B(new_new_n222_), .C(new_new_n37_), .Y(new_new_n284_));
  INV        g0262(.A(new_new_n284_), .Y(new_new_n285_));
  NA2        g0263(.A(i_8_), .B(new_new_n105_), .Y(new_new_n286_));
  NOi21      g0264(.An(new_new_n163_), .B(new_new_n87_), .Y(new_new_n287_));
  NO3        g0265(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n288_));
  AOI220     g0266(.A0(new_new_n288_), .A1(new_new_n193_), .B0(new_new_n287_), .B1(new_new_n230_), .Y(new_new_n289_));
  NO2        g0267(.A(new_new_n289_), .B(new_new_n286_), .Y(new_new_n290_));
  NO3        g0268(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n291_));
  NO2        g0269(.A(new_new_n235_), .B(i_0_), .Y(new_new_n292_));
  AOI220     g0270(.A0(new_new_n292_), .A1(new_new_n191_), .B0(new_new_n291_), .B1(new_new_n146_), .Y(new_new_n293_));
  NA2        g0271(.A(new_new_n277_), .B(new_new_n26_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n294_), .B(new_new_n293_), .Y(new_new_n295_));
  NA2        g0273(.A(i_0_), .B(i_1_), .Y(new_new_n296_));
  NO2        g0274(.A(new_new_n296_), .B(i_2_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n60_), .B(i_6_), .Y(new_new_n298_));
  NA3        g0276(.A(new_new_n298_), .B(new_new_n297_), .C(new_new_n163_), .Y(new_new_n299_));
  INV        g0277(.A(new_new_n299_), .Y(new_new_n300_));
  NO3        g0278(.A(new_new_n300_), .B(new_new_n295_), .C(new_new_n290_), .Y(new_new_n301_));
  NO2        g0279(.A(i_3_), .B(i_10_), .Y(new_new_n302_));
  NA3        g0280(.A(new_new_n302_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n303_));
  NO2        g0281(.A(i_2_), .B(new_new_n105_), .Y(new_new_n304_));
  NA2        g0282(.A(i_1_), .B(new_new_n36_), .Y(new_new_n305_));
  NO2        g0283(.A(new_new_n305_), .B(i_8_), .Y(new_new_n306_));
  NOi21      g0284(.An(new_new_n215_), .B(new_new_n107_), .Y(new_new_n307_));
  NA3        g0285(.A(new_new_n307_), .B(new_new_n306_), .C(new_new_n304_), .Y(new_new_n308_));
  AN2        g0286(.A(i_3_), .B(i_10_), .Y(new_new_n309_));
  NO2        g0287(.A(i_5_), .B(new_new_n37_), .Y(new_new_n310_));
  NO2        g0288(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n311_));
  OR2        g0289(.A(new_new_n308_), .B(new_new_n303_), .Y(new_new_n312_));
  OAI220     g0290(.A0(new_new_n312_), .A1(i_6_), .B0(new_new_n301_), .B1(new_new_n285_), .Y(new_new_n313_));
  NO3        g0291(.A(new_new_n313_), .B(new_new_n283_), .C(new_new_n211_), .Y(new_new_n314_));
  NO3        g0292(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n315_));
  NO2        g0293(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n316_));
  NA2        g0294(.A(new_new_n292_), .B(new_new_n316_), .Y(new_new_n317_));
  NO3        g0295(.A(i_6_), .B(new_new_n190_), .C(i_7_), .Y(new_new_n318_));
  NA2        g0296(.A(new_new_n318_), .B(new_new_n195_), .Y(new_new_n319_));
  AOI210     g0297(.A0(new_new_n319_), .A1(new_new_n317_), .B0(new_new_n166_), .Y(new_new_n320_));
  NO2        g0298(.A(i_2_), .B(i_3_), .Y(new_new_n321_));
  OR2        g0299(.A(i_0_), .B(i_5_), .Y(new_new_n322_));
  NA2        g0300(.A(new_new_n215_), .B(new_new_n322_), .Y(new_new_n323_));
  NA4        g0301(.A(new_new_n323_), .B(new_new_n229_), .C(new_new_n321_), .D(i_1_), .Y(new_new_n324_));
  NA3        g0302(.A(new_new_n292_), .B(new_new_n287_), .C(new_new_n117_), .Y(new_new_n325_));
  NAi21      g0303(.An(i_8_), .B(i_7_), .Y(new_new_n326_));
  NO2        g0304(.A(new_new_n326_), .B(i_6_), .Y(new_new_n327_));
  NO2        g0305(.A(new_new_n157_), .B(new_new_n47_), .Y(new_new_n328_));
  NA2        g0306(.A(new_new_n325_), .B(new_new_n324_), .Y(new_new_n329_));
  OAI210     g0307(.A0(new_new_n329_), .A1(new_new_n320_), .B0(i_4_), .Y(new_new_n330_));
  NO2        g0308(.A(i_12_), .B(i_10_), .Y(new_new_n331_));
  NOi21      g0309(.An(i_5_), .B(i_0_), .Y(new_new_n332_));
  NO3        g0310(.A(new_new_n305_), .B(new_new_n332_), .C(new_new_n132_), .Y(new_new_n333_));
  NA4        g0311(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n334_));
  NA2        g0312(.A(new_new_n333_), .B(new_new_n331_), .Y(new_new_n335_));
  NO2        g0313(.A(i_6_), .B(i_8_), .Y(new_new_n336_));
  NOi21      g0314(.An(i_0_), .B(i_2_), .Y(new_new_n337_));
  AN2        g0315(.A(new_new_n337_), .B(new_new_n336_), .Y(new_new_n338_));
  NO2        g0316(.A(i_1_), .B(i_7_), .Y(new_new_n339_));
  AO220      g0317(.A0(new_new_n339_), .A1(new_new_n338_), .B0(new_new_n327_), .B1(new_new_n230_), .Y(new_new_n340_));
  NA3        g0318(.A(new_new_n340_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n341_));
  NA3        g0319(.A(new_new_n341_), .B(new_new_n335_), .C(new_new_n330_), .Y(new_new_n342_));
  NO3        g0320(.A(new_new_n228_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n343_));
  NO3        g0321(.A(new_new_n326_), .B(i_2_), .C(i_1_), .Y(new_new_n344_));
  OAI210     g0322(.A0(new_new_n344_), .A1(new_new_n343_), .B0(i_6_), .Y(new_new_n345_));
  NO2        g0323(.A(new_new_n345_), .B(new_new_n323_), .Y(new_new_n346_));
  NOi21      g0324(.An(new_new_n155_), .B(new_new_n108_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n347_), .B(new_new_n128_), .Y(new_new_n348_));
  OAI210     g0326(.A0(new_new_n348_), .A1(new_new_n346_), .B0(i_3_), .Y(new_new_n349_));
  INV        g0327(.A(new_new_n85_), .Y(new_new_n350_));
  NO2        g0328(.A(new_new_n296_), .B(new_new_n82_), .Y(new_new_n351_));
  NO2        g0329(.A(new_new_n96_), .B(new_new_n190_), .Y(new_new_n352_));
  NA3        g0330(.A(new_new_n307_), .B(new_new_n352_), .C(new_new_n64_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n353_), .B(new_new_n350_), .Y(new_new_n354_));
  NO2        g0332(.A(new_new_n190_), .B(i_9_), .Y(new_new_n355_));
  NA2        g0333(.A(new_new_n355_), .B(new_new_n201_), .Y(new_new_n356_));
  NO2        g0334(.A(new_new_n356_), .B(new_new_n47_), .Y(new_new_n357_));
  NO3        g0335(.A(new_new_n357_), .B(new_new_n354_), .C(new_new_n295_), .Y(new_new_n358_));
  AOI210     g0336(.A0(new_new_n358_), .A1(new_new_n349_), .B0(new_new_n162_), .Y(new_new_n359_));
  AOI210     g0337(.A0(new_new_n342_), .A1(new_new_n315_), .B0(new_new_n359_), .Y(new_new_n360_));
  NOi32      g0338(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n361_));
  INV        g0339(.A(new_new_n361_), .Y(new_new_n362_));
  NAi21      g0340(.An(i_1_), .B(i_5_), .Y(new_new_n363_));
  NAi41      g0341(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n364_));
  OAI220     g0342(.A0(new_new_n364_), .A1(new_new_n363_), .B0(new_new_n218_), .B1(new_new_n159_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n364_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n366_));
  NOi32      g0344(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n367_));
  NAi21      g0345(.An(i_6_), .B(i_1_), .Y(new_new_n368_));
  NA3        g0346(.A(new_new_n368_), .B(new_new_n367_), .C(new_new_n47_), .Y(new_new_n369_));
  NO2        g0347(.A(new_new_n369_), .B(i_0_), .Y(new_new_n370_));
  OR3        g0348(.A(new_new_n370_), .B(new_new_n366_), .C(new_new_n365_), .Y(new_new_n371_));
  NO2        g0349(.A(i_1_), .B(new_new_n105_), .Y(new_new_n372_));
  NAi21      g0350(.An(i_3_), .B(i_4_), .Y(new_new_n373_));
  NO2        g0351(.A(new_new_n373_), .B(i_9_), .Y(new_new_n374_));
  AN2        g0352(.A(i_6_), .B(i_7_), .Y(new_new_n375_));
  OAI210     g0353(.A0(new_new_n375_), .A1(new_new_n372_), .B0(new_new_n374_), .Y(new_new_n376_));
  NA2        g0354(.A(i_2_), .B(i_7_), .Y(new_new_n377_));
  NO2        g0355(.A(new_new_n373_), .B(i_10_), .Y(new_new_n378_));
  NA3        g0356(.A(new_new_n378_), .B(new_new_n377_), .C(new_new_n240_), .Y(new_new_n379_));
  AOI210     g0357(.A0(new_new_n379_), .A1(new_new_n376_), .B0(new_new_n182_), .Y(new_new_n380_));
  AOI210     g0358(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n381_));
  OAI210     g0359(.A0(new_new_n381_), .A1(new_new_n185_), .B0(new_new_n378_), .Y(new_new_n382_));
  AOI220     g0360(.A0(new_new_n378_), .A1(new_new_n339_), .B0(new_new_n234_), .B1(new_new_n185_), .Y(new_new_n383_));
  AOI210     g0361(.A0(new_new_n383_), .A1(new_new_n382_), .B0(i_5_), .Y(new_new_n384_));
  NO3        g0362(.A(new_new_n384_), .B(new_new_n380_), .C(new_new_n371_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n385_), .B(new_new_n362_), .Y(new_new_n386_));
  NO2        g0364(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n387_));
  AN2        g0365(.A(i_12_), .B(i_5_), .Y(new_new_n388_));
  NO2        g0366(.A(i_4_), .B(new_new_n26_), .Y(new_new_n389_));
  NA2        g0367(.A(new_new_n389_), .B(new_new_n388_), .Y(new_new_n390_));
  NO2        g0368(.A(i_11_), .B(i_6_), .Y(new_new_n391_));
  NA3        g0369(.A(new_new_n391_), .B(new_new_n328_), .C(new_new_n222_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n392_), .B(new_new_n390_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n238_), .B(i_5_), .Y(new_new_n394_));
  NO2        g0372(.A(i_5_), .B(i_10_), .Y(new_new_n395_));
  AOI220     g0373(.A0(new_new_n395_), .A1(new_new_n269_), .B0(new_new_n394_), .B1(new_new_n195_), .Y(new_new_n396_));
  NA2        g0374(.A(new_new_n148_), .B(new_new_n46_), .Y(new_new_n397_));
  NO2        g0375(.A(new_new_n397_), .B(new_new_n396_), .Y(new_new_n398_));
  OAI210     g0376(.A0(new_new_n398_), .A1(new_new_n393_), .B0(new_new_n387_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n400_));
  NA2        g0378(.A(new_new_n393_), .B(new_new_n400_), .Y(new_new_n401_));
  NO3        g0379(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n402_));
  NO2        g0380(.A(i_11_), .B(i_12_), .Y(new_new_n403_));
  NA2        g0381(.A(new_new_n395_), .B(new_new_n232_), .Y(new_new_n404_));
  NA3        g0382(.A(new_new_n117_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n405_));
  OAI220     g0383(.A0(new_new_n405_), .A1(new_new_n218_), .B0(new_new_n404_), .B1(new_new_n334_), .Y(new_new_n406_));
  NAi21      g0384(.An(i_13_), .B(i_0_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(new_new_n235_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n406_), .B(new_new_n408_), .Y(new_new_n409_));
  NA3        g0387(.A(new_new_n409_), .B(new_new_n401_), .C(new_new_n399_), .Y(new_new_n410_));
  NA2        g0388(.A(new_new_n45_), .B(new_new_n222_), .Y(new_new_n411_));
  NO3        g0389(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n412_));
  NO2        g0390(.A(i_0_), .B(i_11_), .Y(new_new_n413_));
  AN2        g0391(.A(i_1_), .B(i_6_), .Y(new_new_n414_));
  NOi21      g0392(.An(i_2_), .B(i_12_), .Y(new_new_n415_));
  NAi21      g0393(.An(i_9_), .B(i_4_), .Y(new_new_n416_));
  OR2        g0394(.A(i_13_), .B(i_10_), .Y(new_new_n417_));
  NO3        g0395(.A(new_new_n417_), .B(new_new_n121_), .C(new_new_n416_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n169_), .B(new_new_n127_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n105_), .B(new_new_n25_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n284_), .B(new_new_n420_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n421_), .B(new_new_n347_), .Y(new_new_n422_));
  INV        g0400(.A(new_new_n422_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n423_), .B(new_new_n26_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n325_), .B(new_new_n324_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n179_), .B(new_new_n87_), .Y(new_new_n426_));
  AOI220     g0404(.A0(new_new_n426_), .A1(new_new_n297_), .B0(new_new_n279_), .B1(new_new_n207_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n427_), .B(new_new_n286_), .Y(new_new_n428_));
  NO2        g0406(.A(new_new_n428_), .B(new_new_n425_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n190_), .B(i_10_), .Y(new_new_n430_));
  NA3        g0408(.A(new_new_n254_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n298_), .B(new_new_n230_), .Y(new_new_n432_));
  OAI220     g0410(.A0(new_new_n432_), .A1(new_new_n179_), .B0(new_new_n431_), .B1(new_new_n430_), .Y(new_new_n433_));
  NO2        g0411(.A(i_3_), .B(new_new_n49_), .Y(new_new_n434_));
  NA3        g0412(.A(new_new_n339_), .B(new_new_n338_), .C(new_new_n434_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n318_), .B(new_new_n323_), .Y(new_new_n436_));
  OAI210     g0414(.A0(new_new_n436_), .A1(new_new_n186_), .B0(new_new_n435_), .Y(new_new_n437_));
  NO2        g0415(.A(new_new_n437_), .B(new_new_n433_), .Y(new_new_n438_));
  AOI210     g0416(.A0(new_new_n438_), .A1(new_new_n429_), .B0(new_new_n271_), .Y(new_new_n439_));
  NO4        g0417(.A(new_new_n439_), .B(new_new_n424_), .C(new_new_n410_), .D(new_new_n386_), .Y(new_new_n440_));
  NO2        g0418(.A(new_new_n64_), .B(i_4_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n74_), .B(i_13_), .Y(new_new_n442_));
  NA3        g0420(.A(new_new_n442_), .B(new_new_n441_), .C(i_2_), .Y(new_new_n443_));
  NO2        g0421(.A(i_10_), .B(i_9_), .Y(new_new_n444_));
  NAi21      g0422(.An(i_12_), .B(i_8_), .Y(new_new_n445_));
  NO2        g0423(.A(new_new_n445_), .B(i_3_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n446_), .B(new_new_n444_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n47_), .B(i_4_), .Y(new_new_n448_));
  NO2        g0426(.A(new_new_n447_), .B(new_new_n443_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n311_), .B(i_0_), .Y(new_new_n450_));
  NO3        g0428(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n266_), .B(new_new_n101_), .Y(new_new_n452_));
  NA2        g0430(.A(new_new_n452_), .B(new_new_n451_), .Y(new_new_n453_));
  NA2        g0431(.A(i_8_), .B(i_9_), .Y(new_new_n454_));
  AOI210     g0432(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n455_));
  OR2        g0433(.A(new_new_n455_), .B(new_new_n454_), .Y(new_new_n456_));
  NA2        g0434(.A(new_new_n284_), .B(new_new_n201_), .Y(new_new_n457_));
  OAI220     g0435(.A0(new_new_n457_), .A1(new_new_n456_), .B0(new_new_n453_), .B1(new_new_n450_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n247_), .B(new_new_n310_), .Y(new_new_n459_));
  NO3        g0437(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n460_));
  INV        g0438(.A(new_new_n460_), .Y(new_new_n461_));
  NA3        g0439(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n462_));
  NA4        g0440(.A(new_new_n149_), .B(new_new_n120_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n463_));
  OAI220     g0441(.A0(new_new_n463_), .A1(new_new_n462_), .B0(new_new_n461_), .B1(new_new_n459_), .Y(new_new_n464_));
  NO3        g0442(.A(new_new_n464_), .B(new_new_n458_), .C(new_new_n449_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n297_), .B(new_new_n112_), .Y(new_new_n466_));
  OR2        g0444(.A(new_new_n466_), .B(new_new_n203_), .Y(new_new_n467_));
  OA210      g0445(.A0(new_new_n356_), .A1(new_new_n105_), .B0(new_new_n299_), .Y(new_new_n468_));
  OA220      g0446(.A0(new_new_n468_), .A1(new_new_n162_), .B0(new_new_n467_), .B1(new_new_n227_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n100_), .B(i_13_), .Y(new_new_n470_));
  NO2        g0448(.A(i_2_), .B(i_13_), .Y(new_new_n471_));
  NO3        g0449(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n472_));
  NO2        g0450(.A(i_6_), .B(i_7_), .Y(new_new_n473_));
  NA2        g0451(.A(new_new_n473_), .B(new_new_n472_), .Y(new_new_n474_));
  NO2        g0452(.A(i_11_), .B(i_1_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n74_), .B(i_3_), .Y(new_new_n476_));
  OR2        g0454(.A(i_11_), .B(i_8_), .Y(new_new_n477_));
  NOi21      g0455(.An(i_2_), .B(i_7_), .Y(new_new_n478_));
  NAi31      g0456(.An(new_new_n477_), .B(new_new_n478_), .C(new_new_n476_), .Y(new_new_n479_));
  NO2        g0457(.A(new_new_n417_), .B(i_6_), .Y(new_new_n480_));
  NA3        g0458(.A(new_new_n480_), .B(new_new_n441_), .C(new_new_n76_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n481_), .B(new_new_n479_), .Y(new_new_n482_));
  NO2        g0460(.A(i_6_), .B(i_10_), .Y(new_new_n483_));
  NA3        g0461(.A(new_new_n241_), .B(new_new_n168_), .C(new_new_n136_), .Y(new_new_n484_));
  NA2        g0462(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n485_));
  NO2        g0463(.A(new_new_n157_), .B(i_3_), .Y(new_new_n486_));
  NAi31      g0464(.An(new_new_n485_), .B(new_new_n486_), .C(new_new_n223_), .Y(new_new_n487_));
  NA3        g0465(.A(new_new_n400_), .B(new_new_n176_), .C(new_new_n153_), .Y(new_new_n488_));
  NA3        g0466(.A(new_new_n488_), .B(new_new_n487_), .C(new_new_n484_), .Y(new_new_n489_));
  NO2        g0467(.A(new_new_n489_), .B(new_new_n482_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n451_), .B(new_new_n388_), .Y(new_new_n491_));
  NA2        g0469(.A(new_new_n460_), .B(new_new_n395_), .Y(new_new_n492_));
  NAi21      g0470(.An(new_new_n213_), .B(new_new_n403_), .Y(new_new_n493_));
  NO2        g0471(.A(new_new_n26_), .B(i_5_), .Y(new_new_n494_));
  NO2        g0472(.A(i_0_), .B(new_new_n87_), .Y(new_new_n495_));
  NA3        g0473(.A(new_new_n495_), .B(new_new_n494_), .C(new_new_n146_), .Y(new_new_n496_));
  OR3        g0474(.A(new_new_n305_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n497_));
  NO2        g0475(.A(new_new_n497_), .B(new_new_n496_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n27_), .B(i_10_), .Y(new_new_n499_));
  NA2        g0477(.A(new_new_n315_), .B(new_new_n234_), .Y(new_new_n500_));
  OAI220     g0478(.A0(new_new_n500_), .A1(new_new_n431_), .B0(new_new_n499_), .B1(new_new_n470_), .Y(new_new_n501_));
  NA4        g0479(.A(new_new_n309_), .B(new_new_n221_), .C(new_new_n74_), .D(new_new_n232_), .Y(new_new_n502_));
  NO2        g0480(.A(new_new_n502_), .B(new_new_n474_), .Y(new_new_n503_));
  NO3        g0481(.A(new_new_n503_), .B(new_new_n501_), .C(new_new_n498_), .Y(new_new_n504_));
  NA4        g0482(.A(new_new_n504_), .B(new_new_n490_), .C(new_new_n469_), .D(new_new_n465_), .Y(new_new_n505_));
  NA3        g0483(.A(new_new_n309_), .B(new_new_n173_), .C(new_new_n171_), .Y(new_new_n506_));
  OAI210     g0484(.A0(new_new_n303_), .A1(i_4_), .B0(new_new_n506_), .Y(new_new_n507_));
  AN2        g0485(.A(new_new_n288_), .B(new_new_n229_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n508_), .B(new_new_n507_), .Y(new_new_n509_));
  NA4        g0487(.A(new_new_n442_), .B(new_new_n441_), .C(new_new_n199_), .D(i_2_), .Y(new_new_n510_));
  INV        g0488(.A(new_new_n510_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n388_), .B(new_new_n222_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n361_), .B(new_new_n74_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n375_), .B(new_new_n367_), .Y(new_new_n514_));
  OR2        g0492(.A(new_new_n512_), .B(new_new_n514_), .Y(new_new_n515_));
  NO2        g0493(.A(new_new_n36_), .B(i_8_), .Y(new_new_n516_));
  NAi41      g0494(.An(new_new_n513_), .B(new_new_n483_), .C(new_new_n516_), .D(new_new_n47_), .Y(new_new_n517_));
  AOI210     g0495(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n418_), .Y(new_new_n518_));
  NA3        g0496(.A(new_new_n518_), .B(new_new_n517_), .C(new_new_n515_), .Y(new_new_n519_));
  AOI210     g0497(.A0(new_new_n511_), .A1(new_new_n200_), .B0(new_new_n519_), .Y(new_new_n520_));
  INV        g0498(.A(new_new_n138_), .Y(new_new_n521_));
  NA2        g0499(.A(new_new_n521_), .B(new_new_n419_), .Y(new_new_n522_));
  NA3        g0500(.A(new_new_n522_), .B(new_new_n520_), .C(new_new_n509_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n394_), .B(new_new_n297_), .Y(new_new_n524_));
  OAI210     g0502(.A0(new_new_n390_), .A1(new_new_n165_), .B0(new_new_n524_), .Y(new_new_n525_));
  NO2        g0503(.A(i_12_), .B(new_new_n190_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n526_), .B(new_new_n222_), .Y(new_new_n527_));
  NA3        g0505(.A(new_new_n483_), .B(new_new_n171_), .C(new_new_n27_), .Y(new_new_n528_));
  NO2        g0506(.A(new_new_n528_), .B(new_new_n527_), .Y(new_new_n529_));
  NOi31      g0507(.An(new_new_n318_), .B(new_new_n417_), .C(new_new_n38_), .Y(new_new_n530_));
  OAI210     g0508(.A0(new_new_n530_), .A1(new_new_n529_), .B0(new_new_n525_), .Y(new_new_n531_));
  NO2        g0509(.A(i_8_), .B(i_7_), .Y(new_new_n532_));
  OAI210     g0510(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n533_));
  NA2        g0511(.A(new_new_n533_), .B(new_new_n221_), .Y(new_new_n534_));
  NO2        g0512(.A(new_new_n534_), .B(new_new_n238_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n45_), .B(i_10_), .Y(new_new_n536_));
  NO2        g0514(.A(new_new_n536_), .B(i_6_), .Y(new_new_n537_));
  NA3        g0515(.A(new_new_n537_), .B(new_new_n535_), .C(new_new_n532_), .Y(new_new_n538_));
  AOI220     g0516(.A0(new_new_n426_), .A1(new_new_n328_), .B0(new_new_n243_), .B1(new_new_n240_), .Y(new_new_n539_));
  OAI220     g0517(.A0(new_new_n539_), .A1(new_new_n262_), .B0(new_new_n470_), .B1(new_new_n137_), .Y(new_new_n540_));
  NA2        g0518(.A(new_new_n540_), .B(new_new_n265_), .Y(new_new_n541_));
  NO2        g0519(.A(new_new_n219_), .B(new_new_n45_), .Y(new_new_n542_));
  NO2        g0520(.A(new_new_n157_), .B(i_5_), .Y(new_new_n543_));
  NA3        g0521(.A(new_new_n543_), .B(new_new_n411_), .C(new_new_n321_), .Y(new_new_n544_));
  NO2        g0522(.A(new_new_n544_), .B(new_new_n542_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n545_), .B(new_new_n460_), .Y(new_new_n546_));
  NA4        g0524(.A(new_new_n546_), .B(new_new_n541_), .C(new_new_n538_), .D(new_new_n531_), .Y(new_new_n547_));
  NA3        g0525(.A(new_new_n215_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n548_));
  NA2        g0526(.A(new_new_n284_), .B(new_new_n85_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n548_), .B(new_new_n549_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n298_), .B(new_new_n288_), .Y(new_new_n551_));
  NO2        g0529(.A(new_new_n551_), .B(new_new_n170_), .Y(new_new_n552_));
  NA2        g0530(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n444_), .B(new_new_n219_), .Y(new_new_n554_));
  NO2        g0532(.A(new_new_n553_), .B(new_new_n554_), .Y(new_new_n555_));
  AOI210     g0533(.A0(new_new_n368_), .A1(new_new_n47_), .B0(new_new_n372_), .Y(new_new_n556_));
  NA2        g0534(.A(i_0_), .B(new_new_n49_), .Y(new_new_n557_));
  NA3        g0535(.A(new_new_n526_), .B(new_new_n275_), .C(new_new_n557_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n556_), .B(new_new_n558_), .Y(new_new_n559_));
  NO4        g0537(.A(new_new_n559_), .B(new_new_n555_), .C(new_new_n552_), .D(new_new_n550_), .Y(new_new_n560_));
  NO4        g0538(.A(new_new_n248_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n561_));
  NO3        g0539(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n562_));
  NO2        g0540(.A(new_new_n228_), .B(new_new_n36_), .Y(new_new_n563_));
  AN2        g0541(.A(new_new_n563_), .B(new_new_n562_), .Y(new_new_n564_));
  OA210      g0542(.A0(new_new_n564_), .A1(new_new_n561_), .B0(new_new_n361_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n417_), .B(i_1_), .Y(new_new_n566_));
  NOi31      g0544(.An(new_new_n566_), .B(new_new_n452_), .C(new_new_n74_), .Y(new_new_n567_));
  INV        g0545(.A(new_new_n565_), .Y(new_new_n568_));
  NOi21      g0546(.An(i_10_), .B(i_6_), .Y(new_new_n569_));
  NO2        g0547(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n570_));
  AOI220     g0548(.A0(new_new_n284_), .A1(new_new_n570_), .B0(new_new_n275_), .B1(new_new_n569_), .Y(new_new_n571_));
  NO2        g0549(.A(new_new_n571_), .B(new_new_n450_), .Y(new_new_n572_));
  NO2        g0550(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n573_));
  NA2        g0551(.A(new_new_n318_), .B(new_new_n164_), .Y(new_new_n574_));
  AOI220     g0552(.A0(new_new_n574_), .A1(new_new_n432_), .B0(new_new_n180_), .B1(new_new_n178_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n195_), .B(new_new_n37_), .Y(new_new_n576_));
  NOi31      g0554(.An(new_new_n150_), .B(new_new_n576_), .C(new_new_n334_), .Y(new_new_n577_));
  NO3        g0555(.A(new_new_n577_), .B(new_new_n575_), .C(new_new_n572_), .Y(new_new_n578_));
  NO2        g0556(.A(new_new_n513_), .B(new_new_n383_), .Y(new_new_n579_));
  INV        g0557(.A(new_new_n321_), .Y(new_new_n580_));
  NO2        g0558(.A(i_12_), .B(new_new_n87_), .Y(new_new_n581_));
  NA2        g0559(.A(new_new_n171_), .B(i_0_), .Y(new_new_n582_));
  NO3        g0560(.A(new_new_n582_), .B(new_new_n345_), .C(new_new_n303_), .Y(new_new_n583_));
  OR2        g0561(.A(i_2_), .B(i_5_), .Y(new_new_n584_));
  OR2        g0562(.A(new_new_n584_), .B(new_new_n414_), .Y(new_new_n585_));
  AOI210     g0563(.A0(new_new_n377_), .A1(new_new_n240_), .B0(new_new_n195_), .Y(new_new_n586_));
  AOI210     g0564(.A0(new_new_n586_), .A1(new_new_n585_), .B0(new_new_n493_), .Y(new_new_n587_));
  NO3        g0565(.A(new_new_n587_), .B(new_new_n583_), .C(new_new_n579_), .Y(new_new_n588_));
  NA4        g0566(.A(new_new_n588_), .B(new_new_n578_), .C(new_new_n568_), .D(new_new_n560_), .Y(new_new_n589_));
  NO4        g0567(.A(new_new_n589_), .B(new_new_n547_), .C(new_new_n523_), .D(new_new_n505_), .Y(new_new_n590_));
  NA4        g0568(.A(new_new_n590_), .B(new_new_n440_), .C(new_new_n360_), .D(new_new_n314_), .Y(mai7));
  NO2        g0569(.A(new_new_n96_), .B(new_new_n55_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n112_), .B(new_new_n93_), .Y(new_new_n593_));
  NA2        g0571(.A(new_new_n389_), .B(new_new_n593_), .Y(new_new_n594_));
  NA2        g0572(.A(new_new_n483_), .B(new_new_n85_), .Y(new_new_n595_));
  NA2        g0573(.A(i_11_), .B(new_new_n190_), .Y(new_new_n596_));
  NA2        g0574(.A(new_new_n148_), .B(new_new_n596_), .Y(new_new_n597_));
  OAI210     g0575(.A0(new_new_n597_), .A1(new_new_n595_), .B0(new_new_n594_), .Y(new_new_n598_));
  NA3        g0576(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n232_), .B(i_4_), .Y(new_new_n600_));
  NA2        g0578(.A(new_new_n600_), .B(i_8_), .Y(new_new_n601_));
  NO2        g0579(.A(new_new_n109_), .B(new_new_n599_), .Y(new_new_n602_));
  NA2        g0580(.A(i_2_), .B(new_new_n87_), .Y(new_new_n603_));
  OAI210     g0581(.A0(new_new_n90_), .A1(new_new_n199_), .B0(new_new_n200_), .Y(new_new_n604_));
  NO2        g0582(.A(i_7_), .B(new_new_n37_), .Y(new_new_n605_));
  NA2        g0583(.A(i_4_), .B(i_8_), .Y(new_new_n606_));
  AOI210     g0584(.A0(new_new_n606_), .A1(new_new_n309_), .B0(new_new_n605_), .Y(new_new_n607_));
  OAI220     g0585(.A0(new_new_n607_), .A1(new_new_n603_), .B0(new_new_n604_), .B1(i_13_), .Y(new_new_n608_));
  NO4        g0586(.A(new_new_n608_), .B(new_new_n602_), .C(new_new_n598_), .D(new_new_n592_), .Y(new_new_n609_));
  AOI210     g0587(.A0(new_new_n132_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n610_));
  AOI210     g0588(.A0(new_new_n610_), .A1(new_new_n232_), .B0(new_new_n161_), .Y(new_new_n611_));
  OR2        g0589(.A(i_6_), .B(i_10_), .Y(new_new_n612_));
  NO2        g0590(.A(new_new_n612_), .B(new_new_n23_), .Y(new_new_n613_));
  OR3        g0591(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n614_));
  NO3        g0592(.A(new_new_n614_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n615_));
  INV        g0593(.A(new_new_n196_), .Y(new_new_n616_));
  NO2        g0594(.A(new_new_n615_), .B(new_new_n613_), .Y(new_new_n617_));
  OA220      g0595(.A0(new_new_n617_), .A1(new_new_n580_), .B0(new_new_n611_), .B1(new_new_n267_), .Y(new_new_n618_));
  AOI210     g0596(.A0(new_new_n618_), .A1(new_new_n609_), .B0(new_new_n64_), .Y(new_new_n619_));
  NOi21      g0597(.An(i_11_), .B(i_7_), .Y(new_new_n620_));
  AO210      g0598(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n621_));
  NO2        g0599(.A(new_new_n621_), .B(new_new_n620_), .Y(new_new_n622_));
  NA2        g0600(.A(new_new_n622_), .B(new_new_n202_), .Y(new_new_n623_));
  NA3        g0601(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n624_));
  NAi31      g0602(.An(new_new_n624_), .B(new_new_n212_), .C(i_11_), .Y(new_new_n625_));
  AOI210     g0603(.A0(new_new_n625_), .A1(new_new_n623_), .B0(new_new_n64_), .Y(new_new_n626_));
  NA2        g0604(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n627_));
  AO210      g0605(.A0(new_new_n627_), .A1(new_new_n383_), .B0(new_new_n41_), .Y(new_new_n628_));
  NO3        g0606(.A(new_new_n256_), .B(new_new_n204_), .C(new_new_n596_), .Y(new_new_n629_));
  OAI210     g0607(.A0(new_new_n629_), .A1(new_new_n223_), .B0(new_new_n64_), .Y(new_new_n630_));
  NA2        g0608(.A(new_new_n415_), .B(new_new_n31_), .Y(new_new_n631_));
  OR2        g0609(.A(new_new_n204_), .B(new_new_n112_), .Y(new_new_n632_));
  NA2        g0610(.A(new_new_n632_), .B(new_new_n631_), .Y(new_new_n633_));
  NO2        g0611(.A(new_new_n64_), .B(i_9_), .Y(new_new_n634_));
  NO2        g0612(.A(new_new_n634_), .B(i_4_), .Y(new_new_n635_));
  NA2        g0613(.A(new_new_n635_), .B(new_new_n633_), .Y(new_new_n636_));
  NO2        g0614(.A(i_1_), .B(i_12_), .Y(new_new_n637_));
  NA3        g0615(.A(new_new_n637_), .B(new_new_n114_), .C(new_new_n24_), .Y(new_new_n638_));
  BUFFER     g0616(.A(new_new_n638_), .Y(new_new_n639_));
  NA4        g0617(.A(new_new_n639_), .B(new_new_n636_), .C(new_new_n630_), .D(new_new_n628_), .Y(new_new_n640_));
  OAI210     g0618(.A0(new_new_n640_), .A1(new_new_n626_), .B0(i_6_), .Y(new_new_n641_));
  NO2        g0619(.A(new_new_n624_), .B(new_new_n112_), .Y(new_new_n642_));
  NA2        g0620(.A(new_new_n642_), .B(new_new_n581_), .Y(new_new_n643_));
  NO2        g0621(.A(i_6_), .B(i_11_), .Y(new_new_n644_));
  NA2        g0622(.A(new_new_n643_), .B(new_new_n453_), .Y(new_new_n645_));
  NO3        g0623(.A(new_new_n612_), .B(new_new_n228_), .C(new_new_n23_), .Y(new_new_n646_));
  AOI210     g0624(.A0(i_1_), .A1(new_new_n257_), .B0(new_new_n646_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n647_), .B(new_new_n45_), .Y(new_new_n648_));
  INV        g0626(.A(i_2_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n142_), .B(i_9_), .Y(new_new_n650_));
  NA3        g0628(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n651_));
  NO2        g0629(.A(new_new_n47_), .B(i_1_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n650_), .B(new_new_n649_), .Y(new_new_n653_));
  NA3        g0631(.A(new_new_n634_), .B(new_new_n321_), .C(i_6_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n654_), .B(new_new_n23_), .Y(new_new_n655_));
  AOI210     g0633(.A0(new_new_n475_), .A1(new_new_n420_), .B0(new_new_n237_), .Y(new_new_n656_));
  NO2        g0634(.A(new_new_n656_), .B(new_new_n603_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n652_), .B(new_new_n266_), .Y(new_new_n658_));
  NO2        g0636(.A(i_11_), .B(new_new_n37_), .Y(new_new_n659_));
  NA2        g0637(.A(new_new_n659_), .B(new_new_n24_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n660_), .B(new_new_n658_), .Y(new_new_n661_));
  OR4        g0639(.A(new_new_n661_), .B(new_new_n657_), .C(new_new_n655_), .D(new_new_n653_), .Y(new_new_n662_));
  NO3        g0640(.A(new_new_n662_), .B(new_new_n648_), .C(new_new_n645_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n232_), .B(new_new_n105_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n664_), .B(new_new_n620_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n665_), .B(i_1_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n666_), .B(new_new_n614_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n416_), .B(new_new_n87_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n667_), .B(new_new_n47_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n228_), .B(new_new_n45_), .Y(new_new_n670_));
  NO3        g0648(.A(new_new_n670_), .B(new_new_n311_), .C(new_new_n233_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n121_), .B(new_new_n37_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n672_), .B(i_6_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n87_), .B(i_9_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n64_), .Y(new_new_n675_));
  NO2        g0653(.A(new_new_n675_), .B(new_new_n637_), .Y(new_new_n676_));
  NO4        g0654(.A(new_new_n676_), .B(new_new_n673_), .C(new_new_n671_), .D(i_4_), .Y(new_new_n677_));
  NA2        g0655(.A(i_1_), .B(i_3_), .Y(new_new_n678_));
  INV        g0656(.A(new_new_n677_), .Y(new_new_n679_));
  NA4        g0657(.A(new_new_n679_), .B(new_new_n669_), .C(new_new_n663_), .D(new_new_n641_), .Y(new_new_n680_));
  NO3        g0658(.A(new_new_n477_), .B(i_3_), .C(i_7_), .Y(new_new_n681_));
  NOi21      g0659(.An(new_new_n681_), .B(i_10_), .Y(new_new_n682_));
  OA210      g0660(.A0(new_new_n682_), .A1(new_new_n241_), .B0(new_new_n87_), .Y(new_new_n683_));
  NA2        g0661(.A(new_new_n375_), .B(new_new_n374_), .Y(new_new_n684_));
  NA3        g0662(.A(new_new_n161_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n685_));
  NA2        g0663(.A(new_new_n685_), .B(new_new_n684_), .Y(new_new_n686_));
  OAI210     g0664(.A0(new_new_n686_), .A1(new_new_n683_), .B0(i_1_), .Y(new_new_n687_));
  AOI210     g0665(.A0(new_new_n266_), .A1(new_new_n101_), .B0(i_1_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n373_), .B(i_2_), .Y(new_new_n689_));
  NA2        g0667(.A(new_new_n689_), .B(new_new_n688_), .Y(new_new_n690_));
  OAI210     g0668(.A0(new_new_n654_), .A1(new_new_n445_), .B0(new_new_n690_), .Y(new_new_n691_));
  INV        g0669(.A(new_new_n691_), .Y(new_new_n692_));
  AOI210     g0670(.A0(new_new_n692_), .A1(new_new_n687_), .B0(i_13_), .Y(new_new_n693_));
  OR2        g0671(.A(i_11_), .B(i_7_), .Y(new_new_n694_));
  NA3        g0672(.A(new_new_n694_), .B(new_new_n110_), .C(new_new_n142_), .Y(new_new_n695_));
  AOI220     g0673(.A0(new_new_n471_), .A1(new_new_n161_), .B0(new_new_n448_), .B1(new_new_n142_), .Y(new_new_n696_));
  OAI210     g0674(.A0(new_new_n696_), .A1(new_new_n45_), .B0(new_new_n695_), .Y(new_new_n697_));
  AOI210     g0675(.A0(new_new_n651_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n698_));
  NO2        g0676(.A(new_new_n478_), .B(new_new_n24_), .Y(new_new_n699_));
  AOI220     g0677(.A0(new_new_n699_), .A1(new_new_n668_), .B0(new_new_n241_), .B1(new_new_n135_), .Y(new_new_n700_));
  OAI220     g0678(.A0(new_new_n700_), .A1(new_new_n41_), .B0(new_new_n1045_), .B1(new_new_n96_), .Y(new_new_n701_));
  AOI210     g0679(.A0(new_new_n697_), .A1(new_new_n336_), .B0(new_new_n701_), .Y(new_new_n702_));
  INV        g0680(.A(new_new_n119_), .Y(new_new_n703_));
  AOI220     g0681(.A0(new_new_n703_), .A1(new_new_n73_), .B0(new_new_n391_), .B1(new_new_n652_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n704_), .B(new_new_n238_), .Y(new_new_n705_));
  AOI210     g0683(.A0(new_new_n445_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n706_));
  NOi31      g0684(.An(new_new_n706_), .B(new_new_n595_), .C(new_new_n45_), .Y(new_new_n707_));
  NA2        g0685(.A(new_new_n131_), .B(i_13_), .Y(new_new_n708_));
  NO2        g0686(.A(new_new_n651_), .B(new_new_n119_), .Y(new_new_n709_));
  INV        g0687(.A(new_new_n709_), .Y(new_new_n710_));
  OAI220     g0688(.A0(new_new_n710_), .A1(new_new_n72_), .B0(new_new_n708_), .B1(new_new_n688_), .Y(new_new_n711_));
  NO3        g0689(.A(new_new_n72_), .B(new_new_n32_), .C(new_new_n105_), .Y(new_new_n712_));
  NA2        g0690(.A(new_new_n26_), .B(new_new_n190_), .Y(new_new_n713_));
  NA2        g0691(.A(new_new_n713_), .B(i_7_), .Y(new_new_n714_));
  NO3        g0692(.A(new_new_n478_), .B(new_new_n232_), .C(new_new_n87_), .Y(new_new_n715_));
  AOI210     g0693(.A0(new_new_n715_), .A1(new_new_n714_), .B0(new_new_n712_), .Y(new_new_n716_));
  AOI220     g0694(.A0(new_new_n391_), .A1(new_new_n652_), .B0(new_new_n95_), .B1(new_new_n106_), .Y(new_new_n717_));
  OAI220     g0695(.A0(new_new_n717_), .A1(new_new_n601_), .B0(new_new_n716_), .B1(new_new_n616_), .Y(new_new_n718_));
  NO4        g0696(.A(new_new_n718_), .B(new_new_n711_), .C(new_new_n707_), .D(new_new_n705_), .Y(new_new_n719_));
  OR2        g0697(.A(i_11_), .B(i_6_), .Y(new_new_n720_));
  NA3        g0698(.A(new_new_n600_), .B(new_new_n713_), .C(i_7_), .Y(new_new_n721_));
  AOI210     g0699(.A0(new_new_n721_), .A1(new_new_n710_), .B0(new_new_n720_), .Y(new_new_n722_));
  NA3        g0700(.A(new_new_n415_), .B(new_new_n605_), .C(new_new_n101_), .Y(new_new_n723_));
  NA2        g0701(.A(new_new_n644_), .B(i_13_), .Y(new_new_n724_));
  NA2        g0702(.A(new_new_n106_), .B(new_new_n713_), .Y(new_new_n725_));
  NAi21      g0703(.An(i_11_), .B(i_12_), .Y(new_new_n726_));
  NOi41      g0704(.An(new_new_n115_), .B(new_new_n726_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n727_));
  NO3        g0705(.A(new_new_n478_), .B(new_new_n581_), .C(new_new_n606_), .Y(new_new_n728_));
  AOI220     g0706(.A0(new_new_n728_), .A1(new_new_n315_), .B0(new_new_n727_), .B1(new_new_n725_), .Y(new_new_n729_));
  NA3        g0707(.A(new_new_n729_), .B(new_new_n724_), .C(new_new_n723_), .Y(new_new_n730_));
  OAI210     g0708(.A0(new_new_n730_), .A1(new_new_n722_), .B0(new_new_n64_), .Y(new_new_n731_));
  NO2        g0709(.A(i_2_), .B(i_12_), .Y(new_new_n732_));
  NA2        g0710(.A(new_new_n372_), .B(new_new_n732_), .Y(new_new_n733_));
  NA2        g0711(.A(new_new_n374_), .B(new_new_n372_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n132_), .B(i_2_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n735_), .B(new_new_n637_), .Y(new_new_n736_));
  NA3        g0714(.A(new_new_n736_), .B(new_new_n734_), .C(new_new_n733_), .Y(new_new_n737_));
  NA3        g0715(.A(new_new_n737_), .B(new_new_n46_), .C(new_new_n222_), .Y(new_new_n738_));
  NA4        g0716(.A(new_new_n738_), .B(new_new_n731_), .C(new_new_n719_), .D(new_new_n702_), .Y(new_new_n739_));
  OR4        g0717(.A(new_new_n739_), .B(new_new_n693_), .C(new_new_n680_), .D(new_new_n619_), .Y(mai5));
  NA2        g0718(.A(new_new_n665_), .B(new_new_n269_), .Y(new_new_n741_));
  AN2        g0719(.A(new_new_n24_), .B(i_10_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n742_), .B(new_new_n732_), .C(new_new_n112_), .Y(new_new_n743_));
  NO2        g0721(.A(new_new_n601_), .B(i_11_), .Y(new_new_n744_));
  NA2        g0722(.A(new_new_n90_), .B(new_new_n744_), .Y(new_new_n745_));
  NA3        g0723(.A(new_new_n745_), .B(new_new_n743_), .C(new_new_n741_), .Y(new_new_n746_));
  NO3        g0724(.A(i_11_), .B(new_new_n232_), .C(i_13_), .Y(new_new_n747_));
  NO2        g0725(.A(new_new_n128_), .B(new_new_n23_), .Y(new_new_n748_));
  NA2        g0726(.A(i_12_), .B(i_8_), .Y(new_new_n749_));
  OAI210     g0727(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n749_), .Y(new_new_n750_));
  INV        g0728(.A(new_new_n444_), .Y(new_new_n751_));
  AOI220     g0729(.A0(new_new_n321_), .A1(new_new_n573_), .B0(new_new_n750_), .B1(new_new_n748_), .Y(new_new_n752_));
  INV        g0730(.A(new_new_n752_), .Y(new_new_n753_));
  NO2        g0731(.A(new_new_n753_), .B(new_new_n746_), .Y(new_new_n754_));
  INV        g0732(.A(new_new_n168_), .Y(new_new_n755_));
  INV        g0733(.A(new_new_n241_), .Y(new_new_n756_));
  OAI210     g0734(.A0(new_new_n689_), .A1(new_new_n446_), .B0(new_new_n115_), .Y(new_new_n757_));
  AOI210     g0735(.A0(new_new_n757_), .A1(new_new_n756_), .B0(new_new_n755_), .Y(new_new_n758_));
  NO2        g0736(.A(new_new_n454_), .B(new_new_n26_), .Y(new_new_n759_));
  NO2        g0737(.A(new_new_n759_), .B(new_new_n420_), .Y(new_new_n760_));
  NA2        g0738(.A(new_new_n760_), .B(i_2_), .Y(new_new_n761_));
  INV        g0739(.A(new_new_n761_), .Y(new_new_n762_));
  AOI210     g0740(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n417_), .Y(new_new_n763_));
  AOI210     g0741(.A0(new_new_n763_), .A1(new_new_n762_), .B0(new_new_n758_), .Y(new_new_n764_));
  NO2        g0742(.A(new_new_n187_), .B(new_new_n129_), .Y(new_new_n765_));
  OAI210     g0743(.A0(new_new_n765_), .A1(new_new_n748_), .B0(i_2_), .Y(new_new_n766_));
  INV        g0744(.A(new_new_n169_), .Y(new_new_n767_));
  NO3        g0745(.A(new_new_n621_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n768_));
  AOI210     g0746(.A0(new_new_n767_), .A1(new_new_n90_), .B0(new_new_n768_), .Y(new_new_n769_));
  AOI210     g0747(.A0(new_new_n769_), .A1(new_new_n766_), .B0(new_new_n190_), .Y(new_new_n770_));
  OA210      g0748(.A0(new_new_n622_), .A1(new_new_n130_), .B0(i_13_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n196_), .B(new_new_n199_), .Y(new_new_n772_));
  NA2        g0750(.A(new_new_n154_), .B(new_new_n596_), .Y(new_new_n773_));
  AOI210     g0751(.A0(new_new_n773_), .A1(new_new_n772_), .B0(new_new_n377_), .Y(new_new_n774_));
  AOI210     g0752(.A0(new_new_n204_), .A1(new_new_n152_), .B0(new_new_n516_), .Y(new_new_n775_));
  NA2        g0753(.A(new_new_n775_), .B(new_new_n420_), .Y(new_new_n776_));
  NO2        g0754(.A(new_new_n106_), .B(new_new_n45_), .Y(new_new_n777_));
  INV        g0755(.A(new_new_n304_), .Y(new_new_n778_));
  NA4        g0756(.A(new_new_n778_), .B(new_new_n309_), .C(new_new_n128_), .D(new_new_n43_), .Y(new_new_n779_));
  OAI210     g0757(.A0(new_new_n779_), .A1(new_new_n777_), .B0(new_new_n776_), .Y(new_new_n780_));
  NO4        g0758(.A(new_new_n780_), .B(new_new_n774_), .C(new_new_n771_), .D(new_new_n770_), .Y(new_new_n781_));
  NA2        g0759(.A(new_new_n573_), .B(new_new_n28_), .Y(new_new_n782_));
  NA2        g0760(.A(new_new_n747_), .B(new_new_n276_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(new_new_n782_), .Y(new_new_n784_));
  NO2        g0762(.A(new_new_n63_), .B(i_12_), .Y(new_new_n785_));
  NO2        g0763(.A(new_new_n785_), .B(new_new_n130_), .Y(new_new_n786_));
  NO2        g0764(.A(new_new_n786_), .B(new_new_n596_), .Y(new_new_n787_));
  AOI220     g0765(.A0(new_new_n787_), .A1(new_new_n36_), .B0(new_new_n784_), .B1(new_new_n47_), .Y(new_new_n788_));
  NA4        g0766(.A(new_new_n788_), .B(new_new_n781_), .C(new_new_n764_), .D(new_new_n754_), .Y(mai6));
  NO3        g0767(.A(new_new_n252_), .B(new_new_n310_), .C(i_1_), .Y(new_new_n790_));
  NO2        g0768(.A(new_new_n182_), .B(new_new_n143_), .Y(new_new_n791_));
  OAI210     g0769(.A0(new_new_n791_), .A1(new_new_n790_), .B0(new_new_n735_), .Y(new_new_n792_));
  NO2        g0770(.A(new_new_n218_), .B(new_new_n485_), .Y(new_new_n793_));
  NO2        g0771(.A(i_11_), .B(i_9_), .Y(new_new_n794_));
  INV        g0772(.A(new_new_n332_), .Y(new_new_n795_));
  AO210      g0773(.A0(new_new_n795_), .A1(new_new_n792_), .B0(i_12_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n378_), .B(new_new_n339_), .Y(new_new_n797_));
  NA2        g0775(.A(new_new_n581_), .B(new_new_n64_), .Y(new_new_n798_));
  NA2        g0776(.A(new_new_n682_), .B(new_new_n72_), .Y(new_new_n799_));
  BUFFER     g0777(.A(new_new_n627_), .Y(new_new_n800_));
  NA4        g0778(.A(new_new_n800_), .B(new_new_n799_), .C(new_new_n798_), .D(new_new_n797_), .Y(new_new_n801_));
  INV        g0779(.A(new_new_n194_), .Y(new_new_n802_));
  AOI220     g0780(.A0(new_new_n802_), .A1(new_new_n794_), .B0(new_new_n801_), .B1(new_new_n74_), .Y(new_new_n803_));
  INV        g0781(.A(new_new_n331_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n76_), .B(new_new_n135_), .Y(new_new_n805_));
  INV        g0783(.A(new_new_n128_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n806_), .B(new_new_n47_), .Y(new_new_n807_));
  AOI210     g0785(.A0(new_new_n807_), .A1(new_new_n805_), .B0(new_new_n804_), .Y(new_new_n808_));
  NO3        g0786(.A(new_new_n248_), .B(new_new_n136_), .C(i_9_), .Y(new_new_n809_));
  NA2        g0787(.A(new_new_n809_), .B(new_new_n785_), .Y(new_new_n810_));
  AOI210     g0788(.A0(new_new_n810_), .A1(new_new_n514_), .B0(new_new_n182_), .Y(new_new_n811_));
  NO2        g0789(.A(new_new_n32_), .B(i_11_), .Y(new_new_n812_));
  NA3        g0790(.A(new_new_n812_), .B(new_new_n473_), .C(new_new_n395_), .Y(new_new_n813_));
  NAi32      g0791(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n814_));
  NO2        g0792(.A(new_new_n720_), .B(new_new_n814_), .Y(new_new_n815_));
  OAI210     g0793(.A0(new_new_n681_), .A1(new_new_n563_), .B0(new_new_n562_), .Y(new_new_n816_));
  NAi31      g0794(.An(new_new_n815_), .B(new_new_n816_), .C(new_new_n813_), .Y(new_new_n817_));
  OR3        g0795(.A(new_new_n817_), .B(new_new_n811_), .C(new_new_n808_), .Y(new_new_n818_));
  NO2        g0796(.A(new_new_n694_), .B(i_2_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n820_));
  NO2        g0798(.A(new_new_n820_), .B(new_new_n414_), .Y(new_new_n821_));
  NA2        g0799(.A(new_new_n821_), .B(new_new_n819_), .Y(new_new_n822_));
  OR2        g0800(.A(new_new_n622_), .B(new_new_n446_), .Y(new_new_n823_));
  NA3        g0801(.A(new_new_n823_), .B(new_new_n151_), .C(new_new_n70_), .Y(new_new_n824_));
  AO210      g0802(.A0(new_new_n492_), .A1(new_new_n751_), .B0(new_new_n36_), .Y(new_new_n825_));
  NA3        g0803(.A(new_new_n825_), .B(new_new_n824_), .C(new_new_n822_), .Y(new_new_n826_));
  OAI210     g0804(.A0(i_6_), .A1(i_11_), .B0(new_new_n88_), .Y(new_new_n827_));
  AOI220     g0805(.A0(new_new_n827_), .A1(new_new_n562_), .B0(new_new_n793_), .B1(new_new_n714_), .Y(new_new_n828_));
  NA3        g0806(.A(new_new_n377_), .B(new_new_n234_), .C(new_new_n151_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n402_), .B(new_new_n71_), .Y(new_new_n830_));
  NA4        g0808(.A(new_new_n830_), .B(new_new_n829_), .C(new_new_n828_), .D(new_new_n604_), .Y(new_new_n831_));
  AO210      g0809(.A0(new_new_n516_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n832_));
  NA3        g0810(.A(new_new_n832_), .B(new_new_n483_), .C(new_new_n215_), .Y(new_new_n833_));
  AOI210     g0811(.A0(new_new_n446_), .A1(new_new_n444_), .B0(new_new_n561_), .Y(new_new_n834_));
  NO2        g0812(.A(new_new_n612_), .B(new_new_n106_), .Y(new_new_n835_));
  OAI210     g0813(.A0(new_new_n835_), .A1(new_new_n116_), .B0(new_new_n413_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n240_), .B(new_new_n47_), .Y(new_new_n837_));
  INV        g0815(.A(new_new_n585_), .Y(new_new_n838_));
  NA3        g0816(.A(new_new_n838_), .B(new_new_n331_), .C(i_7_), .Y(new_new_n839_));
  NA4        g0817(.A(new_new_n839_), .B(new_new_n836_), .C(new_new_n834_), .D(new_new_n833_), .Y(new_new_n840_));
  NO4        g0818(.A(new_new_n840_), .B(new_new_n831_), .C(new_new_n826_), .D(new_new_n818_), .Y(new_new_n841_));
  NA4        g0819(.A(new_new_n841_), .B(new_new_n803_), .C(new_new_n796_), .D(new_new_n385_), .Y(mai3));
  NA2        g0820(.A(i_12_), .B(i_10_), .Y(new_new_n843_));
  NA2        g0821(.A(i_6_), .B(i_7_), .Y(new_new_n844_));
  NO2        g0822(.A(new_new_n844_), .B(i_0_), .Y(new_new_n845_));
  NO2        g0823(.A(i_11_), .B(new_new_n232_), .Y(new_new_n846_));
  OAI210     g0824(.A0(new_new_n845_), .A1(new_new_n292_), .B0(new_new_n846_), .Y(new_new_n847_));
  NO2        g0825(.A(new_new_n847_), .B(new_new_n190_), .Y(new_new_n848_));
  NO3        g0826(.A(new_new_n450_), .B(new_new_n93_), .C(new_new_n45_), .Y(new_new_n849_));
  OA210      g0827(.A0(new_new_n849_), .A1(new_new_n848_), .B0(new_new_n171_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n829_), .B(new_new_n376_), .Y(new_new_n851_));
  NA2        g0829(.A(new_new_n851_), .B(new_new_n40_), .Y(new_new_n852_));
  NOi21      g0830(.An(new_new_n100_), .B(new_new_n760_), .Y(new_new_n853_));
  NO3        g0831(.A(new_new_n632_), .B(new_new_n454_), .C(new_new_n135_), .Y(new_new_n854_));
  NA2        g0832(.A(new_new_n415_), .B(new_new_n46_), .Y(new_new_n855_));
  AN2        g0833(.A(new_new_n452_), .B(new_new_n56_), .Y(new_new_n856_));
  NO3        g0834(.A(new_new_n856_), .B(new_new_n854_), .C(new_new_n853_), .Y(new_new_n857_));
  AOI210     g0835(.A0(new_new_n857_), .A1(new_new_n852_), .B0(new_new_n49_), .Y(new_new_n858_));
  NO4        g0836(.A(new_new_n381_), .B(new_new_n388_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n182_), .B(new_new_n569_), .Y(new_new_n860_));
  NOi21      g0838(.An(new_new_n860_), .B(new_new_n859_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n706_), .B(new_new_n674_), .Y(new_new_n862_));
  NA2        g0840(.A(new_new_n337_), .B(new_new_n434_), .Y(new_new_n863_));
  OAI220     g0841(.A0(new_new_n863_), .A1(new_new_n862_), .B0(new_new_n861_), .B1(new_new_n64_), .Y(new_new_n864_));
  NOi21      g0842(.An(i_5_), .B(i_9_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n865_), .B(new_new_n442_), .Y(new_new_n866_));
  BUFFER     g0844(.A(new_new_n266_), .Y(new_new_n867_));
  NA2        g0845(.A(new_new_n867_), .B(new_new_n475_), .Y(new_new_n868_));
  NO2        g0846(.A(new_new_n172_), .B(new_new_n152_), .Y(new_new_n869_));
  NO2        g0847(.A(new_new_n868_), .B(new_new_n866_), .Y(new_new_n870_));
  NO4        g0848(.A(new_new_n870_), .B(new_new_n864_), .C(new_new_n858_), .D(new_new_n850_), .Y(new_new_n871_));
  NA2        g0849(.A(new_new_n182_), .B(new_new_n24_), .Y(new_new_n872_));
  NO2        g0850(.A(new_new_n672_), .B(new_new_n593_), .Y(new_new_n873_));
  NO2        g0851(.A(new_new_n873_), .B(new_new_n872_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n315_), .B(new_new_n133_), .Y(new_new_n875_));
  NAi21      g0853(.An(new_new_n162_), .B(new_new_n434_), .Y(new_new_n876_));
  OAI220     g0854(.A0(new_new_n876_), .A1(new_new_n837_), .B0(new_new_n875_), .B1(new_new_n404_), .Y(new_new_n877_));
  NO2        g0855(.A(new_new_n877_), .B(new_new_n874_), .Y(new_new_n878_));
  NO2        g0856(.A(new_new_n395_), .B(new_new_n296_), .Y(new_new_n879_));
  NA2        g0857(.A(new_new_n879_), .B(new_new_n709_), .Y(new_new_n880_));
  NA2        g0858(.A(new_new_n570_), .B(i_0_), .Y(new_new_n881_));
  NO3        g0859(.A(new_new_n881_), .B(new_new_n390_), .C(new_new_n90_), .Y(new_new_n882_));
  NO4        g0860(.A(new_new_n584_), .B(new_new_n212_), .C(new_new_n417_), .D(new_new_n414_), .Y(new_new_n883_));
  AOI210     g0861(.A0(new_new_n883_), .A1(i_11_), .B0(new_new_n882_), .Y(new_new_n884_));
  INV        g0862(.A(new_new_n473_), .Y(new_new_n885_));
  AN2        g0863(.A(new_new_n100_), .B(new_new_n239_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n747_), .B(new_new_n332_), .Y(new_new_n887_));
  AOI210     g0865(.A0(new_new_n483_), .A1(new_new_n90_), .B0(new_new_n59_), .Y(new_new_n888_));
  OAI220     g0866(.A0(new_new_n888_), .A1(new_new_n887_), .B0(new_new_n660_), .B1(new_new_n534_), .Y(new_new_n889_));
  NO2        g0867(.A(new_new_n250_), .B(new_new_n155_), .Y(new_new_n890_));
  NA2        g0868(.A(i_0_), .B(i_10_), .Y(new_new_n891_));
  AN2        g0869(.A(new_new_n890_), .B(i_6_), .Y(new_new_n892_));
  NO3        g0870(.A(new_new_n892_), .B(new_new_n889_), .C(new_new_n886_), .Y(new_new_n893_));
  NA4        g0871(.A(new_new_n893_), .B(new_new_n884_), .C(new_new_n880_), .D(new_new_n878_), .Y(new_new_n894_));
  NO2        g0872(.A(new_new_n107_), .B(new_new_n37_), .Y(new_new_n895_));
  NA2        g0873(.A(i_11_), .B(i_9_), .Y(new_new_n896_));
  NO3        g0874(.A(i_12_), .B(new_new_n896_), .C(new_new_n603_), .Y(new_new_n897_));
  AN2        g0875(.A(new_new_n897_), .B(new_new_n895_), .Y(new_new_n898_));
  NO2        g0876(.A(new_new_n49_), .B(i_7_), .Y(new_new_n899_));
  NA2        g0877(.A(new_new_n400_), .B(new_new_n176_), .Y(new_new_n900_));
  NA2        g0878(.A(new_new_n900_), .B(new_new_n160_), .Y(new_new_n901_));
  NO2        g0879(.A(new_new_n896_), .B(new_new_n74_), .Y(new_new_n902_));
  AOI210     g0880(.A0(new_new_n375_), .A1(new_new_n42_), .B0(new_new_n412_), .Y(new_new_n903_));
  NO2        g0881(.A(new_new_n903_), .B(new_new_n866_), .Y(new_new_n904_));
  NO3        g0882(.A(new_new_n904_), .B(new_new_n901_), .C(new_new_n898_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n659_), .B(new_new_n125_), .Y(new_new_n906_));
  NO2        g0884(.A(i_6_), .B(new_new_n906_), .Y(new_new_n907_));
  AOI210     g0885(.A0(new_new_n445_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n908_));
  NA2        g0886(.A(new_new_n168_), .B(new_new_n107_), .Y(new_new_n909_));
  NOi32      g0887(.An(new_new_n908_), .Bn(new_new_n185_), .C(new_new_n909_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n605_), .B(new_new_n332_), .Y(new_new_n911_));
  NO2        g0889(.A(new_new_n911_), .B(new_new_n855_), .Y(new_new_n912_));
  NO3        g0890(.A(new_new_n912_), .B(new_new_n910_), .C(new_new_n907_), .Y(new_new_n913_));
  NOi21      g0891(.An(i_7_), .B(i_5_), .Y(new_new_n914_));
  NOi31      g0892(.An(new_new_n914_), .B(i_0_), .C(new_new_n726_), .Y(new_new_n915_));
  NA3        g0893(.A(new_new_n915_), .B(new_new_n389_), .C(i_6_), .Y(new_new_n916_));
  OA210      g0894(.A0(new_new_n909_), .A1(new_new_n514_), .B0(new_new_n916_), .Y(new_new_n917_));
  NO3        g0895(.A(new_new_n407_), .B(new_new_n364_), .C(new_new_n363_), .Y(new_new_n918_));
  NO2        g0896(.A(new_new_n260_), .B(new_new_n322_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n726_), .B(new_new_n255_), .Y(new_new_n920_));
  AOI210     g0898(.A0(new_new_n920_), .A1(new_new_n919_), .B0(new_new_n918_), .Y(new_new_n921_));
  NA4        g0899(.A(new_new_n921_), .B(new_new_n917_), .C(new_new_n913_), .D(new_new_n905_), .Y(new_new_n922_));
  NO2        g0900(.A(new_new_n872_), .B(new_new_n235_), .Y(new_new_n923_));
  AN2        g0901(.A(new_new_n336_), .B(new_new_n332_), .Y(new_new_n924_));
  AN2        g0902(.A(new_new_n924_), .B(new_new_n869_), .Y(new_new_n925_));
  OAI210     g0903(.A0(new_new_n925_), .A1(new_new_n923_), .B0(i_10_), .Y(new_new_n926_));
  NO2        g0904(.A(new_new_n843_), .B(new_new_n321_), .Y(new_new_n927_));
  OA210      g0905(.A0(new_new_n473_), .A1(new_new_n221_), .B0(new_new_n472_), .Y(new_new_n928_));
  NA2        g0906(.A(new_new_n927_), .B(new_new_n902_), .Y(new_new_n929_));
  NA3        g0907(.A(new_new_n472_), .B(new_new_n415_), .C(new_new_n46_), .Y(new_new_n930_));
  OAI210     g0908(.A0(new_new_n876_), .A1(new_new_n885_), .B0(new_new_n930_), .Y(new_new_n931_));
  NO2        g0909(.A(new_new_n253_), .B(new_new_n47_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n902_), .B(new_new_n309_), .Y(new_new_n933_));
  OAI210     g0911(.A0(new_new_n932_), .A1(new_new_n184_), .B0(new_new_n933_), .Y(new_new_n934_));
  AOI220     g0912(.A0(new_new_n934_), .A1(new_new_n473_), .B0(new_new_n931_), .B1(new_new_n74_), .Y(new_new_n935_));
  NA2        g0913(.A(new_new_n96_), .B(new_new_n45_), .Y(new_new_n936_));
  NO2        g0914(.A(new_new_n76_), .B(new_new_n749_), .Y(new_new_n937_));
  AOI220     g0915(.A0(new_new_n937_), .A1(new_new_n936_), .B0(new_new_n171_), .B1(new_new_n593_), .Y(new_new_n938_));
  NO2        g0916(.A(new_new_n938_), .B(new_new_n48_), .Y(new_new_n939_));
  NA2        g0917(.A(new_new_n699_), .B(new_new_n543_), .Y(new_new_n940_));
  NAi21      g0918(.An(i_9_), .B(i_5_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n941_), .B(new_new_n407_), .Y(new_new_n942_));
  NO2        g0920(.A(new_new_n599_), .B(new_new_n109_), .Y(new_new_n943_));
  AOI220     g0921(.A0(new_new_n943_), .A1(i_0_), .B0(new_new_n942_), .B1(new_new_n622_), .Y(new_new_n944_));
  OAI220     g0922(.A0(new_new_n944_), .A1(new_new_n87_), .B0(new_new_n940_), .B1(new_new_n169_), .Y(new_new_n945_));
  NO3        g0923(.A(new_new_n945_), .B(new_new_n939_), .C(new_new_n519_), .Y(new_new_n946_));
  NA4        g0924(.A(new_new_n946_), .B(new_new_n935_), .C(new_new_n929_), .D(new_new_n926_), .Y(new_new_n947_));
  NO3        g0925(.A(new_new_n947_), .B(new_new_n922_), .C(new_new_n894_), .Y(new_new_n948_));
  NO2        g0926(.A(i_0_), .B(new_new_n726_), .Y(new_new_n949_));
  NA2        g0927(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n950_));
  INV        g0928(.A(new_new_n950_), .Y(new_new_n951_));
  NO3        g0929(.A(new_new_n109_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n952_));
  AO220      g0930(.A0(new_new_n952_), .A1(new_new_n951_), .B0(new_new_n949_), .B1(new_new_n171_), .Y(new_new_n953_));
  AOI210     g0931(.A0(new_new_n798_), .A1(new_new_n684_), .B0(new_new_n909_), .Y(new_new_n954_));
  AOI210     g0932(.A0(new_new_n953_), .A1(new_new_n352_), .B0(new_new_n954_), .Y(new_new_n955_));
  NA2        g0933(.A(new_new_n735_), .B(new_new_n150_), .Y(new_new_n956_));
  INV        g0934(.A(new_new_n956_), .Y(new_new_n957_));
  NA3        g0935(.A(new_new_n957_), .B(new_new_n674_), .C(new_new_n74_), .Y(new_new_n958_));
  NO2        g0936(.A(new_new_n816_), .B(new_new_n407_), .Y(new_new_n959_));
  NA3        g0937(.A(new_new_n845_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n960_));
  NA2        g0938(.A(new_new_n846_), .B(i_9_), .Y(new_new_n961_));
  AOI210     g0939(.A0(new_new_n960_), .A1(new_new_n496_), .B0(new_new_n961_), .Y(new_new_n962_));
  OAI210     g0940(.A0(new_new_n240_), .A1(i_9_), .B0(new_new_n225_), .Y(new_new_n963_));
  AOI210     g0941(.A0(new_new_n963_), .A1(new_new_n881_), .B0(new_new_n155_), .Y(new_new_n964_));
  NO3        g0942(.A(new_new_n964_), .B(new_new_n962_), .C(new_new_n959_), .Y(new_new_n965_));
  NA3        g0943(.A(new_new_n965_), .B(new_new_n958_), .C(new_new_n955_), .Y(new_new_n966_));
  NA3        g0944(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n967_));
  NA2        g0945(.A(new_new_n899_), .B(new_new_n486_), .Y(new_new_n968_));
  AOI210     g0946(.A0(new_new_n967_), .A1(new_new_n162_), .B0(new_new_n968_), .Y(new_new_n969_));
  INV        g0947(.A(new_new_n969_), .Y(new_new_n970_));
  NO3        g0948(.A(new_new_n891_), .B(new_new_n865_), .C(new_new_n187_), .Y(new_new_n971_));
  AOI220     g0949(.A0(new_new_n971_), .A1(i_11_), .B0(new_new_n567_), .B1(new_new_n76_), .Y(new_new_n972_));
  NO3        g0950(.A(new_new_n206_), .B(new_new_n388_), .C(i_0_), .Y(new_new_n973_));
  OAI210     g0951(.A0(new_new_n973_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n974_));
  NA3        g0952(.A(new_new_n974_), .B(new_new_n972_), .C(new_new_n970_), .Y(new_new_n975_));
  NO2        g0953(.A(new_new_n238_), .B(new_new_n96_), .Y(new_new_n976_));
  AOI210     g0954(.A0(new_new_n976_), .A1(new_new_n949_), .B0(new_new_n113_), .Y(new_new_n977_));
  OR2        g0955(.A(new_new_n977_), .B(i_5_), .Y(new_new_n978_));
  AOI210     g0956(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n172_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n979_), .B(new_new_n928_), .Y(new_new_n980_));
  NO3        g0958(.A(new_new_n855_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n491_), .B(new_new_n484_), .Y(new_new_n982_));
  NO2        g0960(.A(new_new_n982_), .B(new_new_n981_), .Y(new_new_n983_));
  NA3        g0961(.A(new_new_n395_), .B(new_new_n168_), .C(new_new_n167_), .Y(new_new_n984_));
  NA3        g0962(.A(new_new_n899_), .B(new_new_n292_), .C(new_new_n225_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n985_), .B(new_new_n984_), .Y(new_new_n986_));
  NOi31      g0964(.An(new_new_n394_), .B(new_new_n950_), .C(new_new_n235_), .Y(new_new_n987_));
  NO3        g0965(.A(new_new_n896_), .B(new_new_n215_), .C(new_new_n187_), .Y(new_new_n988_));
  NO3        g0966(.A(new_new_n988_), .B(new_new_n987_), .C(new_new_n986_), .Y(new_new_n989_));
  NA4        g0967(.A(new_new_n989_), .B(new_new_n983_), .C(new_new_n980_), .D(new_new_n978_), .Y(new_new_n990_));
  INV        g0968(.A(new_new_n615_), .Y(new_new_n991_));
  NO3        g0969(.A(new_new_n991_), .B(new_new_n557_), .C(new_new_n350_), .Y(new_new_n992_));
  NO2        g0970(.A(new_new_n87_), .B(i_5_), .Y(new_new_n993_));
  NA3        g0971(.A(new_new_n846_), .B(new_new_n114_), .C(new_new_n128_), .Y(new_new_n994_));
  INV        g0972(.A(new_new_n994_), .Y(new_new_n995_));
  AOI210     g0973(.A0(new_new_n995_), .A1(new_new_n993_), .B0(new_new_n992_), .Y(new_new_n996_));
  NAi21      g0974(.An(new_new_n237_), .B(new_new_n238_), .Y(new_new_n997_));
  NO4        g0975(.A(new_new_n235_), .B(new_new_n206_), .C(i_0_), .D(i_12_), .Y(new_new_n998_));
  NA2        g0976(.A(new_new_n998_), .B(new_new_n997_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n999_), .B(new_new_n996_), .Y(new_new_n1000_));
  NO4        g0978(.A(new_new_n1000_), .B(new_new_n990_), .C(new_new_n975_), .D(new_new_n966_), .Y(new_new_n1001_));
  OAI210     g0979(.A0(new_new_n819_), .A1(new_new_n812_), .B0(new_new_n37_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n908_), .B(new_new_n372_), .C(i_5_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n1003_), .B(new_new_n1002_), .C(new_new_n611_), .Y(new_new_n1004_));
  NA2        g0982(.A(new_new_n1004_), .B(new_new_n202_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n183_), .B(new_new_n185_), .Y(new_new_n1006_));
  AO210      g0984(.A0(new_new_n694_), .A1(new_new_n33_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  OAI210     g0985(.A0(new_new_n615_), .A1(new_new_n613_), .B0(new_new_n321_), .Y(new_new_n1008_));
  NAi31      g0986(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1009_));
  NO2        g0987(.A(new_new_n71_), .B(new_new_n1009_), .Y(new_new_n1010_));
  INV        g0988(.A(new_new_n1010_), .Y(new_new_n1011_));
  NA3        g0989(.A(new_new_n1011_), .B(new_new_n1008_), .C(new_new_n1007_), .Y(new_new_n1012_));
  NO4        g0990(.A(new_new_n228_), .B(new_new_n149_), .C(new_new_n678_), .D(new_new_n37_), .Y(new_new_n1013_));
  NO2        g0991(.A(new_new_n1013_), .B(new_new_n883_), .Y(new_new_n1014_));
  INV        g0992(.A(new_new_n1014_), .Y(new_new_n1015_));
  AOI210     g0993(.A0(new_new_n1012_), .A1(new_new_n49_), .B0(new_new_n1015_), .Y(new_new_n1016_));
  AOI210     g0994(.A0(new_new_n1016_), .A1(new_new_n1005_), .B0(new_new_n74_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n564_), .B(new_new_n384_), .Y(new_new_n1018_));
  NO2        g0996(.A(new_new_n1018_), .B(new_new_n755_), .Y(new_new_n1019_));
  OAI210     g0997(.A0(new_new_n81_), .A1(new_new_n55_), .B0(new_new_n112_), .Y(new_new_n1020_));
  NA2        g0998(.A(new_new_n1020_), .B(new_new_n77_), .Y(new_new_n1021_));
  AOI210     g0999(.A0(new_new_n979_), .A1(new_new_n899_), .B0(new_new_n915_), .Y(new_new_n1022_));
  AOI210     g1000(.A0(new_new_n1022_), .A1(new_new_n1021_), .B0(new_new_n678_), .Y(new_new_n1023_));
  NA2        g1001(.A(new_new_n260_), .B(new_new_n58_), .Y(new_new_n1024_));
  AOI220     g1002(.A0(new_new_n1024_), .A1(new_new_n77_), .B0(new_new_n351_), .B1(new_new_n252_), .Y(new_new_n1025_));
  NO2        g1003(.A(new_new_n1025_), .B(new_new_n232_), .Y(new_new_n1026_));
  NA3        g1004(.A(new_new_n100_), .B(new_new_n310_), .C(new_new_n31_), .Y(new_new_n1027_));
  INV        g1005(.A(new_new_n1027_), .Y(new_new_n1028_));
  NO3        g1006(.A(new_new_n1028_), .B(new_new_n1026_), .C(new_new_n1023_), .Y(new_new_n1029_));
  OAI210     g1007(.A0(new_new_n268_), .A1(new_new_n158_), .B0(new_new_n90_), .Y(new_new_n1030_));
  NA3        g1008(.A(new_new_n759_), .B(new_new_n292_), .C(new_new_n81_), .Y(new_new_n1031_));
  AOI210     g1009(.A0(new_new_n1031_), .A1(new_new_n1030_), .B0(i_11_), .Y(new_new_n1032_));
  NO3        g1010(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n1033_));
  OAI210     g1011(.A0(new_new_n919_), .A1(new_new_n310_), .B0(new_new_n1033_), .Y(new_new_n1034_));
  NO2        g1012(.A(new_new_n1034_), .B(new_new_n726_), .Y(new_new_n1035_));
  NO4        g1013(.A(new_new_n941_), .B(new_new_n477_), .C(new_new_n249_), .D(new_new_n248_), .Y(new_new_n1036_));
  NO2        g1014(.A(new_new_n1036_), .B(new_new_n561_), .Y(new_new_n1037_));
  NO2        g1015(.A(new_new_n1037_), .B(new_new_n41_), .Y(new_new_n1038_));
  NO3        g1016(.A(new_new_n1038_), .B(new_new_n1035_), .C(new_new_n1032_), .Y(new_new_n1039_));
  OAI210     g1017(.A0(new_new_n1029_), .A1(i_4_), .B0(new_new_n1039_), .Y(new_new_n1040_));
  NO3        g1018(.A(new_new_n1040_), .B(new_new_n1019_), .C(new_new_n1017_), .Y(new_new_n1041_));
  NA4        g1019(.A(new_new_n1041_), .B(new_new_n1001_), .C(new_new_n948_), .D(new_new_n871_), .Y(mai4));
  INV        g1020(.A(new_new_n698_), .Y(new_new_n1045_));
endmodule


