// Benchmark "top" written by ABC on Thu Jun 20 14:59:12 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n141_, new_new_n142_, new_new_n143_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n776_, new_new_n777_,
    new_new_n778_, new_new_n779_, new_new_n780_, new_new_n781_,
    new_new_n782_, new_new_n783_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n825_, new_new_n826_,
    new_new_n827_, new_new_n828_, new_new_n829_, new_new_n830_,
    new_new_n831_, new_new_n832_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n875_,
    new_new_n876_, new_new_n877_, new_new_n878_, new_new_n879_,
    new_new_n880_, new_new_n881_, new_new_n882_, new_new_n883_,
    new_new_n884_, new_new_n885_, new_new_n886_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1100_,
    new_new_n1101_, new_new_n1102_, new_new_n1103_, new_new_n1104_,
    new_new_n1105_, new_new_n1106_, new_new_n1110_, new_new_n1111_,
    new_new_n1112_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  OR4        g0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g0067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  NO2        g0068(.A(new_new_n89_), .B(new_new_n90_), .Y(new_new_n91_));
  OAI210     g0069(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n91_), .Y(new_new_n92_));
  NAi21      g0070(.An(i_6_), .B(i_10_), .Y(new_new_n93_));
  NA2        g0071(.A(i_6_), .B(i_9_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n93_), .B0(new_new_n64_), .Y(new_new_n95_));
  NA2        g0073(.A(i_2_), .B(i_6_), .Y(new_new_n96_));
  NO3        g0074(.A(new_new_n96_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n97_));
  NO2        g0075(.A(new_new_n97_), .B(new_new_n95_), .Y(new_new_n98_));
  AOI210     g0076(.A0(new_new_n98_), .A1(new_new_n92_), .B0(new_new_n81_), .Y(new_new_n99_));
  AN3        g0077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n100_));
  NAi21      g0078(.An(i_6_), .B(i_11_), .Y(new_new_n101_));
  NO2        g0079(.A(i_5_), .B(i_8_), .Y(new_new_n102_));
  NOi21      g0080(.An(new_new_n102_), .B(new_new_n101_), .Y(new_new_n103_));
  AOI220     g0081(.A0(new_new_n103_), .A1(new_new_n63_), .B0(new_new_n100_), .B1(new_new_n32_), .Y(new_new_n104_));
  INV        g0082(.A(i_7_), .Y(new_new_n105_));
  NA2        g0083(.A(new_new_n47_), .B(new_new_n105_), .Y(new_new_n106_));
  NO2        g0084(.A(i_0_), .B(i_5_), .Y(new_new_n107_));
  NO2        g0085(.A(new_new_n107_), .B(new_new_n87_), .Y(new_new_n108_));
  NA2        g0086(.A(i_12_), .B(i_3_), .Y(new_new_n109_));
  INV        g0087(.A(new_new_n109_), .Y(new_new_n110_));
  NA3        g0088(.A(new_new_n110_), .B(new_new_n108_), .C(new_new_n106_), .Y(new_new_n111_));
  NAi21      g0089(.An(i_7_), .B(i_11_), .Y(new_new_n112_));
  AN2        g0090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g0091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g0092(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n115_));
  NO2        g0093(.A(i_8_), .B(new_new_n105_), .Y(new_new_n116_));
  NO3        g0094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g0095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g0097(.A(i_11_), .B(i_12_), .Y(new_new_n120_));
  INV        g0098(.A(new_new_n120_), .Y(new_new_n121_));
  NO2        g0099(.A(new_new_n121_), .B(new_new_n117_), .Y(new_new_n122_));
  NA3        g0100(.A(new_new_n122_), .B(new_new_n111_), .C(new_new_n104_), .Y(new_new_n123_));
  NOi21      g0101(.An(i_1_), .B(i_5_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(i_11_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n126_));
  NA2        g0104(.A(i_7_), .B(new_new_n25_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n127_), .B(new_new_n126_), .Y(new_new_n128_));
  NO2        g0106(.A(new_new_n128_), .B(new_new_n47_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n94_), .B(new_new_n93_), .Y(new_new_n130_));
  NAi21      g0108(.An(i_3_), .B(i_8_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n131_), .B(new_new_n63_), .Y(new_new_n132_));
  NOi31      g0110(.An(new_new_n132_), .B(new_new_n130_), .C(new_new_n129_), .Y(new_new_n133_));
  NO2        g0111(.A(i_1_), .B(new_new_n87_), .Y(new_new_n134_));
  NO2        g0112(.A(i_6_), .B(i_5_), .Y(new_new_n135_));
  NA2        g0113(.A(new_new_n135_), .B(i_3_), .Y(new_new_n136_));
  AO210      g0114(.A0(new_new_n136_), .A1(new_new_n48_), .B0(new_new_n134_), .Y(new_new_n137_));
  OAI220     g0115(.A0(new_new_n137_), .A1(new_new_n112_), .B0(new_new_n133_), .B1(new_new_n125_), .Y(new_new_n138_));
  NO3        g0116(.A(new_new_n138_), .B(new_new_n123_), .C(new_new_n99_), .Y(new_new_n139_));
  NA3        g0117(.A(new_new_n139_), .B(new_new_n80_), .C(new_new_n57_), .Y(men2));
  NO2        g0118(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n141_));
  NA2        g0119(.A(i_6_), .B(new_new_n25_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(new_new_n141_), .Y(new_new_n143_));
  NA4        g0121(.A(new_new_n143_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(men0));
  AN2        g0122(.A(i_8_), .B(i_7_), .Y(new_new_n145_));
  NA2        g0123(.A(new_new_n145_), .B(i_6_), .Y(new_new_n146_));
  NO2        g0124(.A(i_12_), .B(i_13_), .Y(new_new_n147_));
  NAi21      g0125(.An(i_5_), .B(i_11_), .Y(new_new_n148_));
  NOi21      g0126(.An(new_new_n147_), .B(new_new_n148_), .Y(new_new_n149_));
  NO2        g0127(.A(i_0_), .B(i_1_), .Y(new_new_n150_));
  NA2        g0128(.A(i_2_), .B(i_3_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(i_4_), .Y(new_new_n152_));
  NA3        g0130(.A(new_new_n152_), .B(new_new_n150_), .C(new_new_n149_), .Y(new_new_n153_));
  OR2        g0131(.A(new_new_n153_), .B(new_new_n25_), .Y(new_new_n154_));
  AN2        g0132(.A(new_new_n147_), .B(new_new_n84_), .Y(new_new_n155_));
  NO2        g0133(.A(new_new_n155_), .B(new_new_n27_), .Y(new_new_n156_));
  NA2        g0134(.A(i_1_), .B(i_5_), .Y(new_new_n157_));
  NO2        g0135(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n158_));
  NA2        g0136(.A(new_new_n158_), .B(new_new_n36_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n159_), .B(new_new_n157_), .C(new_new_n156_), .Y(new_new_n160_));
  OR2        g0138(.A(i_0_), .B(i_1_), .Y(new_new_n161_));
  NO3        g0139(.A(new_new_n161_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n162_));
  NAi32      g0140(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n163_));
  NAi21      g0141(.An(new_new_n163_), .B(new_new_n162_), .Y(new_new_n164_));
  NOi21      g0142(.An(i_4_), .B(i_10_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n40_), .Y(new_new_n166_));
  NO2        g0144(.A(i_3_), .B(i_5_), .Y(new_new_n167_));
  NO3        g0145(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n168_));
  NA2        g0146(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n169_));
  OAI210     g0147(.A0(new_new_n169_), .A1(new_new_n166_), .B0(new_new_n164_), .Y(new_new_n170_));
  NO2        g0148(.A(new_new_n170_), .B(new_new_n160_), .Y(new_new_n171_));
  AOI210     g0149(.A0(new_new_n171_), .A1(new_new_n154_), .B0(new_new_n146_), .Y(new_new_n172_));
  NA3        g0150(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n173_));
  NA2        g0151(.A(i_3_), .B(new_new_n49_), .Y(new_new_n174_));
  NOi21      g0152(.An(i_4_), .B(i_9_), .Y(new_new_n175_));
  NOi21      g0153(.An(i_11_), .B(i_13_), .Y(new_new_n176_));
  NA2        g0154(.A(new_new_n176_), .B(new_new_n175_), .Y(new_new_n177_));
  OR2        g0155(.A(new_new_n177_), .B(new_new_n174_), .Y(new_new_n178_));
  NO2        g0156(.A(i_4_), .B(i_5_), .Y(new_new_n179_));
  NAi21      g0157(.An(i_12_), .B(i_11_), .Y(new_new_n180_));
  NO2        g0158(.A(new_new_n180_), .B(i_13_), .Y(new_new_n181_));
  NA3        g0159(.A(new_new_n181_), .B(new_new_n179_), .C(new_new_n84_), .Y(new_new_n182_));
  AOI210     g0160(.A0(new_new_n182_), .A1(new_new_n178_), .B0(new_new_n173_), .Y(new_new_n183_));
  NO2        g0161(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n184_));
  NA2        g0162(.A(new_new_n184_), .B(new_new_n47_), .Y(new_new_n185_));
  NA2        g0163(.A(new_new_n36_), .B(i_5_), .Y(new_new_n186_));
  NAi31      g0164(.An(new_new_n186_), .B(new_new_n155_), .C(i_11_), .Y(new_new_n187_));
  NA2        g0165(.A(i_3_), .B(i_5_), .Y(new_new_n188_));
  OR2        g0166(.A(new_new_n188_), .B(new_new_n177_), .Y(new_new_n189_));
  AOI210     g0167(.A0(new_new_n189_), .A1(new_new_n187_), .B0(new_new_n185_), .Y(new_new_n190_));
  NO2        g0168(.A(new_new_n74_), .B(i_5_), .Y(new_new_n191_));
  NO2        g0169(.A(i_13_), .B(i_10_), .Y(new_new_n192_));
  NA3        g0170(.A(new_new_n192_), .B(new_new_n191_), .C(new_new_n45_), .Y(new_new_n193_));
  NO2        g0171(.A(i_2_), .B(i_1_), .Y(new_new_n194_));
  NA2        g0172(.A(new_new_n194_), .B(i_3_), .Y(new_new_n195_));
  NAi21      g0173(.An(i_4_), .B(i_12_), .Y(new_new_n196_));
  NO4        g0174(.A(new_new_n196_), .B(new_new_n195_), .C(new_new_n193_), .D(new_new_n25_), .Y(new_new_n197_));
  NO3        g0175(.A(new_new_n197_), .B(new_new_n190_), .C(new_new_n183_), .Y(new_new_n198_));
  INV        g0176(.A(i_8_), .Y(new_new_n199_));
  NO2        g0177(.A(new_new_n199_), .B(i_7_), .Y(new_new_n200_));
  NA2        g0178(.A(new_new_n200_), .B(i_6_), .Y(new_new_n201_));
  NO3        g0179(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n202_));
  NA2        g0180(.A(new_new_n202_), .B(new_new_n116_), .Y(new_new_n203_));
  NO3        g0181(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n204_));
  NA3        g0182(.A(new_new_n204_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n205_));
  NO3        g0183(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n206_));
  OAI210     g0184(.A0(new_new_n100_), .A1(i_12_), .B0(new_new_n206_), .Y(new_new_n207_));
  AOI210     g0185(.A0(new_new_n207_), .A1(new_new_n205_), .B0(new_new_n203_), .Y(new_new_n208_));
  NO2        g0186(.A(i_3_), .B(i_8_), .Y(new_new_n209_));
  NO3        g0187(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n210_));
  NA3        g0188(.A(new_new_n210_), .B(new_new_n209_), .C(new_new_n40_), .Y(new_new_n211_));
  NO2        g0189(.A(new_new_n107_), .B(new_new_n59_), .Y(new_new_n212_));
  INV        g0190(.A(new_new_n212_), .Y(new_new_n213_));
  NO2        g0191(.A(i_13_), .B(i_9_), .Y(new_new_n214_));
  NA3        g0192(.A(new_new_n214_), .B(i_6_), .C(new_new_n199_), .Y(new_new_n215_));
  NAi21      g0193(.An(i_12_), .B(i_3_), .Y(new_new_n216_));
  OR2        g0194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n45_), .B(i_5_), .Y(new_new_n218_));
  NO3        g0196(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n219_));
  NA3        g0197(.A(new_new_n219_), .B(new_new_n218_), .C(i_10_), .Y(new_new_n220_));
  OAI220     g0198(.A0(new_new_n220_), .A1(new_new_n217_), .B0(new_new_n213_), .B1(new_new_n211_), .Y(new_new_n221_));
  AOI210     g0199(.A0(new_new_n221_), .A1(i_7_), .B0(new_new_n208_), .Y(new_new_n222_));
  OAI220     g0200(.A0(new_new_n222_), .A1(i_4_), .B0(new_new_n201_), .B1(new_new_n198_), .Y(new_new_n223_));
  NAi21      g0201(.An(i_12_), .B(i_7_), .Y(new_new_n224_));
  NA3        g0202(.A(i_13_), .B(new_new_n199_), .C(i_10_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  NA2        g0204(.A(i_0_), .B(i_5_), .Y(new_new_n227_));
  NA2        g0205(.A(new_new_n227_), .B(new_new_n108_), .Y(new_new_n228_));
  OAI220     g0206(.A0(new_new_n228_), .A1(new_new_n195_), .B0(new_new_n185_), .B1(new_new_n136_), .Y(new_new_n229_));
  NAi31      g0207(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n36_), .B(i_13_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n233_));
  NA3        g0211(.A(new_new_n233_), .B(new_new_n232_), .C(new_new_n231_), .Y(new_new_n234_));
  INV        g0212(.A(i_13_), .Y(new_new_n235_));
  NO2        g0213(.A(i_12_), .B(new_new_n235_), .Y(new_new_n236_));
  NA3        g0214(.A(new_new_n236_), .B(new_new_n204_), .C(new_new_n202_), .Y(new_new_n237_));
  OAI210     g0215(.A0(new_new_n234_), .A1(new_new_n230_), .B0(new_new_n237_), .Y(new_new_n238_));
  AOI220     g0216(.A0(new_new_n238_), .A1(new_new_n145_), .B0(new_new_n229_), .B1(new_new_n226_), .Y(new_new_n239_));
  NO2        g0217(.A(i_12_), .B(new_new_n37_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n188_), .B(i_4_), .Y(new_new_n241_));
  NA2        g0219(.A(new_new_n241_), .B(new_new_n240_), .Y(new_new_n242_));
  OR2        g0220(.A(i_8_), .B(i_7_), .Y(new_new_n243_));
  NO2        g0221(.A(new_new_n243_), .B(new_new_n87_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n54_), .B(i_1_), .Y(new_new_n245_));
  NA2        g0223(.A(new_new_n245_), .B(new_new_n244_), .Y(new_new_n246_));
  INV        g0224(.A(i_12_), .Y(new_new_n247_));
  NO2        g0225(.A(new_new_n45_), .B(new_new_n247_), .Y(new_new_n248_));
  NO3        g0226(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n249_));
  NA2        g0227(.A(i_2_), .B(i_1_), .Y(new_new_n250_));
  NO2        g0228(.A(new_new_n246_), .B(new_new_n242_), .Y(new_new_n251_));
  NO3        g0229(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n252_));
  NAi21      g0230(.An(i_4_), .B(i_3_), .Y(new_new_n253_));
  NO2        g0231(.A(new_new_n253_), .B(new_new_n76_), .Y(new_new_n254_));
  NO2        g0232(.A(i_0_), .B(i_6_), .Y(new_new_n255_));
  NOi41      g0233(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n256_), .B(new_new_n255_), .Y(new_new_n257_));
  NO2        g0235(.A(new_new_n250_), .B(new_new_n188_), .Y(new_new_n258_));
  NAi21      g0236(.An(new_new_n257_), .B(new_new_n258_), .Y(new_new_n259_));
  INV        g0237(.A(new_new_n259_), .Y(new_new_n260_));
  AOI220     g0238(.A0(new_new_n260_), .A1(new_new_n40_), .B0(new_new_n251_), .B1(new_new_n214_), .Y(new_new_n261_));
  NO2        g0239(.A(i_11_), .B(new_new_n235_), .Y(new_new_n262_));
  NOi21      g0240(.An(i_1_), .B(i_6_), .Y(new_new_n263_));
  NAi21      g0241(.An(i_3_), .B(i_7_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n247_), .B(i_9_), .Y(new_new_n265_));
  OR4        g0243(.A(new_new_n265_), .B(new_new_n264_), .C(new_new_n263_), .D(new_new_n191_), .Y(new_new_n266_));
  NO2        g0244(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n267_));
  NO2        g0245(.A(i_12_), .B(i_3_), .Y(new_new_n268_));
  NA2        g0246(.A(new_new_n74_), .B(i_5_), .Y(new_new_n269_));
  NA2        g0247(.A(i_3_), .B(i_9_), .Y(new_new_n270_));
  NAi21      g0248(.An(i_7_), .B(i_10_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n271_), .B(new_new_n270_), .Y(new_new_n272_));
  NA3        g0250(.A(new_new_n272_), .B(new_new_n269_), .C(new_new_n65_), .Y(new_new_n273_));
  NA2        g0251(.A(new_new_n273_), .B(new_new_n266_), .Y(new_new_n274_));
  NA3        g0252(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n275_));
  INV        g0253(.A(new_new_n146_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n247_), .B(i_13_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n277_), .B(new_new_n76_), .Y(new_new_n278_));
  AOI220     g0256(.A0(new_new_n278_), .A1(new_new_n276_), .B0(new_new_n274_), .B1(new_new_n262_), .Y(new_new_n279_));
  NO2        g0257(.A(new_new_n243_), .B(new_new_n37_), .Y(new_new_n280_));
  NA2        g0258(.A(i_12_), .B(i_6_), .Y(new_new_n281_));
  OR2        g0259(.A(i_13_), .B(i_9_), .Y(new_new_n282_));
  NO3        g0260(.A(new_new_n282_), .B(new_new_n281_), .C(new_new_n49_), .Y(new_new_n283_));
  NO2        g0261(.A(new_new_n253_), .B(i_2_), .Y(new_new_n284_));
  NA3        g0262(.A(new_new_n284_), .B(new_new_n283_), .C(new_new_n45_), .Y(new_new_n285_));
  NA2        g0263(.A(new_new_n262_), .B(i_9_), .Y(new_new_n286_));
  NA2        g0264(.A(new_new_n269_), .B(new_new_n65_), .Y(new_new_n287_));
  OAI210     g0265(.A0(new_new_n287_), .A1(new_new_n286_), .B0(new_new_n285_), .Y(new_new_n288_));
  NA2        g0266(.A(new_new_n158_), .B(new_new_n64_), .Y(new_new_n289_));
  NO3        g0267(.A(i_11_), .B(new_new_n235_), .C(new_new_n25_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n264_), .B(i_8_), .Y(new_new_n291_));
  NO2        g0269(.A(i_6_), .B(new_new_n49_), .Y(new_new_n292_));
  NA3        g0270(.A(new_new_n292_), .B(new_new_n291_), .C(new_new_n290_), .Y(new_new_n293_));
  NO3        g0271(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n294_));
  NA3        g0272(.A(new_new_n294_), .B(new_new_n280_), .C(new_new_n236_), .Y(new_new_n295_));
  AOI210     g0273(.A0(new_new_n295_), .A1(new_new_n293_), .B0(new_new_n289_), .Y(new_new_n296_));
  AOI210     g0274(.A0(new_new_n288_), .A1(new_new_n280_), .B0(new_new_n296_), .Y(new_new_n297_));
  NA4        g0275(.A(new_new_n297_), .B(new_new_n279_), .C(new_new_n261_), .D(new_new_n239_), .Y(new_new_n298_));
  NO3        g0276(.A(i_12_), .B(new_new_n235_), .C(new_new_n37_), .Y(new_new_n299_));
  INV        g0277(.A(new_new_n299_), .Y(new_new_n300_));
  NA2        g0278(.A(i_8_), .B(new_new_n105_), .Y(new_new_n301_));
  NOi21      g0279(.An(new_new_n167_), .B(new_new_n87_), .Y(new_new_n302_));
  NO3        g0280(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n303_));
  AOI220     g0281(.A0(new_new_n303_), .A1(new_new_n202_), .B0(new_new_n302_), .B1(new_new_n245_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n304_), .B(new_new_n301_), .Y(new_new_n305_));
  NO3        g0283(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n306_));
  NO2        g0284(.A(new_new_n250_), .B(i_0_), .Y(new_new_n307_));
  AOI220     g0285(.A0(new_new_n307_), .A1(new_new_n200_), .B0(new_new_n306_), .B1(new_new_n145_), .Y(new_new_n308_));
  NA2        g0286(.A(new_new_n292_), .B(new_new_n26_), .Y(new_new_n309_));
  NO2        g0287(.A(new_new_n309_), .B(new_new_n308_), .Y(new_new_n310_));
  NA2        g0288(.A(i_0_), .B(i_1_), .Y(new_new_n311_));
  NO2        g0289(.A(new_new_n311_), .B(i_2_), .Y(new_new_n312_));
  NO2        g0290(.A(new_new_n60_), .B(i_6_), .Y(new_new_n313_));
  NA3        g0291(.A(new_new_n313_), .B(new_new_n312_), .C(new_new_n167_), .Y(new_new_n314_));
  OAI210     g0292(.A0(new_new_n169_), .A1(new_new_n146_), .B0(new_new_n314_), .Y(new_new_n315_));
  NO3        g0293(.A(new_new_n315_), .B(new_new_n310_), .C(new_new_n305_), .Y(new_new_n316_));
  NO2        g0294(.A(i_3_), .B(i_10_), .Y(new_new_n317_));
  NA3        g0295(.A(new_new_n317_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n318_));
  NO2        g0296(.A(i_2_), .B(new_new_n105_), .Y(new_new_n319_));
  NA2        g0297(.A(i_1_), .B(new_new_n36_), .Y(new_new_n320_));
  NO2        g0298(.A(new_new_n320_), .B(i_8_), .Y(new_new_n321_));
  NOi21      g0299(.An(new_new_n227_), .B(new_new_n107_), .Y(new_new_n322_));
  NA3        g0300(.A(new_new_n322_), .B(new_new_n321_), .C(new_new_n319_), .Y(new_new_n323_));
  AN2        g0301(.A(i_3_), .B(i_10_), .Y(new_new_n324_));
  NA4        g0302(.A(new_new_n324_), .B(new_new_n204_), .C(new_new_n181_), .D(new_new_n179_), .Y(new_new_n325_));
  NO2        g0303(.A(i_5_), .B(new_new_n37_), .Y(new_new_n326_));
  NO2        g0304(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n327_));
  OR2        g0305(.A(new_new_n323_), .B(new_new_n318_), .Y(new_new_n328_));
  OAI220     g0306(.A0(new_new_n328_), .A1(i_6_), .B0(new_new_n316_), .B1(new_new_n300_), .Y(new_new_n329_));
  NO4        g0307(.A(new_new_n329_), .B(new_new_n298_), .C(new_new_n223_), .D(new_new_n172_), .Y(new_new_n330_));
  NO3        g0308(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n331_));
  NO2        g0309(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n332_));
  NA2        g0310(.A(new_new_n307_), .B(new_new_n332_), .Y(new_new_n333_));
  NO3        g0311(.A(i_6_), .B(new_new_n199_), .C(i_7_), .Y(new_new_n334_));
  NA2        g0312(.A(new_new_n334_), .B(new_new_n204_), .Y(new_new_n335_));
  AOI210     g0313(.A0(new_new_n335_), .A1(new_new_n333_), .B0(new_new_n174_), .Y(new_new_n336_));
  NO2        g0314(.A(i_2_), .B(i_3_), .Y(new_new_n337_));
  OR2        g0315(.A(i_0_), .B(i_5_), .Y(new_new_n338_));
  NA2        g0316(.A(new_new_n227_), .B(new_new_n338_), .Y(new_new_n339_));
  NA4        g0317(.A(new_new_n339_), .B(new_new_n244_), .C(new_new_n337_), .D(i_1_), .Y(new_new_n340_));
  NA3        g0318(.A(new_new_n307_), .B(new_new_n302_), .C(new_new_n116_), .Y(new_new_n341_));
  NAi21      g0319(.An(i_8_), .B(i_7_), .Y(new_new_n342_));
  NO2        g0320(.A(new_new_n342_), .B(i_6_), .Y(new_new_n343_));
  NO2        g0321(.A(new_new_n161_), .B(new_new_n47_), .Y(new_new_n344_));
  NA3        g0322(.A(new_new_n344_), .B(new_new_n343_), .C(new_new_n167_), .Y(new_new_n345_));
  NA3        g0323(.A(new_new_n345_), .B(new_new_n341_), .C(new_new_n340_), .Y(new_new_n346_));
  OAI210     g0324(.A0(new_new_n346_), .A1(new_new_n336_), .B0(i_4_), .Y(new_new_n347_));
  NO2        g0325(.A(i_12_), .B(i_10_), .Y(new_new_n348_));
  NOi21      g0326(.An(i_5_), .B(i_0_), .Y(new_new_n349_));
  NO3        g0327(.A(new_new_n320_), .B(new_new_n349_), .C(new_new_n131_), .Y(new_new_n350_));
  NA4        g0328(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n351_));
  NA2        g0329(.A(new_new_n350_), .B(new_new_n348_), .Y(new_new_n352_));
  NO2        g0330(.A(i_6_), .B(i_8_), .Y(new_new_n353_));
  NOi21      g0331(.An(i_0_), .B(i_2_), .Y(new_new_n354_));
  AN2        g0332(.A(new_new_n354_), .B(new_new_n353_), .Y(new_new_n355_));
  NO2        g0333(.A(i_1_), .B(i_7_), .Y(new_new_n356_));
  AO220      g0334(.A0(new_new_n356_), .A1(new_new_n355_), .B0(new_new_n343_), .B1(new_new_n245_), .Y(new_new_n357_));
  NA3        g0335(.A(new_new_n357_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n358_));
  NA3        g0336(.A(new_new_n358_), .B(new_new_n352_), .C(new_new_n347_), .Y(new_new_n359_));
  NO3        g0337(.A(new_new_n243_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n360_));
  NO3        g0338(.A(new_new_n342_), .B(i_2_), .C(i_1_), .Y(new_new_n361_));
  OAI210     g0339(.A0(new_new_n361_), .A1(new_new_n360_), .B0(i_6_), .Y(new_new_n362_));
  NA3        g0340(.A(new_new_n263_), .B(new_new_n319_), .C(new_new_n199_), .Y(new_new_n363_));
  AOI210     g0341(.A0(new_new_n363_), .A1(new_new_n362_), .B0(new_new_n339_), .Y(new_new_n364_));
  NOi21      g0342(.An(new_new_n157_), .B(new_new_n108_), .Y(new_new_n365_));
  NA2        g0343(.A(new_new_n364_), .B(i_3_), .Y(new_new_n366_));
  INV        g0344(.A(new_new_n85_), .Y(new_new_n367_));
  NO2        g0345(.A(new_new_n311_), .B(new_new_n82_), .Y(new_new_n368_));
  NA2        g0346(.A(new_new_n368_), .B(new_new_n135_), .Y(new_new_n369_));
  NO2        g0347(.A(new_new_n96_), .B(new_new_n199_), .Y(new_new_n370_));
  NA3        g0348(.A(new_new_n322_), .B(new_new_n370_), .C(new_new_n64_), .Y(new_new_n371_));
  AOI210     g0349(.A0(new_new_n371_), .A1(new_new_n369_), .B0(new_new_n367_), .Y(new_new_n372_));
  NO2        g0350(.A(new_new_n199_), .B(i_9_), .Y(new_new_n373_));
  NA2        g0351(.A(new_new_n373_), .B(new_new_n212_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n372_), .B(new_new_n310_), .Y(new_new_n375_));
  AOI210     g0353(.A0(new_new_n375_), .A1(new_new_n366_), .B0(new_new_n166_), .Y(new_new_n376_));
  AOI210     g0354(.A0(new_new_n359_), .A1(new_new_n331_), .B0(new_new_n376_), .Y(new_new_n377_));
  NOi32      g0355(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n378_));
  INV        g0356(.A(new_new_n378_), .Y(new_new_n379_));
  NAi21      g0357(.An(i_0_), .B(i_6_), .Y(new_new_n380_));
  NAi21      g0358(.An(i_1_), .B(i_5_), .Y(new_new_n381_));
  NA2        g0359(.A(new_new_n381_), .B(new_new_n380_), .Y(new_new_n382_));
  NA2        g0360(.A(new_new_n382_), .B(new_new_n25_), .Y(new_new_n383_));
  OAI210     g0361(.A0(new_new_n383_), .A1(new_new_n163_), .B0(new_new_n257_), .Y(new_new_n384_));
  NAi41      g0362(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n385_));
  AOI210     g0363(.A0(new_new_n385_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n386_));
  NOi32      g0364(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n387_));
  NO2        g0365(.A(i_1_), .B(new_new_n105_), .Y(new_new_n388_));
  NAi21      g0366(.An(i_3_), .B(i_4_), .Y(new_new_n389_));
  NO2        g0367(.A(new_new_n389_), .B(i_9_), .Y(new_new_n390_));
  AN2        g0368(.A(i_6_), .B(i_7_), .Y(new_new_n391_));
  OAI210     g0369(.A0(new_new_n391_), .A1(new_new_n388_), .B0(new_new_n390_), .Y(new_new_n392_));
  NA2        g0370(.A(i_2_), .B(i_7_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n389_), .B(i_10_), .Y(new_new_n394_));
  NA3        g0372(.A(new_new_n394_), .B(new_new_n393_), .C(new_new_n255_), .Y(new_new_n395_));
  AOI210     g0373(.A0(new_new_n395_), .A1(new_new_n392_), .B0(new_new_n191_), .Y(new_new_n396_));
  AOI210     g0374(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n397_));
  OAI210     g0375(.A0(new_new_n397_), .A1(new_new_n194_), .B0(new_new_n394_), .Y(new_new_n398_));
  AOI220     g0376(.A0(new_new_n394_), .A1(new_new_n356_), .B0(new_new_n249_), .B1(new_new_n194_), .Y(new_new_n399_));
  AOI210     g0377(.A0(new_new_n399_), .A1(new_new_n398_), .B0(i_5_), .Y(new_new_n400_));
  NO4        g0378(.A(new_new_n400_), .B(new_new_n396_), .C(new_new_n386_), .D(new_new_n384_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n401_), .B(new_new_n379_), .Y(new_new_n402_));
  NO2        g0380(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n403_));
  AN2        g0381(.A(i_12_), .B(i_5_), .Y(new_new_n404_));
  NO2        g0382(.A(i_4_), .B(new_new_n26_), .Y(new_new_n405_));
  NA2        g0383(.A(new_new_n405_), .B(new_new_n404_), .Y(new_new_n406_));
  NO2        g0384(.A(i_11_), .B(i_6_), .Y(new_new_n407_));
  NA3        g0385(.A(new_new_n407_), .B(new_new_n344_), .C(new_new_n235_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n408_), .B(new_new_n406_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n253_), .B(i_5_), .Y(new_new_n410_));
  NO2        g0388(.A(i_5_), .B(i_10_), .Y(new_new_n411_));
  AOI220     g0389(.A0(new_new_n411_), .A1(new_new_n284_), .B0(new_new_n410_), .B1(new_new_n204_), .Y(new_new_n412_));
  NA2        g0390(.A(new_new_n147_), .B(new_new_n46_), .Y(new_new_n413_));
  NO2        g0391(.A(new_new_n413_), .B(new_new_n412_), .Y(new_new_n414_));
  OAI210     g0392(.A0(new_new_n414_), .A1(new_new_n409_), .B0(new_new_n403_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n153_), .B(new_new_n87_), .Y(new_new_n417_));
  OAI210     g0395(.A0(new_new_n417_), .A1(new_new_n409_), .B0(new_new_n416_), .Y(new_new_n418_));
  NO3        g0396(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n419_));
  NO2        g0397(.A(i_11_), .B(i_12_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n411_), .B(new_new_n247_), .Y(new_new_n421_));
  NA3        g0399(.A(new_new_n116_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n422_));
  OAI220     g0400(.A0(new_new_n422_), .A1(new_new_n230_), .B0(new_new_n421_), .B1(new_new_n351_), .Y(new_new_n423_));
  NAi21      g0401(.An(i_13_), .B(i_0_), .Y(new_new_n424_));
  NO2        g0402(.A(new_new_n424_), .B(new_new_n250_), .Y(new_new_n425_));
  NA2        g0403(.A(new_new_n423_), .B(new_new_n425_), .Y(new_new_n426_));
  NA3        g0404(.A(new_new_n426_), .B(new_new_n418_), .C(new_new_n415_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n45_), .B(new_new_n235_), .Y(new_new_n428_));
  NO3        g0406(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n429_));
  NO2        g0407(.A(i_0_), .B(i_11_), .Y(new_new_n430_));
  INV        g0408(.A(i_5_), .Y(new_new_n431_));
  AN2        g0409(.A(i_1_), .B(i_6_), .Y(new_new_n432_));
  NOi21      g0410(.An(i_2_), .B(i_12_), .Y(new_new_n433_));
  NA2        g0411(.A(new_new_n433_), .B(new_new_n432_), .Y(new_new_n434_));
  NO2        g0412(.A(new_new_n434_), .B(new_new_n431_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n145_), .B(i_9_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n436_), .B(i_4_), .Y(new_new_n437_));
  NA2        g0415(.A(new_new_n435_), .B(new_new_n437_), .Y(new_new_n438_));
  NAi21      g0416(.An(i_9_), .B(i_4_), .Y(new_new_n439_));
  OR2        g0417(.A(i_13_), .B(i_10_), .Y(new_new_n440_));
  NO3        g0418(.A(new_new_n440_), .B(new_new_n120_), .C(new_new_n439_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n177_), .B(new_new_n126_), .Y(new_new_n442_));
  OR2        g0420(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n443_));
  NO2        g0421(.A(new_new_n105_), .B(new_new_n25_), .Y(new_new_n444_));
  NA2        g0422(.A(new_new_n299_), .B(new_new_n444_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n292_), .B(new_new_n219_), .Y(new_new_n446_));
  OAI220     g0424(.A0(new_new_n446_), .A1(new_new_n443_), .B0(new_new_n445_), .B1(new_new_n365_), .Y(new_new_n447_));
  INV        g0425(.A(new_new_n447_), .Y(new_new_n448_));
  AOI210     g0426(.A0(new_new_n448_), .A1(new_new_n438_), .B0(new_new_n26_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n341_), .B(new_new_n340_), .Y(new_new_n450_));
  AOI220     g0428(.A0(new_new_n313_), .A1(new_new_n303_), .B0(new_new_n307_), .B1(new_new_n332_), .Y(new_new_n451_));
  NO2        g0429(.A(new_new_n451_), .B(new_new_n174_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n188_), .B(new_new_n87_), .Y(new_new_n453_));
  AOI220     g0431(.A0(new_new_n453_), .A1(new_new_n312_), .B0(new_new_n294_), .B1(new_new_n219_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n454_), .B(new_new_n301_), .Y(new_new_n455_));
  NO3        g0433(.A(new_new_n455_), .B(new_new_n452_), .C(new_new_n450_), .Y(new_new_n456_));
  NA2        g0434(.A(new_new_n202_), .B(new_new_n100_), .Y(new_new_n457_));
  NA3        g0435(.A(new_new_n344_), .B(new_new_n167_), .C(new_new_n87_), .Y(new_new_n458_));
  AOI210     g0436(.A0(new_new_n458_), .A1(new_new_n457_), .B0(new_new_n342_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n313_), .B(new_new_n245_), .Y(new_new_n460_));
  NO2        g0438(.A(new_new_n460_), .B(new_new_n188_), .Y(new_new_n461_));
  NO2        g0439(.A(i_3_), .B(new_new_n49_), .Y(new_new_n462_));
  NA3        g0440(.A(new_new_n356_), .B(new_new_n355_), .C(new_new_n462_), .Y(new_new_n463_));
  NA2        g0441(.A(new_new_n334_), .B(new_new_n339_), .Y(new_new_n464_));
  OAI210     g0442(.A0(new_new_n464_), .A1(new_new_n195_), .B0(new_new_n463_), .Y(new_new_n465_));
  NO3        g0443(.A(new_new_n465_), .B(new_new_n461_), .C(new_new_n459_), .Y(new_new_n466_));
  AOI210     g0444(.A0(new_new_n466_), .A1(new_new_n456_), .B0(new_new_n286_), .Y(new_new_n467_));
  NO4        g0445(.A(new_new_n467_), .B(new_new_n449_), .C(new_new_n427_), .D(new_new_n402_), .Y(new_new_n468_));
  NO2        g0446(.A(new_new_n64_), .B(i_4_), .Y(new_new_n469_));
  NO2        g0447(.A(new_new_n74_), .B(i_13_), .Y(new_new_n470_));
  NO2        g0448(.A(i_10_), .B(i_9_), .Y(new_new_n471_));
  NAi21      g0449(.An(i_12_), .B(i_8_), .Y(new_new_n472_));
  NO2        g0450(.A(new_new_n472_), .B(i_3_), .Y(new_new_n473_));
  NO2        g0451(.A(new_new_n47_), .B(i_4_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n474_), .B(new_new_n108_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n475_), .B(new_new_n211_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n327_), .B(i_0_), .Y(new_new_n477_));
  NO3        g0455(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n478_));
  NA2        g0456(.A(new_new_n281_), .B(new_new_n101_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n479_), .B(new_new_n478_), .Y(new_new_n480_));
  NA2        g0458(.A(i_8_), .B(i_9_), .Y(new_new_n481_));
  AOI210     g0459(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n482_));
  OR2        g0460(.A(new_new_n482_), .B(new_new_n481_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n299_), .B(new_new_n212_), .Y(new_new_n484_));
  OAI220     g0462(.A0(new_new_n484_), .A1(new_new_n483_), .B0(new_new_n480_), .B1(new_new_n477_), .Y(new_new_n485_));
  NA2        g0463(.A(new_new_n262_), .B(new_new_n326_), .Y(new_new_n486_));
  NO3        g0464(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n487_));
  INV        g0465(.A(new_new_n487_), .Y(new_new_n488_));
  NA3        g0466(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n489_));
  NA4        g0467(.A(new_new_n148_), .B(new_new_n119_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n490_));
  OAI220     g0468(.A0(new_new_n490_), .A1(new_new_n489_), .B0(new_new_n488_), .B1(new_new_n486_), .Y(new_new_n491_));
  NO3        g0469(.A(new_new_n491_), .B(new_new_n485_), .C(new_new_n476_), .Y(new_new_n492_));
  NA2        g0470(.A(new_new_n312_), .B(new_new_n112_), .Y(new_new_n493_));
  OR2        g0471(.A(new_new_n493_), .B(new_new_n215_), .Y(new_new_n494_));
  OA210      g0472(.A0(new_new_n374_), .A1(new_new_n105_), .B0(new_new_n314_), .Y(new_new_n495_));
  OA220      g0473(.A0(new_new_n495_), .A1(new_new_n166_), .B0(new_new_n494_), .B1(new_new_n242_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n100_), .B(i_13_), .Y(new_new_n497_));
  NA2        g0475(.A(new_new_n453_), .B(new_new_n403_), .Y(new_new_n498_));
  NO2        g0476(.A(i_2_), .B(i_13_), .Y(new_new_n499_));
  NA3        g0477(.A(new_new_n499_), .B(new_new_n165_), .C(new_new_n103_), .Y(new_new_n500_));
  OAI220     g0478(.A0(new_new_n500_), .A1(new_new_n247_), .B0(new_new_n498_), .B1(new_new_n497_), .Y(new_new_n501_));
  NO3        g0479(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n502_));
  NO2        g0480(.A(i_6_), .B(i_7_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n503_), .B(new_new_n502_), .Y(new_new_n504_));
  NO2        g0482(.A(i_11_), .B(i_1_), .Y(new_new_n505_));
  NO2        g0483(.A(new_new_n74_), .B(i_3_), .Y(new_new_n506_));
  OR2        g0484(.A(i_11_), .B(i_8_), .Y(new_new_n507_));
  NOi21      g0485(.An(i_2_), .B(i_7_), .Y(new_new_n508_));
  NAi31      g0486(.An(new_new_n507_), .B(new_new_n508_), .C(new_new_n506_), .Y(new_new_n509_));
  NO2        g0487(.A(new_new_n440_), .B(i_6_), .Y(new_new_n510_));
  NA3        g0488(.A(new_new_n510_), .B(new_new_n469_), .C(new_new_n76_), .Y(new_new_n511_));
  NO2        g0489(.A(new_new_n511_), .B(new_new_n509_), .Y(new_new_n512_));
  NO2        g0490(.A(i_3_), .B(new_new_n199_), .Y(new_new_n513_));
  NO2        g0491(.A(i_6_), .B(i_10_), .Y(new_new_n514_));
  NA4        g0492(.A(new_new_n514_), .B(new_new_n331_), .C(new_new_n513_), .D(new_new_n247_), .Y(new_new_n515_));
  NO2        g0493(.A(new_new_n515_), .B(new_new_n159_), .Y(new_new_n516_));
  NA3        g0494(.A(new_new_n256_), .B(new_new_n176_), .C(new_new_n135_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n518_));
  NO2        g0496(.A(new_new_n161_), .B(i_3_), .Y(new_new_n519_));
  NAi31      g0497(.An(new_new_n518_), .B(new_new_n519_), .C(new_new_n236_), .Y(new_new_n520_));
  NA3        g0498(.A(new_new_n416_), .B(new_new_n184_), .C(new_new_n152_), .Y(new_new_n521_));
  NA3        g0499(.A(new_new_n521_), .B(new_new_n520_), .C(new_new_n517_), .Y(new_new_n522_));
  NO4        g0500(.A(new_new_n522_), .B(new_new_n516_), .C(new_new_n512_), .D(new_new_n501_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n478_), .B(new_new_n404_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n487_), .B(new_new_n411_), .Y(new_new_n525_));
  NO2        g0503(.A(new_new_n525_), .B(new_new_n234_), .Y(new_new_n526_));
  NAi21      g0504(.An(new_new_n225_), .B(new_new_n420_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n356_), .B(new_new_n227_), .Y(new_new_n528_));
  NO2        g0506(.A(new_new_n26_), .B(i_5_), .Y(new_new_n529_));
  NO2        g0507(.A(i_0_), .B(new_new_n87_), .Y(new_new_n530_));
  NA3        g0508(.A(new_new_n530_), .B(new_new_n529_), .C(new_new_n145_), .Y(new_new_n531_));
  OR3        g0509(.A(new_new_n320_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n532_));
  OAI220     g0510(.A0(new_new_n532_), .A1(new_new_n531_), .B0(new_new_n528_), .B1(new_new_n527_), .Y(new_new_n533_));
  NA2        g0511(.A(new_new_n27_), .B(i_10_), .Y(new_new_n534_));
  NO2        g0512(.A(new_new_n534_), .B(new_new_n497_), .Y(new_new_n535_));
  NA4        g0513(.A(new_new_n324_), .B(new_new_n233_), .C(new_new_n74_), .D(new_new_n247_), .Y(new_new_n536_));
  NO2        g0514(.A(new_new_n536_), .B(new_new_n504_), .Y(new_new_n537_));
  NO4        g0515(.A(new_new_n537_), .B(new_new_n535_), .C(new_new_n533_), .D(new_new_n526_), .Y(new_new_n538_));
  NA4        g0516(.A(new_new_n538_), .B(new_new_n523_), .C(new_new_n496_), .D(new_new_n492_), .Y(new_new_n539_));
  NA3        g0517(.A(new_new_n324_), .B(new_new_n181_), .C(new_new_n179_), .Y(new_new_n540_));
  OAI210     g0518(.A0(new_new_n318_), .A1(new_new_n186_), .B0(new_new_n540_), .Y(new_new_n541_));
  AN2        g0519(.A(new_new_n303_), .B(new_new_n244_), .Y(new_new_n542_));
  NA2        g0520(.A(new_new_n542_), .B(new_new_n541_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n125_), .B(new_new_n115_), .Y(new_new_n544_));
  AO220      g0522(.A0(new_new_n544_), .A1(new_new_n478_), .B0(new_new_n441_), .B1(i_6_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n331_), .B(new_new_n168_), .Y(new_new_n546_));
  OAI210     g0524(.A0(new_new_n546_), .A1(new_new_n242_), .B0(new_new_n325_), .Y(new_new_n547_));
  AOI220     g0525(.A0(new_new_n547_), .A1(new_new_n343_), .B0(new_new_n545_), .B1(new_new_n327_), .Y(new_new_n548_));
  NA2        g0526(.A(new_new_n404_), .B(new_new_n235_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n378_), .B(new_new_n74_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n391_), .B(new_new_n387_), .Y(new_new_n551_));
  AO210      g0529(.A0(new_new_n550_), .A1(new_new_n549_), .B0(new_new_n551_), .Y(new_new_n552_));
  NO2        g0530(.A(new_new_n36_), .B(i_8_), .Y(new_new_n553_));
  AOI210     g0531(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n441_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n554_), .B(new_new_n552_), .Y(new_new_n555_));
  INV        g0533(.A(new_new_n555_), .Y(new_new_n556_));
  NA2        g0534(.A(new_new_n269_), .B(new_new_n65_), .Y(new_new_n557_));
  OAI210     g0535(.A0(i_8_), .A1(new_new_n557_), .B0(new_new_n137_), .Y(new_new_n558_));
  NO2        g0536(.A(i_7_), .B(new_new_n205_), .Y(new_new_n559_));
  OR2        g0537(.A(new_new_n188_), .B(i_4_), .Y(new_new_n560_));
  NO2        g0538(.A(new_new_n560_), .B(new_new_n87_), .Y(new_new_n561_));
  AOI220     g0539(.A0(new_new_n561_), .A1(new_new_n559_), .B0(new_new_n558_), .B1(new_new_n442_), .Y(new_new_n562_));
  NA4        g0540(.A(new_new_n562_), .B(new_new_n556_), .C(new_new_n548_), .D(new_new_n543_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n410_), .B(new_new_n312_), .Y(new_new_n564_));
  OAI210     g0542(.A0(new_new_n406_), .A1(new_new_n173_), .B0(new_new_n564_), .Y(new_new_n565_));
  NO2        g0543(.A(i_12_), .B(new_new_n199_), .Y(new_new_n566_));
  NA2        g0544(.A(new_new_n566_), .B(new_new_n235_), .Y(new_new_n567_));
  NO3        g0545(.A(new_new_n1112_), .B(new_new_n567_), .C(new_new_n493_), .Y(new_new_n568_));
  NOi31      g0546(.An(new_new_n334_), .B(new_new_n440_), .C(new_new_n38_), .Y(new_new_n569_));
  OAI210     g0547(.A0(new_new_n569_), .A1(new_new_n568_), .B0(new_new_n565_), .Y(new_new_n570_));
  NO2        g0548(.A(i_8_), .B(i_7_), .Y(new_new_n571_));
  OAI210     g0549(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n572_));
  NA2        g0550(.A(new_new_n572_), .B(new_new_n233_), .Y(new_new_n573_));
  AOI220     g0551(.A0(new_new_n344_), .A1(new_new_n40_), .B0(new_new_n245_), .B1(new_new_n214_), .Y(new_new_n574_));
  OAI220     g0552(.A0(new_new_n574_), .A1(new_new_n560_), .B0(new_new_n573_), .B1(new_new_n253_), .Y(new_new_n575_));
  NA2        g0553(.A(new_new_n45_), .B(i_10_), .Y(new_new_n576_));
  NO2        g0554(.A(new_new_n576_), .B(i_6_), .Y(new_new_n577_));
  NA3        g0555(.A(new_new_n577_), .B(new_new_n575_), .C(new_new_n571_), .Y(new_new_n578_));
  AOI220     g0556(.A0(new_new_n453_), .A1(new_new_n344_), .B0(new_new_n258_), .B1(new_new_n255_), .Y(new_new_n579_));
  OAI220     g0557(.A0(new_new_n579_), .A1(new_new_n277_), .B0(new_new_n497_), .B1(new_new_n136_), .Y(new_new_n580_));
  NA2        g0558(.A(new_new_n580_), .B(new_new_n280_), .Y(new_new_n581_));
  NOi31      g0559(.An(new_new_n307_), .B(new_new_n318_), .C(new_new_n186_), .Y(new_new_n582_));
  NA3        g0560(.A(new_new_n324_), .B(new_new_n179_), .C(new_new_n100_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n231_), .B(new_new_n45_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n161_), .B(i_5_), .Y(new_new_n585_));
  NA3        g0563(.A(new_new_n585_), .B(new_new_n428_), .C(new_new_n337_), .Y(new_new_n586_));
  OAI210     g0564(.A0(new_new_n586_), .A1(new_new_n584_), .B0(new_new_n583_), .Y(new_new_n587_));
  OAI210     g0565(.A0(new_new_n587_), .A1(new_new_n582_), .B0(new_new_n487_), .Y(new_new_n588_));
  NA4        g0566(.A(new_new_n588_), .B(new_new_n581_), .C(new_new_n578_), .D(new_new_n570_), .Y(new_new_n589_));
  NA3        g0567(.A(new_new_n227_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n590_));
  NA2        g0568(.A(new_new_n299_), .B(new_new_n85_), .Y(new_new_n591_));
  AOI210     g0569(.A0(new_new_n590_), .A1(new_new_n369_), .B0(new_new_n591_), .Y(new_new_n592_));
  NA2        g0570(.A(new_new_n313_), .B(new_new_n303_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n593_), .B(new_new_n178_), .Y(new_new_n594_));
  NA2        g0572(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n595_));
  NA2        g0573(.A(new_new_n471_), .B(new_new_n231_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n595_), .B(new_new_n596_), .Y(new_new_n597_));
  AOI210     g0575(.A0(i_6_), .A1(new_new_n47_), .B0(new_new_n388_), .Y(new_new_n598_));
  NA2        g0576(.A(i_0_), .B(new_new_n49_), .Y(new_new_n599_));
  NA3        g0577(.A(new_new_n566_), .B(new_new_n290_), .C(new_new_n599_), .Y(new_new_n600_));
  NO2        g0578(.A(new_new_n598_), .B(new_new_n600_), .Y(new_new_n601_));
  NO4        g0579(.A(new_new_n601_), .B(new_new_n597_), .C(new_new_n594_), .D(new_new_n592_), .Y(new_new_n602_));
  NO4        g0580(.A(new_new_n263_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n603_));
  NO3        g0581(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n243_), .B(new_new_n36_), .Y(new_new_n605_));
  AN2        g0583(.A(new_new_n605_), .B(new_new_n604_), .Y(new_new_n606_));
  OA210      g0584(.A0(new_new_n606_), .A1(new_new_n603_), .B0(new_new_n378_), .Y(new_new_n607_));
  NO2        g0585(.A(new_new_n440_), .B(i_1_), .Y(new_new_n608_));
  NOi31      g0586(.An(new_new_n608_), .B(new_new_n479_), .C(new_new_n74_), .Y(new_new_n609_));
  AN4        g0587(.A(new_new_n609_), .B(new_new_n437_), .C(new_new_n529_), .D(i_2_), .Y(new_new_n610_));
  NO2        g0588(.A(new_new_n451_), .B(new_new_n182_), .Y(new_new_n611_));
  NO3        g0589(.A(new_new_n611_), .B(new_new_n610_), .C(new_new_n607_), .Y(new_new_n612_));
  NOi21      g0590(.An(i_10_), .B(i_6_), .Y(new_new_n613_));
  NO2        g0591(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n614_));
  AOI220     g0592(.A0(new_new_n299_), .A1(new_new_n614_), .B0(new_new_n290_), .B1(new_new_n613_), .Y(new_new_n615_));
  NO2        g0593(.A(new_new_n615_), .B(new_new_n477_), .Y(new_new_n616_));
  NO2        g0594(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n617_));
  NA2        g0595(.A(new_new_n334_), .B(new_new_n168_), .Y(new_new_n618_));
  AOI220     g0596(.A0(new_new_n618_), .A1(new_new_n460_), .B0(new_new_n189_), .B1(new_new_n187_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n204_), .B(new_new_n37_), .Y(new_new_n620_));
  NOi31      g0598(.An(new_new_n149_), .B(new_new_n620_), .C(new_new_n351_), .Y(new_new_n621_));
  NO3        g0599(.A(new_new_n621_), .B(new_new_n619_), .C(new_new_n616_), .Y(new_new_n622_));
  NO2        g0600(.A(new_new_n550_), .B(new_new_n399_), .Y(new_new_n623_));
  INV        g0601(.A(new_new_n337_), .Y(new_new_n624_));
  NO2        g0602(.A(i_12_), .B(new_new_n87_), .Y(new_new_n625_));
  NA3        g0603(.A(new_new_n625_), .B(new_new_n290_), .C(new_new_n599_), .Y(new_new_n626_));
  NA3        g0604(.A(new_new_n407_), .B(new_new_n299_), .C(new_new_n227_), .Y(new_new_n627_));
  AOI210     g0605(.A0(new_new_n627_), .A1(new_new_n626_), .B0(new_new_n624_), .Y(new_new_n628_));
  NA2        g0606(.A(new_new_n179_), .B(i_0_), .Y(new_new_n629_));
  NO3        g0607(.A(new_new_n629_), .B(new_new_n362_), .C(new_new_n318_), .Y(new_new_n630_));
  OR2        g0608(.A(i_2_), .B(i_5_), .Y(new_new_n631_));
  OR2        g0609(.A(new_new_n631_), .B(new_new_n432_), .Y(new_new_n632_));
  NO2        g0610(.A(new_new_n632_), .B(new_new_n527_), .Y(new_new_n633_));
  NO4        g0611(.A(new_new_n633_), .B(new_new_n630_), .C(new_new_n628_), .D(new_new_n623_), .Y(new_new_n634_));
  NA4        g0612(.A(new_new_n634_), .B(new_new_n622_), .C(new_new_n612_), .D(new_new_n602_), .Y(new_new_n635_));
  NO4        g0613(.A(new_new_n635_), .B(new_new_n589_), .C(new_new_n563_), .D(new_new_n539_), .Y(new_new_n636_));
  NA4        g0614(.A(new_new_n636_), .B(new_new_n468_), .C(new_new_n377_), .D(new_new_n330_), .Y(men7));
  NO2        g0615(.A(new_new_n96_), .B(new_new_n55_), .Y(new_new_n638_));
  NO2        g0616(.A(new_new_n112_), .B(new_new_n93_), .Y(new_new_n639_));
  NA2        g0617(.A(new_new_n405_), .B(new_new_n639_), .Y(new_new_n640_));
  NA2        g0618(.A(new_new_n514_), .B(new_new_n85_), .Y(new_new_n641_));
  NA2        g0619(.A(i_11_), .B(new_new_n199_), .Y(new_new_n642_));
  INV        g0620(.A(new_new_n640_), .Y(new_new_n643_));
  NA3        g0621(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n644_));
  NO2        g0622(.A(new_new_n247_), .B(i_4_), .Y(new_new_n645_));
  NA2        g0623(.A(new_new_n645_), .B(i_8_), .Y(new_new_n646_));
  NO2        g0624(.A(new_new_n109_), .B(new_new_n644_), .Y(new_new_n647_));
  NA2        g0625(.A(i_2_), .B(new_new_n87_), .Y(new_new_n648_));
  OAI210     g0626(.A0(new_new_n90_), .A1(new_new_n209_), .B0(new_new_n210_), .Y(new_new_n649_));
  NO2        g0627(.A(i_7_), .B(new_new_n37_), .Y(new_new_n650_));
  NA2        g0628(.A(i_4_), .B(i_8_), .Y(new_new_n651_));
  AOI210     g0629(.A0(new_new_n651_), .A1(new_new_n324_), .B0(new_new_n650_), .Y(new_new_n652_));
  OAI220     g0630(.A0(new_new_n652_), .A1(new_new_n648_), .B0(new_new_n649_), .B1(i_13_), .Y(new_new_n653_));
  NO4        g0631(.A(new_new_n653_), .B(new_new_n647_), .C(new_new_n643_), .D(new_new_n638_), .Y(new_new_n654_));
  AOI210     g0632(.A0(new_new_n131_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n655_));
  AOI210     g0633(.A0(new_new_n655_), .A1(new_new_n247_), .B0(new_new_n165_), .Y(new_new_n656_));
  OR2        g0634(.A(i_6_), .B(i_10_), .Y(new_new_n657_));
  NO2        g0635(.A(new_new_n657_), .B(new_new_n23_), .Y(new_new_n658_));
  OR3        g0636(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n659_));
  NO3        g0637(.A(new_new_n659_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n660_));
  INV        g0638(.A(new_new_n206_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n660_), .B(new_new_n658_), .Y(new_new_n662_));
  OA220      g0640(.A0(new_new_n662_), .A1(new_new_n624_), .B0(new_new_n656_), .B1(new_new_n282_), .Y(new_new_n663_));
  AOI210     g0641(.A0(new_new_n663_), .A1(new_new_n654_), .B0(new_new_n64_), .Y(new_new_n664_));
  NOi21      g0642(.An(i_11_), .B(i_7_), .Y(new_new_n665_));
  AO210      g0643(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n666_), .B(new_new_n665_), .Y(new_new_n667_));
  NA2        g0645(.A(new_new_n667_), .B(new_new_n214_), .Y(new_new_n668_));
  NA3        g0646(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n669_));
  NAi31      g0647(.An(new_new_n669_), .B(new_new_n224_), .C(i_11_), .Y(new_new_n670_));
  AOI210     g0648(.A0(new_new_n670_), .A1(new_new_n668_), .B0(new_new_n64_), .Y(new_new_n671_));
  NA2        g0649(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n672_));
  AO210      g0650(.A0(new_new_n672_), .A1(new_new_n399_), .B0(new_new_n41_), .Y(new_new_n673_));
  NO3        g0651(.A(new_new_n271_), .B(new_new_n216_), .C(new_new_n642_), .Y(new_new_n674_));
  OAI210     g0652(.A0(new_new_n674_), .A1(new_new_n236_), .B0(new_new_n64_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n433_), .B(new_new_n31_), .Y(new_new_n676_));
  OR2        g0654(.A(new_new_n216_), .B(new_new_n112_), .Y(new_new_n677_));
  NA2        g0655(.A(new_new_n677_), .B(new_new_n676_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n64_), .B(i_9_), .Y(new_new_n679_));
  NO2        g0657(.A(new_new_n679_), .B(i_4_), .Y(new_new_n680_));
  NA2        g0658(.A(new_new_n680_), .B(new_new_n678_), .Y(new_new_n681_));
  NO2        g0659(.A(i_1_), .B(i_12_), .Y(new_new_n682_));
  NA3        g0660(.A(new_new_n682_), .B(new_new_n113_), .C(new_new_n24_), .Y(new_new_n683_));
  NA4        g0661(.A(new_new_n683_), .B(new_new_n681_), .C(new_new_n675_), .D(new_new_n673_), .Y(new_new_n684_));
  OAI210     g0662(.A0(new_new_n684_), .A1(new_new_n671_), .B0(i_6_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n247_), .B(new_new_n87_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n686_), .B(i_11_), .Y(new_new_n687_));
  INV        g0665(.A(new_new_n480_), .Y(new_new_n688_));
  NO4        g0666(.A(new_new_n224_), .B(new_new_n131_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n689_));
  NA2        g0667(.A(new_new_n689_), .B(new_new_n679_), .Y(new_new_n690_));
  NA2        g0668(.A(new_new_n247_), .B(i_6_), .Y(new_new_n691_));
  NO3        g0669(.A(new_new_n657_), .B(new_new_n243_), .C(new_new_n23_), .Y(new_new_n692_));
  AOI210     g0670(.A0(i_1_), .A1(new_new_n272_), .B0(new_new_n692_), .Y(new_new_n693_));
  OAI210     g0671(.A0(new_new_n693_), .A1(new_new_n45_), .B0(new_new_n690_), .Y(new_new_n694_));
  NA3        g0672(.A(new_new_n571_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n695_));
  NA2        g0673(.A(new_new_n141_), .B(i_9_), .Y(new_new_n696_));
  NA3        g0674(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n47_), .B(i_1_), .Y(new_new_n698_));
  NO2        g0676(.A(new_new_n696_), .B(new_new_n1111_), .Y(new_new_n699_));
  NA3        g0677(.A(new_new_n679_), .B(new_new_n337_), .C(i_6_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n700_), .B(new_new_n23_), .Y(new_new_n701_));
  AOI210     g0679(.A0(new_new_n505_), .A1(new_new_n444_), .B0(new_new_n252_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n702_), .B(new_new_n648_), .Y(new_new_n703_));
  NO2        g0681(.A(i_11_), .B(new_new_n37_), .Y(new_new_n704_));
  NA2        g0682(.A(new_new_n704_), .B(new_new_n24_), .Y(new_new_n705_));
  OR3        g0683(.A(new_new_n703_), .B(new_new_n701_), .C(new_new_n699_), .Y(new_new_n706_));
  NO3        g0684(.A(new_new_n706_), .B(new_new_n694_), .C(new_new_n688_), .Y(new_new_n707_));
  NO2        g0685(.A(new_new_n247_), .B(new_new_n105_), .Y(new_new_n708_));
  NO2        g0686(.A(new_new_n708_), .B(new_new_n665_), .Y(new_new_n709_));
  NA2        g0687(.A(new_new_n709_), .B(i_1_), .Y(new_new_n710_));
  NO2        g0688(.A(new_new_n710_), .B(new_new_n659_), .Y(new_new_n711_));
  NO2        g0689(.A(new_new_n439_), .B(new_new_n87_), .Y(new_new_n712_));
  NA2        g0690(.A(new_new_n711_), .B(new_new_n47_), .Y(new_new_n713_));
  NO2        g0691(.A(new_new_n243_), .B(new_new_n45_), .Y(new_new_n714_));
  NO3        g0692(.A(new_new_n714_), .B(new_new_n327_), .C(new_new_n248_), .Y(new_new_n715_));
  NO2        g0693(.A(new_new_n120_), .B(new_new_n37_), .Y(new_new_n716_));
  NO2        g0694(.A(new_new_n716_), .B(i_6_), .Y(new_new_n717_));
  NO2        g0695(.A(new_new_n87_), .B(i_9_), .Y(new_new_n718_));
  NO2        g0696(.A(new_new_n718_), .B(new_new_n64_), .Y(new_new_n719_));
  NO2        g0697(.A(new_new_n719_), .B(new_new_n682_), .Y(new_new_n720_));
  NO4        g0698(.A(new_new_n720_), .B(new_new_n717_), .C(new_new_n715_), .D(i_4_), .Y(new_new_n721_));
  NA2        g0699(.A(i_1_), .B(i_3_), .Y(new_new_n722_));
  INV        g0700(.A(new_new_n721_), .Y(new_new_n723_));
  NA4        g0701(.A(new_new_n723_), .B(new_new_n713_), .C(new_new_n707_), .D(new_new_n685_), .Y(new_new_n724_));
  NO3        g0702(.A(new_new_n507_), .B(i_3_), .C(i_7_), .Y(new_new_n725_));
  NOi21      g0703(.An(new_new_n725_), .B(i_10_), .Y(new_new_n726_));
  OA210      g0704(.A0(new_new_n726_), .A1(new_new_n256_), .B0(new_new_n87_), .Y(new_new_n727_));
  NO3        g0705(.A(new_new_n508_), .B(new_new_n651_), .C(new_new_n87_), .Y(new_new_n728_));
  NA2        g0706(.A(new_new_n728_), .B(new_new_n25_), .Y(new_new_n729_));
  NA3        g0707(.A(new_new_n165_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n730_), .B(new_new_n729_), .Y(new_new_n731_));
  OAI210     g0709(.A0(new_new_n731_), .A1(new_new_n727_), .B0(i_1_), .Y(new_new_n732_));
  AOI210     g0710(.A0(new_new_n281_), .A1(new_new_n101_), .B0(i_1_), .Y(new_new_n733_));
  NO2        g0711(.A(new_new_n389_), .B(i_2_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n734_), .B(new_new_n733_), .Y(new_new_n735_));
  OAI210     g0713(.A0(new_new_n700_), .A1(new_new_n472_), .B0(new_new_n735_), .Y(new_new_n736_));
  INV        g0714(.A(new_new_n736_), .Y(new_new_n737_));
  AOI210     g0715(.A0(new_new_n737_), .A1(new_new_n732_), .B0(i_13_), .Y(new_new_n738_));
  OR2        g0716(.A(i_11_), .B(i_7_), .Y(new_new_n739_));
  NA3        g0717(.A(new_new_n739_), .B(new_new_n110_), .C(new_new_n141_), .Y(new_new_n740_));
  AOI220     g0718(.A0(new_new_n499_), .A1(new_new_n165_), .B0(new_new_n474_), .B1(new_new_n141_), .Y(new_new_n741_));
  OAI210     g0719(.A0(new_new_n741_), .A1(new_new_n45_), .B0(new_new_n740_), .Y(new_new_n742_));
  AOI210     g0720(.A0(new_new_n697_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n743_));
  NO2        g0721(.A(new_new_n508_), .B(new_new_n24_), .Y(new_new_n744_));
  AOI220     g0722(.A0(new_new_n744_), .A1(new_new_n712_), .B0(new_new_n256_), .B1(new_new_n134_), .Y(new_new_n745_));
  OAI220     g0723(.A0(new_new_n745_), .A1(new_new_n41_), .B0(new_new_n1110_), .B1(new_new_n96_), .Y(new_new_n746_));
  AOI210     g0724(.A0(new_new_n742_), .A1(new_new_n353_), .B0(new_new_n746_), .Y(new_new_n747_));
  NA2        g0725(.A(new_new_n407_), .B(new_new_n698_), .Y(new_new_n748_));
  NO2        g0726(.A(new_new_n748_), .B(new_new_n253_), .Y(new_new_n749_));
  AOI210     g0727(.A0(new_new_n472_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n750_));
  NOi31      g0728(.An(new_new_n750_), .B(new_new_n641_), .C(new_new_n45_), .Y(new_new_n751_));
  NA2        g0729(.A(new_new_n130_), .B(i_13_), .Y(new_new_n752_));
  NO2        g0730(.A(new_new_n697_), .B(new_new_n118_), .Y(new_new_n753_));
  INV        g0731(.A(new_new_n753_), .Y(new_new_n754_));
  OAI220     g0732(.A0(new_new_n754_), .A1(new_new_n72_), .B0(new_new_n752_), .B1(new_new_n733_), .Y(new_new_n755_));
  NO3        g0733(.A(new_new_n72_), .B(new_new_n32_), .C(new_new_n105_), .Y(new_new_n756_));
  NA2        g0734(.A(new_new_n26_), .B(new_new_n199_), .Y(new_new_n757_));
  NA2        g0735(.A(new_new_n757_), .B(i_7_), .Y(new_new_n758_));
  INV        g0736(.A(new_new_n756_), .Y(new_new_n759_));
  AOI220     g0737(.A0(new_new_n407_), .A1(new_new_n698_), .B0(new_new_n95_), .B1(new_new_n106_), .Y(new_new_n760_));
  OAI220     g0738(.A0(new_new_n760_), .A1(new_new_n646_), .B0(new_new_n759_), .B1(new_new_n661_), .Y(new_new_n761_));
  NO4        g0739(.A(new_new_n761_), .B(new_new_n755_), .C(new_new_n751_), .D(new_new_n749_), .Y(new_new_n762_));
  OR2        g0740(.A(i_11_), .B(i_6_), .Y(new_new_n763_));
  NA3        g0741(.A(new_new_n645_), .B(new_new_n757_), .C(i_7_), .Y(new_new_n764_));
  AOI210     g0742(.A0(new_new_n764_), .A1(new_new_n754_), .B0(new_new_n763_), .Y(new_new_n765_));
  NA3        g0743(.A(new_new_n433_), .B(new_new_n650_), .C(new_new_n101_), .Y(new_new_n766_));
  NA2        g0744(.A(new_new_n687_), .B(i_13_), .Y(new_new_n767_));
  NA2        g0745(.A(new_new_n106_), .B(new_new_n757_), .Y(new_new_n768_));
  NAi21      g0746(.An(i_11_), .B(i_12_), .Y(new_new_n769_));
  NOi41      g0747(.An(new_new_n114_), .B(new_new_n769_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n770_));
  NA2        g0748(.A(new_new_n770_), .B(new_new_n768_), .Y(new_new_n771_));
  NA3        g0749(.A(new_new_n771_), .B(new_new_n767_), .C(new_new_n766_), .Y(new_new_n772_));
  OAI210     g0750(.A0(new_new_n772_), .A1(new_new_n765_), .B0(new_new_n64_), .Y(new_new_n773_));
  NO2        g0751(.A(i_2_), .B(i_12_), .Y(new_new_n774_));
  NA2        g0752(.A(new_new_n388_), .B(new_new_n774_), .Y(new_new_n775_));
  NA2        g0753(.A(i_8_), .B(new_new_n25_), .Y(new_new_n776_));
  NO3        g0754(.A(new_new_n776_), .B(new_new_n405_), .C(new_new_n645_), .Y(new_new_n777_));
  OAI210     g0755(.A0(new_new_n777_), .A1(new_new_n390_), .B0(new_new_n388_), .Y(new_new_n778_));
  NO2        g0756(.A(new_new_n131_), .B(i_2_), .Y(new_new_n779_));
  NA2        g0757(.A(new_new_n779_), .B(new_new_n682_), .Y(new_new_n780_));
  NA3        g0758(.A(new_new_n780_), .B(new_new_n778_), .C(new_new_n775_), .Y(new_new_n781_));
  NA3        g0759(.A(new_new_n781_), .B(new_new_n46_), .C(new_new_n235_), .Y(new_new_n782_));
  NA4        g0760(.A(new_new_n782_), .B(new_new_n773_), .C(new_new_n762_), .D(new_new_n747_), .Y(new_new_n783_));
  OR4        g0761(.A(new_new_n783_), .B(new_new_n738_), .C(new_new_n724_), .D(new_new_n664_), .Y(men5));
  AOI210     g0762(.A0(new_new_n709_), .A1(new_new_n284_), .B0(new_new_n442_), .Y(new_new_n785_));
  AN2        g0763(.A(new_new_n24_), .B(i_10_), .Y(new_new_n786_));
  NA3        g0764(.A(new_new_n786_), .B(new_new_n774_), .C(new_new_n112_), .Y(new_new_n787_));
  NO2        g0765(.A(new_new_n646_), .B(i_11_), .Y(new_new_n788_));
  NA2        g0766(.A(new_new_n90_), .B(new_new_n788_), .Y(new_new_n789_));
  NA3        g0767(.A(new_new_n789_), .B(new_new_n787_), .C(new_new_n785_), .Y(new_new_n790_));
  NO3        g0768(.A(i_11_), .B(new_new_n247_), .C(i_13_), .Y(new_new_n791_));
  NO2        g0769(.A(new_new_n127_), .B(new_new_n23_), .Y(new_new_n792_));
  NA2        g0770(.A(i_12_), .B(i_8_), .Y(new_new_n793_));
  OAI210     g0771(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n793_), .Y(new_new_n794_));
  INV        g0772(.A(new_new_n471_), .Y(new_new_n795_));
  AOI220     g0773(.A0(new_new_n337_), .A1(new_new_n617_), .B0(new_new_n794_), .B1(new_new_n792_), .Y(new_new_n796_));
  INV        g0774(.A(new_new_n796_), .Y(new_new_n797_));
  NO2        g0775(.A(new_new_n797_), .B(new_new_n790_), .Y(new_new_n798_));
  INV        g0776(.A(new_new_n176_), .Y(new_new_n799_));
  INV        g0777(.A(new_new_n256_), .Y(new_new_n800_));
  OAI210     g0778(.A0(new_new_n734_), .A1(new_new_n473_), .B0(new_new_n114_), .Y(new_new_n801_));
  AOI210     g0779(.A0(new_new_n801_), .A1(new_new_n800_), .B0(new_new_n799_), .Y(new_new_n802_));
  NO2        g0780(.A(new_new_n481_), .B(new_new_n26_), .Y(new_new_n803_));
  NO2        g0781(.A(new_new_n803_), .B(new_new_n444_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n804_), .B(i_2_), .Y(new_new_n805_));
  INV        g0783(.A(new_new_n805_), .Y(new_new_n806_));
  AOI210     g0784(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n440_), .Y(new_new_n807_));
  AOI210     g0785(.A0(new_new_n807_), .A1(new_new_n806_), .B0(new_new_n802_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n196_), .B(new_new_n128_), .Y(new_new_n809_));
  OAI210     g0787(.A0(new_new_n809_), .A1(new_new_n792_), .B0(i_2_), .Y(new_new_n810_));
  INV        g0788(.A(new_new_n177_), .Y(new_new_n811_));
  NO3        g0789(.A(new_new_n666_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n812_));
  AOI210     g0790(.A0(new_new_n811_), .A1(new_new_n90_), .B0(new_new_n812_), .Y(new_new_n813_));
  AOI210     g0791(.A0(new_new_n813_), .A1(new_new_n810_), .B0(new_new_n199_), .Y(new_new_n814_));
  OA210      g0792(.A0(new_new_n667_), .A1(new_new_n129_), .B0(i_13_), .Y(new_new_n815_));
  NA2        g0793(.A(new_new_n206_), .B(new_new_n209_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n155_), .B(new_new_n642_), .Y(new_new_n817_));
  AOI210     g0795(.A0(new_new_n817_), .A1(new_new_n816_), .B0(new_new_n393_), .Y(new_new_n818_));
  AOI210     g0796(.A0(new_new_n216_), .A1(new_new_n151_), .B0(new_new_n553_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n819_), .B(new_new_n444_), .Y(new_new_n820_));
  NO2        g0798(.A(new_new_n106_), .B(new_new_n45_), .Y(new_new_n821_));
  INV        g0799(.A(new_new_n319_), .Y(new_new_n822_));
  NA4        g0800(.A(new_new_n822_), .B(new_new_n324_), .C(new_new_n127_), .D(new_new_n43_), .Y(new_new_n823_));
  OAI210     g0801(.A0(new_new_n823_), .A1(new_new_n821_), .B0(new_new_n820_), .Y(new_new_n824_));
  NO4        g0802(.A(new_new_n824_), .B(new_new_n818_), .C(new_new_n815_), .D(new_new_n814_), .Y(new_new_n825_));
  NA2        g0803(.A(new_new_n617_), .B(new_new_n28_), .Y(new_new_n826_));
  NA2        g0804(.A(new_new_n791_), .B(new_new_n291_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n827_), .B(new_new_n826_), .Y(new_new_n828_));
  NO2        g0806(.A(new_new_n63_), .B(i_12_), .Y(new_new_n829_));
  NO2        g0807(.A(new_new_n829_), .B(new_new_n129_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n830_), .B(new_new_n642_), .Y(new_new_n831_));
  AOI220     g0809(.A0(new_new_n831_), .A1(new_new_n36_), .B0(new_new_n828_), .B1(new_new_n47_), .Y(new_new_n832_));
  NA4        g0810(.A(new_new_n832_), .B(new_new_n825_), .C(new_new_n808_), .D(new_new_n798_), .Y(men6));
  NO3        g0811(.A(new_new_n267_), .B(new_new_n326_), .C(i_1_), .Y(new_new_n834_));
  NO2        g0812(.A(new_new_n191_), .B(new_new_n142_), .Y(new_new_n835_));
  OAI210     g0813(.A0(new_new_n835_), .A1(new_new_n834_), .B0(new_new_n779_), .Y(new_new_n836_));
  NA4        g0814(.A(new_new_n411_), .B(new_new_n513_), .C(new_new_n72_), .D(new_new_n105_), .Y(new_new_n837_));
  INV        g0815(.A(new_new_n837_), .Y(new_new_n838_));
  NO2        g0816(.A(new_new_n230_), .B(new_new_n518_), .Y(new_new_n839_));
  NO2        g0817(.A(new_new_n838_), .B(new_new_n349_), .Y(new_new_n840_));
  AO210      g0818(.A0(new_new_n840_), .A1(new_new_n836_), .B0(i_12_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n625_), .B(new_new_n64_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n726_), .B(new_new_n72_), .Y(new_new_n843_));
  BUFFER     g0821(.A(new_new_n672_), .Y(new_new_n844_));
  NA3        g0822(.A(new_new_n844_), .B(new_new_n843_), .C(new_new_n842_), .Y(new_new_n845_));
  NA2        g0823(.A(new_new_n845_), .B(new_new_n74_), .Y(new_new_n846_));
  INV        g0824(.A(new_new_n348_), .Y(new_new_n847_));
  NA2        g0825(.A(new_new_n76_), .B(new_new_n134_), .Y(new_new_n848_));
  INV        g0826(.A(new_new_n127_), .Y(new_new_n849_));
  NA2        g0827(.A(new_new_n849_), .B(new_new_n47_), .Y(new_new_n850_));
  AOI210     g0828(.A0(new_new_n850_), .A1(new_new_n848_), .B0(new_new_n847_), .Y(new_new_n851_));
  NO3        g0829(.A(new_new_n263_), .B(new_new_n135_), .C(i_9_), .Y(new_new_n852_));
  NA2        g0830(.A(new_new_n852_), .B(new_new_n829_), .Y(new_new_n853_));
  AOI210     g0831(.A0(new_new_n853_), .A1(new_new_n551_), .B0(new_new_n191_), .Y(new_new_n854_));
  NO2        g0832(.A(new_new_n32_), .B(i_11_), .Y(new_new_n855_));
  NA3        g0833(.A(new_new_n855_), .B(new_new_n503_), .C(new_new_n411_), .Y(new_new_n856_));
  NAi32      g0834(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n857_));
  AOI210     g0835(.A0(new_new_n763_), .A1(new_new_n88_), .B0(new_new_n857_), .Y(new_new_n858_));
  OAI210     g0836(.A0(new_new_n725_), .A1(new_new_n605_), .B0(new_new_n604_), .Y(new_new_n859_));
  NAi31      g0837(.An(new_new_n858_), .B(new_new_n859_), .C(new_new_n856_), .Y(new_new_n860_));
  OR3        g0838(.A(new_new_n860_), .B(new_new_n854_), .C(new_new_n851_), .Y(new_new_n861_));
  NO2        g0839(.A(new_new_n739_), .B(i_2_), .Y(new_new_n862_));
  NA2        g0840(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n863_));
  OAI210     g0841(.A0(new_new_n863_), .A1(new_new_n432_), .B0(new_new_n383_), .Y(new_new_n864_));
  NA2        g0842(.A(new_new_n864_), .B(new_new_n862_), .Y(new_new_n865_));
  AO220      g0843(.A0(new_new_n382_), .A1(new_new_n373_), .B0(new_new_n419_), .B1(new_new_n642_), .Y(new_new_n866_));
  NA3        g0844(.A(new_new_n866_), .B(new_new_n268_), .C(i_7_), .Y(new_new_n867_));
  OR2        g0845(.A(new_new_n667_), .B(new_new_n473_), .Y(new_new_n868_));
  NA3        g0846(.A(new_new_n868_), .B(new_new_n150_), .C(new_new_n70_), .Y(new_new_n869_));
  AO210      g0847(.A0(new_new_n525_), .A1(new_new_n795_), .B0(new_new_n36_), .Y(new_new_n870_));
  NA4        g0848(.A(new_new_n870_), .B(new_new_n869_), .C(new_new_n867_), .D(new_new_n865_), .Y(new_new_n871_));
  OAI210     g0849(.A0(new_new_n686_), .A1(i_11_), .B0(new_new_n88_), .Y(new_new_n872_));
  AOI220     g0850(.A0(new_new_n872_), .A1(new_new_n604_), .B0(new_new_n839_), .B1(new_new_n758_), .Y(new_new_n873_));
  NA3        g0851(.A(new_new_n393_), .B(new_new_n249_), .C(new_new_n150_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n419_), .B(new_new_n71_), .Y(new_new_n875_));
  NA4        g0853(.A(new_new_n875_), .B(new_new_n874_), .C(new_new_n873_), .D(new_new_n649_), .Y(new_new_n876_));
  AO210      g0854(.A0(new_new_n553_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n877_));
  NA3        g0855(.A(new_new_n877_), .B(new_new_n514_), .C(new_new_n227_), .Y(new_new_n878_));
  AOI210     g0856(.A0(new_new_n473_), .A1(new_new_n471_), .B0(new_new_n603_), .Y(new_new_n879_));
  NO2        g0857(.A(new_new_n657_), .B(new_new_n106_), .Y(new_new_n880_));
  OAI210     g0858(.A0(new_new_n880_), .A1(new_new_n115_), .B0(new_new_n430_), .Y(new_new_n881_));
  NA2        g0859(.A(new_new_n255_), .B(new_new_n47_), .Y(new_new_n882_));
  INV        g0860(.A(new_new_n632_), .Y(new_new_n883_));
  NA3        g0861(.A(new_new_n883_), .B(new_new_n348_), .C(i_7_), .Y(new_new_n884_));
  NA4        g0862(.A(new_new_n884_), .B(new_new_n881_), .C(new_new_n879_), .D(new_new_n878_), .Y(new_new_n885_));
  NO4        g0863(.A(new_new_n885_), .B(new_new_n876_), .C(new_new_n871_), .D(new_new_n861_), .Y(new_new_n886_));
  NA4        g0864(.A(new_new_n886_), .B(new_new_n846_), .C(new_new_n841_), .D(new_new_n401_), .Y(men3));
  NA2        g0865(.A(i_6_), .B(i_7_), .Y(new_new_n888_));
  NO2        g0866(.A(new_new_n888_), .B(i_0_), .Y(new_new_n889_));
  NO2        g0867(.A(i_11_), .B(new_new_n247_), .Y(new_new_n890_));
  OAI210     g0868(.A0(new_new_n889_), .A1(new_new_n307_), .B0(new_new_n890_), .Y(new_new_n891_));
  NO2        g0869(.A(new_new_n891_), .B(new_new_n199_), .Y(new_new_n892_));
  NO3        g0870(.A(new_new_n477_), .B(new_new_n93_), .C(new_new_n45_), .Y(new_new_n893_));
  OA210      g0871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n179_), .Y(new_new_n894_));
  NA3        g0872(.A(new_new_n874_), .B(new_new_n649_), .C(new_new_n392_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n895_), .B(new_new_n40_), .Y(new_new_n896_));
  NOi21      g0874(.An(new_new_n100_), .B(new_new_n804_), .Y(new_new_n897_));
  NO3        g0875(.A(new_new_n677_), .B(new_new_n481_), .C(new_new_n134_), .Y(new_new_n898_));
  AN2        g0876(.A(new_new_n479_), .B(new_new_n56_), .Y(new_new_n899_));
  NO3        g0877(.A(new_new_n899_), .B(new_new_n898_), .C(new_new_n897_), .Y(new_new_n900_));
  AOI210     g0878(.A0(new_new_n900_), .A1(new_new_n896_), .B0(new_new_n49_), .Y(new_new_n901_));
  NO4        g0879(.A(new_new_n397_), .B(new_new_n404_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n902_));
  NA2        g0880(.A(new_new_n191_), .B(new_new_n613_), .Y(new_new_n903_));
  NOi21      g0881(.An(new_new_n903_), .B(new_new_n902_), .Y(new_new_n904_));
  NA2        g0882(.A(new_new_n750_), .B(new_new_n718_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n354_), .B(new_new_n462_), .Y(new_new_n906_));
  OAI220     g0884(.A0(new_new_n906_), .A1(new_new_n905_), .B0(new_new_n904_), .B1(new_new_n64_), .Y(new_new_n907_));
  NOi21      g0885(.An(i_5_), .B(i_9_), .Y(new_new_n908_));
  NA2        g0886(.A(new_new_n908_), .B(new_new_n470_), .Y(new_new_n909_));
  AOI210     g0887(.A0(new_new_n281_), .A1(new_new_n505_), .B0(new_new_n728_), .Y(new_new_n910_));
  NO3        g0888(.A(new_new_n436_), .B(new_new_n281_), .C(new_new_n74_), .Y(new_new_n911_));
  NO2        g0889(.A(new_new_n180_), .B(new_new_n151_), .Y(new_new_n912_));
  AOI210     g0890(.A0(new_new_n912_), .A1(new_new_n255_), .B0(new_new_n911_), .Y(new_new_n913_));
  OAI220     g0891(.A0(new_new_n913_), .A1(new_new_n186_), .B0(new_new_n910_), .B1(new_new_n909_), .Y(new_new_n914_));
  NO4        g0892(.A(new_new_n914_), .B(new_new_n907_), .C(new_new_n901_), .D(new_new_n894_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n191_), .B(new_new_n24_), .Y(new_new_n916_));
  NO2        g0894(.A(new_new_n716_), .B(new_new_n639_), .Y(new_new_n917_));
  NO2        g0895(.A(new_new_n917_), .B(new_new_n916_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n331_), .B(new_new_n132_), .Y(new_new_n919_));
  NAi21      g0897(.An(new_new_n166_), .B(new_new_n462_), .Y(new_new_n920_));
  OAI220     g0898(.A0(new_new_n920_), .A1(new_new_n882_), .B0(new_new_n919_), .B1(new_new_n421_), .Y(new_new_n921_));
  NO2        g0899(.A(new_new_n921_), .B(new_new_n918_), .Y(new_new_n922_));
  NO2        g0900(.A(new_new_n411_), .B(new_new_n311_), .Y(new_new_n923_));
  NA2        g0901(.A(new_new_n923_), .B(new_new_n753_), .Y(new_new_n924_));
  NA2        g0902(.A(new_new_n614_), .B(i_0_), .Y(new_new_n925_));
  NO3        g0903(.A(new_new_n925_), .B(new_new_n406_), .C(new_new_n90_), .Y(new_new_n926_));
  NO4        g0904(.A(new_new_n631_), .B(new_new_n224_), .C(new_new_n440_), .D(new_new_n432_), .Y(new_new_n927_));
  AOI210     g0905(.A0(new_new_n927_), .A1(i_11_), .B0(new_new_n926_), .Y(new_new_n928_));
  INV        g0906(.A(new_new_n503_), .Y(new_new_n929_));
  AN2        g0907(.A(new_new_n100_), .B(new_new_n254_), .Y(new_new_n930_));
  NA2        g0908(.A(new_new_n791_), .B(new_new_n349_), .Y(new_new_n931_));
  AOI210     g0909(.A0(new_new_n514_), .A1(new_new_n90_), .B0(new_new_n59_), .Y(new_new_n932_));
  OAI220     g0910(.A0(new_new_n932_), .A1(new_new_n931_), .B0(new_new_n705_), .B1(new_new_n573_), .Y(new_new_n933_));
  NO2        g0911(.A(new_new_n265_), .B(new_new_n157_), .Y(new_new_n934_));
  NA2        g0912(.A(i_0_), .B(i_10_), .Y(new_new_n935_));
  AN2        g0913(.A(new_new_n934_), .B(i_6_), .Y(new_new_n936_));
  AOI220     g0914(.A0(new_new_n354_), .A1(new_new_n102_), .B0(new_new_n191_), .B1(new_new_n85_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n608_), .B(i_4_), .Y(new_new_n938_));
  NA2        g0916(.A(new_new_n194_), .B(new_new_n209_), .Y(new_new_n939_));
  OAI220     g0917(.A0(new_new_n939_), .A1(new_new_n931_), .B0(new_new_n938_), .B1(new_new_n937_), .Y(new_new_n940_));
  NO4        g0918(.A(new_new_n940_), .B(new_new_n936_), .C(new_new_n933_), .D(new_new_n930_), .Y(new_new_n941_));
  NA4        g0919(.A(new_new_n941_), .B(new_new_n928_), .C(new_new_n924_), .D(new_new_n922_), .Y(new_new_n942_));
  NO2        g0920(.A(new_new_n107_), .B(new_new_n37_), .Y(new_new_n943_));
  NA2        g0921(.A(i_11_), .B(i_9_), .Y(new_new_n944_));
  NO3        g0922(.A(i_12_), .B(new_new_n944_), .C(new_new_n648_), .Y(new_new_n945_));
  AO220      g0923(.A0(new_new_n945_), .A1(new_new_n943_), .B0(new_new_n283_), .B1(new_new_n89_), .Y(new_new_n946_));
  NO2        g0924(.A(new_new_n49_), .B(i_7_), .Y(new_new_n947_));
  NA2        g0925(.A(new_new_n416_), .B(new_new_n184_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n948_), .B(new_new_n164_), .Y(new_new_n949_));
  NO2        g0927(.A(new_new_n180_), .B(i_0_), .Y(new_new_n950_));
  INV        g0928(.A(new_new_n950_), .Y(new_new_n951_));
  NA2        g0929(.A(new_new_n503_), .B(new_new_n241_), .Y(new_new_n952_));
  AOI210     g0930(.A0(new_new_n391_), .A1(new_new_n42_), .B0(new_new_n429_), .Y(new_new_n953_));
  OAI220     g0931(.A0(new_new_n953_), .A1(new_new_n909_), .B0(new_new_n952_), .B1(new_new_n951_), .Y(new_new_n954_));
  NO3        g0932(.A(new_new_n954_), .B(new_new_n949_), .C(new_new_n946_), .Y(new_new_n955_));
  NA2        g0933(.A(new_new_n704_), .B(new_new_n124_), .Y(new_new_n956_));
  NO2        g0934(.A(i_6_), .B(new_new_n956_), .Y(new_new_n957_));
  AOI210     g0935(.A0(new_new_n472_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n958_));
  NA2        g0936(.A(new_new_n176_), .B(new_new_n107_), .Y(new_new_n959_));
  NOi32      g0937(.An(new_new_n958_), .Bn(new_new_n194_), .C(new_new_n959_), .Y(new_new_n960_));
  NO2        g0938(.A(new_new_n960_), .B(new_new_n957_), .Y(new_new_n961_));
  NOi21      g0939(.An(i_7_), .B(i_5_), .Y(new_new_n962_));
  NOi31      g0940(.An(new_new_n962_), .B(i_0_), .C(new_new_n769_), .Y(new_new_n963_));
  NA3        g0941(.A(new_new_n963_), .B(new_new_n405_), .C(i_6_), .Y(new_new_n964_));
  OA210      g0942(.A0(new_new_n959_), .A1(new_new_n551_), .B0(new_new_n964_), .Y(new_new_n965_));
  NO3        g0943(.A(new_new_n424_), .B(new_new_n385_), .C(new_new_n381_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n275_), .B(new_new_n338_), .Y(new_new_n967_));
  NO2        g0945(.A(new_new_n769_), .B(new_new_n270_), .Y(new_new_n968_));
  AOI210     g0946(.A0(new_new_n968_), .A1(new_new_n967_), .B0(new_new_n966_), .Y(new_new_n969_));
  NA4        g0947(.A(new_new_n969_), .B(new_new_n965_), .C(new_new_n961_), .D(new_new_n955_), .Y(new_new_n970_));
  NO2        g0948(.A(new_new_n916_), .B(new_new_n250_), .Y(new_new_n971_));
  AN2        g0949(.A(new_new_n353_), .B(new_new_n349_), .Y(new_new_n972_));
  AN2        g0950(.A(new_new_n972_), .B(new_new_n912_), .Y(new_new_n973_));
  OAI210     g0951(.A0(new_new_n973_), .A1(new_new_n971_), .B0(i_10_), .Y(new_new_n974_));
  OA210      g0952(.A0(new_new_n503_), .A1(new_new_n233_), .B0(new_new_n502_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n502_), .B(new_new_n433_), .C(new_new_n46_), .Y(new_new_n976_));
  OAI210     g0954(.A0(new_new_n920_), .A1(new_new_n929_), .B0(new_new_n976_), .Y(new_new_n977_));
  NO2        g0955(.A(new_new_n268_), .B(new_new_n47_), .Y(new_new_n978_));
  NO2        g0956(.A(new_new_n978_), .B(new_new_n193_), .Y(new_new_n979_));
  AOI220     g0957(.A0(new_new_n979_), .A1(new_new_n503_), .B0(new_new_n977_), .B1(new_new_n74_), .Y(new_new_n980_));
  NA3        g0958(.A(new_new_n863_), .B(new_new_n403_), .C(new_new_n686_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n96_), .B(new_new_n45_), .Y(new_new_n982_));
  NO2        g0960(.A(new_new_n76_), .B(new_new_n793_), .Y(new_new_n983_));
  AOI220     g0961(.A0(new_new_n983_), .A1(new_new_n982_), .B0(new_new_n179_), .B1(new_new_n639_), .Y(new_new_n984_));
  AOI210     g0962(.A0(new_new_n984_), .A1(new_new_n981_), .B0(new_new_n48_), .Y(new_new_n985_));
  NO3        g0963(.A(new_new_n631_), .B(new_new_n380_), .C(new_new_n24_), .Y(new_new_n986_));
  AOI210     g0964(.A0(new_new_n744_), .A1(new_new_n585_), .B0(new_new_n986_), .Y(new_new_n987_));
  NO2        g0965(.A(new_new_n644_), .B(new_new_n109_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n988_), .B(i_0_), .Y(new_new_n989_));
  OAI220     g0967(.A0(new_new_n989_), .A1(new_new_n87_), .B0(new_new_n987_), .B1(new_new_n177_), .Y(new_new_n990_));
  NO3        g0968(.A(new_new_n990_), .B(new_new_n985_), .C(new_new_n555_), .Y(new_new_n991_));
  NA3        g0969(.A(new_new_n991_), .B(new_new_n980_), .C(new_new_n974_), .Y(new_new_n992_));
  NO3        g0970(.A(new_new_n992_), .B(new_new_n970_), .C(new_new_n942_), .Y(new_new_n993_));
  NO2        g0971(.A(i_0_), .B(new_new_n769_), .Y(new_new_n994_));
  NA2        g0972(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n935_), .B(new_new_n995_), .Y(new_new_n996_));
  NO3        g0974(.A(new_new_n109_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n997_));
  AO220      g0975(.A0(new_new_n997_), .A1(new_new_n996_), .B0(new_new_n994_), .B1(new_new_n179_), .Y(new_new_n998_));
  NO2        g0976(.A(new_new_n842_), .B(new_new_n959_), .Y(new_new_n999_));
  AOI210     g0977(.A0(new_new_n998_), .A1(new_new_n370_), .B0(new_new_n999_), .Y(new_new_n1000_));
  NA2        g0978(.A(new_new_n779_), .B(new_new_n149_), .Y(new_new_n1001_));
  INV        g0979(.A(new_new_n1001_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n1002_), .B(new_new_n718_), .C(new_new_n74_), .Y(new_new_n1003_));
  NO2        g0981(.A(new_new_n859_), .B(new_new_n424_), .Y(new_new_n1004_));
  NA3        g0982(.A(new_new_n889_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n890_), .B(i_9_), .Y(new_new_n1006_));
  AOI210     g0984(.A0(new_new_n1005_), .A1(new_new_n531_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  OAI210     g0985(.A0(new_new_n255_), .A1(i_9_), .B0(new_new_n240_), .Y(new_new_n1008_));
  AOI210     g0986(.A0(new_new_n1008_), .A1(new_new_n925_), .B0(new_new_n157_), .Y(new_new_n1009_));
  NO3        g0987(.A(new_new_n1009_), .B(new_new_n1007_), .C(new_new_n1004_), .Y(new_new_n1010_));
  NA3        g0988(.A(new_new_n1010_), .B(new_new_n1003_), .C(new_new_n1000_), .Y(new_new_n1011_));
  NA2        g0989(.A(new_new_n972_), .B(new_new_n393_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n318_), .A1(new_new_n166_), .B0(new_new_n1012_), .Y(new_new_n1013_));
  NA3        g0991(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n1014_));
  NA2        g0992(.A(new_new_n947_), .B(new_new_n519_), .Y(new_new_n1015_));
  AOI210     g0993(.A0(new_new_n1014_), .A1(new_new_n166_), .B0(new_new_n1015_), .Y(new_new_n1016_));
  NO2        g0994(.A(new_new_n1016_), .B(new_new_n1013_), .Y(new_new_n1017_));
  NO3        g0995(.A(new_new_n935_), .B(new_new_n908_), .C(new_new_n196_), .Y(new_new_n1018_));
  AOI220     g0996(.A0(new_new_n1018_), .A1(i_11_), .B0(new_new_n609_), .B1(new_new_n76_), .Y(new_new_n1019_));
  NO3        g0997(.A(new_new_n218_), .B(new_new_n404_), .C(i_0_), .Y(new_new_n1020_));
  OAI210     g0998(.A0(new_new_n1020_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n1021_));
  INV        g0999(.A(new_new_n227_), .Y(new_new_n1022_));
  OAI220     g1000(.A0(new_new_n567_), .A1(new_new_n142_), .B0(new_new_n691_), .B1(new_new_n661_), .Y(new_new_n1023_));
  NA3        g1001(.A(new_new_n1023_), .B(i_7_), .C(new_new_n1022_), .Y(new_new_n1024_));
  NA4        g1002(.A(new_new_n1024_), .B(new_new_n1021_), .C(new_new_n1019_), .D(new_new_n1017_), .Y(new_new_n1025_));
  NO2        g1003(.A(new_new_n253_), .B(new_new_n96_), .Y(new_new_n1026_));
  NA2        g1004(.A(new_new_n1026_), .B(new_new_n994_), .Y(new_new_n1027_));
  AOI220     g1005(.A0(new_new_n962_), .A1(new_new_n519_), .B0(new_new_n889_), .B1(new_new_n167_), .Y(new_new_n1028_));
  NA2        g1006(.A(new_new_n373_), .B(new_new_n181_), .Y(new_new_n1029_));
  OA220      g1007(.A0(new_new_n1029_), .A1(new_new_n1028_), .B0(new_new_n1027_), .B1(i_5_), .Y(new_new_n1030_));
  AOI210     g1008(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n180_), .Y(new_new_n1031_));
  NA2        g1009(.A(new_new_n1031_), .B(new_new_n975_), .Y(new_new_n1032_));
  NA3        g1010(.A(new_new_n658_), .B(new_new_n191_), .C(new_new_n85_), .Y(new_new_n1033_));
  NA2        g1011(.A(new_new_n1033_), .B(new_new_n583_), .Y(new_new_n1034_));
  NA3        g1012(.A(new_new_n524_), .B(new_new_n517_), .C(new_new_n500_), .Y(new_new_n1035_));
  NO2        g1013(.A(new_new_n1035_), .B(new_new_n1034_), .Y(new_new_n1036_));
  NA3        g1014(.A(new_new_n411_), .B(new_new_n176_), .C(new_new_n175_), .Y(new_new_n1037_));
  NA3        g1015(.A(new_new_n947_), .B(new_new_n307_), .C(new_new_n240_), .Y(new_new_n1038_));
  NA2        g1016(.A(new_new_n1038_), .B(new_new_n1037_), .Y(new_new_n1039_));
  NA3        g1017(.A(new_new_n411_), .B(new_new_n355_), .C(new_new_n231_), .Y(new_new_n1040_));
  INV        g1018(.A(new_new_n1040_), .Y(new_new_n1041_));
  NOi31      g1019(.An(new_new_n410_), .B(new_new_n995_), .C(new_new_n250_), .Y(new_new_n1042_));
  NO3        g1020(.A(new_new_n944_), .B(new_new_n227_), .C(new_new_n196_), .Y(new_new_n1043_));
  NO4        g1021(.A(new_new_n1043_), .B(new_new_n1042_), .C(new_new_n1041_), .D(new_new_n1039_), .Y(new_new_n1044_));
  NA4        g1022(.A(new_new_n1044_), .B(new_new_n1036_), .C(new_new_n1032_), .D(new_new_n1030_), .Y(new_new_n1045_));
  INV        g1023(.A(new_new_n660_), .Y(new_new_n1046_));
  NO3        g1024(.A(new_new_n1046_), .B(new_new_n599_), .C(new_new_n367_), .Y(new_new_n1047_));
  INV        g1025(.A(new_new_n1047_), .Y(new_new_n1048_));
  NA3        g1026(.A(new_new_n324_), .B(i_5_), .C(new_new_n199_), .Y(new_new_n1049_));
  NAi31      g1027(.An(new_new_n252_), .B(new_new_n1049_), .C(new_new_n253_), .Y(new_new_n1050_));
  NO4        g1028(.A(new_new_n250_), .B(new_new_n218_), .C(i_0_), .D(i_12_), .Y(new_new_n1051_));
  AOI220     g1029(.A0(new_new_n1051_), .A1(new_new_n1050_), .B0(new_new_n838_), .B1(new_new_n181_), .Y(new_new_n1052_));
  AN2        g1030(.A(new_new_n935_), .B(new_new_n157_), .Y(new_new_n1053_));
  NO4        g1031(.A(new_new_n1053_), .B(i_12_), .C(new_new_n695_), .D(new_new_n134_), .Y(new_new_n1054_));
  NA2        g1032(.A(new_new_n1054_), .B(new_new_n227_), .Y(new_new_n1055_));
  NA3        g1033(.A(new_new_n102_), .B(new_new_n613_), .C(i_11_), .Y(new_new_n1056_));
  NO2        g1034(.A(new_new_n1056_), .B(new_new_n159_), .Y(new_new_n1057_));
  NA2        g1035(.A(new_new_n962_), .B(new_new_n499_), .Y(new_new_n1058_));
  NA2        g1036(.A(new_new_n65_), .B(new_new_n105_), .Y(new_new_n1059_));
  OAI220     g1037(.A0(new_new_n1059_), .A1(new_new_n1049_), .B0(new_new_n1058_), .B1(new_new_n719_), .Y(new_new_n1060_));
  AOI210     g1038(.A0(new_new_n1060_), .A1(new_new_n950_), .B0(new_new_n1057_), .Y(new_new_n1061_));
  NA4        g1039(.A(new_new_n1061_), .B(new_new_n1055_), .C(new_new_n1052_), .D(new_new_n1048_), .Y(new_new_n1062_));
  NO4        g1040(.A(new_new_n1062_), .B(new_new_n1045_), .C(new_new_n1025_), .D(new_new_n1011_), .Y(new_new_n1063_));
  OAI210     g1041(.A0(new_new_n862_), .A1(new_new_n855_), .B0(new_new_n37_), .Y(new_new_n1064_));
  NA3        g1042(.A(new_new_n958_), .B(new_new_n388_), .C(i_5_), .Y(new_new_n1065_));
  NA3        g1043(.A(new_new_n1065_), .B(new_new_n1064_), .C(new_new_n656_), .Y(new_new_n1066_));
  NA2        g1044(.A(new_new_n1066_), .B(new_new_n214_), .Y(new_new_n1067_));
  AN2        g1045(.A(new_new_n739_), .B(new_new_n389_), .Y(new_new_n1068_));
  NA2        g1046(.A(new_new_n192_), .B(new_new_n194_), .Y(new_new_n1069_));
  AO210      g1047(.A0(new_new_n1068_), .A1(new_new_n33_), .B0(new_new_n1069_), .Y(new_new_n1070_));
  OAI210     g1048(.A0(new_new_n660_), .A1(new_new_n658_), .B0(new_new_n337_), .Y(new_new_n1071_));
  NAi31      g1049(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1072_));
  AOI210     g1050(.A0(new_new_n120_), .A1(new_new_n71_), .B0(new_new_n1072_), .Y(new_new_n1073_));
  NO2        g1051(.A(new_new_n1073_), .B(new_new_n692_), .Y(new_new_n1074_));
  NA3        g1052(.A(new_new_n1074_), .B(new_new_n1071_), .C(new_new_n1070_), .Y(new_new_n1075_));
  NO2        g1053(.A(new_new_n489_), .B(new_new_n281_), .Y(new_new_n1076_));
  NO4        g1054(.A(new_new_n243_), .B(new_new_n148_), .C(new_new_n722_), .D(new_new_n37_), .Y(new_new_n1077_));
  NO3        g1055(.A(new_new_n1077_), .B(new_new_n1076_), .C(new_new_n927_), .Y(new_new_n1078_));
  OAI210     g1056(.A0(new_new_n1056_), .A1(new_new_n151_), .B0(new_new_n1078_), .Y(new_new_n1079_));
  AOI210     g1057(.A0(new_new_n1075_), .A1(new_new_n49_), .B0(new_new_n1079_), .Y(new_new_n1080_));
  AOI210     g1058(.A0(new_new_n1080_), .A1(new_new_n1067_), .B0(new_new_n74_), .Y(new_new_n1081_));
  NO2        g1059(.A(new_new_n606_), .B(new_new_n400_), .Y(new_new_n1082_));
  NO2        g1060(.A(new_new_n1082_), .B(new_new_n799_), .Y(new_new_n1083_));
  OAI210     g1061(.A0(new_new_n81_), .A1(new_new_n55_), .B0(new_new_n112_), .Y(new_new_n1084_));
  NA2        g1062(.A(new_new_n1084_), .B(new_new_n77_), .Y(new_new_n1085_));
  AOI210     g1063(.A0(new_new_n1031_), .A1(new_new_n947_), .B0(new_new_n963_), .Y(new_new_n1086_));
  AOI210     g1064(.A0(new_new_n1086_), .A1(new_new_n1085_), .B0(new_new_n722_), .Y(new_new_n1087_));
  NA2        g1065(.A(new_new_n275_), .B(new_new_n58_), .Y(new_new_n1088_));
  AOI220     g1066(.A0(new_new_n1088_), .A1(new_new_n77_), .B0(new_new_n368_), .B1(new_new_n267_), .Y(new_new_n1089_));
  NO2        g1067(.A(new_new_n1089_), .B(new_new_n247_), .Y(new_new_n1090_));
  NA3        g1068(.A(new_new_n100_), .B(new_new_n326_), .C(new_new_n31_), .Y(new_new_n1091_));
  INV        g1069(.A(new_new_n1091_), .Y(new_new_n1092_));
  NO3        g1070(.A(new_new_n1092_), .B(new_new_n1090_), .C(new_new_n1087_), .Y(new_new_n1093_));
  OAI210     g1071(.A0(new_new_n283_), .A1(new_new_n162_), .B0(new_new_n90_), .Y(new_new_n1094_));
  NA3        g1072(.A(new_new_n803_), .B(new_new_n307_), .C(new_new_n81_), .Y(new_new_n1095_));
  AOI210     g1073(.A0(new_new_n1095_), .A1(new_new_n1094_), .B0(i_11_), .Y(new_new_n1096_));
  NA2        g1074(.A(new_new_n651_), .B(new_new_n224_), .Y(new_new_n1097_));
  OAI210     g1075(.A0(new_new_n1097_), .A1(new_new_n958_), .B0(new_new_n214_), .Y(new_new_n1098_));
  NA2        g1076(.A(new_new_n168_), .B(i_5_), .Y(new_new_n1099_));
  NO2        g1077(.A(new_new_n1098_), .B(new_new_n1099_), .Y(new_new_n1100_));
  NO3        g1078(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n1101_));
  OAI210     g1079(.A0(new_new_n967_), .A1(new_new_n326_), .B0(new_new_n1101_), .Y(new_new_n1102_));
  NO2        g1080(.A(new_new_n1102_), .B(new_new_n769_), .Y(new_new_n1103_));
  NO3        g1081(.A(new_new_n1103_), .B(new_new_n1100_), .C(new_new_n1096_), .Y(new_new_n1104_));
  OAI210     g1082(.A0(new_new_n1093_), .A1(i_4_), .B0(new_new_n1104_), .Y(new_new_n1105_));
  NO3        g1083(.A(new_new_n1105_), .B(new_new_n1083_), .C(new_new_n1081_), .Y(new_new_n1106_));
  NA4        g1084(.A(new_new_n1106_), .B(new_new_n1063_), .C(new_new_n993_), .D(new_new_n915_), .Y(men4));
  INV        g1085(.A(new_new_n743_), .Y(new_new_n1110_));
  INV        g1086(.A(i_2_), .Y(new_new_n1111_));
  INV        g1087(.A(new_new_n514_), .Y(new_new_n1112_));
endmodule


