// Benchmark "data/9sym" written by ABC on Thu Jun 20 14:59:19 2024

module \data/9sym  ( 
    i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_,
    ori00  );
  input  i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;
  output ori00;
  ONE        g0(.Y(ori00));
endmodule


