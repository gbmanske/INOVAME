library verilog;
use verilog.vl_types.all;
entity maquinaVenda_vlg_vec_tst is
end maquinaVenda_vlg_vec_tst;
