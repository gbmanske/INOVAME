//Benchmark atmr_misex3_1774_0.5

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  NOi32      o000(.An(i), .Bn(g), .C(h), .Y(ori_ori_n29_));
  INV        o001(.A(h), .Y(ori_ori_n30_));
  INV        o002(.A(i), .Y(ori_ori_n31_));
  AN2        o003(.A(h), .B(g), .Y(ori_ori_n32_));
  NA2        o004(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NOi32      o005(.An(k), .Bn(h), .C(l), .Y(ori_ori_n34_));
  NOi32      o006(.An(k), .Bn(h), .C(g), .Y(ori_ori_n35_));
  INV        o007(.A(ori_ori_n35_), .Y(ori_ori_n36_));
  NO2        o008(.A(ori_ori_n36_), .B(n), .Y(ori_ori_n37_));
  INV        o009(.A(c), .Y(ori_ori_n38_));
  NA2        o010(.A(e), .B(b), .Y(ori_ori_n39_));
  INV        o011(.A(ori_ori_n39_), .Y(ori_ori_n40_));
  INV        o012(.A(d), .Y(ori_ori_n41_));
  NAi21      o013(.An(i), .B(h), .Y(ori_ori_n42_));
  NAi21      o014(.An(e), .B(h), .Y(ori_ori_n43_));
  INV        o015(.A(m), .Y(ori_ori_n44_));
  NOi21      o016(.An(k), .B(l), .Y(ori_ori_n45_));
  NA2        o017(.A(ori_ori_n45_), .B(ori_ori_n44_), .Y(ori_ori_n46_));
  AN4        o018(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n47_));
  NA2        o019(.A(h), .B(ori_ori_n47_), .Y(ori_ori_n48_));
  NAi32      o020(.An(m), .Bn(k), .C(j), .Y(ori_ori_n49_));
  OR2        o021(.A(ori_ori_n48_), .B(ori_ori_n46_), .Y(ori_ori_n50_));
  INV        o022(.A(ori_ori_n50_), .Y(ori_ori_n51_));
  INV        o023(.A(n), .Y(ori_ori_n52_));
  NOi32      o024(.An(e), .Bn(b), .C(d), .Y(ori_ori_n53_));
  INV        o025(.A(ori_ori_n53_), .Y(ori_ori_n54_));
  INV        o026(.A(j), .Y(ori_ori_n55_));
  AN3        o027(.A(m), .B(k), .C(i), .Y(ori_ori_n56_));
  NA3        o028(.A(ori_ori_n56_), .B(ori_ori_n55_), .C(g), .Y(ori_ori_n57_));
  NO2        o029(.A(ori_ori_n57_), .B(f), .Y(ori_ori_n58_));
  NAi32      o030(.An(g), .Bn(f), .C(h), .Y(ori_ori_n59_));
  NA2        o031(.A(m), .B(l), .Y(ori_ori_n60_));
  NOi32      o032(.An(m), .Bn(l), .C(i), .Y(ori_ori_n61_));
  NOi21      o033(.An(g), .B(i), .Y(ori_ori_n62_));
  NAi41      o034(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n63_));
  AN2        o035(.A(e), .B(b), .Y(ori_ori_n64_));
  NOi31      o036(.An(c), .B(h), .C(f), .Y(ori_ori_n65_));
  NA2        o037(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  NO2        o038(.A(ori_ori_n66_), .B(ori_ori_n63_), .Y(ori_ori_n67_));
  NOi21      o039(.An(i), .B(h), .Y(ori_ori_n68_));
  INV        o040(.A(a), .Y(ori_ori_n69_));
  NA2        o041(.A(ori_ori_n64_), .B(ori_ori_n69_), .Y(ori_ori_n70_));
  INV        o042(.A(l), .Y(ori_ori_n71_));
  NOi21      o043(.An(m), .B(n), .Y(ori_ori_n72_));
  INV        o044(.A(b), .Y(ori_ori_n73_));
  INV        o045(.A(ori_ori_n67_), .Y(ori_ori_n74_));
  OAI210     o046(.A0(ori_ori_n57_), .A1(ori_ori_n54_), .B0(ori_ori_n74_), .Y(ori_ori_n75_));
  NOi31      o047(.An(k), .B(m), .C(j), .Y(ori_ori_n76_));
  NA3        o048(.A(ori_ori_n76_), .B(h), .C(ori_ori_n47_), .Y(ori_ori_n77_));
  NOi31      o049(.An(k), .B(m), .C(i), .Y(ori_ori_n78_));
  INV        o050(.A(ori_ori_n77_), .Y(ori_ori_n79_));
  NOi32      o051(.An(f), .Bn(b), .C(e), .Y(ori_ori_n80_));
  NAi21      o052(.An(m), .B(n), .Y(ori_ori_n81_));
  NAi21      o053(.An(j), .B(k), .Y(ori_ori_n82_));
  NO3        o054(.A(ori_ori_n82_), .B(ori_ori_n81_), .C(g), .Y(ori_ori_n83_));
  NAi31      o055(.An(j), .B(k), .C(h), .Y(ori_ori_n84_));
  NA2        o056(.A(ori_ori_n83_), .B(ori_ori_n80_), .Y(ori_ori_n85_));
  INV        o057(.A(ori_ori_n81_), .Y(ori_ori_n86_));
  AN2        o058(.A(k), .B(j), .Y(ori_ori_n87_));
  NO3        o059(.A(c), .B(ori_ori_n87_), .C(g), .Y(ori_ori_n88_));
  NAi31      o060(.An(f), .B(e), .C(b), .Y(ori_ori_n89_));
  NA2        o061(.A(ori_ori_n88_), .B(ori_ori_n86_), .Y(ori_ori_n90_));
  NA2        o062(.A(d), .B(b), .Y(ori_ori_n91_));
  NAi21      o063(.An(e), .B(f), .Y(ori_ori_n92_));
  NAi21      o064(.An(e), .B(g), .Y(ori_ori_n93_));
  NAi21      o065(.An(c), .B(d), .Y(ori_ori_n94_));
  NAi31      o066(.An(l), .B(k), .C(h), .Y(ori_ori_n95_));
  NAi31      o067(.An(ori_ori_n79_), .B(ori_ori_n90_), .C(ori_ori_n85_), .Y(ori_ori_n96_));
  NAi31      o068(.An(e), .B(f), .C(b), .Y(ori_ori_n97_));
  NOi21      o069(.An(h), .B(i), .Y(ori_ori_n98_));
  NOi21      o070(.An(k), .B(m), .Y(ori_ori_n99_));
  NOi21      o071(.An(h), .B(g), .Y(ori_ori_n100_));
  NAi31      o072(.An(d), .B(f), .C(c), .Y(ori_ori_n101_));
  NAi31      o073(.An(e), .B(f), .C(c), .Y(ori_ori_n102_));
  NA2        o074(.A(j), .B(h), .Y(ori_ori_n103_));
  OR3        o075(.A(n), .B(m), .C(k), .Y(ori_ori_n104_));
  NO2        o076(.A(ori_ori_n104_), .B(ori_ori_n103_), .Y(ori_ori_n105_));
  NAi32      o077(.An(m), .Bn(k), .C(n), .Y(ori_ori_n106_));
  NA2        o078(.A(ori_ori_n105_), .B(f), .Y(ori_ori_n107_));
  NO2        o079(.A(n), .B(m), .Y(ori_ori_n108_));
  NA2        o080(.A(ori_ori_n108_), .B(ori_ori_n34_), .Y(ori_ori_n109_));
  NAi21      o081(.An(f), .B(e), .Y(ori_ori_n110_));
  NAi21      o082(.An(h), .B(f), .Y(ori_ori_n111_));
  INV        o083(.A(ori_ori_n111_), .Y(ori_ori_n112_));
  NO2        o084(.A(m), .B(ori_ori_n94_), .Y(ori_ori_n113_));
  NA2        o085(.A(ori_ori_n113_), .B(ori_ori_n112_), .Y(ori_ori_n114_));
  NOi32      o086(.An(f), .Bn(c), .C(d), .Y(ori_ori_n115_));
  NOi32      o087(.An(f), .Bn(c), .C(e), .Y(ori_ori_n116_));
  NO2        o088(.A(ori_ori_n116_), .B(ori_ori_n115_), .Y(ori_ori_n117_));
  NO3        o089(.A(n), .B(m), .C(j), .Y(ori_ori_n118_));
  NA2        o090(.A(ori_ori_n118_), .B(k), .Y(ori_ori_n119_));
  BUFFER     o091(.A(ori_ori_n109_), .Y(ori_ori_n120_));
  NA3        o092(.A(ori_ori_n120_), .B(ori_ori_n114_), .C(ori_ori_n107_), .Y(ori_ori_n121_));
  OR2        o093(.A(ori_ori_n121_), .B(ori_ori_n96_), .Y(ori_ori_n122_));
  NO3        o094(.A(ori_ori_n122_), .B(ori_ori_n75_), .C(ori_ori_n51_), .Y(ori_ori_n123_));
  NAi31      o095(.An(n), .B(h), .C(g), .Y(ori_ori_n124_));
  NOi32      o096(.An(m), .Bn(k), .C(l), .Y(ori_ori_n125_));
  NA3        o097(.A(ori_ori_n125_), .B(ori_ori_n55_), .C(g), .Y(ori_ori_n126_));
  NOi21      o098(.An(k), .B(j), .Y(ori_ori_n127_));
  NA4        o099(.A(ori_ori_n127_), .B(ori_ori_n72_), .C(i), .D(g), .Y(ori_ori_n128_));
  NAi41      o100(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n129_));
  INV        o101(.A(f), .Y(ori_ori_n130_));
  INV        o102(.A(g), .Y(ori_ori_n131_));
  NOi31      o103(.An(i), .B(j), .C(h), .Y(ori_ori_n132_));
  NOi21      o104(.An(l), .B(m), .Y(ori_ori_n133_));
  NA2        o105(.A(ori_ori_n133_), .B(ori_ori_n132_), .Y(ori_ori_n134_));
  NO3        o106(.A(ori_ori_n134_), .B(ori_ori_n131_), .C(ori_ori_n130_), .Y(ori_ori_n135_));
  NOi21      o107(.An(n), .B(m), .Y(ori_ori_n136_));
  OR2        o108(.A(ori_ori_n49_), .B(ori_ori_n48_), .Y(ori_ori_n137_));
  NAi21      o109(.An(j), .B(h), .Y(ori_ori_n138_));
  NOi31      o110(.An(k), .B(n), .C(m), .Y(ori_ori_n139_));
  NOi21      o111(.An(ori_ori_n139_), .B(ori_ori_n110_), .Y(ori_ori_n140_));
  INV        o112(.A(ori_ori_n140_), .Y(ori_ori_n141_));
  NAi31      o113(.An(f), .B(e), .C(c), .Y(ori_ori_n142_));
  NO4        o114(.A(ori_ori_n142_), .B(ori_ori_n104_), .C(ori_ori_n103_), .D(ori_ori_n41_), .Y(ori_ori_n143_));
  NA3        o115(.A(e), .B(c), .C(b), .Y(ori_ori_n144_));
  NAi32      o116(.An(m), .Bn(i), .C(k), .Y(ori_ori_n145_));
  INV        o117(.A(k), .Y(ori_ori_n146_));
  INV        o118(.A(ori_ori_n143_), .Y(ori_ori_n147_));
  NAi41      o119(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n148_));
  NO2        o120(.A(ori_ori_n148_), .B(e), .Y(ori_ori_n149_));
  AN3        o121(.A(ori_ori_n147_), .B(ori_ori_n141_), .C(ori_ori_n137_), .Y(ori_ori_n150_));
  NO2        o122(.A(h), .B(ori_ori_n63_), .Y(ori_ori_n151_));
  NA2        o123(.A(ori_ori_n151_), .B(ori_ori_n80_), .Y(ori_ori_n152_));
  NAi41      o124(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n153_));
  NO2        o125(.A(ori_ori_n153_), .B(ori_ori_n130_), .Y(ori_ori_n154_));
  NA2        o126(.A(ori_ori_n99_), .B(ori_ori_n68_), .Y(ori_ori_n155_));
  NO2        o127(.A(n), .B(a), .Y(ori_ori_n156_));
  NAi21      o128(.An(h), .B(i), .Y(ori_ori_n157_));
  NA2        o129(.A(ori_ori_n108_), .B(k), .Y(ori_ori_n158_));
  NO2        o130(.A(ori_ori_n158_), .B(ori_ori_n157_), .Y(ori_ori_n159_));
  INV        o131(.A(ori_ori_n159_), .Y(ori_ori_n160_));
  NA2        o132(.A(ori_ori_n160_), .B(ori_ori_n152_), .Y(ori_ori_n161_));
  NOi21      o133(.An(g), .B(e), .Y(ori_ori_n162_));
  NOi21      o134(.An(ori_ori_n150_), .B(ori_ori_n161_), .Y(ori_ori_n163_));
  NA3        o135(.A(ori_ori_n41_), .B(c), .C(b), .Y(ori_ori_n164_));
  NO2        o136(.A(ori_ori_n155_), .B(f), .Y(ori_ori_n165_));
  NAi31      o137(.An(g), .B(k), .C(h), .Y(ori_ori_n166_));
  NA2        o138(.A(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n167_));
  NO2        o139(.A(ori_ori_n167_), .B(ori_ori_n117_), .Y(ori_ori_n168_));
  NA3        o140(.A(e), .B(c), .C(b), .Y(ori_ori_n169_));
  NAi32      o141(.An(j), .Bn(h), .C(i), .Y(ori_ori_n170_));
  NAi21      o142(.An(m), .B(l), .Y(ori_ori_n171_));
  NA2        o143(.A(h), .B(g), .Y(ori_ori_n172_));
  NO2        o144(.A(ori_ori_n89_), .B(d), .Y(ori_ori_n173_));
  NA2        o145(.A(ori_ori_n173_), .B(ori_ori_n37_), .Y(ori_ori_n174_));
  NO2        o146(.A(ori_ori_n66_), .B(ori_ori_n63_), .Y(ori_ori_n175_));
  NAi32      o147(.An(n), .Bn(m), .C(l), .Y(ori_ori_n176_));
  NO2        o148(.A(ori_ori_n176_), .B(ori_ori_n170_), .Y(ori_ori_n177_));
  NA2        o149(.A(ori_ori_n177_), .B(c), .Y(ori_ori_n178_));
  NA2        o150(.A(ori_ori_n178_), .B(ori_ori_n174_), .Y(ori_ori_n179_));
  NO2        o151(.A(ori_ori_n179_), .B(ori_ori_n168_), .Y(ori_ori_n180_));
  NAi21      o152(.An(m), .B(k), .Y(ori_ori_n181_));
  INV        o153(.A(ori_ori_n181_), .Y(ori_ori_n182_));
  NAi41      o154(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n183_));
  NO2        o155(.A(ori_ori_n183_), .B(ori_ori_n93_), .Y(ori_ori_n184_));
  NA2        o156(.A(ori_ori_n184_), .B(ori_ori_n182_), .Y(ori_ori_n185_));
  NOi21      o157(.An(f), .B(h), .Y(ori_ori_n186_));
  NAi31      o158(.An(d), .B(e), .C(b), .Y(ori_ori_n187_));
  NO2        o159(.A(ori_ori_n81_), .B(ori_ori_n187_), .Y(ori_ori_n188_));
  NA2        o160(.A(ori_ori_n188_), .B(ori_ori_n186_), .Y(ori_ori_n189_));
  NA2        o161(.A(ori_ori_n189_), .B(ori_ori_n185_), .Y(ori_ori_n190_));
  NO3        o162(.A(ori_ori_n183_), .B(ori_ori_n49_), .C(ori_ori_n43_), .Y(ori_ori_n191_));
  NA2        o163(.A(ori_ori_n156_), .B(ori_ori_n64_), .Y(ori_ori_n192_));
  OR2        o164(.A(ori_ori_n192_), .B(ori_ori_n126_), .Y(ori_ori_n193_));
  NOi31      o165(.An(l), .B(n), .C(m), .Y(ori_ori_n194_));
  NA2        o166(.A(ori_ori_n194_), .B(ori_ori_n132_), .Y(ori_ori_n195_));
  NAi21      o167(.An(ori_ori_n191_), .B(ori_ori_n193_), .Y(ori_ori_n196_));
  NAi32      o168(.An(m), .Bn(j), .C(k), .Y(ori_ori_n197_));
  NAi41      o169(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n198_));
  NOi31      o170(.An(j), .B(m), .C(k), .Y(ori_ori_n199_));
  NO2        o171(.A(ori_ori_n76_), .B(ori_ori_n199_), .Y(ori_ori_n200_));
  NAi31      o172(.An(ori_ori_n200_), .B(f), .C(e), .Y(ori_ori_n201_));
  NOi32      o173(.An(m), .Bn(j), .C(l), .Y(ori_ori_n202_));
  NO2        o174(.A(ori_ori_n202_), .B(ori_ori_n61_), .Y(ori_ori_n203_));
  NAi32      o175(.An(ori_ori_n203_), .Bn(ori_ori_n124_), .C(ori_ori_n173_), .Y(ori_ori_n204_));
  NO2        o176(.A(ori_ori_n171_), .B(ori_ori_n170_), .Y(ori_ori_n205_));
  NO2        o177(.A(ori_ori_n134_), .B(g), .Y(ori_ori_n206_));
  INV        o178(.A(ori_ori_n97_), .Y(ori_ori_n207_));
  AOI220     o179(.A0(ori_ori_n207_), .A1(ori_ori_n206_), .B0(ori_ori_n154_), .B1(ori_ori_n205_), .Y(ori_ori_n208_));
  NA3        o180(.A(ori_ori_n208_), .B(ori_ori_n204_), .C(ori_ori_n201_), .Y(ori_ori_n209_));
  NA3        o181(.A(h), .B(g), .C(f), .Y(ori_ori_n210_));
  NO2        o182(.A(ori_ori_n210_), .B(ori_ori_n46_), .Y(ori_ori_n211_));
  NA2        o183(.A(ori_ori_n100_), .B(e), .Y(ori_ori_n212_));
  NA2        o184(.A(e), .B(ori_ori_n211_), .Y(ori_ori_n213_));
  NOi32      o185(.An(j), .Bn(g), .C(i), .Y(ori_ori_n214_));
  NOi32      o186(.An(e), .Bn(b), .C(a), .Y(ori_ori_n215_));
  NA2        o187(.A(ori_ori_n35_), .B(ori_ori_n72_), .Y(ori_ori_n216_));
  INV        o188(.A(ori_ori_n213_), .Y(ori_ori_n217_));
  NO4        o189(.A(ori_ori_n217_), .B(ori_ori_n209_), .C(ori_ori_n196_), .D(ori_ori_n190_), .Y(ori_ori_n218_));
  NA4        o190(.A(ori_ori_n218_), .B(ori_ori_n180_), .C(ori_ori_n163_), .D(ori_ori_n123_), .Y(ori10));
  NA3        o191(.A(m), .B(k), .C(i), .Y(ori_ori_n220_));
  NOi21      o192(.An(e), .B(f), .Y(ori_ori_n221_));
  NO3        o193(.A(ori_ori_n94_), .B(n), .C(ori_ori_n69_), .Y(ori_ori_n222_));
  NAi31      o194(.An(b), .B(f), .C(c), .Y(ori_ori_n223_));
  INV        o195(.A(ori_ori_n223_), .Y(ori_ori_n224_));
  NOi32      o196(.An(k), .Bn(h), .C(j), .Y(ori_ori_n225_));
  NA2        o197(.A(ori_ori_n225_), .B(ori_ori_n136_), .Y(ori_ori_n226_));
  AN2        o198(.A(j), .B(h), .Y(ori_ori_n227_));
  NO3        o199(.A(n), .B(m), .C(k), .Y(ori_ori_n228_));
  NA2        o200(.A(ori_ori_n228_), .B(ori_ori_n227_), .Y(ori_ori_n229_));
  NO2        o201(.A(ori_ori_n229_), .B(ori_ori_n94_), .Y(ori_ori_n230_));
  OR2        o202(.A(m), .B(k), .Y(ori_ori_n231_));
  NO2        o203(.A(ori_ori_n103_), .B(ori_ori_n231_), .Y(ori_ori_n232_));
  NA4        o204(.A(n), .B(f), .C(c), .D(ori_ori_n73_), .Y(ori_ori_n233_));
  NOi21      o205(.An(ori_ori_n232_), .B(ori_ori_n233_), .Y(ori_ori_n234_));
  NOi32      o206(.An(d), .Bn(a), .C(c), .Y(ori_ori_n235_));
  NA2        o207(.A(ori_ori_n235_), .B(ori_ori_n110_), .Y(ori_ori_n236_));
  NA2        o208(.A(f), .B(ori_ori_n177_), .Y(ori_ori_n237_));
  NO2        o209(.A(ori_ori_n41_), .B(ori_ori_n73_), .Y(ori_ori_n238_));
  NA2        o210(.A(ori_ori_n156_), .B(ori_ori_n238_), .Y(ori_ori_n239_));
  NA3        o211(.A(m), .B(g), .C(e), .Y(ori_ori_n240_));
  NO2        o212(.A(ori_ori_n240_), .B(ori_ori_n239_), .Y(ori_ori_n241_));
  NA3        o213(.A(ori_ori_n235_), .B(ori_ori_n110_), .C(ori_ori_n52_), .Y(ori_ori_n242_));
  NA2        o214(.A(ori_ori_n35_), .B(m), .Y(ori_ori_n243_));
  NO2        o215(.A(ori_ori_n243_), .B(ori_ori_n92_), .Y(ori_ori_n244_));
  NO3        o216(.A(ori_ori_n244_), .B(ori_ori_n241_), .C(ori_ori_n230_), .Y(ori_ori_n245_));
  NA2        o217(.A(i), .B(g), .Y(ori_ori_n246_));
  OR2        o218(.A(n), .B(m), .Y(ori_ori_n247_));
  NO2        o219(.A(ori_ori_n247_), .B(ori_ori_n95_), .Y(ori_ori_n248_));
  NAi21      o220(.An(k), .B(j), .Y(ori_ori_n249_));
  NOi31      o221(.An(n), .B(m), .C(k), .Y(ori_ori_n250_));
  AOI220     o222(.A0(ori_ori_n250_), .A1(ori_ori_n227_), .B0(ori_ori_n136_), .B1(ori_ori_n34_), .Y(ori_ori_n251_));
  NAi31      o223(.An(g), .B(f), .C(c), .Y(ori_ori_n252_));
  INV        o224(.A(ori_ori_n166_), .Y(ori_ori_n253_));
  NO2        o225(.A(ori_ori_n242_), .B(ori_ori_n126_), .Y(ori_ori_n254_));
  NA2        o226(.A(l), .B(k), .Y(ori_ori_n255_));
  NO2        o227(.A(ori_ori_n673_), .B(ori_ori_n254_), .Y(ori_ori_n256_));
  INV        o228(.A(ori_ori_n111_), .Y(ori_ori_n257_));
  OAI210     o229(.A0(j), .A1(ori_ori_n81_), .B0(ori_ori_n63_), .Y(ori_ori_n258_));
  NA2        o230(.A(ori_ori_n258_), .B(ori_ori_n257_), .Y(ori_ori_n259_));
  NO3        o231(.A(ori_ori_n236_), .B(ori_ori_n203_), .C(ori_ori_n124_), .Y(ori_ori_n260_));
  NO2        o232(.A(ori_ori_n236_), .B(ori_ori_n216_), .Y(ori_ori_n261_));
  NO3        o233(.A(ori_ori_n261_), .B(ori_ori_n260_), .C(ori_ori_n175_), .Y(ori_ori_n262_));
  NA3        o234(.A(ori_ori_n262_), .B(ori_ori_n259_), .C(ori_ori_n150_), .Y(ori_ori_n263_));
  OAI210     o235(.A0(ori_ori_n78_), .A1(ori_ori_n76_), .B0(n), .Y(ori_ori_n264_));
  NO2        o236(.A(ori_ori_n264_), .B(g), .Y(ori_ori_n265_));
  XO2        o237(.A(i), .B(h), .Y(ori_ori_n266_));
  NA3        o238(.A(ori_ori_n266_), .B(ori_ori_n99_), .C(n), .Y(ori_ori_n267_));
  NA3        o239(.A(ori_ori_n267_), .B(ori_ori_n251_), .C(ori_ori_n226_), .Y(ori_ori_n268_));
  AN2        o240(.A(ori_ori_n268_), .B(f), .Y(ori_ori_n269_));
  NAi31      o241(.An(c), .B(f), .C(d), .Y(ori_ori_n270_));
  BUFFER     o242(.A(ori_ori_n50_), .Y(ori_ori_n271_));
  NA2        o243(.A(ori_ori_n139_), .B(ori_ori_n68_), .Y(ori_ori_n272_));
  NA2        o244(.A(ori_ori_n272_), .B(ori_ori_n109_), .Y(ori_ori_n273_));
  INV        o245(.A(ori_ori_n273_), .Y(ori_ori_n274_));
  NA2        o246(.A(ori_ori_n274_), .B(ori_ori_n271_), .Y(ori_ori_n275_));
  NO3        o247(.A(ori_ori_n275_), .B(ori_ori_n269_), .C(ori_ori_n263_), .Y(ori_ori_n276_));
  NA4        o248(.A(ori_ori_n276_), .B(ori_ori_n256_), .C(ori_ori_n195_), .D(ori_ori_n245_), .Y(ori11));
  INV        o249(.A(g), .Y(ori_ori_n278_));
  NAi31      o250(.An(i), .B(m), .C(l), .Y(ori_ori_n279_));
  INV        o251(.A(k), .Y(ori_ori_n280_));
  NOi32      o252(.An(e), .Bn(b), .C(f), .Y(ori_ori_n281_));
  NA2        o253(.A(ori_ori_n32_), .B(j), .Y(ori_ori_n282_));
  NAi31      o254(.An(d), .B(e), .C(a), .Y(ori_ori_n283_));
  NO2        o255(.A(ori_ori_n283_), .B(n), .Y(ori_ori_n284_));
  NA2        o256(.A(j), .B(i), .Y(ori_ori_n285_));
  NA2        o257(.A(ori_ori_n87_), .B(ori_ori_n29_), .Y(ori_ori_n286_));
  OAI220     o258(.A0(ori_ori_n286_), .A1(m), .B0(ori_ori_n282_), .B1(ori_ori_n145_), .Y(ori_ori_n287_));
  NOi41      o259(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n288_));
  NAi32      o260(.An(e), .Bn(b), .C(c), .Y(ori_ori_n289_));
  OR2        o261(.A(ori_ori_n289_), .B(ori_ori_n52_), .Y(ori_ori_n290_));
  AN2        o262(.A(ori_ori_n198_), .B(ori_ori_n183_), .Y(ori_ori_n291_));
  NA2        o263(.A(ori_ori_n291_), .B(ori_ori_n290_), .Y(ori_ori_n292_));
  OA210      o264(.A0(ori_ori_n292_), .A1(ori_ori_n288_), .B0(ori_ori_n287_), .Y(ori_ori_n293_));
  NO2        o265(.A(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n294_));
  NA2        o266(.A(ori_ori_n294_), .B(ori_ori_n40_), .Y(ori_ori_n295_));
  INV        o267(.A(ori_ori_n295_), .Y(ori_ori_n296_));
  AN3        o268(.A(j), .B(h), .C(g), .Y(ori_ori_n297_));
  NO2        o269(.A(ori_ori_n91_), .B(c), .Y(ori_ori_n298_));
  NA3        o270(.A(ori_ori_n298_), .B(ori_ori_n297_), .C(ori_ori_n250_), .Y(ori_ori_n299_));
  NA3        o271(.A(f), .B(d), .C(b), .Y(ori_ori_n300_));
  INV        o272(.A(ori_ori_n299_), .Y(ori_ori_n301_));
  NO3        o273(.A(ori_ori_n301_), .B(ori_ori_n296_), .C(ori_ori_n293_), .Y(ori_ori_n302_));
  INV        o274(.A(k), .Y(ori_ori_n303_));
  NAi41      o275(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n304_));
  OAI210     o276(.A0(ori_ori_n283_), .A1(n), .B0(ori_ori_n304_), .Y(ori_ori_n305_));
  NAi31      o277(.An(f), .B(h), .C(g), .Y(ori_ori_n306_));
  NO3        o278(.A(ori_ori_n181_), .B(ori_ori_n42_), .C(n), .Y(ori_ori_n307_));
  NA3        o279(.A(ori_ori_n270_), .B(ori_ori_n102_), .C(ori_ori_n101_), .Y(ori_ori_n308_));
  NA2        o280(.A(ori_ori_n252_), .B(ori_ori_n142_), .Y(ori_ori_n309_));
  OR2        o281(.A(ori_ori_n309_), .B(ori_ori_n308_), .Y(ori_ori_n310_));
  NA2        o282(.A(ori_ori_n310_), .B(ori_ori_n307_), .Y(ori_ori_n311_));
  INV        o283(.A(ori_ori_n311_), .Y(ori_ori_n312_));
  NA3        o284(.A(ori_ori_n288_), .B(ori_ori_n199_), .C(ori_ori_n32_), .Y(ori_ori_n313_));
  NOi32      o285(.An(e), .Bn(c), .C(f), .Y(ori_ori_n314_));
  INV        o286(.A(ori_ori_n129_), .Y(ori_ori_n315_));
  AOI220     o287(.A0(ori_ori_n315_), .A1(ori_ori_n232_), .B0(ori_ori_n314_), .B1(ori_ori_n105_), .Y(ori_ori_n316_));
  NA3        o288(.A(ori_ori_n316_), .B(ori_ori_n313_), .C(ori_ori_n107_), .Y(ori_ori_n317_));
  INV        o289(.A(m), .Y(ori_ori_n318_));
  NO2        o290(.A(k), .B(ori_ori_n131_), .Y(ori_ori_n319_));
  INV        o291(.A(ori_ori_n215_), .Y(ori_ori_n320_));
  NO2        o292(.A(ori_ori_n320_), .B(n), .Y(ori_ori_n321_));
  NAi31      o293(.An(ori_ori_n318_), .B(ori_ori_n321_), .C(ori_ori_n319_), .Y(ori_ori_n322_));
  NO2        o294(.A(ori_ori_n282_), .B(ori_ori_n106_), .Y(ori_ori_n323_));
  NA2        o295(.A(ori_ori_n266_), .B(ori_ori_n99_), .Y(ori_ori_n324_));
  NA2        o296(.A(c), .B(ori_ori_n323_), .Y(ori_ori_n325_));
  AN3        o297(.A(f), .B(d), .C(b), .Y(ori_ori_n326_));
  OAI210     o298(.A0(ori_ori_n326_), .A1(ori_ori_n80_), .B0(n), .Y(ori_ori_n327_));
  NA2        o299(.A(ori_ori_n266_), .B(ori_ori_n99_), .Y(ori_ori_n328_));
  AOI210     o300(.A0(ori_ori_n327_), .A1(ori_ori_n144_), .B0(ori_ori_n328_), .Y(ori_ori_n329_));
  NAi31      o301(.An(m), .B(n), .C(k), .Y(ori_ori_n330_));
  NA2        o302(.A(ori_ori_n329_), .B(j), .Y(ori_ori_n331_));
  NA3        o303(.A(ori_ori_n331_), .B(ori_ori_n325_), .C(ori_ori_n322_), .Y(ori_ori_n332_));
  NO3        o304(.A(ori_ori_n332_), .B(ori_ori_n317_), .C(ori_ori_n312_), .Y(ori_ori_n333_));
  NA2        o305(.A(ori_ori_n222_), .B(ori_ori_n100_), .Y(ori_ori_n334_));
  NAi31      o306(.An(g), .B(h), .C(f), .Y(ori_ori_n335_));
  OA210      o307(.A0(ori_ori_n283_), .A1(n), .B0(ori_ori_n304_), .Y(ori_ori_n336_));
  NO2        o308(.A(ori_ori_n334_), .B(ori_ori_n280_), .Y(ori_ori_n337_));
  NO3        o309(.A(g), .B(ori_ori_n130_), .C(ori_ori_n38_), .Y(ori_ori_n338_));
  OAI210     o310(.A0(ori_ori_n139_), .A1(ori_ori_n232_), .B0(ori_ori_n338_), .Y(ori_ori_n339_));
  INV        o311(.A(ori_ori_n339_), .Y(ori_ori_n340_));
  NA2        o312(.A(ori_ori_n188_), .B(ori_ori_n87_), .Y(ori_ori_n341_));
  NO2        o313(.A(ori_ori_n341_), .B(ori_ori_n42_), .Y(ori_ori_n342_));
  NO3        o314(.A(ori_ori_n252_), .B(ori_ori_n103_), .C(i), .Y(ori_ori_n343_));
  NO3        o315(.A(ori_ori_n342_), .B(ori_ori_n340_), .C(ori_ori_n337_), .Y(ori_ori_n344_));
  NA3        o316(.A(ori_ori_n344_), .B(ori_ori_n333_), .C(ori_ori_n302_), .Y(ori08));
  NO2        o317(.A(k), .B(h), .Y(ori_ori_n346_));
  OR2        o318(.A(ori_ori_n157_), .B(ori_ori_n346_), .Y(ori_ori_n347_));
  NO2        o319(.A(ori_ori_n347_), .B(ori_ori_n171_), .Y(ori_ori_n348_));
  NA2        o320(.A(ori_ori_n314_), .B(ori_ori_n52_), .Y(ori_ori_n349_));
  NA2        o321(.A(ori_ori_n349_), .B(ori_ori_n252_), .Y(ori_ori_n350_));
  NA2        o322(.A(ori_ori_n350_), .B(ori_ori_n348_), .Y(ori_ori_n351_));
  NA2        o323(.A(ori_ori_n52_), .B(ori_ori_n69_), .Y(ori_ori_n352_));
  NO2        o324(.A(ori_ori_n352_), .B(ori_ori_n39_), .Y(ori_ori_n353_));
  NO3        o325(.A(ori_ori_n220_), .B(j), .C(ori_ori_n131_), .Y(ori_ori_n354_));
  NA2        o326(.A(ori_ori_n354_), .B(ori_ori_n353_), .Y(ori_ori_n355_));
  AOI210     o327(.A0(ori_ori_n300_), .A1(ori_ori_n97_), .B0(ori_ori_n52_), .Y(ori_ori_n356_));
  NA3        o328(.A(ori_ori_n133_), .B(ori_ori_n31_), .C(h), .Y(ori_ori_n357_));
  NA3        o329(.A(l), .B(ori_ori_n68_), .C(ori_ori_n44_), .Y(ori_ori_n358_));
  OAI210     o330(.A0(ori_ori_n357_), .A1(g), .B0(ori_ori_n358_), .Y(ori_ori_n359_));
  NA2        o331(.A(ori_ori_n359_), .B(ori_ori_n356_), .Y(ori_ori_n360_));
  NA4        o332(.A(ori_ori_n360_), .B(ori_ori_n355_), .C(ori_ori_n351_), .D(ori_ori_n208_), .Y(ori_ori_n361_));
  NO3        o333(.A(ori_ori_n103_), .B(ori_ori_n231_), .C(g), .Y(ori_ori_n362_));
  NA2        o334(.A(ori_ori_n362_), .B(e), .Y(ori_ori_n363_));
  NA2        o335(.A(ori_ori_n315_), .B(ori_ori_n205_), .Y(ori_ori_n364_));
  NA2        o336(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n365_));
  NO3        o337(.A(ori_ori_n181_), .B(g), .C(j), .Y(ori_ori_n366_));
  NAi21      o338(.An(ori_ori_n366_), .B(ori_ori_n358_), .Y(ori_ori_n367_));
  NA2        o339(.A(ori_ori_n367_), .B(ori_ori_n47_), .Y(ori_ori_n368_));
  INV        o340(.A(ori_ori_n368_), .Y(ori_ori_n369_));
  NO3        o341(.A(ori_ori_n369_), .B(ori_ori_n365_), .C(ori_ori_n361_), .Y(ori_ori_n370_));
  NA2        o342(.A(ori_ori_n315_), .B(ori_ori_n232_), .Y(ori_ori_n371_));
  INV        o343(.A(ori_ori_n261_), .Y(ori_ori_n372_));
  NA2        o344(.A(ori_ori_n372_), .B(ori_ori_n371_), .Y(ori_ori_n373_));
  INV        o345(.A(ori_ori_n343_), .Y(ori_ori_n374_));
  NO2        o346(.A(ori_ori_n374_), .B(m), .Y(ori_ori_n375_));
  NO2        o347(.A(ori_ori_n373_), .B(ori_ori_n375_), .Y(ori_ori_n376_));
  INV        o348(.A(j), .Y(ori_ori_n377_));
  NO3        o349(.A(ori_ori_n171_), .B(ori_ori_n377_), .C(ori_ori_n30_), .Y(ori_ori_n378_));
  AOI210     o350(.A0(ori_ori_n281_), .A1(n), .B0(ori_ori_n288_), .Y(ori_ori_n379_));
  NA2        o351(.A(ori_ori_n379_), .B(ori_ori_n291_), .Y(ori_ori_n380_));
  AN3        o352(.A(ori_ori_n380_), .B(ori_ori_n378_), .C(ori_ori_n62_), .Y(ori_ori_n381_));
  NA2        o353(.A(ori_ori_n309_), .B(ori_ori_n177_), .Y(ori_ori_n382_));
  INV        o354(.A(ori_ori_n382_), .Y(ori_ori_n383_));
  NO2        o355(.A(ori_ori_n171_), .B(ori_ori_n84_), .Y(ori_ori_n384_));
  AOI220     o356(.A0(ori_ori_n384_), .A1(ori_ori_n315_), .B0(ori_ori_n366_), .B1(ori_ori_n356_), .Y(ori_ori_n385_));
  INV        o357(.A(ori_ori_n59_), .Y(ori_ori_n386_));
  NA2        o358(.A(ori_ori_n386_), .B(ori_ori_n305_), .Y(ori_ori_n387_));
  NA2        o359(.A(ori_ori_n387_), .B(ori_ori_n385_), .Y(ori_ori_n388_));
  OR3        o360(.A(ori_ori_n388_), .B(ori_ori_n383_), .C(ori_ori_n381_), .Y(ori_ori_n389_));
  NA3        o361(.A(ori_ori_n379_), .B(ori_ori_n291_), .C(ori_ori_n290_), .Y(ori_ori_n390_));
  NA3        o362(.A(ori_ori_n390_), .B(ori_ori_n133_), .C(ori_ori_n29_), .Y(ori_ori_n391_));
  NO3        o363(.A(ori_ori_n255_), .B(ori_ori_n246_), .C(f), .Y(ori_ori_n392_));
  NO2        o364(.A(ori_ori_n60_), .B(ori_ori_n33_), .Y(ori_ori_n393_));
  NA2        o365(.A(ori_ori_n393_), .B(ori_ori_n321_), .Y(ori_ori_n394_));
  NA2        o366(.A(ori_ori_n394_), .B(ori_ori_n391_), .Y(ori_ori_n395_));
  NO2        o367(.A(ori_ori_n336_), .B(ori_ori_n44_), .Y(ori_ori_n396_));
  NA2        o368(.A(ori_ori_n392_), .B(ori_ori_n396_), .Y(ori_ori_n397_));
  NA3        o369(.A(ori_ori_n156_), .B(ori_ori_n41_), .C(b), .Y(ori_ori_n398_));
  INV        o370(.A(ori_ori_n397_), .Y(ori_ori_n399_));
  NO3        o371(.A(ori_ori_n399_), .B(ori_ori_n395_), .C(ori_ori_n389_), .Y(ori_ori_n400_));
  NO2        o372(.A(ori_ori_n200_), .B(ori_ori_n172_), .Y(ori_ori_n401_));
  NA2        o373(.A(ori_ori_n401_), .B(ori_ori_n380_), .Y(ori_ori_n402_));
  NO2        o374(.A(ori_ori_n278_), .B(h), .Y(ori_ori_n403_));
  NA2        o375(.A(ori_ori_n403_), .B(ori_ori_n353_), .Y(ori_ori_n404_));
  NA3        o376(.A(ori_ori_n404_), .B(ori_ori_n402_), .C(ori_ori_n237_), .Y(ori_ori_n405_));
  NO2        o377(.A(ori_ori_n289_), .B(ori_ori_n52_), .Y(ori_ori_n406_));
  NA2        o378(.A(ori_ori_n401_), .B(ori_ori_n406_), .Y(ori_ori_n407_));
  OAI210     o379(.A0(ori_ori_n357_), .A1(ori_ori_n233_), .B0(ori_ori_n407_), .Y(ori_ori_n408_));
  BUFFER     o380(.A(ori_ori_n384_), .Y(ori_ori_n409_));
  NA2        o381(.A(ori_ori_n409_), .B(ori_ori_n338_), .Y(ori_ori_n410_));
  INV        o382(.A(ori_ori_n410_), .Y(ori_ori_n411_));
  NO3        o383(.A(ori_ori_n411_), .B(ori_ori_n408_), .C(ori_ori_n405_), .Y(ori_ori_n412_));
  NA4        o384(.A(ori_ori_n412_), .B(ori_ori_n400_), .C(ori_ori_n376_), .D(ori_ori_n370_), .Y(ori09));
  NA3        o385(.A(m), .B(l), .C(i), .Y(ori_ori_n414_));
  NA2        o386(.A(ori_ori_n210_), .B(ori_ori_n414_), .Y(ori_ori_n415_));
  NO2        o387(.A(ori_ori_n78_), .B(ori_ori_n76_), .Y(ori_ori_n416_));
  NOi31      o388(.An(k), .B(m), .C(l), .Y(ori_ori_n417_));
  NO2        o389(.A(ori_ori_n199_), .B(ori_ori_n417_), .Y(ori_ori_n418_));
  AOI210     o390(.A0(ori_ori_n418_), .A1(ori_ori_n416_), .B0(ori_ori_n306_), .Y(ori_ori_n419_));
  NA2        o391(.A(ori_ori_n398_), .B(ori_ori_n192_), .Y(ori_ori_n420_));
  AOI220     o392(.A0(k), .A1(ori_ori_n420_), .B0(ori_ori_n419_), .B1(n), .Y(ori_ori_n421_));
  NA3        o393(.A(ori_ori_n421_), .B(ori_ori_n316_), .C(ori_ori_n50_), .Y(ori_ori_n422_));
  NO3        o394(.A(ori_ori_n81_), .B(ori_ori_n187_), .C(ori_ori_n95_), .Y(ori_ori_n423_));
  NO2        o395(.A(ori_ori_n330_), .B(ori_ori_n187_), .Y(ori_ori_n424_));
  INV        o396(.A(ori_ori_n423_), .Y(ori_ori_n425_));
  NA3        o397(.A(ori_ori_n99_), .B(ori_ori_n68_), .C(g), .Y(ori_ori_n426_));
  NO2        o398(.A(ori_ori_n198_), .B(ori_ori_n426_), .Y(ori_ori_n427_));
  NOi31      o399(.An(ori_ori_n137_), .B(ori_ori_n427_), .C(ori_ori_n175_), .Y(ori_ori_n428_));
  NA3        o400(.A(e), .B(ori_ori_n268_), .C(f), .Y(ori_ori_n429_));
  NA3        o401(.A(ori_ori_n429_), .B(ori_ori_n428_), .C(ori_ori_n425_), .Y(ori_ori_n430_));
  NO2        o402(.A(ori_ori_n430_), .B(ori_ori_n422_), .Y(ori_ori_n431_));
  NO2        o403(.A(ori_ori_n84_), .B(ori_ori_n81_), .Y(ori_ori_n432_));
  INV        o404(.A(ori_ori_n243_), .Y(ori_ori_n433_));
  NA2        o405(.A(ori_ori_n315_), .B(ori_ori_n205_), .Y(ori_ori_n434_));
  NA2        o406(.A(ori_ori_n434_), .B(ori_ori_n158_), .Y(ori_ori_n435_));
  NO2        o407(.A(ori_ori_n435_), .B(ori_ori_n432_), .Y(ori_ori_n436_));
  OAI210     o408(.A0(ori_ori_n172_), .A1(j), .B0(ori_ori_n42_), .Y(ori_ori_n437_));
  AOI220     o409(.A0(ori_ori_n437_), .A1(ori_ori_n424_), .B0(ori_ori_n307_), .B1(ori_ori_n314_), .Y(ori_ori_n438_));
  INV        o410(.A(ori_ori_n438_), .Y(ori_ori_n439_));
  AN2        o411(.A(ori_ori_n420_), .B(ori_ori_n415_), .Y(ori_ori_n440_));
  NO2        o412(.A(ori_ori_n440_), .B(ori_ori_n439_), .Y(ori_ori_n441_));
  AN2        o413(.A(ori_ori_n195_), .B(ori_ori_n441_), .Y(ori_ori_n442_));
  NA3        o414(.A(ori_ori_n442_), .B(ori_ori_n436_), .C(ori_ori_n431_), .Y(ori12));
  NO2        o415(.A(e), .B(c), .Y(ori_ori_n444_));
  NO4        o416(.A(ori_ori_n247_), .B(ori_ori_n157_), .C(ori_ori_n303_), .D(ori_ori_n131_), .Y(ori_ori_n445_));
  NO2        o417(.A(ori_ori_n335_), .B(ori_ori_n220_), .Y(ori_ori_n446_));
  AOI210     o418(.A0(ori_ori_n145_), .A1(ori_ori_n197_), .B0(ori_ori_n124_), .Y(ori_ori_n447_));
  NO2        o419(.A(ori_ori_n229_), .B(ori_ori_n131_), .Y(ori_ori_n448_));
  NA2        o420(.A(ori_ori_n448_), .B(f), .Y(ori_ori_n449_));
  INV        o421(.A(ori_ori_n94_), .Y(ori_ori_n450_));
  NA2        o422(.A(ori_ori_n450_), .B(ori_ori_n149_), .Y(ori_ori_n451_));
  NA2        o423(.A(ori_ori_n451_), .B(ori_ori_n449_), .Y(ori_ori_n452_));
  INV        o424(.A(ori_ori_n211_), .Y(ori_ori_n453_));
  NO3        o425(.A(ori_ori_n81_), .B(ori_ori_n95_), .C(ori_ori_n131_), .Y(ori_ori_n454_));
  NA2        o426(.A(ori_ori_n454_), .B(ori_ori_n281_), .Y(ori_ori_n455_));
  NA3        o427(.A(ori_ori_n248_), .B(d), .C(g), .Y(ori_ori_n456_));
  NA3        o428(.A(ori_ori_n456_), .B(ori_ori_n455_), .C(ori_ori_n453_), .Y(ori_ori_n457_));
  NO3        o429(.A(ori_ori_n457_), .B(ori_ori_n452_), .C(ori_ori_n445_), .Y(ori_ori_n458_));
  NA2        o430(.A(ori_ori_n289_), .B(ori_ori_n89_), .Y(ori_ori_n459_));
  NOi21      o431(.An(ori_ori_n29_), .B(ori_ori_n330_), .Y(ori_ori_n460_));
  NA2        o432(.A(ori_ori_n460_), .B(ori_ori_n459_), .Y(ori_ori_n461_));
  INV        o433(.A(ori_ori_n461_), .Y(ori_ori_n462_));
  INV        o434(.A(ori_ori_n185_), .Y(ori_ori_n463_));
  NO2        o435(.A(ori_ori_n264_), .B(ori_ori_n172_), .Y(ori_ori_n464_));
  NO2        o436(.A(ori_ori_n264_), .B(ori_ori_n89_), .Y(ori_ori_n465_));
  NO3        o437(.A(ori_ori_n465_), .B(ori_ori_n463_), .C(ori_ori_n462_), .Y(ori_ori_n466_));
  NA2        o438(.A(ori_ori_n205_), .B(g), .Y(ori_ori_n467_));
  NA2        o439(.A(ori_ori_n100_), .B(i), .Y(ori_ori_n468_));
  NA2        o440(.A(ori_ori_n32_), .B(i), .Y(ori_ori_n469_));
  NO2        o441(.A(ori_ori_n469_), .B(l), .Y(ori_ori_n470_));
  INV        o442(.A(ori_ori_n470_), .Y(ori_ori_n471_));
  NO2        o443(.A(ori_ori_n89_), .B(ori_ori_n52_), .Y(ori_ori_n472_));
  OR2        o444(.A(ori_ori_n472_), .B(ori_ori_n288_), .Y(ori_ori_n473_));
  NO2        o445(.A(ori_ori_n677_), .B(ori_ori_n473_), .Y(ori_ori_n474_));
  OAI220     o446(.A0(ori_ori_n474_), .A1(ori_ori_n467_), .B0(ori_ori_n471_), .B1(ori_ori_n192_), .Y(ori_ori_n475_));
  NO2        o447(.A(ori_ori_n251_), .B(ori_ori_n131_), .Y(ori_ori_n476_));
  AOI210     o448(.A0(ori_ori_n476_), .A1(ori_ori_n224_), .B0(ori_ori_n135_), .Y(ori_ori_n477_));
  AOI220     o449(.A0(ori_ori_n446_), .A1(ori_ori_n450_), .B0(ori_ori_n305_), .B1(ori_ori_n58_), .Y(ori_ori_n478_));
  NA2        o450(.A(ori_ori_n478_), .B(ori_ori_n477_), .Y(ori_ori_n479_));
  NA2        o451(.A(ori_ori_n323_), .B(ori_ori_n281_), .Y(ori_ori_n480_));
  INV        o452(.A(ori_ori_n480_), .Y(ori_ori_n481_));
  NO3        o453(.A(ori_ori_n481_), .B(ori_ori_n479_), .C(ori_ori_n475_), .Y(ori_ori_n482_));
  NAi31      o454(.An(c), .B(e), .C(n), .Y(ori_ori_n483_));
  NO3        o455(.A(ori_ori_n76_), .B(ori_ori_n199_), .C(ori_ori_n417_), .Y(ori_ori_n484_));
  NO2        o456(.A(ori_ori_n484_), .B(ori_ori_n483_), .Y(ori_ori_n485_));
  NO2        o457(.A(h), .B(c), .Y(ori_ori_n486_));
  AOI210     o458(.A0(ori_ori_n486_), .A1(ori_ori_n258_), .B0(ori_ori_n485_), .Y(ori_ori_n487_));
  INV        o459(.A(ori_ori_n487_), .Y(ori_ori_n488_));
  NO3        o460(.A(ori_ori_n177_), .B(ori_ori_n248_), .C(ori_ori_n105_), .Y(ori_ori_n489_));
  NOi31      o461(.An(e), .B(ori_ori_n489_), .C(ori_ori_n131_), .Y(ori_ori_n490_));
  NAi21      o462(.An(ori_ori_n289_), .B(ori_ori_n476_), .Y(ori_ori_n491_));
  INV        o463(.A(ori_ori_n491_), .Y(ori_ori_n492_));
  NA2        o464(.A(ori_ori_n447_), .B(ori_ori_n444_), .Y(ori_ori_n493_));
  NA2        o465(.A(ori_ori_n493_), .B(ori_ori_n313_), .Y(ori_ori_n494_));
  OR2        o466(.A(ori_ori_n191_), .B(ori_ori_n494_), .Y(ori_ori_n495_));
  NO4        o467(.A(ori_ori_n495_), .B(ori_ori_n492_), .C(ori_ori_n490_), .D(ori_ori_n488_), .Y(ori_ori_n496_));
  NA4        o468(.A(ori_ori_n496_), .B(ori_ori_n482_), .C(ori_ori_n466_), .D(ori_ori_n458_), .Y(ori13));
  NA2        o469(.A(d), .B(ori_ori_n73_), .Y(ori_ori_n498_));
  NAi32      o470(.An(f), .Bn(e), .C(c), .Y(ori_ori_n499_));
  NA3        o471(.A(k), .B(j), .C(i), .Y(ori_ori_n500_));
  NO2        o472(.A(f), .B(c), .Y(ori_ori_n501_));
  NOi21      o473(.An(ori_ori_n501_), .B(ori_ori_n247_), .Y(ori_ori_n502_));
  OR2        o474(.A(m), .B(i), .Y(ori_ori_n503_));
  AN3        o475(.A(g), .B(f), .C(c), .Y(ori_ori_n504_));
  NA3        o476(.A(l), .B(k), .C(j), .Y(ori_ori_n505_));
  NA2        o477(.A(i), .B(h), .Y(ori_ori_n506_));
  NO3        o478(.A(ori_ori_n506_), .B(ori_ori_n505_), .C(ori_ori_n81_), .Y(ori_ori_n507_));
  NO2        o479(.A(ori_ori_n169_), .B(ori_ori_n131_), .Y(ori_ori_n508_));
  NO2        o480(.A(ori_ori_n279_), .B(ori_ori_n306_), .Y(ori_ori_n509_));
  NA4        o481(.A(ori_ori_n56_), .B(ori_ori_n55_), .C(g), .D(ori_ori_n130_), .Y(ori_ori_n510_));
  NA4        o482(.A(ori_ori_n297_), .B(m), .C(ori_ori_n71_), .D(ori_ori_n130_), .Y(ori_ori_n511_));
  NA2        o483(.A(ori_ori_n511_), .B(ori_ori_n510_), .Y(ori_ori_n512_));
  NO2        o484(.A(ori_ori_n512_), .B(ori_ori_n509_), .Y(ori_ori_n513_));
  NO2        o485(.A(ori_ori_n513_), .B(ori_ori_n304_), .Y(ori_ori_n514_));
  NOi31      o486(.An(m), .B(n), .C(f), .Y(ori_ori_n515_));
  NA2        o487(.A(ori_ori_n515_), .B(ori_ori_n35_), .Y(ori_ori_n516_));
  INV        o488(.A(e), .Y(ori_ori_n517_));
  NO2        o489(.A(ori_ori_n517_), .B(ori_ori_n516_), .Y(ori_ori_n518_));
  NO2        o490(.A(ori_ori_n518_), .B(ori_ori_n514_), .Y(ori_ori_n519_));
  NA2        o491(.A(c), .B(b), .Y(ori_ori_n520_));
  NO2        o492(.A(ori_ori_n352_), .B(ori_ori_n520_), .Y(ori_ori_n521_));
  NAi21      o493(.An(ori_ori_n240_), .B(ori_ori_n521_), .Y(ori_ori_n522_));
  NA2        o494(.A(ori_ori_n522_), .B(ori_ori_n519_), .Y(ori00));
  NA2        o495(.A(ori_ori_n433_), .B(ori_ori_n450_), .Y(ori_ori_n524_));
  INV        o496(.A(ori_ori_n524_), .Y(ori_ori_n525_));
  NA2        o497(.A(ori_ori_n268_), .B(f), .Y(ori_ori_n526_));
  OAI210     o498(.A0(ori_ori_n484_), .A1(ori_ori_n30_), .B0(ori_ori_n324_), .Y(ori_ori_n527_));
  NA3        o499(.A(ori_ori_n527_), .B(ori_ori_n162_), .C(n), .Y(ori_ori_n528_));
  AOI210     o500(.A0(ori_ori_n528_), .A1(ori_ori_n526_), .B0(ori_ori_n498_), .Y(ori_ori_n529_));
  NO2        o501(.A(ori_ori_n529_), .B(ori_ori_n525_), .Y(ori_ori_n530_));
  NA3        o502(.A(d), .B(ori_ori_n38_), .C(b), .Y(ori_ori_n531_));
  NO4        o503(.A(ori_ori_n674_), .B(ori_ori_n212_), .C(ori_ori_n520_), .D(ori_ori_n41_), .Y(ori_ori_n532_));
  NA3        o504(.A(ori_ori_n225_), .B(ori_ori_n136_), .C(g), .Y(ori_ori_n533_));
  OR2        o505(.A(ori_ori_n533_), .B(ori_ori_n531_), .Y(ori_ori_n534_));
  NO2        o506(.A(h), .B(g), .Y(ori_ori_n535_));
  NA4        o507(.A(ori_ori_n258_), .B(d), .C(ori_ori_n535_), .D(b), .Y(ori_ori_n536_));
  NO2        o508(.A(ori_ori_n279_), .B(ori_ori_n306_), .Y(ori_ori_n537_));
  AOI220     o509(.A0(ori_ori_n537_), .A1(ori_ori_n284_), .B0(ori_ori_n454_), .B1(ori_ori_n298_), .Y(ori_ori_n538_));
  NA2        o510(.A(ori_ori_n182_), .B(ori_ori_n154_), .Y(ori_ori_n539_));
  NA4        o511(.A(ori_ori_n539_), .B(ori_ori_n538_), .C(ori_ori_n536_), .D(ori_ori_n534_), .Y(ori_ori_n540_));
  NO2        o512(.A(ori_ori_n540_), .B(ori_ori_n532_), .Y(ori_ori_n541_));
  NA2        o513(.A(ori_ori_n154_), .B(ori_ori_n205_), .Y(ori_ori_n542_));
  INV        o514(.A(ori_ori_n542_), .Y(ori_ori_n543_));
  NO2        o515(.A(ori_ori_n148_), .B(ori_ori_n110_), .Y(ori_ori_n544_));
  NO2        o516(.A(ori_ori_n544_), .B(ori_ori_n543_), .Y(ori_ori_n545_));
  AN3        o517(.A(ori_ori_n545_), .B(ori_ori_n541_), .C(ori_ori_n299_), .Y(ori_ori_n546_));
  NA3        o518(.A(ori_ori_n515_), .B(e), .C(ori_ori_n253_), .Y(ori_ori_n547_));
  INV        o519(.A(ori_ori_n547_), .Y(ori_ori_n548_));
  NA2        o520(.A(ori_ori_n512_), .B(ori_ori_n284_), .Y(ori_ori_n549_));
  NA3        o521(.A(ori_ori_n326_), .B(ori_ori_n136_), .C(ori_ori_n100_), .Y(ori_ori_n550_));
  NA2        o522(.A(ori_ori_n550_), .B(ori_ori_n549_), .Y(ori_ori_n551_));
  NA2        o523(.A(n), .B(e), .Y(ori_ori_n552_));
  NO2        o524(.A(ori_ori_n552_), .B(ori_ori_n91_), .Y(ori_ori_n553_));
  NA2        o525(.A(ori_ori_n553_), .B(ori_ori_n165_), .Y(ori_ori_n554_));
  INV        o526(.A(ori_ori_n554_), .Y(ori_ori_n555_));
  NA2        o527(.A(ori_ori_n553_), .B(ori_ori_n419_), .Y(ori_ori_n556_));
  AOI220     o528(.A0(ori_ori_n460_), .A1(ori_ori_n298_), .B0(ori_ori_n326_), .B1(ori_ori_n151_), .Y(ori_ori_n557_));
  NA2        o529(.A(ori_ori_n557_), .B(ori_ori_n556_), .Y(ori_ori_n558_));
  NO4        o530(.A(ori_ori_n558_), .B(ori_ori_n555_), .C(ori_ori_n551_), .D(ori_ori_n548_), .Y(ori_ori_n559_));
  NA3        o531(.A(ori_ori_n559_), .B(ori_ori_n546_), .C(ori_ori_n530_), .Y(ori01));
  NO2        o532(.A(ori_ori_n254_), .B(ori_ori_n168_), .Y(ori_ori_n561_));
  INV        o533(.A(ori_ori_n234_), .Y(ori_ori_n562_));
  NA3        o534(.A(ori_ori_n562_), .B(ori_ori_n561_), .C(ori_ori_n493_), .Y(ori_ori_n563_));
  NA2        o535(.A(ori_ori_n305_), .B(ori_ori_n58_), .Y(ori_ori_n564_));
  NA2        o536(.A(ori_ori_n289_), .B(ori_ori_n164_), .Y(ori_ori_n565_));
  NA2        o537(.A(ori_ori_n464_), .B(ori_ori_n565_), .Y(ori_ori_n566_));
  NA4        o538(.A(ori_ori_n566_), .B(ori_ori_n564_), .C(ori_ori_n438_), .D(ori_ori_n193_), .Y(ori_ori_n567_));
  INV        o539(.A(ori_ori_n85_), .Y(ori_ori_n568_));
  NO3        o540(.A(ori_ori_n568_), .B(ori_ori_n567_), .C(ori_ori_n563_), .Y(ori_ori_n569_));
  INV        o541(.A(ori_ori_n533_), .Y(ori_ori_n570_));
  NA2        o542(.A(ori_ori_n570_), .B(ori_ori_n281_), .Y(ori_ori_n571_));
  OAI210     o543(.A0(ori_ori_n214_), .A1(ori_ori_n29_), .B0(m), .Y(ori_ori_n572_));
  OR2        o544(.A(ori_ori_n572_), .B(ori_ori_n192_), .Y(ori_ori_n573_));
  NA2        o545(.A(ori_ori_n573_), .B(ori_ori_n571_), .Y(ori_ori_n574_));
  NA2        o546(.A(ori_ori_n167_), .B(ori_ori_n119_), .Y(ori_ori_n575_));
  NA2        o547(.A(ori_ori_n575_), .B(ori_ori_n338_), .Y(ori_ori_n576_));
  NA2        o548(.A(ori_ori_n576_), .B(ori_ori_n394_), .Y(ori_ori_n577_));
  NO2        o549(.A(ori_ori_n577_), .B(ori_ori_n574_), .Y(ori_ori_n578_));
  NA2        o550(.A(ori_ori_n265_), .B(ori_ori_n40_), .Y(ori_ori_n579_));
  NO2        o551(.A(ori_ori_n128_), .B(ori_ori_n70_), .Y(ori_ori_n580_));
  INV        o552(.A(ori_ori_n580_), .Y(ori_ori_n581_));
  NA2        o553(.A(ori_ori_n581_), .B(ori_ori_n579_), .Y(ori_ori_n582_));
  INV        o554(.A(ori_ori_n468_), .Y(ori_ori_n583_));
  NO2        o555(.A(ori_ori_n469_), .B(ori_ori_n291_), .Y(ori_ori_n584_));
  OAI210     o556(.A0(ori_ori_n584_), .A1(ori_ori_n583_), .B0(ori_ori_n199_), .Y(ori_ori_n585_));
  NO3        o557(.A(ori_ori_n49_), .B(ori_ori_n172_), .C(ori_ori_n31_), .Y(ori_ori_n586_));
  NA2        o558(.A(ori_ori_n586_), .B(ori_ori_n288_), .Y(ori_ori_n587_));
  INV        o559(.A(ori_ori_n587_), .Y(ori_ori_n588_));
  OR2        o560(.A(ori_ori_n533_), .B(ori_ori_n531_), .Y(ori_ori_n589_));
  NA2        o561(.A(ori_ori_n586_), .B(ori_ori_n406_), .Y(ori_ori_n590_));
  NA2        o562(.A(ori_ori_n590_), .B(ori_ori_n589_), .Y(ori_ori_n591_));
  NOi41      o563(.An(ori_ori_n585_), .B(ori_ori_n591_), .C(ori_ori_n588_), .D(ori_ori_n582_), .Y(ori_ori_n592_));
  NO2        o564(.A(g), .B(ori_ori_n31_), .Y(ori_ori_n593_));
  AO220      o565(.A0(i), .A1(ori_ori_n315_), .B0(ori_ori_n593_), .B1(ori_ori_n356_), .Y(ori_ori_n594_));
  NA2        o566(.A(ori_ori_n594_), .B(ori_ori_n199_), .Y(ori_ori_n595_));
  NO2        o567(.A(ori_ori_n506_), .B(ori_ori_n106_), .Y(ori_ori_n596_));
  NA2        o568(.A(ori_ori_n586_), .B(ori_ori_n472_), .Y(ori_ori_n597_));
  NA2        o569(.A(ori_ori_n597_), .B(ori_ori_n595_), .Y(ori_ori_n598_));
  NO2        o570(.A(ori_ori_n309_), .B(ori_ori_n308_), .Y(ori_ori_n599_));
  NO4        o571(.A(ori_ori_n506_), .B(ori_ori_n599_), .C(ori_ori_n104_), .D(ori_ori_n55_), .Y(ori_ori_n600_));
  NO2        o572(.A(ori_ori_n600_), .B(ori_ori_n598_), .Y(ori_ori_n601_));
  NA4        o573(.A(ori_ori_n601_), .B(ori_ori_n592_), .C(ori_ori_n578_), .D(ori_ori_n569_), .Y(ori06));
  NO2        o574(.A(ori_ori_n138_), .B(ori_ori_n63_), .Y(ori_ori_n603_));
  OAI210     o575(.A0(ori_ori_n603_), .A1(ori_ori_n596_), .B0(ori_ori_n224_), .Y(ori_ori_n604_));
  NA2        o576(.A(ori_ori_n604_), .B(ori_ori_n585_), .Y(ori_ori_n605_));
  NO3        o577(.A(ori_ori_n605_), .B(ori_ori_n588_), .C(ori_ori_n161_), .Y(ori_ori_n606_));
  NA2        o578(.A(i), .B(ori_ori_n473_), .Y(ori_ori_n607_));
  AOI210     o579(.A0(i), .A1(ori_ori_n292_), .B0(ori_ori_n594_), .Y(ori_ori_n608_));
  AOI210     o580(.A0(ori_ori_n608_), .A1(ori_ori_n607_), .B0(ori_ori_n197_), .Y(ori_ori_n609_));
  NA2        o581(.A(ori_ori_n56_), .B(ori_ori_n321_), .Y(ori_ori_n610_));
  NA2        o582(.A(ori_ori_n155_), .B(ori_ori_n610_), .Y(ori_ori_n611_));
  NO3        o583(.A(ori_ori_n460_), .B(ori_ori_n611_), .C(ori_ori_n609_), .Y(ori_ori_n612_));
  NO2        o584(.A(n), .B(ori_ori_n33_), .Y(ori_ori_n613_));
  NA2        o585(.A(ori_ori_n215_), .B(ori_ori_n613_), .Y(ori_ori_n614_));
  INV        o586(.A(k), .Y(ori_ori_n615_));
  NO3        o587(.A(ori_ori_n615_), .B(ori_ori_n306_), .C(j), .Y(ori_ori_n616_));
  INV        o588(.A(ori_ori_n518_), .Y(ori_ori_n617_));
  NA3        o589(.A(ori_ori_n617_), .B(ori_ori_n614_), .C(ori_ori_n557_), .Y(ori_ori_n618_));
  NA2        o590(.A(ori_ori_n616_), .B(ori_ori_n396_), .Y(ori_ori_n619_));
  INV        o591(.A(ori_ori_n619_), .Y(ori_ori_n620_));
  INV        o592(.A(ori_ori_n261_), .Y(ori_ori_n621_));
  NA2        o593(.A(ori_ori_n621_), .B(ori_ori_n590_), .Y(ori_ori_n622_));
  NAi21      o594(.An(j), .B(i), .Y(ori_ori_n623_));
  NO4        o595(.A(ori_ori_n599_), .B(ori_ori_n623_), .C(ori_ori_n247_), .D(ori_ori_n146_), .Y(ori_ori_n624_));
  NO4        o596(.A(ori_ori_n624_), .B(ori_ori_n622_), .C(ori_ori_n620_), .D(ori_ori_n618_), .Y(ori_ori_n625_));
  NA4        o597(.A(ori_ori_n625_), .B(ori_ori_n612_), .C(ori_ori_n606_), .D(ori_ori_n601_), .Y(ori07));
  NOi31      o598(.An(n), .B(m), .C(b), .Y(ori_ori_n627_));
  NO3        o599(.A(ori_ori_n81_), .B(ori_ori_n249_), .C(h), .Y(ori_ori_n628_));
  NO2        o600(.A(m), .B(h), .Y(ori_ori_n629_));
  NO2        o601(.A(ori_ori_n499_), .B(ori_ori_n247_), .Y(ori_ori_n630_));
  NO2        o602(.A(ori_ori_n500_), .B(ori_ori_n176_), .Y(ori_ori_n631_));
  INV        o603(.A(ori_ori_n630_), .Y(ori_ori_n632_));
  NO2        o604(.A(l), .B(k), .Y(ori_ori_n633_));
  NO3        o605(.A(ori_ori_n247_), .B(d), .C(c), .Y(ori_ori_n634_));
  NA2        o606(.A(ori_ori_n504_), .B(d), .Y(ori_ori_n635_));
  NO2        o607(.A(ori_ori_n635_), .B(ori_ori_n247_), .Y(ori_ori_n636_));
  INV        o608(.A(ori_ori_n636_), .Y(ori_ori_n637_));
  NA2        o609(.A(ori_ori_n627_), .B(ori_ori_n221_), .Y(ori_ori_n638_));
  INV        o610(.A(ori_ori_n638_), .Y(ori_ori_n639_));
  INV        o611(.A(ori_ori_n507_), .Y(ori_ori_n640_));
  NAi21      o612(.An(ori_ori_n639_), .B(ori_ori_n640_), .Y(ori_ori_n641_));
  NA2        o613(.A(ori_ori_n629_), .B(ori_ori_n633_), .Y(ori_ori_n642_));
  NO2        o614(.A(ori_ori_n675_), .B(ori_ori_n641_), .Y(ori_ori_n643_));
  NA3        o615(.A(ori_ori_n643_), .B(ori_ori_n637_), .C(ori_ori_n632_), .Y(ori_ori_n644_));
  NO2        o616(.A(ori_ori_n231_), .B(j), .Y(ori_ori_n645_));
  NA2        o617(.A(ori_ori_n502_), .B(ori_ori_n93_), .Y(ori_ori_n646_));
  INV        o618(.A(ori_ori_n646_), .Y(ori_ori_n647_));
  NA2        o619(.A(ori_ori_n645_), .B(ori_ori_n98_), .Y(ori_ori_n648_));
  INV        o620(.A(ori_ori_n648_), .Y(ori_ori_n649_));
  NO2        o621(.A(ori_ori_n649_), .B(ori_ori_n647_), .Y(ori_ori_n650_));
  NO2        o622(.A(ori_ori_n138_), .B(ori_ori_n106_), .Y(ori_ori_n651_));
  NO2        o623(.A(ori_ori_n503_), .B(h), .Y(ori_ori_n652_));
  NO2        o624(.A(ori_ori_n623_), .B(ori_ori_n104_), .Y(ori_ori_n653_));
  NA2        o625(.A(h), .B(ori_ori_n653_), .Y(ori_ori_n654_));
  INV        o626(.A(ori_ori_n654_), .Y(ori_ori_n655_));
  NO3        o627(.A(ori_ori_n655_), .B(ori_ori_n72_), .C(ori_ori_n652_), .Y(ori_ori_n656_));
  NA3        o628(.A(ori_ori_n656_), .B(ori_ori_n676_), .C(ori_ori_n650_), .Y(ori_ori_n657_));
  NA2        o629(.A(h), .B(ori_ori_n631_), .Y(ori_ori_n658_));
  NO2        o630(.A(f), .B(e), .Y(ori_ori_n659_));
  NA2        o631(.A(ori_ori_n659_), .B(ori_ori_n238_), .Y(ori_ori_n660_));
  BUFFER     o632(.A(ori_ori_n81_), .Y(ori_ori_n661_));
  NO2        o633(.A(ori_ori_n661_), .B(ori_ori_n660_), .Y(ori_ori_n662_));
  INV        o634(.A(ori_ori_n662_), .Y(ori_ori_n663_));
  OR2        o635(.A(h), .B(ori_ori_n285_), .Y(ori_ori_n664_));
  NO2        o636(.A(ori_ori_n664_), .B(ori_ori_n104_), .Y(ori_ori_n665_));
  NA2        o637(.A(ori_ori_n508_), .B(ori_ori_n136_), .Y(ori_ori_n666_));
  INV        o638(.A(ori_ori_n666_), .Y(ori_ori_n667_));
  NO3        o639(.A(ori_ori_n667_), .B(ori_ori_n665_), .C(ori_ori_n634_), .Y(ori_ori_n668_));
  NA3        o640(.A(ori_ori_n668_), .B(ori_ori_n663_), .C(ori_ori_n658_), .Y(ori_ori_n669_));
  OR4        o641(.A(ori_ori_n628_), .B(ori_ori_n669_), .C(ori_ori_n657_), .D(ori_ori_n644_), .Y(ori04));
  INV        o642(.A(ori_ori_n77_), .Y(ori_ori_n673_));
  INV        o643(.A(ori_ori_n136_), .Y(ori_ori_n674_));
  INV        o644(.A(ori_ori_n642_), .Y(ori_ori_n675_));
  INV        o645(.A(ori_ori_n651_), .Y(ori_ori_n676_));
  INV        o646(.A(b), .Y(ori_ori_n677_));
  ZERO       o647(.Y(ori02));
  ZERO       o648(.Y(ori03));
  ZERO       o649(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA2        m0003(.A(mai_mai_n30_), .B(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  AN2        m0006(.A(m), .B(l), .Y(mai_mai_n35_));
  NOi32      m0007(.An(j), .Bn(g), .C(k), .Y(mai_mai_n36_));
  NA2        m0008(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n37_));
  NO2        m0009(.A(mai_mai_n37_), .B(n), .Y(mai_mai_n38_));
  NAi21      m0010(.An(j), .B(l), .Y(mai_mai_n39_));
  NAi32      m0011(.An(n), .Bn(g), .C(m), .Y(mai_mai_n40_));
  NO2        m0012(.A(mai_mai_n40_), .B(mai_mai_n39_), .Y(mai_mai_n41_));
  NAi31      m0013(.An(n), .B(m), .C(l), .Y(mai_mai_n42_));
  INV        m0014(.A(i), .Y(mai_mai_n43_));
  AN2        m0015(.A(h), .B(g), .Y(mai_mai_n44_));
  INV        m0016(.A(mai_mai_n42_), .Y(mai_mai_n45_));
  NAi21      m0017(.An(n), .B(m), .Y(mai_mai_n46_));
  NOi32      m0018(.An(k), .Bn(h), .C(g), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n46_), .B(mai_mai_n32_), .Y(mai_mai_n48_));
  INV        m0020(.A(c), .Y(mai_mai_n49_));
  NA2        m0021(.A(e), .B(b), .Y(mai_mai_n50_));
  INV        m0022(.A(d), .Y(mai_mai_n51_));
  NAi21      m0023(.An(i), .B(h), .Y(mai_mai_n52_));
  NAi31      m0024(.An(i), .B(l), .C(j), .Y(mai_mai_n53_));
  OAI220     m0025(.A0(mai_mai_n53_), .A1(mai_mai_n46_), .B0(mai_mai_n52_), .B1(mai_mai_n42_), .Y(mai_mai_n54_));
  NAi31      m0026(.An(d), .B(mai_mai_n54_), .C(c), .Y(mai_mai_n55_));
  NAi41      m0027(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n56_));
  NA2        m0028(.A(g), .B(f), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  NAi21      m0030(.An(i), .B(j), .Y(mai_mai_n59_));
  NAi32      m0031(.An(n), .Bn(k), .C(m), .Y(mai_mai_n60_));
  NAi31      m0032(.An(l), .B(m), .C(k), .Y(mai_mai_n61_));
  NAi41      m0033(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n62_));
  INV        m0034(.A(m), .Y(mai_mai_n63_));
  NOi21      m0035(.An(k), .B(l), .Y(mai_mai_n64_));
  AN4        m0036(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n65_));
  NOi31      m0037(.An(h), .B(g), .C(f), .Y(mai_mai_n66_));
  NA2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NOi32      m0039(.An(h), .Bn(g), .C(f), .Y(mai_mai_n68_));
  INV        m0040(.A(mai_mai_n55_), .Y(mai_mai_n69_));
  INV        m0041(.A(n), .Y(mai_mai_n70_));
  NOi32      m0042(.An(e), .Bn(b), .C(d), .Y(mai_mai_n71_));
  INV        m0043(.A(j), .Y(mai_mai_n72_));
  AN3        m0044(.A(m), .B(k), .C(i), .Y(mai_mai_n73_));
  NA3        m0045(.A(mai_mai_n73_), .B(mai_mai_n72_), .C(g), .Y(mai_mai_n74_));
  NAi32      m0046(.An(g), .Bn(f), .C(h), .Y(mai_mai_n75_));
  NAi31      m0047(.An(j), .B(m), .C(l), .Y(mai_mai_n76_));
  NO2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  NA2        m0049(.A(m), .B(l), .Y(mai_mai_n78_));
  NAi31      m0050(.An(k), .B(j), .C(g), .Y(mai_mai_n79_));
  NO3        m0051(.A(mai_mai_n79_), .B(mai_mai_n78_), .C(f), .Y(mai_mai_n80_));
  NOi32      m0052(.An(m), .Bn(l), .C(i), .Y(mai_mai_n81_));
  NOi21      m0053(.An(g), .B(i), .Y(mai_mai_n82_));
  NOi32      m0054(.An(m), .Bn(j), .C(k), .Y(mai_mai_n83_));
  AOI220     m0055(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n81_), .B1(j), .Y(mai_mai_n84_));
  NO2        m0056(.A(mai_mai_n84_), .B(f), .Y(mai_mai_n85_));
  NAi41      m0057(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n86_));
  AN2        m0058(.A(e), .B(b), .Y(mai_mai_n87_));
  NOi31      m0059(.An(c), .B(h), .C(f), .Y(mai_mai_n88_));
  NA2        m0060(.A(mai_mai_n88_), .B(mai_mai_n87_), .Y(mai_mai_n89_));
  NOi21      m0061(.An(g), .B(f), .Y(mai_mai_n90_));
  NOi21      m0062(.An(i), .B(h), .Y(mai_mai_n91_));
  NA3        m0063(.A(mai_mai_n91_), .B(mai_mai_n90_), .C(mai_mai_n35_), .Y(mai_mai_n92_));
  INV        m0064(.A(a), .Y(mai_mai_n93_));
  NA2        m0065(.A(mai_mai_n87_), .B(mai_mai_n93_), .Y(mai_mai_n94_));
  INV        m0066(.A(l), .Y(mai_mai_n95_));
  NOi21      m0067(.An(m), .B(n), .Y(mai_mai_n96_));
  AN2        m0068(.A(k), .B(h), .Y(mai_mai_n97_));
  INV        m0069(.A(b), .Y(mai_mai_n98_));
  NA2        m0070(.A(l), .B(j), .Y(mai_mai_n99_));
  AN2        m0071(.A(k), .B(i), .Y(mai_mai_n100_));
  NA2        m0072(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  NOi32      m0073(.An(c), .Bn(a), .C(d), .Y(mai_mai_n102_));
  NA2        m0074(.A(mai_mai_n102_), .B(mai_mai_n96_), .Y(mai_mai_n103_));
  NO2        m0075(.A(mai_mai_n103_), .B(mai_mai_n101_), .Y(mai_mai_n104_));
  NOi31      m0076(.An(k), .B(m), .C(j), .Y(mai_mai_n105_));
  NOi31      m0077(.An(k), .B(m), .C(i), .Y(mai_mai_n106_));
  NA3        m0078(.A(mai_mai_n106_), .B(mai_mai_n68_), .C(mai_mai_n65_), .Y(mai_mai_n107_));
  INV        m0079(.A(mai_mai_n107_), .Y(mai_mai_n108_));
  NOi32      m0080(.An(f), .Bn(b), .C(e), .Y(mai_mai_n109_));
  NAi21      m0081(.An(g), .B(h), .Y(mai_mai_n110_));
  NAi21      m0082(.An(m), .B(n), .Y(mai_mai_n111_));
  NAi21      m0083(.An(j), .B(k), .Y(mai_mai_n112_));
  NAi41      m0084(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n113_));
  NAi31      m0085(.An(j), .B(k), .C(h), .Y(mai_mai_n114_));
  NO3        m0086(.A(mai_mai_n114_), .B(mai_mai_n113_), .C(mai_mai_n111_), .Y(mai_mai_n115_));
  INV        m0087(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  NO2        m0088(.A(k), .B(j), .Y(mai_mai_n117_));
  AN2        m0089(.A(k), .B(j), .Y(mai_mai_n118_));
  NAi21      m0090(.An(c), .B(b), .Y(mai_mai_n119_));
  NA2        m0091(.A(f), .B(d), .Y(mai_mai_n120_));
  NA2        m0092(.A(h), .B(c), .Y(mai_mai_n121_));
  NA2        m0093(.A(d), .B(b), .Y(mai_mai_n122_));
  NAi21      m0094(.An(e), .B(f), .Y(mai_mai_n123_));
  NO2        m0095(.A(mai_mai_n123_), .B(mai_mai_n122_), .Y(mai_mai_n124_));
  NA2        m0096(.A(b), .B(a), .Y(mai_mai_n125_));
  NAi21      m0097(.An(c), .B(d), .Y(mai_mai_n126_));
  NAi31      m0098(.An(l), .B(k), .C(h), .Y(mai_mai_n127_));
  NO2        m0099(.A(mai_mai_n111_), .B(mai_mai_n127_), .Y(mai_mai_n128_));
  NA2        m0100(.A(mai_mai_n128_), .B(mai_mai_n124_), .Y(mai_mai_n129_));
  NAi31      m0101(.An(mai_mai_n108_), .B(mai_mai_n129_), .C(mai_mai_n116_), .Y(mai_mai_n130_));
  NAi31      m0102(.An(e), .B(f), .C(b), .Y(mai_mai_n131_));
  INV        m0103(.A(mai_mai_n131_), .Y(mai_mai_n132_));
  NOi21      m0104(.An(h), .B(i), .Y(mai_mai_n133_));
  NOi21      m0105(.An(k), .B(m), .Y(mai_mai_n134_));
  NA3        m0106(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(n), .Y(mai_mai_n135_));
  NOi21      m0107(.An(mai_mai_n132_), .B(mai_mai_n135_), .Y(mai_mai_n136_));
  NOi21      m0108(.An(h), .B(g), .Y(mai_mai_n137_));
  NO2        m0109(.A(mai_mai_n120_), .B(mai_mai_n119_), .Y(mai_mai_n138_));
  NA2        m0110(.A(mai_mai_n138_), .B(mai_mai_n137_), .Y(mai_mai_n139_));
  NAi31      m0111(.An(l), .B(j), .C(h), .Y(mai_mai_n140_));
  INV        m0112(.A(mai_mai_n46_), .Y(mai_mai_n141_));
  NA2        m0113(.A(mai_mai_n141_), .B(mai_mai_n58_), .Y(mai_mai_n142_));
  NOi32      m0114(.An(n), .Bn(k), .C(m), .Y(mai_mai_n143_));
  NA2        m0115(.A(l), .B(i), .Y(mai_mai_n144_));
  NA2        m0116(.A(mai_mai_n144_), .B(mai_mai_n143_), .Y(mai_mai_n145_));
  OAI210     m0117(.A0(mai_mai_n145_), .A1(mai_mai_n139_), .B0(mai_mai_n142_), .Y(mai_mai_n146_));
  NAi31      m0118(.An(d), .B(f), .C(c), .Y(mai_mai_n147_));
  NAi31      m0119(.An(e), .B(f), .C(c), .Y(mai_mai_n148_));
  NA2        m0120(.A(mai_mai_n148_), .B(mai_mai_n147_), .Y(mai_mai_n149_));
  NA2        m0121(.A(j), .B(h), .Y(mai_mai_n150_));
  OR3        m0122(.A(n), .B(m), .C(k), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n151_), .B(mai_mai_n150_), .Y(mai_mai_n152_));
  NAi32      m0124(.An(m), .Bn(k), .C(n), .Y(mai_mai_n153_));
  NO2        m0125(.A(mai_mai_n153_), .B(mai_mai_n150_), .Y(mai_mai_n154_));
  AOI220     m0126(.A0(mai_mai_n154_), .A1(mai_mai_n132_), .B0(mai_mai_n152_), .B1(mai_mai_n149_), .Y(mai_mai_n155_));
  NO2        m0127(.A(n), .B(m), .Y(mai_mai_n156_));
  NAi21      m0128(.An(f), .B(e), .Y(mai_mai_n157_));
  NA2        m0129(.A(d), .B(c), .Y(mai_mai_n158_));
  NAi31      m0130(.An(m), .B(n), .C(b), .Y(mai_mai_n159_));
  NA2        m0131(.A(k), .B(i), .Y(mai_mai_n160_));
  NAi21      m0132(.An(h), .B(f), .Y(mai_mai_n161_));
  NO2        m0133(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n159_), .B(mai_mai_n126_), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  NOi32      m0136(.An(f), .Bn(c), .C(d), .Y(mai_mai_n165_));
  NOi32      m0137(.An(f), .Bn(c), .C(e), .Y(mai_mai_n166_));
  NO2        m0138(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  NO3        m0139(.A(n), .B(m), .C(j), .Y(mai_mai_n168_));
  NA2        m0140(.A(mai_mai_n168_), .B(mai_mai_n97_), .Y(mai_mai_n169_));
  OR2        m0141(.A(mai_mai_n169_), .B(mai_mai_n167_), .Y(mai_mai_n170_));
  NA3        m0142(.A(mai_mai_n170_), .B(mai_mai_n164_), .C(mai_mai_n155_), .Y(mai_mai_n171_));
  OR4        m0143(.A(mai_mai_n171_), .B(mai_mai_n146_), .C(mai_mai_n136_), .D(mai_mai_n130_), .Y(mai_mai_n172_));
  NO4        m0144(.A(mai_mai_n172_), .B(mai_mai_n104_), .C(mai_mai_n69_), .D(mai_mai_n48_), .Y(mai_mai_n173_));
  NA3        m0145(.A(m), .B(mai_mai_n95_), .C(j), .Y(mai_mai_n174_));
  NAi31      m0146(.An(n), .B(h), .C(g), .Y(mai_mai_n175_));
  NO2        m0147(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  NOi32      m0148(.An(m), .Bn(k), .C(l), .Y(mai_mai_n177_));
  NA3        m0149(.A(mai_mai_n177_), .B(mai_mai_n72_), .C(g), .Y(mai_mai_n178_));
  NA4        m0150(.A(k), .B(mai_mai_n96_), .C(i), .D(g), .Y(mai_mai_n179_));
  AN2        m0151(.A(i), .B(g), .Y(mai_mai_n180_));
  NAi41      m0152(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n181_));
  INV        m0153(.A(mai_mai_n181_), .Y(mai_mai_n182_));
  INV        m0154(.A(f), .Y(mai_mai_n183_));
  INV        m0155(.A(g), .Y(mai_mai_n184_));
  NOi31      m0156(.An(i), .B(j), .C(h), .Y(mai_mai_n185_));
  NOi21      m0157(.An(l), .B(m), .Y(mai_mai_n186_));
  NA2        m0158(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  NO2        m0159(.A(mai_mai_n187_), .B(mai_mai_n184_), .Y(mai_mai_n188_));
  NA2        m0160(.A(mai_mai_n188_), .B(mai_mai_n182_), .Y(mai_mai_n189_));
  INV        m0161(.A(mai_mai_n189_), .Y(mai_mai_n190_));
  NOi21      m0162(.An(n), .B(m), .Y(mai_mai_n191_));
  NOi32      m0163(.An(l), .Bn(i), .C(j), .Y(mai_mai_n192_));
  NA2        m0164(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  OA220      m0165(.A0(mai_mai_n193_), .A1(mai_mai_n89_), .B0(m), .B1(mai_mai_n67_), .Y(mai_mai_n194_));
  NAi21      m0166(.An(j), .B(h), .Y(mai_mai_n195_));
  XN2        m0167(.A(i), .B(h), .Y(mai_mai_n196_));
  NA2        m0168(.A(mai_mai_n196_), .B(mai_mai_n195_), .Y(mai_mai_n197_));
  NOi31      m0169(.An(k), .B(n), .C(m), .Y(mai_mai_n198_));
  NOi31      m0170(.An(mai_mai_n198_), .B(mai_mai_n158_), .C(mai_mai_n157_), .Y(mai_mai_n199_));
  NA2        m0171(.A(mai_mai_n199_), .B(mai_mai_n197_), .Y(mai_mai_n200_));
  NAi31      m0172(.An(f), .B(e), .C(c), .Y(mai_mai_n201_));
  NA3        m0173(.A(e), .B(c), .C(b), .Y(mai_mai_n202_));
  NAi32      m0174(.An(m), .Bn(i), .C(k), .Y(mai_mai_n203_));
  NAi21      m0175(.An(n), .B(a), .Y(mai_mai_n204_));
  NO2        m0176(.A(mai_mai_n204_), .B(mai_mai_n122_), .Y(mai_mai_n205_));
  NAi41      m0177(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n206_));
  NO2        m0178(.A(mai_mai_n206_), .B(e), .Y(mai_mai_n207_));
  NA2        m0179(.A(mai_mai_n207_), .B(mai_mai_n205_), .Y(mai_mai_n208_));
  AN3        m0180(.A(mai_mai_n208_), .B(mai_mai_n200_), .C(mai_mai_n194_), .Y(mai_mai_n209_));
  OR2        m0181(.A(h), .B(g), .Y(mai_mai_n210_));
  NO2        m0182(.A(mai_mai_n210_), .B(mai_mai_n86_), .Y(mai_mai_n211_));
  NA2        m0183(.A(mai_mai_n211_), .B(mai_mai_n109_), .Y(mai_mai_n212_));
  NAi41      m0184(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n213_));
  NO2        m0185(.A(mai_mai_n213_), .B(mai_mai_n183_), .Y(mai_mai_n214_));
  NA2        m0186(.A(mai_mai_n134_), .B(mai_mai_n91_), .Y(mai_mai_n215_));
  NAi21      m0187(.An(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n216_));
  NO2        m0188(.A(n), .B(a), .Y(mai_mai_n217_));
  NAi31      m0189(.An(mai_mai_n206_), .B(mai_mai_n217_), .C(mai_mai_n87_), .Y(mai_mai_n218_));
  AN2        m0190(.A(mai_mai_n218_), .B(mai_mai_n216_), .Y(mai_mai_n219_));
  NAi21      m0191(.An(h), .B(i), .Y(mai_mai_n220_));
  NA2        m0192(.A(mai_mai_n156_), .B(k), .Y(mai_mai_n221_));
  NO2        m0193(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  NA2        m0194(.A(mai_mai_n222_), .B(mai_mai_n165_), .Y(mai_mai_n223_));
  NA3        m0195(.A(mai_mai_n223_), .B(mai_mai_n219_), .C(mai_mai_n212_), .Y(mai_mai_n224_));
  NOi21      m0196(.An(g), .B(e), .Y(mai_mai_n225_));
  NO2        m0197(.A(mai_mai_n62_), .B(mai_mai_n63_), .Y(mai_mai_n226_));
  NA2        m0198(.A(mai_mai_n226_), .B(mai_mai_n225_), .Y(mai_mai_n227_));
  NOi32      m0199(.An(l), .Bn(j), .C(i), .Y(mai_mai_n228_));
  AOI210     m0200(.A0(mai_mai_n64_), .A1(mai_mai_n72_), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  NAi21      m0201(.An(f), .B(g), .Y(mai_mai_n230_));
  NO2        m0202(.A(mai_mai_n230_), .B(mai_mai_n56_), .Y(mai_mai_n231_));
  NO2        m0203(.A(mai_mai_n60_), .B(mai_mai_n99_), .Y(mai_mai_n232_));
  NA2        m0204(.A(mai_mai_n232_), .B(mai_mai_n231_), .Y(mai_mai_n233_));
  OAI210     m0205(.A0(mai_mai_n229_), .A1(mai_mai_n227_), .B0(mai_mai_n233_), .Y(mai_mai_n234_));
  NOi41      m0206(.An(mai_mai_n209_), .B(mai_mai_n234_), .C(mai_mai_n224_), .D(mai_mai_n190_), .Y(mai_mai_n235_));
  NO2        m0207(.A(mai_mai_n176_), .B(mai_mai_n45_), .Y(mai_mai_n236_));
  NO2        m0208(.A(mai_mai_n236_), .B(mai_mai_n94_), .Y(mai_mai_n237_));
  NAi21      m0209(.An(h), .B(g), .Y(mai_mai_n238_));
  OR3        m0210(.A(mai_mai_n1232_), .B(mai_mai_n193_), .C(e), .Y(mai_mai_n239_));
  NAi31      m0211(.An(g), .B(k), .C(h), .Y(mai_mai_n240_));
  NO3        m0212(.A(mai_mai_n111_), .B(mai_mai_n240_), .C(l), .Y(mai_mai_n241_));
  NAi31      m0213(.An(e), .B(d), .C(a), .Y(mai_mai_n242_));
  NA2        m0214(.A(mai_mai_n241_), .B(mai_mai_n109_), .Y(mai_mai_n243_));
  NA2        m0215(.A(mai_mai_n243_), .B(mai_mai_n239_), .Y(mai_mai_n244_));
  NA3        m0216(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n70_), .Y(mai_mai_n245_));
  NO2        m0217(.A(mai_mai_n245_), .B(mai_mai_n167_), .Y(mai_mai_n246_));
  INV        m0218(.A(mai_mai_n246_), .Y(mai_mai_n247_));
  NA3        m0219(.A(e), .B(c), .C(b), .Y(mai_mai_n248_));
  NO2        m0220(.A(d), .B(mai_mai_n248_), .Y(mai_mai_n249_));
  NAi32      m0221(.An(k), .Bn(i), .C(j), .Y(mai_mai_n250_));
  NAi31      m0222(.An(h), .B(l), .C(i), .Y(mai_mai_n251_));
  NA3        m0223(.A(mai_mai_n251_), .B(mai_mai_n250_), .C(mai_mai_n140_), .Y(mai_mai_n252_));
  NOi21      m0224(.An(mai_mai_n252_), .B(mai_mai_n46_), .Y(mai_mai_n253_));
  OAI210     m0225(.A0(mai_mai_n231_), .A1(mai_mai_n249_), .B0(mai_mai_n253_), .Y(mai_mai_n254_));
  NAi21      m0226(.An(l), .B(k), .Y(mai_mai_n255_));
  NO2        m0227(.A(mai_mai_n255_), .B(mai_mai_n46_), .Y(mai_mai_n256_));
  NOi21      m0228(.An(l), .B(j), .Y(mai_mai_n257_));
  NA2        m0229(.A(mai_mai_n137_), .B(mai_mai_n257_), .Y(mai_mai_n258_));
  NA3        m0230(.A(mai_mai_n100_), .B(mai_mai_n99_), .C(g), .Y(mai_mai_n259_));
  OR3        m0231(.A(mai_mai_n62_), .B(mai_mai_n63_), .C(e), .Y(mai_mai_n260_));
  AOI210     m0232(.A0(mai_mai_n259_), .A1(mai_mai_n258_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  INV        m0233(.A(mai_mai_n261_), .Y(mai_mai_n262_));
  NAi32      m0234(.An(j), .Bn(h), .C(i), .Y(mai_mai_n263_));
  NAi21      m0235(.An(m), .B(l), .Y(mai_mai_n264_));
  NO3        m0236(.A(mai_mai_n264_), .B(mai_mai_n263_), .C(mai_mai_n70_), .Y(mai_mai_n265_));
  NA2        m0237(.A(h), .B(g), .Y(mai_mai_n266_));
  NA2        m0238(.A(mai_mai_n143_), .B(mai_mai_n43_), .Y(mai_mai_n267_));
  NO2        m0239(.A(mai_mai_n267_), .B(mai_mai_n266_), .Y(mai_mai_n268_));
  OAI210     m0240(.A0(mai_mai_n268_), .A1(mai_mai_n265_), .B0(mai_mai_n138_), .Y(mai_mai_n269_));
  NA4        m0241(.A(mai_mai_n269_), .B(mai_mai_n262_), .C(mai_mai_n254_), .D(mai_mai_n247_), .Y(mai_mai_n270_));
  NAi32      m0242(.An(n), .Bn(m), .C(l), .Y(mai_mai_n271_));
  INV        m0243(.A(mai_mai_n103_), .Y(mai_mai_n272_));
  NAi31      m0244(.An(k), .B(l), .C(j), .Y(mai_mai_n273_));
  OAI210     m0245(.A0(mai_mai_n255_), .A1(j), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  BUFFER     m0246(.A(mai_mai_n274_), .Y(mai_mai_n275_));
  NA2        m0247(.A(mai_mai_n275_), .B(mai_mai_n272_), .Y(mai_mai_n276_));
  INV        m0248(.A(mai_mai_n276_), .Y(mai_mai_n277_));
  NO4        m0249(.A(mai_mai_n277_), .B(mai_mai_n270_), .C(mai_mai_n244_), .D(mai_mai_n237_), .Y(mai_mai_n278_));
  NA2        m0250(.A(mai_mai_n222_), .B(mai_mai_n166_), .Y(mai_mai_n279_));
  NAi21      m0251(.An(m), .B(k), .Y(mai_mai_n280_));
  NAi31      m0252(.An(i), .B(l), .C(h), .Y(mai_mai_n281_));
  NO4        m0253(.A(mai_mai_n281_), .B(e), .C(mai_mai_n62_), .D(mai_mai_n63_), .Y(mai_mai_n282_));
  NA2        m0254(.A(e), .B(c), .Y(mai_mai_n283_));
  NO3        m0255(.A(mai_mai_n283_), .B(n), .C(d), .Y(mai_mai_n284_));
  NA2        m0256(.A(f), .B(mai_mai_n100_), .Y(mai_mai_n285_));
  NO2        m0257(.A(mai_mai_n285_), .B(mai_mai_n184_), .Y(mai_mai_n286_));
  NAi31      m0258(.An(d), .B(e), .C(b), .Y(mai_mai_n287_));
  NO2        m0259(.A(mai_mai_n111_), .B(mai_mai_n287_), .Y(mai_mai_n288_));
  NA2        m0260(.A(mai_mai_n288_), .B(mai_mai_n286_), .Y(mai_mai_n289_));
  NAi31      m0261(.An(mai_mai_n282_), .B(mai_mai_n289_), .C(mai_mai_n279_), .Y(mai_mai_n290_));
  NA2        m0262(.A(mai_mai_n217_), .B(mai_mai_n87_), .Y(mai_mai_n291_));
  OR2        m0263(.A(mai_mai_n291_), .B(mai_mai_n178_), .Y(mai_mai_n292_));
  NOi31      m0264(.An(l), .B(n), .C(m), .Y(mai_mai_n293_));
  INV        m0265(.A(mai_mai_n292_), .Y(mai_mai_n294_));
  NAi32      m0266(.An(m), .Bn(j), .C(k), .Y(mai_mai_n295_));
  NAi41      m0267(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n296_));
  NOi31      m0268(.An(j), .B(m), .C(k), .Y(mai_mai_n297_));
  AN3        m0269(.A(h), .B(g), .C(f), .Y(mai_mai_n298_));
  NOi32      m0270(.An(m), .Bn(j), .C(l), .Y(mai_mai_n299_));
  NO2        m0271(.A(mai_mai_n299_), .B(mai_mai_n81_), .Y(mai_mai_n300_));
  INV        m0272(.A(mai_mai_n131_), .Y(mai_mai_n301_));
  INV        m0273(.A(mai_mai_n203_), .Y(mai_mai_n302_));
  NA3        m0274(.A(mai_mai_n302_), .B(mai_mai_n298_), .C(mai_mai_n182_), .Y(mai_mai_n303_));
  INV        m0275(.A(mai_mai_n303_), .Y(mai_mai_n304_));
  NA3        m0276(.A(h), .B(g), .C(f), .Y(mai_mai_n305_));
  NA2        m0277(.A(mai_mai_n137_), .B(e), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n137_), .B(mai_mai_n272_), .Y(mai_mai_n307_));
  NOi32      m0279(.An(j), .Bn(g), .C(i), .Y(mai_mai_n308_));
  NA3        m0280(.A(mai_mai_n308_), .B(mai_mai_n255_), .C(mai_mai_n96_), .Y(mai_mai_n309_));
  OR2        m0281(.A(mai_mai_n94_), .B(mai_mai_n309_), .Y(mai_mai_n310_));
  NOi32      m0282(.An(e), .Bn(b), .C(a), .Y(mai_mai_n311_));
  AN2        m0283(.A(l), .B(j), .Y(mai_mai_n312_));
  INV        m0284(.A(mai_mai_n179_), .Y(mai_mai_n313_));
  NA2        m0285(.A(mai_mai_n313_), .B(mai_mai_n311_), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n180_), .B(k), .Y(mai_mai_n315_));
  NA3        m0287(.A(m), .B(mai_mai_n95_), .C(mai_mai_n183_), .Y(mai_mai_n316_));
  NA4        m0288(.A(mai_mai_n177_), .B(mai_mai_n72_), .C(g), .D(mai_mai_n183_), .Y(mai_mai_n317_));
  NAi41      m0289(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n318_));
  NA2        m0290(.A(mai_mai_n47_), .B(mai_mai_n96_), .Y(mai_mai_n319_));
  NO2        m0291(.A(mai_mai_n319_), .B(mai_mai_n318_), .Y(mai_mai_n320_));
  NA3        m0292(.A(mai_mai_n314_), .B(mai_mai_n310_), .C(mai_mai_n307_), .Y(mai_mai_n321_));
  NO4        m0293(.A(mai_mai_n321_), .B(mai_mai_n304_), .C(mai_mai_n294_), .D(mai_mai_n290_), .Y(mai_mai_n322_));
  NA4        m0294(.A(mai_mai_n322_), .B(mai_mai_n278_), .C(mai_mai_n235_), .D(mai_mai_n173_), .Y(mai10));
  NA3        m0295(.A(m), .B(k), .C(i), .Y(mai_mai_n324_));
  NO3        m0296(.A(mai_mai_n324_), .B(j), .C(mai_mai_n184_), .Y(mai_mai_n325_));
  NOi21      m0297(.An(e), .B(f), .Y(mai_mai_n326_));
  NO4        m0298(.A(mai_mai_n126_), .B(mai_mai_n326_), .C(n), .D(mai_mai_n93_), .Y(mai_mai_n327_));
  NAi31      m0299(.An(b), .B(f), .C(c), .Y(mai_mai_n328_));
  INV        m0300(.A(mai_mai_n328_), .Y(mai_mai_n329_));
  NOi32      m0301(.An(k), .Bn(h), .C(j), .Y(mai_mai_n330_));
  NA2        m0302(.A(mai_mai_n330_), .B(mai_mai_n191_), .Y(mai_mai_n331_));
  NA2        m0303(.A(mai_mai_n135_), .B(mai_mai_n331_), .Y(mai_mai_n332_));
  AOI220     m0304(.A0(mai_mai_n332_), .A1(mai_mai_n329_), .B0(mai_mai_n327_), .B1(mai_mai_n325_), .Y(mai_mai_n333_));
  OR2        m0305(.A(m), .B(k), .Y(mai_mai_n334_));
  NO2        m0306(.A(mai_mai_n150_), .B(mai_mai_n334_), .Y(mai_mai_n335_));
  NA4        m0307(.A(n), .B(f), .C(c), .D(mai_mai_n98_), .Y(mai_mai_n336_));
  NOi32      m0308(.An(d), .Bn(a), .C(c), .Y(mai_mai_n337_));
  INV        m0309(.A(mai_mai_n337_), .Y(mai_mai_n338_));
  NAi31      m0310(.An(k), .B(m), .C(j), .Y(mai_mai_n339_));
  NO3        m0311(.A(mai_mai_n339_), .B(i), .C(n), .Y(mai_mai_n340_));
  NOi21      m0312(.An(mai_mai_n340_), .B(mai_mai_n338_), .Y(mai_mai_n341_));
  INV        m0313(.A(mai_mai_n341_), .Y(mai_mai_n342_));
  NO2        m0314(.A(mai_mai_n336_), .B(mai_mai_n264_), .Y(mai_mai_n343_));
  NOi32      m0315(.An(f), .Bn(d), .C(c), .Y(mai_mai_n344_));
  NA2        m0316(.A(mai_mai_n343_), .B(mai_mai_n185_), .Y(mai_mai_n345_));
  NA3        m0317(.A(mai_mai_n345_), .B(mai_mai_n342_), .C(mai_mai_n333_), .Y(mai_mai_n346_));
  NA2        m0318(.A(mai_mai_n217_), .B(b), .Y(mai_mai_n347_));
  INV        m0319(.A(e), .Y(mai_mai_n348_));
  NA2        m0320(.A(mai_mai_n44_), .B(e), .Y(mai_mai_n349_));
  OAI220     m0321(.A0(mai_mai_n349_), .A1(mai_mai_n174_), .B0(mai_mai_n178_), .B1(mai_mai_n348_), .Y(mai_mai_n350_));
  NA3        m0322(.A(e), .B(mai_mai_n177_), .C(i), .Y(mai_mai_n351_));
  INV        m0323(.A(mai_mai_n351_), .Y(mai_mai_n352_));
  NO2        m0324(.A(mai_mai_n84_), .B(mai_mai_n348_), .Y(mai_mai_n353_));
  NO3        m0325(.A(mai_mai_n353_), .B(mai_mai_n352_), .C(mai_mai_n350_), .Y(mai_mai_n354_));
  NOi32      m0326(.An(h), .Bn(e), .C(g), .Y(mai_mai_n355_));
  NA3        m0327(.A(mai_mai_n355_), .B(mai_mai_n257_), .C(m), .Y(mai_mai_n356_));
  NOi21      m0328(.An(g), .B(h), .Y(mai_mai_n357_));
  AN3        m0329(.A(m), .B(l), .C(i), .Y(mai_mai_n358_));
  NA3        m0330(.A(mai_mai_n358_), .B(mai_mai_n357_), .C(e), .Y(mai_mai_n359_));
  AN3        m0331(.A(h), .B(g), .C(e), .Y(mai_mai_n360_));
  NA2        m0332(.A(mai_mai_n360_), .B(mai_mai_n81_), .Y(mai_mai_n361_));
  AN3        m0333(.A(mai_mai_n361_), .B(mai_mai_n359_), .C(mai_mai_n356_), .Y(mai_mai_n362_));
  AOI210     m0334(.A0(mai_mai_n362_), .A1(mai_mai_n354_), .B0(mai_mai_n347_), .Y(mai_mai_n363_));
  NA3        m0335(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(e), .Y(mai_mai_n364_));
  NO2        m0336(.A(mai_mai_n364_), .B(mai_mai_n347_), .Y(mai_mai_n365_));
  NA2        m0337(.A(mai_mai_n337_), .B(mai_mai_n70_), .Y(mai_mai_n366_));
  NAi31      m0338(.An(b), .B(c), .C(a), .Y(mai_mai_n367_));
  NO2        m0339(.A(mai_mai_n367_), .B(n), .Y(mai_mai_n368_));
  NO3        m0340(.A(mai_mai_n365_), .B(mai_mai_n363_), .C(mai_mai_n346_), .Y(mai_mai_n369_));
  NA2        m0341(.A(i), .B(g), .Y(mai_mai_n370_));
  NO3        m0342(.A(mai_mai_n242_), .B(mai_mai_n370_), .C(c), .Y(mai_mai_n371_));
  NOi21      m0343(.An(a), .B(n), .Y(mai_mai_n372_));
  NOi21      m0344(.An(d), .B(c), .Y(mai_mai_n373_));
  NA2        m0345(.A(mai_mai_n373_), .B(mai_mai_n372_), .Y(mai_mai_n374_));
  NA3        m0346(.A(i), .B(g), .C(f), .Y(mai_mai_n375_));
  OR2        m0347(.A(mai_mai_n375_), .B(mai_mai_n61_), .Y(mai_mai_n376_));
  NA2        m0348(.A(mai_mai_n358_), .B(mai_mai_n357_), .Y(mai_mai_n377_));
  AOI210     m0349(.A0(mai_mai_n377_), .A1(mai_mai_n376_), .B0(mai_mai_n374_), .Y(mai_mai_n378_));
  AOI210     m0350(.A0(mai_mai_n371_), .A1(mai_mai_n256_), .B0(mai_mai_n378_), .Y(mai_mai_n379_));
  OR2        m0351(.A(n), .B(m), .Y(mai_mai_n380_));
  NO2        m0352(.A(mai_mai_n380_), .B(mai_mai_n127_), .Y(mai_mai_n381_));
  NO2        m0353(.A(mai_mai_n158_), .B(mai_mai_n123_), .Y(mai_mai_n382_));
  OAI210     m0354(.A0(mai_mai_n381_), .A1(mai_mai_n152_), .B0(mai_mai_n382_), .Y(mai_mai_n383_));
  INV        m0355(.A(mai_mai_n319_), .Y(mai_mai_n384_));
  NA2        m0356(.A(mai_mai_n384_), .B(mai_mai_n311_), .Y(mai_mai_n385_));
  NO2        m0357(.A(mai_mai_n367_), .B(mai_mai_n46_), .Y(mai_mai_n386_));
  NAi21      m0358(.An(k), .B(j), .Y(mai_mai_n387_));
  NAi21      m0359(.An(e), .B(d), .Y(mai_mai_n388_));
  INV        m0360(.A(mai_mai_n388_), .Y(mai_mai_n389_));
  NO2        m0361(.A(mai_mai_n221_), .B(mai_mai_n183_), .Y(mai_mai_n390_));
  NA3        m0362(.A(mai_mai_n390_), .B(mai_mai_n389_), .C(mai_mai_n197_), .Y(mai_mai_n391_));
  NA3        m0363(.A(mai_mai_n391_), .B(mai_mai_n385_), .C(mai_mai_n383_), .Y(mai_mai_n392_));
  NAi31      m0364(.An(g), .B(f), .C(c), .Y(mai_mai_n393_));
  NOi31      m0365(.An(mai_mai_n379_), .B(mai_mai_n392_), .C(mai_mai_n234_), .Y(mai_mai_n394_));
  NOi32      m0366(.An(c), .Bn(a), .C(b), .Y(mai_mai_n395_));
  NA2        m0367(.A(mai_mai_n395_), .B(mai_mai_n96_), .Y(mai_mai_n396_));
  AN2        m0368(.A(e), .B(d), .Y(mai_mai_n397_));
  NO2        m0369(.A(mai_mai_n110_), .B(mai_mai_n39_), .Y(mai_mai_n398_));
  NO2        m0370(.A(mai_mai_n57_), .B(e), .Y(mai_mai_n399_));
  NOi31      m0371(.An(j), .B(k), .C(i), .Y(mai_mai_n400_));
  NOi21      m0372(.An(mai_mai_n140_), .B(mai_mai_n400_), .Y(mai_mai_n401_));
  NO2        m0373(.A(e), .B(mai_mai_n396_), .Y(mai_mai_n402_));
  NOi21      m0374(.An(a), .B(b), .Y(mai_mai_n403_));
  NA3        m0375(.A(e), .B(d), .C(c), .Y(mai_mai_n404_));
  NAi21      m0376(.An(mai_mai_n404_), .B(mai_mai_n403_), .Y(mai_mai_n405_));
  NO2        m0377(.A(mai_mai_n1235_), .B(mai_mai_n405_), .Y(mai_mai_n406_));
  NO4        m0378(.A(mai_mai_n161_), .B(mai_mai_n86_), .C(mai_mai_n49_), .D(b), .Y(mai_mai_n407_));
  NA2        m0379(.A(mai_mai_n329_), .B(mai_mai_n128_), .Y(mai_mai_n408_));
  OR2        m0380(.A(k), .B(j), .Y(mai_mai_n409_));
  NA2        m0381(.A(l), .B(k), .Y(mai_mai_n410_));
  NA3        m0382(.A(mai_mai_n410_), .B(mai_mai_n409_), .C(mai_mai_n191_), .Y(mai_mai_n411_));
  AOI210     m0383(.A0(mai_mai_n203_), .A1(mai_mai_n295_), .B0(mai_mai_n70_), .Y(mai_mai_n412_));
  NOi21      m0384(.An(mai_mai_n411_), .B(mai_mai_n412_), .Y(mai_mai_n413_));
  OR3        m0385(.A(mai_mai_n413_), .B(mai_mai_n121_), .C(mai_mai_n113_), .Y(mai_mai_n414_));
  INV        m0386(.A(mai_mai_n107_), .Y(mai_mai_n415_));
  NA2        m0387(.A(mai_mai_n337_), .B(mai_mai_n96_), .Y(mai_mai_n416_));
  NO4        m0388(.A(mai_mai_n416_), .B(mai_mai_n79_), .C(mai_mai_n95_), .D(e), .Y(mai_mai_n417_));
  NO3        m0389(.A(mai_mai_n366_), .B(mai_mai_n76_), .C(mai_mai_n110_), .Y(mai_mai_n418_));
  NO4        m0390(.A(mai_mai_n418_), .B(mai_mai_n417_), .C(mai_mai_n415_), .D(mai_mai_n282_), .Y(mai_mai_n419_));
  NA3        m0391(.A(mai_mai_n419_), .B(mai_mai_n414_), .C(mai_mai_n408_), .Y(mai_mai_n420_));
  NO4        m0392(.A(mai_mai_n420_), .B(mai_mai_n407_), .C(mai_mai_n406_), .D(mai_mai_n402_), .Y(mai_mai_n421_));
  NOi21      m0393(.An(d), .B(e), .Y(mai_mai_n422_));
  NAi31      m0394(.An(j), .B(l), .C(i), .Y(mai_mai_n423_));
  OAI210     m0395(.A0(mai_mai_n423_), .A1(mai_mai_n111_), .B0(mai_mai_n86_), .Y(mai_mai_n424_));
  NO3        m0396(.A(mai_mai_n338_), .B(mai_mai_n300_), .C(mai_mai_n175_), .Y(mai_mai_n425_));
  INV        m0397(.A(mai_mai_n425_), .Y(mai_mai_n426_));
  NA2        m0398(.A(mai_mai_n426_), .B(mai_mai_n209_), .Y(mai_mai_n427_));
  OAI210     m0399(.A0(mai_mai_n106_), .A1(mai_mai_n105_), .B0(n), .Y(mai_mai_n428_));
  NO2        m0400(.A(mai_mai_n428_), .B(mai_mai_n110_), .Y(mai_mai_n429_));
  OA210      m0401(.A0(mai_mai_n211_), .A1(mai_mai_n429_), .B0(mai_mai_n166_), .Y(mai_mai_n430_));
  XO2        m0402(.A(i), .B(h), .Y(mai_mai_n431_));
  BUFFER     m0403(.A(mai_mai_n265_), .Y(mai_mai_n432_));
  NAi31      m0404(.An(c), .B(f), .C(d), .Y(mai_mai_n433_));
  AOI210     m0405(.A0(mai_mai_n245_), .A1(mai_mai_n169_), .B0(mai_mai_n433_), .Y(mai_mai_n434_));
  INV        m0406(.A(mai_mai_n434_), .Y(mai_mai_n435_));
  NA3        m0407(.A(mai_mai_n327_), .B(mai_mai_n81_), .C(j), .Y(mai_mai_n436_));
  NA2        m0408(.A(mai_mai_n198_), .B(mai_mai_n91_), .Y(mai_mai_n437_));
  NO2        m0409(.A(mai_mai_n437_), .B(mai_mai_n433_), .Y(mai_mai_n438_));
  NOi21      m0410(.An(mai_mai_n436_), .B(mai_mai_n438_), .Y(mai_mai_n439_));
  AO220      m0411(.A0(mai_mai_n253_), .A1(mai_mai_n231_), .B0(mai_mai_n141_), .B1(mai_mai_n58_), .Y(mai_mai_n440_));
  NA3        m0412(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(f), .Y(mai_mai_n441_));
  NO2        m0413(.A(mai_mai_n441_), .B(mai_mai_n374_), .Y(mai_mai_n442_));
  NO2        m0414(.A(mai_mai_n442_), .B(mai_mai_n261_), .Y(mai_mai_n443_));
  NAi41      m0415(.An(mai_mai_n440_), .B(mai_mai_n443_), .C(mai_mai_n439_), .D(mai_mai_n435_), .Y(mai_mai_n444_));
  NO3        m0416(.A(mai_mai_n444_), .B(mai_mai_n430_), .C(mai_mai_n427_), .Y(mai_mai_n445_));
  NA4        m0417(.A(mai_mai_n445_), .B(mai_mai_n421_), .C(mai_mai_n394_), .D(mai_mai_n369_), .Y(mai11));
  NO2        m0418(.A(mai_mai_n62_), .B(f), .Y(mai_mai_n447_));
  NA2        m0419(.A(j), .B(g), .Y(mai_mai_n448_));
  NAi31      m0420(.An(i), .B(m), .C(l), .Y(mai_mai_n449_));
  NA3        m0421(.A(m), .B(k), .C(j), .Y(mai_mai_n450_));
  OAI220     m0422(.A0(mai_mai_n450_), .A1(mai_mai_n110_), .B0(mai_mai_n449_), .B1(mai_mai_n448_), .Y(mai_mai_n451_));
  NA2        m0423(.A(mai_mai_n451_), .B(mai_mai_n447_), .Y(mai_mai_n452_));
  NOi32      m0424(.An(e), .Bn(b), .C(f), .Y(mai_mai_n453_));
  NA2        m0425(.A(mai_mai_n44_), .B(j), .Y(mai_mai_n454_));
  NAi31      m0426(.An(d), .B(e), .C(a), .Y(mai_mai_n455_));
  NO2        m0427(.A(mai_mai_n455_), .B(n), .Y(mai_mai_n456_));
  NA2        m0428(.A(mai_mai_n143_), .B(mai_mai_n453_), .Y(mai_mai_n457_));
  NAi41      m0429(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n458_));
  BUFFER     m0430(.A(mai_mai_n318_), .Y(mai_mai_n459_));
  NA2        m0431(.A(j), .B(i), .Y(mai_mai_n460_));
  NAi31      m0432(.An(n), .B(m), .C(k), .Y(mai_mai_n461_));
  NO3        m0433(.A(mai_mai_n461_), .B(mai_mai_n460_), .C(mai_mai_n95_), .Y(mai_mai_n462_));
  NO4        m0434(.A(n), .B(d), .C(mai_mai_n98_), .D(a), .Y(mai_mai_n463_));
  OR2        m0435(.A(n), .B(c), .Y(mai_mai_n464_));
  NO2        m0436(.A(mai_mai_n464_), .B(mai_mai_n125_), .Y(mai_mai_n465_));
  NO2        m0437(.A(mai_mai_n465_), .B(mai_mai_n463_), .Y(mai_mai_n466_));
  NOi32      m0438(.An(g), .Bn(f), .C(i), .Y(mai_mai_n467_));
  AOI220     m0439(.A0(mai_mai_n467_), .A1(mai_mai_n83_), .B0(mai_mai_n451_), .B1(f), .Y(mai_mai_n468_));
  NO2        m0440(.A(mai_mai_n468_), .B(mai_mai_n466_), .Y(mai_mai_n469_));
  INV        m0441(.A(mai_mai_n469_), .Y(mai_mai_n470_));
  NA2        m0442(.A(mai_mai_n118_), .B(mai_mai_n34_), .Y(mai_mai_n471_));
  NAi32      m0443(.An(e), .Bn(b), .C(c), .Y(mai_mai_n472_));
  OAI220     m0444(.A0(mai_mai_n339_), .A1(i), .B0(mai_mai_n449_), .B1(mai_mai_n448_), .Y(mai_mai_n473_));
  NAi31      m0445(.An(d), .B(c), .C(a), .Y(mai_mai_n474_));
  NO2        m0446(.A(mai_mai_n474_), .B(n), .Y(mai_mai_n475_));
  NA3        m0447(.A(mai_mai_n475_), .B(mai_mai_n473_), .C(e), .Y(mai_mai_n476_));
  NO3        m0448(.A(mai_mai_n53_), .B(mai_mai_n46_), .C(mai_mai_n184_), .Y(mai_mai_n477_));
  NA2        m0449(.A(mai_mai_n477_), .B(mai_mai_n1241_), .Y(mai_mai_n478_));
  NA2        m0450(.A(mai_mai_n478_), .B(mai_mai_n476_), .Y(mai_mai_n479_));
  NO2        m0451(.A(mai_mai_n242_), .B(n), .Y(mai_mai_n480_));
  NO2        m0452(.A(mai_mai_n368_), .B(mai_mai_n480_), .Y(mai_mai_n481_));
  NA2        m0453(.A(mai_mai_n473_), .B(f), .Y(mai_mai_n482_));
  NAi32      m0454(.An(d), .Bn(a), .C(b), .Y(mai_mai_n483_));
  NO2        m0455(.A(mai_mai_n483_), .B(mai_mai_n46_), .Y(mai_mai_n484_));
  NA2        m0456(.A(h), .B(f), .Y(mai_mai_n485_));
  NO2        m0457(.A(mai_mai_n485_), .B(mai_mai_n79_), .Y(mai_mai_n486_));
  NA2        m0458(.A(mai_mai_n486_), .B(mai_mai_n484_), .Y(mai_mai_n487_));
  OAI210     m0459(.A0(mai_mai_n482_), .A1(mai_mai_n481_), .B0(mai_mai_n487_), .Y(mai_mai_n488_));
  NO2        m0460(.A(mai_mai_n122_), .B(c), .Y(mai_mai_n489_));
  NA3        m0461(.A(f), .B(d), .C(b), .Y(mai_mai_n490_));
  NO2        m0462(.A(mai_mai_n488_), .B(mai_mai_n479_), .Y(mai_mai_n491_));
  AN4        m0463(.A(mai_mai_n491_), .B(mai_mai_n470_), .C(mai_mai_n457_), .D(mai_mai_n452_), .Y(mai_mai_n492_));
  INV        m0464(.A(k), .Y(mai_mai_n493_));
  NA3        m0465(.A(l), .B(mai_mai_n493_), .C(i), .Y(mai_mai_n494_));
  NA2        m0466(.A(mai_mai_n337_), .B(mai_mai_n96_), .Y(mai_mai_n495_));
  NAi32      m0467(.An(h), .Bn(f), .C(g), .Y(mai_mai_n496_));
  NAi41      m0468(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n497_));
  OAI210     m0469(.A0(mai_mai_n455_), .A1(n), .B0(mai_mai_n497_), .Y(mai_mai_n498_));
  NA2        m0470(.A(mai_mai_n498_), .B(m), .Y(mai_mai_n499_));
  NAi31      m0471(.An(h), .B(g), .C(f), .Y(mai_mai_n500_));
  OR3        m0472(.A(mai_mai_n500_), .B(mai_mai_n242_), .C(mai_mai_n46_), .Y(mai_mai_n501_));
  NA4        m0473(.A(mai_mai_n357_), .B(mai_mai_n102_), .C(mai_mai_n96_), .D(e), .Y(mai_mai_n502_));
  AN2        m0474(.A(mai_mai_n502_), .B(mai_mai_n501_), .Y(mai_mai_n503_));
  OA210      m0475(.A0(mai_mai_n499_), .A1(mai_mai_n496_), .B0(mai_mai_n503_), .Y(mai_mai_n504_));
  NO3        m0476(.A(mai_mai_n496_), .B(mai_mai_n62_), .C(mai_mai_n63_), .Y(mai_mai_n505_));
  NO4        m0477(.A(mai_mai_n500_), .B(mai_mai_n464_), .C(mai_mai_n125_), .D(mai_mai_n63_), .Y(mai_mai_n506_));
  OR2        m0478(.A(mai_mai_n506_), .B(mai_mai_n505_), .Y(mai_mai_n507_));
  NAi31      m0479(.An(mai_mai_n507_), .B(mai_mai_n504_), .C(mai_mai_n495_), .Y(mai_mai_n508_));
  NOi32      m0480(.An(b), .Bn(a), .C(c), .Y(mai_mai_n509_));
  NOi32      m0481(.An(d), .Bn(a), .C(e), .Y(mai_mai_n510_));
  NA2        m0482(.A(mai_mai_n510_), .B(mai_mai_n96_), .Y(mai_mai_n511_));
  NO2        m0483(.A(n), .B(c), .Y(mai_mai_n512_));
  NA3        m0484(.A(mai_mai_n512_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n513_));
  NOi32      m0485(.An(e), .Bn(a), .C(d), .Y(mai_mai_n514_));
  AOI210     m0486(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n514_), .Y(mai_mai_n515_));
  INV        m0487(.A(mai_mai_n471_), .Y(mai_mai_n516_));
  NA2        m0488(.A(mai_mai_n516_), .B(mai_mai_n96_), .Y(mai_mai_n517_));
  NA2        m0489(.A(mai_mai_n216_), .B(mai_mai_n517_), .Y(mai_mai_n518_));
  AOI210     m0490(.A0(mai_mai_n508_), .A1(mai_mai_n493_), .B0(mai_mai_n518_), .Y(mai_mai_n519_));
  NO3        m0491(.A(mai_mai_n280_), .B(mai_mai_n52_), .C(n), .Y(mai_mai_n520_));
  NA3        m0492(.A(mai_mai_n433_), .B(mai_mai_n148_), .C(mai_mai_n147_), .Y(mai_mai_n521_));
  NA2        m0493(.A(mai_mai_n393_), .B(mai_mai_n201_), .Y(mai_mai_n522_));
  OR2        m0494(.A(mai_mai_n522_), .B(mai_mai_n521_), .Y(mai_mai_n523_));
  NA2        m0495(.A(mai_mai_n64_), .B(mai_mai_n96_), .Y(mai_mai_n524_));
  NA2        m0496(.A(mai_mai_n523_), .B(mai_mai_n520_), .Y(mai_mai_n525_));
  NO2        m0497(.A(mai_mai_n525_), .B(mai_mai_n72_), .Y(mai_mai_n526_));
  NOi32      m0498(.An(e), .Bn(c), .C(f), .Y(mai_mai_n527_));
  NOi21      m0499(.An(f), .B(g), .Y(mai_mai_n528_));
  NO2        m0500(.A(mai_mai_n528_), .B(mai_mai_n181_), .Y(mai_mai_n529_));
  INV        m0501(.A(mai_mai_n155_), .Y(mai_mai_n530_));
  AOI210     m0502(.A0(mai_mai_n459_), .A1(mai_mai_n338_), .B0(mai_mai_n266_), .Y(mai_mai_n531_));
  NAi21      m0503(.An(k), .B(h), .Y(mai_mai_n532_));
  NO2        m0504(.A(mai_mai_n532_), .B(mai_mai_n230_), .Y(mai_mai_n533_));
  INV        m0505(.A(mai_mai_n533_), .Y(mai_mai_n534_));
  OR2        m0506(.A(mai_mai_n534_), .B(mai_mai_n499_), .Y(mai_mai_n535_));
  NOi31      m0507(.An(m), .B(n), .C(k), .Y(mai_mai_n536_));
  INV        m0508(.A(mai_mai_n536_), .Y(mai_mai_n537_));
  AOI210     m0509(.A0(mai_mai_n338_), .A1(mai_mai_n318_), .B0(mai_mai_n266_), .Y(mai_mai_n538_));
  NAi21      m0510(.An(mai_mai_n537_), .B(mai_mai_n538_), .Y(mai_mai_n539_));
  NO2        m0511(.A(mai_mai_n242_), .B(mai_mai_n46_), .Y(mai_mai_n540_));
  NO2        m0512(.A(mai_mai_n455_), .B(mai_mai_n46_), .Y(mai_mai_n541_));
  NA2        m0513(.A(mai_mai_n540_), .B(mai_mai_n486_), .Y(mai_mai_n542_));
  NA3        m0514(.A(mai_mai_n542_), .B(mai_mai_n539_), .C(mai_mai_n535_), .Y(mai_mai_n543_));
  NA2        m0515(.A(mai_mai_n91_), .B(mai_mai_n35_), .Y(mai_mai_n544_));
  NO2        m0516(.A(k), .B(mai_mai_n184_), .Y(mai_mai_n545_));
  NO2        m0517(.A(mai_mai_n453_), .B(mai_mai_n311_), .Y(mai_mai_n546_));
  NO2        m0518(.A(mai_mai_n546_), .B(n), .Y(mai_mai_n547_));
  NAi21      m0519(.An(mai_mai_n544_), .B(mai_mai_n547_), .Y(mai_mai_n548_));
  NA2        m0520(.A(mai_mai_n431_), .B(mai_mai_n134_), .Y(mai_mai_n549_));
  NO3        m0521(.A(mai_mai_n336_), .B(mai_mai_n549_), .C(mai_mai_n72_), .Y(mai_mai_n550_));
  INV        m0522(.A(mai_mai_n550_), .Y(mai_mai_n551_));
  AN3        m0523(.A(f), .B(d), .C(b), .Y(mai_mai_n552_));
  OAI210     m0524(.A0(mai_mai_n552_), .A1(mai_mai_n109_), .B0(n), .Y(mai_mai_n553_));
  NA3        m0525(.A(mai_mai_n431_), .B(mai_mai_n134_), .C(mai_mai_n184_), .Y(mai_mai_n554_));
  AOI210     m0526(.A0(mai_mai_n553_), .A1(mai_mai_n202_), .B0(mai_mai_n554_), .Y(mai_mai_n555_));
  NAi31      m0527(.An(m), .B(n), .C(k), .Y(mai_mai_n556_));
  OR2        m0528(.A(mai_mai_n113_), .B(mai_mai_n52_), .Y(mai_mai_n557_));
  OAI210     m0529(.A0(mai_mai_n557_), .A1(mai_mai_n556_), .B0(mai_mai_n218_), .Y(mai_mai_n558_));
  OAI210     m0530(.A0(mai_mai_n558_), .A1(mai_mai_n555_), .B0(j), .Y(mai_mai_n559_));
  NA3        m0531(.A(mai_mai_n559_), .B(mai_mai_n551_), .C(mai_mai_n548_), .Y(mai_mai_n560_));
  NO4        m0532(.A(mai_mai_n560_), .B(mai_mai_n543_), .C(mai_mai_n530_), .D(mai_mai_n526_), .Y(mai_mai_n561_));
  NAi31      m0533(.An(g), .B(h), .C(f), .Y(mai_mai_n562_));
  OR3        m0534(.A(mai_mai_n562_), .B(mai_mai_n242_), .C(n), .Y(mai_mai_n563_));
  OA210      m0535(.A0(mai_mai_n455_), .A1(n), .B0(mai_mai_n497_), .Y(mai_mai_n564_));
  NA3        m0536(.A(mai_mai_n355_), .B(mai_mai_n102_), .C(mai_mai_n70_), .Y(mai_mai_n565_));
  OAI210     m0537(.A0(mai_mai_n564_), .A1(mai_mai_n75_), .B0(mai_mai_n565_), .Y(mai_mai_n566_));
  NOi21      m0538(.An(mai_mai_n563_), .B(mai_mai_n566_), .Y(mai_mai_n567_));
  NO2        m0539(.A(mai_mai_n567_), .B(mai_mai_n450_), .Y(mai_mai_n568_));
  NO3        m0540(.A(g), .B(mai_mai_n183_), .C(mai_mai_n49_), .Y(mai_mai_n569_));
  NO2        m0541(.A(mai_mai_n437_), .B(mai_mai_n72_), .Y(mai_mai_n570_));
  OAI210     m0542(.A0(mai_mai_n570_), .A1(mai_mai_n335_), .B0(mai_mai_n569_), .Y(mai_mai_n571_));
  OR2        m0543(.A(mai_mai_n62_), .B(mai_mai_n63_), .Y(mai_mai_n572_));
  NA2        m0544(.A(mai_mai_n509_), .B(mai_mai_n298_), .Y(mai_mai_n573_));
  OA220      m0545(.A0(mai_mai_n537_), .A1(mai_mai_n573_), .B0(mai_mai_n534_), .B1(mai_mai_n572_), .Y(mai_mai_n574_));
  NA2        m0546(.A(h), .B(mai_mai_n36_), .Y(mai_mai_n575_));
  NA2        m0547(.A(mai_mai_n83_), .B(mai_mai_n44_), .Y(mai_mai_n576_));
  OAI220     m0548(.A0(mai_mai_n576_), .A1(mai_mai_n291_), .B0(mai_mai_n575_), .B1(mai_mai_n396_), .Y(mai_mai_n577_));
  AOI210     m0549(.A0(mai_mai_n483_), .A1(mai_mai_n367_), .B0(mai_mai_n46_), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n500_), .B(mai_mai_n494_), .Y(mai_mai_n579_));
  AOI210     m0551(.A0(mai_mai_n579_), .A1(mai_mai_n578_), .B0(mai_mai_n577_), .Y(mai_mai_n580_));
  NA3        m0552(.A(mai_mai_n580_), .B(mai_mai_n574_), .C(mai_mai_n571_), .Y(mai_mai_n581_));
  NO2        m0553(.A(mai_mai_n220_), .B(f), .Y(mai_mai_n582_));
  INV        m0554(.A(mai_mai_n288_), .Y(mai_mai_n583_));
  OR2        m0555(.A(mai_mai_n309_), .B(mai_mai_n94_), .Y(mai_mai_n584_));
  OAI210     m0556(.A0(mai_mai_n583_), .A1(mai_mai_n528_), .B0(mai_mai_n584_), .Y(mai_mai_n585_));
  NO3        m0557(.A(mai_mai_n344_), .B(mai_mai_n166_), .C(mai_mai_n165_), .Y(mai_mai_n586_));
  NA2        m0558(.A(mai_mai_n586_), .B(mai_mai_n201_), .Y(mai_mai_n587_));
  NA3        m0559(.A(mai_mai_n587_), .B(mai_mai_n222_), .C(j), .Y(mai_mai_n588_));
  NA2        m0560(.A(mai_mai_n395_), .B(mai_mai_n70_), .Y(mai_mai_n589_));
  NO3        m0561(.A(mai_mai_n450_), .B(mai_mai_n589_), .C(mai_mai_n110_), .Y(mai_mai_n590_));
  INV        m0562(.A(mai_mai_n590_), .Y(mai_mai_n591_));
  NA4        m0563(.A(mai_mai_n591_), .B(mai_mai_n588_), .C(mai_mai_n436_), .D(mai_mai_n342_), .Y(mai_mai_n592_));
  NO4        m0564(.A(mai_mai_n592_), .B(mai_mai_n585_), .C(mai_mai_n581_), .D(mai_mai_n568_), .Y(mai_mai_n593_));
  NA4        m0565(.A(mai_mai_n593_), .B(mai_mai_n561_), .C(mai_mai_n519_), .D(mai_mai_n492_), .Y(mai08));
  NO2        m0566(.A(k), .B(h), .Y(mai_mai_n595_));
  AO210      m0567(.A0(mai_mai_n220_), .A1(mai_mai_n387_), .B0(mai_mai_n595_), .Y(mai_mai_n596_));
  NO2        m0568(.A(mai_mai_n596_), .B(mai_mai_n264_), .Y(mai_mai_n597_));
  NA2        m0569(.A(mai_mai_n527_), .B(mai_mai_n70_), .Y(mai_mai_n598_));
  NA2        m0570(.A(mai_mai_n598_), .B(mai_mai_n393_), .Y(mai_mai_n599_));
  AOI210     m0571(.A0(mai_mai_n599_), .A1(mai_mai_n597_), .B0(mai_mai_n418_), .Y(mai_mai_n600_));
  NA2        m0572(.A(mai_mai_n70_), .B(mai_mai_n93_), .Y(mai_mai_n601_));
  NO2        m0573(.A(mai_mai_n601_), .B(mai_mai_n50_), .Y(mai_mai_n602_));
  NA4        m0574(.A(mai_mai_n186_), .B(mai_mai_n118_), .C(mai_mai_n43_), .D(h), .Y(mai_mai_n603_));
  AN2        m0575(.A(l), .B(k), .Y(mai_mai_n604_));
  INV        m0576(.A(mai_mai_n600_), .Y(mai_mai_n605_));
  AN2        m0577(.A(mai_mai_n456_), .B(mai_mai_n80_), .Y(mai_mai_n606_));
  NO4        m0578(.A(mai_mai_n150_), .B(mai_mai_n334_), .C(mai_mai_n95_), .D(g), .Y(mai_mai_n607_));
  INV        m0579(.A(mai_mai_n442_), .Y(mai_mai_n608_));
  INV        m0580(.A(mai_mai_n37_), .Y(mai_mai_n609_));
  NA2        m0581(.A(mai_mai_n609_), .B(mai_mai_n480_), .Y(mai_mai_n610_));
  NA2        m0582(.A(mai_mai_n610_), .B(mai_mai_n608_), .Y(mai_mai_n611_));
  NO2        m0583(.A(mai_mai_n410_), .B(mai_mai_n111_), .Y(mai_mai_n612_));
  NA2        m0584(.A(mai_mai_n612_), .B(mai_mai_n1237_), .Y(mai_mai_n613_));
  NA2        m0585(.A(mai_mai_n596_), .B(mai_mai_n114_), .Y(mai_mai_n614_));
  NA2        m0586(.A(mai_mai_n614_), .B(mai_mai_n343_), .Y(mai_mai_n615_));
  NA2        m0587(.A(mai_mai_n613_), .B(mai_mai_n615_), .Y(mai_mai_n616_));
  NA2        m0588(.A(mai_mai_n311_), .B(mai_mai_n41_), .Y(mai_mai_n617_));
  NA3        m0589(.A(mai_mai_n587_), .B(mai_mai_n293_), .C(mai_mai_n330_), .Y(mai_mai_n618_));
  NA2        m0590(.A(mai_mai_n604_), .B(mai_mai_n191_), .Y(mai_mai_n619_));
  NO2        m0591(.A(mai_mai_n619_), .B(mai_mai_n287_), .Y(mai_mai_n620_));
  AOI210     m0592(.A0(mai_mai_n620_), .A1(mai_mai_n582_), .B0(mai_mai_n417_), .Y(mai_mai_n621_));
  NA3        m0593(.A(m), .B(l), .C(k), .Y(mai_mai_n622_));
  AOI210     m0594(.A0(mai_mai_n565_), .A1(mai_mai_n563_), .B0(mai_mai_n622_), .Y(mai_mai_n623_));
  NO2        m0595(.A(mai_mai_n458_), .B(mai_mai_n238_), .Y(mai_mai_n624_));
  NOi21      m0596(.An(mai_mai_n624_), .B(n), .Y(mai_mai_n625_));
  NA4        m0597(.A(mai_mai_n96_), .B(l), .C(k), .D(mai_mai_n72_), .Y(mai_mai_n626_));
  NA3        m0598(.A(mai_mai_n102_), .B(e), .C(i), .Y(mai_mai_n627_));
  NO2        m0599(.A(mai_mai_n627_), .B(mai_mai_n626_), .Y(mai_mai_n628_));
  NO3        m0600(.A(mai_mai_n628_), .B(mai_mai_n625_), .C(mai_mai_n623_), .Y(mai_mai_n629_));
  NA4        m0601(.A(mai_mai_n629_), .B(mai_mai_n621_), .C(mai_mai_n618_), .D(mai_mai_n617_), .Y(mai_mai_n630_));
  NO4        m0602(.A(mai_mai_n630_), .B(mai_mai_n616_), .C(mai_mai_n611_), .D(mai_mai_n605_), .Y(mai_mai_n631_));
  NA2        m0603(.A(mai_mai_n529_), .B(mai_mai_n335_), .Y(mai_mai_n632_));
  NOi31      m0604(.An(g), .B(h), .C(f), .Y(mai_mai_n633_));
  NA2        m0605(.A(mai_mai_n541_), .B(mai_mai_n633_), .Y(mai_mai_n634_));
  NO3        m0606(.A(mai_mai_n338_), .B(mai_mai_n448_), .C(h), .Y(mai_mai_n635_));
  NA2        m0607(.A(mai_mai_n635_), .B(mai_mai_n96_), .Y(mai_mai_n636_));
  NA4        m0608(.A(mai_mai_n636_), .B(mai_mai_n634_), .C(mai_mai_n632_), .D(mai_mai_n219_), .Y(mai_mai_n637_));
  NA2        m0609(.A(mai_mai_n604_), .B(mai_mai_n63_), .Y(mai_mai_n638_));
  NO3        m0610(.A(mai_mai_n586_), .B(mai_mai_n150_), .C(i), .Y(mai_mai_n639_));
  NOi21      m0611(.An(h), .B(j), .Y(mai_mai_n640_));
  NA2        m0612(.A(mai_mai_n640_), .B(f), .Y(mai_mai_n641_));
  NO2        m0613(.A(mai_mai_n641_), .B(mai_mai_n213_), .Y(mai_mai_n642_));
  NO2        m0614(.A(mai_mai_n642_), .B(mai_mai_n639_), .Y(mai_mai_n643_));
  OAI210     m0615(.A0(mai_mai_n643_), .A1(mai_mai_n638_), .B0(mai_mai_n503_), .Y(mai_mai_n644_));
  AOI210     m0616(.A0(mai_mai_n637_), .A1(l), .B0(mai_mai_n644_), .Y(mai_mai_n645_));
  NO2        m0617(.A(j), .B(i), .Y(mai_mai_n646_));
  NA3        m0618(.A(mai_mai_n646_), .B(mai_mai_n68_), .C(l), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n646_), .B(mai_mai_n33_), .Y(mai_mai_n648_));
  INV        m0620(.A(mai_mai_n360_), .Y(mai_mai_n649_));
  OA220      m0621(.A0(mai_mai_n649_), .A1(mai_mai_n648_), .B0(mai_mai_n647_), .B1(mai_mai_n499_), .Y(mai_mai_n650_));
  NO3        m0622(.A(mai_mai_n126_), .B(mai_mai_n46_), .C(mai_mai_n93_), .Y(mai_mai_n651_));
  NO3        m0623(.A(mai_mai_n464_), .B(mai_mai_n125_), .C(mai_mai_n63_), .Y(mai_mai_n652_));
  NO2        m0624(.A(mai_mai_n410_), .B(mai_mai_n375_), .Y(mai_mai_n653_));
  OAI210     m0625(.A0(mai_mai_n652_), .A1(mai_mai_n651_), .B0(mai_mai_n653_), .Y(mai_mai_n654_));
  INV        m0626(.A(mai_mai_n654_), .Y(mai_mai_n655_));
  NA2        m0627(.A(k), .B(j), .Y(mai_mai_n656_));
  NO3        m0628(.A(mai_mai_n150_), .B(mai_mai_n334_), .C(mai_mai_n95_), .Y(mai_mai_n657_));
  NA2        m0629(.A(mai_mai_n657_), .B(mai_mai_n214_), .Y(mai_mai_n658_));
  NA2        m0630(.A(mai_mai_n77_), .B(mai_mai_n70_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n659_), .B(mai_mai_n658_), .Y(mai_mai_n660_));
  NO2        m0632(.A(mai_mai_n264_), .B(mai_mai_n114_), .Y(mai_mai_n661_));
  NA2        m0633(.A(mai_mai_n661_), .B(mai_mai_n529_), .Y(mai_mai_n662_));
  NO2        m0634(.A(mai_mai_n622_), .B(mai_mai_n75_), .Y(mai_mai_n663_));
  NO2        m0635(.A(mai_mai_n500_), .B(mai_mai_n99_), .Y(mai_mai_n664_));
  OAI210     m0636(.A0(mai_mai_n664_), .A1(mai_mai_n653_), .B0(mai_mai_n578_), .Y(mai_mai_n665_));
  NA2        m0637(.A(mai_mai_n665_), .B(mai_mai_n662_), .Y(mai_mai_n666_));
  OR3        m0638(.A(mai_mai_n666_), .B(mai_mai_n660_), .C(mai_mai_n655_), .Y(mai_mai_n667_));
  NO3        m0639(.A(mai_mai_n370_), .B(j), .C(f), .Y(mai_mai_n668_));
  OAI220     m0640(.A0(mai_mai_n603_), .A1(mai_mai_n598_), .B0(mai_mai_n291_), .B1(mai_mai_n37_), .Y(mai_mai_n669_));
  AOI210     m0641(.A0(mai_mai_n668_), .A1(mai_mai_n226_), .B0(mai_mai_n669_), .Y(mai_mai_n670_));
  NA3        m0642(.A(mai_mai_n467_), .B(mai_mai_n257_), .C(h), .Y(mai_mai_n671_));
  NOi21      m0643(.An(mai_mai_n578_), .B(mai_mai_n671_), .Y(mai_mai_n672_));
  OAI220     m0644(.A0(mai_mai_n671_), .A1(mai_mai_n513_), .B0(mai_mai_n647_), .B1(mai_mai_n572_), .Y(mai_mai_n673_));
  INV        m0645(.A(mai_mai_n673_), .Y(mai_mai_n674_));
  NAi31      m0646(.An(mai_mai_n672_), .B(mai_mai_n674_), .C(mai_mai_n670_), .Y(mai_mai_n675_));
  BUFFER     m0647(.A(mai_mai_n663_), .Y(mai_mai_n676_));
  AOI220     m0648(.A0(mai_mai_n676_), .A1(mai_mai_n205_), .B0(mai_mai_n653_), .B1(mai_mai_n540_), .Y(mai_mai_n677_));
  OAI210     m0649(.A0(mai_mai_n622_), .A1(mai_mai_n562_), .B0(mai_mai_n441_), .Y(mai_mai_n678_));
  NA3        m0650(.A(mai_mai_n217_), .B(mai_mai_n51_), .C(b), .Y(mai_mai_n679_));
  AOI220     m0651(.A0(mai_mai_n512_), .A1(mai_mai_n29_), .B0(mai_mai_n395_), .B1(mai_mai_n70_), .Y(mai_mai_n680_));
  NA2        m0652(.A(mai_mai_n680_), .B(mai_mai_n679_), .Y(mai_mai_n681_));
  NA2        m0653(.A(mai_mai_n681_), .B(mai_mai_n678_), .Y(mai_mai_n682_));
  NA2        m0654(.A(mai_mai_n682_), .B(mai_mai_n677_), .Y(mai_mai_n683_));
  NOi41      m0655(.An(mai_mai_n650_), .B(mai_mai_n683_), .C(mai_mai_n675_), .D(mai_mai_n667_), .Y(mai_mai_n684_));
  OR3        m0656(.A(mai_mai_n603_), .B(mai_mai_n202_), .C(g), .Y(mai_mai_n685_));
  INV        m0657(.A(mai_mai_n44_), .Y(mai_mai_n686_));
  NO3        m0658(.A(mai_mai_n686_), .B(mai_mai_n648_), .C(mai_mai_n242_), .Y(mai_mai_n687_));
  NO3        m0659(.A(mai_mai_n448_), .B(mai_mai_n78_), .C(h), .Y(mai_mai_n688_));
  AOI210     m0660(.A0(mai_mai_n688_), .A1(mai_mai_n602_), .B0(mai_mai_n687_), .Y(mai_mai_n689_));
  NA3        m0661(.A(mai_mai_n689_), .B(mai_mai_n685_), .C(mai_mai_n345_), .Y(mai_mai_n690_));
  OR2        m0662(.A(mai_mai_n562_), .B(mai_mai_n76_), .Y(mai_mai_n691_));
  NOi31      m0663(.An(b), .B(d), .C(a), .Y(mai_mai_n692_));
  NO2        m0664(.A(mai_mai_n692_), .B(mai_mai_n510_), .Y(mai_mai_n693_));
  NO2        m0665(.A(mai_mai_n693_), .B(n), .Y(mai_mai_n694_));
  NOi21      m0666(.An(mai_mai_n680_), .B(mai_mai_n694_), .Y(mai_mai_n695_));
  NO2        m0667(.A(mai_mai_n695_), .B(mai_mai_n691_), .Y(mai_mai_n696_));
  NO3        m0668(.A(mai_mai_n528_), .B(mai_mai_n287_), .C(mai_mai_n99_), .Y(mai_mai_n697_));
  NOi21      m0669(.An(mai_mai_n697_), .B(mai_mai_n135_), .Y(mai_mai_n698_));
  INV        m0670(.A(mai_mai_n698_), .Y(mai_mai_n699_));
  OAI210     m0671(.A0(mai_mai_n603_), .A1(mai_mai_n336_), .B0(mai_mai_n699_), .Y(mai_mai_n700_));
  NO2        m0672(.A(mai_mai_n586_), .B(n), .Y(mai_mai_n701_));
  AOI220     m0673(.A0(mai_mai_n661_), .A1(mai_mai_n569_), .B0(mai_mai_n701_), .B1(mai_mai_n597_), .Y(mai_mai_n702_));
  NA2        m0674(.A(mai_mai_n80_), .B(mai_mai_n1243_), .Y(mai_mai_n703_));
  NA2        m0675(.A(mai_mai_n102_), .B(mai_mai_n70_), .Y(mai_mai_n704_));
  AOI210     m0676(.A0(mai_mai_n364_), .A1(mai_mai_n356_), .B0(mai_mai_n704_), .Y(mai_mai_n705_));
  NAi21      m0677(.An(mai_mai_n705_), .B(mai_mai_n703_), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n620_), .B(mai_mai_n34_), .Y(mai_mai_n707_));
  NAi21      m0679(.An(mai_mai_n626_), .B(mai_mai_n371_), .Y(mai_mai_n708_));
  NO2        m0680(.A(mai_mai_n238_), .B(i), .Y(mai_mai_n709_));
  NA2        m0681(.A(mai_mai_n607_), .B(mai_mai_n301_), .Y(mai_mai_n710_));
  OAI210     m0682(.A0(mai_mai_n506_), .A1(mai_mai_n505_), .B0(mai_mai_n312_), .Y(mai_mai_n711_));
  AN3        m0683(.A(mai_mai_n711_), .B(mai_mai_n710_), .C(mai_mai_n708_), .Y(mai_mai_n712_));
  NAi41      m0684(.An(mai_mai_n706_), .B(mai_mai_n712_), .C(mai_mai_n707_), .D(mai_mai_n702_), .Y(mai_mai_n713_));
  NO4        m0685(.A(mai_mai_n713_), .B(mai_mai_n700_), .C(mai_mai_n696_), .D(mai_mai_n690_), .Y(mai_mai_n714_));
  NA4        m0686(.A(mai_mai_n714_), .B(mai_mai_n684_), .C(mai_mai_n645_), .D(mai_mai_n631_), .Y(mai09));
  INV        m0687(.A(mai_mai_n103_), .Y(mai_mai_n716_));
  NA2        m0688(.A(f), .B(e), .Y(mai_mai_n717_));
  NA4        m0689(.A(mai_mai_n273_), .B(mai_mai_n401_), .C(mai_mai_n229_), .D(mai_mai_n101_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n718_), .B(g), .Y(mai_mai_n719_));
  INV        m0691(.A(mai_mai_n717_), .Y(mai_mai_n720_));
  NA2        m0692(.A(mai_mai_n381_), .B(e), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n720_), .B(mai_mai_n716_), .Y(mai_mai_n722_));
  NO2        m0694(.A(mai_mai_n178_), .B(mai_mai_n183_), .Y(mai_mai_n723_));
  NA3        m0695(.A(m), .B(l), .C(i), .Y(mai_mai_n724_));
  OAI220     m0696(.A0(mai_mai_n500_), .A1(mai_mai_n724_), .B0(mai_mai_n305_), .B1(mai_mai_n449_), .Y(mai_mai_n725_));
  NA4        m0697(.A(mai_mai_n73_), .B(mai_mai_n72_), .C(g), .D(f), .Y(mai_mai_n726_));
  NAi31      m0698(.An(mai_mai_n725_), .B(mai_mai_n726_), .C(mai_mai_n376_), .Y(mai_mai_n727_));
  OR2        m0699(.A(mai_mai_n727_), .B(mai_mai_n723_), .Y(mai_mai_n728_));
  NA3        m0700(.A(mai_mai_n691_), .B(mai_mai_n482_), .C(mai_mai_n441_), .Y(mai_mai_n729_));
  OA210      m0701(.A0(mai_mai_n729_), .A1(mai_mai_n728_), .B0(mai_mai_n694_), .Y(mai_mai_n730_));
  INV        m0702(.A(mai_mai_n296_), .Y(mai_mai_n731_));
  INV        m0703(.A(mai_mai_n106_), .Y(mai_mai_n732_));
  NA2        m0704(.A(mai_mai_n679_), .B(mai_mai_n291_), .Y(mai_mai_n733_));
  NA2        m0705(.A(mai_mai_n298_), .B(mai_mai_n299_), .Y(mai_mai_n734_));
  OAI210     m0706(.A0(mai_mai_n178_), .A1(mai_mai_n183_), .B0(mai_mai_n734_), .Y(mai_mai_n735_));
  NA2        m0707(.A(mai_mai_n735_), .B(mai_mai_n733_), .Y(mai_mai_n736_));
  NA2        m0708(.A(mai_mai_n144_), .B(mai_mai_n97_), .Y(mai_mai_n737_));
  NA2        m0709(.A(mai_mai_n737_), .B(mai_mai_n596_), .Y(mai_mai_n738_));
  NA3        m0710(.A(mai_mai_n738_), .B(mai_mai_n163_), .C(mai_mai_n31_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n739_), .B(mai_mai_n736_), .Y(mai_mai_n740_));
  NO2        m0712(.A(mai_mai_n496_), .B(mai_mai_n423_), .Y(mai_mai_n741_));
  NA2        m0713(.A(mai_mai_n741_), .B(mai_mai_n163_), .Y(mai_mai_n742_));
  NOi21      m0714(.An(f), .B(d), .Y(mai_mai_n743_));
  NA2        m0715(.A(mai_mai_n743_), .B(m), .Y(mai_mai_n744_));
  NO2        m0716(.A(mai_mai_n744_), .B(g), .Y(mai_mai_n745_));
  NOi32      m0717(.An(g), .Bn(f), .C(d), .Y(mai_mai_n746_));
  NA3        m0718(.A(mai_mai_n403_), .B(f), .C(mai_mai_n70_), .Y(mai_mai_n747_));
  NAi21      m0719(.An(mai_mai_n415_), .B(mai_mai_n742_), .Y(mai_mai_n748_));
  NO2        m0720(.A(mai_mai_n556_), .B(mai_mai_n287_), .Y(mai_mai_n749_));
  AN2        m0721(.A(mai_mai_n749_), .B(mai_mai_n582_), .Y(mai_mai_n750_));
  INV        m0722(.A(mai_mai_n750_), .Y(mai_mai_n751_));
  NA2        m0723(.A(mai_mai_n510_), .B(mai_mai_n70_), .Y(mai_mai_n752_));
  NO2        m0724(.A(mai_mai_n734_), .B(mai_mai_n752_), .Y(mai_mai_n753_));
  NA3        m0725(.A(mai_mai_n134_), .B(mai_mai_n91_), .C(mai_mai_n90_), .Y(mai_mai_n754_));
  OAI220     m0726(.A0(mai_mai_n747_), .A1(mai_mai_n1242_), .B0(mai_mai_n296_), .B1(mai_mai_n754_), .Y(mai_mai_n755_));
  NOi31      m0727(.An(mai_mai_n194_), .B(mai_mai_n755_), .C(mai_mai_n753_), .Y(mai_mai_n756_));
  NA2        m0728(.A(c), .B(mai_mai_n98_), .Y(mai_mai_n757_));
  INV        m0729(.A(mai_mai_n757_), .Y(mai_mai_n758_));
  NA2        m0730(.A(mai_mai_n758_), .B(mai_mai_n432_), .Y(mai_mai_n759_));
  OR2        m0731(.A(mai_mai_n562_), .B(mai_mai_n461_), .Y(mai_mai_n760_));
  INV        m0732(.A(mai_mai_n760_), .Y(mai_mai_n761_));
  NA2        m0733(.A(mai_mai_n693_), .B(mai_mai_n94_), .Y(mai_mai_n762_));
  NA2        m0734(.A(mai_mai_n762_), .B(mai_mai_n761_), .Y(mai_mai_n763_));
  NA4        m0735(.A(mai_mai_n763_), .B(mai_mai_n759_), .C(mai_mai_n756_), .D(mai_mai_n751_), .Y(mai_mai_n764_));
  NO4        m0736(.A(mai_mai_n764_), .B(mai_mai_n748_), .C(mai_mai_n740_), .D(mai_mai_n730_), .Y(mai_mai_n765_));
  NO2        m0737(.A(mai_mai_n291_), .B(mai_mai_n726_), .Y(mai_mai_n766_));
  NO2        m0738(.A(mai_mai_n201_), .B(mai_mai_n195_), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n767_), .B(mai_mai_n198_), .Y(mai_mai_n768_));
  INV        m0740(.A(mai_mai_n768_), .Y(mai_mai_n769_));
  NA2        m0741(.A(e), .B(d), .Y(mai_mai_n770_));
  OAI220     m0742(.A0(mai_mai_n770_), .A1(c), .B0(mai_mai_n283_), .B1(d), .Y(mai_mai_n771_));
  NA3        m0743(.A(mai_mai_n771_), .B(mai_mai_n390_), .C(mai_mai_n431_), .Y(mai_mai_n772_));
  NO2        m0744(.A(mai_mai_n437_), .B(mai_mai_n201_), .Y(mai_mai_n773_));
  INV        m0745(.A(mai_mai_n773_), .Y(mai_mai_n774_));
  NA3        m0746(.A(mai_mai_n143_), .B(mai_mai_n71_), .C(mai_mai_n34_), .Y(mai_mai_n775_));
  NA3        m0747(.A(mai_mai_n775_), .B(mai_mai_n774_), .C(mai_mai_n772_), .Y(mai_mai_n776_));
  NO3        m0748(.A(mai_mai_n776_), .B(mai_mai_n769_), .C(mai_mai_n766_), .Y(mai_mai_n777_));
  NA2        m0749(.A(mai_mai_n731_), .B(mai_mai_n31_), .Y(mai_mai_n778_));
  OR2        m0750(.A(mai_mai_n778_), .B(mai_mai_n187_), .Y(mai_mai_n779_));
  OAI220     m0751(.A0(mai_mai_n528_), .A1(mai_mai_n52_), .B0(mai_mai_n266_), .B1(j), .Y(mai_mai_n780_));
  AOI220     m0752(.A0(mai_mai_n780_), .A1(mai_mai_n749_), .B0(mai_mai_n520_), .B1(mai_mai_n527_), .Y(mai_mai_n781_));
  OAI210     m0753(.A0(mai_mai_n721_), .A1(mai_mai_n147_), .B0(mai_mai_n781_), .Y(mai_mai_n782_));
  AN2        m0754(.A(mai_mai_n733_), .B(mai_mai_n725_), .Y(mai_mai_n783_));
  NOi21      m0755(.An(mai_mai_n465_), .B(mai_mai_n744_), .Y(mai_mai_n784_));
  NO3        m0756(.A(mai_mai_n784_), .B(mai_mai_n783_), .C(mai_mai_n782_), .Y(mai_mai_n785_));
  AO220      m0757(.A0(mai_mai_n390_), .A1(mai_mai_n640_), .B0(mai_mai_n152_), .B1(f), .Y(mai_mai_n786_));
  NA2        m0758(.A(mai_mai_n786_), .B(mai_mai_n771_), .Y(mai_mai_n787_));
  NO2        m0759(.A(mai_mai_n375_), .B(mai_mai_n61_), .Y(mai_mai_n788_));
  OAI210     m0760(.A0(mai_mai_n729_), .A1(mai_mai_n788_), .B0(mai_mai_n602_), .Y(mai_mai_n789_));
  AN4        m0761(.A(mai_mai_n789_), .B(mai_mai_n787_), .C(mai_mai_n785_), .D(mai_mai_n779_), .Y(mai_mai_n790_));
  NA4        m0762(.A(mai_mai_n790_), .B(mai_mai_n777_), .C(mai_mai_n765_), .D(mai_mai_n722_), .Y(mai12));
  NO4        m0763(.A(mai_mai_n380_), .B(mai_mai_n220_), .C(mai_mai_n493_), .D(mai_mai_n184_), .Y(mai_mai_n792_));
  NA2        m0764(.A(mai_mai_n465_), .B(mai_mai_n788_), .Y(mai_mai_n793_));
  NO2        m0765(.A(mai_mai_n388_), .B(mai_mai_n98_), .Y(mai_mai_n794_));
  NO2        m0766(.A(mai_mai_n732_), .B(mai_mai_n305_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n562_), .B(mai_mai_n324_), .Y(mai_mai_n796_));
  NA2        m0768(.A(mai_mai_n795_), .B(mai_mai_n794_), .Y(mai_mai_n797_));
  NA3        m0769(.A(mai_mai_n797_), .B(mai_mai_n793_), .C(mai_mai_n379_), .Y(mai_mai_n798_));
  AOI210     m0770(.A0(mai_mai_n203_), .A1(mai_mai_n295_), .B0(mai_mai_n175_), .Y(mai_mai_n799_));
  OR2        m0771(.A(mai_mai_n799_), .B(mai_mai_n792_), .Y(mai_mai_n800_));
  NA2        m0772(.A(mai_mai_n800_), .B(mai_mai_n344_), .Y(mai_mai_n801_));
  NO2        m0773(.A(mai_mai_n544_), .B(mai_mai_n230_), .Y(mai_mai_n802_));
  NO2        m0774(.A(mai_mai_n500_), .B(mai_mai_n724_), .Y(mai_mai_n803_));
  AOI220     m0775(.A0(mai_mai_n803_), .A1(mai_mai_n480_), .B0(mai_mai_n1243_), .B1(mai_mai_n802_), .Y(mai_mai_n804_));
  NA2        m0776(.A(mai_mai_n804_), .B(mai_mai_n801_), .Y(mai_mai_n805_));
  NO3        m0777(.A(mai_mai_n567_), .B(mai_mai_n76_), .C(mai_mai_n43_), .Y(mai_mai_n806_));
  NO3        m0778(.A(mai_mai_n806_), .B(mai_mai_n805_), .C(mai_mai_n798_), .Y(mai_mai_n807_));
  NO2        m0779(.A(mai_mai_n316_), .B(mai_mai_n315_), .Y(mai_mai_n808_));
  NOi21      m0780(.An(mai_mai_n34_), .B(mai_mai_n556_), .Y(mai_mai_n809_));
  NA2        m0781(.A(mai_mai_n1239_), .B(mai_mai_n808_), .Y(mai_mai_n810_));
  NA2        m0782(.A(mai_mai_n218_), .B(mai_mai_n810_), .Y(mai_mai_n811_));
  NO3        m0783(.A(mai_mai_n704_), .B(mai_mai_n74_), .C(mai_mai_n348_), .Y(mai_mai_n812_));
  NO2        m0784(.A(mai_mai_n46_), .B(mai_mai_n43_), .Y(mai_mai_n813_));
  INV        m0785(.A(mai_mai_n314_), .Y(mai_mai_n814_));
  NO2        m0786(.A(mai_mai_n814_), .B(mai_mai_n811_), .Y(mai_mai_n815_));
  NA2        m0787(.A(mai_mai_n472_), .B(mai_mai_n328_), .Y(mai_mai_n816_));
  NO2        m0788(.A(mai_mai_n1236_), .B(mai_mai_n291_), .Y(mai_mai_n817_));
  NO2        m0789(.A(mai_mai_n562_), .B(mai_mai_n423_), .Y(mai_mai_n818_));
  NA3        m0790(.A(mai_mai_n298_), .B(j), .C(i), .Y(mai_mai_n819_));
  INV        m0791(.A(mai_mai_n819_), .Y(mai_mai_n820_));
  OAI220     m0792(.A0(mai_mai_n820_), .A1(mai_mai_n818_), .B0(mai_mai_n578_), .B1(mai_mai_n652_), .Y(mai_mai_n821_));
  INV        m0793(.A(mai_mai_n96_), .Y(mai_mai_n822_));
  NA3        m0794(.A(j), .B(mai_mai_n68_), .C(i), .Y(mai_mai_n823_));
  OR2        m0795(.A(mai_mai_n823_), .B(mai_mai_n822_), .Y(mai_mai_n824_));
  NA3        m0796(.A(f), .B(mai_mai_n100_), .C(g), .Y(mai_mai_n825_));
  AOI210     m0797(.A0(mai_mai_n575_), .A1(mai_mai_n825_), .B0(m), .Y(mai_mai_n826_));
  OAI210     m0798(.A0(mai_mai_n826_), .A1(mai_mai_n795_), .B0(mai_mai_n284_), .Y(mai_mai_n827_));
  NA2        m0799(.A(mai_mai_n589_), .B(mai_mai_n752_), .Y(mai_mai_n828_));
  NA2        m0800(.A(mai_mai_n192_), .B(mai_mai_n66_), .Y(mai_mai_n829_));
  NA2        m0801(.A(mai_mai_n829_), .B(mai_mai_n823_), .Y(mai_mai_n830_));
  AOI220     m0802(.A0(mai_mai_n830_), .A1(mai_mai_n226_), .B0(mai_mai_n73_), .B1(mai_mai_n828_), .Y(mai_mai_n831_));
  NA4        m0803(.A(mai_mai_n831_), .B(mai_mai_n827_), .C(mai_mai_n824_), .D(mai_mai_n821_), .Y(mai_mai_n832_));
  NO2        m0804(.A(mai_mai_n324_), .B(mai_mai_n75_), .Y(mai_mai_n833_));
  OAI210     m0805(.A0(mai_mai_n833_), .A1(mai_mai_n802_), .B0(mai_mai_n205_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n566_), .B(mai_mai_n73_), .Y(mai_mai_n835_));
  NA2        m0807(.A(mai_mai_n835_), .B(mai_mai_n834_), .Y(mai_mai_n836_));
  OAI210     m0808(.A0(mai_mai_n73_), .A1(mai_mai_n803_), .B0(mai_mai_n463_), .Y(mai_mai_n837_));
  AOI210     m0809(.A0(mai_mai_n359_), .A1(mai_mai_n351_), .B0(mai_mai_n704_), .Y(mai_mai_n838_));
  OAI210     m0810(.A0(mai_mai_n316_), .A1(mai_mai_n315_), .B0(mai_mai_n92_), .Y(mai_mai_n839_));
  AOI210     m0811(.A0(mai_mai_n839_), .A1(mai_mai_n456_), .B0(mai_mai_n838_), .Y(mai_mai_n840_));
  NA2        m0812(.A(mai_mai_n826_), .B(mai_mai_n794_), .Y(mai_mai_n841_));
  NO2        m0813(.A(mai_mai_n46_), .B(mai_mai_n43_), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n842_), .B(mai_mai_n531_), .Y(mai_mai_n843_));
  NA4        m0815(.A(mai_mai_n843_), .B(mai_mai_n841_), .C(mai_mai_n840_), .D(mai_mai_n837_), .Y(mai_mai_n844_));
  NO4        m0816(.A(mai_mai_n844_), .B(mai_mai_n836_), .C(mai_mai_n832_), .D(mai_mai_n817_), .Y(mai_mai_n845_));
  NAi31      m0817(.An(mai_mai_n119_), .B(mai_mai_n360_), .C(n), .Y(mai_mai_n846_));
  NO3        m0818(.A(mai_mai_n238_), .B(mai_mai_n119_), .C(mai_mai_n348_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n847_), .B(mai_mai_n424_), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n418_), .B(i), .Y(mai_mai_n849_));
  NA2        m0821(.A(mai_mai_n849_), .B(mai_mai_n848_), .Y(mai_mai_n850_));
  NA2        m0822(.A(mai_mai_n201_), .B(mai_mai_n148_), .Y(mai_mai_n851_));
  OAI220     m0823(.A0(mai_mai_n846_), .A1(mai_mai_n203_), .B0(mai_mai_n819_), .B1(mai_mai_n511_), .Y(mai_mai_n852_));
  NO2        m0824(.A(mai_mai_n464_), .B(mai_mai_n125_), .Y(mai_mai_n853_));
  OAI210     m0825(.A0(mai_mai_n853_), .A1(mai_mai_n447_), .B0(mai_mai_n325_), .Y(mai_mai_n854_));
  OAI220     m0826(.A0(mai_mai_n796_), .A1(mai_mai_n803_), .B0(mai_mai_n465_), .B1(mai_mai_n368_), .Y(mai_mai_n855_));
  NA2        m0827(.A(mai_mai_n855_), .B(mai_mai_n854_), .Y(mai_mai_n856_));
  OAI210     m0828(.A0(mai_mai_n799_), .A1(mai_mai_n792_), .B0(mai_mai_n851_), .Y(mai_mai_n857_));
  NA3        m0829(.A(mai_mai_n816_), .B(mai_mai_n412_), .C(mai_mai_n44_), .Y(mai_mai_n858_));
  NA3        m0830(.A(mai_mai_n858_), .B(mai_mai_n857_), .C(mai_mai_n239_), .Y(mai_mai_n859_));
  OR3        m0831(.A(mai_mai_n859_), .B(mai_mai_n856_), .C(mai_mai_n852_), .Y(mai_mai_n860_));
  NO3        m0832(.A(mai_mai_n860_), .B(mai_mai_n407_), .C(mai_mai_n850_), .Y(mai_mai_n861_));
  NA4        m0833(.A(mai_mai_n861_), .B(mai_mai_n845_), .C(mai_mai_n815_), .D(mai_mai_n807_), .Y(mai13));
  NA2        m0834(.A(mai_mai_n422_), .B(f), .Y(mai_mai_n863_));
  NO3        m0835(.A(mai_mai_n863_), .B(j), .C(mai_mai_n494_), .Y(mai_mai_n864_));
  NO3        m0836(.A(mai_mai_n60_), .B(mai_mai_n863_), .C(g), .Y(mai_mai_n865_));
  NA2        m0837(.A(mai_mai_n118_), .B(mai_mai_n43_), .Y(mai_mai_n866_));
  NO4        m0838(.A(mai_mai_n866_), .B(c), .C(mai_mai_n500_), .D(mai_mai_n271_), .Y(mai_mai_n867_));
  NA2        m0839(.A(c), .B(mai_mai_n98_), .Y(mai_mai_n868_));
  NO4        m0840(.A(mai_mai_n868_), .B(f), .C(mai_mai_n153_), .D(mai_mai_n144_), .Y(mai_mai_n869_));
  NO3        m0841(.A(mai_mai_n866_), .B(mai_mai_n496_), .C(mai_mai_n271_), .Y(mai_mai_n870_));
  OR2        m0842(.A(mai_mai_n869_), .B(mai_mai_n870_), .Y(mai_mai_n871_));
  OR4        m0843(.A(mai_mai_n871_), .B(mai_mai_n867_), .C(mai_mai_n865_), .D(mai_mai_n864_), .Y(mai_mai_n872_));
  NAi32      m0844(.An(f), .Bn(e), .C(c), .Y(mai_mai_n873_));
  OR3        m0845(.A(mai_mai_n195_), .B(mai_mai_n153_), .C(mai_mai_n144_), .Y(mai_mai_n874_));
  NO2        m0846(.A(mai_mai_n874_), .B(mai_mai_n873_), .Y(mai_mai_n875_));
  NO2        m0847(.A(e), .B(mai_mai_n271_), .Y(mai_mai_n876_));
  NA2        m0848(.A(mai_mai_n533_), .B(mai_mai_n1231_), .Y(mai_mai_n877_));
  NOi21      m0849(.An(mai_mai_n876_), .B(mai_mai_n877_), .Y(mai_mai_n878_));
  NO2        m0850(.A(mai_mai_n656_), .B(mai_mai_n95_), .Y(mai_mai_n879_));
  NOi41      m0851(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n880_));
  NA2        m0852(.A(mai_mai_n880_), .B(mai_mai_n879_), .Y(mai_mai_n881_));
  NO2        m0853(.A(mai_mai_n881_), .B(mai_mai_n873_), .Y(mai_mai_n882_));
  NA3        m0854(.A(k), .B(j), .C(i), .Y(mai_mai_n883_));
  NO2        m0855(.A(mai_mai_n271_), .B(mai_mai_n75_), .Y(mai_mai_n884_));
  BUFFER     m0856(.A(mai_mai_n884_), .Y(mai_mai_n885_));
  OR4        m0857(.A(mai_mai_n885_), .B(mai_mai_n882_), .C(mai_mai_n878_), .D(mai_mai_n875_), .Y(mai_mai_n886_));
  NA2        m0858(.A(mai_mai_n397_), .B(mai_mai_n293_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n887_), .B(mai_mai_n877_), .Y(mai_mai_n888_));
  NO3        m0860(.A(mai_mai_n887_), .B(mai_mai_n496_), .C(mai_mai_n387_), .Y(mai_mai_n889_));
  NO2        m0861(.A(f), .B(c), .Y(mai_mai_n890_));
  NOi21      m0862(.An(mai_mai_n890_), .B(mai_mai_n380_), .Y(mai_mai_n891_));
  INV        m0863(.A(mai_mai_n891_), .Y(mai_mai_n892_));
  OR2        m0864(.A(k), .B(i), .Y(mai_mai_n893_));
  NO3        m0865(.A(mai_mai_n893_), .B(mai_mai_n210_), .C(l), .Y(mai_mai_n894_));
  NOi21      m0866(.An(mai_mai_n894_), .B(j), .Y(mai_mai_n895_));
  OR3        m0867(.A(mai_mai_n895_), .B(mai_mai_n889_), .C(mai_mai_n888_), .Y(mai_mai_n896_));
  OR3        m0868(.A(mai_mai_n896_), .B(mai_mai_n886_), .C(mai_mai_n872_), .Y(mai02));
  OR2        m0869(.A(l), .B(k), .Y(mai_mai_n898_));
  OR3        m0870(.A(h), .B(g), .C(f), .Y(mai_mai_n899_));
  NO4        m0871(.A(n), .B(mai_mai_n899_), .C(mai_mai_n898_), .D(e), .Y(mai_mai_n900_));
  NO2        m0872(.A(mai_mai_n884_), .B(mai_mai_n867_), .Y(mai_mai_n901_));
  AN3        m0873(.A(g), .B(f), .C(c), .Y(mai_mai_n902_));
  NA3        m0874(.A(mai_mai_n902_), .B(mai_mai_n397_), .C(h), .Y(mai_mai_n903_));
  OR2        m0875(.A(mai_mai_n271_), .B(mai_mai_n903_), .Y(mai_mai_n904_));
  NO3        m0876(.A(mai_mai_n887_), .B(mai_mai_n866_), .C(mai_mai_n496_), .Y(mai_mai_n905_));
  NO2        m0877(.A(mai_mai_n905_), .B(mai_mai_n875_), .Y(mai_mai_n906_));
  NA3        m0878(.A(l), .B(k), .C(j), .Y(mai_mai_n907_));
  NA2        m0879(.A(i), .B(h), .Y(mai_mai_n908_));
  NO3        m0880(.A(mai_mai_n908_), .B(mai_mai_n907_), .C(mai_mai_n111_), .Y(mai_mai_n909_));
  NO3        m0881(.A(mai_mai_n120_), .B(mai_mai_n248_), .C(mai_mai_n184_), .Y(mai_mai_n910_));
  AOI210     m0882(.A0(mai_mai_n910_), .A1(mai_mai_n909_), .B0(mai_mai_n878_), .Y(mai_mai_n911_));
  NA3        m0883(.A(c), .B(b), .C(a), .Y(mai_mai_n912_));
  NO3        m0884(.A(mai_mai_n912_), .B(mai_mai_n770_), .C(mai_mai_n183_), .Y(mai_mai_n913_));
  NO3        m0885(.A(mai_mai_n266_), .B(mai_mai_n46_), .C(mai_mai_n95_), .Y(mai_mai_n914_));
  AOI210     m0886(.A0(mai_mai_n914_), .A1(mai_mai_n913_), .B0(mai_mai_n888_), .Y(mai_mai_n915_));
  AN4        m0887(.A(mai_mai_n915_), .B(mai_mai_n911_), .C(mai_mai_n906_), .D(mai_mai_n904_), .Y(mai_mai_n916_));
  NA2        m0888(.A(mai_mai_n881_), .B(mai_mai_n874_), .Y(mai_mai_n917_));
  AOI210     m0889(.A0(mai_mai_n917_), .A1(c), .B0(mai_mai_n864_), .Y(mai_mai_n918_));
  NAi41      m0890(.An(mai_mai_n900_), .B(mai_mai_n918_), .C(mai_mai_n916_), .D(mai_mai_n901_), .Y(mai03));
  INV        m0891(.A(mai_mai_n317_), .Y(mai_mai_n920_));
  INV        m0892(.A(mai_mai_n589_), .Y(mai_mai_n921_));
  NOi31      m0893(.An(i), .B(k), .C(j), .Y(mai_mai_n922_));
  NA4        m0894(.A(mai_mai_n922_), .B(e), .C(mai_mai_n298_), .D(mai_mai_n293_), .Y(mai_mai_n923_));
  OAI210     m0895(.A0(mai_mai_n704_), .A1(mai_mai_n361_), .B0(mai_mai_n923_), .Y(mai_mai_n924_));
  NOi31      m0896(.An(m), .B(n), .C(f), .Y(mai_mai_n925_));
  NA2        m0897(.A(mai_mai_n925_), .B(mai_mai_n47_), .Y(mai_mai_n926_));
  NA2        m0898(.A(mai_mai_n431_), .B(l), .Y(mai_mai_n927_));
  NOi31      m0899(.An(mai_mai_n746_), .B(mai_mai_n1244_), .C(mai_mai_n927_), .Y(mai_mai_n928_));
  NO3        m0900(.A(mai_mai_n928_), .B(mai_mai_n924_), .C(mai_mai_n838_), .Y(mai_mai_n929_));
  NO2        m0901(.A(mai_mai_n248_), .B(a), .Y(mai_mai_n930_));
  INV        m0902(.A(mai_mai_n867_), .Y(mai_mai_n931_));
  NO2        m0903(.A(mai_mai_n908_), .B(mai_mai_n410_), .Y(mai_mai_n932_));
  NO2        m0904(.A(mai_mai_n72_), .B(g), .Y(mai_mai_n933_));
  NO2        m0905(.A(mai_mai_n932_), .B(mai_mai_n894_), .Y(mai_mai_n934_));
  OR2        m0906(.A(mai_mai_n934_), .B(mai_mai_n892_), .Y(mai_mai_n935_));
  NA3        m0907(.A(mai_mai_n935_), .B(mai_mai_n931_), .C(mai_mai_n929_), .Y(mai_mai_n936_));
  NO4        m0908(.A(mai_mai_n936_), .B(mai_mai_n921_), .C(mai_mai_n706_), .D(mai_mai_n479_), .Y(mai_mai_n937_));
  NA2        m0909(.A(c), .B(b), .Y(mai_mai_n938_));
  NO2        m0910(.A(mai_mai_n601_), .B(mai_mai_n938_), .Y(mai_mai_n939_));
  OAI210     m0911(.A0(mai_mai_n744_), .A1(mai_mai_n719_), .B0(mai_mai_n354_), .Y(mai_mai_n940_));
  OAI210     m0912(.A0(mai_mai_n940_), .A1(mai_mai_n745_), .B0(mai_mai_n939_), .Y(mai_mai_n941_));
  NAi21      m0913(.An(mai_mai_n362_), .B(mai_mai_n939_), .Y(mai_mai_n942_));
  OAI210     m0914(.A0(mai_mai_n1246_), .A1(mai_mai_n38_), .B0(mai_mai_n930_), .Y(mai_mai_n943_));
  NA2        m0915(.A(mai_mai_n943_), .B(mai_mai_n942_), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n229_), .B(mai_mai_n101_), .Y(mai_mai_n945_));
  OAI210     m0917(.A0(mai_mai_n945_), .A1(mai_mai_n252_), .B0(g), .Y(mai_mai_n946_));
  NO2        m0918(.A(mai_mai_n946_), .B(f), .Y(mai_mai_n947_));
  AOI210     m0919(.A0(mai_mai_n947_), .A1(mai_mai_n96_), .B0(mai_mai_n944_), .Y(mai_mai_n948_));
  INV        m0920(.A(mai_mai_n398_), .Y(mai_mai_n949_));
  NO2        m0921(.A(mai_mai_n158_), .B(mai_mai_n204_), .Y(mai_mai_n950_));
  NA2        m0922(.A(mai_mai_n950_), .B(m), .Y(mai_mai_n951_));
  AOI210     m0923(.A0(mai_mai_n1233_), .A1(mai_mai_n949_), .B0(mai_mai_n951_), .Y(mai_mai_n952_));
  NA2        m0924(.A(mai_mai_n475_), .B(mai_mai_n350_), .Y(mai_mai_n953_));
  NA2        m0925(.A(mai_mai_n133_), .B(mai_mai_n33_), .Y(mai_mai_n954_));
  NO2        m0926(.A(mai_mai_n954_), .B(mai_mai_n184_), .Y(mai_mai_n955_));
  NA2        m0927(.A(mai_mai_n955_), .B(mai_mai_n1245_), .Y(mai_mai_n956_));
  NO2        m0928(.A(mai_mai_n319_), .B(mai_mai_n318_), .Y(mai_mai_n957_));
  AOI210     m0929(.A0(mai_mai_n950_), .A1(mai_mai_n47_), .B0(mai_mai_n812_), .Y(mai_mai_n958_));
  NAi41      m0930(.An(mai_mai_n957_), .B(mai_mai_n958_), .C(mai_mai_n956_), .D(mai_mai_n953_), .Y(mai_mai_n959_));
  NO2        m0931(.A(mai_mai_n959_), .B(mai_mai_n952_), .Y(mai_mai_n960_));
  NA4        m0932(.A(mai_mai_n960_), .B(mai_mai_n948_), .C(mai_mai_n941_), .D(mai_mai_n937_), .Y(mai00));
  AOI210     m0933(.A0(mai_mai_n265_), .A1(mai_mai_n184_), .B0(mai_mai_n241_), .Y(mai_mai_n962_));
  NO2        m0934(.A(mai_mai_n962_), .B(mai_mai_n490_), .Y(mai_mai_n963_));
  INV        m0935(.A(mai_mai_n924_), .Y(mai_mai_n964_));
  NO2        m0936(.A(mai_mai_n812_), .B(mai_mai_n606_), .Y(mai_mai_n965_));
  NA3        m0937(.A(mai_mai_n965_), .B(mai_mai_n964_), .C(mai_mai_n840_), .Y(mai_mai_n966_));
  NO3        m0938(.A(mai_mai_n966_), .B(mai_mai_n963_), .C(mai_mai_n886_), .Y(mai_mai_n967_));
  NA3        m0939(.A(mai_mai_n143_), .B(mai_mai_n44_), .C(mai_mai_n43_), .Y(mai_mai_n968_));
  NA3        m0940(.A(d), .B(mai_mai_n49_), .C(b), .Y(mai_mai_n969_));
  NOi31      m0941(.An(n), .B(m), .C(i), .Y(mai_mai_n970_));
  NA3        m0942(.A(mai_mai_n970_), .B(mai_mai_n552_), .C(mai_mai_n47_), .Y(mai_mai_n971_));
  OAI210     m0943(.A0(mai_mai_n969_), .A1(mai_mai_n968_), .B0(mai_mai_n971_), .Y(mai_mai_n972_));
  NO3        m0944(.A(mai_mai_n972_), .B(mai_mai_n957_), .C(mai_mai_n784_), .Y(mai_mai_n973_));
  NO3        m0945(.A(mai_mai_n413_), .B(mai_mai_n306_), .C(mai_mai_n938_), .Y(mai_mai_n974_));
  OR2        m0946(.A(mai_mai_n331_), .B(mai_mai_n113_), .Y(mai_mai_n975_));
  NO2        m0947(.A(h), .B(g), .Y(mai_mai_n976_));
  NO2        m0948(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n977_));
  NA2        m0949(.A(mai_mai_n977_), .B(mai_mai_n456_), .Y(mai_mai_n978_));
  NA2        m0950(.A(mai_mai_n154_), .B(mai_mai_n124_), .Y(mai_mai_n979_));
  NA3        m0951(.A(mai_mai_n979_), .B(mai_mai_n978_), .C(mai_mai_n975_), .Y(mai_mai_n980_));
  NO3        m0952(.A(mai_mai_n980_), .B(mai_mai_n974_), .C(mai_mai_n234_), .Y(mai_mai_n981_));
  INV        m0953(.A(mai_mai_n282_), .Y(mai_mai_n982_));
  NA2        m0954(.A(mai_mai_n982_), .B(mai_mai_n129_), .Y(mai_mai_n983_));
  NA3        m0955(.A(mai_mai_n156_), .B(mai_mai_n95_), .C(g), .Y(mai_mai_n984_));
  NA2        m0956(.A(mai_mai_n397_), .B(f), .Y(mai_mai_n985_));
  NOi31      m0957(.An(mai_mai_n1240_), .B(mai_mai_n985_), .C(mai_mai_n984_), .Y(mai_mai_n986_));
  NAi31      m0958(.An(mai_mai_n159_), .B(mai_mai_n741_), .C(mai_mai_n397_), .Y(mai_mai_n987_));
  NAi21      m0959(.An(mai_mai_n986_), .B(mai_mai_n987_), .Y(mai_mai_n988_));
  INV        m0960(.A(mai_mai_n900_), .Y(mai_mai_n989_));
  NAi21      m0961(.An(mai_mai_n870_), .B(mai_mai_n989_), .Y(mai_mai_n990_));
  NO4        m0962(.A(mai_mai_n990_), .B(mai_mai_n988_), .C(mai_mai_n983_), .D(mai_mai_n440_), .Y(mai_mai_n991_));
  AN3        m0963(.A(mai_mai_n991_), .B(mai_mai_n981_), .C(mai_mai_n973_), .Y(mai_mai_n992_));
  NA2        m0964(.A(mai_mai_n456_), .B(mai_mai_n85_), .Y(mai_mai_n993_));
  NA3        m0965(.A(mai_mai_n476_), .B(mai_mai_n993_), .C(mai_mai_n208_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n920_), .B(mai_mai_n456_), .Y(mai_mai_n995_));
  NA2        m0967(.A(mai_mai_n995_), .B(mai_mai_n262_), .Y(mai_mai_n996_));
  INV        m0968(.A(mai_mai_n396_), .Y(mai_mai_n997_));
  AOI210     m0969(.A0(mai_mai_n475_), .A1(mai_mai_n350_), .B0(mai_mai_n997_), .Y(mai_mai_n998_));
  OR2        m0970(.A(mai_mai_n868_), .B(mai_mai_n193_), .Y(mai_mai_n999_));
  NO2        m0971(.A(mai_mai_n187_), .B(mai_mai_n184_), .Y(mai_mai_n1000_));
  NA2        m0972(.A(mai_mai_n731_), .B(mai_mai_n1000_), .Y(mai_mai_n1001_));
  NA3        m0973(.A(mai_mai_n1001_), .B(mai_mai_n999_), .C(mai_mai_n998_), .Y(mai_mai_n1002_));
  INV        m0974(.A(mai_mai_n705_), .Y(mai_mai_n1003_));
  AOI220     m0975(.A0(mai_mai_n809_), .A1(mai_mai_n489_), .B0(mai_mai_n552_), .B1(mai_mai_n211_), .Y(mai_mai_n1004_));
  NO2        m0976(.A(mai_mai_n59_), .B(h), .Y(mai_mai_n1005_));
  NO3        m0977(.A(mai_mai_n868_), .B(f), .C(mai_mai_n619_), .Y(mai_mai_n1006_));
  NO2        m0978(.A(mai_mai_n898_), .B(mai_mai_n111_), .Y(mai_mai_n1007_));
  AN2        m0979(.A(mai_mai_n1007_), .B(mai_mai_n910_), .Y(mai_mai_n1008_));
  OAI210     m0980(.A0(mai_mai_n1008_), .A1(mai_mai_n1006_), .B0(mai_mai_n1005_), .Y(mai_mai_n1009_));
  NA3        m0981(.A(mai_mai_n1009_), .B(mai_mai_n1004_), .C(mai_mai_n1003_), .Y(mai_mai_n1010_));
  NO4        m0982(.A(mai_mai_n1010_), .B(mai_mai_n1002_), .C(mai_mai_n996_), .D(mai_mai_n994_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(mai_mai_n720_), .B(mai_mai_n651_), .Y(mai_mai_n1012_));
  NA4        m0984(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .C(mai_mai_n992_), .D(mai_mai_n967_), .Y(mai01));
  NO2        m0985(.A(mai_mai_n687_), .B(mai_mai_n246_), .Y(mai_mai_n1014_));
  NA2        m0986(.A(mai_mai_n1014_), .B(mai_mai_n854_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(mai_mai_n781_), .B(mai_mai_n292_), .Y(mai_mai_n1016_));
  INV        m0988(.A(mai_mai_n100_), .Y(mai_mai_n1017_));
  OA220      m0989(.A0(mai_mai_n1017_), .A1(mai_mai_n495_), .B0(mai_mai_n564_), .B1(mai_mai_n317_), .Y(mai_mai_n1018_));
  NAi31      m0990(.An(mai_mai_n136_), .B(mai_mai_n1018_), .C(mai_mai_n768_), .Y(mai_mai_n1019_));
  NO3        m0991(.A(mai_mai_n672_), .B(mai_mai_n577_), .C(mai_mai_n434_), .Y(mai_mai_n1020_));
  OR2        m0992(.A(mai_mai_n169_), .B(mai_mai_n167_), .Y(mai_mai_n1021_));
  NA3        m0993(.A(mai_mai_n1021_), .B(mai_mai_n1020_), .C(mai_mai_n116_), .Y(mai_mai_n1022_));
  NO4        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1019_), .C(mai_mai_n1016_), .D(mai_mai_n1015_), .Y(mai_mai_n1023_));
  NA2        m0995(.A(mai_mai_n268_), .B(mai_mai_n453_), .Y(mai_mai_n1024_));
  NOi21      m0996(.An(mai_mai_n477_), .B(mai_mai_n493_), .Y(mai_mai_n1025_));
  INV        m0997(.A(mai_mai_n1025_), .Y(mai_mai_n1026_));
  AOI210     m0998(.A0(mai_mai_n178_), .A1(mai_mai_n74_), .B0(mai_mai_n183_), .Y(mai_mai_n1027_));
  OAI210     m0999(.A0(mai_mai_n694_), .A1(mai_mai_n368_), .B0(mai_mai_n1027_), .Y(mai_mai_n1028_));
  AN3        m1000(.A(m), .B(l), .C(k), .Y(mai_mai_n1029_));
  OAI210     m1001(.A0(mai_mai_n308_), .A1(mai_mai_n34_), .B0(mai_mai_n1029_), .Y(mai_mai_n1030_));
  NA2        m1002(.A(mai_mai_n177_), .B(mai_mai_n34_), .Y(mai_mai_n1031_));
  AO210      m1003(.A0(mai_mai_n1031_), .A1(mai_mai_n1030_), .B0(mai_mai_n291_), .Y(mai_mai_n1032_));
  NA4        m1004(.A(mai_mai_n1032_), .B(mai_mai_n1028_), .C(mai_mai_n1026_), .D(mai_mai_n1024_), .Y(mai_mai_n1033_));
  NA2        m1005(.A(mai_mai_n507_), .B(mai_mai_n100_), .Y(mai_mai_n1034_));
  OAI210     m1006(.A0(mai_mai_n1017_), .A1(mai_mai_n504_), .B0(mai_mai_n1034_), .Y(mai_mai_n1035_));
  NA2        m1007(.A(mai_mai_n245_), .B(mai_mai_n169_), .Y(mai_mai_n1036_));
  NA2        m1008(.A(mai_mai_n1036_), .B(mai_mai_n569_), .Y(mai_mai_n1037_));
  NO3        m1009(.A(mai_mai_n704_), .B(mai_mai_n178_), .C(mai_mai_n348_), .Y(mai_mai_n1038_));
  NO2        m1010(.A(mai_mai_n1038_), .B(mai_mai_n812_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n286_), .B(mai_mai_n578_), .Y(mai_mai_n1040_));
  NA4        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1039_), .C(mai_mai_n1037_), .D(mai_mai_n674_), .Y(mai_mai_n1041_));
  NO3        m1013(.A(mai_mai_n1041_), .B(mai_mai_n1035_), .C(mai_mai_n1033_), .Y(mai_mai_n1042_));
  NA3        m1014(.A(mai_mai_n512_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1043_));
  NO2        m1015(.A(mai_mai_n1043_), .B(mai_mai_n178_), .Y(mai_mai_n1044_));
  AOI210     m1016(.A0(mai_mai_n429_), .A1(c), .B0(mai_mai_n1044_), .Y(mai_mai_n1045_));
  INV        m1017(.A(mai_mai_n972_), .Y(mai_mai_n1046_));
  NA3        m1018(.A(mai_mai_n1046_), .B(mai_mai_n1045_), .C(mai_mai_n650_), .Y(mai_mai_n1047_));
  NA2        m1019(.A(mai_mai_n486_), .B(mai_mai_n484_), .Y(mai_mai_n1048_));
  NA2        m1020(.A(mai_mai_n1048_), .B(mai_mai_n574_), .Y(mai_mai_n1049_));
  NO2        m1021(.A(mai_mai_n317_), .B(mai_mai_n62_), .Y(mai_mai_n1050_));
  INV        m1022(.A(mai_mai_n1050_), .Y(mai_mai_n1051_));
  NA2        m1023(.A(mai_mai_n1051_), .B(mai_mai_n333_), .Y(mai_mai_n1052_));
  NO3        m1024(.A(mai_mai_n1052_), .B(mai_mai_n1049_), .C(mai_mai_n1047_), .Y(mai_mai_n1053_));
  AN2        m1025(.A(h), .B(mai_mai_n529_), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n1054_), .B(mai_mai_n297_), .Y(mai_mai_n1055_));
  INV        m1027(.A(mai_mai_n113_), .Y(mai_mai_n1056_));
  NO2        m1028(.A(mai_mai_n908_), .B(mai_mai_n153_), .Y(mai_mai_n1057_));
  NA2        m1029(.A(mai_mai_n1057_), .B(mai_mai_n1056_), .Y(mai_mai_n1058_));
  NA2        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1055_), .Y(mai_mai_n1059_));
  NO2        m1031(.A(mai_mai_n522_), .B(mai_mai_n521_), .Y(mai_mai_n1060_));
  NO4        m1032(.A(mai_mai_n908_), .B(mai_mai_n1060_), .C(mai_mai_n151_), .D(mai_mai_n72_), .Y(mai_mai_n1061_));
  NO3        m1033(.A(mai_mai_n1061_), .B(mai_mai_n1059_), .C(mai_mai_n543_), .Y(mai_mai_n1062_));
  NA4        m1034(.A(mai_mai_n1062_), .B(mai_mai_n1053_), .C(mai_mai_n1042_), .D(mai_mai_n1023_), .Y(mai06));
  NO2        m1035(.A(mai_mai_n349_), .B(mai_mai_n474_), .Y(mai_mai_n1064_));
  NA2        m1036(.A(mai_mai_n96_), .B(mai_mai_n1064_), .Y(mai_mai_n1065_));
  NO2        m1037(.A(mai_mai_n195_), .B(mai_mai_n86_), .Y(mai_mai_n1066_));
  NA2        m1038(.A(mai_mai_n1066_), .B(mai_mai_n329_), .Y(mai_mai_n1067_));
  NO3        m1039(.A(mai_mai_n509_), .B(mai_mai_n692_), .C(mai_mai_n510_), .Y(mai_mai_n1068_));
  OR2        m1040(.A(mai_mai_n1068_), .B(mai_mai_n760_), .Y(mai_mai_n1069_));
  NA3        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1067_), .C(mai_mai_n1065_), .Y(mai_mai_n1070_));
  NO3        m1042(.A(mai_mai_n1070_), .B(mai_mai_n1049_), .C(mai_mai_n224_), .Y(mai_mai_n1071_));
  INV        m1043(.A(mai_mai_n1054_), .Y(mai_mai_n1072_));
  NO2        m1044(.A(mai_mai_n1072_), .B(mai_mai_n295_), .Y(mai_mai_n1073_));
  NA2        m1045(.A(mai_mai_n83_), .B(mai_mai_n547_), .Y(mai_mai_n1074_));
  NO2        m1046(.A(mai_mai_n437_), .B(mai_mai_n148_), .Y(mai_mai_n1075_));
  NOi21      m1047(.An(mai_mai_n115_), .B(mai_mai_n43_), .Y(mai_mai_n1076_));
  NO2        m1048(.A(mai_mai_n515_), .B(mai_mai_n926_), .Y(mai_mai_n1077_));
  OAI210     m1049(.A0(mai_mai_n393_), .A1(mai_mai_n215_), .B0(mai_mai_n775_), .Y(mai_mai_n1078_));
  NO4        m1050(.A(mai_mai_n1078_), .B(mai_mai_n1077_), .C(mai_mai_n1076_), .D(mai_mai_n1075_), .Y(mai_mai_n1079_));
  NA2        m1051(.A(mai_mai_n1079_), .B(mai_mai_n1074_), .Y(mai_mai_n1080_));
  NO2        m1052(.A(mai_mai_n641_), .B(mai_mai_n315_), .Y(mai_mai_n1081_));
  NO3        m1053(.A(mai_mai_n578_), .B(mai_mai_n652_), .C(mai_mai_n540_), .Y(mai_mai_n1082_));
  NOi21      m1054(.An(mai_mai_n1081_), .B(mai_mai_n1082_), .Y(mai_mai_n1083_));
  NO3        m1055(.A(mai_mai_n1083_), .B(mai_mai_n1080_), .C(mai_mai_n1073_), .Y(mai_mai_n1084_));
  OAI220     m1056(.A0(mai_mai_n626_), .A1(mai_mai_n1238_), .B0(mai_mai_n195_), .B1(mai_mai_n524_), .Y(mai_mai_n1085_));
  OAI210     m1057(.A0(mai_mai_n242_), .A1(c), .B0(mai_mai_n546_), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n1085_), .Y(mai_mai_n1087_));
  OAI220     m1059(.A0(mai_mai_n598_), .A1(mai_mai_n215_), .B0(mai_mai_n433_), .B1(mai_mai_n437_), .Y(mai_mai_n1088_));
  NO2        m1060(.A(f), .B(j), .Y(mai_mai_n1089_));
  NOi21      m1061(.An(mai_mai_n1089_), .B(mai_mai_n572_), .Y(mai_mai_n1090_));
  NO2        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1088_), .Y(mai_mai_n1091_));
  NA4        m1063(.A(mai_mai_n680_), .B(mai_mai_n679_), .C(mai_mai_n374_), .D(mai_mai_n752_), .Y(mai_mai_n1092_));
  NAi31      m1064(.An(mai_mai_n641_), .B(mai_mai_n1092_), .C(mai_mai_n177_), .Y(mai_mai_n1093_));
  NA4        m1065(.A(mai_mai_n1093_), .B(mai_mai_n1091_), .C(mai_mai_n1087_), .D(mai_mai_n1004_), .Y(mai_mai_n1094_));
  NOi31      m1066(.An(mai_mai_n1068_), .B(mai_mai_n395_), .C(mai_mai_n337_), .Y(mai_mai_n1095_));
  OR3        m1067(.A(mai_mai_n1095_), .B(mai_mai_n671_), .C(mai_mai_n461_), .Y(mai_mai_n1096_));
  NO2        m1068(.A(mai_mai_n386_), .B(mai_mai_n320_), .Y(mai_mai_n1097_));
  NA2        m1069(.A(mai_mai_n1097_), .B(mai_mai_n1096_), .Y(mai_mai_n1098_));
  NA2        m1070(.A(mai_mai_n1081_), .B(mai_mai_n651_), .Y(mai_mai_n1099_));
  NO2        m1071(.A(mai_mai_n750_), .B(mai_mai_n407_), .Y(mai_mai_n1100_));
  NA2        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1099_), .Y(mai_mai_n1101_));
  NAi21      m1073(.An(j), .B(i), .Y(mai_mai_n1102_));
  NO3        m1074(.A(mai_mai_n1060_), .B(mai_mai_n1102_), .C(mai_mai_n380_), .Y(mai_mai_n1103_));
  NO4        m1075(.A(mai_mai_n1103_), .B(mai_mai_n1101_), .C(mai_mai_n1098_), .D(mai_mai_n1094_), .Y(mai_mai_n1104_));
  NA4        m1076(.A(mai_mai_n1104_), .B(mai_mai_n1084_), .C(mai_mai_n1071_), .D(mai_mai_n1062_), .Y(mai07));
  NOi21      m1077(.An(j), .B(k), .Y(mai_mai_n1106_));
  NA4        m1078(.A(mai_mai_n156_), .B(mai_mai_n91_), .C(mai_mai_n1106_), .D(f), .Y(mai_mai_n1107_));
  NAi21      m1079(.An(f), .B(c), .Y(mai_mai_n1108_));
  OR2        m1080(.A(e), .B(d), .Y(mai_mai_n1109_));
  OAI220     m1081(.A0(mai_mai_n1109_), .A1(mai_mai_n1108_), .B0(mai_mai_n532_), .B1(mai_mai_n283_), .Y(mai_mai_n1110_));
  NA3        m1082(.A(mai_mai_n1110_), .B(mai_mai_n1231_), .C(mai_mai_n156_), .Y(mai_mai_n1111_));
  NOi31      m1083(.An(n), .B(m), .C(b), .Y(mai_mai_n1112_));
  NO3        m1084(.A(mai_mai_n111_), .B(mai_mai_n387_), .C(h), .Y(mai_mai_n1113_));
  NA2        m1085(.A(mai_mai_n1111_), .B(mai_mai_n1107_), .Y(mai_mai_n1114_));
  NA2        m1086(.A(mai_mai_n72_), .B(mai_mai_n43_), .Y(mai_mai_n1115_));
  NO2        m1087(.A(mai_mai_n873_), .B(mai_mai_n380_), .Y(mai_mai_n1116_));
  NA3        m1088(.A(mai_mai_n1116_), .B(mai_mai_n1115_), .C(mai_mai_n184_), .Y(mai_mai_n1117_));
  NO2        m1089(.A(mai_mai_n883_), .B(mai_mai_n271_), .Y(mai_mai_n1118_));
  NA2        m1090(.A(mai_mai_n462_), .B(mai_mai_n68_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n1005_), .B(mai_mai_n256_), .Y(mai_mai_n1120_));
  NA3        m1092(.A(mai_mai_n1120_), .B(mai_mai_n1119_), .C(mai_mai_n1117_), .Y(mai_mai_n1121_));
  NO2        m1093(.A(mai_mai_n1121_), .B(mai_mai_n1114_), .Y(mai_mai_n1122_));
  NO3        m1094(.A(e), .B(d), .C(c), .Y(mai_mai_n1123_));
  NA2        m1095(.A(mai_mai_n1228_), .B(mai_mai_n1123_), .Y(mai_mai_n1124_));
  NO2        m1096(.A(mai_mai_n1124_), .B(mai_mai_n184_), .Y(mai_mai_n1125_));
  NA3        m1097(.A(mai_mai_n595_), .B(mai_mai_n1234_), .C(mai_mai_n95_), .Y(mai_mai_n1126_));
  NO2        m1098(.A(mai_mai_n1126_), .B(mai_mai_n43_), .Y(mai_mai_n1127_));
  NO2        m1099(.A(l), .B(k), .Y(mai_mai_n1128_));
  NOi41      m1100(.An(mai_mai_n467_), .B(mai_mai_n1128_), .C(mai_mai_n404_), .D(mai_mai_n380_), .Y(mai_mai_n1129_));
  NO3        m1101(.A(mai_mai_n1129_), .B(mai_mai_n1127_), .C(mai_mai_n1125_), .Y(mai_mai_n1130_));
  NO2        m1102(.A(mai_mai_n123_), .B(h), .Y(mai_mai_n1131_));
  NO2        m1103(.A(g), .B(c), .Y(mai_mai_n1132_));
  NA2        m1104(.A(mai_mai_n1132_), .B(mai_mai_n160_), .Y(mai_mai_n1133_));
  NO2        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1227_), .Y(mai_mai_n1134_));
  NA2        m1106(.A(mai_mai_n1134_), .B(mai_mai_n156_), .Y(mai_mai_n1135_));
  NO2        m1107(.A(mai_mai_n388_), .B(a), .Y(mai_mai_n1136_));
  NA3        m1108(.A(mai_mai_n1136_), .B(mai_mai_n1230_), .C(mai_mai_n96_), .Y(mai_mai_n1137_));
  NO2        m1109(.A(i), .B(h), .Y(mai_mai_n1138_));
  NO2        m1110(.A(mai_mai_n648_), .B(mai_mai_n161_), .Y(mai_mai_n1139_));
  NOi31      m1111(.An(m), .B(n), .C(b), .Y(mai_mai_n1140_));
  INV        m1112(.A(mai_mai_n1139_), .Y(mai_mai_n1141_));
  NA2        m1113(.A(mai_mai_n902_), .B(mai_mai_n397_), .Y(mai_mai_n1142_));
  NO4        m1114(.A(mai_mai_n1142_), .B(mai_mai_n879_), .C(mai_mai_n380_), .D(mai_mai_n43_), .Y(mai_mai_n1143_));
  NO3        m1115(.A(mai_mai_n39_), .B(i), .C(h), .Y(mai_mai_n1144_));
  INV        m1116(.A(mai_mai_n1143_), .Y(mai_mai_n1145_));
  AN4        m1117(.A(mai_mai_n1145_), .B(mai_mai_n1141_), .C(mai_mai_n1137_), .D(mai_mai_n1135_), .Y(mai_mai_n1146_));
  NA2        m1118(.A(mai_mai_n1112_), .B(mai_mai_n326_), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n161_), .B(b), .Y(mai_mai_n1148_));
  AOI220     m1120(.A0(mai_mai_n970_), .A1(mai_mai_n1148_), .B0(mai_mai_n909_), .B1(mai_mai_n1142_), .Y(mai_mai_n1149_));
  NO4        m1121(.A(mai_mai_n111_), .B(g), .C(f), .D(e), .Y(mai_mai_n1150_));
  OR2        m1122(.A(e), .B(a), .Y(mai_mai_n1151_));
  NA4        m1123(.A(mai_mai_n1149_), .B(mai_mai_n1146_), .C(mai_mai_n1130_), .D(mai_mai_n1122_), .Y(mai_mai_n1152_));
  NO2        m1124(.A(mai_mai_n334_), .B(j), .Y(mai_mai_n1153_));
  NA3        m1125(.A(mai_mai_n1144_), .B(mai_mai_n1109_), .C(mai_mai_n925_), .Y(mai_mai_n1154_));
  NAi31      m1126(.An(mai_mai_n1138_), .B(mai_mai_n891_), .C(mai_mai_n144_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n1155_), .B(mai_mai_n1154_), .Y(mai_mai_n1156_));
  NA3        m1128(.A(g), .B(mai_mai_n1153_), .C(mai_mai_n133_), .Y(mai_mai_n1157_));
  INV        m1129(.A(mai_mai_n1157_), .Y(mai_mai_n1158_));
  NO2        m1130(.A(mai_mai_n1158_), .B(mai_mai_n1156_), .Y(mai_mai_n1159_));
  OR2        m1131(.A(n), .B(i), .Y(mai_mai_n1160_));
  OAI210     m1132(.A0(mai_mai_n1160_), .A1(mai_mai_n890_), .B0(mai_mai_n46_), .Y(mai_mai_n1161_));
  AOI220     m1133(.A0(mai_mai_n1161_), .A1(mai_mai_n976_), .B0(mai_mai_n709_), .B1(mai_mai_n168_), .Y(mai_mai_n1162_));
  NO2        m1134(.A(mai_mai_n195_), .B(k), .Y(mai_mai_n1163_));
  NO3        m1135(.A(mai_mai_n912_), .B(mai_mai_n1109_), .C(mai_mai_n46_), .Y(mai_mai_n1164_));
  NOi21      m1136(.An(d), .B(f), .Y(mai_mai_n1165_));
  NO2        m1137(.A(mai_mai_n1109_), .B(f), .Y(mai_mai_n1166_));
  NA2        m1138(.A(mai_mai_n1162_), .B(mai_mai_n1159_), .Y(mai_mai_n1167_));
  OAI220     m1139(.A0(mai_mai_n397_), .A1(mai_mai_n266_), .B0(mai_mai_n110_), .B1(mai_mai_n51_), .Y(mai_mai_n1168_));
  NA2        m1140(.A(mai_mai_n1168_), .B(mai_mai_n1118_), .Y(mai_mai_n1169_));
  OAI210     m1141(.A0(mai_mai_n1150_), .A1(mai_mai_n1112_), .B0(mai_mai_n757_), .Y(mai_mai_n1170_));
  NO2        m1142(.A(c), .B(mai_mai_n111_), .Y(mai_mai_n1171_));
  NA2        m1143(.A(mai_mai_n1171_), .B(mai_mai_n528_), .Y(mai_mai_n1172_));
  NA3        m1144(.A(mai_mai_n1172_), .B(mai_mai_n1170_), .C(mai_mai_n1169_), .Y(mai_mai_n1173_));
  NA2        m1145(.A(mai_mai_n1132_), .B(mai_mai_n1165_), .Y(mai_mai_n1174_));
  NO2        m1146(.A(mai_mai_n1174_), .B(m), .Y(mai_mai_n1175_));
  OAI220     m1147(.A0(mai_mai_n126_), .A1(mai_mai_n157_), .B0(mai_mai_n387_), .B1(g), .Y(mai_mai_n1176_));
  OAI210     m1148(.A0(mai_mai_n1176_), .A1(mai_mai_n93_), .B0(mai_mai_n1140_), .Y(mai_mai_n1177_));
  INV        m1149(.A(mai_mai_n1177_), .Y(mai_mai_n1178_));
  NO3        m1150(.A(mai_mai_n1178_), .B(mai_mai_n1175_), .C(mai_mai_n1173_), .Y(mai_mai_n1179_));
  NO2        m1151(.A(mai_mai_n1108_), .B(e), .Y(mai_mai_n1180_));
  INV        m1152(.A(mai_mai_n1180_), .Y(mai_mai_n1181_));
  OAI210     m1153(.A0(mai_mai_n1166_), .A1(mai_mai_n933_), .B0(mai_mai_n536_), .Y(mai_mai_n1182_));
  OR3        m1154(.A(mai_mai_n1163_), .B(mai_mai_n1005_), .C(mai_mai_n111_), .Y(mai_mai_n1183_));
  OAI220     m1155(.A0(mai_mai_n1183_), .A1(mai_mai_n1181_), .B0(mai_mai_n1182_), .B1(mai_mai_n382_), .Y(mai_mai_n1184_));
  INV        m1156(.A(mai_mai_n1184_), .Y(mai_mai_n1185_));
  NA2        m1157(.A(mai_mai_n1180_), .B(mai_mai_n156_), .Y(mai_mai_n1186_));
  AOI220     m1158(.A0(mai_mai_n1186_), .A1(mai_mai_n892_), .B0(mai_mai_n454_), .B1(mai_mai_n315_), .Y(mai_mai_n1187_));
  NO2        m1159(.A(mai_mai_n1151_), .B(f), .Y(mai_mai_n1188_));
  NA2        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1115_), .Y(mai_mai_n1189_));
  OAI220     m1161(.A0(mai_mai_n1189_), .A1(mai_mai_n46_), .B0(mai_mai_n1229_), .B1(mai_mai_n151_), .Y(mai_mai_n1190_));
  NA4        m1162(.A(mai_mai_n910_), .B(mai_mai_n907_), .C(mai_mai_n191_), .D(mai_mai_n59_), .Y(mai_mai_n1191_));
  NA2        m1163(.A(mai_mai_n1113_), .B(mai_mai_n158_), .Y(mai_mai_n1192_));
  NO2        m1164(.A(mai_mai_n46_), .B(l), .Y(mai_mai_n1193_));
  OAI210     m1165(.A0(mai_mai_n1151_), .A1(mai_mai_n743_), .B0(mai_mai_n409_), .Y(mai_mai_n1194_));
  OAI210     m1166(.A0(mai_mai_n1194_), .A1(mai_mai_n913_), .B0(mai_mai_n1193_), .Y(mai_mai_n1195_));
  NO2        m1167(.A(mai_mai_n220_), .B(g), .Y(mai_mai_n1196_));
  NO2        m1168(.A(m), .B(i), .Y(mai_mai_n1197_));
  BUFFER     m1169(.A(mai_mai_n1197_), .Y(mai_mai_n1198_));
  AOI220     m1170(.A0(mai_mai_n1198_), .A1(mai_mai_n1131_), .B0(mai_mai_n891_), .B1(mai_mai_n1196_), .Y(mai_mai_n1199_));
  NA4        m1171(.A(mai_mai_n1199_), .B(mai_mai_n1195_), .C(mai_mai_n1192_), .D(mai_mai_n1191_), .Y(mai_mai_n1200_));
  NO4        m1172(.A(mai_mai_n1200_), .B(mai_mai_n1190_), .C(mai_mai_n1164_), .D(mai_mai_n1187_), .Y(mai_mai_n1201_));
  NA3        m1173(.A(mai_mai_n1201_), .B(mai_mai_n1185_), .C(mai_mai_n1179_), .Y(mai_mai_n1202_));
  NA3        m1174(.A(mai_mai_n813_), .B(mai_mai_n117_), .C(mai_mai_n44_), .Y(mai_mai_n1203_));
  AOI210     m1175(.A0(mai_mai_n124_), .A1(c), .B0(mai_mai_n1203_), .Y(mai_mai_n1204_));
  AO210      m1176(.A0(mai_mai_n112_), .A1(l), .B0(mai_mai_n1147_), .Y(mai_mai_n1205_));
  INV        m1177(.A(mai_mai_n1205_), .Y(mai_mai_n1206_));
  NO2        m1178(.A(mai_mai_n1206_), .B(mai_mai_n1204_), .Y(mai_mai_n1207_));
  NO4        m1179(.A(mai_mai_n195_), .B(mai_mai_n159_), .C(mai_mai_n225_), .D(k), .Y(mai_mai_n1208_));
  NOi21      m1180(.An(mai_mai_n1113_), .B(e), .Y(mai_mai_n1209_));
  NO2        m1181(.A(mai_mai_n1209_), .B(mai_mai_n1208_), .Y(mai_mai_n1210_));
  AN2        m1182(.A(mai_mai_n910_), .B(mai_mai_n898_), .Y(mai_mai_n1211_));
  AOI220     m1183(.A0(mai_mai_n1197_), .A1(mai_mai_n545_), .B0(mai_mai_n1231_), .B1(mai_mai_n134_), .Y(mai_mai_n1212_));
  NOi21      m1184(.An(mai_mai_n30_), .B(mai_mai_n1212_), .Y(mai_mai_n1213_));
  AOI210     m1185(.A0(mai_mai_n1211_), .A1(mai_mai_n970_), .B0(mai_mai_n1213_), .Y(mai_mai_n1214_));
  NA3        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1210_), .C(mai_mai_n1207_), .Y(mai_mai_n1215_));
  OR4        m1187(.A(mai_mai_n1215_), .B(mai_mai_n1202_), .C(mai_mai_n1167_), .D(mai_mai_n1152_), .Y(mai04));
  NA2        m1188(.A(mai_mai_n1166_), .B(mai_mai_n709_), .Y(mai_mai_n1217_));
  NO2        m1189(.A(mai_mai_n1217_), .B(j), .Y(mai_mai_n1218_));
  OR3        m1190(.A(mai_mai_n1218_), .B(mai_mai_n1150_), .C(mai_mai_n882_), .Y(mai_mai_n1219_));
  NO2        m1191(.A(mai_mai_n1115_), .B(mai_mai_n75_), .Y(mai_mai_n1220_));
  AOI210     m1192(.A0(mai_mai_n1220_), .A1(mai_mai_n876_), .B0(mai_mai_n986_), .Y(mai_mai_n1221_));
  NA2        m1193(.A(mai_mai_n1221_), .B(mai_mai_n1009_), .Y(mai_mai_n1222_));
  NO4        m1194(.A(mai_mai_n1222_), .B(mai_mai_n1219_), .C(mai_mai_n889_), .D(mai_mai_n872_), .Y(mai_mai_n1223_));
  NA4        m1195(.A(mai_mai_n1223_), .B(mai_mai_n935_), .C(mai_mai_n923_), .D(mai_mai_n916_), .Y(mai05));
  INV        m1196(.A(l), .Y(mai_mai_n1227_));
  INV        m1197(.A(m), .Y(mai_mai_n1228_));
  INV        m1198(.A(mai_mai_n88_), .Y(mai_mai_n1229_));
  INV        m1199(.A(i), .Y(mai_mai_n1230_));
  INV        m1200(.A(j), .Y(mai_mai_n1231_));
  INV        m1201(.A(c), .Y(mai_mai_n1232_));
  INV        m1202(.A(mai_mai_n399_), .Y(mai_mai_n1233_));
  INV        m1203(.A(m), .Y(mai_mai_n1234_));
  INV        m1204(.A(mai_mai_n96_), .Y(mai_mai_n1235_));
  INV        m1205(.A(mai_mai_n358_), .Y(mai_mai_n1236_));
  INV        m1206(.A(mai_mai_n472_), .Y(mai_mai_n1237_));
  INV        m1207(.A(h), .Y(mai_mai_n1238_));
  INV        m1208(.A(n), .Y(mai_mai_n1239_));
  INV        m1209(.A(k), .Y(mai_mai_n1240_));
  INV        m1210(.A(f), .Y(mai_mai_n1241_));
  INV        m1211(.A(m), .Y(mai_mai_n1242_));
  INV        m1212(.A(n), .Y(mai_mai_n1243_));
  INV        m1213(.A(m), .Y(mai_mai_n1244_));
  INV        m1214(.A(f), .Y(mai_mai_n1245_));
  INV        m1215(.A(g), .Y(mai_mai_n1246_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA2        u0003(.A(men_men_n31_), .B(men_men_n30_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO2        u0025(.A(men_men_n53_), .B(men_men_n48_), .Y(men_men_n54_));
  NO2        u0026(.A(men_men_n54_), .B(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  INV        u0028(.A(d), .Y(men_men_n57_));
  NA2        u0029(.A(g), .B(a), .Y(men_men_n58_));
  NAi21      u0030(.An(i), .B(h), .Y(men_men_n59_));
  NAi31      u0031(.An(i), .B(l), .C(j), .Y(men_men_n60_));
  NAi41      u0032(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n61_));
  NA2        u0033(.A(g), .B(f), .Y(men_men_n62_));
  NO2        u0034(.A(men_men_n62_), .B(men_men_n61_), .Y(men_men_n63_));
  NAi21      u0035(.An(i), .B(j), .Y(men_men_n64_));
  NAi32      u0036(.An(n), .Bn(k), .C(m), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi31      u0038(.An(l), .B(m), .C(k), .Y(men_men_n67_));
  NAi21      u0039(.An(e), .B(h), .Y(men_men_n68_));
  NAi41      u0040(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n69_));
  NA2        u0041(.A(men_men_n66_), .B(men_men_n63_), .Y(men_men_n70_));
  INV        u0042(.A(m), .Y(men_men_n71_));
  NOi21      u0043(.An(k), .B(l), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n73_));
  AN4        u0045(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n74_));
  NOi31      u0046(.An(h), .B(g), .C(f), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  NAi32      u0048(.An(m), .Bn(k), .C(j), .Y(men_men_n77_));
  NOi32      u0049(.An(h), .Bn(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n78_), .B(men_men_n74_), .Y(men_men_n79_));
  OA220      u0051(.A0(men_men_n79_), .A1(men_men_n77_), .B0(men_men_n76_), .B1(men_men_n73_), .Y(men_men_n80_));
  NA2        u0052(.A(men_men_n80_), .B(men_men_n70_), .Y(men_men_n81_));
  INV        u0053(.A(n), .Y(men_men_n82_));
  NOi32      u0054(.An(e), .Bn(b), .C(d), .Y(men_men_n83_));
  NA2        u0055(.A(men_men_n83_), .B(men_men_n82_), .Y(men_men_n84_));
  INV        u0056(.A(j), .Y(men_men_n85_));
  AN3        u0057(.A(m), .B(k), .C(i), .Y(men_men_n86_));
  NA3        u0058(.A(men_men_n86_), .B(men_men_n85_), .C(g), .Y(men_men_n87_));
  NO2        u0059(.A(men_men_n87_), .B(f), .Y(men_men_n88_));
  NAi32      u0060(.An(g), .Bn(f), .C(h), .Y(men_men_n89_));
  NAi31      u0061(.An(j), .B(m), .C(l), .Y(men_men_n90_));
  NO2        u0062(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n91_));
  NA2        u0063(.A(m), .B(l), .Y(men_men_n92_));
  NAi31      u0064(.An(k), .B(j), .C(g), .Y(men_men_n93_));
  NO3        u0065(.A(men_men_n93_), .B(men_men_n92_), .C(f), .Y(men_men_n94_));
  AN2        u0066(.A(j), .B(g), .Y(men_men_n95_));
  NOi32      u0067(.An(m), .Bn(l), .C(i), .Y(men_men_n96_));
  NOi21      u0068(.An(g), .B(i), .Y(men_men_n97_));
  NOi32      u0069(.An(m), .Bn(j), .C(k), .Y(men_men_n98_));
  AOI220     u0070(.A0(men_men_n98_), .A1(men_men_n97_), .B0(men_men_n96_), .B1(men_men_n95_), .Y(men_men_n99_));
  NO2        u0071(.A(men_men_n99_), .B(f), .Y(men_men_n100_));
  NAi41      u0072(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n101_));
  AN2        u0073(.A(e), .B(b), .Y(men_men_n102_));
  NOi31      u0074(.An(c), .B(h), .C(f), .Y(men_men_n103_));
  NA2        u0075(.A(men_men_n103_), .B(men_men_n102_), .Y(men_men_n104_));
  NOi21      u0076(.An(i), .B(h), .Y(men_men_n105_));
  NA3        u0077(.A(men_men_n105_), .B(g), .C(men_men_n36_), .Y(men_men_n106_));
  INV        u0078(.A(a), .Y(men_men_n107_));
  INV        u0079(.A(men_men_n102_), .Y(men_men_n108_));
  INV        u0080(.A(l), .Y(men_men_n109_));
  NOi21      u0081(.An(m), .B(n), .Y(men_men_n110_));
  NO2        u0082(.A(men_men_n106_), .B(men_men_n84_), .Y(men_men_n111_));
  INV        u0083(.A(b), .Y(men_men_n112_));
  NA2        u0084(.A(l), .B(j), .Y(men_men_n113_));
  AN2        u0085(.A(k), .B(i), .Y(men_men_n114_));
  NA2        u0086(.A(men_men_n114_), .B(men_men_n113_), .Y(men_men_n115_));
  NA2        u0087(.A(g), .B(e), .Y(men_men_n116_));
  NOi32      u0088(.An(c), .Bn(a), .C(d), .Y(men_men_n117_));
  NA2        u0089(.A(men_men_n117_), .B(men_men_n110_), .Y(men_men_n118_));
  INV        u0090(.A(men_men_n111_), .Y(men_men_n119_));
  OAI210     u0091(.A0(men_men_n87_), .A1(men_men_n84_), .B0(men_men_n119_), .Y(men_men_n120_));
  NOi31      u0092(.An(k), .B(m), .C(j), .Y(men_men_n121_));
  NA3        u0093(.A(men_men_n121_), .B(men_men_n75_), .C(men_men_n74_), .Y(men_men_n122_));
  NOi31      u0094(.An(k), .B(m), .C(i), .Y(men_men_n123_));
  NA3        u0095(.A(men_men_n123_), .B(men_men_n78_), .C(men_men_n74_), .Y(men_men_n124_));
  NA2        u0096(.A(men_men_n124_), .B(men_men_n122_), .Y(men_men_n125_));
  NAi21      u0097(.An(g), .B(h), .Y(men_men_n126_));
  NAi21      u0098(.An(m), .B(n), .Y(men_men_n127_));
  NAi21      u0099(.An(j), .B(k), .Y(men_men_n128_));
  NAi41      u0100(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n129_));
  NAi31      u0101(.An(j), .B(k), .C(h), .Y(men_men_n130_));
  NO2        u0102(.A(k), .B(j), .Y(men_men_n131_));
  NO2        u0103(.A(men_men_n131_), .B(men_men_n127_), .Y(men_men_n132_));
  AN2        u0104(.A(k), .B(j), .Y(men_men_n133_));
  NAi21      u0105(.An(c), .B(b), .Y(men_men_n134_));
  NA2        u0106(.A(f), .B(d), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n126_), .Y(men_men_n136_));
  NA2        u0108(.A(h), .B(c), .Y(men_men_n137_));
  NAi31      u0109(.An(f), .B(e), .C(b), .Y(men_men_n138_));
  NA2        u0110(.A(men_men_n136_), .B(men_men_n132_), .Y(men_men_n139_));
  NA2        u0111(.A(d), .B(b), .Y(men_men_n140_));
  NAi21      u0112(.An(e), .B(f), .Y(men_men_n141_));
  NO2        u0113(.A(men_men_n141_), .B(men_men_n140_), .Y(men_men_n142_));
  NA2        u0114(.A(b), .B(a), .Y(men_men_n143_));
  NAi21      u0115(.An(e), .B(g), .Y(men_men_n144_));
  NAi21      u0116(.An(c), .B(d), .Y(men_men_n145_));
  NAi31      u0117(.An(l), .B(k), .C(h), .Y(men_men_n146_));
  NO2        u0118(.A(men_men_n127_), .B(men_men_n146_), .Y(men_men_n147_));
  NA2        u0119(.A(men_men_n147_), .B(men_men_n142_), .Y(men_men_n148_));
  NAi31      u0120(.An(men_men_n125_), .B(men_men_n148_), .C(men_men_n139_), .Y(men_men_n149_));
  NAi31      u0121(.An(e), .B(f), .C(b), .Y(men_men_n150_));
  NOi21      u0122(.An(g), .B(d), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n151_), .B(men_men_n150_), .Y(men_men_n152_));
  NOi21      u0124(.An(k), .B(m), .Y(men_men_n153_));
  NA3        u0125(.A(men_men_n153_), .B(h), .C(n), .Y(men_men_n154_));
  NOi21      u0126(.An(men_men_n152_), .B(men_men_n154_), .Y(men_men_n155_));
  NOi21      u0127(.An(h), .B(g), .Y(men_men_n156_));
  NO2        u0128(.A(men_men_n135_), .B(men_men_n134_), .Y(men_men_n157_));
  NAi31      u0129(.An(l), .B(j), .C(h), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n158_), .B(men_men_n49_), .Y(men_men_n159_));
  NA2        u0131(.A(men_men_n159_), .B(men_men_n63_), .Y(men_men_n160_));
  INV        u0132(.A(men_men_n160_), .Y(men_men_n161_));
  NAi31      u0133(.An(e), .B(f), .C(c), .Y(men_men_n162_));
  NA2        u0134(.A(j), .B(h), .Y(men_men_n163_));
  OR3        u0135(.A(n), .B(m), .C(k), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  NAi32      u0137(.An(m), .Bn(k), .C(n), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n166_), .B(men_men_n163_), .Y(men_men_n167_));
  NA2        u0139(.A(men_men_n167_), .B(men_men_n152_), .Y(men_men_n168_));
  NO2        u0140(.A(n), .B(m), .Y(men_men_n169_));
  NA2        u0141(.A(men_men_n169_), .B(men_men_n50_), .Y(men_men_n170_));
  NAi21      u0142(.An(f), .B(e), .Y(men_men_n171_));
  NA2        u0143(.A(d), .B(c), .Y(men_men_n172_));
  NO2        u0144(.A(men_men_n172_), .B(men_men_n171_), .Y(men_men_n173_));
  NOi21      u0145(.An(men_men_n173_), .B(men_men_n170_), .Y(men_men_n174_));
  NAi21      u0146(.An(d), .B(c), .Y(men_men_n175_));
  NAi31      u0147(.An(m), .B(n), .C(b), .Y(men_men_n176_));
  NAi21      u0148(.An(h), .B(f), .Y(men_men_n177_));
  NO2        u0149(.A(men_men_n176_), .B(men_men_n145_), .Y(men_men_n178_));
  NOi32      u0150(.An(f), .Bn(c), .C(d), .Y(men_men_n179_));
  NOi32      u0151(.An(f), .Bn(c), .C(e), .Y(men_men_n180_));
  NO2        u0152(.A(men_men_n180_), .B(men_men_n179_), .Y(men_men_n181_));
  NO3        u0153(.A(n), .B(m), .C(j), .Y(men_men_n182_));
  NA2        u0154(.A(men_men_n182_), .B(h), .Y(men_men_n183_));
  AO210      u0155(.A0(men_men_n183_), .A1(men_men_n170_), .B0(men_men_n181_), .Y(men_men_n184_));
  NAi31      u0156(.An(men_men_n174_), .B(men_men_n184_), .C(men_men_n168_), .Y(men_men_n185_));
  OR4        u0157(.A(men_men_n185_), .B(men_men_n161_), .C(men_men_n155_), .D(men_men_n149_), .Y(men_men_n186_));
  NO4        u0158(.A(men_men_n186_), .B(men_men_n120_), .C(men_men_n81_), .D(men_men_n55_), .Y(men_men_n187_));
  NA3        u0159(.A(m), .B(men_men_n109_), .C(j), .Y(men_men_n188_));
  NAi31      u0160(.An(n), .B(h), .C(g), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NOi32      u0162(.An(m), .Bn(k), .C(l), .Y(men_men_n191_));
  NA3        u0163(.A(men_men_n191_), .B(men_men_n85_), .C(g), .Y(men_men_n192_));
  NO2        u0164(.A(men_men_n192_), .B(n), .Y(men_men_n193_));
  NOi21      u0165(.An(k), .B(j), .Y(men_men_n194_));
  NA4        u0166(.A(men_men_n194_), .B(men_men_n110_), .C(i), .D(g), .Y(men_men_n195_));
  AN2        u0167(.A(i), .B(g), .Y(men_men_n196_));
  NA3        u0168(.A(men_men_n72_), .B(men_men_n196_), .C(men_men_n110_), .Y(men_men_n197_));
  NA2        u0169(.A(men_men_n197_), .B(men_men_n195_), .Y(men_men_n198_));
  NO2        u0170(.A(men_men_n198_), .B(men_men_n193_), .Y(men_men_n199_));
  NAi41      u0171(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n200_));
  INV        u0172(.A(men_men_n200_), .Y(men_men_n201_));
  INV        u0173(.A(f), .Y(men_men_n202_));
  INV        u0174(.A(g), .Y(men_men_n203_));
  NOi31      u0175(.An(i), .B(j), .C(h), .Y(men_men_n204_));
  NOi21      u0176(.An(l), .B(m), .Y(men_men_n205_));
  NA2        u0177(.A(men_men_n205_), .B(men_men_n204_), .Y(men_men_n206_));
  NO3        u0178(.A(men_men_n206_), .B(men_men_n203_), .C(men_men_n202_), .Y(men_men_n207_));
  NA2        u0179(.A(men_men_n207_), .B(men_men_n201_), .Y(men_men_n208_));
  OAI210     u0180(.A0(men_men_n199_), .A1(men_men_n32_), .B0(men_men_n208_), .Y(men_men_n209_));
  NOi21      u0181(.An(n), .B(m), .Y(men_men_n210_));
  NA2        u0182(.A(i), .B(men_men_n210_), .Y(men_men_n211_));
  OR2        u0183(.A(men_men_n211_), .B(men_men_n104_), .Y(men_men_n212_));
  NAi21      u0184(.An(j), .B(h), .Y(men_men_n213_));
  XN2        u0185(.A(i), .B(h), .Y(men_men_n214_));
  NOi31      u0186(.An(k), .B(n), .C(m), .Y(men_men_n215_));
  NAi31      u0187(.An(f), .B(e), .C(c), .Y(men_men_n216_));
  NO3        u0188(.A(men_men_n216_), .B(men_men_n164_), .C(men_men_n163_), .Y(men_men_n217_));
  NA4        u0189(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n218_));
  NAi32      u0190(.An(m), .Bn(i), .C(k), .Y(men_men_n219_));
  NO3        u0191(.A(men_men_n219_), .B(men_men_n89_), .C(men_men_n218_), .Y(men_men_n220_));
  NO2        u0192(.A(men_men_n220_), .B(men_men_n217_), .Y(men_men_n221_));
  NAi21      u0193(.An(n), .B(a), .Y(men_men_n222_));
  NO2        u0194(.A(men_men_n222_), .B(men_men_n140_), .Y(men_men_n223_));
  NAi41      u0195(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n224_));
  NO2        u0196(.A(men_men_n224_), .B(e), .Y(men_men_n225_));
  NO3        u0197(.A(men_men_n141_), .B(men_men_n93_), .C(men_men_n92_), .Y(men_men_n226_));
  OAI210     u0198(.A0(men_men_n226_), .A1(men_men_n225_), .B0(men_men_n223_), .Y(men_men_n227_));
  AN3        u0199(.A(men_men_n227_), .B(men_men_n221_), .C(men_men_n212_), .Y(men_men_n228_));
  NAi41      u0200(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n229_));
  NO2        u0201(.A(men_men_n229_), .B(men_men_n202_), .Y(men_men_n230_));
  NA2        u0202(.A(men_men_n153_), .B(men_men_n105_), .Y(men_men_n231_));
  NAi21      u0203(.An(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  NO2        u0204(.A(n), .B(a), .Y(men_men_n233_));
  NAi31      u0205(.An(men_men_n224_), .B(men_men_n233_), .C(men_men_n102_), .Y(men_men_n234_));
  AN2        u0206(.A(men_men_n234_), .B(men_men_n232_), .Y(men_men_n235_));
  NAi21      u0207(.An(h), .B(i), .Y(men_men_n236_));
  NA2        u0208(.A(men_men_n169_), .B(k), .Y(men_men_n237_));
  NO2        u0209(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  INV        u0210(.A(men_men_n235_), .Y(men_men_n239_));
  NOi21      u0211(.An(g), .B(e), .Y(men_men_n240_));
  NO2        u0212(.A(men_men_n69_), .B(men_men_n71_), .Y(men_men_n241_));
  NA2        u0213(.A(men_men_n241_), .B(men_men_n240_), .Y(men_men_n242_));
  NOi32      u0214(.An(l), .Bn(j), .C(i), .Y(men_men_n243_));
  AOI210     u0215(.A0(men_men_n72_), .A1(men_men_n85_), .B0(men_men_n243_), .Y(men_men_n244_));
  NO2        u0216(.A(men_men_n236_), .B(men_men_n44_), .Y(men_men_n245_));
  NAi21      u0217(.An(f), .B(g), .Y(men_men_n246_));
  NO2        u0218(.A(men_men_n246_), .B(men_men_n61_), .Y(men_men_n247_));
  NO2        u0219(.A(men_men_n65_), .B(men_men_n113_), .Y(men_men_n248_));
  AOI220     u0220(.A0(men_men_n248_), .A1(men_men_n247_), .B0(men_men_n245_), .B1(men_men_n63_), .Y(men_men_n249_));
  OAI210     u0221(.A0(men_men_n244_), .A1(men_men_n242_), .B0(men_men_n249_), .Y(men_men_n250_));
  NO3        u0222(.A(men_men_n128_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n251_));
  NOi41      u0223(.An(men_men_n228_), .B(men_men_n250_), .C(men_men_n239_), .D(men_men_n209_), .Y(men_men_n252_));
  NO4        u0224(.A(men_men_n190_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n253_));
  NO2        u0225(.A(men_men_n253_), .B(men_men_n108_), .Y(men_men_n254_));
  NA3        u0226(.A(men_men_n57_), .B(c), .C(b), .Y(men_men_n255_));
  NAi21      u0227(.An(h), .B(g), .Y(men_men_n256_));
  OR4        u0228(.A(men_men_n256_), .B(men_men_n255_), .C(men_men_n211_), .D(e), .Y(men_men_n257_));
  NAi31      u0229(.An(g), .B(k), .C(h), .Y(men_men_n258_));
  NO3        u0230(.A(men_men_n127_), .B(men_men_n258_), .C(l), .Y(men_men_n259_));
  NAi31      u0231(.An(e), .B(d), .C(a), .Y(men_men_n260_));
  INV        u0232(.A(men_men_n257_), .Y(men_men_n261_));
  NA4        u0233(.A(men_men_n153_), .B(men_men_n78_), .C(men_men_n74_), .D(men_men_n113_), .Y(men_men_n262_));
  NA3        u0234(.A(men_men_n153_), .B(h), .C(men_men_n82_), .Y(men_men_n263_));
  NA3        u0235(.A(e), .B(c), .C(b), .Y(men_men_n264_));
  NO2        u0236(.A(men_men_n58_), .B(men_men_n264_), .Y(men_men_n265_));
  NAi32      u0237(.An(k), .Bn(i), .C(j), .Y(men_men_n266_));
  INV        u0238(.A(men_men_n49_), .Y(men_men_n267_));
  OAI210     u0239(.A0(men_men_n247_), .A1(men_men_n265_), .B0(men_men_n267_), .Y(men_men_n268_));
  NAi21      u0240(.An(l), .B(k), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n269_), .B(men_men_n49_), .Y(men_men_n270_));
  NOi21      u0242(.An(l), .B(j), .Y(men_men_n271_));
  NA2        u0243(.A(men_men_n156_), .B(men_men_n271_), .Y(men_men_n272_));
  NA3        u0244(.A(men_men_n114_), .B(men_men_n113_), .C(g), .Y(men_men_n273_));
  OR3        u0245(.A(men_men_n69_), .B(men_men_n71_), .C(e), .Y(men_men_n274_));
  AOI210     u0246(.A0(men_men_n273_), .A1(men_men_n272_), .B0(men_men_n274_), .Y(men_men_n275_));
  INV        u0247(.A(men_men_n275_), .Y(men_men_n276_));
  NAi32      u0248(.An(j), .Bn(h), .C(i), .Y(men_men_n277_));
  NAi21      u0249(.An(m), .B(l), .Y(men_men_n278_));
  NO3        u0250(.A(men_men_n278_), .B(men_men_n277_), .C(men_men_n82_), .Y(men_men_n279_));
  NA2        u0251(.A(h), .B(g), .Y(men_men_n280_));
  NA2        u0252(.A(men_men_n279_), .B(men_men_n157_), .Y(men_men_n281_));
  NA4        u0253(.A(men_men_n281_), .B(men_men_n276_), .C(men_men_n268_), .D(men_men_n262_), .Y(men_men_n282_));
  NO2        u0254(.A(men_men_n138_), .B(d), .Y(men_men_n283_));
  NA2        u0255(.A(men_men_n283_), .B(men_men_n53_), .Y(men_men_n284_));
  NAi32      u0256(.An(n), .Bn(m), .C(l), .Y(men_men_n285_));
  NO2        u0257(.A(men_men_n285_), .B(men_men_n277_), .Y(men_men_n286_));
  NA2        u0258(.A(men_men_n286_), .B(men_men_n173_), .Y(men_men_n287_));
  NAi31      u0259(.An(k), .B(l), .C(j), .Y(men_men_n288_));
  OAI210     u0260(.A0(men_men_n269_), .A1(j), .B0(men_men_n288_), .Y(men_men_n289_));
  NOi21      u0261(.An(men_men_n289_), .B(men_men_n116_), .Y(men_men_n290_));
  NA2        u0262(.A(men_men_n287_), .B(men_men_n284_), .Y(men_men_n291_));
  NO4        u0263(.A(men_men_n291_), .B(men_men_n282_), .C(men_men_n261_), .D(men_men_n254_), .Y(men_men_n292_));
  NA2        u0264(.A(men_men_n238_), .B(men_men_n180_), .Y(men_men_n293_));
  NAi21      u0265(.An(m), .B(k), .Y(men_men_n294_));
  NO2        u0266(.A(men_men_n214_), .B(men_men_n294_), .Y(men_men_n295_));
  NAi41      u0267(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n296_));
  NO2        u0268(.A(men_men_n296_), .B(men_men_n144_), .Y(men_men_n297_));
  NA2        u0269(.A(men_men_n297_), .B(men_men_n295_), .Y(men_men_n298_));
  NAi31      u0270(.An(i), .B(l), .C(h), .Y(men_men_n299_));
  NO4        u0271(.A(men_men_n299_), .B(men_men_n144_), .C(men_men_n69_), .D(men_men_n71_), .Y(men_men_n300_));
  NA2        u0272(.A(e), .B(c), .Y(men_men_n301_));
  NO3        u0273(.A(men_men_n301_), .B(n), .C(d), .Y(men_men_n302_));
  NOi21      u0274(.An(f), .B(h), .Y(men_men_n303_));
  NA2        u0275(.A(men_men_n303_), .B(men_men_n114_), .Y(men_men_n304_));
  NO2        u0276(.A(men_men_n304_), .B(men_men_n203_), .Y(men_men_n305_));
  NAi31      u0277(.An(d), .B(e), .C(b), .Y(men_men_n306_));
  NO2        u0278(.A(men_men_n127_), .B(men_men_n306_), .Y(men_men_n307_));
  NAi31      u0279(.An(men_men_n300_), .B(men_men_n298_), .C(men_men_n293_), .Y(men_men_n308_));
  NO4        u0280(.A(men_men_n296_), .B(men_men_n77_), .C(men_men_n68_), .D(men_men_n203_), .Y(men_men_n309_));
  NA2        u0281(.A(men_men_n233_), .B(men_men_n102_), .Y(men_men_n310_));
  NOi31      u0282(.An(l), .B(n), .C(m), .Y(men_men_n311_));
  NA2        u0283(.A(men_men_n311_), .B(men_men_n204_), .Y(men_men_n312_));
  NO2        u0284(.A(men_men_n312_), .B(men_men_n181_), .Y(men_men_n313_));
  OR2        u0285(.A(men_men_n313_), .B(men_men_n309_), .Y(men_men_n314_));
  NAi32      u0286(.An(m), .Bn(j), .C(k), .Y(men_men_n315_));
  NAi41      u0287(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n316_));
  INV        u0288(.A(men_men_n316_), .Y(men_men_n317_));
  NOi31      u0289(.An(j), .B(m), .C(k), .Y(men_men_n318_));
  NO2        u0290(.A(men_men_n121_), .B(men_men_n318_), .Y(men_men_n319_));
  AN3        u0291(.A(h), .B(g), .C(f), .Y(men_men_n320_));
  NA2        u0292(.A(men_men_n320_), .B(men_men_n317_), .Y(men_men_n321_));
  NOi32      u0293(.An(m), .Bn(j), .C(l), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n278_), .B(men_men_n277_), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n206_), .B(g), .Y(men_men_n324_));
  NO2        u0296(.A(men_men_n150_), .B(men_men_n82_), .Y(men_men_n325_));
  AOI220     u0297(.A0(men_men_n325_), .A1(men_men_n324_), .B0(men_men_n230_), .B1(men_men_n323_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n219_), .B(men_men_n77_), .Y(men_men_n327_));
  NA3        u0299(.A(men_men_n327_), .B(men_men_n320_), .C(men_men_n201_), .Y(men_men_n328_));
  NA3        u0300(.A(men_men_n328_), .B(men_men_n326_), .C(men_men_n321_), .Y(men_men_n329_));
  NA3        u0301(.A(h), .B(g), .C(f), .Y(men_men_n330_));
  NA2        u0302(.A(men_men_n156_), .B(e), .Y(men_men_n331_));
  NO2        u0303(.A(men_men_n331_), .B(men_men_n41_), .Y(men_men_n332_));
  NOi32      u0304(.An(j), .Bn(g), .C(i), .Y(men_men_n333_));
  NA3        u0305(.A(men_men_n333_), .B(men_men_n269_), .C(men_men_n110_), .Y(men_men_n334_));
  AO210      u0306(.A0(men_men_n108_), .A1(men_men_n32_), .B0(men_men_n334_), .Y(men_men_n335_));
  NOi32      u0307(.An(e), .Bn(b), .C(a), .Y(men_men_n336_));
  AN2        u0308(.A(l), .B(j), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n294_), .B(men_men_n337_), .Y(men_men_n338_));
  NO3        u0310(.A(men_men_n296_), .B(men_men_n68_), .C(men_men_n203_), .Y(men_men_n339_));
  NA3        u0311(.A(men_men_n197_), .B(men_men_n195_), .C(men_men_n35_), .Y(men_men_n340_));
  AOI220     u0312(.A0(men_men_n340_), .A1(men_men_n336_), .B0(men_men_n339_), .B1(men_men_n338_), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n306_), .B(n), .Y(men_men_n342_));
  NA2        u0314(.A(men_men_n196_), .B(k), .Y(men_men_n343_));
  NA3        u0315(.A(m), .B(men_men_n109_), .C(men_men_n202_), .Y(men_men_n344_));
  NA4        u0316(.A(men_men_n191_), .B(men_men_n85_), .C(g), .D(men_men_n202_), .Y(men_men_n345_));
  OAI210     u0317(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n345_), .Y(men_men_n346_));
  NAi41      u0318(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n347_));
  NA2        u0319(.A(men_men_n51_), .B(men_men_n110_), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n348_), .B(men_men_n347_), .Y(men_men_n349_));
  AOI220     u0321(.A0(men_men_n349_), .A1(b), .B0(men_men_n346_), .B1(men_men_n342_), .Y(men_men_n350_));
  NA3        u0322(.A(men_men_n350_), .B(men_men_n341_), .C(men_men_n335_), .Y(men_men_n351_));
  NO4        u0323(.A(men_men_n351_), .B(men_men_n329_), .C(men_men_n314_), .D(men_men_n308_), .Y(men_men_n352_));
  NA4        u0324(.A(men_men_n352_), .B(men_men_n292_), .C(men_men_n252_), .D(men_men_n187_), .Y(men10));
  NA3        u0325(.A(m), .B(k), .C(i), .Y(men_men_n354_));
  NO3        u0326(.A(men_men_n354_), .B(j), .C(men_men_n203_), .Y(men_men_n355_));
  NOi21      u0327(.An(e), .B(f), .Y(men_men_n356_));
  NO4        u0328(.A(men_men_n145_), .B(men_men_n356_), .C(n), .D(men_men_n107_), .Y(men_men_n357_));
  NAi31      u0329(.An(b), .B(f), .C(c), .Y(men_men_n358_));
  INV        u0330(.A(men_men_n358_), .Y(men_men_n359_));
  NOi32      u0331(.An(k), .Bn(h), .C(j), .Y(men_men_n360_));
  NA2        u0332(.A(men_men_n360_), .B(men_men_n210_), .Y(men_men_n361_));
  NA2        u0333(.A(men_men_n154_), .B(men_men_n361_), .Y(men_men_n362_));
  AOI220     u0334(.A0(men_men_n362_), .A1(men_men_n359_), .B0(men_men_n357_), .B1(men_men_n355_), .Y(men_men_n363_));
  NO3        u0335(.A(n), .B(m), .C(k), .Y(men_men_n364_));
  NA2        u0336(.A(men_men_n364_), .B(j), .Y(men_men_n365_));
  NO3        u0337(.A(men_men_n365_), .B(men_men_n145_), .C(men_men_n202_), .Y(men_men_n366_));
  NO2        u0338(.A(men_men_n163_), .B(k), .Y(men_men_n367_));
  NA4        u0339(.A(n), .B(f), .C(c), .D(men_men_n112_), .Y(men_men_n368_));
  NOi21      u0340(.An(men_men_n367_), .B(men_men_n368_), .Y(men_men_n369_));
  NOi32      u0341(.An(d), .Bn(a), .C(c), .Y(men_men_n370_));
  NA2        u0342(.A(men_men_n370_), .B(men_men_n171_), .Y(men_men_n371_));
  NAi21      u0343(.An(i), .B(g), .Y(men_men_n372_));
  NAi31      u0344(.An(k), .B(m), .C(j), .Y(men_men_n373_));
  NO3        u0345(.A(men_men_n373_), .B(men_men_n372_), .C(n), .Y(men_men_n374_));
  NOi21      u0346(.An(men_men_n374_), .B(men_men_n371_), .Y(men_men_n375_));
  NO3        u0347(.A(men_men_n375_), .B(men_men_n369_), .C(men_men_n366_), .Y(men_men_n376_));
  NO2        u0348(.A(men_men_n368_), .B(men_men_n278_), .Y(men_men_n377_));
  NOi32      u0349(.An(f), .Bn(d), .C(c), .Y(men_men_n378_));
  AOI220     u0350(.A0(men_men_n378_), .A1(men_men_n286_), .B0(men_men_n377_), .B1(men_men_n204_), .Y(men_men_n379_));
  NA3        u0351(.A(men_men_n379_), .B(men_men_n376_), .C(men_men_n363_), .Y(men_men_n380_));
  NA2        u0352(.A(men_men_n233_), .B(d), .Y(men_men_n381_));
  INV        u0353(.A(e), .Y(men_men_n382_));
  NA2        u0354(.A(men_men_n46_), .B(e), .Y(men_men_n383_));
  OAI220     u0355(.A0(men_men_n383_), .A1(men_men_n188_), .B0(men_men_n192_), .B1(men_men_n382_), .Y(men_men_n384_));
  AN2        u0356(.A(g), .B(e), .Y(men_men_n385_));
  NA3        u0357(.A(men_men_n385_), .B(men_men_n191_), .C(i), .Y(men_men_n386_));
  OAI210     u0358(.A0(men_men_n87_), .A1(men_men_n382_), .B0(men_men_n386_), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n387_), .B(men_men_n384_), .Y(men_men_n388_));
  NOi32      u0360(.An(h), .Bn(e), .C(g), .Y(men_men_n389_));
  NA3        u0361(.A(men_men_n389_), .B(men_men_n271_), .C(m), .Y(men_men_n390_));
  NOi21      u0362(.An(g), .B(h), .Y(men_men_n391_));
  AN3        u0363(.A(m), .B(l), .C(i), .Y(men_men_n392_));
  AN3        u0364(.A(h), .B(g), .C(e), .Y(men_men_n393_));
  NA2        u0365(.A(men_men_n393_), .B(men_men_n96_), .Y(men_men_n394_));
  AOI210     u0366(.A0(men_men_n390_), .A1(men_men_n388_), .B0(men_men_n381_), .Y(men_men_n395_));
  NA3        u0367(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n396_));
  NO2        u0368(.A(men_men_n396_), .B(men_men_n381_), .Y(men_men_n397_));
  NA3        u0369(.A(men_men_n370_), .B(men_men_n171_), .C(men_men_n82_), .Y(men_men_n398_));
  NAi31      u0370(.An(b), .B(c), .C(a), .Y(men_men_n399_));
  NO2        u0371(.A(men_men_n399_), .B(n), .Y(men_men_n400_));
  OAI210     u0372(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n401_));
  NO2        u0373(.A(men_men_n401_), .B(men_men_n141_), .Y(men_men_n402_));
  NO3        u0374(.A(men_men_n397_), .B(men_men_n395_), .C(men_men_n380_), .Y(men_men_n403_));
  NA2        u0375(.A(i), .B(g), .Y(men_men_n404_));
  NO3        u0376(.A(men_men_n260_), .B(men_men_n404_), .C(c), .Y(men_men_n405_));
  NOi21      u0377(.An(d), .B(c), .Y(men_men_n406_));
  NA2        u0378(.A(men_men_n406_), .B(a), .Y(men_men_n407_));
  NA3        u0379(.A(i), .B(g), .C(f), .Y(men_men_n408_));
  OR2        u0380(.A(men_men_n408_), .B(men_men_n67_), .Y(men_men_n409_));
  NA3        u0381(.A(men_men_n392_), .B(men_men_n391_), .C(men_men_n171_), .Y(men_men_n410_));
  AOI210     u0382(.A0(men_men_n410_), .A1(men_men_n409_), .B0(men_men_n407_), .Y(men_men_n411_));
  AOI210     u0383(.A0(men_men_n405_), .A1(men_men_n270_), .B0(men_men_n411_), .Y(men_men_n412_));
  OR2        u0384(.A(n), .B(m), .Y(men_men_n413_));
  NO2        u0385(.A(men_men_n413_), .B(men_men_n146_), .Y(men_men_n414_));
  NA2        u0386(.A(men_men_n165_), .B(c), .Y(men_men_n415_));
  INV        u0387(.A(men_men_n348_), .Y(men_men_n416_));
  NA3        u0388(.A(men_men_n416_), .B(men_men_n336_), .C(d), .Y(men_men_n417_));
  NO2        u0389(.A(men_men_n399_), .B(men_men_n49_), .Y(men_men_n418_));
  NO3        u0390(.A(men_men_n62_), .B(men_men_n109_), .C(e), .Y(men_men_n419_));
  NAi21      u0391(.An(k), .B(j), .Y(men_men_n420_));
  NA2        u0392(.A(men_men_n236_), .B(men_men_n420_), .Y(men_men_n421_));
  NA3        u0393(.A(men_men_n421_), .B(men_men_n419_), .C(men_men_n418_), .Y(men_men_n422_));
  NAi21      u0394(.An(e), .B(d), .Y(men_men_n423_));
  INV        u0395(.A(men_men_n423_), .Y(men_men_n424_));
  NO2        u0396(.A(men_men_n237_), .B(men_men_n202_), .Y(men_men_n425_));
  NA2        u0397(.A(men_men_n425_), .B(men_men_n424_), .Y(men_men_n426_));
  NA4        u0398(.A(men_men_n426_), .B(men_men_n422_), .C(men_men_n417_), .D(men_men_n415_), .Y(men_men_n427_));
  NO2        u0399(.A(men_men_n312_), .B(men_men_n202_), .Y(men_men_n428_));
  NA2        u0400(.A(men_men_n428_), .B(men_men_n424_), .Y(men_men_n429_));
  NOi31      u0401(.An(n), .B(m), .C(k), .Y(men_men_n430_));
  AOI220     u0402(.A0(men_men_n430_), .A1(j), .B0(men_men_n210_), .B1(men_men_n50_), .Y(men_men_n431_));
  NAi31      u0403(.An(g), .B(f), .C(c), .Y(men_men_n432_));
  OR3        u0404(.A(men_men_n432_), .B(men_men_n431_), .C(e), .Y(men_men_n433_));
  NA3        u0405(.A(men_men_n433_), .B(men_men_n429_), .C(men_men_n287_), .Y(men_men_n434_));
  NOi41      u0406(.An(men_men_n412_), .B(men_men_n434_), .C(men_men_n427_), .D(men_men_n250_), .Y(men_men_n435_));
  NOi32      u0407(.An(c), .Bn(a), .C(b), .Y(men_men_n436_));
  NA2        u0408(.A(men_men_n436_), .B(men_men_n110_), .Y(men_men_n437_));
  INV        u0409(.A(men_men_n258_), .Y(men_men_n438_));
  AN2        u0410(.A(e), .B(d), .Y(men_men_n439_));
  NA2        u0411(.A(men_men_n439_), .B(men_men_n438_), .Y(men_men_n440_));
  INV        u0412(.A(men_men_n141_), .Y(men_men_n441_));
  NO2        u0413(.A(men_men_n126_), .B(men_men_n41_), .Y(men_men_n442_));
  NO2        u0414(.A(men_men_n62_), .B(e), .Y(men_men_n443_));
  NOi31      u0415(.An(j), .B(k), .C(i), .Y(men_men_n444_));
  NOi21      u0416(.An(men_men_n158_), .B(men_men_n444_), .Y(men_men_n445_));
  NA4        u0417(.A(men_men_n299_), .B(men_men_n445_), .C(men_men_n244_), .D(men_men_n115_), .Y(men_men_n446_));
  AOI220     u0418(.A0(men_men_n446_), .A1(men_men_n443_), .B0(men_men_n442_), .B1(men_men_n441_), .Y(men_men_n447_));
  AOI210     u0419(.A0(men_men_n447_), .A1(men_men_n440_), .B0(men_men_n437_), .Y(men_men_n448_));
  NO2        u0420(.A(men_men_n198_), .B(men_men_n193_), .Y(men_men_n449_));
  NA3        u0421(.A(e), .B(d), .C(c), .Y(men_men_n450_));
  NO2        u0422(.A(men_men_n398_), .B(men_men_n192_), .Y(men_men_n451_));
  NOi21      u0423(.An(men_men_n450_), .B(men_men_n451_), .Y(men_men_n452_));
  AOI210     u0424(.A0(men_men_n253_), .A1(men_men_n449_), .B0(men_men_n452_), .Y(men_men_n453_));
  NO4        u0425(.A(men_men_n177_), .B(men_men_n101_), .C(men_men_n56_), .D(b), .Y(men_men_n454_));
  OR2        u0426(.A(k), .B(j), .Y(men_men_n455_));
  NA2        u0427(.A(l), .B(k), .Y(men_men_n456_));
  AOI210     u0428(.A0(men_men_n219_), .A1(men_men_n315_), .B0(men_men_n82_), .Y(men_men_n457_));
  OR3        u0429(.A(m), .B(men_men_n137_), .C(men_men_n129_), .Y(men_men_n458_));
  NA3        u0430(.A(men_men_n262_), .B(men_men_n124_), .C(men_men_n122_), .Y(men_men_n459_));
  NA2        u0431(.A(men_men_n370_), .B(men_men_n110_), .Y(men_men_n460_));
  NO4        u0432(.A(men_men_n460_), .B(men_men_n93_), .C(men_men_n109_), .D(e), .Y(men_men_n461_));
  NO3        u0433(.A(men_men_n398_), .B(men_men_n90_), .C(men_men_n126_), .Y(men_men_n462_));
  NO4        u0434(.A(men_men_n462_), .B(men_men_n461_), .C(men_men_n459_), .D(men_men_n300_), .Y(men_men_n463_));
  NA2        u0435(.A(men_men_n463_), .B(men_men_n458_), .Y(men_men_n464_));
  NO4        u0436(.A(men_men_n464_), .B(men_men_n454_), .C(men_men_n453_), .D(men_men_n448_), .Y(men_men_n465_));
  NA2        u0437(.A(men_men_n66_), .B(men_men_n63_), .Y(men_men_n466_));
  NOi21      u0438(.An(d), .B(e), .Y(men_men_n467_));
  NAi31      u0439(.An(j), .B(l), .C(i), .Y(men_men_n468_));
  OAI210     u0440(.A0(men_men_n468_), .A1(men_men_n127_), .B0(men_men_n101_), .Y(men_men_n469_));
  NA3        u0441(.A(men_men_n469_), .B(c), .C(men_men_n467_), .Y(men_men_n470_));
  NO2        u0442(.A(men_men_n371_), .B(men_men_n348_), .Y(men_men_n471_));
  NO2        u0443(.A(men_men_n471_), .B(men_men_n174_), .Y(men_men_n472_));
  NA4        u0444(.A(men_men_n472_), .B(men_men_n470_), .C(men_men_n466_), .D(men_men_n228_), .Y(men_men_n473_));
  OAI210     u0445(.A0(men_men_n123_), .A1(men_men_n121_), .B0(n), .Y(men_men_n474_));
  AN2        u0446(.A(men_men_n279_), .B(men_men_n180_), .Y(men_men_n475_));
  XO2        u0447(.A(i), .B(h), .Y(men_men_n476_));
  NA3        u0448(.A(men_men_n476_), .B(men_men_n153_), .C(n), .Y(men_men_n477_));
  NAi41      u0449(.An(men_men_n279_), .B(men_men_n477_), .C(men_men_n431_), .D(men_men_n361_), .Y(men_men_n478_));
  NOi32      u0450(.An(men_men_n478_), .Bn(men_men_n443_), .C(men_men_n255_), .Y(men_men_n479_));
  NAi31      u0451(.An(c), .B(f), .C(d), .Y(men_men_n480_));
  AOI210     u0452(.A0(men_men_n263_), .A1(men_men_n183_), .B0(men_men_n480_), .Y(men_men_n481_));
  NOi21      u0453(.An(men_men_n80_), .B(men_men_n481_), .Y(men_men_n482_));
  NA3        u0454(.A(men_men_n357_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n483_));
  NA2        u0455(.A(men_men_n215_), .B(men_men_n105_), .Y(men_men_n484_));
  AOI210     u0456(.A0(men_men_n334_), .A1(men_men_n35_), .B0(men_men_n450_), .Y(men_men_n485_));
  NOi21      u0457(.An(men_men_n483_), .B(men_men_n485_), .Y(men_men_n486_));
  AO220      u0458(.A0(men_men_n267_), .A1(men_men_n247_), .B0(men_men_n159_), .B1(men_men_n63_), .Y(men_men_n487_));
  NA3        u0459(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n488_));
  NO2        u0460(.A(men_men_n488_), .B(men_men_n407_), .Y(men_men_n489_));
  NO2        u0461(.A(men_men_n489_), .B(men_men_n275_), .Y(men_men_n490_));
  NAi41      u0462(.An(men_men_n487_), .B(men_men_n490_), .C(men_men_n486_), .D(men_men_n482_), .Y(men_men_n491_));
  NO4        u0463(.A(men_men_n491_), .B(men_men_n479_), .C(men_men_n475_), .D(men_men_n473_), .Y(men_men_n492_));
  NA4        u0464(.A(men_men_n492_), .B(men_men_n465_), .C(men_men_n435_), .D(men_men_n403_), .Y(men11));
  NO2        u0465(.A(men_men_n69_), .B(f), .Y(men_men_n494_));
  NA2        u0466(.A(j), .B(g), .Y(men_men_n495_));
  NAi31      u0467(.An(i), .B(m), .C(l), .Y(men_men_n496_));
  NA3        u0468(.A(m), .B(k), .C(j), .Y(men_men_n497_));
  OAI220     u0469(.A0(men_men_n497_), .A1(men_men_n126_), .B0(men_men_n496_), .B1(men_men_n495_), .Y(men_men_n498_));
  NA2        u0470(.A(men_men_n498_), .B(men_men_n494_), .Y(men_men_n499_));
  NOi32      u0471(.An(e), .Bn(b), .C(f), .Y(men_men_n500_));
  NA2        u0472(.A(men_men_n243_), .B(men_men_n110_), .Y(men_men_n501_));
  NA2        u0473(.A(men_men_n46_), .B(j), .Y(men_men_n502_));
  NO2        u0474(.A(men_men_n502_), .B(i), .Y(men_men_n503_));
  NAi31      u0475(.An(d), .B(e), .C(a), .Y(men_men_n504_));
  NO2        u0476(.A(men_men_n504_), .B(n), .Y(men_men_n505_));
  AOI220     u0477(.A0(men_men_n505_), .A1(men_men_n100_), .B0(men_men_n503_), .B1(men_men_n500_), .Y(men_men_n506_));
  NAi41      u0478(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n507_));
  AN2        u0479(.A(men_men_n507_), .B(men_men_n347_), .Y(men_men_n508_));
  AOI210     u0480(.A0(men_men_n508_), .A1(men_men_n371_), .B0(men_men_n256_), .Y(men_men_n509_));
  NA2        u0481(.A(j), .B(i), .Y(men_men_n510_));
  NAi31      u0482(.An(n), .B(m), .C(k), .Y(men_men_n511_));
  NO3        u0483(.A(men_men_n511_), .B(men_men_n510_), .C(men_men_n109_), .Y(men_men_n512_));
  NO2        u0484(.A(n), .B(men_men_n143_), .Y(men_men_n513_));
  NOi32      u0485(.An(g), .Bn(f), .C(i), .Y(men_men_n514_));
  AOI220     u0486(.A0(men_men_n514_), .A1(men_men_n98_), .B0(men_men_n498_), .B1(f), .Y(men_men_n515_));
  NO2        u0487(.A(men_men_n515_), .B(n), .Y(men_men_n516_));
  AOI210     u0488(.A0(men_men_n512_), .A1(men_men_n509_), .B0(men_men_n516_), .Y(men_men_n517_));
  NA2        u0489(.A(men_men_n133_), .B(men_men_n34_), .Y(men_men_n518_));
  OAI220     u0490(.A0(men_men_n518_), .A1(m), .B0(men_men_n502_), .B1(men_men_n219_), .Y(men_men_n519_));
  NOi41      u0491(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n520_));
  NAi32      u0492(.An(e), .Bn(b), .C(c), .Y(men_men_n521_));
  AN2        u0493(.A(men_men_n316_), .B(men_men_n296_), .Y(men_men_n522_));
  NA2        u0494(.A(men_men_n522_), .B(men_men_n521_), .Y(men_men_n523_));
  OA210      u0495(.A0(men_men_n523_), .A1(men_men_n520_), .B0(men_men_n519_), .Y(men_men_n524_));
  OAI220     u0496(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n496_), .B1(men_men_n495_), .Y(men_men_n525_));
  NAi31      u0497(.An(d), .B(c), .C(a), .Y(men_men_n526_));
  NO2        u0498(.A(men_men_n526_), .B(n), .Y(men_men_n527_));
  NA3        u0499(.A(men_men_n527_), .B(men_men_n525_), .C(e), .Y(men_men_n528_));
  NO3        u0500(.A(men_men_n60_), .B(men_men_n49_), .C(men_men_n203_), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n216_), .B(men_men_n107_), .Y(men_men_n530_));
  OAI210     u0502(.A0(men_men_n529_), .A1(men_men_n374_), .B0(men_men_n530_), .Y(men_men_n531_));
  NA2        u0503(.A(men_men_n531_), .B(men_men_n528_), .Y(men_men_n532_));
  NA2        u0504(.A(men_men_n525_), .B(f), .Y(men_men_n533_));
  NAi32      u0505(.An(d), .Bn(a), .C(b), .Y(men_men_n534_));
  NA2        u0506(.A(h), .B(f), .Y(men_men_n535_));
  NO2        u0507(.A(men_men_n535_), .B(men_men_n93_), .Y(men_men_n536_));
  NO3        u0508(.A(men_men_n166_), .B(men_men_n163_), .C(g), .Y(men_men_n537_));
  AOI220     u0509(.A0(men_men_n537_), .A1(c), .B0(men_men_n536_), .B1(m), .Y(men_men_n538_));
  INV        u0510(.A(men_men_n538_), .Y(men_men_n539_));
  AN3        u0511(.A(j), .B(h), .C(g), .Y(men_men_n540_));
  NO2        u0512(.A(men_men_n140_), .B(c), .Y(men_men_n541_));
  NA3        u0513(.A(men_men_n541_), .B(men_men_n540_), .C(men_men_n430_), .Y(men_men_n542_));
  NA3        u0514(.A(f), .B(d), .C(b), .Y(men_men_n543_));
  NO4        u0515(.A(men_men_n543_), .B(men_men_n166_), .C(men_men_n163_), .D(g), .Y(men_men_n544_));
  NAi21      u0516(.An(men_men_n544_), .B(men_men_n542_), .Y(men_men_n545_));
  NO4        u0517(.A(men_men_n545_), .B(men_men_n539_), .C(men_men_n532_), .D(men_men_n524_), .Y(men_men_n546_));
  AN4        u0518(.A(men_men_n546_), .B(men_men_n517_), .C(men_men_n506_), .D(men_men_n499_), .Y(men_men_n547_));
  INV        u0519(.A(k), .Y(men_men_n548_));
  NA3        u0520(.A(l), .B(men_men_n548_), .C(i), .Y(men_men_n549_));
  INV        u0521(.A(men_men_n549_), .Y(men_men_n550_));
  NA4        u0522(.A(men_men_n370_), .B(men_men_n391_), .C(men_men_n171_), .D(men_men_n110_), .Y(men_men_n551_));
  NAi32      u0523(.An(h), .Bn(f), .C(g), .Y(men_men_n552_));
  NAi41      u0524(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n553_));
  OAI210     u0525(.A0(men_men_n504_), .A1(n), .B0(men_men_n553_), .Y(men_men_n554_));
  NA2        u0526(.A(men_men_n554_), .B(m), .Y(men_men_n555_));
  NAi31      u0527(.An(h), .B(g), .C(f), .Y(men_men_n556_));
  OR2        u0528(.A(men_men_n555_), .B(men_men_n552_), .Y(men_men_n557_));
  NO3        u0529(.A(men_men_n552_), .B(men_men_n69_), .C(men_men_n71_), .Y(men_men_n558_));
  NO4        u0530(.A(men_men_n556_), .B(n), .C(men_men_n143_), .D(men_men_n71_), .Y(men_men_n559_));
  OR2        u0531(.A(men_men_n559_), .B(men_men_n558_), .Y(men_men_n560_));
  NAi31      u0532(.An(men_men_n560_), .B(men_men_n557_), .C(men_men_n551_), .Y(men_men_n561_));
  NAi31      u0533(.An(f), .B(h), .C(g), .Y(men_men_n562_));
  NO4        u0534(.A(men_men_n288_), .B(men_men_n562_), .C(men_men_n69_), .D(men_men_n71_), .Y(men_men_n563_));
  NOi32      u0535(.An(d), .Bn(a), .C(e), .Y(men_men_n564_));
  NA2        u0536(.A(men_men_n564_), .B(men_men_n110_), .Y(men_men_n565_));
  NO2        u0537(.A(n), .B(c), .Y(men_men_n566_));
  NA3        u0538(.A(men_men_n566_), .B(men_men_n29_), .C(m), .Y(men_men_n567_));
  NAi32      u0539(.An(n), .Bn(f), .C(m), .Y(men_men_n568_));
  NA3        u0540(.A(men_men_n568_), .B(men_men_n567_), .C(men_men_n565_), .Y(men_men_n569_));
  NOi32      u0541(.An(e), .Bn(a), .C(d), .Y(men_men_n570_));
  AOI210     u0542(.A0(men_men_n29_), .A1(d), .B0(men_men_n570_), .Y(men_men_n571_));
  AOI210     u0543(.A0(men_men_n571_), .A1(men_men_n202_), .B0(men_men_n518_), .Y(men_men_n572_));
  AOI210     u0544(.A0(men_men_n572_), .A1(men_men_n569_), .B0(men_men_n563_), .Y(men_men_n573_));
  INV        u0545(.A(men_men_n573_), .Y(men_men_n574_));
  AOI210     u0546(.A0(men_men_n561_), .A1(men_men_n550_), .B0(men_men_n574_), .Y(men_men_n575_));
  NA2        u0547(.A(men_men_n432_), .B(men_men_n216_), .Y(men_men_n576_));
  NA2        u0548(.A(men_men_n72_), .B(men_men_n110_), .Y(men_men_n577_));
  NO2        u0549(.A(men_men_n577_), .B(men_men_n45_), .Y(men_men_n578_));
  NA2        u0550(.A(men_men_n578_), .B(men_men_n509_), .Y(men_men_n579_));
  INV        u0551(.A(men_men_n579_), .Y(men_men_n580_));
  NA3        u0552(.A(men_men_n520_), .B(men_men_n318_), .C(men_men_n46_), .Y(men_men_n581_));
  NOi32      u0553(.An(e), .Bn(c), .C(f), .Y(men_men_n582_));
  NOi21      u0554(.An(f), .B(g), .Y(men_men_n583_));
  NO2        u0555(.A(men_men_n583_), .B(men_men_n200_), .Y(men_men_n584_));
  AOI220     u0556(.A0(men_men_n584_), .A1(men_men_n367_), .B0(men_men_n582_), .B1(men_men_n165_), .Y(men_men_n585_));
  NA3        u0557(.A(men_men_n585_), .B(men_men_n581_), .C(men_men_n168_), .Y(men_men_n586_));
  AOI210     u0558(.A0(men_men_n508_), .A1(men_men_n371_), .B0(men_men_n280_), .Y(men_men_n587_));
  NA2        u0559(.A(men_men_n587_), .B(men_men_n248_), .Y(men_men_n588_));
  NOi21      u0560(.An(j), .B(l), .Y(men_men_n589_));
  NAi21      u0561(.An(k), .B(h), .Y(men_men_n590_));
  NO2        u0562(.A(men_men_n590_), .B(men_men_n246_), .Y(men_men_n591_));
  NA2        u0563(.A(men_men_n591_), .B(men_men_n589_), .Y(men_men_n592_));
  OR2        u0564(.A(men_men_n592_), .B(men_men_n555_), .Y(men_men_n593_));
  NOi31      u0565(.An(m), .B(n), .C(k), .Y(men_men_n594_));
  NA2        u0566(.A(men_men_n589_), .B(men_men_n594_), .Y(men_men_n595_));
  NO2        u0567(.A(men_men_n371_), .B(men_men_n280_), .Y(men_men_n596_));
  NAi21      u0568(.An(men_men_n595_), .B(men_men_n596_), .Y(men_men_n597_));
  NO2        u0569(.A(men_men_n260_), .B(men_men_n49_), .Y(men_men_n598_));
  NO2        u0570(.A(men_men_n288_), .B(men_men_n562_), .Y(men_men_n599_));
  NO2        u0571(.A(men_men_n504_), .B(men_men_n49_), .Y(men_men_n600_));
  NA2        u0572(.A(men_men_n600_), .B(men_men_n599_), .Y(men_men_n601_));
  NA4        u0573(.A(men_men_n601_), .B(men_men_n597_), .C(men_men_n593_), .D(men_men_n588_), .Y(men_men_n602_));
  NA2        u0574(.A(men_men_n105_), .B(men_men_n36_), .Y(men_men_n603_));
  NO2        u0575(.A(k), .B(men_men_n203_), .Y(men_men_n604_));
  NO2        u0576(.A(men_men_n502_), .B(men_men_n166_), .Y(men_men_n605_));
  NA3        u0577(.A(men_men_n521_), .B(men_men_n255_), .C(men_men_n138_), .Y(men_men_n606_));
  NO3        u0578(.A(men_men_n368_), .B(m), .C(men_men_n85_), .Y(men_men_n607_));
  AOI210     u0579(.A0(men_men_n606_), .A1(men_men_n605_), .B0(men_men_n607_), .Y(men_men_n608_));
  AN3        u0580(.A(f), .B(d), .C(b), .Y(men_men_n609_));
  NAi31      u0581(.An(m), .B(n), .C(k), .Y(men_men_n610_));
  OAI210     u0582(.A0(men_men_n129_), .A1(men_men_n610_), .B0(men_men_n234_), .Y(men_men_n611_));
  NA2        u0583(.A(men_men_n611_), .B(j), .Y(men_men_n612_));
  NA2        u0584(.A(men_men_n612_), .B(men_men_n608_), .Y(men_men_n613_));
  NO4        u0585(.A(men_men_n613_), .B(men_men_n602_), .C(men_men_n586_), .D(men_men_n580_), .Y(men_men_n614_));
  NA2        u0586(.A(men_men_n357_), .B(men_men_n156_), .Y(men_men_n615_));
  NAi31      u0587(.An(g), .B(h), .C(f), .Y(men_men_n616_));
  OA210      u0588(.A0(men_men_n504_), .A1(n), .B0(men_men_n553_), .Y(men_men_n617_));
  NO2        u0589(.A(men_men_n617_), .B(men_men_n89_), .Y(men_men_n618_));
  INV        u0590(.A(men_men_n618_), .Y(men_men_n619_));
  AOI210     u0591(.A0(men_men_n619_), .A1(men_men_n615_), .B0(men_men_n497_), .Y(men_men_n620_));
  NAi21      u0592(.An(h), .B(j), .Y(men_men_n621_));
  OR2        u0593(.A(men_men_n592_), .B(men_men_n69_), .Y(men_men_n622_));
  NA3        u0594(.A(men_men_n494_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n623_));
  AN2        u0595(.A(h), .B(f), .Y(men_men_n624_));
  NA2        u0596(.A(men_men_n624_), .B(men_men_n37_), .Y(men_men_n625_));
  NA2        u0597(.A(men_men_n98_), .B(men_men_n46_), .Y(men_men_n626_));
  OAI220     u0598(.A0(men_men_n626_), .A1(men_men_n310_), .B0(men_men_n625_), .B1(men_men_n437_), .Y(men_men_n627_));
  AOI210     u0599(.A0(men_men_n534_), .A1(men_men_n399_), .B0(men_men_n49_), .Y(men_men_n628_));
  OAI220     u0600(.A0(men_men_n556_), .A1(men_men_n549_), .B0(men_men_n304_), .B1(men_men_n495_), .Y(men_men_n629_));
  AOI210     u0601(.A0(men_men_n629_), .A1(men_men_n628_), .B0(men_men_n627_), .Y(men_men_n630_));
  NA3        u0602(.A(men_men_n630_), .B(men_men_n623_), .C(men_men_n622_), .Y(men_men_n631_));
  NO2        u0603(.A(men_men_n236_), .B(f), .Y(men_men_n632_));
  NA2        u0604(.A(men_men_n307_), .B(men_men_n133_), .Y(men_men_n633_));
  AOI210     u0605(.A0(men_men_n336_), .A1(men_men_n110_), .B0(men_men_n500_), .Y(men_men_n634_));
  OA220      u0606(.A0(men_men_n634_), .A1(men_men_n518_), .B0(men_men_n334_), .B1(men_men_n108_), .Y(men_men_n635_));
  OAI210     u0607(.A0(men_men_n633_), .A1(men_men_n236_), .B0(men_men_n635_), .Y(men_men_n636_));
  NO3        u0608(.A(men_men_n378_), .B(men_men_n180_), .C(men_men_n179_), .Y(men_men_n637_));
  NA2        u0609(.A(men_men_n637_), .B(men_men_n216_), .Y(men_men_n638_));
  NA3        u0610(.A(men_men_n638_), .B(men_men_n238_), .C(j), .Y(men_men_n639_));
  NO3        u0611(.A(men_men_n432_), .B(men_men_n163_), .C(i), .Y(men_men_n640_));
  NA2        u0612(.A(men_men_n436_), .B(men_men_n82_), .Y(men_men_n641_));
  NA3        u0613(.A(men_men_n639_), .B(men_men_n483_), .C(men_men_n376_), .Y(men_men_n642_));
  NO4        u0614(.A(men_men_n642_), .B(men_men_n636_), .C(men_men_n631_), .D(men_men_n620_), .Y(men_men_n643_));
  NA4        u0615(.A(men_men_n643_), .B(men_men_n614_), .C(men_men_n575_), .D(men_men_n547_), .Y(men08));
  NO2        u0616(.A(k), .B(h), .Y(men_men_n645_));
  AO210      u0617(.A0(men_men_n236_), .A1(men_men_n420_), .B0(men_men_n645_), .Y(men_men_n646_));
  NO2        u0618(.A(men_men_n646_), .B(men_men_n278_), .Y(men_men_n647_));
  NA2        u0619(.A(men_men_n582_), .B(men_men_n82_), .Y(men_men_n648_));
  INV        u0620(.A(men_men_n462_), .Y(men_men_n649_));
  NA2        u0621(.A(men_men_n82_), .B(men_men_n107_), .Y(men_men_n650_));
  NO4        u0622(.A(men_men_n354_), .B(men_men_n109_), .C(j), .D(men_men_n203_), .Y(men_men_n651_));
  NA2        u0623(.A(men_men_n543_), .B(men_men_n218_), .Y(men_men_n652_));
  AOI210     u0624(.A0(men_men_n652_), .A1(men_men_n324_), .B0(men_men_n651_), .Y(men_men_n653_));
  AOI210     u0625(.A0(men_men_n543_), .A1(men_men_n150_), .B0(men_men_n82_), .Y(men_men_n654_));
  NA4        u0626(.A(men_men_n205_), .B(men_men_n133_), .C(men_men_n45_), .D(h), .Y(men_men_n655_));
  AN2        u0627(.A(l), .B(k), .Y(men_men_n656_));
  NA4        u0628(.A(men_men_n656_), .B(men_men_n105_), .C(men_men_n71_), .D(men_men_n203_), .Y(men_men_n657_));
  OAI210     u0629(.A0(men_men_n655_), .A1(g), .B0(men_men_n657_), .Y(men_men_n658_));
  NA2        u0630(.A(men_men_n658_), .B(men_men_n654_), .Y(men_men_n659_));
  NA4        u0631(.A(men_men_n659_), .B(men_men_n653_), .C(men_men_n649_), .D(men_men_n326_), .Y(men_men_n660_));
  AN2        u0632(.A(men_men_n505_), .B(men_men_n94_), .Y(men_men_n661_));
  NO4        u0633(.A(men_men_n163_), .B(k), .C(men_men_n109_), .D(g), .Y(men_men_n662_));
  AOI210     u0634(.A0(men_men_n662_), .A1(men_men_n652_), .B0(men_men_n489_), .Y(men_men_n663_));
  NO2        u0635(.A(men_men_n38_), .B(men_men_n202_), .Y(men_men_n664_));
  NA2        u0636(.A(men_men_n584_), .B(men_men_n323_), .Y(men_men_n665_));
  NAi31      u0637(.An(men_men_n661_), .B(men_men_n665_), .C(men_men_n663_), .Y(men_men_n666_));
  NO2        u0638(.A(men_men_n508_), .B(men_men_n35_), .Y(men_men_n667_));
  OAI210     u0639(.A0(men_men_n521_), .A1(men_men_n47_), .B0(men_men_n129_), .Y(men_men_n668_));
  NO2        u0640(.A(men_men_n456_), .B(men_men_n127_), .Y(men_men_n669_));
  AOI210     u0641(.A0(men_men_n669_), .A1(men_men_n668_), .B0(men_men_n667_), .Y(men_men_n670_));
  NO3        u0642(.A(men_men_n294_), .B(men_men_n126_), .C(men_men_n41_), .Y(men_men_n671_));
  NAi21      u0643(.An(men_men_n671_), .B(men_men_n657_), .Y(men_men_n672_));
  NA2        u0644(.A(men_men_n646_), .B(men_men_n130_), .Y(men_men_n673_));
  AOI220     u0645(.A0(men_men_n673_), .A1(men_men_n377_), .B0(men_men_n672_), .B1(men_men_n74_), .Y(men_men_n674_));
  OAI210     u0646(.A0(men_men_n670_), .A1(men_men_n85_), .B0(men_men_n674_), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n336_), .B(men_men_n43_), .Y(men_men_n676_));
  NA3        u0648(.A(men_men_n638_), .B(men_men_n311_), .C(men_men_n360_), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n656_), .B(men_men_n210_), .Y(men_men_n678_));
  NO2        u0650(.A(men_men_n678_), .B(men_men_n306_), .Y(men_men_n679_));
  AOI210     u0651(.A0(men_men_n679_), .A1(men_men_n632_), .B0(men_men_n461_), .Y(men_men_n680_));
  NA3        u0652(.A(m), .B(l), .C(k), .Y(men_men_n681_));
  NO2        u0653(.A(men_men_n507_), .B(men_men_n256_), .Y(men_men_n682_));
  NOi21      u0654(.An(men_men_n682_), .B(men_men_n501_), .Y(men_men_n683_));
  INV        u0655(.A(men_men_n683_), .Y(men_men_n684_));
  NA4        u0656(.A(men_men_n684_), .B(men_men_n680_), .C(men_men_n677_), .D(men_men_n676_), .Y(men_men_n685_));
  NO4        u0657(.A(men_men_n685_), .B(men_men_n675_), .C(men_men_n666_), .D(men_men_n660_), .Y(men_men_n686_));
  NOi31      u0658(.An(g), .B(h), .C(f), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n600_), .B(men_men_n687_), .Y(men_men_n688_));
  OR2        u0660(.A(men_men_n688_), .B(men_men_n510_), .Y(men_men_n689_));
  NO3        u0661(.A(men_men_n371_), .B(men_men_n495_), .C(h), .Y(men_men_n690_));
  AOI210     u0662(.A0(men_men_n690_), .A1(men_men_n110_), .B0(men_men_n471_), .Y(men_men_n691_));
  NA3        u0663(.A(men_men_n691_), .B(men_men_n689_), .C(men_men_n235_), .Y(men_men_n692_));
  NA2        u0664(.A(men_men_n656_), .B(men_men_n71_), .Y(men_men_n693_));
  NO4        u0665(.A(men_men_n637_), .B(men_men_n163_), .C(n), .D(i), .Y(men_men_n694_));
  NOi21      u0666(.An(h), .B(j), .Y(men_men_n695_));
  NA2        u0667(.A(men_men_n695_), .B(f), .Y(men_men_n696_));
  NO2        u0668(.A(men_men_n694_), .B(men_men_n640_), .Y(men_men_n697_));
  NO2        u0669(.A(men_men_n697_), .B(men_men_n693_), .Y(men_men_n698_));
  AOI210     u0670(.A0(men_men_n692_), .A1(l), .B0(men_men_n698_), .Y(men_men_n699_));
  NO2        u0671(.A(j), .B(i), .Y(men_men_n700_));
  NA3        u0672(.A(men_men_n700_), .B(men_men_n78_), .C(l), .Y(men_men_n701_));
  NA2        u0673(.A(men_men_n700_), .B(men_men_n33_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n393_), .B(men_men_n117_), .Y(men_men_n703_));
  OA220      u0675(.A0(men_men_n703_), .A1(men_men_n702_), .B0(men_men_n701_), .B1(men_men_n555_), .Y(men_men_n704_));
  NO2        u0676(.A(men_men_n49_), .B(men_men_n107_), .Y(men_men_n705_));
  NO3        u0677(.A(n), .B(men_men_n143_), .C(men_men_n71_), .Y(men_men_n706_));
  NO2        u0678(.A(men_men_n688_), .B(men_men_n60_), .Y(men_men_n707_));
  NO2        u0679(.A(men_men_n278_), .B(men_men_n40_), .Y(men_men_n708_));
  AOI210     u0680(.A0(men_men_n500_), .A1(n), .B0(men_men_n520_), .Y(men_men_n709_));
  NA2        u0681(.A(men_men_n709_), .B(men_men_n522_), .Y(men_men_n710_));
  AN3        u0682(.A(men_men_n710_), .B(men_men_n708_), .C(men_men_n97_), .Y(men_men_n711_));
  NA2        u0683(.A(men_men_n576_), .B(men_men_n286_), .Y(men_men_n712_));
  NAi21      u0684(.An(men_men_n571_), .B(men_men_n91_), .Y(men_men_n713_));
  NA2        u0685(.A(men_men_n713_), .B(men_men_n712_), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n671_), .B(men_men_n654_), .Y(men_men_n715_));
  NO2        u0687(.A(men_men_n681_), .B(men_men_n89_), .Y(men_men_n716_));
  NA2        u0688(.A(men_men_n716_), .B(men_men_n554_), .Y(men_men_n717_));
  NO2        u0689(.A(men_men_n556_), .B(men_men_n113_), .Y(men_men_n718_));
  NA2        u0690(.A(men_men_n718_), .B(men_men_n628_), .Y(men_men_n719_));
  NA3        u0691(.A(men_men_n719_), .B(men_men_n717_), .C(men_men_n715_), .Y(men_men_n720_));
  OR4        u0692(.A(men_men_n720_), .B(men_men_n714_), .C(men_men_n711_), .D(men_men_n707_), .Y(men_men_n721_));
  NA3        u0693(.A(men_men_n709_), .B(men_men_n522_), .C(men_men_n521_), .Y(men_men_n722_));
  NA4        u0694(.A(men_men_n722_), .B(men_men_n205_), .C(men_men_n420_), .D(men_men_n34_), .Y(men_men_n723_));
  OAI220     u0695(.A0(men_men_n655_), .A1(men_men_n648_), .B0(men_men_n310_), .B1(men_men_n38_), .Y(men_men_n724_));
  INV        u0696(.A(men_men_n724_), .Y(men_men_n725_));
  NA3        u0697(.A(men_men_n514_), .B(men_men_n271_), .C(h), .Y(men_men_n726_));
  NOi21      u0698(.An(men_men_n628_), .B(men_men_n726_), .Y(men_men_n727_));
  OAI220     u0699(.A0(men_men_n726_), .A1(men_men_n567_), .B0(men_men_n701_), .B1(men_men_n69_), .Y(men_men_n728_));
  INV        u0700(.A(men_men_n728_), .Y(men_men_n729_));
  NAi41      u0701(.An(men_men_n727_), .B(men_men_n729_), .C(men_men_n725_), .D(men_men_n723_), .Y(men_men_n730_));
  OR2        u0702(.A(men_men_n716_), .B(men_men_n94_), .Y(men_men_n731_));
  NA2        u0703(.A(men_men_n731_), .B(men_men_n223_), .Y(men_men_n732_));
  INV        u0704(.A(men_men_n617_), .Y(men_men_n733_));
  INV        u0705(.A(men_men_n313_), .Y(men_men_n734_));
  OAI210     u0706(.A0(men_men_n681_), .A1(men_men_n616_), .B0(men_men_n488_), .Y(men_men_n735_));
  NO2        u0707(.A(men_men_n726_), .B(men_men_n460_), .Y(men_men_n736_));
  NO2        u0708(.A(men_men_n735_), .B(men_men_n736_), .Y(men_men_n737_));
  NA3        u0709(.A(men_men_n737_), .B(men_men_n734_), .C(men_men_n732_), .Y(men_men_n738_));
  NOi41      u0710(.An(men_men_n704_), .B(men_men_n738_), .C(men_men_n730_), .D(men_men_n721_), .Y(men_men_n739_));
  OR2        u0711(.A(men_men_n655_), .B(men_men_n218_), .Y(men_men_n740_));
  NO3        u0712(.A(men_men_n319_), .B(men_men_n280_), .C(men_men_n109_), .Y(men_men_n741_));
  INV        u0713(.A(men_men_n741_), .Y(men_men_n742_));
  NA2        u0714(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n743_));
  NO3        u0715(.A(men_men_n743_), .B(men_men_n702_), .C(men_men_n260_), .Y(men_men_n744_));
  INV        u0716(.A(men_men_n744_), .Y(men_men_n745_));
  NA4        u0717(.A(men_men_n745_), .B(men_men_n742_), .C(men_men_n740_), .D(men_men_n379_), .Y(men_men_n746_));
  OR2        u0718(.A(men_men_n616_), .B(men_men_n90_), .Y(men_men_n747_));
  NO2        u0719(.A(men_men_n1368_), .B(n), .Y(men_men_n748_));
  OAI220     u0720(.A0(n), .A1(men_men_n747_), .B0(men_men_n726_), .B1(men_men_n565_), .Y(men_men_n749_));
  NO2        u0721(.A(men_men_n306_), .B(men_men_n113_), .Y(men_men_n750_));
  NOi21      u0722(.An(men_men_n750_), .B(men_men_n154_), .Y(men_men_n751_));
  NO2        u0723(.A(men_men_n637_), .B(n), .Y(men_men_n752_));
  NA2        u0724(.A(men_men_n752_), .B(men_men_n647_), .Y(men_men_n753_));
  NO2        u0725(.A(men_men_n301_), .B(men_men_n222_), .Y(men_men_n754_));
  OAI210     u0726(.A0(men_men_n94_), .A1(men_men_n91_), .B0(men_men_n754_), .Y(men_men_n755_));
  NA2        u0727(.A(men_men_n117_), .B(men_men_n82_), .Y(men_men_n756_));
  AOI210     u0728(.A0(men_men_n396_), .A1(men_men_n390_), .B0(men_men_n756_), .Y(men_men_n757_));
  NAi21      u0729(.An(men_men_n757_), .B(men_men_n755_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n679_), .B(men_men_n34_), .Y(men_men_n759_));
  NA2        u0731(.A(men_men_n662_), .B(men_men_n325_), .Y(men_men_n760_));
  OAI210     u0732(.A0(men_men_n559_), .A1(men_men_n558_), .B0(men_men_n337_), .Y(men_men_n761_));
  AN2        u0733(.A(men_men_n761_), .B(men_men_n760_), .Y(men_men_n762_));
  NAi41      u0734(.An(men_men_n758_), .B(men_men_n762_), .C(men_men_n759_), .D(men_men_n753_), .Y(men_men_n763_));
  NO4        u0735(.A(men_men_n763_), .B(men_men_n751_), .C(men_men_n749_), .D(men_men_n746_), .Y(men_men_n764_));
  NA4        u0736(.A(men_men_n764_), .B(men_men_n739_), .C(men_men_n699_), .D(men_men_n686_), .Y(men09));
  INV        u0737(.A(men_men_n118_), .Y(men_men_n766_));
  NA2        u0738(.A(f), .B(e), .Y(men_men_n767_));
  NO2        u0739(.A(men_men_n214_), .B(men_men_n109_), .Y(men_men_n768_));
  NA2        u0740(.A(men_men_n768_), .B(g), .Y(men_men_n769_));
  NA4        u0741(.A(men_men_n288_), .B(men_men_n445_), .C(men_men_n244_), .D(men_men_n115_), .Y(men_men_n770_));
  AOI210     u0742(.A0(men_men_n770_), .A1(g), .B0(men_men_n442_), .Y(men_men_n771_));
  AOI210     u0743(.A0(men_men_n771_), .A1(men_men_n769_), .B0(men_men_n767_), .Y(men_men_n772_));
  NA2        u0744(.A(men_men_n414_), .B(e), .Y(men_men_n773_));
  NO2        u0745(.A(men_men_n773_), .B(men_men_n480_), .Y(men_men_n774_));
  AOI210     u0746(.A0(men_men_n772_), .A1(men_men_n766_), .B0(men_men_n774_), .Y(men_men_n775_));
  NO2        u0747(.A(men_men_n192_), .B(men_men_n202_), .Y(men_men_n776_));
  NA3        u0748(.A(m), .B(l), .C(i), .Y(men_men_n777_));
  OAI220     u0749(.A0(men_men_n556_), .A1(men_men_n777_), .B0(men_men_n330_), .B1(men_men_n496_), .Y(men_men_n778_));
  NA4        u0750(.A(men_men_n86_), .B(men_men_n85_), .C(g), .D(f), .Y(men_men_n779_));
  NAi31      u0751(.An(men_men_n778_), .B(men_men_n779_), .C(men_men_n409_), .Y(men_men_n780_));
  OR2        u0752(.A(men_men_n780_), .B(men_men_n776_), .Y(men_men_n781_));
  NA3        u0753(.A(men_men_n747_), .B(men_men_n533_), .C(men_men_n488_), .Y(men_men_n782_));
  OA210      u0754(.A0(men_men_n782_), .A1(men_men_n781_), .B0(men_men_n748_), .Y(men_men_n783_));
  INV        u0755(.A(men_men_n316_), .Y(men_men_n784_));
  NO2        u0756(.A(men_men_n123_), .B(men_men_n121_), .Y(men_men_n785_));
  NO2        u0757(.A(m), .B(men_men_n562_), .Y(men_men_n786_));
  NA2        u0758(.A(men_men_n320_), .B(men_men_n322_), .Y(men_men_n787_));
  OAI210     u0759(.A0(men_men_n192_), .A1(men_men_n202_), .B0(men_men_n787_), .Y(men_men_n788_));
  NA2        u0760(.A(men_men_n786_), .B(men_men_n784_), .Y(men_men_n789_));
  NA2        u0761(.A(men_men_n178_), .B(men_men_n31_), .Y(men_men_n790_));
  NA4        u0762(.A(men_men_n790_), .B(men_men_n789_), .C(men_men_n585_), .D(men_men_n80_), .Y(men_men_n791_));
  INV        u0763(.A(men_men_n552_), .Y(men_men_n792_));
  NA2        u0764(.A(men_men_n792_), .B(men_men_n178_), .Y(men_men_n793_));
  NA2        u0765(.A(f), .B(m), .Y(men_men_n794_));
  NO2        u0766(.A(men_men_n794_), .B(men_men_n52_), .Y(men_men_n795_));
  NOi32      u0767(.An(g), .Bn(f), .C(d), .Y(men_men_n796_));
  NA3        u0768(.A(men_men_n796_), .B(men_men_n566_), .C(m), .Y(men_men_n797_));
  NOi21      u0769(.An(men_men_n289_), .B(men_men_n797_), .Y(men_men_n798_));
  AOI210     u0770(.A0(men_men_n795_), .A1(men_men_n513_), .B0(men_men_n798_), .Y(men_men_n799_));
  NA3        u0771(.A(men_men_n288_), .B(men_men_n244_), .C(men_men_n115_), .Y(men_men_n800_));
  AN2        u0772(.A(f), .B(d), .Y(men_men_n801_));
  NA3        u0773(.A(a), .B(men_men_n801_), .C(men_men_n82_), .Y(men_men_n802_));
  NO3        u0774(.A(men_men_n802_), .B(men_men_n71_), .C(men_men_n203_), .Y(men_men_n803_));
  NO2        u0775(.A(men_men_n266_), .B(men_men_n56_), .Y(men_men_n804_));
  NA2        u0776(.A(men_men_n800_), .B(men_men_n803_), .Y(men_men_n805_));
  NAi31      u0777(.An(men_men_n459_), .B(men_men_n805_), .C(men_men_n793_), .Y(men_men_n806_));
  NO4        u0778(.A(men_men_n583_), .B(men_men_n127_), .C(men_men_n306_), .D(men_men_n146_), .Y(men_men_n807_));
  NO2        u0779(.A(men_men_n610_), .B(men_men_n306_), .Y(men_men_n808_));
  AN2        u0780(.A(men_men_n808_), .B(men_men_n632_), .Y(men_men_n809_));
  NO3        u0781(.A(men_men_n809_), .B(men_men_n807_), .C(men_men_n220_), .Y(men_men_n810_));
  NO2        u0782(.A(men_men_n802_), .B(men_men_n401_), .Y(men_men_n811_));
  NOi21      u0783(.An(men_men_n212_), .B(men_men_n811_), .Y(men_men_n812_));
  NA2        u0784(.A(c), .B(men_men_n112_), .Y(men_men_n813_));
  NO2        u0785(.A(men_men_n813_), .B(men_men_n382_), .Y(men_men_n814_));
  NA3        u0786(.A(men_men_n814_), .B(men_men_n478_), .C(f), .Y(men_men_n815_));
  OR2        u0787(.A(men_men_n616_), .B(men_men_n511_), .Y(men_men_n816_));
  INV        u0788(.A(men_men_n816_), .Y(men_men_n817_));
  NA2        u0789(.A(b), .B(men_men_n817_), .Y(men_men_n818_));
  NA4        u0790(.A(men_men_n818_), .B(men_men_n815_), .C(men_men_n812_), .D(men_men_n810_), .Y(men_men_n819_));
  NO4        u0791(.A(men_men_n819_), .B(men_men_n806_), .C(men_men_n791_), .D(men_men_n783_), .Y(men_men_n820_));
  OR2        u0792(.A(men_men_n802_), .B(men_men_n71_), .Y(men_men_n821_));
  NA2        u0793(.A(men_men_n109_), .B(j), .Y(men_men_n822_));
  NA2        u0794(.A(men_men_n768_), .B(g), .Y(men_men_n823_));
  AOI210     u0795(.A0(men_men_n823_), .A1(men_men_n272_), .B0(men_men_n821_), .Y(men_men_n824_));
  NO2        u0796(.A(men_men_n130_), .B(men_men_n127_), .Y(men_men_n825_));
  NO2        u0797(.A(men_men_n216_), .B(men_men_n213_), .Y(men_men_n826_));
  AOI220     u0798(.A0(men_men_n826_), .A1(men_men_n215_), .B0(men_men_n283_), .B1(men_men_n825_), .Y(men_men_n827_));
  NO2        u0799(.A(men_men_n401_), .B(men_men_n767_), .Y(men_men_n828_));
  NA2        u0800(.A(men_men_n828_), .B(men_men_n527_), .Y(men_men_n829_));
  NA2        u0801(.A(men_men_n829_), .B(men_men_n827_), .Y(men_men_n830_));
  NA2        u0802(.A(e), .B(d), .Y(men_men_n831_));
  OAI220     u0803(.A0(men_men_n831_), .A1(c), .B0(men_men_n301_), .B1(d), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n170_), .B(men_men_n216_), .Y(men_men_n833_));
  AOI210     u0805(.A0(men_men_n584_), .A1(men_men_n323_), .B0(men_men_n833_), .Y(men_men_n834_));
  NA2        u0806(.A(men_men_n266_), .B(men_men_n158_), .Y(men_men_n835_));
  NA2        u0807(.A(men_men_n803_), .B(men_men_n835_), .Y(men_men_n836_));
  NA2        u0808(.A(men_men_n836_), .B(men_men_n834_), .Y(men_men_n837_));
  NO3        u0809(.A(men_men_n837_), .B(men_men_n830_), .C(men_men_n824_), .Y(men_men_n838_));
  OR2        u0810(.A(men_men_n648_), .B(men_men_n206_), .Y(men_men_n839_));
  OAI210     u0811(.A0(men_men_n768_), .A1(men_men_n835_), .B0(men_men_n796_), .Y(men_men_n840_));
  NO2        u0812(.A(men_men_n840_), .B(men_men_n567_), .Y(men_men_n841_));
  AOI210     u0813(.A0(men_men_n114_), .A1(men_men_n113_), .B0(men_men_n243_), .Y(men_men_n842_));
  NOi31      u0814(.An(men_men_n513_), .B(men_men_n794_), .C(men_men_n272_), .Y(men_men_n843_));
  INV        u0815(.A(men_men_n841_), .Y(men_men_n844_));
  AO210      u0816(.A0(men_men_n425_), .A1(men_men_n695_), .B0(men_men_n165_), .Y(men_men_n845_));
  OAI210     u0817(.A0(men_men_n845_), .A1(men_men_n428_), .B0(men_men_n832_), .Y(men_men_n846_));
  AN3        u0818(.A(men_men_n846_), .B(men_men_n844_), .C(men_men_n839_), .Y(men_men_n847_));
  NA4        u0819(.A(men_men_n847_), .B(men_men_n838_), .C(men_men_n820_), .D(men_men_n775_), .Y(men12));
  NO2        u0820(.A(men_men_n423_), .B(c), .Y(men_men_n849_));
  NO4        u0821(.A(men_men_n413_), .B(men_men_n236_), .C(men_men_n548_), .D(men_men_n203_), .Y(men_men_n850_));
  NA2        u0822(.A(men_men_n850_), .B(men_men_n849_), .Y(men_men_n851_));
  NO2        u0823(.A(men_men_n423_), .B(men_men_n112_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n785_), .B(men_men_n330_), .Y(men_men_n853_));
  NO2        u0825(.A(men_men_n616_), .B(men_men_n354_), .Y(men_men_n854_));
  AOI220     u0826(.A0(men_men_n854_), .A1(men_men_n1373_), .B0(men_men_n853_), .B1(men_men_n852_), .Y(men_men_n855_));
  NA3        u0827(.A(men_men_n855_), .B(men_men_n851_), .C(men_men_n412_), .Y(men_men_n856_));
  AOI210     u0828(.A0(men_men_n219_), .A1(men_men_n315_), .B0(men_men_n189_), .Y(men_men_n857_));
  BUFFER     u0829(.A(men_men_n857_), .Y(men_men_n858_));
  AOI210     u0830(.A0(men_men_n312_), .A1(men_men_n365_), .B0(men_men_n203_), .Y(men_men_n859_));
  OAI210     u0831(.A0(men_men_n859_), .A1(men_men_n858_), .B0(men_men_n378_), .Y(men_men_n860_));
  NO2        u0832(.A(men_men_n603_), .B(men_men_n246_), .Y(men_men_n861_));
  NO2        u0833(.A(men_men_n556_), .B(men_men_n777_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n754_), .B(men_men_n861_), .Y(men_men_n863_));
  NO2        u0835(.A(men_men_n145_), .B(men_men_n222_), .Y(men_men_n864_));
  NA3        u0836(.A(men_men_n864_), .B(men_men_n225_), .C(i), .Y(men_men_n865_));
  NA3        u0837(.A(men_men_n865_), .B(men_men_n863_), .C(men_men_n860_), .Y(men_men_n866_));
  OR2        u0838(.A(men_men_n302_), .B(men_men_n852_), .Y(men_men_n867_));
  NO3        u0839(.A(men_men_n127_), .B(men_men_n146_), .C(men_men_n203_), .Y(men_men_n868_));
  NA2        u0840(.A(men_men_n868_), .B(men_men_n500_), .Y(men_men_n869_));
  NA4        u0841(.A(men_men_n414_), .B(men_men_n406_), .C(men_men_n171_), .D(g), .Y(men_men_n870_));
  NA2        u0842(.A(men_men_n870_), .B(men_men_n869_), .Y(men_men_n871_));
  NO4        u0843(.A(men_men_n618_), .B(men_men_n871_), .C(men_men_n866_), .D(men_men_n856_), .Y(men_men_n872_));
  NO2        u0844(.A(men_men_n344_), .B(men_men_n343_), .Y(men_men_n873_));
  NA2        u0845(.A(men_men_n553_), .B(men_men_n69_), .Y(men_men_n874_));
  NA2        u0846(.A(men_men_n521_), .B(men_men_n138_), .Y(men_men_n875_));
  NOi21      u0847(.An(men_men_n34_), .B(men_men_n610_), .Y(men_men_n876_));
  AOI220     u0848(.A0(men_men_n876_), .A1(men_men_n875_), .B0(men_men_n874_), .B1(men_men_n873_), .Y(men_men_n877_));
  OAI210     u0849(.A0(men_men_n234_), .A1(men_men_n45_), .B0(men_men_n877_), .Y(men_men_n878_));
  NA2        u0850(.A(men_men_n405_), .B(men_men_n248_), .Y(men_men_n879_));
  NO3        u0851(.A(men_men_n756_), .B(men_men_n87_), .C(men_men_n382_), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n879_), .B(men_men_n298_), .Y(men_men_n881_));
  NO2        u0853(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n882_));
  NO2        u0854(.A(men_men_n474_), .B(men_men_n280_), .Y(men_men_n883_));
  NO2        u0855(.A(men_men_n883_), .B(men_men_n340_), .Y(men_men_n884_));
  NO2        u0856(.A(men_men_n884_), .B(men_men_n138_), .Y(men_men_n885_));
  INV        u0857(.A(men_men_n341_), .Y(men_men_n886_));
  NO4        u0858(.A(men_men_n886_), .B(men_men_n885_), .C(men_men_n881_), .D(men_men_n878_), .Y(men_men_n887_));
  NA2        u0859(.A(men_men_n323_), .B(g), .Y(men_men_n888_));
  NA2        u0860(.A(men_men_n156_), .B(i), .Y(men_men_n889_));
  NA2        u0861(.A(men_men_n46_), .B(i), .Y(men_men_n890_));
  OAI220     u0862(.A0(men_men_n890_), .A1(men_men_n188_), .B0(men_men_n889_), .B1(men_men_n90_), .Y(men_men_n891_));
  AOI210     u0863(.A0(men_men_n392_), .A1(men_men_n37_), .B0(men_men_n891_), .Y(men_men_n892_));
  NO2        u0864(.A(men_men_n138_), .B(men_men_n82_), .Y(men_men_n893_));
  OR2        u0865(.A(men_men_n893_), .B(men_men_n520_), .Y(men_men_n894_));
  NA2        u0866(.A(men_men_n521_), .B(men_men_n358_), .Y(men_men_n895_));
  AOI210     u0867(.A0(men_men_n895_), .A1(n), .B0(men_men_n894_), .Y(men_men_n896_));
  OAI220     u0868(.A0(men_men_n896_), .A1(men_men_n888_), .B0(men_men_n892_), .B1(men_men_n310_), .Y(men_men_n897_));
  NO2        u0869(.A(men_men_n616_), .B(men_men_n468_), .Y(men_men_n898_));
  NA3        u0870(.A(men_men_n320_), .B(men_men_n589_), .C(i), .Y(men_men_n899_));
  OAI210     u0871(.A0(men_men_n408_), .A1(men_men_n288_), .B0(men_men_n899_), .Y(men_men_n900_));
  OAI220     u0872(.A0(men_men_n900_), .A1(men_men_n898_), .B0(men_men_n628_), .B1(men_men_n706_), .Y(men_men_n901_));
  NA2        u0873(.A(men_men_n570_), .B(men_men_n110_), .Y(men_men_n902_));
  NA3        u0874(.A(men_men_n589_), .B(men_men_n78_), .C(i), .Y(men_men_n903_));
  OA220      u0875(.A0(men_men_n903_), .A1(men_men_n902_), .B0(men_men_n288_), .B1(men_men_n555_), .Y(men_men_n904_));
  NA3        u0876(.A(men_men_n303_), .B(men_men_n114_), .C(g), .Y(men_men_n905_));
  AOI210     u0877(.A0(men_men_n625_), .A1(men_men_n905_), .B0(m), .Y(men_men_n906_));
  OAI210     u0878(.A0(men_men_n906_), .A1(men_men_n853_), .B0(men_men_n302_), .Y(men_men_n907_));
  NA2        u0879(.A(men_men_n779_), .B(men_men_n409_), .Y(men_men_n908_));
  NA2        u0880(.A(i), .B(men_men_n75_), .Y(men_men_n909_));
  NA3        u0881(.A(men_men_n909_), .B(men_men_n903_), .C(men_men_n288_), .Y(men_men_n910_));
  AOI210     u0882(.A0(men_men_n910_), .A1(men_men_n241_), .B0(men_men_n908_), .Y(men_men_n911_));
  NA4        u0883(.A(men_men_n911_), .B(men_men_n907_), .C(men_men_n904_), .D(men_men_n901_), .Y(men_men_n912_));
  NA2        u0884(.A(men_men_n861_), .B(men_men_n223_), .Y(men_men_n913_));
  NO2        u0885(.A(men_men_n431_), .B(men_men_n203_), .Y(men_men_n914_));
  AOI220     u0886(.A0(men_men_n914_), .A1(men_men_n359_), .B0(men_men_n867_), .B1(men_men_n207_), .Y(men_men_n915_));
  AOI220     u0887(.A0(men_men_n854_), .A1(men_men_n864_), .B0(men_men_n554_), .B1(men_men_n88_), .Y(men_men_n916_));
  NA3        u0888(.A(men_men_n916_), .B(men_men_n915_), .C(men_men_n913_), .Y(men_men_n917_));
  INV        u0889(.A(men_men_n862_), .Y(men_men_n918_));
  NO2        u0890(.A(men_men_n386_), .B(men_men_n756_), .Y(men_men_n919_));
  OAI210     u0891(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n106_), .Y(men_men_n920_));
  AOI210     u0892(.A0(men_men_n920_), .A1(men_men_n505_), .B0(men_men_n919_), .Y(men_men_n921_));
  NA2        u0893(.A(men_men_n906_), .B(men_men_n852_), .Y(men_men_n922_));
  NO3        u0894(.A(men_men_n822_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n923_));
  AOI220     u0895(.A0(men_men_n923_), .A1(men_men_n587_), .B0(men_men_n605_), .B1(men_men_n500_), .Y(men_men_n924_));
  NA4        u0896(.A(men_men_n924_), .B(men_men_n922_), .C(men_men_n921_), .D(men_men_n918_), .Y(men_men_n925_));
  NO4        u0897(.A(men_men_n925_), .B(men_men_n917_), .C(men_men_n912_), .D(men_men_n897_), .Y(men_men_n926_));
  NAi31      u0898(.An(men_men_n134_), .B(men_men_n393_), .C(n), .Y(men_men_n927_));
  NO3        u0899(.A(men_men_n121_), .B(men_men_n318_), .C(k), .Y(men_men_n928_));
  NA2        u0900(.A(men_men_n462_), .B(i), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n929_), .B(men_men_n927_), .Y(men_men_n930_));
  NA2        u0902(.A(men_men_n216_), .B(men_men_n162_), .Y(men_men_n931_));
  NO3        u0903(.A(men_men_n286_), .B(men_men_n414_), .C(men_men_n165_), .Y(men_men_n932_));
  NOi21      u0904(.An(men_men_n931_), .B(men_men_n932_), .Y(men_men_n933_));
  NAi21      u0905(.An(men_men_n521_), .B(men_men_n914_), .Y(men_men_n934_));
  NO3        u0906(.A(men_men_n408_), .B(men_men_n288_), .C(men_men_n71_), .Y(men_men_n935_));
  AOI220     u0907(.A0(men_men_n935_), .A1(a), .B0(men_men_n454_), .B1(g), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n936_), .B(men_men_n934_), .Y(men_men_n937_));
  NA2        u0909(.A(men_men_n857_), .B(men_men_n849_), .Y(men_men_n938_));
  NA2        u0910(.A(men_men_n494_), .B(men_men_n355_), .Y(men_men_n939_));
  OAI220     u0911(.A0(men_men_n854_), .A1(men_men_n862_), .B0(men_men_n513_), .B1(men_men_n400_), .Y(men_men_n940_));
  NA4        u0912(.A(men_men_n940_), .B(men_men_n939_), .C(men_men_n938_), .D(men_men_n581_), .Y(men_men_n941_));
  OAI210     u0913(.A0(men_men_n857_), .A1(men_men_n850_), .B0(men_men_n931_), .Y(men_men_n942_));
  NA3        u0914(.A(men_men_n895_), .B(men_men_n457_), .C(men_men_n46_), .Y(men_men_n943_));
  AOI210     u0915(.A0(men_men_n357_), .A1(men_men_n355_), .B0(men_men_n309_), .Y(men_men_n944_));
  NA4        u0916(.A(men_men_n944_), .B(men_men_n943_), .C(men_men_n942_), .D(men_men_n257_), .Y(men_men_n945_));
  OR2        u0917(.A(men_men_n945_), .B(men_men_n941_), .Y(men_men_n946_));
  NO4        u0918(.A(men_men_n946_), .B(men_men_n937_), .C(men_men_n933_), .D(men_men_n930_), .Y(men_men_n947_));
  NA4        u0919(.A(men_men_n947_), .B(men_men_n926_), .C(men_men_n887_), .D(men_men_n872_), .Y(men13));
  NA2        u0920(.A(men_men_n46_), .B(men_men_n85_), .Y(men_men_n949_));
  AN2        u0921(.A(c), .B(b), .Y(men_men_n950_));
  NA3        u0922(.A(men_men_n233_), .B(men_men_n950_), .C(m), .Y(men_men_n951_));
  NO2        u0923(.A(men_men_n951_), .B(men_men_n949_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n248_), .B(men_men_n950_), .Y(men_men_n953_));
  NO4        u0925(.A(men_men_n953_), .B(e), .C(men_men_n889_), .D(a), .Y(men_men_n954_));
  NAi32      u0926(.An(d), .Bn(c), .C(e), .Y(men_men_n955_));
  NO3        u0927(.A(men_men_n955_), .B(men_men_n556_), .C(men_men_n285_), .Y(men_men_n956_));
  NA2        u0928(.A(men_men_n621_), .B(men_men_n213_), .Y(men_men_n957_));
  NA2        u0929(.A(men_men_n385_), .B(men_men_n202_), .Y(men_men_n958_));
  AN2        u0930(.A(d), .B(c), .Y(men_men_n959_));
  NA2        u0931(.A(men_men_n959_), .B(men_men_n112_), .Y(men_men_n960_));
  NO3        u0932(.A(men_men_n960_), .B(men_men_n958_), .C(men_men_n166_), .Y(men_men_n961_));
  NA2        u0933(.A(men_men_n467_), .B(c), .Y(men_men_n962_));
  NO4        u0934(.A(men_men_n1371_), .B(men_men_n552_), .C(men_men_n962_), .D(men_men_n285_), .Y(men_men_n963_));
  AO210      u0935(.A0(men_men_n961_), .A1(men_men_n957_), .B0(men_men_n963_), .Y(men_men_n964_));
  OR4        u0936(.A(men_men_n964_), .B(men_men_n956_), .C(men_men_n954_), .D(men_men_n952_), .Y(men_men_n965_));
  NAi32      u0937(.An(f), .Bn(e), .C(c), .Y(men_men_n966_));
  NO2        u0938(.A(men_men_n966_), .B(men_men_n140_), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n967_), .B(g), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n166_), .B(men_men_n968_), .Y(men_men_n969_));
  NO2        u0941(.A(men_men_n962_), .B(men_men_n285_), .Y(men_men_n970_));
  NA2        u0942(.A(men_men_n591_), .B(i), .Y(men_men_n971_));
  NOi21      u0943(.An(men_men_n970_), .B(men_men_n971_), .Y(men_men_n972_));
  NOi41      u0944(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n973_));
  NO2        u0945(.A(men_men_n1375_), .B(men_men_n968_), .Y(men_men_n974_));
  OR3        u0946(.A(e), .B(d), .C(c), .Y(men_men_n975_));
  NA3        u0947(.A(k), .B(j), .C(i), .Y(men_men_n976_));
  NO3        u0948(.A(men_men_n976_), .B(men_men_n285_), .C(men_men_n89_), .Y(men_men_n977_));
  NOi21      u0949(.An(men_men_n977_), .B(men_men_n975_), .Y(men_men_n978_));
  OR4        u0950(.A(men_men_n978_), .B(men_men_n974_), .C(men_men_n972_), .D(men_men_n969_), .Y(men_men_n979_));
  NA3        u0951(.A(men_men_n439_), .B(men_men_n311_), .C(men_men_n56_), .Y(men_men_n980_));
  NO2        u0952(.A(men_men_n980_), .B(men_men_n971_), .Y(men_men_n981_));
  NO3        u0953(.A(men_men_n980_), .B(men_men_n552_), .C(men_men_n45_), .Y(men_men_n982_));
  NO2        u0954(.A(f), .B(c), .Y(men_men_n983_));
  NOi21      u0955(.An(men_men_n983_), .B(men_men_n413_), .Y(men_men_n984_));
  NA2        u0956(.A(men_men_n984_), .B(men_men_n57_), .Y(men_men_n985_));
  NO3        u0957(.A(i), .B(g), .C(l), .Y(men_men_n986_));
  NOi21      u0958(.An(men_men_n986_), .B(men_men_n985_), .Y(men_men_n987_));
  OR3        u0959(.A(men_men_n987_), .B(men_men_n982_), .C(men_men_n981_), .Y(men_men_n988_));
  OR3        u0960(.A(men_men_n988_), .B(men_men_n979_), .C(men_men_n965_), .Y(men02));
  OR3        u0961(.A(n), .B(m), .C(i), .Y(men_men_n990_));
  NO4        u0962(.A(men_men_n990_), .B(h), .C(l), .D(men_men_n975_), .Y(men_men_n991_));
  NOi31      u0963(.An(e), .B(d), .C(c), .Y(men_men_n992_));
  AOI210     u0964(.A0(men_men_n977_), .A1(men_men_n992_), .B0(men_men_n956_), .Y(men_men_n993_));
  AN3        u0965(.A(g), .B(f), .C(c), .Y(men_men_n994_));
  NA3        u0966(.A(men_men_n994_), .B(men_men_n439_), .C(h), .Y(men_men_n995_));
  OR2        u0967(.A(men_men_n976_), .B(men_men_n995_), .Y(men_men_n996_));
  NO3        u0968(.A(men_men_n980_), .B(men_men_n1371_), .C(men_men_n552_), .Y(men_men_n997_));
  NO2        u0969(.A(men_men_n997_), .B(men_men_n969_), .Y(men_men_n998_));
  NO3        u0970(.A(men_men_n135_), .B(men_men_n264_), .C(men_men_n203_), .Y(men_men_n999_));
  INV        u0971(.A(men_men_n972_), .Y(men_men_n1000_));
  NA3        u0972(.A(c), .B(b), .C(a), .Y(men_men_n1001_));
  NO3        u0973(.A(men_men_n1001_), .B(men_men_n831_), .C(men_men_n202_), .Y(men_men_n1002_));
  INV        u0974(.A(men_men_n981_), .Y(men_men_n1003_));
  AN4        u0975(.A(men_men_n1003_), .B(men_men_n1000_), .C(men_men_n998_), .D(men_men_n996_), .Y(men_men_n1004_));
  NO2        u0976(.A(men_men_n960_), .B(men_men_n958_), .Y(men_men_n1005_));
  INV        u0977(.A(men_men_n1375_), .Y(men_men_n1006_));
  AOI210     u0978(.A0(men_men_n1006_), .A1(men_men_n1005_), .B0(men_men_n952_), .Y(men_men_n1007_));
  NAi41      u0979(.An(men_men_n991_), .B(men_men_n1007_), .C(men_men_n1004_), .D(men_men_n993_), .Y(men03));
  NO2        u0980(.A(men_men_n496_), .B(men_men_n562_), .Y(men_men_n1009_));
  NA4        u0981(.A(men_men_n86_), .B(men_men_n85_), .C(g), .D(men_men_n202_), .Y(men_men_n1010_));
  NA4        u0982(.A(men_men_n540_), .B(m), .C(men_men_n109_), .D(men_men_n202_), .Y(men_men_n1011_));
  NA3        u0983(.A(men_men_n1011_), .B(men_men_n345_), .C(men_men_n1010_), .Y(men_men_n1012_));
  NO3        u0984(.A(men_men_n1012_), .B(men_men_n1009_), .C(men_men_n920_), .Y(men_men_n1013_));
  NOi41      u0985(.An(men_men_n747_), .B(men_men_n788_), .C(men_men_n780_), .D(men_men_n664_), .Y(men_men_n1014_));
  OAI220     u0986(.A0(men_men_n1014_), .A1(men_men_n641_), .B0(men_men_n1013_), .B1(men_men_n553_), .Y(men_men_n1015_));
  NA4        u0987(.A(i), .B(men_men_n992_), .C(men_men_n320_), .D(men_men_n311_), .Y(men_men_n1016_));
  OAI210     u0988(.A0(men_men_n756_), .A1(men_men_n394_), .B0(men_men_n1016_), .Y(men_men_n1017_));
  NOi31      u0989(.An(m), .B(n), .C(f), .Y(men_men_n1018_));
  NA2        u0990(.A(men_men_n1018_), .B(men_men_n51_), .Y(men_men_n1019_));
  AN2        u0991(.A(e), .B(c), .Y(men_men_n1020_));
  NA2        u0992(.A(men_men_n1020_), .B(a), .Y(men_men_n1021_));
  OAI220     u0993(.A0(men_men_n1021_), .A1(men_men_n1019_), .B0(men_men_n816_), .B1(men_men_n399_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n476_), .B(l), .Y(men_men_n1023_));
  NOi31      u0995(.An(men_men_n796_), .B(men_men_n951_), .C(men_men_n1023_), .Y(men_men_n1024_));
  NO4        u0996(.A(men_men_n1024_), .B(men_men_n1022_), .C(men_men_n1017_), .D(men_men_n919_), .Y(men_men_n1025_));
  NO2        u0997(.A(men_men_n264_), .B(a), .Y(men_men_n1026_));
  INV        u0998(.A(men_men_n956_), .Y(men_men_n1027_));
  NO2        u0999(.A(men_men_n85_), .B(g), .Y(men_men_n1028_));
  AOI210     u1000(.A0(men_men_n1028_), .A1(i), .B0(men_men_n986_), .Y(men_men_n1029_));
  OR2        u1001(.A(men_men_n1029_), .B(men_men_n985_), .Y(men_men_n1030_));
  NA3        u1002(.A(men_men_n1030_), .B(men_men_n1027_), .C(men_men_n1025_), .Y(men_men_n1031_));
  NO4        u1003(.A(men_men_n1031_), .B(men_men_n1015_), .C(men_men_n758_), .D(men_men_n532_), .Y(men_men_n1032_));
  NA2        u1004(.A(c), .B(b), .Y(men_men_n1033_));
  NO2        u1005(.A(men_men_n650_), .B(men_men_n1033_), .Y(men_men_n1034_));
  OAI210     u1006(.A0(men_men_n794_), .A1(men_men_n771_), .B0(men_men_n388_), .Y(men_men_n1035_));
  OAI210     u1007(.A0(men_men_n1035_), .A1(men_men_n795_), .B0(men_men_n1034_), .Y(men_men_n1036_));
  NAi21      u1008(.An(men_men_n390_), .B(men_men_n1034_), .Y(men_men_n1037_));
  NA3        u1009(.A(men_men_n400_), .B(men_men_n525_), .C(f), .Y(men_men_n1038_));
  NA2        u1010(.A(men_men_n39_), .B(men_men_n1026_), .Y(men_men_n1039_));
  NA3        u1011(.A(men_men_n1039_), .B(men_men_n1038_), .C(men_men_n1037_), .Y(men_men_n1040_));
  NAi21      u1012(.An(f), .B(d), .Y(men_men_n1041_));
  NO2        u1013(.A(men_men_n1041_), .B(men_men_n1001_), .Y(men_men_n1042_));
  AOI210     u1014(.A0(men_men_n1042_), .A1(men_men_n110_), .B0(men_men_n1040_), .Y(men_men_n1043_));
  NA2        u1015(.A(men_men_n442_), .B(men_men_n441_), .Y(men_men_n1044_));
  NO2        u1016(.A(men_men_n172_), .B(men_men_n222_), .Y(men_men_n1045_));
  NA2        u1017(.A(men_men_n1045_), .B(m), .Y(men_men_n1046_));
  NA3        u1018(.A(men_men_n842_), .B(men_men_n1023_), .C(men_men_n445_), .Y(men_men_n1047_));
  OAI210     u1019(.A0(men_men_n1047_), .A1(men_men_n289_), .B0(men_men_n443_), .Y(men_men_n1048_));
  AOI210     u1020(.A0(men_men_n1048_), .A1(men_men_n1044_), .B0(men_men_n1046_), .Y(men_men_n1049_));
  NA2        u1021(.A(men_men_n527_), .B(men_men_n384_), .Y(men_men_n1050_));
  NO2        u1022(.A(men_men_n348_), .B(men_men_n347_), .Y(men_men_n1051_));
  NO2        u1023(.A(men_men_n402_), .B(men_men_n880_), .Y(men_men_n1052_));
  NAi31      u1024(.An(men_men_n1051_), .B(men_men_n1052_), .C(men_men_n1050_), .Y(men_men_n1053_));
  NO2        u1025(.A(men_men_n1053_), .B(men_men_n1049_), .Y(men_men_n1054_));
  NA4        u1026(.A(men_men_n1054_), .B(men_men_n1043_), .C(men_men_n1036_), .D(men_men_n1032_), .Y(men00));
  AOI210     u1027(.A0(men_men_n279_), .A1(men_men_n203_), .B0(men_men_n259_), .Y(men_men_n1056_));
  NO2        u1028(.A(men_men_n1056_), .B(men_men_n543_), .Y(men_men_n1057_));
  AOI210     u1029(.A0(men_men_n828_), .A1(men_men_n864_), .B0(men_men_n1017_), .Y(men_men_n1058_));
  NO3        u1030(.A(men_men_n997_), .B(men_men_n880_), .C(men_men_n661_), .Y(men_men_n1059_));
  NA3        u1031(.A(men_men_n1059_), .B(men_men_n1058_), .C(men_men_n921_), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n478_), .B(f), .Y(men_men_n1061_));
  NO2        u1033(.A(men_men_n928_), .B(men_men_n40_), .Y(men_men_n1062_));
  NA3        u1034(.A(men_men_n1062_), .B(men_men_n240_), .C(n), .Y(men_men_n1063_));
  AOI210     u1035(.A0(men_men_n1063_), .A1(men_men_n1061_), .B0(men_men_n960_), .Y(men_men_n1064_));
  NO4        u1036(.A(men_men_n1064_), .B(men_men_n1060_), .C(men_men_n1057_), .D(men_men_n979_), .Y(men_men_n1065_));
  NA3        u1037(.A(n), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1066_));
  NA3        u1038(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1067_));
  NOi31      u1039(.An(n), .B(m), .C(i), .Y(men_men_n1068_));
  NA3        u1040(.A(men_men_n1068_), .B(men_men_n609_), .C(men_men_n51_), .Y(men_men_n1069_));
  OAI210     u1041(.A0(men_men_n1067_), .A1(men_men_n1066_), .B0(men_men_n1069_), .Y(men_men_n1070_));
  INV        u1042(.A(men_men_n542_), .Y(men_men_n1071_));
  NO4        u1043(.A(men_men_n1071_), .B(men_men_n1070_), .C(men_men_n1051_), .D(men_men_n843_), .Y(men_men_n1072_));
  NA3        u1044(.A(men_men_n360_), .B(men_men_n210_), .C(g), .Y(men_men_n1073_));
  OA220      u1045(.A0(men_men_n1073_), .A1(men_men_n1067_), .B0(men_men_n361_), .B1(men_men_n129_), .Y(men_men_n1074_));
  NO2        u1046(.A(h), .B(g), .Y(men_men_n1075_));
  NA4        u1047(.A(men_men_n469_), .B(men_men_n439_), .C(men_men_n1075_), .D(men_men_n950_), .Y(men_men_n1076_));
  OAI220     u1048(.A0(men_men_n496_), .A1(men_men_n562_), .B0(men_men_n90_), .B1(men_men_n89_), .Y(men_men_n1077_));
  AOI220     u1049(.A0(men_men_n1077_), .A1(men_men_n505_), .B0(men_men_n868_), .B1(men_men_n541_), .Y(men_men_n1078_));
  AOI220     u1050(.A0(men_men_n295_), .A1(men_men_n230_), .B0(men_men_n167_), .B1(men_men_n142_), .Y(men_men_n1079_));
  NA4        u1051(.A(men_men_n1079_), .B(men_men_n1078_), .C(men_men_n1076_), .D(men_men_n1074_), .Y(men_men_n1080_));
  NO2        u1052(.A(men_men_n1080_), .B(men_men_n250_), .Y(men_men_n1081_));
  INV        u1053(.A(men_men_n300_), .Y(men_men_n1082_));
  AOI210     u1054(.A0(men_men_n230_), .A1(men_men_n323_), .B0(men_men_n544_), .Y(men_men_n1083_));
  NA3        u1055(.A(men_men_n1083_), .B(men_men_n1082_), .C(men_men_n148_), .Y(men_men_n1084_));
  NO2        u1056(.A(men_men_n224_), .B(men_men_n171_), .Y(men_men_n1085_));
  NA2        u1057(.A(men_men_n1085_), .B(men_men_n400_), .Y(men_men_n1086_));
  NA3        u1058(.A(men_men_n169_), .B(men_men_n109_), .C(g), .Y(men_men_n1087_));
  NOi31      u1059(.An(men_men_n804_), .B(h), .C(men_men_n1087_), .Y(men_men_n1088_));
  NAi21      u1060(.An(men_men_n1088_), .B(men_men_n1086_), .Y(men_men_n1089_));
  NO2        u1061(.A(men_men_n258_), .B(men_men_n71_), .Y(men_men_n1090_));
  NO3        u1062(.A(men_men_n399_), .B(men_men_n767_), .C(n), .Y(men_men_n1091_));
  AOI210     u1063(.A0(men_men_n1091_), .A1(men_men_n1090_), .B0(men_men_n991_), .Y(men_men_n1092_));
  NAi31      u1064(.An(men_men_n963_), .B(men_men_n1092_), .C(men_men_n70_), .Y(men_men_n1093_));
  NO4        u1065(.A(men_men_n1093_), .B(men_men_n1089_), .C(men_men_n1084_), .D(men_men_n487_), .Y(men_men_n1094_));
  AN3        u1066(.A(men_men_n1094_), .B(men_men_n1081_), .C(men_men_n1072_), .Y(men_men_n1095_));
  NA2        u1067(.A(men_men_n505_), .B(men_men_n100_), .Y(men_men_n1096_));
  NA3        u1068(.A(men_men_n1018_), .B(men_men_n570_), .C(men_men_n438_), .Y(men_men_n1097_));
  NA3        u1069(.A(men_men_n1097_), .B(men_men_n1096_), .C(men_men_n227_), .Y(men_men_n1098_));
  NA2        u1070(.A(men_men_n1012_), .B(men_men_n505_), .Y(men_men_n1099_));
  NA4        u1071(.A(men_men_n609_), .B(men_men_n194_), .C(men_men_n210_), .D(men_men_n156_), .Y(men_men_n1100_));
  NA3        u1072(.A(men_men_n1100_), .B(men_men_n1099_), .C(men_men_n276_), .Y(men_men_n1101_));
  OAI210     u1073(.A0(men_men_n437_), .A1(men_men_n116_), .B0(men_men_n797_), .Y(men_men_n1102_));
  NA2        u1074(.A(men_men_n1102_), .B(men_men_n1047_), .Y(men_men_n1103_));
  OR4        u1075(.A(men_men_n960_), .B(men_men_n256_), .C(men_men_n211_), .D(e), .Y(men_men_n1104_));
  NO2        u1076(.A(men_men_n206_), .B(men_men_n203_), .Y(men_men_n1105_));
  NA2        u1077(.A(n), .B(e), .Y(men_men_n1106_));
  NO2        u1078(.A(men_men_n1106_), .B(men_men_n140_), .Y(men_men_n1107_));
  AOI220     u1079(.A0(men_men_n1107_), .A1(men_men_n1374_), .B0(men_men_n784_), .B1(men_men_n1105_), .Y(men_men_n1108_));
  OAI210     u1080(.A0(men_men_n332_), .A1(men_men_n290_), .B0(men_men_n418_), .Y(men_men_n1109_));
  NA4        u1081(.A(men_men_n1109_), .B(men_men_n1108_), .C(men_men_n1104_), .D(men_men_n1103_), .Y(men_men_n1110_));
  NO2        u1082(.A(men_men_n64_), .B(h), .Y(men_men_n1111_));
  NO3        u1083(.A(men_men_n960_), .B(men_men_n958_), .C(men_men_n678_), .Y(men_men_n1112_));
  OAI210     u1084(.A0(men_men_n999_), .A1(men_men_n1112_), .B0(men_men_n1111_), .Y(men_men_n1113_));
  NA2        u1085(.A(men_men_n1113_), .B(men_men_n799_), .Y(men_men_n1114_));
  NO4        u1086(.A(men_men_n1114_), .B(men_men_n1110_), .C(men_men_n1101_), .D(men_men_n1098_), .Y(men_men_n1115_));
  NA2        u1087(.A(men_men_n772_), .B(men_men_n705_), .Y(men_men_n1116_));
  NA4        u1088(.A(men_men_n1116_), .B(men_men_n1115_), .C(men_men_n1095_), .D(men_men_n1065_), .Y(men01));
  AN2        u1089(.A(men_men_n939_), .B(men_men_n938_), .Y(men_men_n1118_));
  NO3        u1090(.A(men_men_n744_), .B(men_men_n736_), .C(men_men_n451_), .Y(men_men_n1119_));
  NA2        u1091(.A(men_men_n369_), .B(i), .Y(men_men_n1120_));
  NA3        u1092(.A(men_men_n1120_), .B(men_men_n1119_), .C(men_men_n1118_), .Y(men_men_n1121_));
  NA2        u1093(.A(men_men_n554_), .B(men_men_n88_), .Y(men_men_n1122_));
  NA2        u1094(.A(men_men_n883_), .B(c), .Y(men_men_n1123_));
  NA2        u1095(.A(men_men_n1123_), .B(men_men_n1122_), .Y(men_men_n1124_));
  NA2        u1096(.A(men_men_n45_), .B(f), .Y(men_men_n1125_));
  NA2        u1097(.A(men_men_n656_), .B(men_men_n95_), .Y(men_men_n1126_));
  NO2        u1098(.A(men_men_n1126_), .B(men_men_n1125_), .Y(men_men_n1127_));
  OAI210     u1099(.A0(men_men_n726_), .A1(men_men_n565_), .B0(men_men_n1100_), .Y(men_men_n1128_));
  AOI210     u1100(.A0(men_men_n1127_), .A1(men_men_n598_), .B0(men_men_n1128_), .Y(men_men_n1129_));
  OA210      u1101(.A0(men_men_n617_), .A1(men_men_n345_), .B0(men_men_n551_), .Y(men_men_n1130_));
  NAi41      u1102(.An(men_men_n155_), .B(men_men_n1130_), .C(men_men_n1129_), .D(men_men_n827_), .Y(men_men_n1131_));
  NO3        u1103(.A(men_men_n727_), .B(men_men_n627_), .C(men_men_n481_), .Y(men_men_n1132_));
  NA4        u1104(.A(men_men_n656_), .B(men_men_n95_), .C(men_men_n45_), .D(men_men_n202_), .Y(men_men_n1133_));
  OA220      u1105(.A0(men_men_n1133_), .A1(men_men_n69_), .B0(men_men_n183_), .B1(men_men_n181_), .Y(men_men_n1134_));
  NA2        u1106(.A(men_men_n1134_), .B(men_men_n1132_), .Y(men_men_n1135_));
  NO4        u1107(.A(men_men_n1135_), .B(men_men_n1131_), .C(men_men_n1124_), .D(men_men_n1121_), .Y(men_men_n1136_));
  NA2        u1108(.A(men_men_n1073_), .B(men_men_n195_), .Y(men_men_n1137_));
  NA2        u1109(.A(men_men_n1137_), .B(men_men_n500_), .Y(men_men_n1138_));
  NA2        u1110(.A(men_men_n508_), .B(men_men_n371_), .Y(men_men_n1139_));
  NA2        u1111(.A(men_men_n529_), .B(men_men_n1139_), .Y(men_men_n1140_));
  AOI210     u1112(.A0(men_men_n192_), .A1(men_men_n87_), .B0(men_men_n202_), .Y(men_men_n1141_));
  OAI210     u1113(.A0(men_men_n748_), .A1(men_men_n400_), .B0(men_men_n1141_), .Y(men_men_n1142_));
  NA2        u1114(.A(men_men_n191_), .B(men_men_n34_), .Y(men_men_n1143_));
  OR2        u1115(.A(men_men_n1143_), .B(men_men_n310_), .Y(men_men_n1144_));
  NA4        u1116(.A(men_men_n1144_), .B(men_men_n1142_), .C(men_men_n1140_), .D(men_men_n1138_), .Y(men_men_n1145_));
  AOI210     u1117(.A0(men_men_n560_), .A1(men_men_n114_), .B0(men_men_n563_), .Y(men_men_n1146_));
  NA2        u1118(.A(men_men_n557_), .B(men_men_n1146_), .Y(men_men_n1147_));
  OAI210     u1119(.A0(men_men_n1127_), .A1(men_men_n305_), .B0(men_men_n628_), .Y(men_men_n1148_));
  NA2        u1120(.A(men_men_n1148_), .B(men_men_n729_), .Y(men_men_n1149_));
  NO3        u1121(.A(men_men_n1149_), .B(men_men_n1147_), .C(men_men_n1145_), .Y(men_men_n1150_));
  OR3        u1122(.A(men_men_n1126_), .B(men_men_n567_), .C(men_men_n1125_), .Y(men_men_n1151_));
  NO2        u1123(.A(men_men_n1133_), .B(men_men_n902_), .Y(men_men_n1152_));
  NO2        u1124(.A(men_men_n1152_), .B(men_men_n1070_), .Y(men_men_n1153_));
  NA3        u1125(.A(men_men_n1153_), .B(men_men_n1151_), .C(men_men_n704_), .Y(men_men_n1154_));
  NO2        u1126(.A(men_men_n889_), .B(men_men_n218_), .Y(men_men_n1155_));
  INV        u1127(.A(men_men_n890_), .Y(men_men_n1156_));
  OAI210     u1128(.A0(men_men_n1156_), .A1(men_men_n1155_), .B0(men_men_n318_), .Y(men_men_n1157_));
  NA2        u1129(.A(men_men_n536_), .B(m), .Y(men_men_n1158_));
  NA2        u1130(.A(men_men_n1158_), .B(men_men_n622_), .Y(men_men_n1159_));
  OR2        u1131(.A(men_men_n1073_), .B(men_men_n1067_), .Y(men_men_n1160_));
  NO2        u1132(.A(men_men_n345_), .B(men_men_n69_), .Y(men_men_n1161_));
  INV        u1133(.A(men_men_n1161_), .Y(men_men_n1162_));
  NA3        u1134(.A(men_men_n1162_), .B(men_men_n1160_), .C(men_men_n363_), .Y(men_men_n1163_));
  NOi41      u1135(.An(men_men_n1157_), .B(men_men_n1163_), .C(men_men_n1159_), .D(men_men_n1154_), .Y(men_men_n1164_));
  AN2        u1136(.A(h), .B(men_men_n654_), .Y(men_men_n1165_));
  NA2        u1137(.A(men_men_n1165_), .B(men_men_n318_), .Y(men_men_n1166_));
  NO2        u1138(.A(men_men_n166_), .B(men_men_n85_), .Y(men_men_n1167_));
  INV        u1139(.A(men_men_n1166_), .Y(men_men_n1168_));
  NO2        u1140(.A(men_men_n1168_), .B(men_men_n602_), .Y(men_men_n1169_));
  NA4        u1141(.A(men_men_n1169_), .B(men_men_n1164_), .C(men_men_n1150_), .D(men_men_n1136_), .Y(men06));
  NA2        u1142(.A(men_men_n1167_), .B(men_men_n359_), .Y(men_men_n1171_));
  NA3        u1143(.A(men_men_n816_), .B(men_men_n1171_), .C(men_men_n1157_), .Y(men_men_n1172_));
  NO3        u1144(.A(men_men_n1172_), .B(men_men_n1159_), .C(men_men_n239_), .Y(men_men_n1173_));
  NO2        u1145(.A(men_men_n280_), .B(men_men_n45_), .Y(men_men_n1174_));
  INV        u1146(.A(men_men_n1165_), .Y(men_men_n1175_));
  AOI210     u1147(.A0(men_men_n1175_), .A1(men_men_n1370_), .B0(men_men_n315_), .Y(men_men_n1176_));
  OAI210     u1148(.A0(men_men_n87_), .A1(men_men_n40_), .B0(men_men_n626_), .Y(men_men_n1177_));
  NA2        u1149(.A(men_men_n1177_), .B(men_men_n336_), .Y(men_men_n1178_));
  NO2        u1150(.A(men_men_n484_), .B(men_men_n162_), .Y(men_men_n1179_));
  NO2        u1151(.A(men_men_n571_), .B(men_men_n1019_), .Y(men_men_n1180_));
  NO2        u1152(.A(men_men_n1180_), .B(men_men_n1179_), .Y(men_men_n1181_));
  NO2        u1153(.A(men_men_n344_), .B(men_men_n130_), .Y(men_men_n1182_));
  AOI210     u1154(.A0(men_men_n1182_), .A1(men_men_n554_), .B0(men_men_n563_), .Y(men_men_n1183_));
  NA3        u1155(.A(men_men_n1183_), .B(men_men_n1181_), .C(men_men_n1178_), .Y(men_men_n1184_));
  NO2        u1156(.A(men_men_n696_), .B(men_men_n343_), .Y(men_men_n1185_));
  AN2        u1157(.A(men_men_n876_), .B(men_men_n606_), .Y(men_men_n1186_));
  NO4        u1158(.A(men_men_n1186_), .B(men_men_n1185_), .C(men_men_n1184_), .D(men_men_n1176_), .Y(men_men_n1187_));
  NO2        u1159(.A(men_men_n743_), .B(men_men_n260_), .Y(men_men_n1188_));
  NO2        u1160(.A(men_men_n1372_), .B(men_men_n47_), .Y(men_men_n1189_));
  NO2        u1161(.A(men_men_n260_), .B(c), .Y(men_men_n1190_));
  AOI220     u1162(.A0(men_men_n1190_), .A1(men_men_n1189_), .B0(men_men_n1188_), .B1(men_men_n251_), .Y(men_men_n1191_));
  NO3        u1163(.A(g), .B(men_men_n101_), .C(men_men_n264_), .Y(men_men_n1192_));
  OAI210     u1164(.A0(l), .A1(i), .B0(k), .Y(men_men_n1193_));
  NO3        u1165(.A(men_men_n1193_), .B(men_men_n562_), .C(j), .Y(men_men_n1194_));
  NOi21      u1166(.An(men_men_n1194_), .B(men_men_n69_), .Y(men_men_n1195_));
  NO3        u1167(.A(men_men_n1195_), .B(men_men_n1192_), .C(men_men_n1022_), .Y(men_men_n1196_));
  NAi31      u1168(.An(men_men_n696_), .B(men_men_n82_), .C(men_men_n191_), .Y(men_men_n1197_));
  NA3        u1169(.A(men_men_n1197_), .B(men_men_n1196_), .C(men_men_n1191_), .Y(men_men_n1198_));
  OR2        u1170(.A(men_men_n726_), .B(men_men_n511_), .Y(men_men_n1199_));
  NA2        u1171(.A(men_men_n1194_), .B(men_men_n733_), .Y(men_men_n1200_));
  NA2        u1172(.A(men_men_n1200_), .B(men_men_n1199_), .Y(men_men_n1201_));
  NA2        u1173(.A(men_men_n1182_), .B(men_men_n223_), .Y(men_men_n1202_));
  AN2        u1174(.A(men_men_n850_), .B(men_men_n849_), .Y(men_men_n1203_));
  NO4        u1175(.A(men_men_n1203_), .B(men_men_n809_), .C(men_men_n471_), .D(men_men_n454_), .Y(men_men_n1204_));
  NA2        u1176(.A(men_men_n1204_), .B(men_men_n1202_), .Y(men_men_n1205_));
  NO3        u1177(.A(men_men_n1205_), .B(men_men_n1201_), .C(men_men_n1198_), .Y(men_men_n1206_));
  NA4        u1178(.A(men_men_n1206_), .B(men_men_n1187_), .C(men_men_n1173_), .D(men_men_n1169_), .Y(men07));
  NOi21      u1179(.An(j), .B(k), .Y(men_men_n1208_));
  NAi32      u1180(.An(m), .Bn(b), .C(n), .Y(men_men_n1209_));
  NO3        u1181(.A(men_men_n1209_), .B(g), .C(f), .Y(men_men_n1210_));
  OAI210     u1182(.A0(men_men_n299_), .A1(men_men_n455_), .B0(men_men_n1210_), .Y(men_men_n1211_));
  NAi21      u1183(.An(f), .B(c), .Y(men_men_n1212_));
  NOi31      u1184(.An(n), .B(m), .C(b), .Y(men_men_n1213_));
  INV        u1185(.A(men_men_n1211_), .Y(men_men_n1214_));
  NOi41      u1186(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1215_));
  NA3        u1187(.A(men_men_n1215_), .B(men_men_n801_), .C(men_men_n385_), .Y(men_men_n1216_));
  INV        u1188(.A(men_men_n1216_), .Y(men_men_n1217_));
  NA2        u1189(.A(men_men_n999_), .B(men_men_n210_), .Y(men_men_n1218_));
  NO2        u1190(.A(men_men_n1218_), .B(men_men_n59_), .Y(men_men_n1219_));
  NO2        u1191(.A(k), .B(i), .Y(men_men_n1220_));
  NO2        u1192(.A(men_men_n976_), .B(men_men_n285_), .Y(men_men_n1221_));
  NA2        u1193(.A(men_men_n1111_), .B(men_men_n270_), .Y(men_men_n1222_));
  INV        u1194(.A(men_men_n1222_), .Y(men_men_n1223_));
  NO4        u1195(.A(men_men_n1223_), .B(men_men_n1219_), .C(men_men_n1217_), .D(men_men_n1214_), .Y(men_men_n1224_));
  NO3        u1196(.A(e), .B(d), .C(c), .Y(men_men_n1225_));
  OAI210     u1197(.A0(men_men_n127_), .A1(men_men_n203_), .B0(men_men_n568_), .Y(men_men_n1226_));
  NA2        u1198(.A(men_men_n1226_), .B(men_men_n1225_), .Y(men_men_n1227_));
  INV        u1199(.A(men_men_n1227_), .Y(men_men_n1228_));
  OR2        u1200(.A(h), .B(f), .Y(men_men_n1229_));
  NO3        u1201(.A(n), .B(m), .C(i), .Y(men_men_n1230_));
  OAI210     u1202(.A0(men_men_n1020_), .A1(men_men_n151_), .B0(men_men_n1230_), .Y(men_men_n1231_));
  NO2        u1203(.A(i), .B(g), .Y(men_men_n1232_));
  OR3        u1204(.A(men_men_n1232_), .B(men_men_n1209_), .C(men_men_n68_), .Y(men_men_n1233_));
  OAI220     u1205(.A0(men_men_n1233_), .A1(men_men_n455_), .B0(men_men_n1231_), .B1(men_men_n1229_), .Y(men_men_n1234_));
  NA2        u1206(.A(men_men_n645_), .B(men_men_n109_), .Y(men_men_n1235_));
  NA3        u1207(.A(men_men_n1213_), .B(l), .C(men_men_n624_), .Y(men_men_n1236_));
  AOI210     u1208(.A0(men_men_n1236_), .A1(men_men_n1235_), .B0(men_men_n45_), .Y(men_men_n1237_));
  NA2        u1209(.A(men_men_n1230_), .B(men_men_n604_), .Y(men_men_n1238_));
  NO3        u1210(.A(men_men_n413_), .B(d), .C(c), .Y(men_men_n1239_));
  NO3        u1211(.A(men_men_n1237_), .B(men_men_n1234_), .C(men_men_n1228_), .Y(men_men_n1240_));
  NO2        u1212(.A(g), .B(c), .Y(men_men_n1241_));
  NO2        u1213(.A(men_men_n423_), .B(a), .Y(men_men_n1242_));
  NA3        u1214(.A(men_men_n1242_), .B(k), .C(men_men_n110_), .Y(men_men_n1243_));
  NO2        u1215(.A(i), .B(h), .Y(men_men_n1244_));
  NA2        u1216(.A(men_men_n1244_), .B(men_men_n210_), .Y(men_men_n1245_));
  NA2        u1217(.A(men_men_n1041_), .B(h), .Y(men_men_n1246_));
  NA2        u1218(.A(men_men_n131_), .B(men_men_n210_), .Y(men_men_n1247_));
  AOI210     u1219(.A0(men_men_n240_), .A1(men_men_n112_), .B0(men_men_n500_), .Y(men_men_n1248_));
  OAI220     u1220(.A0(men_men_n1248_), .A1(men_men_n1245_), .B0(men_men_n1247_), .B1(men_men_n1246_), .Y(men_men_n1249_));
  NO2        u1221(.A(men_men_n702_), .B(men_men_n177_), .Y(men_men_n1250_));
  NOi31      u1222(.An(m), .B(n), .C(b), .Y(men_men_n1251_));
  NOi31      u1223(.An(f), .B(d), .C(c), .Y(men_men_n1252_));
  NA2        u1224(.A(men_men_n1252_), .B(men_men_n1251_), .Y(men_men_n1253_));
  INV        u1225(.A(men_men_n1253_), .Y(men_men_n1254_));
  NO3        u1226(.A(men_men_n1254_), .B(men_men_n1250_), .C(men_men_n1249_), .Y(men_men_n1255_));
  OAI210     u1227(.A0(men_men_n172_), .A1(men_men_n495_), .B0(men_men_n973_), .Y(men_men_n1256_));
  AN3        u1228(.A(men_men_n1256_), .B(men_men_n1255_), .C(men_men_n1243_), .Y(men_men_n1257_));
  NA2        u1229(.A(men_men_n1213_), .B(men_men_n356_), .Y(men_men_n1258_));
  NO2        u1230(.A(men_men_n1258_), .B(men_men_n957_), .Y(men_men_n1259_));
  NA2        u1231(.A(men_men_n1239_), .B(men_men_n204_), .Y(men_men_n1260_));
  NO2        u1232(.A(men_men_n177_), .B(b), .Y(men_men_n1261_));
  NO2        u1233(.A(i), .B(men_men_n202_), .Y(men_men_n1262_));
  NA4        u1234(.A(men_men_n1045_), .B(men_men_n1262_), .C(men_men_n102_), .D(m), .Y(men_men_n1263_));
  NAi31      u1235(.An(men_men_n1259_), .B(men_men_n1263_), .C(men_men_n1260_), .Y(men_men_n1264_));
  NO4        u1236(.A(men_men_n127_), .B(g), .C(f), .D(e), .Y(men_men_n1265_));
  NA3        u1237(.A(men_men_n1220_), .B(men_men_n271_), .C(h), .Y(men_men_n1266_));
  NA2        u1238(.A(men_men_n182_), .B(men_men_n97_), .Y(men_men_n1267_));
  NA2        u1239(.A(men_men_n30_), .B(h), .Y(men_men_n1268_));
  NO2        u1240(.A(men_men_n1268_), .B(men_men_n990_), .Y(men_men_n1269_));
  NOi41      u1241(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1270_));
  NA2        u1242(.A(men_men_n1270_), .B(men_men_n110_), .Y(men_men_n1271_));
  INV        u1243(.A(men_men_n1271_), .Y(men_men_n1272_));
  OR3        u1244(.A(men_men_n511_), .B(men_men_n510_), .C(men_men_n109_), .Y(men_men_n1273_));
  NA2        u1245(.A(men_men_n1018_), .B(men_men_n382_), .Y(men_men_n1274_));
  OAI220     u1246(.A0(men_men_n1274_), .A1(men_men_n406_), .B0(men_men_n1273_), .B1(men_men_n280_), .Y(men_men_n1275_));
  AO210      u1247(.A0(men_men_n1275_), .A1(men_men_n112_), .B0(men_men_n1272_), .Y(men_men_n1276_));
  NO3        u1248(.A(men_men_n1276_), .B(men_men_n1269_), .C(men_men_n1264_), .Y(men_men_n1277_));
  NA4        u1249(.A(men_men_n1277_), .B(men_men_n1257_), .C(men_men_n1240_), .D(men_men_n1224_), .Y(men_men_n1278_));
  NO2        u1250(.A(men_men_n1033_), .B(men_men_n107_), .Y(men_men_n1279_));
  NA2        u1251(.A(men_men_n356_), .B(men_men_n56_), .Y(men_men_n1280_));
  NO2        u1252(.A(men_men_n1280_), .B(men_men_n1238_), .Y(men_men_n1281_));
  NA2        u1253(.A(men_men_n204_), .B(men_men_n169_), .Y(men_men_n1282_));
  AOI210     u1254(.A0(men_men_n1282_), .A1(men_men_n1087_), .B0(men_men_n1280_), .Y(men_men_n1283_));
  NO2        u1255(.A(men_men_n995_), .B(men_men_n990_), .Y(men_men_n1284_));
  NO3        u1256(.A(men_men_n1284_), .B(men_men_n1283_), .C(men_men_n1281_), .Y(men_men_n1285_));
  NO3        u1257(.A(men_men_n990_), .B(men_men_n548_), .C(g), .Y(men_men_n1286_));
  NOi21      u1258(.An(men_men_n1282_), .B(men_men_n1286_), .Y(men_men_n1287_));
  AOI210     u1259(.A0(men_men_n1287_), .A1(men_men_n1267_), .B0(men_men_n966_), .Y(men_men_n1288_));
  OAI220     u1260(.A0(men_men_n621_), .A1(g), .B0(men_men_n213_), .B1(c), .Y(men_men_n1289_));
  AOI210     u1261(.A0(men_men_n1261_), .A1(men_men_n41_), .B0(men_men_n1289_), .Y(men_men_n1290_));
  NO2        u1262(.A(men_men_n127_), .B(l), .Y(men_men_n1291_));
  NO2        u1263(.A(men_men_n213_), .B(k), .Y(men_men_n1292_));
  OAI210     u1264(.A0(men_men_n1292_), .A1(men_men_n1244_), .B0(men_men_n1291_), .Y(men_men_n1293_));
  OAI220     u1265(.A0(men_men_n1293_), .A1(men_men_n31_), .B0(men_men_n1290_), .B1(men_men_n166_), .Y(men_men_n1294_));
  NO3        u1266(.A(men_men_n1273_), .B(men_men_n439_), .C(men_men_n330_), .Y(men_men_n1295_));
  NO3        u1267(.A(men_men_n1295_), .B(men_men_n1294_), .C(men_men_n1288_), .Y(men_men_n1296_));
  INV        u1268(.A(men_men_n1002_), .Y(men_men_n1297_));
  NO2        u1269(.A(men_men_n990_), .B(h), .Y(men_men_n1298_));
  NA3        u1270(.A(men_men_n1298_), .B(d), .C(men_men_n958_), .Y(men_men_n1299_));
  OAI220     u1271(.A0(men_men_n1299_), .A1(c), .B0(men_men_n1297_), .B1(j), .Y(men_men_n1300_));
  NA3        u1272(.A(men_men_n1279_), .B(men_men_n439_), .C(f), .Y(men_men_n1301_));
  NA2        u1273(.A(men_men_n169_), .B(men_men_n109_), .Y(men_men_n1302_));
  NO2        u1274(.A(men_men_n1208_), .B(men_men_n42_), .Y(men_men_n1303_));
  AOI210     u1275(.A0(men_men_n110_), .A1(men_men_n40_), .B0(men_men_n1303_), .Y(men_men_n1304_));
  NO2        u1276(.A(men_men_n1304_), .B(men_men_n1301_), .Y(men_men_n1305_));
  AOI210     u1277(.A0(men_men_n495_), .A1(h), .B0(men_men_n65_), .Y(men_men_n1306_));
  NA2        u1278(.A(men_men_n1306_), .B(men_men_n1242_), .Y(men_men_n1307_));
  NO2        u1279(.A(j), .B(men_men_n164_), .Y(men_men_n1308_));
  NOi21      u1280(.An(d), .B(f), .Y(men_men_n1309_));
  NO3        u1281(.A(men_men_n1252_), .B(men_men_n1309_), .C(men_men_n40_), .Y(men_men_n1310_));
  NA2        u1282(.A(men_men_n1310_), .B(men_men_n1308_), .Y(men_men_n1311_));
  NA2        u1283(.A(men_men_n1242_), .B(men_men_n1303_), .Y(men_men_n1312_));
  NO2        u1284(.A(men_men_n280_), .B(c), .Y(men_men_n1313_));
  NA2        u1285(.A(men_men_n1313_), .B(men_men_n512_), .Y(men_men_n1314_));
  NA4        u1286(.A(men_men_n1314_), .B(men_men_n1312_), .C(men_men_n1311_), .D(men_men_n1307_), .Y(men_men_n1315_));
  NO3        u1287(.A(men_men_n1315_), .B(men_men_n1305_), .C(men_men_n1300_), .Y(men_men_n1316_));
  NA3        u1288(.A(men_men_n1316_), .B(men_men_n1296_), .C(men_men_n1285_), .Y(men_men_n1317_));
  NO3        u1289(.A(men_men_n994_), .B(men_men_n983_), .C(men_men_n40_), .Y(men_men_n1318_));
  NA2        u1290(.A(men_men_n1318_), .B(men_men_n1221_), .Y(men_men_n1319_));
  OAI210     u1291(.A0(men_men_n1265_), .A1(men_men_n1213_), .B0(men_men_n813_), .Y(men_men_n1320_));
  NO2        u1292(.A(men_men_n955_), .B(men_men_n127_), .Y(men_men_n1321_));
  NA2        u1293(.A(men_men_n1321_), .B(men_men_n583_), .Y(men_men_n1322_));
  NA3        u1294(.A(men_men_n1322_), .B(men_men_n1320_), .C(men_men_n1319_), .Y(men_men_n1323_));
  NA2        u1295(.A(men_men_n1241_), .B(men_men_n1309_), .Y(men_men_n1324_));
  NO2        u1296(.A(men_men_n1324_), .B(m), .Y(men_men_n1325_));
  NA3        u1297(.A(men_men_n999_), .B(men_men_n105_), .C(men_men_n210_), .Y(men_men_n1326_));
  INV        u1298(.A(men_men_n1326_), .Y(men_men_n1327_));
  NO3        u1299(.A(men_men_n1327_), .B(men_men_n1325_), .C(men_men_n1323_), .Y(men_men_n1328_));
  NO2        u1300(.A(men_men_n1212_), .B(e), .Y(men_men_n1329_));
  NO3        u1301(.A(men_men_n1273_), .B(men_men_n330_), .C(a), .Y(men_men_n1330_));
  NA2        u1302(.A(men_men_n510_), .B(g), .Y(men_men_n1331_));
  NA2        u1303(.A(men_men_n1331_), .B(men_men_n1239_), .Y(men_men_n1332_));
  NA2        u1304(.A(men_men_n1028_), .B(a), .Y(men_men_n1333_));
  OAI220     u1305(.A0(men_men_n1333_), .A1(men_men_n65_), .B0(men_men_n1332_), .B1(men_men_n202_), .Y(men_men_n1334_));
  NA2        u1306(.A(men_men_n831_), .B(men_men_n391_), .Y(men_men_n1335_));
  OR2        u1307(.A(men_men_n1335_), .B(men_men_n510_), .Y(men_men_n1336_));
  NO2        u1308(.A(men_men_n1336_), .B(men_men_n164_), .Y(men_men_n1337_));
  NO2        u1309(.A(men_men_n1337_), .B(men_men_n1334_), .Y(men_men_n1338_));
  NA3        u1310(.A(men_men_n1338_), .B(men_men_n1369_), .C(men_men_n1328_), .Y(men_men_n1339_));
  NA3        u1311(.A(men_men_n882_), .B(men_men_n131_), .C(men_men_n46_), .Y(men_men_n1340_));
  OAI210     u1312(.A0(men_men_n548_), .A1(g), .B0(men_men_n175_), .Y(men_men_n1341_));
  NA2        u1313(.A(men_men_n1341_), .B(men_men_n1298_), .Y(men_men_n1342_));
  NO2        u1314(.A(men_men_n68_), .B(c), .Y(men_men_n1343_));
  NO4        u1315(.A(men_men_n1229_), .B(men_men_n176_), .C(men_men_n420_), .D(men_men_n45_), .Y(men_men_n1344_));
  AOI210     u1316(.A0(men_men_n1308_), .A1(men_men_n1343_), .B0(men_men_n1344_), .Y(men_men_n1345_));
  NA2        u1317(.A(men_men_n1345_), .B(men_men_n1342_), .Y(men_men_n1346_));
  INV        u1318(.A(men_men_n1346_), .Y(men_men_n1347_));
  NO2        u1319(.A(men_men_n151_), .B(men_men_n1329_), .Y(men_men_n1348_));
  NO2        u1320(.A(men_men_n1348_), .B(men_men_n1302_), .Y(men_men_n1349_));
  NO2        u1321(.A(men_men_n1340_), .B(men_men_n107_), .Y(men_men_n1350_));
  NO2        u1322(.A(men_men_n1350_), .B(men_men_n1349_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n1301_), .B(men_men_n65_), .Y(men_men_n1352_));
  NO2        u1324(.A(men_men_n1220_), .B(men_men_n114_), .Y(men_men_n1353_));
  NO2        u1325(.A(men_men_n1353_), .B(men_men_n1258_), .Y(men_men_n1354_));
  NO2        u1326(.A(men_men_n1354_), .B(men_men_n1352_), .Y(men_men_n1355_));
  NA3        u1327(.A(men_men_n1355_), .B(men_men_n1351_), .C(men_men_n1347_), .Y(men_men_n1356_));
  OR4        u1328(.A(men_men_n1356_), .B(men_men_n1339_), .C(men_men_n1317_), .D(men_men_n1278_), .Y(men04));
  NOi31      u1329(.An(men_men_n1265_), .B(men_men_n1266_), .C(men_men_n960_), .Y(men_men_n1358_));
  NO3        u1330(.A(men_men_n951_), .B(men_men_n456_), .C(j), .Y(men_men_n1359_));
  OR3        u1331(.A(men_men_n1359_), .B(men_men_n1358_), .C(men_men_n974_), .Y(men_men_n1360_));
  NO2        u1332(.A(men_men_n89_), .B(k), .Y(men_men_n1361_));
  AOI210     u1333(.A0(men_men_n1361_), .A1(men_men_n970_), .B0(men_men_n1088_), .Y(men_men_n1362_));
  NA2        u1334(.A(men_men_n1362_), .B(men_men_n1113_), .Y(men_men_n1363_));
  NO4        u1335(.A(men_men_n1363_), .B(men_men_n1360_), .C(men_men_n982_), .D(men_men_n965_), .Y(men_men_n1364_));
  NA4        u1336(.A(men_men_n1364_), .B(men_men_n1030_), .C(men_men_n1016_), .D(men_men_n1004_), .Y(men05));
  INV        u1337(.A(b), .Y(men_men_n1368_));
  INV        u1338(.A(men_men_n1330_), .Y(men_men_n1369_));
  INV        u1339(.A(men_men_n1174_), .Y(men_men_n1370_));
  INV        u1340(.A(k), .Y(men_men_n1371_));
  INV        u1341(.A(k), .Y(men_men_n1372_));
  INV        u1342(.A(d), .Y(men_men_n1373_));
  INV        u1343(.A(men_men_n246_), .Y(men_men_n1374_));
  INV        u1344(.A(n), .Y(men_men_n1375_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule