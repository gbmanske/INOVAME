//Benchmark atmr_misex3_1774_0.25

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n33_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1606_, men_men_n1607_, men_men_n1608_, men_men_n1610_, men_men_n1611_, men_men_n1612_, men_men_n1613_, men_men_n1614_, men_men_n1615_, men_men_n1616_, men_men_n1617_, men_men_n1621_, men_men_n1622_, men_men_n1623_, men_men_n1624_, men_men_n1625_, men_men_n1626_, men_men_n1627_, men_men_n1628_, men_men_n1629_, men_men_n1630_, men_men_n1631_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  INV        o00(.A(n), .Y(ori_ori_n29_));
  OR2        o01(.A(ori_ori_n33_), .B(ori_ori_n29_), .Y(ori04));
  INV        o02(.A(m), .Y(ori_ori_n33_));
  ZERO       o03(.Y(ori10));
  ZERO       o04(.Y(ori11));
  ZERO       o05(.Y(ori08));
  ZERO       o06(.Y(ori09));
  ZERO       o07(.Y(ori12));
  ZERO       o08(.Y(ori13));
  ZERO       o09(.Y(ori02));
  ZERO       o10(.Y(ori03));
  ZERO       o11(.Y(ori00));
  ZERO       o12(.Y(ori01));
  ZERO       o13(.Y(ori06));
  ZERO       o14(.Y(ori07));
  ZERO       o15(.Y(ori05));
  NO2        m0000(.A(d), .B(c), .Y(mai_mai_n29_));
  AN2        m0001(.A(f), .B(e), .Y(mai_mai_n30_));
  NA3        m0002(.A(mai_mai_n30_), .B(mai_mai_n29_), .C(a), .Y(mai_mai_n31_));
  NOi32      m0003(.An(m), .Bn(l), .C(n), .Y(mai_mai_n32_));
  NOi32      m0004(.An(i), .Bn(g), .C(h), .Y(mai_mai_n33_));
  NA2        m0005(.A(mai_mai_n33_), .B(mai_mai_n32_), .Y(mai_mai_n34_));
  AN2        m0006(.A(m), .B(l), .Y(mai_mai_n35_));
  NOi32      m0007(.An(j), .Bn(g), .C(k), .Y(mai_mai_n36_));
  NA2        m0008(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n37_));
  NO2        m0009(.A(mai_mai_n37_), .B(n), .Y(mai_mai_n38_));
  INV        m0010(.A(h), .Y(mai_mai_n39_));
  NAi21      m0011(.An(j), .B(l), .Y(mai_mai_n40_));
  NAi32      m0012(.An(n), .Bn(g), .C(m), .Y(mai_mai_n41_));
  NO3        m0013(.A(mai_mai_n41_), .B(mai_mai_n40_), .C(mai_mai_n39_), .Y(mai_mai_n42_));
  NAi31      m0014(.An(n), .B(m), .C(l), .Y(mai_mai_n43_));
  INV        m0015(.A(i), .Y(mai_mai_n44_));
  AN2        m0016(.A(h), .B(g), .Y(mai_mai_n45_));
  NO2        m0017(.A(mai_mai_n1368_), .B(mai_mai_n43_), .Y(mai_mai_n46_));
  NAi21      m0018(.An(n), .B(m), .Y(mai_mai_n47_));
  NOi32      m0019(.An(k), .Bn(h), .C(l), .Y(mai_mai_n48_));
  NOi32      m0020(.An(k), .Bn(h), .C(g), .Y(mai_mai_n49_));
  NO2        m0021(.A(mai_mai_n49_), .B(mai_mai_n48_), .Y(mai_mai_n50_));
  NO2        m0022(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n51_));
  AOI210     m0023(.A0(mai_mai_n47_), .A1(mai_mai_n34_), .B0(mai_mai_n31_), .Y(mai_mai_n52_));
  INV        m0024(.A(c), .Y(mai_mai_n53_));
  NA2        m0025(.A(e), .B(b), .Y(mai_mai_n54_));
  NO2        m0026(.A(mai_mai_n54_), .B(mai_mai_n53_), .Y(mai_mai_n55_));
  INV        m0027(.A(d), .Y(mai_mai_n56_));
  NAi21      m0028(.An(i), .B(h), .Y(mai_mai_n57_));
  NAi31      m0029(.An(i), .B(l), .C(j), .Y(mai_mai_n58_));
  NAi41      m0030(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n59_));
  NA2        m0031(.A(g), .B(f), .Y(mai_mai_n60_));
  NO2        m0032(.A(mai_mai_n60_), .B(mai_mai_n59_), .Y(mai_mai_n61_));
  NAi21      m0033(.An(i), .B(j), .Y(mai_mai_n62_));
  NAi32      m0034(.An(n), .Bn(k), .C(m), .Y(mai_mai_n63_));
  NO2        m0035(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n64_));
  NAi31      m0036(.An(l), .B(m), .C(k), .Y(mai_mai_n65_));
  NAi21      m0037(.An(e), .B(h), .Y(mai_mai_n66_));
  NAi41      m0038(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n67_));
  NA2        m0039(.A(mai_mai_n64_), .B(mai_mai_n61_), .Y(mai_mai_n68_));
  INV        m0040(.A(m), .Y(mai_mai_n69_));
  NA2        m0041(.A(k), .B(mai_mai_n69_), .Y(mai_mai_n70_));
  AN4        m0042(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n71_));
  NA2        m0043(.A(h), .B(mai_mai_n71_), .Y(mai_mai_n72_));
  NAi32      m0044(.An(m), .Bn(k), .C(j), .Y(mai_mai_n73_));
  NOi32      m0045(.An(h), .Bn(g), .C(f), .Y(mai_mai_n74_));
  NA2        m0046(.A(mai_mai_n74_), .B(mai_mai_n71_), .Y(mai_mai_n75_));
  OA220      m0047(.A0(mai_mai_n75_), .A1(mai_mai_n73_), .B0(mai_mai_n72_), .B1(mai_mai_n70_), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n68_), .Y(mai_mai_n77_));
  INV        m0049(.A(n), .Y(mai_mai_n78_));
  NOi32      m0050(.An(e), .Bn(b), .C(d), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  INV        m0052(.A(j), .Y(mai_mai_n81_));
  AN3        m0053(.A(m), .B(k), .C(i), .Y(mai_mai_n82_));
  NA3        m0054(.A(mai_mai_n82_), .B(mai_mai_n81_), .C(g), .Y(mai_mai_n83_));
  NO2        m0055(.A(mai_mai_n83_), .B(f), .Y(mai_mai_n84_));
  NAi32      m0056(.An(g), .Bn(f), .C(h), .Y(mai_mai_n85_));
  NAi31      m0057(.An(j), .B(m), .C(l), .Y(mai_mai_n86_));
  NO2        m0058(.A(mai_mai_n86_), .B(mai_mai_n85_), .Y(mai_mai_n87_));
  NA2        m0059(.A(m), .B(l), .Y(mai_mai_n88_));
  NAi31      m0060(.An(k), .B(j), .C(g), .Y(mai_mai_n89_));
  NO3        m0061(.A(mai_mai_n89_), .B(mai_mai_n88_), .C(f), .Y(mai_mai_n90_));
  AN2        m0062(.A(j), .B(g), .Y(mai_mai_n91_));
  NOi21      m0063(.An(g), .B(i), .Y(mai_mai_n92_));
  NOi32      m0064(.An(m), .Bn(j), .C(k), .Y(mai_mai_n93_));
  AOI220     m0065(.A0(mai_mai_n93_), .A1(mai_mai_n92_), .B0(m), .B1(mai_mai_n91_), .Y(mai_mai_n94_));
  NO2        m0066(.A(mai_mai_n94_), .B(f), .Y(mai_mai_n95_));
  NO4        m0067(.A(mai_mai_n95_), .B(mai_mai_n90_), .C(mai_mai_n87_), .D(mai_mai_n84_), .Y(mai_mai_n96_));
  NAi41      m0068(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n97_));
  AN2        m0069(.A(e), .B(b), .Y(mai_mai_n98_));
  NOi31      m0070(.An(c), .B(h), .C(f), .Y(mai_mai_n99_));
  NA2        m0071(.A(mai_mai_n99_), .B(mai_mai_n98_), .Y(mai_mai_n100_));
  NO3        m0072(.A(mai_mai_n100_), .B(mai_mai_n97_), .C(g), .Y(mai_mai_n101_));
  NOi21      m0073(.An(i), .B(h), .Y(mai_mai_n102_));
  NA3        m0074(.A(mai_mai_n102_), .B(g), .C(mai_mai_n35_), .Y(mai_mai_n103_));
  INV        m0075(.A(a), .Y(mai_mai_n104_));
  NA2        m0076(.A(mai_mai_n98_), .B(mai_mai_n104_), .Y(mai_mai_n105_));
  INV        m0077(.A(l), .Y(mai_mai_n106_));
  NOi21      m0078(.An(m), .B(n), .Y(mai_mai_n107_));
  AN2        m0079(.A(k), .B(h), .Y(mai_mai_n108_));
  NO2        m0080(.A(mai_mai_n103_), .B(mai_mai_n80_), .Y(mai_mai_n109_));
  INV        m0081(.A(b), .Y(mai_mai_n110_));
  NA2        m0082(.A(l), .B(j), .Y(mai_mai_n111_));
  AN2        m0083(.A(k), .B(i), .Y(mai_mai_n112_));
  NA2        m0084(.A(g), .B(e), .Y(mai_mai_n113_));
  NOi32      m0085(.An(c), .Bn(a), .C(d), .Y(mai_mai_n114_));
  NA2        m0086(.A(mai_mai_n114_), .B(mai_mai_n107_), .Y(mai_mai_n115_));
  NO4        m0087(.A(mai_mai_n115_), .B(mai_mai_n113_), .C(mai_mai_n111_), .D(mai_mai_n110_), .Y(mai_mai_n116_));
  NO3        m0088(.A(mai_mai_n116_), .B(mai_mai_n109_), .C(mai_mai_n101_), .Y(mai_mai_n117_));
  OAI210     m0089(.A0(mai_mai_n96_), .A1(mai_mai_n80_), .B0(mai_mai_n117_), .Y(mai_mai_n118_));
  NOi31      m0090(.An(k), .B(m), .C(j), .Y(mai_mai_n119_));
  NA3        m0091(.A(mai_mai_n119_), .B(h), .C(mai_mai_n71_), .Y(mai_mai_n120_));
  NOi31      m0092(.An(k), .B(m), .C(i), .Y(mai_mai_n121_));
  NA3        m0093(.A(mai_mai_n121_), .B(mai_mai_n74_), .C(mai_mai_n71_), .Y(mai_mai_n122_));
  NA2        m0094(.A(mai_mai_n122_), .B(mai_mai_n120_), .Y(mai_mai_n123_));
  NOi32      m0095(.An(f), .Bn(b), .C(e), .Y(mai_mai_n124_));
  NAi21      m0096(.An(g), .B(h), .Y(mai_mai_n125_));
  NAi21      m0097(.An(m), .B(n), .Y(mai_mai_n126_));
  NAi21      m0098(.An(j), .B(k), .Y(mai_mai_n127_));
  NO3        m0099(.A(mai_mai_n127_), .B(mai_mai_n126_), .C(mai_mai_n125_), .Y(mai_mai_n128_));
  NAi41      m0100(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n129_));
  NAi31      m0101(.An(j), .B(k), .C(h), .Y(mai_mai_n130_));
  NO3        m0102(.A(mai_mai_n130_), .B(mai_mai_n129_), .C(mai_mai_n126_), .Y(mai_mai_n131_));
  AOI210     m0103(.A0(mai_mai_n128_), .A1(mai_mai_n124_), .B0(mai_mai_n131_), .Y(mai_mai_n132_));
  NO2        m0104(.A(k), .B(j), .Y(mai_mai_n133_));
  INV        m0105(.A(mai_mai_n126_), .Y(mai_mai_n134_));
  AN2        m0106(.A(k), .B(j), .Y(mai_mai_n135_));
  NAi21      m0107(.An(c), .B(b), .Y(mai_mai_n136_));
  NA2        m0108(.A(f), .B(d), .Y(mai_mai_n137_));
  NO3        m0109(.A(mai_mai_n137_), .B(mai_mai_n136_), .C(mai_mai_n125_), .Y(mai_mai_n138_));
  NA2        m0110(.A(h), .B(c), .Y(mai_mai_n139_));
  NAi31      m0111(.An(f), .B(e), .C(b), .Y(mai_mai_n140_));
  NA2        m0112(.A(mai_mai_n138_), .B(mai_mai_n134_), .Y(mai_mai_n141_));
  NA2        m0113(.A(d), .B(b), .Y(mai_mai_n142_));
  NAi21      m0114(.An(e), .B(f), .Y(mai_mai_n143_));
  NO2        m0115(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NA2        m0116(.A(b), .B(a), .Y(mai_mai_n145_));
  NAi21      m0117(.An(e), .B(g), .Y(mai_mai_n146_));
  NAi21      m0118(.An(c), .B(d), .Y(mai_mai_n147_));
  NAi31      m0119(.An(l), .B(k), .C(h), .Y(mai_mai_n148_));
  NO2        m0120(.A(mai_mai_n126_), .B(mai_mai_n148_), .Y(mai_mai_n149_));
  NA2        m0121(.A(mai_mai_n149_), .B(mai_mai_n144_), .Y(mai_mai_n150_));
  NAi41      m0122(.An(mai_mai_n123_), .B(mai_mai_n150_), .C(mai_mai_n141_), .D(mai_mai_n132_), .Y(mai_mai_n151_));
  NAi31      m0123(.An(e), .B(f), .C(b), .Y(mai_mai_n152_));
  INV        m0124(.A(mai_mai_n152_), .Y(mai_mai_n153_));
  NOi21      m0125(.An(h), .B(i), .Y(mai_mai_n154_));
  NOi21      m0126(.An(k), .B(m), .Y(mai_mai_n155_));
  NA3        m0127(.A(mai_mai_n155_), .B(mai_mai_n154_), .C(n), .Y(mai_mai_n156_));
  NOi21      m0128(.An(mai_mai_n153_), .B(mai_mai_n156_), .Y(mai_mai_n157_));
  NO2        m0129(.A(mai_mai_n137_), .B(mai_mai_n136_), .Y(mai_mai_n158_));
  NA2        m0130(.A(mai_mai_n158_), .B(h), .Y(mai_mai_n159_));
  INV        m0131(.A(mai_mai_n47_), .Y(mai_mai_n160_));
  NA2        m0132(.A(mai_mai_n160_), .B(mai_mai_n61_), .Y(mai_mai_n161_));
  NOi32      m0133(.An(n), .Bn(k), .C(m), .Y(mai_mai_n162_));
  NA2        m0134(.A(l), .B(i), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  OAI210     m0136(.A0(mai_mai_n164_), .A1(mai_mai_n159_), .B0(mai_mai_n161_), .Y(mai_mai_n165_));
  NAi31      m0137(.An(d), .B(f), .C(c), .Y(mai_mai_n166_));
  NAi31      m0138(.An(e), .B(f), .C(c), .Y(mai_mai_n167_));
  NA2        m0139(.A(mai_mai_n167_), .B(mai_mai_n166_), .Y(mai_mai_n168_));
  NA2        m0140(.A(j), .B(h), .Y(mai_mai_n169_));
  OR3        m0141(.A(n), .B(m), .C(k), .Y(mai_mai_n170_));
  NO2        m0142(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n171_));
  NAi32      m0143(.An(m), .Bn(k), .C(n), .Y(mai_mai_n172_));
  NO2        m0144(.A(mai_mai_n172_), .B(mai_mai_n169_), .Y(mai_mai_n173_));
  AOI220     m0145(.A0(mai_mai_n173_), .A1(mai_mai_n153_), .B0(mai_mai_n171_), .B1(mai_mai_n168_), .Y(mai_mai_n174_));
  NO2        m0146(.A(n), .B(m), .Y(mai_mai_n175_));
  NA2        m0147(.A(mai_mai_n175_), .B(mai_mai_n48_), .Y(mai_mai_n176_));
  NAi21      m0148(.An(f), .B(e), .Y(mai_mai_n177_));
  NA2        m0149(.A(d), .B(c), .Y(mai_mai_n178_));
  NO2        m0150(.A(mai_mai_n178_), .B(mai_mai_n177_), .Y(mai_mai_n179_));
  NOi21      m0151(.An(mai_mai_n179_), .B(mai_mai_n176_), .Y(mai_mai_n180_));
  NAi31      m0152(.An(m), .B(n), .C(b), .Y(mai_mai_n181_));
  NA2        m0153(.A(k), .B(i), .Y(mai_mai_n182_));
  NAi21      m0154(.An(h), .B(f), .Y(mai_mai_n183_));
  NO2        m0155(.A(mai_mai_n183_), .B(mai_mai_n182_), .Y(mai_mai_n184_));
  NO2        m0156(.A(mai_mai_n181_), .B(mai_mai_n147_), .Y(mai_mai_n185_));
  NA2        m0157(.A(mai_mai_n185_), .B(mai_mai_n184_), .Y(mai_mai_n186_));
  NOi32      m0158(.An(f), .Bn(c), .C(d), .Y(mai_mai_n187_));
  NOi32      m0159(.An(f), .Bn(c), .C(e), .Y(mai_mai_n188_));
  NO2        m0160(.A(mai_mai_n188_), .B(mai_mai_n187_), .Y(mai_mai_n189_));
  NO3        m0161(.A(n), .B(m), .C(j), .Y(mai_mai_n190_));
  NA2        m0162(.A(mai_mai_n190_), .B(mai_mai_n108_), .Y(mai_mai_n191_));
  AO210      m0163(.A0(mai_mai_n191_), .A1(mai_mai_n176_), .B0(mai_mai_n189_), .Y(mai_mai_n192_));
  NAi41      m0164(.An(mai_mai_n180_), .B(mai_mai_n192_), .C(mai_mai_n186_), .D(mai_mai_n174_), .Y(mai_mai_n193_));
  OR4        m0165(.A(mai_mai_n193_), .B(mai_mai_n165_), .C(mai_mai_n157_), .D(mai_mai_n151_), .Y(mai_mai_n194_));
  NO4        m0166(.A(mai_mai_n194_), .B(mai_mai_n118_), .C(mai_mai_n77_), .D(mai_mai_n52_), .Y(mai_mai_n195_));
  NAi31      m0167(.An(n), .B(h), .C(g), .Y(mai_mai_n196_));
  NO2        m0168(.A(mai_mai_n196_), .B(mai_mai_n1358_), .Y(mai_mai_n197_));
  NOi32      m0169(.An(m), .Bn(k), .C(l), .Y(mai_mai_n198_));
  NA3        m0170(.A(mai_mai_n198_), .B(mai_mai_n81_), .C(g), .Y(mai_mai_n199_));
  NO2        m0171(.A(mai_mai_n199_), .B(n), .Y(mai_mai_n200_));
  NOi21      m0172(.An(k), .B(j), .Y(mai_mai_n201_));
  NA4        m0173(.A(mai_mai_n201_), .B(mai_mai_n107_), .C(i), .D(g), .Y(mai_mai_n202_));
  AN2        m0174(.A(i), .B(g), .Y(mai_mai_n203_));
  NA3        m0175(.A(k), .B(mai_mai_n203_), .C(mai_mai_n107_), .Y(mai_mai_n204_));
  NA2        m0176(.A(mai_mai_n204_), .B(mai_mai_n202_), .Y(mai_mai_n205_));
  NAi41      m0177(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n206_));
  INV        m0178(.A(mai_mai_n206_), .Y(mai_mai_n207_));
  INV        m0179(.A(f), .Y(mai_mai_n208_));
  INV        m0180(.A(g), .Y(mai_mai_n209_));
  NOi31      m0181(.An(i), .B(j), .C(h), .Y(mai_mai_n210_));
  NOi21      m0182(.An(l), .B(m), .Y(mai_mai_n211_));
  NA2        m0183(.A(mai_mai_n211_), .B(mai_mai_n210_), .Y(mai_mai_n212_));
  NO3        m0184(.A(mai_mai_n212_), .B(mai_mai_n209_), .C(mai_mai_n208_), .Y(mai_mai_n213_));
  NA2        m0185(.A(mai_mai_n213_), .B(mai_mai_n207_), .Y(mai_mai_n214_));
  INV        m0186(.A(mai_mai_n214_), .Y(mai_mai_n215_));
  NOi21      m0187(.An(n), .B(m), .Y(mai_mai_n216_));
  NOi32      m0188(.An(l), .Bn(i), .C(j), .Y(mai_mai_n217_));
  NA2        m0189(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  OA220      m0190(.A0(mai_mai_n218_), .A1(mai_mai_n100_), .B0(mai_mai_n73_), .B1(mai_mai_n72_), .Y(mai_mai_n219_));
  NAi21      m0191(.An(j), .B(h), .Y(mai_mai_n220_));
  NOi31      m0192(.An(k), .B(n), .C(m), .Y(mai_mai_n221_));
  NOi31      m0193(.An(mai_mai_n221_), .B(mai_mai_n178_), .C(mai_mai_n177_), .Y(mai_mai_n222_));
  INV        m0194(.A(mai_mai_n222_), .Y(mai_mai_n223_));
  NAi31      m0195(.An(f), .B(e), .C(c), .Y(mai_mai_n224_));
  NO4        m0196(.A(mai_mai_n224_), .B(mai_mai_n170_), .C(mai_mai_n169_), .D(mai_mai_n56_), .Y(mai_mai_n225_));
  NA4        m0197(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n226_));
  NAi32      m0198(.An(m), .Bn(i), .C(k), .Y(mai_mai_n227_));
  NO3        m0199(.A(mai_mai_n227_), .B(mai_mai_n85_), .C(mai_mai_n226_), .Y(mai_mai_n228_));
  NA2        m0200(.A(k), .B(h), .Y(mai_mai_n229_));
  NO2        m0201(.A(mai_mai_n228_), .B(mai_mai_n225_), .Y(mai_mai_n230_));
  NAi21      m0202(.An(n), .B(a), .Y(mai_mai_n231_));
  NO2        m0203(.A(mai_mai_n231_), .B(mai_mai_n142_), .Y(mai_mai_n232_));
  NAi41      m0204(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n233_));
  NO2        m0205(.A(mai_mai_n233_), .B(e), .Y(mai_mai_n234_));
  NO3        m0206(.A(mai_mai_n143_), .B(mai_mai_n89_), .C(mai_mai_n88_), .Y(mai_mai_n235_));
  OAI210     m0207(.A0(mai_mai_n235_), .A1(mai_mai_n234_), .B0(mai_mai_n232_), .Y(mai_mai_n236_));
  AN4        m0208(.A(mai_mai_n236_), .B(mai_mai_n230_), .C(mai_mai_n223_), .D(mai_mai_n219_), .Y(mai_mai_n237_));
  OR2        m0209(.A(h), .B(g), .Y(mai_mai_n238_));
  NO2        m0210(.A(mai_mai_n238_), .B(mai_mai_n97_), .Y(mai_mai_n239_));
  NA2        m0211(.A(mai_mai_n239_), .B(mai_mai_n124_), .Y(mai_mai_n240_));
  NAi41      m0212(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n241_), .B(mai_mai_n208_), .Y(mai_mai_n242_));
  NA2        m0214(.A(mai_mai_n155_), .B(mai_mai_n102_), .Y(mai_mai_n243_));
  NAi21      m0215(.An(mai_mai_n243_), .B(mai_mai_n242_), .Y(mai_mai_n244_));
  NO2        m0216(.A(n), .B(a), .Y(mai_mai_n245_));
  NAi31      m0217(.An(mai_mai_n233_), .B(mai_mai_n245_), .C(mai_mai_n98_), .Y(mai_mai_n246_));
  AN2        m0218(.A(mai_mai_n246_), .B(mai_mai_n244_), .Y(mai_mai_n247_));
  NAi21      m0219(.An(h), .B(i), .Y(mai_mai_n248_));
  NA2        m0220(.A(mai_mai_n175_), .B(k), .Y(mai_mai_n249_));
  NO2        m0221(.A(mai_mai_n249_), .B(mai_mai_n248_), .Y(mai_mai_n250_));
  NA2        m0222(.A(mai_mai_n250_), .B(mai_mai_n187_), .Y(mai_mai_n251_));
  NA3        m0223(.A(mai_mai_n251_), .B(mai_mai_n247_), .C(mai_mai_n240_), .Y(mai_mai_n252_));
  NOi21      m0224(.An(g), .B(e), .Y(mai_mai_n253_));
  NO2        m0225(.A(mai_mai_n67_), .B(mai_mai_n69_), .Y(mai_mai_n254_));
  NA2        m0226(.A(mai_mai_n254_), .B(mai_mai_n253_), .Y(mai_mai_n255_));
  NO2        m0227(.A(mai_mai_n248_), .B(mai_mai_n43_), .Y(mai_mai_n256_));
  NAi21      m0228(.An(f), .B(g), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n257_), .B(mai_mai_n59_), .Y(mai_mai_n258_));
  NO2        m0230(.A(mai_mai_n63_), .B(mai_mai_n111_), .Y(mai_mai_n259_));
  AOI220     m0231(.A0(mai_mai_n259_), .A1(mai_mai_n258_), .B0(mai_mai_n256_), .B1(mai_mai_n61_), .Y(mai_mai_n260_));
  NA2        m0232(.A(mai_mai_n255_), .B(mai_mai_n260_), .Y(mai_mai_n261_));
  NO3        m0233(.A(mai_mai_n127_), .B(mai_mai_n47_), .C(mai_mai_n44_), .Y(mai_mai_n262_));
  NOi41      m0234(.An(mai_mai_n237_), .B(mai_mai_n261_), .C(mai_mai_n252_), .D(mai_mai_n215_), .Y(mai_mai_n263_));
  NO4        m0235(.A(mai_mai_n197_), .B(mai_mai_n46_), .C(mai_mai_n42_), .D(mai_mai_n38_), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n264_), .B(mai_mai_n105_), .Y(mai_mai_n265_));
  NAi21      m0237(.An(h), .B(g), .Y(mai_mai_n266_));
  OR4        m0238(.A(mai_mai_n266_), .B(mai_mai_n1366_), .C(mai_mai_n218_), .D(e), .Y(mai_mai_n267_));
  NO2        m0239(.A(mai_mai_n243_), .B(mai_mai_n257_), .Y(mai_mai_n268_));
  NA2        m0240(.A(mai_mai_n268_), .B(mai_mai_n71_), .Y(mai_mai_n269_));
  NAi31      m0241(.An(g), .B(k), .C(h), .Y(mai_mai_n270_));
  NO3        m0242(.A(mai_mai_n126_), .B(mai_mai_n270_), .C(l), .Y(mai_mai_n271_));
  NAi31      m0243(.An(e), .B(d), .C(a), .Y(mai_mai_n272_));
  NA2        m0244(.A(mai_mai_n271_), .B(mai_mai_n124_), .Y(mai_mai_n273_));
  NA3        m0245(.A(mai_mai_n273_), .B(mai_mai_n269_), .C(mai_mai_n267_), .Y(mai_mai_n274_));
  NA4        m0246(.A(mai_mai_n155_), .B(mai_mai_n74_), .C(mai_mai_n71_), .D(mai_mai_n111_), .Y(mai_mai_n275_));
  NA3        m0247(.A(mai_mai_n155_), .B(mai_mai_n154_), .C(mai_mai_n78_), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n276_), .B(mai_mai_n189_), .Y(mai_mai_n277_));
  NOi21      m0249(.An(mai_mai_n275_), .B(mai_mai_n277_), .Y(mai_mai_n278_));
  NA3        m0250(.A(e), .B(c), .C(b), .Y(mai_mai_n279_));
  NAi32      m0251(.An(k), .Bn(i), .C(j), .Y(mai_mai_n280_));
  INV        m0252(.A(mai_mai_n47_), .Y(mai_mai_n281_));
  NA2        m0253(.A(mai_mai_n258_), .B(mai_mai_n281_), .Y(mai_mai_n282_));
  NAi21      m0254(.An(l), .B(k), .Y(mai_mai_n283_));
  NO2        m0255(.A(mai_mai_n283_), .B(mai_mai_n47_), .Y(mai_mai_n284_));
  NOi21      m0256(.An(l), .B(j), .Y(mai_mai_n285_));
  NA2        m0257(.A(h), .B(mai_mai_n285_), .Y(mai_mai_n286_));
  OR3        m0258(.A(mai_mai_n67_), .B(mai_mai_n69_), .C(e), .Y(mai_mai_n287_));
  NO2        m0259(.A(mai_mai_n286_), .B(mai_mai_n287_), .Y(mai_mai_n288_));
  INV        m0260(.A(mai_mai_n288_), .Y(mai_mai_n289_));
  NAi32      m0261(.An(j), .Bn(h), .C(i), .Y(mai_mai_n290_));
  NAi21      m0262(.An(m), .B(l), .Y(mai_mai_n291_));
  NO3        m0263(.A(mai_mai_n291_), .B(mai_mai_n290_), .C(mai_mai_n78_), .Y(mai_mai_n292_));
  NA2        m0264(.A(h), .B(g), .Y(mai_mai_n293_));
  NA2        m0265(.A(mai_mai_n162_), .B(mai_mai_n44_), .Y(mai_mai_n294_));
  NA2        m0266(.A(mai_mai_n292_), .B(mai_mai_n158_), .Y(mai_mai_n295_));
  NA4        m0267(.A(mai_mai_n295_), .B(mai_mai_n289_), .C(mai_mai_n282_), .D(mai_mai_n278_), .Y(mai_mai_n296_));
  NO2        m0268(.A(mai_mai_n140_), .B(d), .Y(mai_mai_n297_));
  NA2        m0269(.A(mai_mai_n297_), .B(mai_mai_n51_), .Y(mai_mai_n298_));
  NO2        m0270(.A(mai_mai_n100_), .B(mai_mai_n97_), .Y(mai_mai_n299_));
  NAi32      m0271(.An(n), .Bn(m), .C(l), .Y(mai_mai_n300_));
  NO2        m0272(.A(mai_mai_n300_), .B(mai_mai_n290_), .Y(mai_mai_n301_));
  AOI220     m0273(.A0(mai_mai_n301_), .A1(mai_mai_n179_), .B0(mai_mai_n299_), .B1(mai_mai_n56_), .Y(mai_mai_n302_));
  NO2        m0274(.A(mai_mai_n115_), .B(mai_mai_n110_), .Y(mai_mai_n303_));
  INV        m0275(.A(mai_mai_n113_), .Y(mai_mai_n304_));
  NA2        m0276(.A(mai_mai_n304_), .B(mai_mai_n303_), .Y(mai_mai_n305_));
  NA3        m0277(.A(mai_mai_n305_), .B(mai_mai_n302_), .C(mai_mai_n298_), .Y(mai_mai_n306_));
  NO4        m0278(.A(mai_mai_n306_), .B(mai_mai_n296_), .C(mai_mai_n274_), .D(mai_mai_n265_), .Y(mai_mai_n307_));
  NA2        m0279(.A(mai_mai_n250_), .B(mai_mai_n188_), .Y(mai_mai_n308_));
  NAi21      m0280(.An(m), .B(k), .Y(mai_mai_n309_));
  INV        m0281(.A(mai_mai_n309_), .Y(mai_mai_n310_));
  NAi41      m0282(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n311_));
  NO2        m0283(.A(mai_mai_n311_), .B(mai_mai_n146_), .Y(mai_mai_n312_));
  NA2        m0284(.A(mai_mai_n312_), .B(mai_mai_n310_), .Y(mai_mai_n313_));
  NO4        m0285(.A(i), .B(mai_mai_n146_), .C(mai_mai_n67_), .D(mai_mai_n69_), .Y(mai_mai_n314_));
  NA2        m0286(.A(e), .B(c), .Y(mai_mai_n315_));
  NO3        m0287(.A(mai_mai_n315_), .B(n), .C(d), .Y(mai_mai_n316_));
  NA2        m0288(.A(f), .B(mai_mai_n112_), .Y(mai_mai_n317_));
  NO2        m0289(.A(mai_mai_n317_), .B(mai_mai_n209_), .Y(mai_mai_n318_));
  NAi31      m0290(.An(d), .B(e), .C(b), .Y(mai_mai_n319_));
  NO2        m0291(.A(mai_mai_n126_), .B(mai_mai_n319_), .Y(mai_mai_n320_));
  NA2        m0292(.A(mai_mai_n320_), .B(mai_mai_n318_), .Y(mai_mai_n321_));
  NAi41      m0293(.An(mai_mai_n314_), .B(mai_mai_n321_), .C(mai_mai_n313_), .D(mai_mai_n308_), .Y(mai_mai_n322_));
  NO4        m0294(.A(mai_mai_n311_), .B(mai_mai_n73_), .C(mai_mai_n66_), .D(mai_mai_n209_), .Y(mai_mai_n323_));
  NA2        m0295(.A(mai_mai_n245_), .B(mai_mai_n98_), .Y(mai_mai_n324_));
  OR2        m0296(.A(mai_mai_n324_), .B(mai_mai_n199_), .Y(mai_mai_n325_));
  NOi31      m0297(.An(l), .B(n), .C(m), .Y(mai_mai_n326_));
  NA2        m0298(.A(mai_mai_n326_), .B(mai_mai_n210_), .Y(mai_mai_n327_));
  NO2        m0299(.A(mai_mai_n327_), .B(mai_mai_n189_), .Y(mai_mai_n328_));
  NAi32      m0300(.An(mai_mai_n328_), .Bn(mai_mai_n323_), .C(mai_mai_n325_), .Y(mai_mai_n329_));
  NAi32      m0301(.An(m), .Bn(j), .C(k), .Y(mai_mai_n330_));
  NAi41      m0302(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n331_));
  NA2        m0303(.A(mai_mai_n206_), .B(mai_mai_n331_), .Y(mai_mai_n332_));
  NOi31      m0304(.An(j), .B(m), .C(k), .Y(mai_mai_n333_));
  NO2        m0305(.A(mai_mai_n119_), .B(mai_mai_n333_), .Y(mai_mai_n334_));
  AN3        m0306(.A(h), .B(g), .C(f), .Y(mai_mai_n335_));
  NAi31      m0307(.An(mai_mai_n334_), .B(mai_mai_n335_), .C(mai_mai_n332_), .Y(mai_mai_n336_));
  NAi32      m0308(.An(mai_mai_n1357_), .Bn(mai_mai_n196_), .C(mai_mai_n297_), .Y(mai_mai_n337_));
  NO2        m0309(.A(mai_mai_n291_), .B(mai_mai_n290_), .Y(mai_mai_n338_));
  NO2        m0310(.A(mai_mai_n212_), .B(g), .Y(mai_mai_n339_));
  NO2        m0311(.A(mai_mai_n152_), .B(mai_mai_n78_), .Y(mai_mai_n340_));
  AOI220     m0312(.A0(mai_mai_n340_), .A1(mai_mai_n339_), .B0(mai_mai_n242_), .B1(mai_mai_n338_), .Y(mai_mai_n341_));
  NA3        m0313(.A(mai_mai_n341_), .B(mai_mai_n337_), .C(mai_mai_n336_), .Y(mai_mai_n342_));
  NA3        m0314(.A(h), .B(g), .C(f), .Y(mai_mai_n343_));
  NO2        m0315(.A(mai_mai_n343_), .B(mai_mai_n70_), .Y(mai_mai_n344_));
  NA2        m0316(.A(mai_mai_n331_), .B(mai_mai_n206_), .Y(mai_mai_n345_));
  NA2        m0317(.A(h), .B(e), .Y(mai_mai_n346_));
  NO2        m0318(.A(mai_mai_n346_), .B(mai_mai_n40_), .Y(mai_mai_n347_));
  AOI220     m0319(.A0(mai_mai_n347_), .A1(mai_mai_n303_), .B0(mai_mai_n345_), .B1(mai_mai_n344_), .Y(mai_mai_n348_));
  NA3        m0320(.A(g), .B(mai_mai_n283_), .C(mai_mai_n107_), .Y(mai_mai_n349_));
  AO210      m0321(.A0(mai_mai_n105_), .A1(mai_mai_n31_), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  NOi32      m0322(.An(e), .Bn(b), .C(a), .Y(mai_mai_n351_));
  AN2        m0323(.A(l), .B(j), .Y(mai_mai_n352_));
  INV        m0324(.A(mai_mai_n309_), .Y(mai_mai_n353_));
  NO3        m0325(.A(mai_mai_n311_), .B(mai_mai_n66_), .C(mai_mai_n209_), .Y(mai_mai_n354_));
  NA3        m0326(.A(mai_mai_n204_), .B(mai_mai_n202_), .C(mai_mai_n34_), .Y(mai_mai_n355_));
  AOI220     m0327(.A0(mai_mai_n355_), .A1(mai_mai_n351_), .B0(mai_mai_n354_), .B1(mai_mai_n353_), .Y(mai_mai_n356_));
  NO2        m0328(.A(mai_mai_n319_), .B(n), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n203_), .B(k), .Y(mai_mai_n358_));
  NA4        m0330(.A(mai_mai_n198_), .B(mai_mai_n81_), .C(g), .D(mai_mai_n208_), .Y(mai_mai_n359_));
  INV        m0331(.A(mai_mai_n359_), .Y(mai_mai_n360_));
  NAi41      m0332(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n361_));
  NA2        m0333(.A(mai_mai_n49_), .B(mai_mai_n107_), .Y(mai_mai_n362_));
  NO2        m0334(.A(mai_mai_n362_), .B(mai_mai_n361_), .Y(mai_mai_n363_));
  AOI220     m0335(.A0(mai_mai_n363_), .A1(b), .B0(mai_mai_n360_), .B1(mai_mai_n357_), .Y(mai_mai_n364_));
  NA4        m0336(.A(mai_mai_n364_), .B(mai_mai_n356_), .C(mai_mai_n350_), .D(mai_mai_n348_), .Y(mai_mai_n365_));
  NO4        m0337(.A(mai_mai_n365_), .B(mai_mai_n342_), .C(mai_mai_n329_), .D(mai_mai_n322_), .Y(mai_mai_n366_));
  NA4        m0338(.A(mai_mai_n366_), .B(mai_mai_n307_), .C(mai_mai_n263_), .D(mai_mai_n195_), .Y(mai10));
  NA3        m0339(.A(m), .B(k), .C(i), .Y(mai_mai_n368_));
  NO3        m0340(.A(mai_mai_n368_), .B(j), .C(mai_mai_n209_), .Y(mai_mai_n369_));
  NO3        m0341(.A(mai_mai_n147_), .B(n), .C(mai_mai_n104_), .Y(mai_mai_n370_));
  NAi31      m0342(.An(b), .B(f), .C(c), .Y(mai_mai_n371_));
  INV        m0343(.A(mai_mai_n371_), .Y(mai_mai_n372_));
  NOi32      m0344(.An(k), .Bn(h), .C(j), .Y(mai_mai_n373_));
  NA2        m0345(.A(mai_mai_n373_), .B(mai_mai_n216_), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n156_), .B(mai_mai_n374_), .Y(mai_mai_n375_));
  AOI220     m0347(.A0(mai_mai_n375_), .A1(mai_mai_n372_), .B0(mai_mai_n370_), .B1(mai_mai_n369_), .Y(mai_mai_n376_));
  AN2        m0348(.A(j), .B(h), .Y(mai_mai_n377_));
  NO3        m0349(.A(n), .B(m), .C(k), .Y(mai_mai_n378_));
  NA2        m0350(.A(mai_mai_n378_), .B(mai_mai_n377_), .Y(mai_mai_n379_));
  NO3        m0351(.A(mai_mai_n379_), .B(mai_mai_n147_), .C(mai_mai_n208_), .Y(mai_mai_n380_));
  OR2        m0352(.A(m), .B(k), .Y(mai_mai_n381_));
  NO2        m0353(.A(mai_mai_n169_), .B(mai_mai_n381_), .Y(mai_mai_n382_));
  NA4        m0354(.A(n), .B(f), .C(c), .D(mai_mai_n110_), .Y(mai_mai_n383_));
  NOi21      m0355(.An(mai_mai_n382_), .B(mai_mai_n383_), .Y(mai_mai_n384_));
  NOi32      m0356(.An(d), .Bn(a), .C(c), .Y(mai_mai_n385_));
  NA2        m0357(.A(mai_mai_n385_), .B(mai_mai_n177_), .Y(mai_mai_n386_));
  NAi21      m0358(.An(i), .B(g), .Y(mai_mai_n387_));
  NAi31      m0359(.An(k), .B(m), .C(j), .Y(mai_mai_n388_));
  NO3        m0360(.A(mai_mai_n388_), .B(mai_mai_n387_), .C(n), .Y(mai_mai_n389_));
  NOi21      m0361(.An(mai_mai_n389_), .B(mai_mai_n386_), .Y(mai_mai_n390_));
  NO3        m0362(.A(mai_mai_n390_), .B(mai_mai_n384_), .C(mai_mai_n380_), .Y(mai_mai_n391_));
  NO2        m0363(.A(mai_mai_n383_), .B(mai_mai_n291_), .Y(mai_mai_n392_));
  NOi32      m0364(.An(f), .Bn(d), .C(c), .Y(mai_mai_n393_));
  AOI220     m0365(.A0(mai_mai_n393_), .A1(mai_mai_n301_), .B0(mai_mai_n392_), .B1(mai_mai_n210_), .Y(mai_mai_n394_));
  NA3        m0366(.A(mai_mai_n394_), .B(mai_mai_n391_), .C(mai_mai_n376_), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n56_), .B(mai_mai_n110_), .Y(mai_mai_n396_));
  NA2        m0368(.A(mai_mai_n245_), .B(mai_mai_n396_), .Y(mai_mai_n397_));
  INV        m0369(.A(e), .Y(mai_mai_n398_));
  NA2        m0370(.A(mai_mai_n45_), .B(e), .Y(mai_mai_n399_));
  OAI210     m0371(.A0(mai_mai_n399_), .A1(mai_mai_n1358_), .B0(mai_mai_n199_), .Y(mai_mai_n400_));
  AN2        m0372(.A(g), .B(e), .Y(mai_mai_n401_));
  NA3        m0373(.A(mai_mai_n401_), .B(mai_mai_n198_), .C(i), .Y(mai_mai_n402_));
  NA2        m0374(.A(mai_mai_n83_), .B(mai_mai_n402_), .Y(mai_mai_n403_));
  NO2        m0375(.A(mai_mai_n94_), .B(mai_mai_n398_), .Y(mai_mai_n404_));
  NO3        m0376(.A(mai_mai_n404_), .B(mai_mai_n403_), .C(mai_mai_n400_), .Y(mai_mai_n405_));
  NOi32      m0377(.An(h), .Bn(e), .C(g), .Y(mai_mai_n406_));
  NA3        m0378(.A(mai_mai_n406_), .B(mai_mai_n285_), .C(m), .Y(mai_mai_n407_));
  NOi21      m0379(.An(g), .B(h), .Y(mai_mai_n408_));
  NA3        m0380(.A(m), .B(mai_mai_n408_), .C(e), .Y(mai_mai_n409_));
  AN3        m0381(.A(h), .B(g), .C(e), .Y(mai_mai_n410_));
  NA2        m0382(.A(mai_mai_n410_), .B(m), .Y(mai_mai_n411_));
  AN3        m0383(.A(mai_mai_n411_), .B(mai_mai_n409_), .C(mai_mai_n407_), .Y(mai_mai_n412_));
  AOI210     m0384(.A0(mai_mai_n412_), .A1(mai_mai_n405_), .B0(mai_mai_n397_), .Y(mai_mai_n413_));
  NA3        m0385(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(e), .Y(mai_mai_n414_));
  NO2        m0386(.A(mai_mai_n414_), .B(mai_mai_n397_), .Y(mai_mai_n415_));
  NA3        m0387(.A(mai_mai_n385_), .B(mai_mai_n177_), .C(mai_mai_n78_), .Y(mai_mai_n416_));
  NAi31      m0388(.An(b), .B(c), .C(a), .Y(mai_mai_n417_));
  NO2        m0389(.A(mai_mai_n417_), .B(n), .Y(mai_mai_n418_));
  OAI210     m0390(.A0(mai_mai_n49_), .A1(mai_mai_n48_), .B0(m), .Y(mai_mai_n419_));
  NO2        m0391(.A(mai_mai_n419_), .B(mai_mai_n143_), .Y(mai_mai_n420_));
  NA2        m0392(.A(mai_mai_n420_), .B(mai_mai_n418_), .Y(mai_mai_n421_));
  INV        m0393(.A(mai_mai_n421_), .Y(mai_mai_n422_));
  NO4        m0394(.A(mai_mai_n422_), .B(mai_mai_n415_), .C(mai_mai_n413_), .D(mai_mai_n395_), .Y(mai_mai_n423_));
  NA2        m0395(.A(i), .B(g), .Y(mai_mai_n424_));
  NO3        m0396(.A(mai_mai_n272_), .B(mai_mai_n424_), .C(c), .Y(mai_mai_n425_));
  NOi21      m0397(.An(a), .B(n), .Y(mai_mai_n426_));
  NA2        m0398(.A(d), .B(mai_mai_n426_), .Y(mai_mai_n427_));
  NA3        m0399(.A(i), .B(g), .C(f), .Y(mai_mai_n428_));
  OR2        m0400(.A(mai_mai_n428_), .B(mai_mai_n65_), .Y(mai_mai_n429_));
  NA3        m0401(.A(m), .B(mai_mai_n408_), .C(mai_mai_n177_), .Y(mai_mai_n430_));
  AOI210     m0402(.A0(mai_mai_n430_), .A1(mai_mai_n429_), .B0(mai_mai_n427_), .Y(mai_mai_n431_));
  AOI210     m0403(.A0(mai_mai_n425_), .A1(mai_mai_n284_), .B0(mai_mai_n431_), .Y(mai_mai_n432_));
  OR2        m0404(.A(n), .B(m), .Y(mai_mai_n433_));
  NO2        m0405(.A(mai_mai_n433_), .B(mai_mai_n148_), .Y(mai_mai_n434_));
  NO2        m0406(.A(mai_mai_n178_), .B(mai_mai_n143_), .Y(mai_mai_n435_));
  OAI210     m0407(.A0(mai_mai_n434_), .A1(mai_mai_n171_), .B0(mai_mai_n435_), .Y(mai_mai_n436_));
  INV        m0408(.A(mai_mai_n362_), .Y(mai_mai_n437_));
  NA3        m0409(.A(mai_mai_n437_), .B(mai_mai_n351_), .C(d), .Y(mai_mai_n438_));
  NO2        m0410(.A(mai_mai_n417_), .B(mai_mai_n47_), .Y(mai_mai_n439_));
  NAi21      m0411(.An(k), .B(j), .Y(mai_mai_n440_));
  NA3        m0412(.A(i), .B(g), .C(mai_mai_n439_), .Y(mai_mai_n441_));
  NAi21      m0413(.An(e), .B(d), .Y(mai_mai_n442_));
  NO2        m0414(.A(mai_mai_n442_), .B(mai_mai_n53_), .Y(mai_mai_n443_));
  NO2        m0415(.A(mai_mai_n249_), .B(mai_mai_n208_), .Y(mai_mai_n444_));
  NA2        m0416(.A(mai_mai_n444_), .B(mai_mai_n443_), .Y(mai_mai_n445_));
  NA4        m0417(.A(mai_mai_n445_), .B(mai_mai_n441_), .C(mai_mai_n438_), .D(mai_mai_n436_), .Y(mai_mai_n446_));
  NO2        m0418(.A(mai_mai_n327_), .B(mai_mai_n208_), .Y(mai_mai_n447_));
  NA2        m0419(.A(mai_mai_n447_), .B(mai_mai_n443_), .Y(mai_mai_n448_));
  NOi31      m0420(.An(n), .B(m), .C(k), .Y(mai_mai_n449_));
  AOI220     m0421(.A0(mai_mai_n449_), .A1(mai_mai_n377_), .B0(mai_mai_n216_), .B1(mai_mai_n48_), .Y(mai_mai_n450_));
  NAi31      m0422(.An(g), .B(f), .C(c), .Y(mai_mai_n451_));
  OR3        m0423(.A(mai_mai_n451_), .B(mai_mai_n450_), .C(e), .Y(mai_mai_n452_));
  NA3        m0424(.A(mai_mai_n452_), .B(mai_mai_n448_), .C(mai_mai_n302_), .Y(mai_mai_n453_));
  NOi41      m0425(.An(mai_mai_n432_), .B(mai_mai_n453_), .C(mai_mai_n446_), .D(mai_mai_n261_), .Y(mai_mai_n454_));
  NOi32      m0426(.An(c), .Bn(a), .C(b), .Y(mai_mai_n455_));
  NA2        m0427(.A(mai_mai_n455_), .B(mai_mai_n107_), .Y(mai_mai_n456_));
  AN2        m0428(.A(e), .B(d), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n125_), .B(mai_mai_n40_), .Y(mai_mai_n458_));
  NO2        m0430(.A(mai_mai_n60_), .B(e), .Y(mai_mai_n459_));
  AOI210     m0431(.A0(mai_mai_n458_), .A1(f), .B0(mai_mai_n459_), .Y(mai_mai_n460_));
  AOI210     m0432(.A0(mai_mai_n460_), .A1(mai_mai_n270_), .B0(mai_mai_n456_), .Y(mai_mai_n461_));
  NO2        m0433(.A(mai_mai_n205_), .B(mai_mai_n200_), .Y(mai_mai_n462_));
  NA3        m0434(.A(e), .B(d), .C(c), .Y(mai_mai_n463_));
  NAi21      m0435(.An(mai_mai_n463_), .B(a), .Y(mai_mai_n464_));
  NO2        m0436(.A(mai_mai_n416_), .B(mai_mai_n199_), .Y(mai_mai_n465_));
  NOi21      m0437(.An(mai_mai_n464_), .B(mai_mai_n465_), .Y(mai_mai_n466_));
  AOI210     m0438(.A0(mai_mai_n264_), .A1(mai_mai_n462_), .B0(mai_mai_n466_), .Y(mai_mai_n467_));
  NO4        m0439(.A(mai_mai_n183_), .B(mai_mai_n97_), .C(mai_mai_n53_), .D(b), .Y(mai_mai_n468_));
  NA2        m0440(.A(mai_mai_n372_), .B(mai_mai_n149_), .Y(mai_mai_n469_));
  NA2        m0441(.A(l), .B(k), .Y(mai_mai_n470_));
  AOI210     m0442(.A0(mai_mai_n227_), .A1(mai_mai_n330_), .B0(mai_mai_n78_), .Y(mai_mai_n471_));
  OR3        m0443(.A(mai_mai_n1362_), .B(mai_mai_n139_), .C(mai_mai_n129_), .Y(mai_mai_n472_));
  NA3        m0444(.A(mai_mai_n275_), .B(mai_mai_n122_), .C(mai_mai_n120_), .Y(mai_mai_n473_));
  NA2        m0445(.A(mai_mai_n385_), .B(mai_mai_n107_), .Y(mai_mai_n474_));
  NO4        m0446(.A(mai_mai_n474_), .B(mai_mai_n89_), .C(mai_mai_n106_), .D(e), .Y(mai_mai_n475_));
  NO3        m0447(.A(mai_mai_n416_), .B(mai_mai_n86_), .C(mai_mai_n125_), .Y(mai_mai_n476_));
  NO4        m0448(.A(mai_mai_n476_), .B(mai_mai_n475_), .C(mai_mai_n473_), .D(mai_mai_n314_), .Y(mai_mai_n477_));
  NA3        m0449(.A(mai_mai_n477_), .B(mai_mai_n472_), .C(mai_mai_n469_), .Y(mai_mai_n478_));
  NO4        m0450(.A(mai_mai_n478_), .B(mai_mai_n468_), .C(mai_mai_n467_), .D(mai_mai_n461_), .Y(mai_mai_n479_));
  NA2        m0451(.A(mai_mai_n64_), .B(mai_mai_n61_), .Y(mai_mai_n480_));
  NOi21      m0452(.An(d), .B(e), .Y(mai_mai_n481_));
  NO2        m0453(.A(mai_mai_n183_), .B(mai_mai_n53_), .Y(mai_mai_n482_));
  NAi31      m0454(.An(j), .B(l), .C(i), .Y(mai_mai_n483_));
  OAI210     m0455(.A0(mai_mai_n483_), .A1(mai_mai_n126_), .B0(mai_mai_n97_), .Y(mai_mai_n484_));
  NA3        m0456(.A(mai_mai_n484_), .B(mai_mai_n482_), .C(b), .Y(mai_mai_n485_));
  NO3        m0457(.A(mai_mai_n386_), .B(mai_mai_n1357_), .C(mai_mai_n196_), .Y(mai_mai_n486_));
  NO2        m0458(.A(mai_mai_n386_), .B(mai_mai_n362_), .Y(mai_mai_n487_));
  NO4        m0459(.A(mai_mai_n487_), .B(mai_mai_n486_), .C(mai_mai_n180_), .D(mai_mai_n299_), .Y(mai_mai_n488_));
  NA4        m0460(.A(mai_mai_n488_), .B(mai_mai_n485_), .C(mai_mai_n480_), .D(mai_mai_n237_), .Y(mai_mai_n489_));
  OAI210     m0461(.A0(mai_mai_n121_), .A1(mai_mai_n119_), .B0(n), .Y(mai_mai_n490_));
  NO2        m0462(.A(mai_mai_n490_), .B(mai_mai_n125_), .Y(mai_mai_n491_));
  AO210      m0463(.A0(mai_mai_n292_), .A1(mai_mai_n209_), .B0(mai_mai_n239_), .Y(mai_mai_n492_));
  OA210      m0464(.A0(mai_mai_n492_), .A1(mai_mai_n491_), .B0(mai_mai_n188_), .Y(mai_mai_n493_));
  XO2        m0465(.A(i), .B(h), .Y(mai_mai_n494_));
  NA3        m0466(.A(mai_mai_n494_), .B(mai_mai_n155_), .C(n), .Y(mai_mai_n495_));
  NAi41      m0467(.An(mai_mai_n292_), .B(mai_mai_n495_), .C(mai_mai_n450_), .D(mai_mai_n374_), .Y(mai_mai_n496_));
  NOi32      m0468(.An(mai_mai_n496_), .Bn(mai_mai_n459_), .C(mai_mai_n1366_), .Y(mai_mai_n497_));
  NAi31      m0469(.An(c), .B(f), .C(d), .Y(mai_mai_n498_));
  AOI210     m0470(.A0(mai_mai_n276_), .A1(mai_mai_n191_), .B0(mai_mai_n498_), .Y(mai_mai_n499_));
  NOi21      m0471(.An(mai_mai_n76_), .B(mai_mai_n499_), .Y(mai_mai_n500_));
  NA3        m0472(.A(mai_mai_n370_), .B(m), .C(mai_mai_n91_), .Y(mai_mai_n501_));
  NA2        m0473(.A(mai_mai_n221_), .B(mai_mai_n102_), .Y(mai_mai_n502_));
  AOI210     m0474(.A0(mai_mai_n502_), .A1(mai_mai_n176_), .B0(mai_mai_n498_), .Y(mai_mai_n503_));
  AOI210     m0475(.A0(mai_mai_n349_), .A1(mai_mai_n34_), .B0(mai_mai_n464_), .Y(mai_mai_n504_));
  NOi31      m0476(.An(mai_mai_n501_), .B(mai_mai_n504_), .C(mai_mai_n503_), .Y(mai_mai_n505_));
  AO220      m0477(.A0(mai_mai_n281_), .A1(mai_mai_n258_), .B0(mai_mai_n160_), .B1(mai_mai_n61_), .Y(mai_mai_n506_));
  NA3        m0478(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(f), .Y(mai_mai_n507_));
  NO2        m0479(.A(mai_mai_n507_), .B(mai_mai_n427_), .Y(mai_mai_n508_));
  NO2        m0480(.A(mai_mai_n508_), .B(mai_mai_n288_), .Y(mai_mai_n509_));
  NAi41      m0481(.An(mai_mai_n506_), .B(mai_mai_n509_), .C(mai_mai_n505_), .D(mai_mai_n500_), .Y(mai_mai_n510_));
  NO4        m0482(.A(mai_mai_n510_), .B(mai_mai_n497_), .C(mai_mai_n493_), .D(mai_mai_n489_), .Y(mai_mai_n511_));
  NA4        m0483(.A(mai_mai_n511_), .B(mai_mai_n479_), .C(mai_mai_n454_), .D(mai_mai_n423_), .Y(mai11));
  NO2        m0484(.A(mai_mai_n67_), .B(f), .Y(mai_mai_n513_));
  NA2        m0485(.A(j), .B(g), .Y(mai_mai_n514_));
  NAi31      m0486(.An(i), .B(m), .C(l), .Y(mai_mai_n515_));
  NA3        m0487(.A(m), .B(k), .C(j), .Y(mai_mai_n516_));
  OAI220     m0488(.A0(mai_mai_n516_), .A1(mai_mai_n125_), .B0(mai_mai_n515_), .B1(mai_mai_n514_), .Y(mai_mai_n517_));
  NA2        m0489(.A(mai_mai_n517_), .B(mai_mai_n513_), .Y(mai_mai_n518_));
  NOi32      m0490(.An(e), .Bn(b), .C(f), .Y(mai_mai_n519_));
  NA2        m0491(.A(j), .B(mai_mai_n107_), .Y(mai_mai_n520_));
  NA2        m0492(.A(mai_mai_n45_), .B(j), .Y(mai_mai_n521_));
  OAI220     m0493(.A0(mai_mai_n521_), .A1(mai_mai_n294_), .B0(mai_mai_n520_), .B1(mai_mai_n209_), .Y(mai_mai_n522_));
  NAi31      m0494(.An(d), .B(e), .C(a), .Y(mai_mai_n523_));
  NO2        m0495(.A(mai_mai_n523_), .B(n), .Y(mai_mai_n524_));
  AOI220     m0496(.A0(mai_mai_n524_), .A1(mai_mai_n95_), .B0(mai_mai_n522_), .B1(mai_mai_n519_), .Y(mai_mai_n525_));
  NAi41      m0497(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n526_));
  NO2        m0498(.A(mai_mai_n386_), .B(mai_mai_n266_), .Y(mai_mai_n527_));
  NA2        m0499(.A(j), .B(i), .Y(mai_mai_n528_));
  NAi31      m0500(.An(n), .B(m), .C(k), .Y(mai_mai_n529_));
  NO3        m0501(.A(mai_mai_n529_), .B(mai_mai_n528_), .C(mai_mai_n106_), .Y(mai_mai_n530_));
  NO4        m0502(.A(n), .B(d), .C(mai_mai_n110_), .D(a), .Y(mai_mai_n531_));
  OR2        m0503(.A(n), .B(c), .Y(mai_mai_n532_));
  NO2        m0504(.A(mai_mai_n532_), .B(mai_mai_n145_), .Y(mai_mai_n533_));
  NO2        m0505(.A(mai_mai_n533_), .B(mai_mai_n531_), .Y(mai_mai_n534_));
  NOi32      m0506(.An(g), .Bn(f), .C(i), .Y(mai_mai_n535_));
  AOI220     m0507(.A0(mai_mai_n535_), .A1(mai_mai_n93_), .B0(mai_mai_n517_), .B1(f), .Y(mai_mai_n536_));
  NO2        m0508(.A(mai_mai_n270_), .B(mai_mai_n47_), .Y(mai_mai_n537_));
  NO2        m0509(.A(mai_mai_n536_), .B(mai_mai_n534_), .Y(mai_mai_n538_));
  AOI210     m0510(.A0(mai_mai_n530_), .A1(mai_mai_n527_), .B0(mai_mai_n538_), .Y(mai_mai_n539_));
  NA2        m0511(.A(mai_mai_n135_), .B(mai_mai_n33_), .Y(mai_mai_n540_));
  OAI220     m0512(.A0(mai_mai_n540_), .A1(m), .B0(mai_mai_n521_), .B1(mai_mai_n227_), .Y(mai_mai_n541_));
  NOi41      m0513(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n542_));
  NAi32      m0514(.An(e), .Bn(b), .C(c), .Y(mai_mai_n543_));
  AN2        m0515(.A(mai_mai_n331_), .B(mai_mai_n311_), .Y(mai_mai_n544_));
  NA2        m0516(.A(mai_mai_n544_), .B(mai_mai_n543_), .Y(mai_mai_n545_));
  OA210      m0517(.A0(mai_mai_n545_), .A1(mai_mai_n542_), .B0(mai_mai_n541_), .Y(mai_mai_n546_));
  OAI220     m0518(.A0(mai_mai_n388_), .A1(mai_mai_n387_), .B0(mai_mai_n515_), .B1(mai_mai_n514_), .Y(mai_mai_n547_));
  NAi31      m0519(.An(d), .B(c), .C(a), .Y(mai_mai_n548_));
  NO2        m0520(.A(mai_mai_n548_), .B(n), .Y(mai_mai_n549_));
  NA3        m0521(.A(mai_mai_n549_), .B(mai_mai_n547_), .C(e), .Y(mai_mai_n550_));
  NO3        m0522(.A(mai_mai_n58_), .B(mai_mai_n47_), .C(mai_mai_n209_), .Y(mai_mai_n551_));
  NO2        m0523(.A(mai_mai_n224_), .B(mai_mai_n104_), .Y(mai_mai_n552_));
  OAI210     m0524(.A0(mai_mai_n551_), .A1(mai_mai_n389_), .B0(mai_mai_n552_), .Y(mai_mai_n553_));
  NA2        m0525(.A(mai_mai_n553_), .B(mai_mai_n550_), .Y(mai_mai_n554_));
  NO2        m0526(.A(mai_mai_n272_), .B(n), .Y(mai_mai_n555_));
  NO2        m0527(.A(mai_mai_n418_), .B(mai_mai_n555_), .Y(mai_mai_n556_));
  NA2        m0528(.A(mai_mai_n547_), .B(f), .Y(mai_mai_n557_));
  NAi32      m0529(.An(d), .Bn(a), .C(b), .Y(mai_mai_n558_));
  NO2        m0530(.A(mai_mai_n558_), .B(mai_mai_n47_), .Y(mai_mai_n559_));
  INV        m0531(.A(mai_mai_n89_), .Y(mai_mai_n560_));
  NO3        m0532(.A(mai_mai_n172_), .B(mai_mai_n169_), .C(g), .Y(mai_mai_n561_));
  AOI220     m0533(.A0(mai_mai_n561_), .A1(mai_mai_n55_), .B0(mai_mai_n560_), .B1(mai_mai_n559_), .Y(mai_mai_n562_));
  OAI210     m0534(.A0(mai_mai_n557_), .A1(mai_mai_n556_), .B0(mai_mai_n562_), .Y(mai_mai_n563_));
  NO2        m0535(.A(mai_mai_n142_), .B(c), .Y(mai_mai_n564_));
  NA3        m0536(.A(mai_mai_n564_), .B(h), .C(mai_mai_n449_), .Y(mai_mai_n565_));
  NA3        m0537(.A(f), .B(d), .C(b), .Y(mai_mai_n566_));
  NO4        m0538(.A(mai_mai_n566_), .B(mai_mai_n172_), .C(mai_mai_n169_), .D(g), .Y(mai_mai_n567_));
  NAi21      m0539(.An(mai_mai_n567_), .B(mai_mai_n565_), .Y(mai_mai_n568_));
  NO4        m0540(.A(mai_mai_n568_), .B(mai_mai_n563_), .C(mai_mai_n554_), .D(mai_mai_n546_), .Y(mai_mai_n569_));
  AN4        m0541(.A(mai_mai_n569_), .B(mai_mai_n539_), .C(mai_mai_n525_), .D(mai_mai_n518_), .Y(mai_mai_n570_));
  INV        m0542(.A(k), .Y(mai_mai_n571_));
  INV        m0543(.A(k), .Y(mai_mai_n572_));
  NA4        m0544(.A(mai_mai_n385_), .B(mai_mai_n408_), .C(mai_mai_n177_), .D(mai_mai_n107_), .Y(mai_mai_n573_));
  NAi32      m0545(.An(h), .Bn(f), .C(g), .Y(mai_mai_n574_));
  NAi41      m0546(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n575_));
  OAI210     m0547(.A0(mai_mai_n523_), .A1(n), .B0(mai_mai_n575_), .Y(mai_mai_n576_));
  NA2        m0548(.A(mai_mai_n576_), .B(m), .Y(mai_mai_n577_));
  NAi31      m0549(.An(h), .B(g), .C(f), .Y(mai_mai_n578_));
  OR3        m0550(.A(mai_mai_n578_), .B(mai_mai_n272_), .C(mai_mai_n47_), .Y(mai_mai_n579_));
  NA4        m0551(.A(mai_mai_n408_), .B(mai_mai_n114_), .C(mai_mai_n107_), .D(e), .Y(mai_mai_n580_));
  AN2        m0552(.A(mai_mai_n580_), .B(mai_mai_n579_), .Y(mai_mai_n581_));
  OA210      m0553(.A0(mai_mai_n577_), .A1(mai_mai_n574_), .B0(mai_mai_n581_), .Y(mai_mai_n582_));
  NO3        m0554(.A(mai_mai_n574_), .B(mai_mai_n67_), .C(mai_mai_n69_), .Y(mai_mai_n583_));
  NO4        m0555(.A(mai_mai_n578_), .B(mai_mai_n532_), .C(mai_mai_n145_), .D(mai_mai_n69_), .Y(mai_mai_n584_));
  OR2        m0556(.A(mai_mai_n584_), .B(mai_mai_n583_), .Y(mai_mai_n585_));
  NAi31      m0557(.An(mai_mai_n585_), .B(mai_mai_n582_), .C(mai_mai_n573_), .Y(mai_mai_n586_));
  NAi31      m0558(.An(f), .B(h), .C(g), .Y(mai_mai_n587_));
  NO4        m0559(.A(k), .B(mai_mai_n587_), .C(mai_mai_n67_), .D(mai_mai_n69_), .Y(mai_mai_n588_));
  NOi41      m0560(.An(b), .B(mai_mai_n343_), .C(mai_mai_n63_), .D(mai_mai_n111_), .Y(mai_mai_n589_));
  OR2        m0561(.A(mai_mai_n589_), .B(mai_mai_n588_), .Y(mai_mai_n590_));
  NA2        m0562(.A(a), .B(mai_mai_n107_), .Y(mai_mai_n591_));
  NO2        m0563(.A(n), .B(c), .Y(mai_mai_n592_));
  NA3        m0564(.A(mai_mai_n592_), .B(a), .C(m), .Y(mai_mai_n593_));
  NOi32      m0565(.An(e), .Bn(a), .C(d), .Y(mai_mai_n594_));
  AOI210     m0566(.A0(a), .A1(d), .B0(mai_mai_n594_), .Y(mai_mai_n595_));
  INV        m0567(.A(mai_mai_n540_), .Y(mai_mai_n596_));
  AOI210     m0568(.A0(mai_mai_n596_), .A1(mai_mai_n107_), .B0(mai_mai_n590_), .Y(mai_mai_n597_));
  OAI210     m0569(.A0(mai_mai_n244_), .A1(mai_mai_n81_), .B0(mai_mai_n597_), .Y(mai_mai_n598_));
  AOI210     m0570(.A0(mai_mai_n586_), .A1(mai_mai_n572_), .B0(mai_mai_n598_), .Y(mai_mai_n599_));
  NO3        m0571(.A(mai_mai_n309_), .B(mai_mai_n57_), .C(n), .Y(mai_mai_n600_));
  NA3        m0572(.A(mai_mai_n498_), .B(mai_mai_n167_), .C(mai_mai_n166_), .Y(mai_mai_n601_));
  NA2        m0573(.A(mai_mai_n451_), .B(mai_mai_n224_), .Y(mai_mai_n602_));
  OR2        m0574(.A(mai_mai_n602_), .B(mai_mai_n601_), .Y(mai_mai_n603_));
  NA2        m0575(.A(k), .B(mai_mai_n107_), .Y(mai_mai_n604_));
  AOI220     m0576(.A0(mai_mai_n107_), .A1(mai_mai_n527_), .B0(mai_mai_n603_), .B1(mai_mai_n600_), .Y(mai_mai_n605_));
  NO2        m0577(.A(mai_mai_n605_), .B(mai_mai_n81_), .Y(mai_mai_n606_));
  NA3        m0578(.A(mai_mai_n542_), .B(mai_mai_n333_), .C(mai_mai_n45_), .Y(mai_mai_n607_));
  NOi32      m0579(.An(e), .Bn(c), .C(f), .Y(mai_mai_n608_));
  INV        m0580(.A(mai_mai_n206_), .Y(mai_mai_n609_));
  AOI220     m0581(.A0(mai_mai_n609_), .A1(mai_mai_n382_), .B0(mai_mai_n608_), .B1(mai_mai_n171_), .Y(mai_mai_n610_));
  NA3        m0582(.A(mai_mai_n610_), .B(mai_mai_n607_), .C(mai_mai_n174_), .Y(mai_mai_n611_));
  AOI210     m0583(.A0(mai_mai_n1370_), .A1(mai_mai_n386_), .B0(mai_mai_n293_), .Y(mai_mai_n612_));
  NA2        m0584(.A(mai_mai_n612_), .B(mai_mai_n259_), .Y(mai_mai_n613_));
  NAi21      m0585(.An(k), .B(h), .Y(mai_mai_n614_));
  NO2        m0586(.A(mai_mai_n614_), .B(mai_mai_n257_), .Y(mai_mai_n615_));
  NA2        m0587(.A(mai_mai_n615_), .B(j), .Y(mai_mai_n616_));
  OR2        m0588(.A(mai_mai_n616_), .B(mai_mai_n577_), .Y(mai_mai_n617_));
  NOi31      m0589(.An(m), .B(n), .C(k), .Y(mai_mai_n618_));
  NA2        m0590(.A(j), .B(mai_mai_n618_), .Y(mai_mai_n619_));
  AOI210     m0591(.A0(mai_mai_n386_), .A1(mai_mai_n361_), .B0(mai_mai_n293_), .Y(mai_mai_n620_));
  NAi21      m0592(.An(mai_mai_n619_), .B(mai_mai_n620_), .Y(mai_mai_n621_));
  NO2        m0593(.A(mai_mai_n272_), .B(mai_mai_n47_), .Y(mai_mai_n622_));
  NO2        m0594(.A(k), .B(mai_mai_n587_), .Y(mai_mai_n623_));
  NO2        m0595(.A(mai_mai_n523_), .B(mai_mai_n47_), .Y(mai_mai_n624_));
  AOI220     m0596(.A0(mai_mai_n624_), .A1(mai_mai_n623_), .B0(mai_mai_n622_), .B1(mai_mai_n560_), .Y(mai_mai_n625_));
  NA4        m0597(.A(mai_mai_n625_), .B(mai_mai_n621_), .C(mai_mai_n617_), .D(mai_mai_n613_), .Y(mai_mai_n626_));
  NA2        m0598(.A(mai_mai_n102_), .B(mai_mai_n35_), .Y(mai_mai_n627_));
  NO2        m0599(.A(k), .B(mai_mai_n209_), .Y(mai_mai_n628_));
  NO2        m0600(.A(mai_mai_n519_), .B(mai_mai_n351_), .Y(mai_mai_n629_));
  NO2        m0601(.A(mai_mai_n629_), .B(n), .Y(mai_mai_n630_));
  NAi31      m0602(.An(mai_mai_n627_), .B(mai_mai_n630_), .C(mai_mai_n628_), .Y(mai_mai_n631_));
  NO2        m0603(.A(mai_mai_n521_), .B(mai_mai_n172_), .Y(mai_mai_n632_));
  NA2        m0604(.A(mai_mai_n494_), .B(mai_mai_n155_), .Y(mai_mai_n633_));
  NO3        m0605(.A(mai_mai_n383_), .B(mai_mai_n633_), .C(mai_mai_n81_), .Y(mai_mai_n634_));
  AOI210     m0606(.A0(c), .A1(mai_mai_n632_), .B0(mai_mai_n634_), .Y(mai_mai_n635_));
  AN3        m0607(.A(f), .B(d), .C(b), .Y(mai_mai_n636_));
  OAI210     m0608(.A0(mai_mai_n636_), .A1(mai_mai_n124_), .B0(n), .Y(mai_mai_n637_));
  NA3        m0609(.A(mai_mai_n494_), .B(mai_mai_n155_), .C(mai_mai_n209_), .Y(mai_mai_n638_));
  AOI210     m0610(.A0(mai_mai_n637_), .A1(mai_mai_n226_), .B0(mai_mai_n638_), .Y(mai_mai_n639_));
  NAi31      m0611(.An(m), .B(n), .C(k), .Y(mai_mai_n640_));
  OAI210     m0612(.A0(mai_mai_n129_), .A1(mai_mai_n640_), .B0(mai_mai_n246_), .Y(mai_mai_n641_));
  OAI210     m0613(.A0(mai_mai_n641_), .A1(mai_mai_n639_), .B0(j), .Y(mai_mai_n642_));
  NA3        m0614(.A(mai_mai_n642_), .B(mai_mai_n635_), .C(mai_mai_n631_), .Y(mai_mai_n643_));
  NO4        m0615(.A(mai_mai_n643_), .B(mai_mai_n626_), .C(mai_mai_n611_), .D(mai_mai_n606_), .Y(mai_mai_n644_));
  NA2        m0616(.A(mai_mai_n370_), .B(h), .Y(mai_mai_n645_));
  NAi31      m0617(.An(g), .B(h), .C(f), .Y(mai_mai_n646_));
  OR3        m0618(.A(mai_mai_n646_), .B(mai_mai_n272_), .C(n), .Y(mai_mai_n647_));
  OA210      m0619(.A0(mai_mai_n523_), .A1(n), .B0(mai_mai_n575_), .Y(mai_mai_n648_));
  NA3        m0620(.A(mai_mai_n406_), .B(mai_mai_n114_), .C(mai_mai_n78_), .Y(mai_mai_n649_));
  OAI210     m0621(.A0(mai_mai_n648_), .A1(mai_mai_n85_), .B0(mai_mai_n649_), .Y(mai_mai_n650_));
  NOi21      m0622(.An(mai_mai_n647_), .B(mai_mai_n650_), .Y(mai_mai_n651_));
  AOI210     m0623(.A0(mai_mai_n651_), .A1(mai_mai_n645_), .B0(mai_mai_n516_), .Y(mai_mai_n652_));
  NO3        m0624(.A(g), .B(mai_mai_n208_), .C(mai_mai_n53_), .Y(mai_mai_n653_));
  NAi21      m0625(.An(h), .B(j), .Y(mai_mai_n654_));
  OAI220     m0626(.A0(mai_mai_n654_), .A1(mai_mai_n97_), .B0(mai_mai_n502_), .B1(mai_mai_n81_), .Y(mai_mai_n655_));
  OAI210     m0627(.A0(mai_mai_n655_), .A1(mai_mai_n382_), .B0(mai_mai_n653_), .Y(mai_mai_n656_));
  NA2        m0628(.A(b), .B(mai_mai_n335_), .Y(mai_mai_n657_));
  OA220      m0629(.A0(mai_mai_n619_), .A1(mai_mai_n657_), .B0(mai_mai_n616_), .B1(mai_mai_n67_), .Y(mai_mai_n658_));
  NA3        m0630(.A(mai_mai_n513_), .B(mai_mai_n93_), .C(mai_mai_n92_), .Y(mai_mai_n659_));
  NA2        m0631(.A(h), .B(mai_mai_n36_), .Y(mai_mai_n660_));
  NA2        m0632(.A(mai_mai_n93_), .B(mai_mai_n45_), .Y(mai_mai_n661_));
  OAI220     m0633(.A0(mai_mai_n661_), .A1(mai_mai_n324_), .B0(mai_mai_n660_), .B1(mai_mai_n456_), .Y(mai_mai_n662_));
  AOI210     m0634(.A0(mai_mai_n558_), .A1(mai_mai_n417_), .B0(mai_mai_n47_), .Y(mai_mai_n663_));
  AOI210     m0635(.A0(mai_mai_n1365_), .A1(mai_mai_n663_), .B0(mai_mai_n662_), .Y(mai_mai_n664_));
  NA4        m0636(.A(mai_mai_n664_), .B(mai_mai_n659_), .C(mai_mai_n658_), .D(mai_mai_n656_), .Y(mai_mai_n665_));
  NA2        m0637(.A(mai_mai_n320_), .B(mai_mai_n135_), .Y(mai_mai_n666_));
  NA2        m0638(.A(mai_mai_n126_), .B(mai_mai_n47_), .Y(mai_mai_n667_));
  AOI220     m0639(.A0(mai_mai_n667_), .A1(mai_mai_n519_), .B0(mai_mai_n351_), .B1(mai_mai_n107_), .Y(mai_mai_n668_));
  OA220      m0640(.A0(mai_mai_n668_), .A1(mai_mai_n540_), .B0(mai_mai_n349_), .B1(mai_mai_n105_), .Y(mai_mai_n669_));
  NA2        m0641(.A(mai_mai_n666_), .B(mai_mai_n669_), .Y(mai_mai_n670_));
  NO3        m0642(.A(mai_mai_n393_), .B(mai_mai_n188_), .C(mai_mai_n187_), .Y(mai_mai_n671_));
  NA2        m0643(.A(mai_mai_n671_), .B(mai_mai_n224_), .Y(mai_mai_n672_));
  NA3        m0644(.A(mai_mai_n672_), .B(mai_mai_n250_), .C(j), .Y(mai_mai_n673_));
  NO3        m0645(.A(mai_mai_n451_), .B(mai_mai_n169_), .C(i), .Y(mai_mai_n674_));
  NA2        m0646(.A(mai_mai_n455_), .B(mai_mai_n78_), .Y(mai_mai_n675_));
  NO4        m0647(.A(mai_mai_n516_), .B(mai_mai_n675_), .C(mai_mai_n125_), .D(mai_mai_n208_), .Y(mai_mai_n676_));
  INV        m0648(.A(mai_mai_n676_), .Y(mai_mai_n677_));
  NA4        m0649(.A(mai_mai_n677_), .B(mai_mai_n673_), .C(mai_mai_n501_), .D(mai_mai_n391_), .Y(mai_mai_n678_));
  NO4        m0650(.A(mai_mai_n678_), .B(mai_mai_n670_), .C(mai_mai_n665_), .D(mai_mai_n652_), .Y(mai_mai_n679_));
  NA4        m0651(.A(mai_mai_n679_), .B(mai_mai_n644_), .C(mai_mai_n599_), .D(mai_mai_n570_), .Y(mai08));
  NO2        m0652(.A(k), .B(h), .Y(mai_mai_n681_));
  AO210      m0653(.A0(mai_mai_n248_), .A1(mai_mai_n440_), .B0(mai_mai_n681_), .Y(mai_mai_n682_));
  NO2        m0654(.A(mai_mai_n682_), .B(mai_mai_n291_), .Y(mai_mai_n683_));
  NA2        m0655(.A(mai_mai_n608_), .B(mai_mai_n78_), .Y(mai_mai_n684_));
  NA2        m0656(.A(mai_mai_n684_), .B(mai_mai_n451_), .Y(mai_mai_n685_));
  AOI210     m0657(.A0(mai_mai_n685_), .A1(mai_mai_n683_), .B0(mai_mai_n476_), .Y(mai_mai_n686_));
  NO2        m0658(.A(n), .B(mai_mai_n54_), .Y(mai_mai_n687_));
  NO4        m0659(.A(mai_mai_n368_), .B(mai_mai_n106_), .C(j), .D(mai_mai_n209_), .Y(mai_mai_n688_));
  OAI210     m0660(.A0(mai_mai_n566_), .A1(mai_mai_n78_), .B0(mai_mai_n226_), .Y(mai_mai_n689_));
  AOI220     m0661(.A0(mai_mai_n689_), .A1(mai_mai_n339_), .B0(mai_mai_n688_), .B1(mai_mai_n687_), .Y(mai_mai_n690_));
  AOI210     m0662(.A0(mai_mai_n566_), .A1(mai_mai_n152_), .B0(mai_mai_n78_), .Y(mai_mai_n691_));
  NA4        m0663(.A(mai_mai_n211_), .B(mai_mai_n135_), .C(mai_mai_n44_), .D(h), .Y(mai_mai_n692_));
  NA4        m0664(.A(l), .B(mai_mai_n102_), .C(mai_mai_n69_), .D(mai_mai_n209_), .Y(mai_mai_n693_));
  OAI210     m0665(.A0(mai_mai_n692_), .A1(g), .B0(mai_mai_n693_), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n694_), .B(mai_mai_n691_), .Y(mai_mai_n695_));
  NA4        m0667(.A(mai_mai_n695_), .B(mai_mai_n690_), .C(mai_mai_n686_), .D(mai_mai_n341_), .Y(mai_mai_n696_));
  AN2        m0668(.A(mai_mai_n524_), .B(mai_mai_n90_), .Y(mai_mai_n697_));
  NO4        m0669(.A(mai_mai_n169_), .B(mai_mai_n381_), .C(mai_mai_n106_), .D(g), .Y(mai_mai_n698_));
  AOI210     m0670(.A0(mai_mai_n698_), .A1(mai_mai_n689_), .B0(mai_mai_n508_), .Y(mai_mai_n699_));
  NO2        m0671(.A(mai_mai_n37_), .B(mai_mai_n208_), .Y(mai_mai_n700_));
  AOI220     m0672(.A0(mai_mai_n609_), .A1(mai_mai_n338_), .B0(mai_mai_n700_), .B1(mai_mai_n555_), .Y(mai_mai_n701_));
  NAi31      m0673(.An(mai_mai_n697_), .B(mai_mai_n701_), .C(mai_mai_n699_), .Y(mai_mai_n702_));
  NO2        m0674(.A(mai_mai_n1370_), .B(mai_mai_n34_), .Y(mai_mai_n703_));
  NO2        m0675(.A(mai_mai_n470_), .B(mai_mai_n126_), .Y(mai_mai_n704_));
  AOI210     m0676(.A0(mai_mai_n704_), .A1(mai_mai_n45_), .B0(mai_mai_n703_), .Y(mai_mai_n705_));
  NO3        m0677(.A(mai_mai_n309_), .B(mai_mai_n125_), .C(mai_mai_n40_), .Y(mai_mai_n706_));
  NAi21      m0678(.An(mai_mai_n706_), .B(mai_mai_n693_), .Y(mai_mai_n707_));
  NA2        m0679(.A(mai_mai_n682_), .B(mai_mai_n130_), .Y(mai_mai_n708_));
  AOI220     m0680(.A0(mai_mai_n708_), .A1(mai_mai_n392_), .B0(mai_mai_n707_), .B1(mai_mai_n71_), .Y(mai_mai_n709_));
  OAI210     m0681(.A0(mai_mai_n705_), .A1(mai_mai_n81_), .B0(mai_mai_n709_), .Y(mai_mai_n710_));
  NA2        m0682(.A(mai_mai_n351_), .B(mai_mai_n42_), .Y(mai_mai_n711_));
  NA3        m0683(.A(mai_mai_n672_), .B(mai_mai_n326_), .C(mai_mai_n373_), .Y(mai_mai_n712_));
  NA2        m0684(.A(l), .B(mai_mai_n216_), .Y(mai_mai_n713_));
  NO2        m0685(.A(mai_mai_n713_), .B(mai_mai_n319_), .Y(mai_mai_n714_));
  AOI210     m0686(.A0(mai_mai_n714_), .A1(i), .B0(mai_mai_n475_), .Y(mai_mai_n715_));
  NA3        m0687(.A(m), .B(l), .C(k), .Y(mai_mai_n716_));
  AOI210     m0688(.A0(mai_mai_n649_), .A1(mai_mai_n647_), .B0(mai_mai_n716_), .Y(mai_mai_n717_));
  NO2        m0689(.A(mai_mai_n526_), .B(mai_mai_n266_), .Y(mai_mai_n718_));
  NOi21      m0690(.An(mai_mai_n718_), .B(mai_mai_n520_), .Y(mai_mai_n719_));
  NA4        m0691(.A(mai_mai_n107_), .B(l), .C(k), .D(mai_mai_n81_), .Y(mai_mai_n720_));
  NA3        m0692(.A(mai_mai_n114_), .B(mai_mai_n401_), .C(i), .Y(mai_mai_n721_));
  NO2        m0693(.A(mai_mai_n721_), .B(mai_mai_n720_), .Y(mai_mai_n722_));
  NO3        m0694(.A(mai_mai_n722_), .B(mai_mai_n719_), .C(mai_mai_n717_), .Y(mai_mai_n723_));
  NA4        m0695(.A(mai_mai_n723_), .B(mai_mai_n715_), .C(mai_mai_n712_), .D(mai_mai_n711_), .Y(mai_mai_n724_));
  NO4        m0696(.A(mai_mai_n724_), .B(mai_mai_n710_), .C(mai_mai_n702_), .D(mai_mai_n696_), .Y(mai_mai_n725_));
  NA2        m0697(.A(mai_mai_n609_), .B(mai_mai_n382_), .Y(mai_mai_n726_));
  NA2        m0698(.A(mai_mai_n624_), .B(g), .Y(mai_mai_n727_));
  AO210      m0699(.A0(mai_mai_n727_), .A1(mai_mai_n579_), .B0(mai_mai_n528_), .Y(mai_mai_n728_));
  NO3        m0700(.A(mai_mai_n386_), .B(mai_mai_n514_), .C(h), .Y(mai_mai_n729_));
  AOI210     m0701(.A0(mai_mai_n729_), .A1(mai_mai_n107_), .B0(mai_mai_n487_), .Y(mai_mai_n730_));
  NA4        m0702(.A(mai_mai_n730_), .B(mai_mai_n728_), .C(mai_mai_n726_), .D(mai_mai_n247_), .Y(mai_mai_n731_));
  NA2        m0703(.A(l), .B(mai_mai_n69_), .Y(mai_mai_n732_));
  NO4        m0704(.A(mai_mai_n671_), .B(mai_mai_n169_), .C(n), .D(i), .Y(mai_mai_n733_));
  NOi21      m0705(.An(h), .B(j), .Y(mai_mai_n734_));
  NA2        m0706(.A(mai_mai_n734_), .B(f), .Y(mai_mai_n735_));
  NO2        m0707(.A(mai_mai_n735_), .B(mai_mai_n241_), .Y(mai_mai_n736_));
  NO3        m0708(.A(mai_mai_n736_), .B(mai_mai_n733_), .C(mai_mai_n674_), .Y(mai_mai_n737_));
  OAI210     m0709(.A0(mai_mai_n737_), .A1(mai_mai_n732_), .B0(mai_mai_n581_), .Y(mai_mai_n738_));
  AOI210     m0710(.A0(mai_mai_n731_), .A1(l), .B0(mai_mai_n738_), .Y(mai_mai_n739_));
  NO2        m0711(.A(j), .B(i), .Y(mai_mai_n740_));
  NA3        m0712(.A(mai_mai_n740_), .B(mai_mai_n74_), .C(l), .Y(mai_mai_n741_));
  NA2        m0713(.A(mai_mai_n740_), .B(mai_mai_n32_), .Y(mai_mai_n742_));
  NA2        m0714(.A(mai_mai_n410_), .B(mai_mai_n114_), .Y(mai_mai_n743_));
  OA220      m0715(.A0(mai_mai_n743_), .A1(mai_mai_n742_), .B0(mai_mai_n741_), .B1(mai_mai_n577_), .Y(mai_mai_n744_));
  NO3        m0716(.A(mai_mai_n147_), .B(mai_mai_n47_), .C(mai_mai_n104_), .Y(mai_mai_n745_));
  NO3        m0717(.A(mai_mai_n532_), .B(mai_mai_n145_), .C(mai_mai_n69_), .Y(mai_mai_n746_));
  NO3        m0718(.A(mai_mai_n470_), .B(mai_mai_n428_), .C(j), .Y(mai_mai_n747_));
  OAI210     m0719(.A0(mai_mai_n746_), .A1(mai_mai_n745_), .B0(mai_mai_n747_), .Y(mai_mai_n748_));
  OAI210     m0720(.A0(mai_mai_n727_), .A1(mai_mai_n58_), .B0(mai_mai_n748_), .Y(mai_mai_n749_));
  NA2        m0721(.A(k), .B(j), .Y(mai_mai_n750_));
  NO3        m0722(.A(mai_mai_n291_), .B(mai_mai_n750_), .C(mai_mai_n39_), .Y(mai_mai_n751_));
  AOI210     m0723(.A0(mai_mai_n519_), .A1(n), .B0(mai_mai_n542_), .Y(mai_mai_n752_));
  NA2        m0724(.A(mai_mai_n752_), .B(mai_mai_n544_), .Y(mai_mai_n753_));
  AN3        m0725(.A(mai_mai_n753_), .B(mai_mai_n751_), .C(mai_mai_n92_), .Y(mai_mai_n754_));
  NO3        m0726(.A(mai_mai_n169_), .B(mai_mai_n381_), .C(mai_mai_n106_), .Y(mai_mai_n755_));
  AOI220     m0727(.A0(mai_mai_n755_), .A1(mai_mai_n242_), .B0(mai_mai_n602_), .B1(mai_mai_n301_), .Y(mai_mai_n756_));
  NAi31      m0728(.An(mai_mai_n595_), .B(mai_mai_n87_), .C(mai_mai_n78_), .Y(mai_mai_n757_));
  NA2        m0729(.A(mai_mai_n757_), .B(mai_mai_n756_), .Y(mai_mai_n758_));
  NO2        m0730(.A(mai_mai_n291_), .B(mai_mai_n130_), .Y(mai_mai_n759_));
  AOI220     m0731(.A0(mai_mai_n759_), .A1(mai_mai_n609_), .B0(mai_mai_n706_), .B1(mai_mai_n691_), .Y(mai_mai_n760_));
  NO2        m0732(.A(mai_mai_n716_), .B(mai_mai_n85_), .Y(mai_mai_n761_));
  NA2        m0733(.A(mai_mai_n761_), .B(mai_mai_n576_), .Y(mai_mai_n762_));
  NO2        m0734(.A(mai_mai_n578_), .B(mai_mai_n111_), .Y(mai_mai_n763_));
  OAI210     m0735(.A0(mai_mai_n763_), .A1(mai_mai_n747_), .B0(mai_mai_n663_), .Y(mai_mai_n764_));
  NA3        m0736(.A(mai_mai_n764_), .B(mai_mai_n762_), .C(mai_mai_n760_), .Y(mai_mai_n765_));
  OR4        m0737(.A(mai_mai_n765_), .B(mai_mai_n758_), .C(mai_mai_n754_), .D(mai_mai_n749_), .Y(mai_mai_n766_));
  NA3        m0738(.A(mai_mai_n752_), .B(mai_mai_n544_), .C(mai_mai_n543_), .Y(mai_mai_n767_));
  NA4        m0739(.A(mai_mai_n767_), .B(mai_mai_n211_), .C(mai_mai_n440_), .D(mai_mai_n33_), .Y(mai_mai_n768_));
  NO4        m0740(.A(mai_mai_n470_), .B(mai_mai_n424_), .C(j), .D(f), .Y(mai_mai_n769_));
  OAI220     m0741(.A0(mai_mai_n692_), .A1(mai_mai_n684_), .B0(mai_mai_n324_), .B1(mai_mai_n37_), .Y(mai_mai_n770_));
  AOI210     m0742(.A0(mai_mai_n769_), .A1(mai_mai_n254_), .B0(mai_mai_n770_), .Y(mai_mai_n771_));
  NA3        m0743(.A(mai_mai_n535_), .B(mai_mai_n285_), .C(h), .Y(mai_mai_n772_));
  NOi21      m0744(.An(mai_mai_n663_), .B(mai_mai_n772_), .Y(mai_mai_n773_));
  NO2        m0745(.A(mai_mai_n86_), .B(mai_mai_n1368_), .Y(mai_mai_n774_));
  OAI220     m0746(.A0(mai_mai_n772_), .A1(mai_mai_n593_), .B0(mai_mai_n741_), .B1(mai_mai_n67_), .Y(mai_mai_n775_));
  AOI210     m0747(.A0(mai_mai_n774_), .A1(mai_mai_n630_), .B0(mai_mai_n775_), .Y(mai_mai_n776_));
  NAi41      m0748(.An(mai_mai_n773_), .B(mai_mai_n776_), .C(mai_mai_n771_), .D(mai_mai_n768_), .Y(mai_mai_n777_));
  OR2        m0749(.A(mai_mai_n761_), .B(mai_mai_n90_), .Y(mai_mai_n778_));
  AOI220     m0750(.A0(mai_mai_n778_), .A1(mai_mai_n232_), .B0(mai_mai_n747_), .B1(mai_mai_n622_), .Y(mai_mai_n779_));
  NO2        m0751(.A(mai_mai_n648_), .B(mai_mai_n69_), .Y(mai_mai_n780_));
  AOI210     m0752(.A0(mai_mai_n769_), .A1(mai_mai_n780_), .B0(mai_mai_n328_), .Y(mai_mai_n781_));
  OAI210     m0753(.A0(mai_mai_n716_), .A1(mai_mai_n646_), .B0(mai_mai_n507_), .Y(mai_mai_n782_));
  NA3        m0754(.A(mai_mai_n245_), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n783_));
  NO2        m0755(.A(mai_mai_n772_), .B(mai_mai_n474_), .Y(mai_mai_n784_));
  AOI210     m0756(.A0(mai_mai_n78_), .A1(mai_mai_n782_), .B0(mai_mai_n784_), .Y(mai_mai_n785_));
  NA3        m0757(.A(mai_mai_n785_), .B(mai_mai_n781_), .C(mai_mai_n779_), .Y(mai_mai_n786_));
  NOi41      m0758(.An(mai_mai_n744_), .B(mai_mai_n786_), .C(mai_mai_n777_), .D(mai_mai_n766_), .Y(mai_mai_n787_));
  OR3        m0759(.A(mai_mai_n692_), .B(mai_mai_n226_), .C(g), .Y(mai_mai_n788_));
  NO3        m0760(.A(mai_mai_n334_), .B(mai_mai_n293_), .C(mai_mai_n106_), .Y(mai_mai_n789_));
  NA2        m0761(.A(mai_mai_n789_), .B(mai_mai_n753_), .Y(mai_mai_n790_));
  NO3        m0762(.A(mai_mai_n1367_), .B(mai_mai_n742_), .C(mai_mai_n272_), .Y(mai_mai_n791_));
  NO3        m0763(.A(mai_mai_n514_), .B(mai_mai_n88_), .C(h), .Y(mai_mai_n792_));
  AOI210     m0764(.A0(mai_mai_n792_), .A1(mai_mai_n687_), .B0(mai_mai_n791_), .Y(mai_mai_n793_));
  NA4        m0765(.A(mai_mai_n793_), .B(mai_mai_n790_), .C(mai_mai_n788_), .D(mai_mai_n394_), .Y(mai_mai_n794_));
  OR2        m0766(.A(mai_mai_n646_), .B(mai_mai_n86_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n1364_), .B(n), .Y(mai_mai_n796_));
  OAI220     m0768(.A0(n), .A1(mai_mai_n795_), .B0(mai_mai_n772_), .B1(mai_mai_n591_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n543_), .B(mai_mai_n78_), .Y(mai_mai_n798_));
  NO2        m0770(.A(mai_mai_n319_), .B(mai_mai_n111_), .Y(mai_mai_n799_));
  NOi21      m0771(.An(mai_mai_n799_), .B(mai_mai_n156_), .Y(mai_mai_n800_));
  AOI210     m0772(.A0(mai_mai_n789_), .A1(mai_mai_n798_), .B0(mai_mai_n800_), .Y(mai_mai_n801_));
  OAI210     m0773(.A0(mai_mai_n692_), .A1(mai_mai_n383_), .B0(mai_mai_n801_), .Y(mai_mai_n802_));
  NO2        m0774(.A(mai_mai_n671_), .B(n), .Y(mai_mai_n803_));
  AOI220     m0775(.A0(mai_mai_n759_), .A1(mai_mai_n653_), .B0(mai_mai_n803_), .B1(mai_mai_n683_), .Y(mai_mai_n804_));
  NO2        m0776(.A(mai_mai_n315_), .B(mai_mai_n231_), .Y(mai_mai_n805_));
  OAI210     m0777(.A0(mai_mai_n90_), .A1(mai_mai_n87_), .B0(mai_mai_n805_), .Y(mai_mai_n806_));
  NA2        m0778(.A(mai_mai_n114_), .B(mai_mai_n78_), .Y(mai_mai_n807_));
  AOI210     m0779(.A0(mai_mai_n414_), .A1(mai_mai_n407_), .B0(mai_mai_n807_), .Y(mai_mai_n808_));
  NAi21      m0780(.An(mai_mai_n808_), .B(mai_mai_n806_), .Y(mai_mai_n809_));
  NA2        m0781(.A(mai_mai_n714_), .B(mai_mai_n33_), .Y(mai_mai_n810_));
  NAi21      m0782(.An(mai_mai_n720_), .B(mai_mai_n425_), .Y(mai_mai_n811_));
  NO2        m0783(.A(mai_mai_n266_), .B(i), .Y(mai_mai_n812_));
  NA2        m0784(.A(mai_mai_n698_), .B(mai_mai_n340_), .Y(mai_mai_n813_));
  OAI210     m0785(.A0(mai_mai_n584_), .A1(mai_mai_n583_), .B0(mai_mai_n352_), .Y(mai_mai_n814_));
  AN3        m0786(.A(mai_mai_n814_), .B(mai_mai_n813_), .C(mai_mai_n811_), .Y(mai_mai_n815_));
  NAi41      m0787(.An(mai_mai_n809_), .B(mai_mai_n815_), .C(mai_mai_n810_), .D(mai_mai_n804_), .Y(mai_mai_n816_));
  NO4        m0788(.A(mai_mai_n816_), .B(mai_mai_n802_), .C(mai_mai_n797_), .D(mai_mai_n794_), .Y(mai_mai_n817_));
  NA4        m0789(.A(mai_mai_n817_), .B(mai_mai_n787_), .C(mai_mai_n739_), .D(mai_mai_n725_), .Y(mai09));
  INV        m0790(.A(mai_mai_n115_), .Y(mai_mai_n819_));
  NA2        m0791(.A(f), .B(e), .Y(mai_mai_n820_));
  NA2        m0792(.A(l), .B(g), .Y(mai_mai_n821_));
  NO2        m0793(.A(g), .B(mai_mai_n458_), .Y(mai_mai_n822_));
  AOI210     m0794(.A0(mai_mai_n822_), .A1(mai_mai_n821_), .B0(mai_mai_n820_), .Y(mai_mai_n823_));
  NA2        m0795(.A(mai_mai_n434_), .B(e), .Y(mai_mai_n824_));
  NO2        m0796(.A(mai_mai_n824_), .B(mai_mai_n498_), .Y(mai_mai_n825_));
  AOI210     m0797(.A0(mai_mai_n823_), .A1(mai_mai_n819_), .B0(mai_mai_n825_), .Y(mai_mai_n826_));
  NA3        m0798(.A(m), .B(l), .C(i), .Y(mai_mai_n827_));
  OAI220     m0799(.A0(mai_mai_n578_), .A1(mai_mai_n827_), .B0(mai_mai_n343_), .B1(mai_mai_n515_), .Y(mai_mai_n828_));
  NA4        m0800(.A(mai_mai_n82_), .B(mai_mai_n81_), .C(g), .D(f), .Y(mai_mai_n829_));
  NAi31      m0801(.An(mai_mai_n828_), .B(mai_mai_n829_), .C(mai_mai_n429_), .Y(mai_mai_n830_));
  NA3        m0802(.A(mai_mai_n795_), .B(mai_mai_n557_), .C(mai_mai_n507_), .Y(mai_mai_n831_));
  OA210      m0803(.A0(mai_mai_n831_), .A1(n), .B0(mai_mai_n796_), .Y(mai_mai_n832_));
  INV        m0804(.A(mai_mai_n331_), .Y(mai_mai_n833_));
  AOI210     m0805(.A0(m), .A1(m), .B0(mai_mai_n587_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n783_), .B(mai_mai_n324_), .Y(mai_mai_n835_));
  NA2        m0807(.A(mai_mai_n335_), .B(m), .Y(mai_mai_n836_));
  OAI210     m0808(.A0(mai_mai_n199_), .A1(mai_mai_n208_), .B0(mai_mai_n836_), .Y(mai_mai_n837_));
  AOI220     m0809(.A0(mai_mai_n837_), .A1(mai_mai_n835_), .B0(mai_mai_n834_), .B1(mai_mai_n833_), .Y(mai_mai_n838_));
  NA3        m0810(.A(mai_mai_n1361_), .B(mai_mai_n185_), .C(mai_mai_n30_), .Y(mai_mai_n839_));
  NA4        m0811(.A(mai_mai_n839_), .B(mai_mai_n838_), .C(mai_mai_n610_), .D(mai_mai_n76_), .Y(mai_mai_n840_));
  NO2        m0812(.A(mai_mai_n574_), .B(mai_mai_n483_), .Y(mai_mai_n841_));
  NA2        m0813(.A(mai_mai_n841_), .B(mai_mai_n185_), .Y(mai_mai_n842_));
  NA2        m0814(.A(f), .B(m), .Y(mai_mai_n843_));
  NO2        m0815(.A(mai_mai_n843_), .B(mai_mai_n50_), .Y(mai_mai_n844_));
  NOi32      m0816(.An(g), .Bn(f), .C(d), .Y(mai_mai_n845_));
  NA4        m0817(.A(mai_mai_n845_), .B(mai_mai_n592_), .C(a), .D(m), .Y(mai_mai_n846_));
  INV        m0818(.A(mai_mai_n846_), .Y(mai_mai_n847_));
  AOI210     m0819(.A0(mai_mai_n844_), .A1(mai_mai_n533_), .B0(mai_mai_n847_), .Y(mai_mai_n848_));
  AN2        m0820(.A(f), .B(d), .Y(mai_mai_n849_));
  NA3        m0821(.A(a), .B(mai_mai_n849_), .C(mai_mai_n78_), .Y(mai_mai_n850_));
  NO3        m0822(.A(mai_mai_n850_), .B(mai_mai_n69_), .C(mai_mai_n209_), .Y(mai_mai_n851_));
  NO2        m0823(.A(mai_mai_n280_), .B(mai_mai_n53_), .Y(mai_mai_n852_));
  OAI210     m0824(.A0(mai_mai_n852_), .A1(k), .B0(mai_mai_n851_), .Y(mai_mai_n853_));
  NAi41      m0825(.An(mai_mai_n473_), .B(mai_mai_n853_), .C(mai_mai_n848_), .D(mai_mai_n842_), .Y(mai_mai_n854_));
  NO3        m0826(.A(mai_mai_n126_), .B(mai_mai_n319_), .C(mai_mai_n148_), .Y(mai_mai_n855_));
  NO2        m0827(.A(mai_mai_n640_), .B(mai_mai_n319_), .Y(mai_mai_n856_));
  AN2        m0828(.A(mai_mai_n856_), .B(i), .Y(mai_mai_n857_));
  NO3        m0829(.A(mai_mai_n857_), .B(mai_mai_n855_), .C(mai_mai_n228_), .Y(mai_mai_n858_));
  NA2        m0830(.A(a), .B(mai_mai_n78_), .Y(mai_mai_n859_));
  OAI220     m0831(.A0(mai_mai_n836_), .A1(mai_mai_n859_), .B0(mai_mai_n783_), .B1(mai_mai_n429_), .Y(mai_mai_n860_));
  NA3        m0832(.A(mai_mai_n155_), .B(mai_mai_n102_), .C(g), .Y(mai_mai_n861_));
  OAI220     m0833(.A0(mai_mai_n850_), .A1(mai_mai_n419_), .B0(mai_mai_n331_), .B1(mai_mai_n861_), .Y(mai_mai_n862_));
  NOi41      m0834(.An(mai_mai_n219_), .B(mai_mai_n862_), .C(mai_mai_n860_), .D(mai_mai_n299_), .Y(mai_mai_n863_));
  NA2        m0835(.A(c), .B(mai_mai_n110_), .Y(mai_mai_n864_));
  NO2        m0836(.A(mai_mai_n864_), .B(mai_mai_n398_), .Y(mai_mai_n865_));
  NA3        m0837(.A(mai_mai_n865_), .B(mai_mai_n496_), .C(f), .Y(mai_mai_n866_));
  OR2        m0838(.A(mai_mai_n646_), .B(mai_mai_n529_), .Y(mai_mai_n867_));
  NA4        m0839(.A(mai_mai_n867_), .B(mai_mai_n866_), .C(mai_mai_n863_), .D(mai_mai_n858_), .Y(mai_mai_n868_));
  NO4        m0840(.A(mai_mai_n868_), .B(mai_mai_n854_), .C(mai_mai_n840_), .D(mai_mai_n832_), .Y(mai_mai_n869_));
  OR2        m0841(.A(mai_mai_n850_), .B(mai_mai_n69_), .Y(mai_mai_n870_));
  OAI210     m0842(.A0(j), .A1(l), .B0(g), .Y(mai_mai_n871_));
  AOI210     m0843(.A0(mai_mai_n871_), .A1(mai_mai_n286_), .B0(mai_mai_n870_), .Y(mai_mai_n872_));
  AOI210     m0844(.A0(mai_mai_n783_), .A1(mai_mai_n324_), .B0(mai_mai_n829_), .Y(mai_mai_n873_));
  NO2        m0845(.A(mai_mai_n130_), .B(mai_mai_n126_), .Y(mai_mai_n874_));
  NO2        m0846(.A(mai_mai_n224_), .B(mai_mai_n220_), .Y(mai_mai_n875_));
  AOI220     m0847(.A0(mai_mai_n875_), .A1(mai_mai_n221_), .B0(mai_mai_n297_), .B1(mai_mai_n874_), .Y(mai_mai_n876_));
  NO2        m0848(.A(mai_mai_n419_), .B(mai_mai_n820_), .Y(mai_mai_n877_));
  NA2        m0849(.A(mai_mai_n877_), .B(mai_mai_n549_), .Y(mai_mai_n878_));
  NA2        m0850(.A(mai_mai_n878_), .B(mai_mai_n876_), .Y(mai_mai_n879_));
  NA2        m0851(.A(e), .B(d), .Y(mai_mai_n880_));
  OAI220     m0852(.A0(mai_mai_n880_), .A1(c), .B0(mai_mai_n315_), .B1(d), .Y(mai_mai_n881_));
  NA3        m0853(.A(mai_mai_n881_), .B(mai_mai_n444_), .C(mai_mai_n494_), .Y(mai_mai_n882_));
  AOI210     m0854(.A0(mai_mai_n502_), .A1(mai_mai_n176_), .B0(mai_mai_n224_), .Y(mai_mai_n883_));
  AOI210     m0855(.A0(mai_mai_n609_), .A1(mai_mai_n338_), .B0(mai_mai_n883_), .Y(mai_mai_n884_));
  NA3        m0856(.A(mai_mai_n851_), .B(j), .C(mai_mai_n53_), .Y(mai_mai_n885_));
  NA3        m0857(.A(mai_mai_n162_), .B(mai_mai_n79_), .C(mai_mai_n33_), .Y(mai_mai_n886_));
  NA4        m0858(.A(mai_mai_n886_), .B(mai_mai_n885_), .C(mai_mai_n884_), .D(mai_mai_n882_), .Y(mai_mai_n887_));
  NO4        m0859(.A(mai_mai_n887_), .B(mai_mai_n879_), .C(mai_mai_n873_), .D(mai_mai_n872_), .Y(mai_mai_n888_));
  AO210      m0860(.A0(mai_mai_n331_), .A1(mai_mai_n684_), .B0(mai_mai_n212_), .Y(mai_mai_n889_));
  AOI220     m0861(.A0(h), .A1(mai_mai_n856_), .B0(mai_mai_n600_), .B1(mai_mai_n608_), .Y(mai_mai_n890_));
  OAI210     m0862(.A0(mai_mai_n824_), .A1(mai_mai_n166_), .B0(mai_mai_n890_), .Y(mai_mai_n891_));
  INV        m0863(.A(mai_mai_n845_), .Y(mai_mai_n892_));
  NO2        m0864(.A(mai_mai_n892_), .B(mai_mai_n593_), .Y(mai_mai_n893_));
  INV        m0865(.A(mai_mai_n846_), .Y(mai_mai_n894_));
  AO210      m0866(.A0(mai_mai_n835_), .A1(mai_mai_n828_), .B0(mai_mai_n894_), .Y(mai_mai_n895_));
  NOi31      m0867(.An(mai_mai_n533_), .B(mai_mai_n843_), .C(mai_mai_n286_), .Y(mai_mai_n896_));
  NO4        m0868(.A(mai_mai_n896_), .B(mai_mai_n895_), .C(mai_mai_n893_), .D(mai_mai_n891_), .Y(mai_mai_n897_));
  AO220      m0869(.A0(mai_mai_n444_), .A1(mai_mai_n734_), .B0(mai_mai_n171_), .B1(f), .Y(mai_mai_n898_));
  OAI210     m0870(.A0(mai_mai_n898_), .A1(mai_mai_n447_), .B0(mai_mai_n881_), .Y(mai_mai_n899_));
  NO2        m0871(.A(mai_mai_n428_), .B(mai_mai_n65_), .Y(mai_mai_n900_));
  OAI210     m0872(.A0(mai_mai_n831_), .A1(mai_mai_n900_), .B0(mai_mai_n687_), .Y(mai_mai_n901_));
  AN4        m0873(.A(mai_mai_n901_), .B(mai_mai_n899_), .C(mai_mai_n897_), .D(mai_mai_n889_), .Y(mai_mai_n902_));
  NA4        m0874(.A(mai_mai_n902_), .B(mai_mai_n888_), .C(mai_mai_n869_), .D(mai_mai_n826_), .Y(mai12));
  NO2        m0875(.A(mai_mai_n442_), .B(c), .Y(mai_mai_n904_));
  NO4        m0876(.A(mai_mai_n433_), .B(mai_mai_n248_), .C(mai_mai_n571_), .D(mai_mai_n209_), .Y(mai_mai_n905_));
  NA2        m0877(.A(mai_mai_n905_), .B(mai_mai_n904_), .Y(mai_mai_n906_));
  NA2        m0878(.A(mai_mai_n533_), .B(mai_mai_n900_), .Y(mai_mai_n907_));
  NO3        m0879(.A(mai_mai_n442_), .B(mai_mai_n78_), .C(mai_mai_n110_), .Y(mai_mai_n908_));
  NO2        m0880(.A(m), .B(mai_mai_n343_), .Y(mai_mai_n909_));
  NO2        m0881(.A(mai_mai_n646_), .B(mai_mai_n368_), .Y(mai_mai_n910_));
  AOI220     m0882(.A0(mai_mai_n910_), .A1(mai_mai_n531_), .B0(mai_mai_n909_), .B1(mai_mai_n908_), .Y(mai_mai_n911_));
  NA4        m0883(.A(mai_mai_n911_), .B(mai_mai_n907_), .C(mai_mai_n906_), .D(mai_mai_n432_), .Y(mai_mai_n912_));
  AOI210     m0884(.A0(mai_mai_n227_), .A1(mai_mai_n330_), .B0(mai_mai_n196_), .Y(mai_mai_n913_));
  OR2        m0885(.A(mai_mai_n913_), .B(mai_mai_n905_), .Y(mai_mai_n914_));
  AOI210     m0886(.A0(mai_mai_n327_), .A1(mai_mai_n379_), .B0(mai_mai_n209_), .Y(mai_mai_n915_));
  OAI210     m0887(.A0(mai_mai_n915_), .A1(mai_mai_n914_), .B0(mai_mai_n393_), .Y(mai_mai_n916_));
  NO2        m0888(.A(mai_mai_n627_), .B(mai_mai_n257_), .Y(mai_mai_n917_));
  NO2        m0889(.A(mai_mai_n578_), .B(mai_mai_n827_), .Y(mai_mai_n918_));
  AOI220     m0890(.A0(mai_mai_n918_), .A1(mai_mai_n555_), .B0(mai_mai_n805_), .B1(mai_mai_n917_), .Y(mai_mai_n919_));
  NO2        m0891(.A(mai_mai_n147_), .B(mai_mai_n231_), .Y(mai_mai_n920_));
  NA3        m0892(.A(mai_mai_n920_), .B(mai_mai_n234_), .C(i), .Y(mai_mai_n921_));
  NA3        m0893(.A(mai_mai_n921_), .B(mai_mai_n919_), .C(mai_mai_n916_), .Y(mai_mai_n922_));
  OR2        m0894(.A(mai_mai_n316_), .B(mai_mai_n908_), .Y(mai_mai_n923_));
  NA2        m0895(.A(mai_mai_n923_), .B(mai_mai_n344_), .Y(mai_mai_n924_));
  NO3        m0896(.A(mai_mai_n126_), .B(mai_mai_n148_), .C(mai_mai_n209_), .Y(mai_mai_n925_));
  NA2        m0897(.A(mai_mai_n925_), .B(mai_mai_n519_), .Y(mai_mai_n926_));
  NA4        m0898(.A(mai_mai_n434_), .B(d), .C(mai_mai_n177_), .D(g), .Y(mai_mai_n927_));
  NA3        m0899(.A(mai_mai_n927_), .B(mai_mai_n926_), .C(mai_mai_n924_), .Y(mai_mai_n928_));
  NO3        m0900(.A(mai_mai_n651_), .B(mai_mai_n86_), .C(mai_mai_n44_), .Y(mai_mai_n929_));
  NO4        m0901(.A(mai_mai_n929_), .B(mai_mai_n928_), .C(mai_mai_n922_), .D(mai_mai_n912_), .Y(mai_mai_n930_));
  NO2        m0902(.A(mai_mai_n1363_), .B(mai_mai_n358_), .Y(mai_mai_n931_));
  NA2        m0903(.A(mai_mai_n575_), .B(mai_mai_n67_), .Y(mai_mai_n932_));
  NOi21      m0904(.An(mai_mai_n33_), .B(mai_mai_n640_), .Y(mai_mai_n933_));
  AOI220     m0905(.A0(mai_mai_n933_), .A1(c), .B0(mai_mai_n932_), .B1(mai_mai_n931_), .Y(mai_mai_n934_));
  OAI210     m0906(.A0(mai_mai_n246_), .A1(mai_mai_n44_), .B0(mai_mai_n934_), .Y(mai_mai_n935_));
  NA2        m0907(.A(mai_mai_n425_), .B(mai_mai_n259_), .Y(mai_mai_n936_));
  NO2        m0908(.A(mai_mai_n807_), .B(mai_mai_n83_), .Y(mai_mai_n937_));
  NAi31      m0909(.An(mai_mai_n937_), .B(mai_mai_n936_), .C(mai_mai_n313_), .Y(mai_mai_n938_));
  NO2        m0910(.A(mai_mai_n490_), .B(mai_mai_n293_), .Y(mai_mai_n939_));
  NO2        m0911(.A(mai_mai_n204_), .B(mai_mai_n140_), .Y(mai_mai_n940_));
  OAI210     m0912(.A0(mai_mai_n721_), .A1(n), .B0(mai_mai_n356_), .Y(mai_mai_n941_));
  NO4        m0913(.A(mai_mai_n941_), .B(mai_mai_n940_), .C(mai_mai_n938_), .D(mai_mai_n935_), .Y(mai_mai_n942_));
  NA2        m0914(.A(mai_mai_n338_), .B(g), .Y(mai_mai_n943_));
  NA2        m0915(.A(h), .B(i), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n45_), .B(i), .Y(mai_mai_n945_));
  OAI220     m0917(.A0(mai_mai_n945_), .A1(mai_mai_n1358_), .B0(mai_mai_n944_), .B1(mai_mai_n86_), .Y(mai_mai_n946_));
  AOI210     m0918(.A0(m), .A1(mai_mai_n36_), .B0(mai_mai_n946_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n140_), .B(mai_mai_n78_), .Y(mai_mai_n948_));
  OR2        m0920(.A(mai_mai_n948_), .B(mai_mai_n542_), .Y(mai_mai_n949_));
  AOI210     m0921(.A0(c), .A1(n), .B0(mai_mai_n949_), .Y(mai_mai_n950_));
  OAI220     m0922(.A0(mai_mai_n950_), .A1(mai_mai_n943_), .B0(mai_mai_n947_), .B1(mai_mai_n324_), .Y(mai_mai_n951_));
  NO2        m0923(.A(mai_mai_n646_), .B(mai_mai_n483_), .Y(mai_mai_n952_));
  NA3        m0924(.A(mai_mai_n335_), .B(j), .C(i), .Y(mai_mai_n953_));
  OAI220     m0925(.A0(mai_mai_n1356_), .A1(mai_mai_n952_), .B0(mai_mai_n663_), .B1(mai_mai_n746_), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n594_), .B(mai_mai_n107_), .Y(mai_mai_n955_));
  NA3        m0927(.A(j), .B(mai_mai_n74_), .C(i), .Y(mai_mai_n956_));
  OR2        m0928(.A(mai_mai_n956_), .B(mai_mai_n955_), .Y(mai_mai_n957_));
  NA3        m0929(.A(f), .B(mai_mai_n112_), .C(g), .Y(mai_mai_n958_));
  AOI210     m0930(.A0(mai_mai_n660_), .A1(mai_mai_n958_), .B0(m), .Y(mai_mai_n959_));
  OAI210     m0931(.A0(mai_mai_n959_), .A1(mai_mai_n909_), .B0(mai_mai_n316_), .Y(mai_mai_n960_));
  NA2        m0932(.A(mai_mai_n829_), .B(mai_mai_n429_), .Y(mai_mai_n961_));
  NA2        m0933(.A(mai_mai_n217_), .B(h), .Y(mai_mai_n962_));
  NA2        m0934(.A(mai_mai_n962_), .B(mai_mai_n956_), .Y(mai_mai_n963_));
  AOI220     m0935(.A0(mai_mai_n963_), .A1(mai_mai_n254_), .B0(mai_mai_n961_), .B1(mai_mai_n78_), .Y(mai_mai_n964_));
  NA4        m0936(.A(mai_mai_n964_), .B(mai_mai_n960_), .C(mai_mai_n957_), .D(mai_mai_n954_), .Y(mai_mai_n965_));
  NO2        m0937(.A(mai_mai_n368_), .B(mai_mai_n85_), .Y(mai_mai_n966_));
  OAI210     m0938(.A0(mai_mai_n966_), .A1(mai_mai_n917_), .B0(mai_mai_n232_), .Y(mai_mai_n967_));
  NA2        m0939(.A(mai_mai_n650_), .B(mai_mai_n82_), .Y(mai_mai_n968_));
  NO2        m0940(.A(mai_mai_n450_), .B(mai_mai_n209_), .Y(mai_mai_n969_));
  AOI220     m0941(.A0(mai_mai_n969_), .A1(mai_mai_n372_), .B0(mai_mai_n923_), .B1(mai_mai_n213_), .Y(mai_mai_n970_));
  AOI220     m0942(.A0(mai_mai_n910_), .A1(mai_mai_n920_), .B0(mai_mai_n576_), .B1(mai_mai_n84_), .Y(mai_mai_n971_));
  NA4        m0943(.A(mai_mai_n971_), .B(mai_mai_n970_), .C(mai_mai_n968_), .D(mai_mai_n967_), .Y(mai_mai_n972_));
  OAI210     m0944(.A0(mai_mai_n961_), .A1(mai_mai_n918_), .B0(mai_mai_n531_), .Y(mai_mai_n973_));
  AOI210     m0945(.A0(mai_mai_n409_), .A1(mai_mai_n402_), .B0(mai_mai_n807_), .Y(mai_mai_n974_));
  OAI210     m0946(.A0(mai_mai_n1363_), .A1(mai_mai_n358_), .B0(mai_mai_n103_), .Y(mai_mai_n975_));
  AOI210     m0947(.A0(mai_mai_n975_), .A1(mai_mai_n524_), .B0(mai_mai_n974_), .Y(mai_mai_n976_));
  NA2        m0948(.A(mai_mai_n959_), .B(mai_mai_n908_), .Y(mai_mai_n977_));
  NO2        m0949(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n978_));
  AOI220     m0950(.A0(mai_mai_n978_), .A1(mai_mai_n612_), .B0(mai_mai_n632_), .B1(mai_mai_n519_), .Y(mai_mai_n979_));
  NA4        m0951(.A(mai_mai_n979_), .B(mai_mai_n977_), .C(mai_mai_n976_), .D(mai_mai_n973_), .Y(mai_mai_n980_));
  NO4        m0952(.A(mai_mai_n980_), .B(mai_mai_n972_), .C(mai_mai_n965_), .D(mai_mai_n951_), .Y(mai_mai_n981_));
  NAi31      m0953(.An(mai_mai_n136_), .B(mai_mai_n410_), .C(n), .Y(mai_mai_n982_));
  NO2        m0954(.A(m), .B(mai_mai_n982_), .Y(mai_mai_n983_));
  NO3        m0955(.A(mai_mai_n266_), .B(mai_mai_n136_), .C(mai_mai_n398_), .Y(mai_mai_n984_));
  AOI210     m0956(.A0(mai_mai_n984_), .A1(mai_mai_n484_), .B0(mai_mai_n983_), .Y(mai_mai_n985_));
  NA2        m0957(.A(mai_mai_n476_), .B(i), .Y(mai_mai_n986_));
  NA2        m0958(.A(mai_mai_n986_), .B(mai_mai_n985_), .Y(mai_mai_n987_));
  NA2        m0959(.A(mai_mai_n224_), .B(mai_mai_n167_), .Y(mai_mai_n988_));
  NO3        m0960(.A(mai_mai_n301_), .B(mai_mai_n434_), .C(mai_mai_n171_), .Y(mai_mai_n989_));
  NOi31      m0961(.An(mai_mai_n988_), .B(mai_mai_n989_), .C(mai_mai_n209_), .Y(mai_mai_n990_));
  NAi21      m0962(.An(mai_mai_n543_), .B(mai_mai_n969_), .Y(mai_mai_n991_));
  NO3        m0963(.A(mai_mai_n428_), .B(k), .C(mai_mai_n69_), .Y(mai_mai_n992_));
  AOI220     m0964(.A0(mai_mai_n992_), .A1(mai_mai_n426_), .B0(mai_mai_n468_), .B1(g), .Y(mai_mai_n993_));
  NA2        m0965(.A(mai_mai_n993_), .B(mai_mai_n991_), .Y(mai_mai_n994_));
  OAI220     m0966(.A0(mai_mai_n982_), .A1(mai_mai_n227_), .B0(mai_mai_n953_), .B1(mai_mai_n591_), .Y(mai_mai_n995_));
  NO2        m0967(.A(mai_mai_n647_), .B(mai_mai_n368_), .Y(mai_mai_n996_));
  NA2        m0968(.A(mai_mai_n913_), .B(mai_mai_n904_), .Y(mai_mai_n997_));
  NA2        m0969(.A(mai_mai_n513_), .B(mai_mai_n369_), .Y(mai_mai_n998_));
  OAI220     m0970(.A0(mai_mai_n910_), .A1(mai_mai_n918_), .B0(mai_mai_n533_), .B1(mai_mai_n418_), .Y(mai_mai_n999_));
  NA4        m0971(.A(mai_mai_n999_), .B(mai_mai_n998_), .C(mai_mai_n997_), .D(mai_mai_n607_), .Y(mai_mai_n1000_));
  OAI210     m0972(.A0(mai_mai_n913_), .A1(mai_mai_n905_), .B0(mai_mai_n988_), .Y(mai_mai_n1001_));
  NA3        m0973(.A(c), .B(mai_mai_n471_), .C(mai_mai_n45_), .Y(mai_mai_n1002_));
  AOI210     m0974(.A0(mai_mai_n370_), .A1(mai_mai_n369_), .B0(mai_mai_n323_), .Y(mai_mai_n1003_));
  NA4        m0975(.A(mai_mai_n1003_), .B(mai_mai_n1002_), .C(mai_mai_n1001_), .D(mai_mai_n267_), .Y(mai_mai_n1004_));
  OR4        m0976(.A(mai_mai_n1004_), .B(mai_mai_n1000_), .C(mai_mai_n996_), .D(mai_mai_n995_), .Y(mai_mai_n1005_));
  NO4        m0977(.A(mai_mai_n1005_), .B(mai_mai_n994_), .C(mai_mai_n990_), .D(mai_mai_n987_), .Y(mai_mai_n1006_));
  NA4        m0978(.A(mai_mai_n1006_), .B(mai_mai_n981_), .C(mai_mai_n942_), .D(mai_mai_n930_), .Y(mai13));
  AN2        m0979(.A(c), .B(b), .Y(mai_mai_n1008_));
  NA3        m0980(.A(mai_mai_n245_), .B(mai_mai_n1008_), .C(m), .Y(mai_mai_n1009_));
  NA2        m0981(.A(mai_mai_n481_), .B(f), .Y(mai_mai_n1010_));
  NO4        m0982(.A(mai_mai_n1010_), .B(mai_mai_n1009_), .C(j), .D(k), .Y(mai_mai_n1011_));
  NO4        m0983(.A(mai_mai_n63_), .B(mai_mai_n1010_), .C(mai_mai_n944_), .D(a), .Y(mai_mai_n1012_));
  NAi32      m0984(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1013_));
  NA2        m0985(.A(mai_mai_n135_), .B(mai_mai_n44_), .Y(mai_mai_n1014_));
  NO4        m0986(.A(mai_mai_n1014_), .B(mai_mai_n1013_), .C(mai_mai_n578_), .D(mai_mai_n300_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(mai_mai_n401_), .B(mai_mai_n208_), .Y(mai_mai_n1016_));
  AN2        m0988(.A(d), .B(c), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n1017_), .B(mai_mai_n110_), .Y(mai_mai_n1018_));
  NO3        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1016_), .C(mai_mai_n172_), .Y(mai_mai_n1019_));
  NA2        m0991(.A(mai_mai_n481_), .B(c), .Y(mai_mai_n1020_));
  NO3        m0992(.A(mai_mai_n1014_), .B(mai_mai_n574_), .C(mai_mai_n300_), .Y(mai_mai_n1021_));
  OR2        m0993(.A(mai_mai_n1019_), .B(mai_mai_n1021_), .Y(mai_mai_n1022_));
  OR4        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1015_), .C(mai_mai_n1012_), .D(mai_mai_n1011_), .Y(mai_mai_n1023_));
  OR3        m0995(.A(mai_mai_n220_), .B(mai_mai_n172_), .C(mai_mai_n163_), .Y(mai_mai_n1024_));
  NO2        m0996(.A(mai_mai_n1024_), .B(mai_mai_n142_), .Y(mai_mai_n1025_));
  NO2        m0997(.A(mai_mai_n1020_), .B(mai_mai_n300_), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n615_), .B(mai_mai_n1359_), .Y(mai_mai_n1027_));
  NOi21      m0999(.An(mai_mai_n1026_), .B(mai_mai_n1027_), .Y(mai_mai_n1028_));
  NO2        m1000(.A(mai_mai_n750_), .B(mai_mai_n106_), .Y(mai_mai_n1029_));
  NOi41      m1001(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1030_));
  NA2        m1002(.A(mai_mai_n1030_), .B(mai_mai_n1029_), .Y(mai_mai_n1031_));
  NO2        m1003(.A(mai_mai_n1031_), .B(mai_mai_n142_), .Y(mai_mai_n1032_));
  OR3        m1004(.A(e), .B(d), .C(c), .Y(mai_mai_n1033_));
  NA3        m1005(.A(k), .B(j), .C(i), .Y(mai_mai_n1034_));
  NO3        m1006(.A(mai_mai_n1034_), .B(mai_mai_n300_), .C(mai_mai_n85_), .Y(mai_mai_n1035_));
  OR4        m1007(.A(mai_mai_n1035_), .B(mai_mai_n1032_), .C(mai_mai_n1028_), .D(mai_mai_n1025_), .Y(mai_mai_n1036_));
  NA3        m1008(.A(mai_mai_n457_), .B(mai_mai_n326_), .C(mai_mai_n53_), .Y(mai_mai_n1037_));
  NO2        m1009(.A(mai_mai_n1037_), .B(mai_mai_n1027_), .Y(mai_mai_n1038_));
  NO4        m1010(.A(mai_mai_n1037_), .B(mai_mai_n574_), .C(mai_mai_n440_), .D(mai_mai_n44_), .Y(mai_mai_n1039_));
  NO2        m1011(.A(f), .B(c), .Y(mai_mai_n1040_));
  NOi21      m1012(.An(mai_mai_n1040_), .B(mai_mai_n433_), .Y(mai_mai_n1041_));
  NA2        m1013(.A(mai_mai_n1041_), .B(mai_mai_n56_), .Y(mai_mai_n1042_));
  OR2        m1014(.A(k), .B(i), .Y(mai_mai_n1043_));
  NO3        m1015(.A(mai_mai_n1043_), .B(mai_mai_n238_), .C(l), .Y(mai_mai_n1044_));
  NOi31      m1016(.An(mai_mai_n1044_), .B(mai_mai_n1042_), .C(j), .Y(mai_mai_n1045_));
  OR3        m1017(.A(mai_mai_n1045_), .B(mai_mai_n1039_), .C(mai_mai_n1038_), .Y(mai_mai_n1046_));
  OR3        m1018(.A(mai_mai_n1046_), .B(mai_mai_n1036_), .C(mai_mai_n1023_), .Y(mai02));
  OR2        m1019(.A(l), .B(k), .Y(mai_mai_n1048_));
  OR3        m1020(.A(n), .B(m), .C(i), .Y(mai_mai_n1049_));
  NO4        m1021(.A(mai_mai_n1049_), .B(h), .C(mai_mai_n1048_), .D(mai_mai_n1033_), .Y(mai_mai_n1050_));
  NO2        m1022(.A(mai_mai_n1035_), .B(mai_mai_n1015_), .Y(mai_mai_n1051_));
  AN3        m1023(.A(g), .B(f), .C(c), .Y(mai_mai_n1052_));
  NA3        m1024(.A(mai_mai_n1052_), .B(mai_mai_n457_), .C(h), .Y(mai_mai_n1053_));
  OR2        m1025(.A(mai_mai_n1034_), .B(mai_mai_n300_), .Y(mai_mai_n1054_));
  OR2        m1026(.A(mai_mai_n1054_), .B(mai_mai_n1053_), .Y(mai_mai_n1055_));
  NO3        m1027(.A(mai_mai_n1037_), .B(mai_mai_n1014_), .C(mai_mai_n574_), .Y(mai_mai_n1056_));
  NO2        m1028(.A(mai_mai_n1056_), .B(mai_mai_n1025_), .Y(mai_mai_n1057_));
  NA3        m1029(.A(l), .B(k), .C(j), .Y(mai_mai_n1058_));
  NA2        m1030(.A(i), .B(h), .Y(mai_mai_n1059_));
  NO3        m1031(.A(mai_mai_n1059_), .B(mai_mai_n1058_), .C(mai_mai_n126_), .Y(mai_mai_n1060_));
  NO3        m1032(.A(mai_mai_n137_), .B(mai_mai_n279_), .C(mai_mai_n209_), .Y(mai_mai_n1061_));
  AOI210     m1033(.A0(mai_mai_n1061_), .A1(mai_mai_n1060_), .B0(mai_mai_n1028_), .Y(mai_mai_n1062_));
  NA3        m1034(.A(c), .B(b), .C(a), .Y(mai_mai_n1063_));
  NO3        m1035(.A(mai_mai_n1063_), .B(mai_mai_n880_), .C(mai_mai_n208_), .Y(mai_mai_n1064_));
  NO4        m1036(.A(mai_mai_n1034_), .B(mai_mai_n293_), .C(mai_mai_n47_), .D(mai_mai_n106_), .Y(mai_mai_n1065_));
  AOI210     m1037(.A0(mai_mai_n1065_), .A1(mai_mai_n1064_), .B0(mai_mai_n1038_), .Y(mai_mai_n1066_));
  AN4        m1038(.A(mai_mai_n1066_), .B(mai_mai_n1062_), .C(mai_mai_n1057_), .D(mai_mai_n1055_), .Y(mai_mai_n1067_));
  INV        m1039(.A(mai_mai_n1016_), .Y(mai_mai_n1068_));
  NA2        m1040(.A(mai_mai_n1031_), .B(mai_mai_n1024_), .Y(mai_mai_n1069_));
  AOI210     m1041(.A0(mai_mai_n1069_), .A1(mai_mai_n1068_), .B0(mai_mai_n1011_), .Y(mai_mai_n1070_));
  NAi41      m1042(.An(mai_mai_n1050_), .B(mai_mai_n1070_), .C(mai_mai_n1067_), .D(mai_mai_n1051_), .Y(mai03));
  NO2        m1043(.A(mai_mai_n515_), .B(mai_mai_n587_), .Y(mai_mai_n1072_));
  NA4        m1044(.A(mai_mai_n82_), .B(mai_mai_n81_), .C(g), .D(mai_mai_n208_), .Y(mai_mai_n1073_));
  NA4        m1045(.A(h), .B(m), .C(mai_mai_n106_), .D(mai_mai_n208_), .Y(mai_mai_n1074_));
  NA3        m1046(.A(mai_mai_n1074_), .B(mai_mai_n359_), .C(mai_mai_n1073_), .Y(mai_mai_n1075_));
  NO3        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1072_), .C(mai_mai_n975_), .Y(mai_mai_n1076_));
  NOi41      m1048(.An(mai_mai_n795_), .B(mai_mai_n837_), .C(mai_mai_n830_), .D(mai_mai_n700_), .Y(mai_mai_n1077_));
  OAI220     m1049(.A0(mai_mai_n1077_), .A1(mai_mai_n675_), .B0(mai_mai_n1076_), .B1(mai_mai_n575_), .Y(mai_mai_n1078_));
  NA4        m1050(.A(i), .B(e), .C(mai_mai_n335_), .D(mai_mai_n326_), .Y(mai_mai_n1079_));
  OAI210     m1051(.A0(mai_mai_n807_), .A1(mai_mai_n411_), .B0(mai_mai_n1079_), .Y(mai_mai_n1080_));
  NOi31      m1052(.An(m), .B(n), .C(f), .Y(mai_mai_n1081_));
  NA2        m1053(.A(mai_mai_n1081_), .B(mai_mai_n49_), .Y(mai_mai_n1082_));
  OAI220     m1054(.A0(mai_mai_n1369_), .A1(mai_mai_n1082_), .B0(mai_mai_n867_), .B1(mai_mai_n417_), .Y(mai_mai_n1083_));
  NOi21      m1055(.An(mai_mai_n845_), .B(mai_mai_n1009_), .Y(mai_mai_n1084_));
  NO4        m1056(.A(mai_mai_n1084_), .B(mai_mai_n1083_), .C(mai_mai_n1080_), .D(mai_mai_n974_), .Y(mai_mai_n1085_));
  INV        m1057(.A(mai_mai_n1015_), .Y(mai_mai_n1086_));
  NO2        m1058(.A(mai_mai_n81_), .B(g), .Y(mai_mai_n1087_));
  AOI210     m1059(.A0(mai_mai_n1087_), .A1(i), .B0(mai_mai_n1044_), .Y(mai_mai_n1088_));
  OR2        m1060(.A(mai_mai_n1088_), .B(mai_mai_n1042_), .Y(mai_mai_n1089_));
  NA3        m1061(.A(mai_mai_n1089_), .B(mai_mai_n1086_), .C(mai_mai_n1085_), .Y(mai_mai_n1090_));
  NO4        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1078_), .C(mai_mai_n809_), .D(mai_mai_n554_), .Y(mai_mai_n1091_));
  NA2        m1063(.A(c), .B(b), .Y(mai_mai_n1092_));
  NO2        m1064(.A(n), .B(mai_mai_n1092_), .Y(mai_mai_n1093_));
  OAI210     m1065(.A0(mai_mai_n843_), .A1(mai_mai_n822_), .B0(mai_mai_n405_), .Y(mai_mai_n1094_));
  OAI210     m1066(.A0(mai_mai_n1094_), .A1(mai_mai_n844_), .B0(mai_mai_n1093_), .Y(mai_mai_n1095_));
  NAi21      m1067(.An(mai_mai_n412_), .B(mai_mai_n1093_), .Y(mai_mai_n1096_));
  NA3        m1068(.A(mai_mai_n418_), .B(mai_mai_n547_), .C(f), .Y(mai_mai_n1097_));
  OAI210     m1069(.A0(mai_mai_n537_), .A1(mai_mai_n38_), .B0(c), .Y(mai_mai_n1098_));
  NA3        m1070(.A(mai_mai_n1098_), .B(mai_mai_n1097_), .C(mai_mai_n1096_), .Y(mai_mai_n1099_));
  NAi21      m1071(.An(f), .B(d), .Y(mai_mai_n1100_));
  NO2        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1063_), .Y(mai_mai_n1101_));
  AOI210     m1073(.A0(mai_mai_n1101_), .A1(mai_mai_n107_), .B0(mai_mai_n1099_), .Y(mai_mai_n1102_));
  NO2        m1074(.A(mai_mai_n178_), .B(mai_mai_n231_), .Y(mai_mai_n1103_));
  NA2        m1075(.A(mai_mai_n1103_), .B(m), .Y(mai_mai_n1104_));
  NO2        m1076(.A(mai_mai_n60_), .B(mai_mai_n1104_), .Y(mai_mai_n1105_));
  NA2        m1077(.A(mai_mai_n549_), .B(mai_mai_n400_), .Y(mai_mai_n1106_));
  NA2        m1078(.A(mai_mai_n437_), .B(mai_mai_n1101_), .Y(mai_mai_n1107_));
  NO2        m1079(.A(mai_mai_n362_), .B(mai_mai_n361_), .Y(mai_mai_n1108_));
  AOI210     m1080(.A0(mai_mai_n1103_), .A1(mai_mai_n420_), .B0(mai_mai_n937_), .Y(mai_mai_n1109_));
  NAi41      m1081(.An(mai_mai_n1108_), .B(mai_mai_n1109_), .C(mai_mai_n1107_), .D(mai_mai_n1106_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(mai_mai_n1110_), .B(mai_mai_n1105_), .Y(mai_mai_n1111_));
  NA4        m1083(.A(mai_mai_n1111_), .B(mai_mai_n1102_), .C(mai_mai_n1095_), .D(mai_mai_n1091_), .Y(mai00));
  AOI210     m1084(.A0(mai_mai_n292_), .A1(mai_mai_n209_), .B0(mai_mai_n271_), .Y(mai_mai_n1113_));
  NO2        m1085(.A(mai_mai_n1113_), .B(mai_mai_n566_), .Y(mai_mai_n1114_));
  AOI210     m1086(.A0(mai_mai_n877_), .A1(mai_mai_n920_), .B0(mai_mai_n1080_), .Y(mai_mai_n1115_));
  NO3        m1087(.A(mai_mai_n1056_), .B(mai_mai_n937_), .C(mai_mai_n697_), .Y(mai_mai_n1116_));
  NA3        m1088(.A(mai_mai_n1116_), .B(mai_mai_n1115_), .C(mai_mai_n976_), .Y(mai_mai_n1117_));
  NA2        m1089(.A(mai_mai_n496_), .B(f), .Y(mai_mai_n1118_));
  OAI210     m1090(.A0(m), .A1(mai_mai_n39_), .B0(mai_mai_n633_), .Y(mai_mai_n1119_));
  NA3        m1091(.A(mai_mai_n1119_), .B(mai_mai_n253_), .C(n), .Y(mai_mai_n1120_));
  AOI210     m1092(.A0(mai_mai_n1120_), .A1(mai_mai_n1118_), .B0(mai_mai_n1018_), .Y(mai_mai_n1121_));
  NO4        m1093(.A(mai_mai_n1121_), .B(mai_mai_n1117_), .C(mai_mai_n1114_), .D(mai_mai_n1036_), .Y(mai_mai_n1122_));
  NA3        m1094(.A(mai_mai_n162_), .B(mai_mai_n45_), .C(mai_mai_n44_), .Y(mai_mai_n1123_));
  NA3        m1095(.A(d), .B(mai_mai_n53_), .C(b), .Y(mai_mai_n1124_));
  NOi31      m1096(.An(n), .B(m), .C(i), .Y(mai_mai_n1125_));
  NA3        m1097(.A(mai_mai_n1125_), .B(mai_mai_n636_), .C(mai_mai_n49_), .Y(mai_mai_n1126_));
  OAI210     m1098(.A0(mai_mai_n1124_), .A1(mai_mai_n1123_), .B0(mai_mai_n1126_), .Y(mai_mai_n1127_));
  INV        m1099(.A(mai_mai_n565_), .Y(mai_mai_n1128_));
  NO4        m1100(.A(mai_mai_n1128_), .B(mai_mai_n1127_), .C(mai_mai_n1108_), .D(mai_mai_n896_), .Y(mai_mai_n1129_));
  NO4        m1101(.A(mai_mai_n1362_), .B(mai_mai_n346_), .C(mai_mai_n1092_), .D(mai_mai_n56_), .Y(mai_mai_n1130_));
  NA3        m1102(.A(mai_mai_n373_), .B(mai_mai_n216_), .C(g), .Y(mai_mai_n1131_));
  OA220      m1103(.A0(mai_mai_n1131_), .A1(mai_mai_n1124_), .B0(mai_mai_n374_), .B1(mai_mai_n129_), .Y(mai_mai_n1132_));
  NO2        m1104(.A(h), .B(g), .Y(mai_mai_n1133_));
  NA4        m1105(.A(mai_mai_n484_), .B(mai_mai_n457_), .C(mai_mai_n1133_), .D(mai_mai_n1008_), .Y(mai_mai_n1134_));
  OAI220     m1106(.A0(mai_mai_n515_), .A1(mai_mai_n587_), .B0(mai_mai_n86_), .B1(mai_mai_n85_), .Y(mai_mai_n1135_));
  AOI220     m1107(.A0(mai_mai_n1135_), .A1(mai_mai_n524_), .B0(mai_mai_n925_), .B1(mai_mai_n564_), .Y(mai_mai_n1136_));
  AOI220     m1108(.A0(mai_mai_n310_), .A1(mai_mai_n242_), .B0(mai_mai_n173_), .B1(mai_mai_n144_), .Y(mai_mai_n1137_));
  NA4        m1109(.A(mai_mai_n1137_), .B(mai_mai_n1136_), .C(mai_mai_n1134_), .D(mai_mai_n1132_), .Y(mai_mai_n1138_));
  NO3        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1130_), .C(mai_mai_n261_), .Y(mai_mai_n1139_));
  INV        m1111(.A(mai_mai_n314_), .Y(mai_mai_n1140_));
  AOI210     m1112(.A0(mai_mai_n242_), .A1(mai_mai_n338_), .B0(mai_mai_n567_), .Y(mai_mai_n1141_));
  NA3        m1113(.A(mai_mai_n1141_), .B(mai_mai_n1140_), .C(mai_mai_n150_), .Y(mai_mai_n1142_));
  NO2        m1114(.A(mai_mai_n233_), .B(mai_mai_n177_), .Y(mai_mai_n1143_));
  NA2        m1115(.A(mai_mai_n1143_), .B(mai_mai_n418_), .Y(mai_mai_n1144_));
  NA3        m1116(.A(mai_mai_n175_), .B(mai_mai_n106_), .C(g), .Y(mai_mai_n1145_));
  NOi31      m1117(.An(mai_mai_n852_), .B(h), .C(mai_mai_n1145_), .Y(mai_mai_n1146_));
  NAi31      m1118(.An(mai_mai_n181_), .B(mai_mai_n841_), .C(mai_mai_n457_), .Y(mai_mai_n1147_));
  NAi31      m1119(.An(mai_mai_n1146_), .B(mai_mai_n1147_), .C(mai_mai_n1144_), .Y(mai_mai_n1148_));
  NO2        m1120(.A(mai_mai_n270_), .B(mai_mai_n69_), .Y(mai_mai_n1149_));
  NO3        m1121(.A(mai_mai_n417_), .B(mai_mai_n820_), .C(n), .Y(mai_mai_n1150_));
  AOI210     m1122(.A0(mai_mai_n1150_), .A1(mai_mai_n1149_), .B0(mai_mai_n1050_), .Y(mai_mai_n1151_));
  NAi31      m1123(.An(mai_mai_n1021_), .B(mai_mai_n1151_), .C(mai_mai_n68_), .Y(mai_mai_n1152_));
  NO4        m1124(.A(mai_mai_n1152_), .B(mai_mai_n1148_), .C(mai_mai_n1142_), .D(mai_mai_n506_), .Y(mai_mai_n1153_));
  AN3        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1139_), .C(mai_mai_n1129_), .Y(mai_mai_n1154_));
  NA2        m1126(.A(mai_mai_n524_), .B(mai_mai_n95_), .Y(mai_mai_n1155_));
  NA3        m1127(.A(mai_mai_n1081_), .B(mai_mai_n594_), .C(h), .Y(mai_mai_n1156_));
  NA4        m1128(.A(mai_mai_n1156_), .B(mai_mai_n550_), .C(mai_mai_n1155_), .D(mai_mai_n236_), .Y(mai_mai_n1157_));
  NA2        m1129(.A(mai_mai_n1075_), .B(mai_mai_n524_), .Y(mai_mai_n1158_));
  NA4        m1130(.A(mai_mai_n636_), .B(mai_mai_n201_), .C(mai_mai_n216_), .D(h), .Y(mai_mai_n1159_));
  NA3        m1131(.A(mai_mai_n1159_), .B(mai_mai_n1158_), .C(mai_mai_n289_), .Y(mai_mai_n1160_));
  OAI210     m1132(.A0(mai_mai_n456_), .A1(mai_mai_n113_), .B0(mai_mai_n846_), .Y(mai_mai_n1161_));
  AOI210     m1133(.A0(mai_mai_n549_), .A1(mai_mai_n400_), .B0(mai_mai_n1161_), .Y(mai_mai_n1162_));
  OR4        m1134(.A(mai_mai_n1018_), .B(mai_mai_n266_), .C(mai_mai_n218_), .D(e), .Y(mai_mai_n1163_));
  NO2        m1135(.A(mai_mai_n212_), .B(mai_mai_n209_), .Y(mai_mai_n1164_));
  NA2        m1136(.A(n), .B(e), .Y(mai_mai_n1165_));
  NO2        m1137(.A(mai_mai_n1165_), .B(mai_mai_n142_), .Y(mai_mai_n1166_));
  AOI220     m1138(.A0(mai_mai_n1166_), .A1(mai_mai_n268_), .B0(mai_mai_n833_), .B1(mai_mai_n1164_), .Y(mai_mai_n1167_));
  OAI210     m1139(.A0(mai_mai_n347_), .A1(mai_mai_n304_), .B0(mai_mai_n439_), .Y(mai_mai_n1168_));
  NA4        m1140(.A(mai_mai_n1168_), .B(mai_mai_n1167_), .C(mai_mai_n1163_), .D(mai_mai_n1162_), .Y(mai_mai_n1169_));
  AOI210     m1141(.A0(mai_mai_n1166_), .A1(mai_mai_n834_), .B0(mai_mai_n808_), .Y(mai_mai_n1170_));
  AOI220     m1142(.A0(mai_mai_n933_), .A1(mai_mai_n564_), .B0(mai_mai_n636_), .B1(mai_mai_n239_), .Y(mai_mai_n1171_));
  NO2        m1143(.A(mai_mai_n62_), .B(h), .Y(mai_mai_n1172_));
  NO2        m1144(.A(mai_mai_n1016_), .B(mai_mai_n713_), .Y(mai_mai_n1173_));
  OAI210     m1145(.A0(mai_mai_n1061_), .A1(mai_mai_n1173_), .B0(mai_mai_n1172_), .Y(mai_mai_n1174_));
  NA4        m1146(.A(mai_mai_n1174_), .B(mai_mai_n1171_), .C(mai_mai_n1170_), .D(mai_mai_n848_), .Y(mai_mai_n1175_));
  NO4        m1147(.A(mai_mai_n1175_), .B(mai_mai_n1169_), .C(mai_mai_n1160_), .D(mai_mai_n1157_), .Y(mai_mai_n1176_));
  NA2        m1148(.A(mai_mai_n823_), .B(mai_mai_n745_), .Y(mai_mai_n1177_));
  NA4        m1149(.A(mai_mai_n1177_), .B(mai_mai_n1176_), .C(mai_mai_n1154_), .D(mai_mai_n1122_), .Y(mai01));
  AN2        m1150(.A(mai_mai_n998_), .B(mai_mai_n997_), .Y(mai_mai_n1179_));
  NO4        m1151(.A(mai_mai_n791_), .B(mai_mai_n784_), .C(mai_mai_n465_), .D(mai_mai_n277_), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n580_), .B(mai_mai_n283_), .Y(mai_mai_n1181_));
  OAI210     m1153(.A0(mai_mai_n1181_), .A1(mai_mai_n384_), .B0(i), .Y(mai_mai_n1182_));
  NA3        m1154(.A(mai_mai_n1182_), .B(mai_mai_n1180_), .C(mai_mai_n1179_), .Y(mai_mai_n1183_));
  NA2        m1155(.A(mai_mai_n576_), .B(mai_mai_n84_), .Y(mai_mai_n1184_));
  NA2        m1156(.A(mai_mai_n939_), .B(c), .Y(mai_mai_n1185_));
  NA4        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1184_), .C(mai_mai_n890_), .D(mai_mai_n325_), .Y(mai_mai_n1186_));
  NA2        m1158(.A(l), .B(mai_mai_n91_), .Y(mai_mai_n1187_));
  OAI210     m1159(.A0(mai_mai_n772_), .A1(mai_mai_n591_), .B0(mai_mai_n1159_), .Y(mai_mai_n1188_));
  AOI210     m1160(.A0(mai_mai_n91_), .A1(mai_mai_n622_), .B0(mai_mai_n1188_), .Y(mai_mai_n1189_));
  OA210      m1161(.A0(mai_mai_n648_), .A1(mai_mai_n359_), .B0(mai_mai_n573_), .Y(mai_mai_n1190_));
  NAi41      m1162(.An(mai_mai_n157_), .B(mai_mai_n1190_), .C(mai_mai_n1189_), .D(mai_mai_n876_), .Y(mai_mai_n1191_));
  NO3        m1163(.A(mai_mai_n773_), .B(mai_mai_n662_), .C(mai_mai_n499_), .Y(mai_mai_n1192_));
  OR2        m1164(.A(mai_mai_n191_), .B(mai_mai_n189_), .Y(mai_mai_n1193_));
  NA3        m1165(.A(mai_mai_n1193_), .B(mai_mai_n1192_), .C(mai_mai_n132_), .Y(mai_mai_n1194_));
  NO4        m1166(.A(mai_mai_n1194_), .B(mai_mai_n1191_), .C(mai_mai_n1186_), .D(mai_mai_n1183_), .Y(mai_mai_n1195_));
  NA2        m1167(.A(mai_mai_n579_), .B(mai_mai_n573_), .Y(mai_mai_n1196_));
  AOI210     m1168(.A0(mai_mai_n551_), .A1(a), .B0(mai_mai_n1196_), .Y(mai_mai_n1197_));
  AOI210     m1169(.A0(mai_mai_n199_), .A1(mai_mai_n83_), .B0(mai_mai_n208_), .Y(mai_mai_n1198_));
  OAI210     m1170(.A0(mai_mai_n796_), .A1(mai_mai_n418_), .B0(mai_mai_n1198_), .Y(mai_mai_n1199_));
  OAI210     m1171(.A0(g), .A1(mai_mai_n33_), .B0(m), .Y(mai_mai_n1200_));
  NA2        m1172(.A(mai_mai_n198_), .B(mai_mai_n33_), .Y(mai_mai_n1201_));
  AO210      m1173(.A0(mai_mai_n1201_), .A1(mai_mai_n1200_), .B0(mai_mai_n324_), .Y(mai_mai_n1202_));
  NA4        m1174(.A(mai_mai_n1202_), .B(mai_mai_n1199_), .C(mai_mai_n1197_), .D(mai_mai_n202_), .Y(mai_mai_n1203_));
  AOI210     m1175(.A0(mai_mai_n585_), .A1(mai_mai_n112_), .B0(mai_mai_n590_), .Y(mai_mai_n1204_));
  NA2        m1176(.A(mai_mai_n582_), .B(mai_mai_n1204_), .Y(mai_mai_n1205_));
  NA2        m1177(.A(mai_mai_n276_), .B(mai_mai_n191_), .Y(mai_mai_n1206_));
  OAI210     m1178(.A0(mai_mai_n1206_), .A1(mai_mai_n375_), .B0(mai_mai_n653_), .Y(mai_mai_n1207_));
  NO2        m1179(.A(mai_mai_n807_), .B(mai_mai_n199_), .Y(mai_mai_n1208_));
  NO2        m1180(.A(mai_mai_n1208_), .B(mai_mai_n937_), .Y(mai_mai_n1209_));
  OAI210     m1181(.A0(mai_mai_n91_), .A1(mai_mai_n318_), .B0(mai_mai_n663_), .Y(mai_mai_n1210_));
  NA4        m1182(.A(mai_mai_n1210_), .B(mai_mai_n1209_), .C(mai_mai_n1207_), .D(mai_mai_n776_), .Y(mai_mai_n1211_));
  NO3        m1183(.A(mai_mai_n1211_), .B(mai_mai_n1205_), .C(mai_mai_n1203_), .Y(mai_mai_n1212_));
  NA2        m1184(.A(mai_mai_n592_), .B(f), .Y(mai_mai_n1213_));
  NO2        m1185(.A(mai_mai_n1213_), .B(mai_mai_n199_), .Y(mai_mai_n1214_));
  AOI210     m1186(.A0(mai_mai_n491_), .A1(mai_mai_n55_), .B0(mai_mai_n1214_), .Y(mai_mai_n1215_));
  OR2        m1187(.A(mai_mai_n1187_), .B(mai_mai_n593_), .Y(mai_mai_n1216_));
  NA3        m1188(.A(g), .B(k), .C(i), .Y(mai_mai_n1217_));
  NO2        m1189(.A(mai_mai_n1217_), .B(mai_mai_n955_), .Y(mai_mai_n1218_));
  NO2        m1190(.A(mai_mai_n202_), .B(mai_mai_n105_), .Y(mai_mai_n1219_));
  NO3        m1191(.A(mai_mai_n1219_), .B(mai_mai_n1218_), .C(mai_mai_n1127_), .Y(mai_mai_n1220_));
  NA4        m1192(.A(mai_mai_n1220_), .B(mai_mai_n1216_), .C(mai_mai_n1215_), .D(mai_mai_n744_), .Y(mai_mai_n1221_));
  NO2        m1193(.A(mai_mai_n944_), .B(mai_mai_n226_), .Y(mai_mai_n1222_));
  NO2        m1194(.A(mai_mai_n945_), .B(mai_mai_n544_), .Y(mai_mai_n1223_));
  OAI210     m1195(.A0(mai_mai_n1223_), .A1(mai_mai_n1222_), .B0(mai_mai_n333_), .Y(mai_mai_n1224_));
  NA2        m1196(.A(mai_mai_n560_), .B(mai_mai_n559_), .Y(mai_mai_n1225_));
  NO3        m1197(.A(mai_mai_n73_), .B(mai_mai_n293_), .C(mai_mai_n44_), .Y(mai_mai_n1226_));
  NA2        m1198(.A(mai_mai_n1226_), .B(mai_mai_n542_), .Y(mai_mai_n1227_));
  NA3        m1199(.A(mai_mai_n1227_), .B(mai_mai_n1225_), .C(mai_mai_n658_), .Y(mai_mai_n1228_));
  OR2        m1200(.A(mai_mai_n1131_), .B(mai_mai_n1124_), .Y(mai_mai_n1229_));
  NO2        m1201(.A(mai_mai_n359_), .B(mai_mai_n67_), .Y(mai_mai_n1230_));
  AOI210     m1202(.A0(mai_mai_n718_), .A1(mai_mai_n107_), .B0(mai_mai_n1230_), .Y(mai_mai_n1231_));
  NA2        m1203(.A(mai_mai_n1226_), .B(mai_mai_n798_), .Y(mai_mai_n1232_));
  NA4        m1204(.A(mai_mai_n1232_), .B(mai_mai_n1231_), .C(mai_mai_n1229_), .D(mai_mai_n376_), .Y(mai_mai_n1233_));
  NOi41      m1205(.An(mai_mai_n1224_), .B(mai_mai_n1233_), .C(mai_mai_n1228_), .D(mai_mai_n1221_), .Y(mai_mai_n1234_));
  NO2        m1206(.A(mai_mai_n125_), .B(mai_mai_n44_), .Y(mai_mai_n1235_));
  AO220      m1207(.A0(i), .A1(mai_mai_n609_), .B0(mai_mai_n1235_), .B1(mai_mai_n691_), .Y(mai_mai_n1236_));
  NO3        m1208(.A(mai_mai_n1059_), .B(mai_mai_n172_), .C(mai_mai_n81_), .Y(mai_mai_n1237_));
  NO2        m1209(.A(mai_mai_n602_), .B(mai_mai_n601_), .Y(mai_mai_n1238_));
  NO4        m1210(.A(mai_mai_n1059_), .B(mai_mai_n1238_), .C(mai_mai_n170_), .D(mai_mai_n81_), .Y(mai_mai_n1239_));
  NO3        m1211(.A(mai_mai_n1239_), .B(mai_mai_n1237_), .C(mai_mai_n626_), .Y(mai_mai_n1240_));
  NA4        m1212(.A(mai_mai_n1240_), .B(mai_mai_n1234_), .C(mai_mai_n1212_), .D(mai_mai_n1195_), .Y(mai06));
  NO2        m1213(.A(mai_mai_n399_), .B(mai_mai_n548_), .Y(mai_mai_n1242_));
  OAI210     m1214(.A0(mai_mai_n107_), .A1(mai_mai_n262_), .B0(mai_mai_n1242_), .Y(mai_mai_n1243_));
  NO2        m1215(.A(mai_mai_n220_), .B(mai_mai_n97_), .Y(mai_mai_n1244_));
  OAI210     m1216(.A0(mai_mai_n1244_), .A1(mai_mai_n1237_), .B0(mai_mai_n372_), .Y(mai_mai_n1245_));
  NA4        m1217(.A(mai_mai_n867_), .B(mai_mai_n1245_), .C(mai_mai_n1243_), .D(mai_mai_n1224_), .Y(mai_mai_n1246_));
  NO3        m1218(.A(mai_mai_n1246_), .B(mai_mai_n1228_), .C(mai_mai_n252_), .Y(mai_mai_n1247_));
  NO2        m1219(.A(mai_mai_n293_), .B(mai_mai_n44_), .Y(mai_mai_n1248_));
  AOI210     m1220(.A0(mai_mai_n1248_), .A1(mai_mai_n949_), .B0(mai_mai_n1222_), .Y(mai_mai_n1249_));
  AOI210     m1221(.A0(mai_mai_n1248_), .A1(mai_mai_n545_), .B0(mai_mai_n1236_), .Y(mai_mai_n1250_));
  AOI210     m1222(.A0(mai_mai_n1250_), .A1(mai_mai_n1249_), .B0(mai_mai_n330_), .Y(mai_mai_n1251_));
  OAI210     m1223(.A0(mai_mai_n83_), .A1(mai_mai_n39_), .B0(mai_mai_n661_), .Y(mai_mai_n1252_));
  NA2        m1224(.A(mai_mai_n1252_), .B(mai_mai_n630_), .Y(mai_mai_n1253_));
  NO2        m1225(.A(mai_mai_n502_), .B(mai_mai_n167_), .Y(mai_mai_n1254_));
  AOI210     m1226(.A0(mai_mai_n595_), .A1(mai_mai_n54_), .B0(mai_mai_n1082_), .Y(mai_mai_n1255_));
  OAI210     m1227(.A0(mai_mai_n451_), .A1(mai_mai_n243_), .B0(mai_mai_n886_), .Y(mai_mai_n1256_));
  NO4        m1228(.A(mai_mai_n1256_), .B(mai_mai_n1255_), .C(mai_mai_n131_), .D(mai_mai_n1254_), .Y(mai_mai_n1257_));
  OR2        m1229(.A(mai_mai_n589_), .B(mai_mai_n588_), .Y(mai_mai_n1258_));
  NO2        m1230(.A(mai_mai_n1363_), .B(mai_mai_n130_), .Y(mai_mai_n1259_));
  AOI210     m1231(.A0(mai_mai_n1259_), .A1(mai_mai_n576_), .B0(mai_mai_n1258_), .Y(mai_mai_n1260_));
  NA3        m1232(.A(mai_mai_n1260_), .B(mai_mai_n1257_), .C(mai_mai_n1253_), .Y(mai_mai_n1261_));
  NO2        m1233(.A(mai_mai_n735_), .B(mai_mai_n358_), .Y(mai_mai_n1262_));
  NOi21      m1234(.An(mai_mai_n1262_), .B(mai_mai_n47_), .Y(mai_mai_n1263_));
  AN2        m1235(.A(mai_mai_n933_), .B(c), .Y(mai_mai_n1264_));
  NO4        m1236(.A(mai_mai_n1264_), .B(mai_mai_n1263_), .C(mai_mai_n1261_), .D(mai_mai_n1251_), .Y(mai_mai_n1265_));
  NO2        m1237(.A(mai_mai_n220_), .B(mai_mai_n604_), .Y(mai_mai_n1266_));
  OAI210     m1238(.A0(mai_mai_n272_), .A1(c), .B0(mai_mai_n629_), .Y(mai_mai_n1267_));
  AOI220     m1239(.A0(mai_mai_n1267_), .A1(mai_mai_n1266_), .B0(mai_mai_n45_), .B1(mai_mai_n262_), .Y(mai_mai_n1268_));
  NO3        m1240(.A(mai_mai_n238_), .B(mai_mai_n97_), .C(mai_mai_n279_), .Y(mai_mai_n1269_));
  OAI220     m1241(.A0(mai_mai_n684_), .A1(mai_mai_n243_), .B0(mai_mai_n498_), .B1(mai_mai_n502_), .Y(mai_mai_n1270_));
  NO2        m1242(.A(mai_mai_n587_), .B(j), .Y(mai_mai_n1271_));
  NOi21      m1243(.An(mai_mai_n1271_), .B(mai_mai_n67_), .Y(mai_mai_n1272_));
  NO4        m1244(.A(mai_mai_n1272_), .B(mai_mai_n1270_), .C(mai_mai_n1269_), .D(mai_mai_n1083_), .Y(mai_mai_n1273_));
  NAi31      m1245(.An(mai_mai_n735_), .B(mai_mai_n78_), .C(mai_mai_n198_), .Y(mai_mai_n1274_));
  NA4        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1273_), .C(mai_mai_n1268_), .D(mai_mai_n1171_), .Y(mai_mai_n1275_));
  OR2        m1247(.A(mai_mai_n772_), .B(mai_mai_n529_), .Y(mai_mai_n1276_));
  OR3        m1248(.A(mai_mai_n361_), .B(mai_mai_n220_), .C(mai_mai_n604_), .Y(mai_mai_n1277_));
  AOI210     m1249(.A0(mai_mai_n560_), .A1(mai_mai_n439_), .B0(mai_mai_n363_), .Y(mai_mai_n1278_));
  NA2        m1250(.A(mai_mai_n1271_), .B(mai_mai_n780_), .Y(mai_mai_n1279_));
  NA4        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1278_), .C(mai_mai_n1277_), .D(mai_mai_n1276_), .Y(mai_mai_n1280_));
  AOI220     m1252(.A0(mai_mai_n1262_), .A1(mai_mai_n745_), .B0(mai_mai_n1259_), .B1(mai_mai_n232_), .Y(mai_mai_n1281_));
  AO220      m1253(.A0(mai_mai_n1244_), .A1(mai_mai_n653_), .B0(mai_mai_n905_), .B1(mai_mai_n904_), .Y(mai_mai_n1282_));
  NO4        m1254(.A(mai_mai_n1282_), .B(mai_mai_n857_), .C(mai_mai_n487_), .D(mai_mai_n468_), .Y(mai_mai_n1283_));
  NA3        m1255(.A(mai_mai_n1283_), .B(mai_mai_n1281_), .C(mai_mai_n1232_), .Y(mai_mai_n1284_));
  NAi21      m1256(.An(j), .B(i), .Y(mai_mai_n1285_));
  NO4        m1257(.A(mai_mai_n1238_), .B(mai_mai_n1285_), .C(mai_mai_n433_), .D(mai_mai_n229_), .Y(mai_mai_n1286_));
  NO4        m1258(.A(mai_mai_n1286_), .B(mai_mai_n1284_), .C(mai_mai_n1280_), .D(mai_mai_n1275_), .Y(mai_mai_n1287_));
  NA4        m1259(.A(mai_mai_n1287_), .B(mai_mai_n1265_), .C(mai_mai_n1247_), .D(mai_mai_n1240_), .Y(mai07));
  NAi21      m1260(.An(f), .B(c), .Y(mai_mai_n1289_));
  OR2        m1261(.A(e), .B(d), .Y(mai_mai_n1290_));
  OAI220     m1262(.A0(mai_mai_n1290_), .A1(mai_mai_n1289_), .B0(mai_mai_n614_), .B1(mai_mai_n315_), .Y(mai_mai_n1291_));
  NA3        m1263(.A(mai_mai_n1291_), .B(mai_mai_n1359_), .C(mai_mai_n175_), .Y(mai_mai_n1292_));
  NOi31      m1264(.An(n), .B(m), .C(b), .Y(mai_mai_n1293_));
  NOi41      m1265(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1294_));
  NA3        m1266(.A(mai_mai_n681_), .B(mai_mai_n667_), .C(mai_mai_n106_), .Y(mai_mai_n1295_));
  NO2        m1267(.A(mai_mai_n1295_), .B(mai_mai_n44_), .Y(mai_mai_n1296_));
  NO2        m1268(.A(l), .B(k), .Y(mai_mai_n1297_));
  NO3        m1269(.A(mai_mai_n433_), .B(d), .C(c), .Y(mai_mai_n1298_));
  INV        m1270(.A(mai_mai_n1296_), .Y(mai_mai_n1299_));
  NO2        m1271(.A(g), .B(c), .Y(mai_mai_n1300_));
  NA2        m1272(.A(mai_mai_n1100_), .B(h), .Y(mai_mai_n1301_));
  NA2        m1273(.A(mai_mai_n133_), .B(mai_mai_n216_), .Y(mai_mai_n1302_));
  NO2        m1274(.A(mai_mai_n1302_), .B(mai_mai_n1301_), .Y(mai_mai_n1303_));
  NOi31      m1275(.An(m), .B(n), .C(b), .Y(mai_mai_n1304_));
  INV        m1276(.A(mai_mai_n1303_), .Y(mai_mai_n1305_));
  OAI210     m1277(.A0(mai_mai_n178_), .A1(mai_mai_n514_), .B0(mai_mai_n1030_), .Y(mai_mai_n1306_));
  AN2        m1278(.A(mai_mai_n1306_), .B(mai_mai_n1305_), .Y(mai_mai_n1307_));
  NA2        m1279(.A(mai_mai_n1298_), .B(mai_mai_n210_), .Y(mai_mai_n1308_));
  INV        m1280(.A(mai_mai_n1308_), .Y(mai_mai_n1309_));
  NO4        m1281(.A(mai_mai_n126_), .B(g), .C(f), .D(e), .Y(mai_mai_n1310_));
  NA2        m1282(.A(mai_mai_n29_), .B(h), .Y(mai_mai_n1311_));
  NO2        m1283(.A(mai_mai_n1311_), .B(mai_mai_n1049_), .Y(mai_mai_n1312_));
  NA2        m1284(.A(mai_mai_n1294_), .B(mai_mai_n1297_), .Y(mai_mai_n1313_));
  NA2        m1285(.A(mai_mai_n1081_), .B(mai_mai_n398_), .Y(mai_mai_n1314_));
  NO3        m1286(.A(mai_mai_n1360_), .B(mai_mai_n1312_), .C(mai_mai_n1309_), .Y(mai_mai_n1315_));
  NA4        m1287(.A(mai_mai_n1315_), .B(mai_mai_n1307_), .C(mai_mai_n1299_), .D(mai_mai_n1292_), .Y(mai_mai_n1316_));
  NO3        m1288(.A(mai_mai_n735_), .B(mai_mai_n170_), .C(mai_mai_n401_), .Y(mai_mai_n1317_));
  INV        m1289(.A(mai_mai_n1317_), .Y(mai_mai_n1318_));
  OR2        m1290(.A(n), .B(i), .Y(mai_mai_n1319_));
  OAI210     m1291(.A0(mai_mai_n1319_), .A1(mai_mai_n1040_), .B0(mai_mai_n47_), .Y(mai_mai_n1320_));
  AOI220     m1292(.A0(mai_mai_n1320_), .A1(mai_mai_n1133_), .B0(mai_mai_n812_), .B1(mai_mai_n190_), .Y(mai_mai_n1321_));
  NOi21      m1293(.An(d), .B(f), .Y(mai_mai_n1322_));
  NA2        m1294(.A(mai_mai_n1321_), .B(mai_mai_n1318_), .Y(mai_mai_n1323_));
  OAI210     m1295(.A0(mai_mai_n1310_), .A1(mai_mai_n1293_), .B0(mai_mai_n864_), .Y(mai_mai_n1324_));
  INV        m1296(.A(mai_mai_n1324_), .Y(mai_mai_n1325_));
  NA2        m1297(.A(mai_mai_n1300_), .B(mai_mai_n1322_), .Y(mai_mai_n1326_));
  NO2        m1298(.A(mai_mai_n1326_), .B(m), .Y(mai_mai_n1327_));
  NA2        m1299(.A(mai_mai_n104_), .B(mai_mai_n1304_), .Y(mai_mai_n1328_));
  INV        m1300(.A(mai_mai_n1328_), .Y(mai_mai_n1329_));
  NO3        m1301(.A(mai_mai_n1329_), .B(mai_mai_n1327_), .C(mai_mai_n1325_), .Y(mai_mai_n1330_));
  NO2        m1302(.A(mai_mai_n1289_), .B(e), .Y(mai_mai_n1331_));
  NA2        m1303(.A(mai_mai_n1087_), .B(mai_mai_n618_), .Y(mai_mai_n1332_));
  NO2        m1304(.A(mai_mai_n1332_), .B(mai_mai_n435_), .Y(mai_mai_n1333_));
  INV        m1305(.A(mai_mai_n1333_), .Y(mai_mai_n1334_));
  NO2        m1306(.A(mai_mai_n177_), .B(c), .Y(mai_mai_n1335_));
  OAI210     m1307(.A0(mai_mai_n1335_), .A1(mai_mai_n1331_), .B0(mai_mai_n175_), .Y(mai_mai_n1336_));
  AOI220     m1308(.A0(mai_mai_n1336_), .A1(mai_mai_n1042_), .B0(mai_mai_n521_), .B1(mai_mai_n358_), .Y(mai_mai_n1337_));
  NA2        m1309(.A(mai_mai_n528_), .B(g), .Y(mai_mai_n1338_));
  NA2        m1310(.A(mai_mai_n1338_), .B(mai_mai_n1298_), .Y(mai_mai_n1339_));
  NO2        m1311(.A(mai_mai_n1339_), .B(mai_mai_n208_), .Y(mai_mai_n1340_));
  NO2        m1312(.A(mai_mai_n1340_), .B(mai_mai_n1337_), .Y(mai_mai_n1341_));
  NA3        m1313(.A(mai_mai_n1341_), .B(mai_mai_n1334_), .C(mai_mai_n1330_), .Y(mai_mai_n1342_));
  NA2        m1314(.A(mai_mai_n56_), .B(a), .Y(mai_mai_n1343_));
  NO2        m1315(.A(mai_mai_n1314_), .B(mai_mai_n1343_), .Y(mai_mai_n1344_));
  OR4        m1316(.A(mai_mai_n1344_), .B(mai_mai_n1342_), .C(mai_mai_n1323_), .D(mai_mai_n1316_), .Y(mai04));
  NOi31      m1317(.An(mai_mai_n1310_), .B(k), .C(mai_mai_n1018_), .Y(mai_mai_n1346_));
  NO4        m1318(.A(mai_mai_n1290_), .B(mai_mai_n1009_), .C(mai_mai_n470_), .D(j), .Y(mai_mai_n1347_));
  OR3        m1319(.A(mai_mai_n1347_), .B(mai_mai_n1346_), .C(mai_mai_n1032_), .Y(mai_mai_n1348_));
  NO2        m1320(.A(mai_mai_n85_), .B(k), .Y(mai_mai_n1349_));
  AOI210     m1321(.A0(mai_mai_n1349_), .A1(mai_mai_n1026_), .B0(mai_mai_n1146_), .Y(mai_mai_n1350_));
  NA2        m1322(.A(mai_mai_n1350_), .B(mai_mai_n1174_), .Y(mai_mai_n1351_));
  NO4        m1323(.A(mai_mai_n1351_), .B(mai_mai_n1348_), .C(mai_mai_n1039_), .D(mai_mai_n1023_), .Y(mai_mai_n1352_));
  NA4        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1089_), .C(mai_mai_n1079_), .D(mai_mai_n1067_), .Y(mai05));
  INV        m1325(.A(mai_mai_n428_), .Y(mai_mai_n1356_));
  INV        m1326(.A(m), .Y(mai_mai_n1357_));
  INV        m1327(.A(m), .Y(mai_mai_n1358_));
  INV        m1328(.A(j), .Y(mai_mai_n1359_));
  INV        m1329(.A(mai_mai_n1313_), .Y(mai_mai_n1360_));
  INV        m1330(.A(mai_mai_n681_), .Y(mai_mai_n1361_));
  INV        m1331(.A(mai_mai_n216_), .Y(mai_mai_n1362_));
  INV        m1332(.A(m), .Y(mai_mai_n1363_));
  INV        m1333(.A(b), .Y(mai_mai_n1364_));
  INV        m1334(.A(mai_mai_n578_), .Y(mai_mai_n1365_));
  INV        m1335(.A(c), .Y(mai_mai_n1366_));
  INV        m1336(.A(g), .Y(mai_mai_n1367_));
  INV        m1337(.A(g), .Y(mai_mai_n1368_));
  INV        m1338(.A(c), .Y(mai_mai_n1369_));
  INV        m1339(.A(a), .Y(mai_mai_n1370_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NAi21      u0031(.An(i), .B(h), .Y(men_men_n60_));
  NAi31      u0032(.An(i), .B(l), .C(j), .Y(men_men_n61_));
  OAI220     u0033(.A0(men_men_n61_), .A1(men_men_n49_), .B0(men_men_n60_), .B1(men_men_n44_), .Y(men_men_n62_));
  NAi31      u0034(.An(d), .B(men_men_n62_), .C(men_men_n58_), .Y(men_men_n63_));
  NAi41      u0035(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n64_));
  NA2        u0036(.A(g), .B(f), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi21      u0038(.An(i), .B(j), .Y(men_men_n67_));
  NAi32      u0039(.An(n), .Bn(k), .C(m), .Y(men_men_n68_));
  NO2        u0040(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi31      u0041(.An(l), .B(m), .C(k), .Y(men_men_n70_));
  NAi21      u0042(.An(e), .B(h), .Y(men_men_n71_));
  NAi41      u0043(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n73_));
  INV        u0045(.A(m), .Y(men_men_n74_));
  NOi21      u0046(.An(k), .B(l), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  AN4        u0048(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n77_));
  NOi31      u0049(.An(h), .B(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n78_), .B(men_men_n77_), .Y(men_men_n79_));
  NAi32      u0051(.An(m), .Bn(k), .C(j), .Y(men_men_n80_));
  NOi32      u0052(.An(h), .Bn(g), .C(f), .Y(men_men_n81_));
  NA2        u0053(.A(men_men_n81_), .B(men_men_n77_), .Y(men_men_n82_));
  OA220      u0054(.A0(men_men_n82_), .A1(men_men_n80_), .B0(men_men_n79_), .B1(men_men_n76_), .Y(men_men_n83_));
  NA3        u0055(.A(men_men_n83_), .B(men_men_n73_), .C(men_men_n63_), .Y(men_men_n84_));
  INV        u0056(.A(n), .Y(men_men_n85_));
  NOi32      u0057(.An(e), .Bn(b), .C(d), .Y(men_men_n86_));
  NA2        u0058(.A(men_men_n86_), .B(men_men_n85_), .Y(men_men_n87_));
  INV        u0059(.A(j), .Y(men_men_n88_));
  AN3        u0060(.A(m), .B(k), .C(i), .Y(men_men_n89_));
  NA3        u0061(.A(men_men_n89_), .B(men_men_n88_), .C(g), .Y(men_men_n90_));
  NO2        u0062(.A(men_men_n90_), .B(f), .Y(men_men_n91_));
  NAi32      u0063(.An(g), .Bn(f), .C(h), .Y(men_men_n92_));
  NAi31      u0064(.An(j), .B(m), .C(l), .Y(men_men_n93_));
  NO2        u0065(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NA2        u0066(.A(m), .B(l), .Y(men_men_n95_));
  NAi31      u0067(.An(k), .B(j), .C(g), .Y(men_men_n96_));
  NO3        u0068(.A(men_men_n96_), .B(men_men_n95_), .C(f), .Y(men_men_n97_));
  AN2        u0069(.A(j), .B(g), .Y(men_men_n98_));
  NOi32      u0070(.An(m), .Bn(l), .C(i), .Y(men_men_n99_));
  NOi21      u0071(.An(g), .B(i), .Y(men_men_n100_));
  NOi32      u0072(.An(m), .Bn(j), .C(k), .Y(men_men_n101_));
  AOI220     u0073(.A0(men_men_n101_), .A1(men_men_n100_), .B0(men_men_n99_), .B1(men_men_n98_), .Y(men_men_n102_));
  NO2        u0074(.A(men_men_n102_), .B(f), .Y(men_men_n103_));
  NO4        u0075(.A(men_men_n103_), .B(men_men_n97_), .C(men_men_n94_), .D(men_men_n91_), .Y(men_men_n104_));
  NAi41      u0076(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n105_));
  AN2        u0077(.A(e), .B(b), .Y(men_men_n106_));
  NOi31      u0078(.An(c), .B(h), .C(f), .Y(men_men_n107_));
  NA2        u0079(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NO3        u0080(.A(men_men_n108_), .B(men_men_n105_), .C(g), .Y(men_men_n109_));
  NOi21      u0081(.An(g), .B(f), .Y(men_men_n110_));
  NOi21      u0082(.An(i), .B(h), .Y(men_men_n111_));
  NA3        u0083(.A(men_men_n111_), .B(men_men_n110_), .C(men_men_n36_), .Y(men_men_n112_));
  INV        u0084(.A(a), .Y(men_men_n113_));
  NA2        u0085(.A(men_men_n106_), .B(men_men_n113_), .Y(men_men_n114_));
  INV        u0086(.A(l), .Y(men_men_n115_));
  NOi21      u0087(.An(m), .B(n), .Y(men_men_n116_));
  AN2        u0088(.A(k), .B(h), .Y(men_men_n117_));
  NO2        u0089(.A(men_men_n112_), .B(men_men_n87_), .Y(men_men_n118_));
  INV        u0090(.A(b), .Y(men_men_n119_));
  NA2        u0091(.A(l), .B(j), .Y(men_men_n120_));
  AN2        u0092(.A(k), .B(i), .Y(men_men_n121_));
  NA2        u0093(.A(men_men_n121_), .B(men_men_n120_), .Y(men_men_n122_));
  NA2        u0094(.A(g), .B(e), .Y(men_men_n123_));
  NOi32      u0095(.An(c), .Bn(a), .C(d), .Y(men_men_n124_));
  NA2        u0096(.A(men_men_n124_), .B(men_men_n116_), .Y(men_men_n125_));
  NO4        u0097(.A(men_men_n125_), .B(men_men_n123_), .C(men_men_n122_), .D(men_men_n119_), .Y(men_men_n126_));
  NO3        u0098(.A(men_men_n126_), .B(men_men_n118_), .C(men_men_n109_), .Y(men_men_n127_));
  OAI210     u0099(.A0(men_men_n104_), .A1(men_men_n87_), .B0(men_men_n127_), .Y(men_men_n128_));
  NOi31      u0100(.An(k), .B(m), .C(j), .Y(men_men_n129_));
  NA3        u0101(.A(men_men_n129_), .B(men_men_n78_), .C(men_men_n77_), .Y(men_men_n130_));
  NOi31      u0102(.An(k), .B(m), .C(i), .Y(men_men_n131_));
  NA3        u0103(.A(men_men_n131_), .B(men_men_n81_), .C(men_men_n77_), .Y(men_men_n132_));
  NA2        u0104(.A(men_men_n132_), .B(men_men_n130_), .Y(men_men_n133_));
  NOi32      u0105(.An(f), .Bn(b), .C(e), .Y(men_men_n134_));
  NAi21      u0106(.An(g), .B(h), .Y(men_men_n135_));
  NAi21      u0107(.An(m), .B(n), .Y(men_men_n136_));
  NAi21      u0108(.An(j), .B(k), .Y(men_men_n137_));
  NO3        u0109(.A(men_men_n137_), .B(men_men_n136_), .C(men_men_n135_), .Y(men_men_n138_));
  NAi41      u0110(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n139_));
  NAi31      u0111(.An(j), .B(k), .C(h), .Y(men_men_n140_));
  NO3        u0112(.A(men_men_n140_), .B(men_men_n139_), .C(men_men_n136_), .Y(men_men_n141_));
  AOI210     u0113(.A0(men_men_n138_), .A1(men_men_n134_), .B0(men_men_n141_), .Y(men_men_n142_));
  NO2        u0114(.A(k), .B(j), .Y(men_men_n143_));
  NO2        u0115(.A(men_men_n143_), .B(men_men_n136_), .Y(men_men_n144_));
  AN2        u0116(.A(k), .B(j), .Y(men_men_n145_));
  NAi21      u0117(.An(c), .B(b), .Y(men_men_n146_));
  NA2        u0118(.A(f), .B(d), .Y(men_men_n147_));
  NO4        u0119(.A(men_men_n147_), .B(men_men_n146_), .C(men_men_n145_), .D(men_men_n135_), .Y(men_men_n148_));
  NA2        u0120(.A(h), .B(c), .Y(men_men_n149_));
  NAi31      u0121(.An(f), .B(e), .C(b), .Y(men_men_n150_));
  NA2        u0122(.A(men_men_n148_), .B(men_men_n144_), .Y(men_men_n151_));
  NA2        u0123(.A(d), .B(b), .Y(men_men_n152_));
  NAi21      u0124(.An(e), .B(f), .Y(men_men_n153_));
  NO2        u0125(.A(men_men_n153_), .B(men_men_n152_), .Y(men_men_n154_));
  NA2        u0126(.A(b), .B(a), .Y(men_men_n155_));
  NAi21      u0127(.An(e), .B(g), .Y(men_men_n156_));
  NAi21      u0128(.An(c), .B(d), .Y(men_men_n157_));
  NAi31      u0129(.An(l), .B(k), .C(h), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n136_), .B(men_men_n158_), .Y(men_men_n159_));
  NA2        u0131(.A(men_men_n159_), .B(men_men_n154_), .Y(men_men_n160_));
  NAi41      u0132(.An(men_men_n133_), .B(men_men_n160_), .C(men_men_n151_), .D(men_men_n142_), .Y(men_men_n161_));
  NAi31      u0133(.An(e), .B(f), .C(b), .Y(men_men_n162_));
  NOi21      u0134(.An(g), .B(d), .Y(men_men_n163_));
  NO2        u0135(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  NOi21      u0136(.An(h), .B(i), .Y(men_men_n165_));
  NOi21      u0137(.An(k), .B(m), .Y(men_men_n166_));
  NA3        u0138(.A(men_men_n166_), .B(men_men_n165_), .C(n), .Y(men_men_n167_));
  NOi21      u0139(.An(men_men_n164_), .B(men_men_n167_), .Y(men_men_n168_));
  NOi21      u0140(.An(h), .B(g), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n147_), .B(men_men_n146_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  NAi31      u0143(.An(l), .B(j), .C(h), .Y(men_men_n172_));
  NO2        u0144(.A(men_men_n172_), .B(men_men_n49_), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n66_), .Y(men_men_n174_));
  NOi32      u0146(.An(n), .Bn(k), .C(m), .Y(men_men_n175_));
  NA2        u0147(.A(l), .B(i), .Y(men_men_n176_));
  NA2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  OAI210     u0149(.A0(men_men_n177_), .A1(men_men_n171_), .B0(men_men_n174_), .Y(men_men_n178_));
  NAi31      u0150(.An(d), .B(f), .C(c), .Y(men_men_n179_));
  NAi31      u0151(.An(e), .B(f), .C(c), .Y(men_men_n180_));
  NA2        u0152(.A(j), .B(h), .Y(men_men_n181_));
  OR3        u0153(.A(n), .B(m), .C(k), .Y(men_men_n182_));
  NO2        u0154(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  NAi32      u0155(.An(m), .Bn(k), .C(n), .Y(men_men_n184_));
  NO2        u0156(.A(men_men_n184_), .B(men_men_n181_), .Y(men_men_n185_));
  AOI220     u0157(.A0(men_men_n185_), .A1(men_men_n164_), .B0(men_men_n183_), .B1(f), .Y(men_men_n186_));
  NO2        u0158(.A(n), .B(m), .Y(men_men_n187_));
  NA2        u0159(.A(men_men_n187_), .B(men_men_n50_), .Y(men_men_n188_));
  NAi21      u0160(.An(f), .B(e), .Y(men_men_n189_));
  NA2        u0161(.A(d), .B(c), .Y(men_men_n190_));
  NOi21      u0162(.An(d), .B(men_men_n188_), .Y(men_men_n191_));
  NAi21      u0163(.An(d), .B(c), .Y(men_men_n192_));
  NAi31      u0164(.An(m), .B(n), .C(b), .Y(men_men_n193_));
  NA2        u0165(.A(k), .B(i), .Y(men_men_n194_));
  NAi21      u0166(.An(h), .B(f), .Y(men_men_n195_));
  INV        u0167(.A(men_men_n195_), .Y(men_men_n196_));
  NO2        u0168(.A(men_men_n193_), .B(men_men_n157_), .Y(men_men_n197_));
  NA2        u0169(.A(men_men_n197_), .B(men_men_n196_), .Y(men_men_n198_));
  NOi32      u0170(.An(f), .Bn(c), .C(e), .Y(men_men_n199_));
  NO3        u0171(.A(n), .B(m), .C(j), .Y(men_men_n200_));
  NA2        u0172(.A(men_men_n200_), .B(men_men_n117_), .Y(men_men_n201_));
  AO210      u0173(.A0(men_men_n201_), .A1(men_men_n188_), .B0(men_men_n1626_), .Y(men_men_n202_));
  NAi41      u0174(.An(men_men_n191_), .B(men_men_n202_), .C(men_men_n198_), .D(men_men_n186_), .Y(men_men_n203_));
  OR4        u0175(.A(men_men_n203_), .B(men_men_n178_), .C(men_men_n168_), .D(men_men_n161_), .Y(men_men_n204_));
  NO4        u0176(.A(men_men_n204_), .B(men_men_n128_), .C(men_men_n84_), .D(men_men_n55_), .Y(men_men_n205_));
  NA3        u0177(.A(m), .B(men_men_n115_), .C(j), .Y(men_men_n206_));
  NAi31      u0178(.An(n), .B(h), .C(g), .Y(men_men_n207_));
  NO2        u0179(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  NOi32      u0180(.An(m), .Bn(k), .C(l), .Y(men_men_n209_));
  NA3        u0181(.A(men_men_n209_), .B(men_men_n88_), .C(g), .Y(men_men_n210_));
  NO2        u0182(.A(men_men_n210_), .B(n), .Y(men_men_n211_));
  NOi21      u0183(.An(k), .B(j), .Y(men_men_n212_));
  NA4        u0184(.A(men_men_n212_), .B(men_men_n116_), .C(i), .D(g), .Y(men_men_n213_));
  AN2        u0185(.A(i), .B(g), .Y(men_men_n214_));
  NA3        u0186(.A(men_men_n75_), .B(men_men_n214_), .C(men_men_n116_), .Y(men_men_n215_));
  NA2        u0187(.A(men_men_n215_), .B(men_men_n213_), .Y(men_men_n216_));
  NO3        u0188(.A(men_men_n216_), .B(men_men_n211_), .C(men_men_n208_), .Y(men_men_n217_));
  NAi41      u0189(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n218_));
  INV        u0190(.A(men_men_n218_), .Y(men_men_n219_));
  INV        u0191(.A(f), .Y(men_men_n220_));
  INV        u0192(.A(g), .Y(men_men_n221_));
  NOi31      u0193(.An(i), .B(j), .C(h), .Y(men_men_n222_));
  NOi21      u0194(.An(l), .B(m), .Y(men_men_n223_));
  NA2        u0195(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n224_));
  NO3        u0196(.A(men_men_n224_), .B(men_men_n221_), .C(men_men_n220_), .Y(men_men_n225_));
  NA2        u0197(.A(men_men_n225_), .B(men_men_n219_), .Y(men_men_n226_));
  OAI210     u0198(.A0(men_men_n217_), .A1(men_men_n32_), .B0(men_men_n226_), .Y(men_men_n227_));
  NOi21      u0199(.An(n), .B(m), .Y(men_men_n228_));
  NA2        u0200(.A(i), .B(men_men_n228_), .Y(men_men_n229_));
  OA220      u0201(.A0(men_men_n229_), .A1(men_men_n108_), .B0(men_men_n80_), .B1(men_men_n79_), .Y(men_men_n230_));
  NAi21      u0202(.An(j), .B(h), .Y(men_men_n231_));
  XN2        u0203(.A(i), .B(h), .Y(men_men_n232_));
  NA2        u0204(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n233_));
  NOi31      u0205(.An(k), .B(n), .C(m), .Y(men_men_n234_));
  NOi31      u0206(.An(men_men_n234_), .B(men_men_n190_), .C(men_men_n189_), .Y(men_men_n235_));
  NA2        u0207(.A(men_men_n235_), .B(men_men_n233_), .Y(men_men_n236_));
  NAi31      u0208(.An(f), .B(e), .C(c), .Y(men_men_n237_));
  NO4        u0209(.A(men_men_n237_), .B(men_men_n182_), .C(men_men_n181_), .D(men_men_n59_), .Y(men_men_n238_));
  NA4        u0210(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n239_));
  NAi32      u0211(.An(m), .Bn(i), .C(k), .Y(men_men_n240_));
  NO3        u0212(.A(men_men_n240_), .B(men_men_n92_), .C(men_men_n239_), .Y(men_men_n241_));
  NA2        u0213(.A(k), .B(h), .Y(men_men_n242_));
  NO2        u0214(.A(men_men_n241_), .B(men_men_n238_), .Y(men_men_n243_));
  NAi21      u0215(.An(n), .B(a), .Y(men_men_n244_));
  NO2        u0216(.A(men_men_n244_), .B(men_men_n152_), .Y(men_men_n245_));
  NAi41      u0217(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n246_));
  NO2        u0218(.A(men_men_n246_), .B(e), .Y(men_men_n247_));
  NO3        u0219(.A(men_men_n153_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n248_));
  OAI210     u0220(.A0(men_men_n248_), .A1(men_men_n247_), .B0(men_men_n245_), .Y(men_men_n249_));
  AN4        u0221(.A(men_men_n249_), .B(men_men_n243_), .C(men_men_n236_), .D(men_men_n230_), .Y(men_men_n250_));
  OR2        u0222(.A(h), .B(g), .Y(men_men_n251_));
  NO2        u0223(.A(men_men_n251_), .B(men_men_n105_), .Y(men_men_n252_));
  NA2        u0224(.A(men_men_n252_), .B(men_men_n134_), .Y(men_men_n253_));
  NAi41      u0225(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n254_));
  NO2        u0226(.A(men_men_n254_), .B(men_men_n220_), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n166_), .B(men_men_n111_), .Y(men_men_n256_));
  NAi21      u0228(.An(men_men_n256_), .B(men_men_n255_), .Y(men_men_n257_));
  NO2        u0229(.A(n), .B(a), .Y(men_men_n258_));
  NAi31      u0230(.An(men_men_n246_), .B(men_men_n258_), .C(men_men_n106_), .Y(men_men_n259_));
  AN2        u0231(.A(men_men_n259_), .B(men_men_n257_), .Y(men_men_n260_));
  NAi21      u0232(.An(h), .B(i), .Y(men_men_n261_));
  NA2        u0233(.A(men_men_n187_), .B(k), .Y(men_men_n262_));
  NO2        u0234(.A(men_men_n262_), .B(men_men_n261_), .Y(men_men_n263_));
  NA2        u0235(.A(men_men_n263_), .B(f), .Y(men_men_n264_));
  NA3        u0236(.A(men_men_n264_), .B(men_men_n260_), .C(men_men_n253_), .Y(men_men_n265_));
  NOi21      u0237(.An(g), .B(e), .Y(men_men_n266_));
  NO2        u0238(.A(men_men_n72_), .B(men_men_n74_), .Y(men_men_n267_));
  NA2        u0239(.A(men_men_n267_), .B(men_men_n266_), .Y(men_men_n268_));
  NOi32      u0240(.An(l), .Bn(j), .C(i), .Y(men_men_n269_));
  AOI210     u0241(.A0(men_men_n75_), .A1(men_men_n88_), .B0(men_men_n269_), .Y(men_men_n270_));
  NO2        u0242(.A(men_men_n261_), .B(men_men_n44_), .Y(men_men_n271_));
  NAi21      u0243(.An(f), .B(g), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n272_), .B(men_men_n64_), .Y(men_men_n273_));
  NO2        u0245(.A(men_men_n68_), .B(men_men_n120_), .Y(men_men_n274_));
  AOI220     u0246(.A0(men_men_n274_), .A1(men_men_n273_), .B0(men_men_n271_), .B1(men_men_n66_), .Y(men_men_n275_));
  OAI210     u0247(.A0(men_men_n270_), .A1(men_men_n268_), .B0(men_men_n275_), .Y(men_men_n276_));
  NO3        u0248(.A(men_men_n137_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n277_));
  NOi41      u0249(.An(men_men_n250_), .B(men_men_n276_), .C(men_men_n265_), .D(men_men_n227_), .Y(men_men_n278_));
  NO4        u0250(.A(men_men_n208_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n279_));
  NO2        u0251(.A(men_men_n279_), .B(men_men_n114_), .Y(men_men_n280_));
  NA3        u0252(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n281_));
  NAi21      u0253(.An(h), .B(g), .Y(men_men_n282_));
  OR4        u0254(.A(men_men_n282_), .B(men_men_n281_), .C(men_men_n229_), .D(e), .Y(men_men_n283_));
  NO2        u0255(.A(men_men_n256_), .B(men_men_n272_), .Y(men_men_n284_));
  NA2        u0256(.A(men_men_n284_), .B(men_men_n77_), .Y(men_men_n285_));
  NAi31      u0257(.An(g), .B(k), .C(h), .Y(men_men_n286_));
  NO3        u0258(.A(men_men_n136_), .B(men_men_n286_), .C(l), .Y(men_men_n287_));
  NAi31      u0259(.An(e), .B(d), .C(a), .Y(men_men_n288_));
  NA2        u0260(.A(men_men_n287_), .B(men_men_n134_), .Y(men_men_n289_));
  NA3        u0261(.A(men_men_n289_), .B(men_men_n285_), .C(men_men_n283_), .Y(men_men_n290_));
  NA4        u0262(.A(men_men_n166_), .B(men_men_n81_), .C(men_men_n77_), .D(men_men_n120_), .Y(men_men_n291_));
  NA3        u0263(.A(men_men_n166_), .B(men_men_n165_), .C(men_men_n85_), .Y(men_men_n292_));
  NO2        u0264(.A(men_men_n292_), .B(men_men_n1626_), .Y(men_men_n293_));
  NOi21      u0265(.An(men_men_n291_), .B(men_men_n293_), .Y(men_men_n294_));
  NA3        u0266(.A(e), .B(c), .C(b), .Y(men_men_n295_));
  NO2        u0267(.A(d), .B(men_men_n295_), .Y(men_men_n296_));
  NAi32      u0268(.An(k), .Bn(i), .C(j), .Y(men_men_n297_));
  NAi31      u0269(.An(h), .B(l), .C(i), .Y(men_men_n298_));
  NA3        u0270(.A(men_men_n298_), .B(men_men_n297_), .C(men_men_n172_), .Y(men_men_n299_));
  NOi21      u0271(.An(men_men_n299_), .B(men_men_n49_), .Y(men_men_n300_));
  OAI210     u0272(.A0(men_men_n273_), .A1(men_men_n296_), .B0(men_men_n300_), .Y(men_men_n301_));
  NAi21      u0273(.An(l), .B(k), .Y(men_men_n302_));
  NO2        u0274(.A(men_men_n302_), .B(men_men_n49_), .Y(men_men_n303_));
  NOi21      u0275(.An(l), .B(j), .Y(men_men_n304_));
  NA2        u0276(.A(men_men_n169_), .B(men_men_n304_), .Y(men_men_n305_));
  NA3        u0277(.A(men_men_n121_), .B(men_men_n120_), .C(g), .Y(men_men_n306_));
  OR3        u0278(.A(men_men_n72_), .B(men_men_n74_), .C(e), .Y(men_men_n307_));
  AOI210     u0279(.A0(men_men_n306_), .A1(men_men_n305_), .B0(men_men_n307_), .Y(men_men_n308_));
  INV        u0280(.A(men_men_n308_), .Y(men_men_n309_));
  NAi32      u0281(.An(j), .Bn(h), .C(i), .Y(men_men_n310_));
  NAi21      u0282(.An(m), .B(l), .Y(men_men_n311_));
  NO3        u0283(.A(men_men_n311_), .B(men_men_n310_), .C(men_men_n85_), .Y(men_men_n312_));
  NA2        u0284(.A(h), .B(g), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n175_), .B(men_men_n45_), .Y(men_men_n314_));
  NO2        u0286(.A(men_men_n314_), .B(men_men_n313_), .Y(men_men_n315_));
  OAI210     u0287(.A0(men_men_n315_), .A1(men_men_n312_), .B0(men_men_n170_), .Y(men_men_n316_));
  NA4        u0288(.A(men_men_n316_), .B(men_men_n309_), .C(men_men_n301_), .D(men_men_n294_), .Y(men_men_n317_));
  NO2        u0289(.A(men_men_n150_), .B(d), .Y(men_men_n318_));
  NA2        u0290(.A(men_men_n318_), .B(men_men_n53_), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n108_), .B(men_men_n105_), .Y(men_men_n320_));
  NAi32      u0292(.An(n), .Bn(m), .C(l), .Y(men_men_n321_));
  NO2        u0293(.A(men_men_n321_), .B(men_men_n310_), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n125_), .B(men_men_n119_), .Y(men_men_n323_));
  NAi31      u0295(.An(k), .B(l), .C(j), .Y(men_men_n324_));
  OAI210     u0296(.A0(men_men_n302_), .A1(j), .B0(men_men_n324_), .Y(men_men_n325_));
  NOi21      u0297(.An(men_men_n325_), .B(men_men_n123_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n326_), .B(men_men_n323_), .Y(men_men_n327_));
  NA3        u0299(.A(men_men_n327_), .B(men_men_n1627_), .C(men_men_n319_), .Y(men_men_n328_));
  NO4        u0300(.A(men_men_n328_), .B(men_men_n317_), .C(men_men_n290_), .D(men_men_n280_), .Y(men_men_n329_));
  NA2        u0301(.A(men_men_n263_), .B(men_men_n199_), .Y(men_men_n330_));
  NAi21      u0302(.An(m), .B(k), .Y(men_men_n331_));
  NO2        u0303(.A(men_men_n232_), .B(men_men_n331_), .Y(men_men_n332_));
  NAi41      u0304(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n333_));
  NO2        u0305(.A(men_men_n333_), .B(men_men_n156_), .Y(men_men_n334_));
  NA2        u0306(.A(men_men_n334_), .B(men_men_n332_), .Y(men_men_n335_));
  NAi31      u0307(.An(i), .B(l), .C(h), .Y(men_men_n336_));
  NO4        u0308(.A(men_men_n336_), .B(men_men_n156_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n337_));
  NA2        u0309(.A(e), .B(c), .Y(men_men_n338_));
  NO3        u0310(.A(men_men_n338_), .B(n), .C(d), .Y(men_men_n339_));
  NOi21      u0311(.An(f), .B(h), .Y(men_men_n340_));
  NA2        u0312(.A(men_men_n340_), .B(men_men_n121_), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n341_), .B(men_men_n221_), .Y(men_men_n342_));
  NAi31      u0314(.An(d), .B(e), .C(b), .Y(men_men_n343_));
  NO2        u0315(.A(men_men_n136_), .B(men_men_n343_), .Y(men_men_n344_));
  NA2        u0316(.A(men_men_n344_), .B(men_men_n342_), .Y(men_men_n345_));
  NAi41      u0317(.An(men_men_n337_), .B(men_men_n345_), .C(men_men_n335_), .D(men_men_n330_), .Y(men_men_n346_));
  NO4        u0318(.A(men_men_n333_), .B(men_men_n80_), .C(men_men_n71_), .D(men_men_n221_), .Y(men_men_n347_));
  NA2        u0319(.A(men_men_n258_), .B(men_men_n106_), .Y(men_men_n348_));
  OR2        u0320(.A(men_men_n348_), .B(men_men_n210_), .Y(men_men_n349_));
  NOi31      u0321(.An(l), .B(n), .C(m), .Y(men_men_n350_));
  NA2        u0322(.A(men_men_n350_), .B(men_men_n222_), .Y(men_men_n351_));
  NO2        u0323(.A(men_men_n351_), .B(men_men_n1626_), .Y(men_men_n352_));
  NAi32      u0324(.An(men_men_n352_), .Bn(men_men_n347_), .C(men_men_n349_), .Y(men_men_n353_));
  NAi32      u0325(.An(m), .Bn(j), .C(k), .Y(men_men_n354_));
  NAi41      u0326(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n355_));
  OAI210     u0327(.A0(men_men_n218_), .A1(men_men_n354_), .B0(men_men_n355_), .Y(men_men_n356_));
  NOi31      u0328(.An(j), .B(m), .C(k), .Y(men_men_n357_));
  NO2        u0329(.A(men_men_n129_), .B(men_men_n357_), .Y(men_men_n358_));
  AN3        u0330(.A(h), .B(g), .C(f), .Y(men_men_n359_));
  NAi31      u0331(.An(men_men_n358_), .B(men_men_n359_), .C(men_men_n356_), .Y(men_men_n360_));
  NOi32      u0332(.An(m), .Bn(j), .C(l), .Y(men_men_n361_));
  NO2        u0333(.A(men_men_n361_), .B(men_men_n99_), .Y(men_men_n362_));
  NAi32      u0334(.An(men_men_n362_), .Bn(men_men_n207_), .C(men_men_n318_), .Y(men_men_n363_));
  NO2        u0335(.A(men_men_n311_), .B(men_men_n310_), .Y(men_men_n364_));
  NO2        u0336(.A(men_men_n224_), .B(g), .Y(men_men_n365_));
  NO2        u0337(.A(men_men_n162_), .B(men_men_n85_), .Y(men_men_n366_));
  AOI220     u0338(.A0(men_men_n366_), .A1(men_men_n365_), .B0(men_men_n255_), .B1(men_men_n364_), .Y(men_men_n367_));
  NA2        u0339(.A(men_men_n240_), .B(men_men_n80_), .Y(men_men_n368_));
  NA3        u0340(.A(men_men_n368_), .B(men_men_n359_), .C(men_men_n219_), .Y(men_men_n369_));
  NA4        u0341(.A(men_men_n369_), .B(men_men_n367_), .C(men_men_n363_), .D(men_men_n360_), .Y(men_men_n370_));
  NA3        u0342(.A(h), .B(g), .C(f), .Y(men_men_n371_));
  NO2        u0343(.A(men_men_n371_), .B(men_men_n76_), .Y(men_men_n372_));
  NA2        u0344(.A(men_men_n355_), .B(men_men_n218_), .Y(men_men_n373_));
  NA2        u0345(.A(men_men_n169_), .B(e), .Y(men_men_n374_));
  NO2        u0346(.A(men_men_n374_), .B(men_men_n41_), .Y(men_men_n375_));
  AOI220     u0347(.A0(men_men_n375_), .A1(men_men_n323_), .B0(men_men_n373_), .B1(men_men_n372_), .Y(men_men_n376_));
  NOi32      u0348(.An(j), .Bn(g), .C(i), .Y(men_men_n377_));
  NA3        u0349(.A(men_men_n377_), .B(men_men_n302_), .C(men_men_n116_), .Y(men_men_n378_));
  AO210      u0350(.A0(men_men_n114_), .A1(men_men_n32_), .B0(men_men_n378_), .Y(men_men_n379_));
  NOi32      u0351(.An(e), .Bn(b), .C(a), .Y(men_men_n380_));
  AN2        u0352(.A(l), .B(j), .Y(men_men_n381_));
  NO2        u0353(.A(men_men_n331_), .B(men_men_n381_), .Y(men_men_n382_));
  NO3        u0354(.A(men_men_n333_), .B(men_men_n71_), .C(men_men_n221_), .Y(men_men_n383_));
  NA3        u0355(.A(men_men_n215_), .B(men_men_n213_), .C(men_men_n35_), .Y(men_men_n384_));
  AOI220     u0356(.A0(men_men_n384_), .A1(men_men_n380_), .B0(men_men_n383_), .B1(men_men_n382_), .Y(men_men_n385_));
  NO2        u0357(.A(men_men_n343_), .B(n), .Y(men_men_n386_));
  NA2        u0358(.A(men_men_n214_), .B(k), .Y(men_men_n387_));
  NA3        u0359(.A(m), .B(men_men_n115_), .C(men_men_n220_), .Y(men_men_n388_));
  NA4        u0360(.A(men_men_n209_), .B(men_men_n88_), .C(g), .D(men_men_n220_), .Y(men_men_n389_));
  OAI210     u0361(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n389_), .Y(men_men_n390_));
  NAi41      u0362(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n391_));
  NA2        u0363(.A(men_men_n51_), .B(men_men_n116_), .Y(men_men_n392_));
  NO2        u0364(.A(men_men_n392_), .B(men_men_n391_), .Y(men_men_n393_));
  AOI220     u0365(.A0(men_men_n393_), .A1(b), .B0(men_men_n390_), .B1(men_men_n386_), .Y(men_men_n394_));
  NA4        u0366(.A(men_men_n394_), .B(men_men_n385_), .C(men_men_n379_), .D(men_men_n376_), .Y(men_men_n395_));
  NO4        u0367(.A(men_men_n395_), .B(men_men_n370_), .C(men_men_n353_), .D(men_men_n346_), .Y(men_men_n396_));
  NA4        u0368(.A(men_men_n396_), .B(men_men_n329_), .C(men_men_n278_), .D(men_men_n205_), .Y(men10));
  NA3        u0369(.A(m), .B(k), .C(i), .Y(men_men_n398_));
  NO3        u0370(.A(men_men_n398_), .B(j), .C(men_men_n221_), .Y(men_men_n399_));
  NOi21      u0371(.An(e), .B(f), .Y(men_men_n400_));
  NO4        u0372(.A(men_men_n157_), .B(men_men_n400_), .C(n), .D(men_men_n113_), .Y(men_men_n401_));
  NAi31      u0373(.An(b), .B(f), .C(c), .Y(men_men_n402_));
  INV        u0374(.A(men_men_n402_), .Y(men_men_n403_));
  NOi32      u0375(.An(k), .Bn(h), .C(j), .Y(men_men_n404_));
  NA2        u0376(.A(men_men_n404_), .B(men_men_n228_), .Y(men_men_n405_));
  NA2        u0377(.A(men_men_n167_), .B(men_men_n405_), .Y(men_men_n406_));
  AOI220     u0378(.A0(men_men_n406_), .A1(men_men_n403_), .B0(men_men_n401_), .B1(men_men_n399_), .Y(men_men_n407_));
  NO3        u0379(.A(n), .B(m), .C(k), .Y(men_men_n408_));
  NA2        u0380(.A(men_men_n408_), .B(j), .Y(men_men_n409_));
  NO3        u0381(.A(men_men_n409_), .B(men_men_n157_), .C(men_men_n220_), .Y(men_men_n410_));
  OR2        u0382(.A(m), .B(k), .Y(men_men_n411_));
  NO2        u0383(.A(men_men_n181_), .B(men_men_n411_), .Y(men_men_n412_));
  NA4        u0384(.A(n), .B(f), .C(c), .D(men_men_n119_), .Y(men_men_n413_));
  NOi21      u0385(.An(men_men_n412_), .B(men_men_n413_), .Y(men_men_n414_));
  NOi32      u0386(.An(d), .Bn(a), .C(c), .Y(men_men_n415_));
  NA2        u0387(.A(men_men_n415_), .B(men_men_n189_), .Y(men_men_n416_));
  NAi21      u0388(.An(i), .B(g), .Y(men_men_n417_));
  NAi31      u0389(.An(k), .B(m), .C(j), .Y(men_men_n418_));
  NO3        u0390(.A(men_men_n418_), .B(men_men_n417_), .C(n), .Y(men_men_n419_));
  NOi21      u0391(.An(men_men_n419_), .B(men_men_n416_), .Y(men_men_n420_));
  NO3        u0392(.A(men_men_n420_), .B(men_men_n414_), .C(men_men_n410_), .Y(men_men_n421_));
  NO2        u0393(.A(men_men_n413_), .B(men_men_n311_), .Y(men_men_n422_));
  NOi32      u0394(.An(f), .Bn(d), .C(c), .Y(men_men_n423_));
  AOI220     u0395(.A0(men_men_n423_), .A1(men_men_n322_), .B0(men_men_n422_), .B1(men_men_n222_), .Y(men_men_n424_));
  NA3        u0396(.A(men_men_n424_), .B(men_men_n421_), .C(men_men_n407_), .Y(men_men_n425_));
  NO2        u0397(.A(men_men_n59_), .B(men_men_n119_), .Y(men_men_n426_));
  NA2        u0398(.A(men_men_n258_), .B(men_men_n426_), .Y(men_men_n427_));
  INV        u0399(.A(e), .Y(men_men_n428_));
  NA2        u0400(.A(men_men_n46_), .B(e), .Y(men_men_n429_));
  OAI220     u0401(.A0(men_men_n429_), .A1(men_men_n206_), .B0(men_men_n210_), .B1(men_men_n428_), .Y(men_men_n430_));
  AN2        u0402(.A(g), .B(e), .Y(men_men_n431_));
  NA3        u0403(.A(men_men_n431_), .B(men_men_n209_), .C(i), .Y(men_men_n432_));
  OAI210     u0404(.A0(men_men_n90_), .A1(men_men_n428_), .B0(men_men_n432_), .Y(men_men_n433_));
  NO2        u0405(.A(men_men_n102_), .B(men_men_n428_), .Y(men_men_n434_));
  NO3        u0406(.A(men_men_n434_), .B(men_men_n433_), .C(men_men_n430_), .Y(men_men_n435_));
  NOi32      u0407(.An(h), .Bn(e), .C(g), .Y(men_men_n436_));
  NA3        u0408(.A(men_men_n436_), .B(men_men_n304_), .C(m), .Y(men_men_n437_));
  NOi21      u0409(.An(g), .B(h), .Y(men_men_n438_));
  AN3        u0410(.A(m), .B(l), .C(i), .Y(men_men_n439_));
  NA3        u0411(.A(men_men_n439_), .B(men_men_n438_), .C(e), .Y(men_men_n440_));
  AN3        u0412(.A(h), .B(g), .C(e), .Y(men_men_n441_));
  NA2        u0413(.A(men_men_n441_), .B(men_men_n99_), .Y(men_men_n442_));
  AN3        u0414(.A(men_men_n442_), .B(men_men_n440_), .C(men_men_n437_), .Y(men_men_n443_));
  AOI210     u0415(.A0(men_men_n443_), .A1(men_men_n435_), .B0(men_men_n427_), .Y(men_men_n444_));
  NA3        u0416(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n445_));
  NO2        u0417(.A(men_men_n445_), .B(men_men_n427_), .Y(men_men_n446_));
  NA3        u0418(.A(men_men_n415_), .B(men_men_n189_), .C(men_men_n85_), .Y(men_men_n447_));
  NAi31      u0419(.An(b), .B(c), .C(a), .Y(men_men_n448_));
  NO2        u0420(.A(men_men_n448_), .B(n), .Y(men_men_n449_));
  OAI210     u0421(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n450_));
  NO2        u0422(.A(men_men_n450_), .B(men_men_n153_), .Y(men_men_n451_));
  NA2        u0423(.A(men_men_n451_), .B(men_men_n449_), .Y(men_men_n452_));
  INV        u0424(.A(men_men_n452_), .Y(men_men_n453_));
  NO4        u0425(.A(men_men_n453_), .B(men_men_n446_), .C(men_men_n444_), .D(men_men_n425_), .Y(men_men_n454_));
  NA2        u0426(.A(i), .B(g), .Y(men_men_n455_));
  NO3        u0427(.A(men_men_n288_), .B(men_men_n455_), .C(c), .Y(men_men_n456_));
  NOi21      u0428(.An(d), .B(c), .Y(men_men_n457_));
  NA2        u0429(.A(men_men_n457_), .B(a), .Y(men_men_n458_));
  NA3        u0430(.A(i), .B(g), .C(f), .Y(men_men_n459_));
  OR2        u0431(.A(men_men_n459_), .B(men_men_n70_), .Y(men_men_n460_));
  NA3        u0432(.A(men_men_n439_), .B(men_men_n438_), .C(men_men_n189_), .Y(men_men_n461_));
  AOI210     u0433(.A0(men_men_n461_), .A1(men_men_n460_), .B0(men_men_n458_), .Y(men_men_n462_));
  AOI210     u0434(.A0(men_men_n456_), .A1(men_men_n303_), .B0(men_men_n462_), .Y(men_men_n463_));
  OR2        u0435(.A(n), .B(m), .Y(men_men_n464_));
  NO2        u0436(.A(men_men_n464_), .B(men_men_n158_), .Y(men_men_n465_));
  OAI210     u0437(.A0(men_men_n465_), .A1(men_men_n183_), .B0(d), .Y(men_men_n466_));
  INV        u0438(.A(men_men_n392_), .Y(men_men_n467_));
  NA3        u0439(.A(men_men_n467_), .B(men_men_n380_), .C(d), .Y(men_men_n468_));
  NO2        u0440(.A(men_men_n448_), .B(men_men_n49_), .Y(men_men_n469_));
  NO3        u0441(.A(men_men_n65_), .B(men_men_n115_), .C(e), .Y(men_men_n470_));
  NAi21      u0442(.An(k), .B(j), .Y(men_men_n471_));
  NA2        u0443(.A(men_men_n261_), .B(men_men_n471_), .Y(men_men_n472_));
  NA3        u0444(.A(men_men_n472_), .B(men_men_n470_), .C(men_men_n469_), .Y(men_men_n473_));
  NAi21      u0445(.An(e), .B(d), .Y(men_men_n474_));
  NO2        u0446(.A(men_men_n262_), .B(men_men_n220_), .Y(men_men_n475_));
  NA3        u0447(.A(men_men_n475_), .B(d), .C(men_men_n233_), .Y(men_men_n476_));
  NA4        u0448(.A(men_men_n476_), .B(men_men_n473_), .C(men_men_n468_), .D(men_men_n466_), .Y(men_men_n477_));
  NO2        u0449(.A(men_men_n351_), .B(men_men_n220_), .Y(men_men_n478_));
  NOi31      u0450(.An(n), .B(m), .C(k), .Y(men_men_n479_));
  AOI220     u0451(.A0(men_men_n479_), .A1(j), .B0(men_men_n228_), .B1(men_men_n50_), .Y(men_men_n480_));
  NAi31      u0452(.An(g), .B(f), .C(c), .Y(men_men_n481_));
  OR3        u0453(.A(men_men_n481_), .B(men_men_n480_), .C(e), .Y(men_men_n482_));
  NA3        u0454(.A(men_men_n482_), .B(men_men_n351_), .C(men_men_n1627_), .Y(men_men_n483_));
  NOi41      u0455(.An(men_men_n463_), .B(men_men_n483_), .C(men_men_n477_), .D(men_men_n276_), .Y(men_men_n484_));
  NOi32      u0456(.An(c), .Bn(a), .C(b), .Y(men_men_n485_));
  NA2        u0457(.A(men_men_n485_), .B(men_men_n116_), .Y(men_men_n486_));
  NA2        u0458(.A(men_men_n286_), .B(men_men_n158_), .Y(men_men_n487_));
  AN2        u0459(.A(e), .B(d), .Y(men_men_n488_));
  NA2        u0460(.A(men_men_n488_), .B(men_men_n487_), .Y(men_men_n489_));
  INV        u0461(.A(men_men_n153_), .Y(men_men_n490_));
  NO2        u0462(.A(men_men_n135_), .B(men_men_n41_), .Y(men_men_n491_));
  NO2        u0463(.A(men_men_n65_), .B(e), .Y(men_men_n492_));
  NOi31      u0464(.An(j), .B(k), .C(i), .Y(men_men_n493_));
  NOi21      u0465(.An(men_men_n172_), .B(men_men_n493_), .Y(men_men_n494_));
  NA4        u0466(.A(men_men_n336_), .B(men_men_n494_), .C(men_men_n270_), .D(men_men_n122_), .Y(men_men_n495_));
  AOI220     u0467(.A0(men_men_n495_), .A1(men_men_n492_), .B0(men_men_n491_), .B1(men_men_n490_), .Y(men_men_n496_));
  AOI210     u0468(.A0(men_men_n496_), .A1(men_men_n489_), .B0(men_men_n486_), .Y(men_men_n497_));
  NO2        u0469(.A(men_men_n216_), .B(men_men_n211_), .Y(men_men_n498_));
  NOi21      u0470(.An(a), .B(b), .Y(men_men_n499_));
  NA3        u0471(.A(e), .B(d), .C(c), .Y(men_men_n500_));
  NAi21      u0472(.An(men_men_n500_), .B(men_men_n499_), .Y(men_men_n501_));
  NO2        u0473(.A(men_men_n447_), .B(men_men_n210_), .Y(men_men_n502_));
  NOi21      u0474(.An(men_men_n501_), .B(men_men_n502_), .Y(men_men_n503_));
  AOI210     u0475(.A0(men_men_n279_), .A1(men_men_n498_), .B0(men_men_n503_), .Y(men_men_n504_));
  NO4        u0476(.A(men_men_n195_), .B(men_men_n105_), .C(men_men_n56_), .D(b), .Y(men_men_n505_));
  NA2        u0477(.A(men_men_n403_), .B(men_men_n159_), .Y(men_men_n506_));
  OR2        u0478(.A(k), .B(j), .Y(men_men_n507_));
  NA2        u0479(.A(l), .B(k), .Y(men_men_n508_));
  NA3        u0480(.A(men_men_n508_), .B(men_men_n507_), .C(men_men_n228_), .Y(men_men_n509_));
  AOI210     u0481(.A0(men_men_n240_), .A1(men_men_n354_), .B0(men_men_n85_), .Y(men_men_n510_));
  NOi21      u0482(.An(men_men_n509_), .B(men_men_n510_), .Y(men_men_n511_));
  OR3        u0483(.A(men_men_n511_), .B(men_men_n149_), .C(men_men_n139_), .Y(men_men_n512_));
  NA3        u0484(.A(men_men_n291_), .B(men_men_n132_), .C(men_men_n130_), .Y(men_men_n513_));
  NA2        u0485(.A(men_men_n415_), .B(men_men_n116_), .Y(men_men_n514_));
  NO4        u0486(.A(men_men_n514_), .B(men_men_n96_), .C(men_men_n115_), .D(e), .Y(men_men_n515_));
  NO3        u0487(.A(men_men_n447_), .B(men_men_n93_), .C(men_men_n135_), .Y(men_men_n516_));
  NO4        u0488(.A(men_men_n516_), .B(men_men_n515_), .C(men_men_n513_), .D(men_men_n337_), .Y(men_men_n517_));
  NA3        u0489(.A(men_men_n517_), .B(men_men_n512_), .C(men_men_n506_), .Y(men_men_n518_));
  NO4        u0490(.A(men_men_n518_), .B(men_men_n505_), .C(men_men_n504_), .D(men_men_n497_), .Y(men_men_n519_));
  NA2        u0491(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n520_));
  NOi21      u0492(.An(d), .B(e), .Y(men_men_n521_));
  NO2        u0493(.A(men_men_n195_), .B(men_men_n56_), .Y(men_men_n522_));
  OAI210     u0494(.A0(j), .A1(men_men_n136_), .B0(men_men_n105_), .Y(men_men_n523_));
  NA4        u0495(.A(men_men_n523_), .B(men_men_n522_), .C(men_men_n521_), .D(b), .Y(men_men_n524_));
  NO3        u0496(.A(men_men_n416_), .B(men_men_n362_), .C(men_men_n207_), .Y(men_men_n525_));
  NO2        u0497(.A(men_men_n416_), .B(men_men_n392_), .Y(men_men_n526_));
  NO4        u0498(.A(men_men_n526_), .B(men_men_n525_), .C(men_men_n191_), .D(men_men_n320_), .Y(men_men_n527_));
  NA4        u0499(.A(men_men_n527_), .B(men_men_n524_), .C(men_men_n520_), .D(men_men_n250_), .Y(men_men_n528_));
  OAI210     u0500(.A0(men_men_n131_), .A1(men_men_n129_), .B0(n), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n529_), .B(men_men_n135_), .Y(men_men_n530_));
  AO210      u0502(.A0(men_men_n312_), .A1(men_men_n221_), .B0(men_men_n252_), .Y(men_men_n531_));
  OA210      u0503(.A0(men_men_n531_), .A1(men_men_n530_), .B0(men_men_n199_), .Y(men_men_n532_));
  XO2        u0504(.A(i), .B(h), .Y(men_men_n533_));
  NA3        u0505(.A(men_men_n533_), .B(men_men_n166_), .C(n), .Y(men_men_n534_));
  NAi41      u0506(.An(men_men_n312_), .B(men_men_n534_), .C(men_men_n480_), .D(men_men_n405_), .Y(men_men_n535_));
  NOi32      u0507(.An(men_men_n535_), .Bn(men_men_n492_), .C(men_men_n281_), .Y(men_men_n536_));
  NAi31      u0508(.An(c), .B(f), .C(d), .Y(men_men_n537_));
  AOI210     u0509(.A0(men_men_n292_), .A1(men_men_n201_), .B0(men_men_n537_), .Y(men_men_n538_));
  NOi21      u0510(.An(men_men_n83_), .B(men_men_n538_), .Y(men_men_n539_));
  NA3        u0511(.A(men_men_n401_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n540_));
  NA2        u0512(.A(men_men_n234_), .B(men_men_n111_), .Y(men_men_n541_));
  AOI210     u0513(.A0(men_men_n541_), .A1(men_men_n188_), .B0(men_men_n537_), .Y(men_men_n542_));
  AOI210     u0514(.A0(men_men_n378_), .A1(men_men_n35_), .B0(men_men_n501_), .Y(men_men_n543_));
  NOi31      u0515(.An(men_men_n540_), .B(men_men_n543_), .C(men_men_n542_), .Y(men_men_n544_));
  AO220      u0516(.A0(men_men_n300_), .A1(men_men_n273_), .B0(men_men_n173_), .B1(men_men_n66_), .Y(men_men_n545_));
  NA3        u0517(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n546_));
  NO2        u0518(.A(men_men_n546_), .B(men_men_n458_), .Y(men_men_n547_));
  NO2        u0519(.A(men_men_n547_), .B(men_men_n308_), .Y(men_men_n548_));
  NAi41      u0520(.An(men_men_n545_), .B(men_men_n548_), .C(men_men_n544_), .D(men_men_n539_), .Y(men_men_n549_));
  NO4        u0521(.A(men_men_n549_), .B(men_men_n536_), .C(men_men_n532_), .D(men_men_n528_), .Y(men_men_n550_));
  NA4        u0522(.A(men_men_n550_), .B(men_men_n519_), .C(men_men_n484_), .D(men_men_n454_), .Y(men11));
  NO2        u0523(.A(men_men_n72_), .B(f), .Y(men_men_n552_));
  NA2        u0524(.A(j), .B(g), .Y(men_men_n553_));
  NAi31      u0525(.An(i), .B(m), .C(l), .Y(men_men_n554_));
  NA3        u0526(.A(m), .B(k), .C(j), .Y(men_men_n555_));
  OAI220     u0527(.A0(men_men_n555_), .A1(men_men_n135_), .B0(men_men_n554_), .B1(men_men_n553_), .Y(men_men_n556_));
  NA2        u0528(.A(men_men_n556_), .B(men_men_n552_), .Y(men_men_n557_));
  NOi32      u0529(.An(e), .Bn(b), .C(f), .Y(men_men_n558_));
  NA2        u0530(.A(men_men_n269_), .B(men_men_n116_), .Y(men_men_n559_));
  NA2        u0531(.A(men_men_n46_), .B(j), .Y(men_men_n560_));
  OAI220     u0532(.A0(men_men_n560_), .A1(men_men_n314_), .B0(men_men_n559_), .B1(men_men_n221_), .Y(men_men_n561_));
  NAi31      u0533(.An(d), .B(e), .C(a), .Y(men_men_n562_));
  NO2        u0534(.A(men_men_n562_), .B(n), .Y(men_men_n563_));
  AOI220     u0535(.A0(men_men_n563_), .A1(men_men_n103_), .B0(men_men_n561_), .B1(men_men_n558_), .Y(men_men_n564_));
  NAi41      u0536(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n565_));
  AN2        u0537(.A(men_men_n565_), .B(men_men_n391_), .Y(men_men_n566_));
  AOI210     u0538(.A0(men_men_n566_), .A1(men_men_n416_), .B0(men_men_n282_), .Y(men_men_n567_));
  NA2        u0539(.A(j), .B(i), .Y(men_men_n568_));
  NAi31      u0540(.An(n), .B(m), .C(k), .Y(men_men_n569_));
  NO3        u0541(.A(men_men_n569_), .B(men_men_n568_), .C(men_men_n115_), .Y(men_men_n570_));
  NO4        u0542(.A(n), .B(d), .C(men_men_n119_), .D(a), .Y(men_men_n571_));
  NO2        u0543(.A(c), .B(men_men_n155_), .Y(men_men_n572_));
  NO2        u0544(.A(men_men_n572_), .B(men_men_n571_), .Y(men_men_n573_));
  NOi32      u0545(.An(g), .Bn(f), .C(i), .Y(men_men_n574_));
  AOI220     u0546(.A0(men_men_n574_), .A1(men_men_n101_), .B0(men_men_n556_), .B1(f), .Y(men_men_n575_));
  NO2        u0547(.A(men_men_n286_), .B(men_men_n49_), .Y(men_men_n576_));
  NO2        u0548(.A(men_men_n575_), .B(men_men_n573_), .Y(men_men_n577_));
  AOI210     u0549(.A0(men_men_n570_), .A1(men_men_n567_), .B0(men_men_n577_), .Y(men_men_n578_));
  NA2        u0550(.A(men_men_n145_), .B(men_men_n34_), .Y(men_men_n579_));
  OAI220     u0551(.A0(men_men_n579_), .A1(m), .B0(men_men_n560_), .B1(men_men_n240_), .Y(men_men_n580_));
  NOi41      u0552(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n581_));
  NAi32      u0553(.An(e), .Bn(b), .C(c), .Y(men_men_n582_));
  OR2        u0554(.A(men_men_n582_), .B(men_men_n85_), .Y(men_men_n583_));
  AN2        u0555(.A(men_men_n355_), .B(men_men_n333_), .Y(men_men_n584_));
  NA2        u0556(.A(men_men_n584_), .B(men_men_n583_), .Y(men_men_n585_));
  OA210      u0557(.A0(men_men_n585_), .A1(men_men_n581_), .B0(men_men_n580_), .Y(men_men_n586_));
  OAI220     u0558(.A0(men_men_n418_), .A1(men_men_n417_), .B0(men_men_n554_), .B1(men_men_n553_), .Y(men_men_n587_));
  NAi31      u0559(.An(d), .B(c), .C(a), .Y(men_men_n588_));
  NO2        u0560(.A(men_men_n588_), .B(n), .Y(men_men_n589_));
  NA3        u0561(.A(men_men_n589_), .B(men_men_n587_), .C(e), .Y(men_men_n590_));
  NO3        u0562(.A(men_men_n61_), .B(men_men_n49_), .C(men_men_n221_), .Y(men_men_n591_));
  NO2        u0563(.A(men_men_n237_), .B(men_men_n113_), .Y(men_men_n592_));
  OAI210     u0564(.A0(men_men_n591_), .A1(men_men_n419_), .B0(men_men_n592_), .Y(men_men_n593_));
  NA2        u0565(.A(men_men_n593_), .B(men_men_n590_), .Y(men_men_n594_));
  NO2        u0566(.A(men_men_n288_), .B(n), .Y(men_men_n595_));
  NO2        u0567(.A(men_men_n449_), .B(men_men_n595_), .Y(men_men_n596_));
  NA2        u0568(.A(men_men_n587_), .B(f), .Y(men_men_n597_));
  NAi32      u0569(.An(d), .Bn(a), .C(b), .Y(men_men_n598_));
  NO2        u0570(.A(men_men_n598_), .B(men_men_n49_), .Y(men_men_n599_));
  NA2        u0571(.A(h), .B(f), .Y(men_men_n600_));
  NO2        u0572(.A(men_men_n600_), .B(men_men_n96_), .Y(men_men_n601_));
  NO3        u0573(.A(men_men_n184_), .B(men_men_n181_), .C(g), .Y(men_men_n602_));
  AOI220     u0574(.A0(men_men_n602_), .A1(men_men_n58_), .B0(men_men_n601_), .B1(men_men_n599_), .Y(men_men_n603_));
  OAI210     u0575(.A0(men_men_n597_), .A1(men_men_n596_), .B0(men_men_n603_), .Y(men_men_n604_));
  AN3        u0576(.A(j), .B(h), .C(g), .Y(men_men_n605_));
  NO2        u0577(.A(men_men_n152_), .B(c), .Y(men_men_n606_));
  NA3        u0578(.A(men_men_n606_), .B(men_men_n605_), .C(men_men_n479_), .Y(men_men_n607_));
  NA3        u0579(.A(f), .B(d), .C(b), .Y(men_men_n608_));
  NO4        u0580(.A(men_men_n608_), .B(men_men_n184_), .C(men_men_n181_), .D(g), .Y(men_men_n609_));
  NAi21      u0581(.An(men_men_n609_), .B(men_men_n607_), .Y(men_men_n610_));
  NO4        u0582(.A(men_men_n610_), .B(men_men_n604_), .C(men_men_n594_), .D(men_men_n586_), .Y(men_men_n611_));
  AN4        u0583(.A(men_men_n611_), .B(men_men_n578_), .C(men_men_n564_), .D(men_men_n557_), .Y(men_men_n612_));
  INV        u0584(.A(k), .Y(men_men_n613_));
  NA3        u0585(.A(l), .B(men_men_n613_), .C(i), .Y(men_men_n614_));
  INV        u0586(.A(men_men_n614_), .Y(men_men_n615_));
  NA4        u0587(.A(men_men_n415_), .B(men_men_n438_), .C(men_men_n189_), .D(men_men_n116_), .Y(men_men_n616_));
  NAi32      u0588(.An(h), .Bn(f), .C(g), .Y(men_men_n617_));
  NAi41      u0589(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n618_));
  OAI210     u0590(.A0(men_men_n562_), .A1(n), .B0(men_men_n618_), .Y(men_men_n619_));
  NA2        u0591(.A(men_men_n619_), .B(m), .Y(men_men_n620_));
  NAi31      u0592(.An(h), .B(g), .C(f), .Y(men_men_n621_));
  OR3        u0593(.A(men_men_n621_), .B(men_men_n288_), .C(men_men_n49_), .Y(men_men_n622_));
  NA4        u0594(.A(men_men_n438_), .B(men_men_n124_), .C(men_men_n116_), .D(e), .Y(men_men_n623_));
  AN2        u0595(.A(men_men_n623_), .B(men_men_n622_), .Y(men_men_n624_));
  OA210      u0596(.A0(men_men_n620_), .A1(men_men_n617_), .B0(men_men_n624_), .Y(men_men_n625_));
  NO3        u0597(.A(men_men_n617_), .B(men_men_n72_), .C(men_men_n74_), .Y(men_men_n626_));
  NO4        u0598(.A(men_men_n621_), .B(c), .C(men_men_n155_), .D(men_men_n74_), .Y(men_men_n627_));
  OR2        u0599(.A(men_men_n627_), .B(men_men_n626_), .Y(men_men_n628_));
  NAi31      u0600(.An(men_men_n628_), .B(men_men_n625_), .C(men_men_n616_), .Y(men_men_n629_));
  NAi31      u0601(.An(f), .B(h), .C(g), .Y(men_men_n630_));
  NO4        u0602(.A(men_men_n324_), .B(men_men_n630_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n631_));
  NOi32      u0603(.An(b), .Bn(a), .C(c), .Y(men_men_n632_));
  NOi41      u0604(.An(men_men_n632_), .B(men_men_n371_), .C(men_men_n68_), .D(men_men_n120_), .Y(men_men_n633_));
  OR2        u0605(.A(men_men_n633_), .B(men_men_n631_), .Y(men_men_n634_));
  NOi32      u0606(.An(d), .Bn(a), .C(e), .Y(men_men_n635_));
  NA2        u0607(.A(men_men_n635_), .B(men_men_n116_), .Y(men_men_n636_));
  NO2        u0608(.A(n), .B(c), .Y(men_men_n637_));
  NA3        u0609(.A(men_men_n637_), .B(men_men_n29_), .C(m), .Y(men_men_n638_));
  NAi32      u0610(.An(n), .Bn(f), .C(m), .Y(men_men_n639_));
  NA3        u0611(.A(men_men_n639_), .B(men_men_n638_), .C(men_men_n636_), .Y(men_men_n640_));
  NOi32      u0612(.An(e), .Bn(a), .C(d), .Y(men_men_n641_));
  AOI210     u0613(.A0(men_men_n29_), .A1(d), .B0(men_men_n641_), .Y(men_men_n642_));
  AOI210     u0614(.A0(men_men_n642_), .A1(men_men_n220_), .B0(men_men_n579_), .Y(men_men_n643_));
  AOI210     u0615(.A0(men_men_n643_), .A1(men_men_n640_), .B0(men_men_n634_), .Y(men_men_n644_));
  OAI210     u0616(.A0(men_men_n257_), .A1(men_men_n88_), .B0(men_men_n644_), .Y(men_men_n645_));
  AOI210     u0617(.A0(men_men_n629_), .A1(men_men_n615_), .B0(men_men_n645_), .Y(men_men_n646_));
  NO3        u0618(.A(men_men_n331_), .B(men_men_n60_), .C(n), .Y(men_men_n647_));
  NA2        u0619(.A(men_men_n481_), .B(men_men_n237_), .Y(men_men_n648_));
  OR2        u0620(.A(men_men_n648_), .B(f), .Y(men_men_n649_));
  NA2        u0621(.A(men_men_n75_), .B(men_men_n116_), .Y(men_men_n650_));
  NO2        u0622(.A(men_men_n650_), .B(men_men_n45_), .Y(men_men_n651_));
  AOI220     u0623(.A0(men_men_n651_), .A1(men_men_n567_), .B0(men_men_n649_), .B1(men_men_n647_), .Y(men_men_n652_));
  NO2        u0624(.A(men_men_n652_), .B(men_men_n88_), .Y(men_men_n653_));
  NA3        u0625(.A(men_men_n581_), .B(men_men_n357_), .C(men_men_n46_), .Y(men_men_n654_));
  NOi32      u0626(.An(e), .Bn(c), .C(f), .Y(men_men_n655_));
  NOi21      u0627(.An(f), .B(g), .Y(men_men_n656_));
  NO2        u0628(.A(men_men_n656_), .B(men_men_n218_), .Y(men_men_n657_));
  AOI220     u0629(.A0(men_men_n657_), .A1(men_men_n412_), .B0(men_men_n655_), .B1(men_men_n183_), .Y(men_men_n658_));
  NA3        u0630(.A(men_men_n658_), .B(men_men_n654_), .C(men_men_n186_), .Y(men_men_n659_));
  AOI210     u0631(.A0(men_men_n566_), .A1(men_men_n416_), .B0(men_men_n313_), .Y(men_men_n660_));
  NA2        u0632(.A(men_men_n660_), .B(men_men_n274_), .Y(men_men_n661_));
  NOi21      u0633(.An(j), .B(l), .Y(men_men_n662_));
  NAi21      u0634(.An(k), .B(h), .Y(men_men_n663_));
  NO2        u0635(.A(men_men_n663_), .B(men_men_n272_), .Y(men_men_n664_));
  NA2        u0636(.A(men_men_n664_), .B(men_men_n662_), .Y(men_men_n665_));
  OR2        u0637(.A(men_men_n665_), .B(men_men_n620_), .Y(men_men_n666_));
  NOi31      u0638(.An(m), .B(n), .C(k), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n662_), .B(men_men_n667_), .Y(men_men_n668_));
  AOI210     u0640(.A0(men_men_n416_), .A1(men_men_n391_), .B0(men_men_n313_), .Y(men_men_n669_));
  NAi21      u0641(.An(men_men_n668_), .B(men_men_n669_), .Y(men_men_n670_));
  NO2        u0642(.A(men_men_n288_), .B(men_men_n49_), .Y(men_men_n671_));
  NO2        u0643(.A(men_men_n324_), .B(men_men_n630_), .Y(men_men_n672_));
  NO2        u0644(.A(men_men_n562_), .B(men_men_n49_), .Y(men_men_n673_));
  AOI220     u0645(.A0(men_men_n673_), .A1(men_men_n672_), .B0(men_men_n671_), .B1(men_men_n601_), .Y(men_men_n674_));
  NA4        u0646(.A(men_men_n674_), .B(men_men_n670_), .C(men_men_n666_), .D(men_men_n661_), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n111_), .B(men_men_n36_), .Y(men_men_n676_));
  NO2        u0648(.A(k), .B(men_men_n221_), .Y(men_men_n677_));
  NO2        u0649(.A(men_men_n558_), .B(men_men_n380_), .Y(men_men_n678_));
  NAi31      u0650(.An(men_men_n676_), .B(men_men_n380_), .C(men_men_n677_), .Y(men_men_n679_));
  NO2        u0651(.A(men_men_n560_), .B(men_men_n184_), .Y(men_men_n680_));
  NA3        u0652(.A(men_men_n582_), .B(men_men_n281_), .C(men_men_n150_), .Y(men_men_n681_));
  NA2        u0653(.A(men_men_n533_), .B(men_men_n166_), .Y(men_men_n682_));
  NO3        u0654(.A(men_men_n413_), .B(men_men_n682_), .C(men_men_n88_), .Y(men_men_n683_));
  AOI210     u0655(.A0(men_men_n681_), .A1(men_men_n680_), .B0(men_men_n683_), .Y(men_men_n684_));
  OAI210     u0656(.A0(d), .A1(men_men_n134_), .B0(n), .Y(men_men_n685_));
  NA3        u0657(.A(men_men_n533_), .B(men_men_n166_), .C(men_men_n221_), .Y(men_men_n686_));
  AOI210     u0658(.A0(men_men_n685_), .A1(men_men_n239_), .B0(men_men_n686_), .Y(men_men_n687_));
  NAi31      u0659(.An(m), .B(n), .C(k), .Y(men_men_n688_));
  OR2        u0660(.A(men_men_n139_), .B(men_men_n60_), .Y(men_men_n689_));
  OAI210     u0661(.A0(men_men_n689_), .A1(men_men_n688_), .B0(men_men_n259_), .Y(men_men_n690_));
  OAI210     u0662(.A0(men_men_n690_), .A1(men_men_n687_), .B0(j), .Y(men_men_n691_));
  NA3        u0663(.A(men_men_n691_), .B(men_men_n684_), .C(men_men_n679_), .Y(men_men_n692_));
  NO4        u0664(.A(men_men_n692_), .B(men_men_n675_), .C(men_men_n659_), .D(men_men_n653_), .Y(men_men_n693_));
  NA2        u0665(.A(men_men_n401_), .B(men_men_n169_), .Y(men_men_n694_));
  NAi31      u0666(.An(g), .B(h), .C(f), .Y(men_men_n695_));
  OR3        u0667(.A(men_men_n695_), .B(men_men_n288_), .C(n), .Y(men_men_n696_));
  OA210      u0668(.A0(men_men_n562_), .A1(n), .B0(men_men_n618_), .Y(men_men_n697_));
  NA3        u0669(.A(men_men_n436_), .B(men_men_n124_), .C(men_men_n85_), .Y(men_men_n698_));
  OAI210     u0670(.A0(men_men_n697_), .A1(men_men_n92_), .B0(men_men_n698_), .Y(men_men_n699_));
  NOi21      u0671(.An(men_men_n696_), .B(men_men_n699_), .Y(men_men_n700_));
  AOI210     u0672(.A0(men_men_n700_), .A1(men_men_n694_), .B0(men_men_n555_), .Y(men_men_n701_));
  NO3        u0673(.A(g), .B(men_men_n220_), .C(men_men_n56_), .Y(men_men_n702_));
  NAi21      u0674(.An(h), .B(j), .Y(men_men_n703_));
  OAI210     u0675(.A0(men_men_n234_), .A1(men_men_n412_), .B0(men_men_n702_), .Y(men_men_n704_));
  OR2        u0676(.A(men_men_n72_), .B(men_men_n74_), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n632_), .B(men_men_n359_), .Y(men_men_n706_));
  OA220      u0678(.A0(men_men_n668_), .A1(men_men_n706_), .B0(men_men_n665_), .B1(men_men_n705_), .Y(men_men_n707_));
  NA3        u0679(.A(men_men_n552_), .B(men_men_n101_), .C(men_men_n100_), .Y(men_men_n708_));
  AN2        u0680(.A(h), .B(f), .Y(men_men_n709_));
  NA2        u0681(.A(men_men_n709_), .B(men_men_n37_), .Y(men_men_n710_));
  NA2        u0682(.A(men_men_n101_), .B(men_men_n46_), .Y(men_men_n711_));
  OAI220     u0683(.A0(men_men_n711_), .A1(men_men_n348_), .B0(men_men_n710_), .B1(men_men_n486_), .Y(men_men_n712_));
  AOI210     u0684(.A0(men_men_n598_), .A1(men_men_n448_), .B0(men_men_n49_), .Y(men_men_n713_));
  OAI220     u0685(.A0(men_men_n621_), .A1(men_men_n614_), .B0(men_men_n341_), .B1(men_men_n553_), .Y(men_men_n714_));
  AOI210     u0686(.A0(men_men_n714_), .A1(men_men_n713_), .B0(men_men_n712_), .Y(men_men_n715_));
  NA4        u0687(.A(men_men_n715_), .B(men_men_n708_), .C(men_men_n707_), .D(men_men_n704_), .Y(men_men_n716_));
  NO2        u0688(.A(men_men_n261_), .B(f), .Y(men_men_n717_));
  NO2        u0689(.A(men_men_n656_), .B(men_men_n60_), .Y(men_men_n718_));
  NO3        u0690(.A(men_men_n718_), .B(men_men_n717_), .C(men_men_n34_), .Y(men_men_n719_));
  NA2        u0691(.A(men_men_n344_), .B(men_men_n145_), .Y(men_men_n720_));
  AOI210     u0692(.A0(men_men_n380_), .A1(men_men_n116_), .B0(men_men_n558_), .Y(men_men_n721_));
  OA220      u0693(.A0(men_men_n721_), .A1(men_men_n579_), .B0(men_men_n378_), .B1(men_men_n114_), .Y(men_men_n722_));
  OAI210     u0694(.A0(men_men_n720_), .A1(men_men_n719_), .B0(men_men_n722_), .Y(men_men_n723_));
  NA2        u0695(.A(men_men_n1622_), .B(men_men_n237_), .Y(men_men_n724_));
  NA3        u0696(.A(men_men_n724_), .B(men_men_n263_), .C(j), .Y(men_men_n725_));
  NO3        u0697(.A(men_men_n481_), .B(men_men_n181_), .C(i), .Y(men_men_n726_));
  NA2        u0698(.A(men_men_n485_), .B(men_men_n85_), .Y(men_men_n727_));
  NO4        u0699(.A(men_men_n555_), .B(men_men_n727_), .C(men_men_n135_), .D(men_men_n220_), .Y(men_men_n728_));
  AOI210     u0700(.A0(men_men_n726_), .A1(men_men_n175_), .B0(men_men_n728_), .Y(men_men_n729_));
  NA4        u0701(.A(men_men_n729_), .B(men_men_n725_), .C(men_men_n540_), .D(men_men_n421_), .Y(men_men_n730_));
  NO4        u0702(.A(men_men_n730_), .B(men_men_n723_), .C(men_men_n716_), .D(men_men_n701_), .Y(men_men_n731_));
  NA4        u0703(.A(men_men_n731_), .B(men_men_n693_), .C(men_men_n646_), .D(men_men_n612_), .Y(men08));
  NO2        u0704(.A(k), .B(h), .Y(men_men_n733_));
  AO210      u0705(.A0(men_men_n261_), .A1(men_men_n471_), .B0(men_men_n733_), .Y(men_men_n734_));
  NO2        u0706(.A(men_men_n734_), .B(men_men_n311_), .Y(men_men_n735_));
  NA2        u0707(.A(men_men_n655_), .B(men_men_n85_), .Y(men_men_n736_));
  NA2        u0708(.A(men_men_n736_), .B(men_men_n481_), .Y(men_men_n737_));
  AOI210     u0709(.A0(men_men_n737_), .A1(men_men_n735_), .B0(men_men_n516_), .Y(men_men_n738_));
  NA2        u0710(.A(men_men_n85_), .B(men_men_n113_), .Y(men_men_n739_));
  NO2        u0711(.A(men_men_n739_), .B(men_men_n57_), .Y(men_men_n740_));
  NO4        u0712(.A(men_men_n398_), .B(men_men_n115_), .C(j), .D(men_men_n221_), .Y(men_men_n741_));
  OAI210     u0713(.A0(men_men_n608_), .A1(men_men_n85_), .B0(men_men_n239_), .Y(men_men_n742_));
  AOI220     u0714(.A0(men_men_n742_), .A1(men_men_n365_), .B0(men_men_n741_), .B1(men_men_n740_), .Y(men_men_n743_));
  AOI210     u0715(.A0(men_men_n608_), .A1(men_men_n162_), .B0(men_men_n85_), .Y(men_men_n744_));
  NA4        u0716(.A(men_men_n223_), .B(men_men_n145_), .C(men_men_n45_), .D(h), .Y(men_men_n745_));
  AN2        u0717(.A(l), .B(k), .Y(men_men_n746_));
  NA4        u0718(.A(men_men_n746_), .B(men_men_n111_), .C(men_men_n74_), .D(men_men_n221_), .Y(men_men_n747_));
  OAI210     u0719(.A0(men_men_n745_), .A1(g), .B0(men_men_n747_), .Y(men_men_n748_));
  NA2        u0720(.A(men_men_n748_), .B(men_men_n744_), .Y(men_men_n749_));
  NA4        u0721(.A(men_men_n749_), .B(men_men_n743_), .C(men_men_n738_), .D(men_men_n367_), .Y(men_men_n750_));
  AN2        u0722(.A(men_men_n563_), .B(men_men_n97_), .Y(men_men_n751_));
  NO4        u0723(.A(men_men_n181_), .B(men_men_n411_), .C(men_men_n115_), .D(g), .Y(men_men_n752_));
  AOI210     u0724(.A0(men_men_n752_), .A1(men_men_n742_), .B0(men_men_n547_), .Y(men_men_n753_));
  NO2        u0725(.A(men_men_n38_), .B(men_men_n220_), .Y(men_men_n754_));
  AOI220     u0726(.A0(men_men_n657_), .A1(men_men_n364_), .B0(men_men_n754_), .B1(men_men_n595_), .Y(men_men_n755_));
  NAi31      u0727(.An(men_men_n751_), .B(men_men_n755_), .C(men_men_n753_), .Y(men_men_n756_));
  NO2        u0728(.A(men_men_n566_), .B(men_men_n35_), .Y(men_men_n757_));
  OAI210     u0729(.A0(men_men_n582_), .A1(men_men_n47_), .B0(men_men_n689_), .Y(men_men_n758_));
  AOI210     u0730(.A0(men_men_n1631_), .A1(men_men_n758_), .B0(men_men_n757_), .Y(men_men_n759_));
  NO3        u0731(.A(men_men_n331_), .B(men_men_n135_), .C(men_men_n41_), .Y(men_men_n760_));
  NAi21      u0732(.An(men_men_n760_), .B(men_men_n747_), .Y(men_men_n761_));
  NA2        u0733(.A(men_men_n734_), .B(men_men_n140_), .Y(men_men_n762_));
  AOI220     u0734(.A0(men_men_n762_), .A1(men_men_n422_), .B0(men_men_n761_), .B1(men_men_n77_), .Y(men_men_n763_));
  OAI210     u0735(.A0(men_men_n759_), .A1(men_men_n88_), .B0(men_men_n763_), .Y(men_men_n764_));
  NA2        u0736(.A(men_men_n380_), .B(men_men_n43_), .Y(men_men_n765_));
  NA3        u0737(.A(men_men_n724_), .B(men_men_n350_), .C(men_men_n404_), .Y(men_men_n766_));
  NA2        u0738(.A(men_men_n746_), .B(men_men_n228_), .Y(men_men_n767_));
  NO2        u0739(.A(men_men_n767_), .B(men_men_n343_), .Y(men_men_n768_));
  AOI210     u0740(.A0(men_men_n768_), .A1(men_men_n717_), .B0(men_men_n515_), .Y(men_men_n769_));
  NA3        u0741(.A(m), .B(l), .C(k), .Y(men_men_n770_));
  AOI210     u0742(.A0(men_men_n698_), .A1(men_men_n696_), .B0(men_men_n770_), .Y(men_men_n771_));
  NO2        u0743(.A(men_men_n565_), .B(men_men_n282_), .Y(men_men_n772_));
  NOi21      u0744(.An(men_men_n772_), .B(men_men_n559_), .Y(men_men_n773_));
  NA4        u0745(.A(men_men_n116_), .B(l), .C(k), .D(men_men_n88_), .Y(men_men_n774_));
  NA3        u0746(.A(men_men_n124_), .B(men_men_n431_), .C(i), .Y(men_men_n775_));
  NO2        u0747(.A(men_men_n775_), .B(men_men_n774_), .Y(men_men_n776_));
  NO3        u0748(.A(men_men_n776_), .B(men_men_n773_), .C(men_men_n771_), .Y(men_men_n777_));
  NA4        u0749(.A(men_men_n777_), .B(men_men_n769_), .C(men_men_n766_), .D(men_men_n765_), .Y(men_men_n778_));
  NO4        u0750(.A(men_men_n778_), .B(men_men_n764_), .C(men_men_n756_), .D(men_men_n750_), .Y(men_men_n779_));
  NA2        u0751(.A(men_men_n657_), .B(men_men_n412_), .Y(men_men_n780_));
  NOi31      u0752(.An(g), .B(h), .C(f), .Y(men_men_n781_));
  NA2        u0753(.A(men_men_n673_), .B(men_men_n781_), .Y(men_men_n782_));
  AO210      u0754(.A0(men_men_n782_), .A1(men_men_n622_), .B0(men_men_n568_), .Y(men_men_n783_));
  NO3        u0755(.A(men_men_n416_), .B(men_men_n553_), .C(h), .Y(men_men_n784_));
  AOI210     u0756(.A0(men_men_n784_), .A1(men_men_n116_), .B0(men_men_n526_), .Y(men_men_n785_));
  NA4        u0757(.A(men_men_n785_), .B(men_men_n783_), .C(men_men_n780_), .D(men_men_n260_), .Y(men_men_n786_));
  NA2        u0758(.A(men_men_n746_), .B(men_men_n74_), .Y(men_men_n787_));
  NO3        u0759(.A(men_men_n181_), .B(n), .C(i), .Y(men_men_n788_));
  NOi21      u0760(.An(h), .B(j), .Y(men_men_n789_));
  NA2        u0761(.A(men_men_n789_), .B(f), .Y(men_men_n790_));
  NO2        u0762(.A(men_men_n790_), .B(men_men_n254_), .Y(men_men_n791_));
  NO3        u0763(.A(men_men_n791_), .B(men_men_n788_), .C(men_men_n726_), .Y(men_men_n792_));
  OAI220     u0764(.A0(men_men_n792_), .A1(men_men_n787_), .B0(men_men_n624_), .B1(men_men_n61_), .Y(men_men_n793_));
  AOI210     u0765(.A0(men_men_n786_), .A1(l), .B0(men_men_n793_), .Y(men_men_n794_));
  NO2        u0766(.A(j), .B(i), .Y(men_men_n795_));
  NA3        u0767(.A(men_men_n795_), .B(men_men_n81_), .C(l), .Y(men_men_n796_));
  NA2        u0768(.A(men_men_n795_), .B(men_men_n33_), .Y(men_men_n797_));
  NA2        u0769(.A(men_men_n441_), .B(men_men_n124_), .Y(men_men_n798_));
  OA220      u0770(.A0(men_men_n798_), .A1(men_men_n797_), .B0(men_men_n796_), .B1(men_men_n620_), .Y(men_men_n799_));
  NO3        u0771(.A(men_men_n157_), .B(men_men_n49_), .C(men_men_n113_), .Y(men_men_n800_));
  NO3        u0772(.A(c), .B(men_men_n155_), .C(men_men_n74_), .Y(men_men_n801_));
  NO3        u0773(.A(men_men_n508_), .B(men_men_n459_), .C(j), .Y(men_men_n802_));
  OAI210     u0774(.A0(men_men_n801_), .A1(men_men_n800_), .B0(men_men_n802_), .Y(men_men_n803_));
  OAI210     u0775(.A0(men_men_n782_), .A1(men_men_n61_), .B0(men_men_n803_), .Y(men_men_n804_));
  NA2        u0776(.A(k), .B(j), .Y(men_men_n805_));
  NO3        u0777(.A(men_men_n311_), .B(men_men_n805_), .C(men_men_n40_), .Y(men_men_n806_));
  AOI210     u0778(.A0(men_men_n558_), .A1(n), .B0(men_men_n581_), .Y(men_men_n807_));
  NA2        u0779(.A(men_men_n807_), .B(men_men_n584_), .Y(men_men_n808_));
  AN3        u0780(.A(men_men_n808_), .B(men_men_n806_), .C(men_men_n100_), .Y(men_men_n809_));
  NO3        u0781(.A(men_men_n181_), .B(men_men_n411_), .C(men_men_n115_), .Y(men_men_n810_));
  AOI220     u0782(.A0(men_men_n810_), .A1(men_men_n255_), .B0(men_men_n648_), .B1(men_men_n322_), .Y(men_men_n811_));
  NAi31      u0783(.An(men_men_n642_), .B(men_men_n94_), .C(men_men_n85_), .Y(men_men_n812_));
  NA2        u0784(.A(men_men_n812_), .B(men_men_n811_), .Y(men_men_n813_));
  NO2        u0785(.A(men_men_n311_), .B(men_men_n140_), .Y(men_men_n814_));
  AOI220     u0786(.A0(men_men_n814_), .A1(men_men_n657_), .B0(men_men_n760_), .B1(men_men_n744_), .Y(men_men_n815_));
  NO2        u0787(.A(men_men_n770_), .B(men_men_n92_), .Y(men_men_n816_));
  NA2        u0788(.A(men_men_n816_), .B(men_men_n619_), .Y(men_men_n817_));
  NO2        u0789(.A(men_men_n621_), .B(men_men_n120_), .Y(men_men_n818_));
  OAI210     u0790(.A0(men_men_n818_), .A1(men_men_n802_), .B0(men_men_n713_), .Y(men_men_n819_));
  NA3        u0791(.A(men_men_n819_), .B(men_men_n817_), .C(men_men_n815_), .Y(men_men_n820_));
  OR4        u0792(.A(men_men_n820_), .B(men_men_n813_), .C(men_men_n809_), .D(men_men_n804_), .Y(men_men_n821_));
  NA3        u0793(.A(men_men_n807_), .B(men_men_n584_), .C(men_men_n583_), .Y(men_men_n822_));
  NA4        u0794(.A(men_men_n822_), .B(men_men_n223_), .C(men_men_n471_), .D(men_men_n34_), .Y(men_men_n823_));
  NO4        u0795(.A(men_men_n508_), .B(men_men_n455_), .C(j), .D(f), .Y(men_men_n824_));
  OAI220     u0796(.A0(men_men_n745_), .A1(men_men_n736_), .B0(men_men_n348_), .B1(men_men_n38_), .Y(men_men_n825_));
  AOI210     u0797(.A0(men_men_n824_), .A1(men_men_n267_), .B0(men_men_n825_), .Y(men_men_n826_));
  NA3        u0798(.A(men_men_n574_), .B(men_men_n304_), .C(h), .Y(men_men_n827_));
  NOi21      u0799(.An(men_men_n713_), .B(men_men_n827_), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n93_), .B(men_men_n47_), .Y(men_men_n829_));
  OAI220     u0801(.A0(men_men_n827_), .A1(men_men_n638_), .B0(men_men_n796_), .B1(men_men_n705_), .Y(men_men_n830_));
  AOI210     u0802(.A0(men_men_n829_), .A1(men_men_n380_), .B0(men_men_n830_), .Y(men_men_n831_));
  NAi41      u0803(.An(men_men_n828_), .B(men_men_n831_), .C(men_men_n826_), .D(men_men_n823_), .Y(men_men_n832_));
  OR2        u0804(.A(men_men_n816_), .B(men_men_n97_), .Y(men_men_n833_));
  AOI220     u0805(.A0(men_men_n833_), .A1(men_men_n245_), .B0(men_men_n802_), .B1(men_men_n671_), .Y(men_men_n834_));
  NO2        u0806(.A(men_men_n697_), .B(men_men_n74_), .Y(men_men_n835_));
  AOI210     u0807(.A0(men_men_n824_), .A1(men_men_n835_), .B0(men_men_n352_), .Y(men_men_n836_));
  NA2        u0808(.A(men_men_n695_), .B(men_men_n546_), .Y(men_men_n837_));
  NA3        u0809(.A(men_men_n258_), .B(men_men_n59_), .C(b), .Y(men_men_n838_));
  AOI220     u0810(.A0(men_men_n637_), .A1(men_men_n29_), .B0(men_men_n485_), .B1(men_men_n85_), .Y(men_men_n839_));
  NA2        u0811(.A(men_men_n839_), .B(men_men_n838_), .Y(men_men_n840_));
  NO2        u0812(.A(men_men_n827_), .B(men_men_n514_), .Y(men_men_n841_));
  AOI210     u0813(.A0(men_men_n840_), .A1(men_men_n837_), .B0(men_men_n841_), .Y(men_men_n842_));
  NA3        u0814(.A(men_men_n842_), .B(men_men_n836_), .C(men_men_n834_), .Y(men_men_n843_));
  NOi41      u0815(.An(men_men_n799_), .B(men_men_n843_), .C(men_men_n832_), .D(men_men_n821_), .Y(men_men_n844_));
  OR3        u0816(.A(men_men_n745_), .B(men_men_n239_), .C(g), .Y(men_men_n845_));
  NO3        u0817(.A(men_men_n358_), .B(men_men_n313_), .C(men_men_n115_), .Y(men_men_n846_));
  NA2        u0818(.A(men_men_n846_), .B(men_men_n808_), .Y(men_men_n847_));
  NA2        u0819(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n848_));
  NO3        u0820(.A(men_men_n848_), .B(men_men_n797_), .C(men_men_n288_), .Y(men_men_n849_));
  NO3        u0821(.A(men_men_n553_), .B(men_men_n95_), .C(h), .Y(men_men_n850_));
  AOI210     u0822(.A0(men_men_n850_), .A1(men_men_n740_), .B0(men_men_n849_), .Y(men_men_n851_));
  NA4        u0823(.A(men_men_n851_), .B(men_men_n847_), .C(men_men_n845_), .D(men_men_n424_), .Y(men_men_n852_));
  NOi31      u0824(.An(b), .B(d), .C(a), .Y(men_men_n853_));
  NO2        u0825(.A(men_men_n853_), .B(men_men_n635_), .Y(men_men_n854_));
  NO2        u0826(.A(men_men_n854_), .B(n), .Y(men_men_n855_));
  NOi21      u0827(.An(men_men_n839_), .B(men_men_n855_), .Y(men_men_n856_));
  OAI220     u0828(.A0(men_men_n856_), .A1(men_men_n695_), .B0(men_men_n827_), .B1(men_men_n636_), .Y(men_men_n857_));
  NO2        u0829(.A(men_men_n582_), .B(men_men_n85_), .Y(men_men_n858_));
  NO3        u0830(.A(men_men_n656_), .B(men_men_n343_), .C(men_men_n120_), .Y(men_men_n859_));
  NOi21      u0831(.An(men_men_n859_), .B(men_men_n167_), .Y(men_men_n860_));
  AOI210     u0832(.A0(men_men_n846_), .A1(men_men_n858_), .B0(men_men_n860_), .Y(men_men_n861_));
  OAI210     u0833(.A0(men_men_n745_), .A1(men_men_n413_), .B0(men_men_n861_), .Y(men_men_n862_));
  NO2        u0834(.A(men_men_n1622_), .B(n), .Y(men_men_n863_));
  AOI220     u0835(.A0(men_men_n814_), .A1(men_men_n702_), .B0(men_men_n863_), .B1(men_men_n735_), .Y(men_men_n864_));
  NO2        u0836(.A(men_men_n338_), .B(men_men_n244_), .Y(men_men_n865_));
  OAI210     u0837(.A0(men_men_n97_), .A1(men_men_n94_), .B0(men_men_n865_), .Y(men_men_n866_));
  NA2        u0838(.A(men_men_n124_), .B(men_men_n85_), .Y(men_men_n867_));
  AOI210     u0839(.A0(men_men_n445_), .A1(men_men_n437_), .B0(men_men_n867_), .Y(men_men_n868_));
  NAi21      u0840(.An(men_men_n868_), .B(men_men_n866_), .Y(men_men_n869_));
  NA2        u0841(.A(men_men_n768_), .B(men_men_n34_), .Y(men_men_n870_));
  NAi21      u0842(.An(men_men_n774_), .B(men_men_n456_), .Y(men_men_n871_));
  NO2        u0843(.A(men_men_n282_), .B(i), .Y(men_men_n872_));
  NA2        u0844(.A(men_men_n752_), .B(men_men_n366_), .Y(men_men_n873_));
  OAI210     u0845(.A0(men_men_n627_), .A1(men_men_n626_), .B0(men_men_n381_), .Y(men_men_n874_));
  AN3        u0846(.A(men_men_n874_), .B(men_men_n873_), .C(men_men_n871_), .Y(men_men_n875_));
  NAi41      u0847(.An(men_men_n869_), .B(men_men_n875_), .C(men_men_n870_), .D(men_men_n864_), .Y(men_men_n876_));
  NO4        u0848(.A(men_men_n876_), .B(men_men_n862_), .C(men_men_n857_), .D(men_men_n852_), .Y(men_men_n877_));
  NA4        u0849(.A(men_men_n877_), .B(men_men_n844_), .C(men_men_n794_), .D(men_men_n779_), .Y(men09));
  INV        u0850(.A(men_men_n125_), .Y(men_men_n879_));
  NA2        u0851(.A(f), .B(e), .Y(men_men_n880_));
  NO2        u0852(.A(men_men_n232_), .B(men_men_n115_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n881_), .B(g), .Y(men_men_n882_));
  NA4        u0854(.A(men_men_n324_), .B(men_men_n494_), .C(men_men_n270_), .D(men_men_n122_), .Y(men_men_n883_));
  AOI210     u0855(.A0(men_men_n883_), .A1(g), .B0(men_men_n491_), .Y(men_men_n884_));
  AOI210     u0856(.A0(men_men_n884_), .A1(men_men_n882_), .B0(men_men_n880_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n465_), .B(e), .Y(men_men_n886_));
  NO2        u0858(.A(men_men_n886_), .B(men_men_n537_), .Y(men_men_n887_));
  AOI210     u0859(.A0(men_men_n885_), .A1(men_men_n879_), .B0(men_men_n887_), .Y(men_men_n888_));
  NO2        u0860(.A(men_men_n210_), .B(men_men_n220_), .Y(men_men_n889_));
  NA3        u0861(.A(m), .B(l), .C(i), .Y(men_men_n890_));
  OAI220     u0862(.A0(men_men_n621_), .A1(men_men_n890_), .B0(men_men_n371_), .B1(men_men_n554_), .Y(men_men_n891_));
  NA4        u0863(.A(men_men_n89_), .B(men_men_n88_), .C(g), .D(f), .Y(men_men_n892_));
  NAi31      u0864(.An(men_men_n891_), .B(men_men_n892_), .C(men_men_n460_), .Y(men_men_n893_));
  OA210      u0865(.A0(men_men_n893_), .A1(men_men_n889_), .B0(men_men_n595_), .Y(men_men_n894_));
  NA3        u0866(.A(men_men_n695_), .B(men_men_n597_), .C(men_men_n546_), .Y(men_men_n895_));
  OA210      u0867(.A0(men_men_n895_), .A1(men_men_n894_), .B0(men_men_n855_), .Y(men_men_n896_));
  INV        u0868(.A(men_men_n355_), .Y(men_men_n897_));
  NO2        u0869(.A(men_men_n131_), .B(men_men_n129_), .Y(men_men_n898_));
  NOi31      u0870(.An(k), .B(m), .C(l), .Y(men_men_n899_));
  NO2        u0871(.A(men_men_n357_), .B(men_men_n899_), .Y(men_men_n900_));
  AOI210     u0872(.A0(men_men_n900_), .A1(men_men_n898_), .B0(men_men_n630_), .Y(men_men_n901_));
  NA2        u0873(.A(men_men_n838_), .B(men_men_n348_), .Y(men_men_n902_));
  NA2        u0874(.A(men_men_n359_), .B(men_men_n361_), .Y(men_men_n903_));
  OAI210     u0875(.A0(men_men_n210_), .A1(men_men_n220_), .B0(men_men_n903_), .Y(men_men_n904_));
  AOI220     u0876(.A0(men_men_n904_), .A1(men_men_n902_), .B0(men_men_n901_), .B1(men_men_n897_), .Y(men_men_n905_));
  NA2        u0877(.A(men_men_n176_), .B(men_men_n117_), .Y(men_men_n906_));
  NA3        u0878(.A(men_men_n906_), .B(men_men_n734_), .C(men_men_n140_), .Y(men_men_n907_));
  NA3        u0879(.A(men_men_n907_), .B(men_men_n197_), .C(men_men_n31_), .Y(men_men_n908_));
  NA4        u0880(.A(men_men_n908_), .B(men_men_n905_), .C(men_men_n658_), .D(men_men_n83_), .Y(men_men_n909_));
  NO2        u0881(.A(men_men_n617_), .B(j), .Y(men_men_n910_));
  NA2        u0882(.A(men_men_n910_), .B(men_men_n197_), .Y(men_men_n911_));
  NOi21      u0883(.An(f), .B(d), .Y(men_men_n912_));
  NA2        u0884(.A(men_men_n912_), .B(m), .Y(men_men_n913_));
  NO2        u0885(.A(men_men_n913_), .B(men_men_n52_), .Y(men_men_n914_));
  NOi32      u0886(.An(g), .Bn(f), .C(d), .Y(men_men_n915_));
  NA4        u0887(.A(men_men_n915_), .B(men_men_n637_), .C(men_men_n29_), .D(m), .Y(men_men_n916_));
  NOi21      u0888(.An(men_men_n325_), .B(men_men_n916_), .Y(men_men_n917_));
  AOI210     u0889(.A0(men_men_n914_), .A1(men_men_n572_), .B0(men_men_n917_), .Y(men_men_n918_));
  NA3        u0890(.A(men_men_n324_), .B(men_men_n270_), .C(men_men_n122_), .Y(men_men_n919_));
  AN2        u0891(.A(f), .B(d), .Y(men_men_n920_));
  NA3        u0892(.A(men_men_n499_), .B(men_men_n920_), .C(men_men_n85_), .Y(men_men_n921_));
  NO3        u0893(.A(men_men_n921_), .B(men_men_n74_), .C(men_men_n221_), .Y(men_men_n922_));
  NO2        u0894(.A(men_men_n297_), .B(men_men_n56_), .Y(men_men_n923_));
  OAI210     u0895(.A0(men_men_n923_), .A1(men_men_n919_), .B0(men_men_n922_), .Y(men_men_n924_));
  NAi41      u0896(.An(men_men_n513_), .B(men_men_n924_), .C(men_men_n918_), .D(men_men_n911_), .Y(men_men_n925_));
  NO4        u0897(.A(men_men_n656_), .B(men_men_n136_), .C(men_men_n343_), .D(men_men_n158_), .Y(men_men_n926_));
  NO2        u0898(.A(men_men_n688_), .B(men_men_n343_), .Y(men_men_n927_));
  AN2        u0899(.A(men_men_n927_), .B(men_men_n717_), .Y(men_men_n928_));
  NO3        u0900(.A(men_men_n928_), .B(men_men_n926_), .C(men_men_n241_), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n635_), .B(men_men_n85_), .Y(men_men_n930_));
  OAI220     u0902(.A0(men_men_n903_), .A1(men_men_n930_), .B0(men_men_n838_), .B1(men_men_n460_), .Y(men_men_n931_));
  NA3        u0903(.A(men_men_n166_), .B(men_men_n111_), .C(men_men_n110_), .Y(men_men_n932_));
  OAI220     u0904(.A0(men_men_n921_), .A1(men_men_n450_), .B0(men_men_n355_), .B1(men_men_n932_), .Y(men_men_n933_));
  NOi41      u0905(.An(men_men_n230_), .B(men_men_n933_), .C(men_men_n931_), .D(men_men_n320_), .Y(men_men_n934_));
  NA2        u0906(.A(c), .B(men_men_n119_), .Y(men_men_n935_));
  NO2        u0907(.A(men_men_n935_), .B(men_men_n428_), .Y(men_men_n936_));
  NA3        u0908(.A(men_men_n936_), .B(men_men_n535_), .C(f), .Y(men_men_n937_));
  OR2        u0909(.A(men_men_n695_), .B(men_men_n569_), .Y(men_men_n938_));
  OAI210     u0910(.A0(men_men_n600_), .A1(men_men_n650_), .B0(men_men_n938_), .Y(men_men_n939_));
  NA2        u0911(.A(men_men_n854_), .B(men_men_n114_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n940_), .B(men_men_n939_), .Y(men_men_n941_));
  NA4        u0913(.A(men_men_n941_), .B(men_men_n937_), .C(men_men_n934_), .D(men_men_n929_), .Y(men_men_n942_));
  NO4        u0914(.A(men_men_n942_), .B(men_men_n925_), .C(men_men_n909_), .D(men_men_n896_), .Y(men_men_n943_));
  NA2        u0915(.A(men_men_n115_), .B(j), .Y(men_men_n944_));
  NO2        u0916(.A(men_men_n944_), .B(men_men_n149_), .Y(men_men_n945_));
  OAI210     u0917(.A0(men_men_n945_), .A1(men_men_n881_), .B0(g), .Y(men_men_n946_));
  AOI210     u0918(.A0(men_men_n946_), .A1(men_men_n305_), .B0(men_men_n921_), .Y(men_men_n947_));
  AOI210     u0919(.A0(men_men_n838_), .A1(men_men_n348_), .B0(men_men_n892_), .Y(men_men_n948_));
  NO2        u0920(.A(men_men_n140_), .B(men_men_n136_), .Y(men_men_n949_));
  NO2        u0921(.A(men_men_n237_), .B(men_men_n231_), .Y(men_men_n950_));
  AOI220     u0922(.A0(men_men_n950_), .A1(men_men_n234_), .B0(men_men_n318_), .B1(men_men_n949_), .Y(men_men_n951_));
  NO2        u0923(.A(men_men_n450_), .B(men_men_n880_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n952_), .B(men_men_n589_), .Y(men_men_n953_));
  NA2        u0925(.A(men_men_n953_), .B(men_men_n951_), .Y(men_men_n954_));
  NA2        u0926(.A(e), .B(d), .Y(men_men_n955_));
  NA3        u0927(.A(e), .B(men_men_n475_), .C(men_men_n533_), .Y(men_men_n956_));
  AOI210     u0928(.A0(men_men_n541_), .A1(men_men_n188_), .B0(men_men_n237_), .Y(men_men_n957_));
  AOI210     u0929(.A0(men_men_n657_), .A1(men_men_n364_), .B0(men_men_n957_), .Y(men_men_n958_));
  NA2        u0930(.A(men_men_n297_), .B(men_men_n172_), .Y(men_men_n959_));
  NA3        u0931(.A(men_men_n922_), .B(men_men_n959_), .C(men_men_n56_), .Y(men_men_n960_));
  NA3        u0932(.A(men_men_n175_), .B(men_men_n86_), .C(men_men_n34_), .Y(men_men_n961_));
  NA4        u0933(.A(men_men_n961_), .B(men_men_n960_), .C(men_men_n958_), .D(men_men_n956_), .Y(men_men_n962_));
  NO4        u0934(.A(men_men_n962_), .B(men_men_n954_), .C(men_men_n948_), .D(men_men_n947_), .Y(men_men_n963_));
  NA2        u0935(.A(men_men_n897_), .B(men_men_n31_), .Y(men_men_n964_));
  AO210      u0936(.A0(men_men_n964_), .A1(men_men_n736_), .B0(men_men_n224_), .Y(men_men_n965_));
  OAI220     u0937(.A0(men_men_n656_), .A1(men_men_n60_), .B0(men_men_n313_), .B1(j), .Y(men_men_n966_));
  AOI220     u0938(.A0(men_men_n966_), .A1(men_men_n927_), .B0(men_men_n647_), .B1(men_men_n655_), .Y(men_men_n967_));
  OAI210     u0939(.A0(men_men_n886_), .A1(men_men_n179_), .B0(men_men_n967_), .Y(men_men_n968_));
  OAI210     u0940(.A0(men_men_n881_), .A1(men_men_n959_), .B0(men_men_n915_), .Y(men_men_n969_));
  NO2        u0941(.A(men_men_n969_), .B(men_men_n638_), .Y(men_men_n970_));
  AOI210     u0942(.A0(men_men_n121_), .A1(men_men_n120_), .B0(men_men_n269_), .Y(men_men_n971_));
  NO2        u0943(.A(men_men_n971_), .B(men_men_n916_), .Y(men_men_n972_));
  AO210      u0944(.A0(men_men_n902_), .A1(men_men_n891_), .B0(men_men_n972_), .Y(men_men_n973_));
  NOi31      u0945(.An(men_men_n572_), .B(men_men_n913_), .C(men_men_n305_), .Y(men_men_n974_));
  NO4        u0946(.A(men_men_n974_), .B(men_men_n973_), .C(men_men_n970_), .D(men_men_n968_), .Y(men_men_n975_));
  AO220      u0947(.A0(men_men_n475_), .A1(men_men_n789_), .B0(men_men_n183_), .B1(f), .Y(men_men_n976_));
  OAI210     u0948(.A0(men_men_n976_), .A1(men_men_n478_), .B0(e), .Y(men_men_n977_));
  NO2        u0949(.A(men_men_n459_), .B(men_men_n70_), .Y(men_men_n978_));
  OAI210     u0950(.A0(men_men_n895_), .A1(men_men_n978_), .B0(men_men_n740_), .Y(men_men_n979_));
  AN4        u0951(.A(men_men_n979_), .B(men_men_n977_), .C(men_men_n975_), .D(men_men_n965_), .Y(men_men_n980_));
  NA4        u0952(.A(men_men_n980_), .B(men_men_n963_), .C(men_men_n943_), .D(men_men_n888_), .Y(men12));
  NO2        u0953(.A(men_men_n474_), .B(c), .Y(men_men_n982_));
  NO4        u0954(.A(men_men_n464_), .B(men_men_n261_), .C(men_men_n613_), .D(men_men_n221_), .Y(men_men_n983_));
  NA2        u0955(.A(men_men_n983_), .B(men_men_n982_), .Y(men_men_n984_));
  NA2        u0956(.A(men_men_n572_), .B(men_men_n978_), .Y(men_men_n985_));
  NO2        u0957(.A(men_men_n898_), .B(men_men_n371_), .Y(men_men_n986_));
  NO2        u0958(.A(men_men_n695_), .B(men_men_n398_), .Y(men_men_n987_));
  AOI220     u0959(.A0(men_men_n987_), .A1(men_men_n571_), .B0(men_men_n986_), .B1(men_men_n1629_), .Y(men_men_n988_));
  NA4        u0960(.A(men_men_n988_), .B(men_men_n985_), .C(men_men_n984_), .D(men_men_n463_), .Y(men_men_n989_));
  AOI210     u0961(.A0(men_men_n240_), .A1(men_men_n354_), .B0(men_men_n207_), .Y(men_men_n990_));
  OAI210     u0962(.A0(men_men_n408_), .A1(men_men_n1628_), .B0(men_men_n423_), .Y(men_men_n991_));
  NO2        u0963(.A(men_men_n676_), .B(men_men_n272_), .Y(men_men_n992_));
  NO2        u0964(.A(men_men_n621_), .B(men_men_n890_), .Y(men_men_n993_));
  AOI220     u0965(.A0(men_men_n993_), .A1(men_men_n595_), .B0(men_men_n865_), .B1(men_men_n992_), .Y(men_men_n994_));
  NO2        u0966(.A(men_men_n157_), .B(men_men_n244_), .Y(men_men_n995_));
  NA3        u0967(.A(men_men_n995_), .B(men_men_n247_), .C(i), .Y(men_men_n996_));
  NA3        u0968(.A(men_men_n996_), .B(men_men_n994_), .C(men_men_n991_), .Y(men_men_n997_));
  OR2        u0969(.A(men_men_n339_), .B(men_men_n1629_), .Y(men_men_n998_));
  NA2        u0970(.A(men_men_n998_), .B(men_men_n372_), .Y(men_men_n999_));
  NO3        u0971(.A(men_men_n136_), .B(men_men_n158_), .C(men_men_n221_), .Y(men_men_n1000_));
  NA2        u0972(.A(men_men_n1000_), .B(men_men_n558_), .Y(men_men_n1001_));
  NA4        u0973(.A(men_men_n465_), .B(men_men_n457_), .C(men_men_n189_), .D(g), .Y(men_men_n1002_));
  NA3        u0974(.A(men_men_n1002_), .B(men_men_n1001_), .C(men_men_n999_), .Y(men_men_n1003_));
  NO3        u0975(.A(men_men_n700_), .B(men_men_n93_), .C(men_men_n45_), .Y(men_men_n1004_));
  NO4        u0976(.A(men_men_n1004_), .B(men_men_n1003_), .C(men_men_n997_), .D(men_men_n989_), .Y(men_men_n1005_));
  NO2        u0977(.A(men_men_n388_), .B(men_men_n387_), .Y(men_men_n1006_));
  NA2        u0978(.A(men_men_n618_), .B(men_men_n72_), .Y(men_men_n1007_));
  NA2        u0979(.A(men_men_n582_), .B(men_men_n150_), .Y(men_men_n1008_));
  NOi21      u0980(.An(men_men_n34_), .B(men_men_n688_), .Y(men_men_n1009_));
  AOI220     u0981(.A0(men_men_n1009_), .A1(men_men_n1008_), .B0(men_men_n1007_), .B1(men_men_n1006_), .Y(men_men_n1010_));
  OAI210     u0982(.A0(men_men_n259_), .A1(men_men_n45_), .B0(men_men_n1010_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n456_), .B(men_men_n274_), .Y(men_men_n1012_));
  NO3        u0984(.A(men_men_n867_), .B(men_men_n90_), .C(men_men_n428_), .Y(men_men_n1013_));
  NAi31      u0985(.An(men_men_n1013_), .B(men_men_n1012_), .C(men_men_n335_), .Y(men_men_n1014_));
  NO2        u0986(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n1015_));
  NO2        u0987(.A(men_men_n529_), .B(men_men_n313_), .Y(men_men_n1016_));
  NO2        u0988(.A(men_men_n529_), .B(men_men_n150_), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n667_), .B(men_men_n381_), .Y(men_men_n1018_));
  OAI210     u0990(.A0(men_men_n775_), .A1(men_men_n1018_), .B0(men_men_n385_), .Y(men_men_n1019_));
  NO4        u0991(.A(men_men_n1019_), .B(men_men_n1017_), .C(men_men_n1014_), .D(men_men_n1011_), .Y(men_men_n1020_));
  NA2        u0992(.A(men_men_n364_), .B(g), .Y(men_men_n1021_));
  NA2        u0993(.A(men_men_n46_), .B(i), .Y(men_men_n1022_));
  OAI220     u0994(.A0(men_men_n1022_), .A1(men_men_n206_), .B0(g), .B1(men_men_n93_), .Y(men_men_n1023_));
  AOI210     u0995(.A0(men_men_n439_), .A1(men_men_n37_), .B0(men_men_n1023_), .Y(men_men_n1024_));
  NO2        u0996(.A(men_men_n150_), .B(men_men_n85_), .Y(men_men_n1025_));
  OR2        u0997(.A(men_men_n1025_), .B(men_men_n581_), .Y(men_men_n1026_));
  NA2        u0998(.A(men_men_n582_), .B(men_men_n402_), .Y(men_men_n1027_));
  AOI210     u0999(.A0(men_men_n1027_), .A1(n), .B0(men_men_n1026_), .Y(men_men_n1028_));
  OAI220     u1000(.A0(men_men_n1028_), .A1(men_men_n1021_), .B0(men_men_n1024_), .B1(men_men_n348_), .Y(men_men_n1029_));
  NO2        u1001(.A(men_men_n695_), .B(j), .Y(men_men_n1030_));
  NA3        u1002(.A(men_men_n359_), .B(men_men_n662_), .C(i), .Y(men_men_n1031_));
  OAI210     u1003(.A0(men_men_n459_), .A1(men_men_n324_), .B0(men_men_n1031_), .Y(men_men_n1032_));
  OAI220     u1004(.A0(men_men_n1032_), .A1(men_men_n1030_), .B0(men_men_n713_), .B1(men_men_n801_), .Y(men_men_n1033_));
  NA2        u1005(.A(men_men_n641_), .B(men_men_n116_), .Y(men_men_n1034_));
  OR3        u1006(.A(men_men_n324_), .B(men_men_n455_), .C(f), .Y(men_men_n1035_));
  NA3        u1007(.A(men_men_n662_), .B(men_men_n81_), .C(i), .Y(men_men_n1036_));
  OA220      u1008(.A0(men_men_n1036_), .A1(men_men_n1034_), .B0(men_men_n1035_), .B1(men_men_n620_), .Y(men_men_n1037_));
  NA3        u1009(.A(men_men_n340_), .B(men_men_n121_), .C(g), .Y(men_men_n1038_));
  AOI210     u1010(.A0(men_men_n710_), .A1(men_men_n1038_), .B0(m), .Y(men_men_n1039_));
  OAI210     u1011(.A0(men_men_n1039_), .A1(men_men_n986_), .B0(men_men_n339_), .Y(men_men_n1040_));
  NA2        u1012(.A(men_men_n727_), .B(men_men_n930_), .Y(men_men_n1041_));
  NA2        u1013(.A(men_men_n892_), .B(men_men_n460_), .Y(men_men_n1042_));
  NA2        u1014(.A(i), .B(men_men_n78_), .Y(men_men_n1043_));
  NA3        u1015(.A(men_men_n1043_), .B(men_men_n1036_), .C(men_men_n1035_), .Y(men_men_n1044_));
  AOI220     u1016(.A0(men_men_n1044_), .A1(men_men_n267_), .B0(men_men_n1042_), .B1(men_men_n1041_), .Y(men_men_n1045_));
  NA4        u1017(.A(men_men_n1045_), .B(men_men_n1040_), .C(men_men_n1037_), .D(men_men_n1033_), .Y(men_men_n1046_));
  NO2        u1018(.A(men_men_n398_), .B(men_men_n92_), .Y(men_men_n1047_));
  OAI210     u1019(.A0(men_men_n1047_), .A1(men_men_n992_), .B0(men_men_n245_), .Y(men_men_n1048_));
  NA2        u1020(.A(men_men_n699_), .B(men_men_n89_), .Y(men_men_n1049_));
  NO2        u1021(.A(men_men_n480_), .B(men_men_n221_), .Y(men_men_n1050_));
  AOI220     u1022(.A0(men_men_n1050_), .A1(men_men_n403_), .B0(men_men_n998_), .B1(men_men_n225_), .Y(men_men_n1051_));
  AOI220     u1023(.A0(men_men_n987_), .A1(men_men_n995_), .B0(men_men_n619_), .B1(men_men_n91_), .Y(men_men_n1052_));
  NA4        u1024(.A(men_men_n1052_), .B(men_men_n1051_), .C(men_men_n1049_), .D(men_men_n1048_), .Y(men_men_n1053_));
  OAI210     u1025(.A0(men_men_n1042_), .A1(men_men_n993_), .B0(men_men_n571_), .Y(men_men_n1054_));
  AOI210     u1026(.A0(men_men_n440_), .A1(men_men_n432_), .B0(men_men_n867_), .Y(men_men_n1055_));
  OAI210     u1027(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n112_), .Y(men_men_n1056_));
  AOI210     u1028(.A0(men_men_n1056_), .A1(men_men_n563_), .B0(men_men_n1055_), .Y(men_men_n1057_));
  NA2        u1029(.A(men_men_n1039_), .B(men_men_n1629_), .Y(men_men_n1058_));
  NO3        u1030(.A(men_men_n944_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1059_));
  AOI220     u1031(.A0(men_men_n1059_), .A1(men_men_n660_), .B0(men_men_n680_), .B1(men_men_n558_), .Y(men_men_n1060_));
  NA4        u1032(.A(men_men_n1060_), .B(men_men_n1058_), .C(men_men_n1057_), .D(men_men_n1054_), .Y(men_men_n1061_));
  NO4        u1033(.A(men_men_n1061_), .B(men_men_n1053_), .C(men_men_n1046_), .D(men_men_n1029_), .Y(men_men_n1062_));
  NAi31      u1034(.An(men_men_n146_), .B(men_men_n441_), .C(n), .Y(men_men_n1063_));
  NO3        u1035(.A(men_men_n129_), .B(men_men_n357_), .C(men_men_n899_), .Y(men_men_n1064_));
  NO2        u1036(.A(men_men_n1064_), .B(men_men_n1063_), .Y(men_men_n1065_));
  NO3        u1037(.A(men_men_n282_), .B(men_men_n146_), .C(men_men_n428_), .Y(men_men_n1066_));
  AOI210     u1038(.A0(men_men_n1066_), .A1(men_men_n523_), .B0(men_men_n1065_), .Y(men_men_n1067_));
  NA2        u1039(.A(men_men_n516_), .B(i), .Y(men_men_n1068_));
  NA2        u1040(.A(men_men_n1068_), .B(men_men_n1067_), .Y(men_men_n1069_));
  NA2        u1041(.A(men_men_n237_), .B(men_men_n180_), .Y(men_men_n1070_));
  NO3        u1042(.A(men_men_n322_), .B(men_men_n465_), .C(men_men_n183_), .Y(men_men_n1071_));
  NOi31      u1043(.An(men_men_n1070_), .B(men_men_n1071_), .C(men_men_n221_), .Y(men_men_n1072_));
  NAi21      u1044(.An(men_men_n582_), .B(men_men_n1050_), .Y(men_men_n1073_));
  NA2        u1045(.A(men_men_n458_), .B(men_men_n930_), .Y(men_men_n1074_));
  NO3        u1046(.A(men_men_n459_), .B(men_men_n324_), .C(men_men_n74_), .Y(men_men_n1075_));
  AOI220     u1047(.A0(men_men_n1075_), .A1(men_men_n1074_), .B0(men_men_n505_), .B1(g), .Y(men_men_n1076_));
  NA2        u1048(.A(men_men_n1076_), .B(men_men_n1073_), .Y(men_men_n1077_));
  OAI220     u1049(.A0(men_men_n1063_), .A1(men_men_n240_), .B0(men_men_n1031_), .B1(men_men_n636_), .Y(men_men_n1078_));
  NO2        u1050(.A(men_men_n696_), .B(men_men_n398_), .Y(men_men_n1079_));
  NA2        u1051(.A(men_men_n990_), .B(men_men_n982_), .Y(men_men_n1080_));
  NO3        u1052(.A(c), .B(men_men_n155_), .C(men_men_n220_), .Y(men_men_n1081_));
  OAI210     u1053(.A0(men_men_n1081_), .A1(men_men_n552_), .B0(men_men_n399_), .Y(men_men_n1082_));
  OAI220     u1054(.A0(men_men_n987_), .A1(men_men_n993_), .B0(men_men_n572_), .B1(men_men_n449_), .Y(men_men_n1083_));
  NA4        u1055(.A(men_men_n1083_), .B(men_men_n1082_), .C(men_men_n1080_), .D(men_men_n654_), .Y(men_men_n1084_));
  OAI210     u1056(.A0(men_men_n990_), .A1(men_men_n983_), .B0(men_men_n1070_), .Y(men_men_n1085_));
  NA3        u1057(.A(men_men_n1027_), .B(men_men_n510_), .C(men_men_n46_), .Y(men_men_n1086_));
  AOI210     u1058(.A0(men_men_n401_), .A1(men_men_n399_), .B0(men_men_n347_), .Y(men_men_n1087_));
  NA4        u1059(.A(men_men_n1087_), .B(men_men_n1086_), .C(men_men_n1085_), .D(men_men_n283_), .Y(men_men_n1088_));
  OR4        u1060(.A(men_men_n1088_), .B(men_men_n1084_), .C(men_men_n1079_), .D(men_men_n1078_), .Y(men_men_n1089_));
  NO4        u1061(.A(men_men_n1089_), .B(men_men_n1077_), .C(men_men_n1072_), .D(men_men_n1069_), .Y(men_men_n1090_));
  NA4        u1062(.A(men_men_n1090_), .B(men_men_n1062_), .C(men_men_n1020_), .D(men_men_n1005_), .Y(men13));
  NA2        u1063(.A(men_men_n46_), .B(men_men_n88_), .Y(men_men_n1092_));
  AN2        u1064(.A(c), .B(b), .Y(men_men_n1093_));
  NA3        u1065(.A(men_men_n258_), .B(men_men_n1093_), .C(m), .Y(men_men_n1094_));
  NO4        u1066(.A(e), .B(men_men_n1094_), .C(men_men_n1092_), .D(men_men_n614_), .Y(men_men_n1095_));
  NA2        u1067(.A(men_men_n274_), .B(men_men_n1093_), .Y(men_men_n1096_));
  NO4        u1068(.A(men_men_n1096_), .B(e), .C(g), .D(a), .Y(men_men_n1097_));
  NAi32      u1069(.An(d), .Bn(c), .C(e), .Y(men_men_n1098_));
  NO3        u1070(.A(men_men_n1098_), .B(men_men_n621_), .C(men_men_n321_), .Y(men_men_n1099_));
  NA2        u1071(.A(men_men_n703_), .B(men_men_n231_), .Y(men_men_n1100_));
  NA2        u1072(.A(men_men_n431_), .B(men_men_n220_), .Y(men_men_n1101_));
  AN2        u1073(.A(d), .B(c), .Y(men_men_n1102_));
  NA2        u1074(.A(men_men_n1102_), .B(men_men_n119_), .Y(men_men_n1103_));
  NO4        u1075(.A(men_men_n1103_), .B(men_men_n1101_), .C(men_men_n184_), .D(men_men_n176_), .Y(men_men_n1104_));
  NA2        u1076(.A(men_men_n521_), .B(c), .Y(men_men_n1105_));
  NO3        u1077(.A(men_men_n617_), .B(men_men_n1105_), .C(men_men_n321_), .Y(men_men_n1106_));
  AO210      u1078(.A0(men_men_n1104_), .A1(men_men_n1100_), .B0(men_men_n1106_), .Y(men_men_n1107_));
  OR4        u1079(.A(men_men_n1107_), .B(men_men_n1099_), .C(men_men_n1097_), .D(men_men_n1095_), .Y(men_men_n1108_));
  NAi32      u1080(.An(f), .Bn(e), .C(c), .Y(men_men_n1109_));
  NO2        u1081(.A(men_men_n1109_), .B(men_men_n152_), .Y(men_men_n1110_));
  NA2        u1082(.A(men_men_n1110_), .B(g), .Y(men_men_n1111_));
  NO2        u1083(.A(men_men_n184_), .B(men_men_n1111_), .Y(men_men_n1112_));
  NO2        u1084(.A(j), .B(men_men_n45_), .Y(men_men_n1113_));
  NA2        u1085(.A(men_men_n664_), .B(men_men_n1113_), .Y(men_men_n1114_));
  NOi21      u1086(.An(men_men_n1625_), .B(men_men_n1114_), .Y(men_men_n1115_));
  NO2        u1087(.A(men_men_n805_), .B(men_men_n115_), .Y(men_men_n1116_));
  NO2        u1088(.A(men_men_n1623_), .B(men_men_n1111_), .Y(men_men_n1117_));
  OR3        u1089(.A(e), .B(d), .C(c), .Y(men_men_n1118_));
  NA3        u1090(.A(k), .B(j), .C(i), .Y(men_men_n1119_));
  NO3        u1091(.A(men_men_n1119_), .B(men_men_n321_), .C(men_men_n92_), .Y(men_men_n1120_));
  NOi21      u1092(.An(men_men_n1120_), .B(men_men_n1118_), .Y(men_men_n1121_));
  OR4        u1093(.A(men_men_n1121_), .B(men_men_n1117_), .C(men_men_n1115_), .D(men_men_n1112_), .Y(men_men_n1122_));
  NA3        u1094(.A(men_men_n488_), .B(men_men_n350_), .C(men_men_n56_), .Y(men_men_n1123_));
  NO2        u1095(.A(men_men_n1123_), .B(men_men_n1114_), .Y(men_men_n1124_));
  NO4        u1096(.A(men_men_n1123_), .B(men_men_n617_), .C(men_men_n471_), .D(men_men_n45_), .Y(men_men_n1125_));
  NO2        u1097(.A(f), .B(c), .Y(men_men_n1126_));
  NOi21      u1098(.An(men_men_n1126_), .B(men_men_n464_), .Y(men_men_n1127_));
  NA2        u1099(.A(men_men_n1127_), .B(men_men_n59_), .Y(men_men_n1128_));
  OR2        u1100(.A(k), .B(i), .Y(men_men_n1129_));
  NO3        u1101(.A(men_men_n1129_), .B(men_men_n251_), .C(l), .Y(men_men_n1130_));
  NOi31      u1102(.An(men_men_n1130_), .B(men_men_n1128_), .C(j), .Y(men_men_n1131_));
  OR3        u1103(.A(men_men_n1131_), .B(men_men_n1125_), .C(men_men_n1124_), .Y(men_men_n1132_));
  OR3        u1104(.A(men_men_n1132_), .B(men_men_n1122_), .C(men_men_n1108_), .Y(men02));
  OR2        u1105(.A(l), .B(k), .Y(men_men_n1134_));
  OR3        u1106(.A(h), .B(g), .C(f), .Y(men_men_n1135_));
  OR3        u1107(.A(n), .B(m), .C(i), .Y(men_men_n1136_));
  NO4        u1108(.A(men_men_n1136_), .B(men_men_n1135_), .C(men_men_n1134_), .D(men_men_n1118_), .Y(men_men_n1137_));
  NOi31      u1109(.An(e), .B(d), .C(c), .Y(men_men_n1138_));
  AOI210     u1110(.A0(men_men_n1120_), .A1(men_men_n1138_), .B0(men_men_n1099_), .Y(men_men_n1139_));
  AN3        u1111(.A(g), .B(f), .C(c), .Y(men_men_n1140_));
  NA3        u1112(.A(men_men_n1140_), .B(men_men_n488_), .C(h), .Y(men_men_n1141_));
  OR2        u1113(.A(men_men_n1119_), .B(men_men_n321_), .Y(men_men_n1142_));
  OR2        u1114(.A(men_men_n1142_), .B(men_men_n1141_), .Y(men_men_n1143_));
  NO2        u1115(.A(men_men_n1123_), .B(men_men_n617_), .Y(men_men_n1144_));
  NO2        u1116(.A(men_men_n1144_), .B(men_men_n1112_), .Y(men_men_n1145_));
  NA3        u1117(.A(l), .B(k), .C(j), .Y(men_men_n1146_));
  NA2        u1118(.A(i), .B(h), .Y(men_men_n1147_));
  NO3        u1119(.A(men_men_n1147_), .B(men_men_n1146_), .C(men_men_n136_), .Y(men_men_n1148_));
  NO3        u1120(.A(men_men_n147_), .B(men_men_n295_), .C(men_men_n221_), .Y(men_men_n1149_));
  AOI210     u1121(.A0(men_men_n1149_), .A1(men_men_n1148_), .B0(men_men_n1115_), .Y(men_men_n1150_));
  NA3        u1122(.A(c), .B(b), .C(a), .Y(men_men_n1151_));
  NO3        u1123(.A(men_men_n1151_), .B(men_men_n955_), .C(men_men_n220_), .Y(men_men_n1152_));
  NO4        u1124(.A(men_men_n1119_), .B(men_men_n313_), .C(men_men_n49_), .D(men_men_n115_), .Y(men_men_n1153_));
  AOI210     u1125(.A0(men_men_n1153_), .A1(men_men_n1152_), .B0(men_men_n1124_), .Y(men_men_n1154_));
  AN4        u1126(.A(men_men_n1154_), .B(men_men_n1150_), .C(men_men_n1145_), .D(men_men_n1143_), .Y(men_men_n1155_));
  NO2        u1127(.A(men_men_n1103_), .B(men_men_n1101_), .Y(men_men_n1156_));
  AOI210     u1128(.A0(men_men_n1624_), .A1(men_men_n1156_), .B0(men_men_n1095_), .Y(men_men_n1157_));
  NAi41      u1129(.An(men_men_n1137_), .B(men_men_n1157_), .C(men_men_n1155_), .D(men_men_n1139_), .Y(men03));
  NO2        u1130(.A(men_men_n554_), .B(men_men_n630_), .Y(men_men_n1159_));
  NA4        u1131(.A(men_men_n89_), .B(men_men_n88_), .C(g), .D(men_men_n220_), .Y(men_men_n1160_));
  NA4        u1132(.A(men_men_n605_), .B(m), .C(men_men_n115_), .D(men_men_n220_), .Y(men_men_n1161_));
  NA3        u1133(.A(men_men_n1161_), .B(men_men_n389_), .C(men_men_n1160_), .Y(men_men_n1162_));
  NO3        u1134(.A(men_men_n1162_), .B(men_men_n1159_), .C(men_men_n1056_), .Y(men_men_n1163_));
  NOi41      u1135(.An(men_men_n695_), .B(men_men_n904_), .C(men_men_n893_), .D(men_men_n754_), .Y(men_men_n1164_));
  OAI220     u1136(.A0(men_men_n1164_), .A1(men_men_n727_), .B0(men_men_n1163_), .B1(men_men_n618_), .Y(men_men_n1165_));
  NOi31      u1137(.An(i), .B(k), .C(j), .Y(men_men_n1166_));
  NA4        u1138(.A(men_men_n1166_), .B(men_men_n1138_), .C(men_men_n359_), .D(men_men_n350_), .Y(men_men_n1167_));
  OAI210     u1139(.A0(men_men_n867_), .A1(men_men_n442_), .B0(men_men_n1167_), .Y(men_men_n1168_));
  NOi31      u1140(.An(m), .B(n), .C(f), .Y(men_men_n1169_));
  NA2        u1141(.A(men_men_n1169_), .B(men_men_n51_), .Y(men_men_n1170_));
  AN2        u1142(.A(e), .B(c), .Y(men_men_n1171_));
  NA2        u1143(.A(men_men_n1171_), .B(a), .Y(men_men_n1172_));
  OAI220     u1144(.A0(men_men_n1172_), .A1(men_men_n1170_), .B0(men_men_n938_), .B1(men_men_n448_), .Y(men_men_n1173_));
  NA2        u1145(.A(men_men_n533_), .B(l), .Y(men_men_n1174_));
  NOi31      u1146(.An(men_men_n915_), .B(men_men_n1094_), .C(men_men_n1174_), .Y(men_men_n1175_));
  NO4        u1147(.A(men_men_n1175_), .B(men_men_n1173_), .C(men_men_n1168_), .D(men_men_n1055_), .Y(men_men_n1176_));
  NO2        u1148(.A(men_men_n295_), .B(a), .Y(men_men_n1177_));
  INV        u1149(.A(men_men_n1099_), .Y(men_men_n1178_));
  NO2        u1150(.A(men_men_n1147_), .B(men_men_n508_), .Y(men_men_n1179_));
  NO2        u1151(.A(men_men_n88_), .B(g), .Y(men_men_n1180_));
  AOI210     u1152(.A0(men_men_n1180_), .A1(men_men_n1179_), .B0(men_men_n1130_), .Y(men_men_n1181_));
  OR2        u1153(.A(men_men_n1181_), .B(men_men_n1128_), .Y(men_men_n1182_));
  NA3        u1154(.A(men_men_n1182_), .B(men_men_n1178_), .C(men_men_n1176_), .Y(men_men_n1183_));
  NO4        u1155(.A(men_men_n1183_), .B(men_men_n1165_), .C(men_men_n869_), .D(men_men_n594_), .Y(men_men_n1184_));
  NA2        u1156(.A(c), .B(b), .Y(men_men_n1185_));
  NO2        u1157(.A(men_men_n739_), .B(men_men_n1185_), .Y(men_men_n1186_));
  OAI210     u1158(.A0(men_men_n913_), .A1(men_men_n884_), .B0(men_men_n435_), .Y(men_men_n1187_));
  OAI210     u1159(.A0(men_men_n1187_), .A1(men_men_n914_), .B0(men_men_n1186_), .Y(men_men_n1188_));
  NAi21      u1160(.An(men_men_n443_), .B(men_men_n1186_), .Y(men_men_n1189_));
  NA3        u1161(.A(men_men_n449_), .B(men_men_n587_), .C(f), .Y(men_men_n1190_));
  OAI210     u1162(.A0(men_men_n576_), .A1(men_men_n39_), .B0(men_men_n1177_), .Y(men_men_n1191_));
  NA3        u1163(.A(men_men_n1191_), .B(men_men_n1190_), .C(men_men_n1189_), .Y(men_men_n1192_));
  NA2        u1164(.A(men_men_n270_), .B(men_men_n122_), .Y(men_men_n1193_));
  OAI210     u1165(.A0(men_men_n1193_), .A1(men_men_n299_), .B0(g), .Y(men_men_n1194_));
  NAi21      u1166(.An(f), .B(d), .Y(men_men_n1195_));
  NO2        u1167(.A(men_men_n1195_), .B(men_men_n1151_), .Y(men_men_n1196_));
  INV        u1168(.A(men_men_n1196_), .Y(men_men_n1197_));
  AOI210     u1169(.A0(men_men_n1194_), .A1(men_men_n305_), .B0(men_men_n1197_), .Y(men_men_n1198_));
  AOI210     u1170(.A0(men_men_n1198_), .A1(men_men_n116_), .B0(men_men_n1192_), .Y(men_men_n1199_));
  NA2        u1171(.A(men_men_n491_), .B(men_men_n490_), .Y(men_men_n1200_));
  NO2        u1172(.A(men_men_n190_), .B(men_men_n244_), .Y(men_men_n1201_));
  NA2        u1173(.A(men_men_n1201_), .B(m), .Y(men_men_n1202_));
  NA3        u1174(.A(men_men_n971_), .B(men_men_n1174_), .C(men_men_n494_), .Y(men_men_n1203_));
  OAI210     u1175(.A0(men_men_n1203_), .A1(men_men_n325_), .B0(men_men_n492_), .Y(men_men_n1204_));
  AOI210     u1176(.A0(men_men_n1204_), .A1(men_men_n1200_), .B0(men_men_n1202_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n589_), .B(men_men_n430_), .Y(men_men_n1206_));
  NA2        u1178(.A(men_men_n165_), .B(men_men_n33_), .Y(men_men_n1207_));
  AOI210     u1179(.A0(men_men_n1018_), .A1(men_men_n1207_), .B0(men_men_n221_), .Y(men_men_n1208_));
  OAI210     u1180(.A0(men_men_n1208_), .A1(men_men_n467_), .B0(men_men_n1196_), .Y(men_men_n1209_));
  NO2        u1181(.A(men_men_n392_), .B(men_men_n391_), .Y(men_men_n1210_));
  AOI210     u1182(.A0(men_men_n1201_), .A1(men_men_n451_), .B0(men_men_n1013_), .Y(men_men_n1211_));
  NAi41      u1183(.An(men_men_n1210_), .B(men_men_n1211_), .C(men_men_n1209_), .D(men_men_n1206_), .Y(men_men_n1212_));
  NO2        u1184(.A(men_men_n1212_), .B(men_men_n1205_), .Y(men_men_n1213_));
  NA4        u1185(.A(men_men_n1213_), .B(men_men_n1199_), .C(men_men_n1188_), .D(men_men_n1184_), .Y(men00));
  AOI210     u1186(.A0(men_men_n312_), .A1(men_men_n221_), .B0(men_men_n287_), .Y(men_men_n1215_));
  NO2        u1187(.A(men_men_n1215_), .B(men_men_n608_), .Y(men_men_n1216_));
  AOI210     u1188(.A0(men_men_n952_), .A1(men_men_n995_), .B0(men_men_n1168_), .Y(men_men_n1217_));
  NO3        u1189(.A(men_men_n1144_), .B(men_men_n1013_), .C(men_men_n751_), .Y(men_men_n1218_));
  NA3        u1190(.A(men_men_n1218_), .B(men_men_n1217_), .C(men_men_n1057_), .Y(men_men_n1219_));
  NA2        u1191(.A(men_men_n535_), .B(f), .Y(men_men_n1220_));
  OAI210     u1192(.A0(men_men_n1064_), .A1(men_men_n40_), .B0(men_men_n682_), .Y(men_men_n1221_));
  NA3        u1193(.A(men_men_n1221_), .B(men_men_n266_), .C(n), .Y(men_men_n1222_));
  AOI210     u1194(.A0(men_men_n1222_), .A1(men_men_n1220_), .B0(men_men_n1103_), .Y(men_men_n1223_));
  NO4        u1195(.A(men_men_n1223_), .B(men_men_n1219_), .C(men_men_n1216_), .D(men_men_n1122_), .Y(men_men_n1224_));
  NA3        u1196(.A(men_men_n175_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1225_));
  NA3        u1197(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1226_));
  NOi31      u1198(.An(n), .B(m), .C(i), .Y(men_men_n1227_));
  NA3        u1199(.A(men_men_n1227_), .B(d), .C(men_men_n51_), .Y(men_men_n1228_));
  OAI210     u1200(.A0(men_men_n1226_), .A1(men_men_n1225_), .B0(men_men_n1228_), .Y(men_men_n1229_));
  INV        u1201(.A(men_men_n607_), .Y(men_men_n1230_));
  NO4        u1202(.A(men_men_n1230_), .B(men_men_n1229_), .C(men_men_n1210_), .D(men_men_n974_), .Y(men_men_n1231_));
  NO4        u1203(.A(men_men_n511_), .B(men_men_n374_), .C(men_men_n1185_), .D(men_men_n59_), .Y(men_men_n1232_));
  NA3        u1204(.A(men_men_n404_), .B(men_men_n228_), .C(g), .Y(men_men_n1233_));
  OA220      u1205(.A0(men_men_n1233_), .A1(men_men_n1226_), .B0(men_men_n405_), .B1(men_men_n139_), .Y(men_men_n1234_));
  NO2        u1206(.A(h), .B(g), .Y(men_men_n1235_));
  NA4        u1207(.A(men_men_n523_), .B(men_men_n488_), .C(men_men_n1235_), .D(men_men_n1093_), .Y(men_men_n1236_));
  OAI220     u1208(.A0(men_men_n554_), .A1(men_men_n630_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n1237_));
  AOI220     u1209(.A0(men_men_n1237_), .A1(men_men_n563_), .B0(men_men_n1000_), .B1(men_men_n606_), .Y(men_men_n1238_));
  AOI220     u1210(.A0(men_men_n332_), .A1(men_men_n255_), .B0(men_men_n185_), .B1(men_men_n154_), .Y(men_men_n1239_));
  NA4        u1211(.A(men_men_n1239_), .B(men_men_n1238_), .C(men_men_n1236_), .D(men_men_n1234_), .Y(men_men_n1240_));
  NO3        u1212(.A(men_men_n1240_), .B(men_men_n1232_), .C(men_men_n276_), .Y(men_men_n1241_));
  INV        u1213(.A(men_men_n337_), .Y(men_men_n1242_));
  AOI210     u1214(.A0(men_men_n255_), .A1(men_men_n364_), .B0(men_men_n609_), .Y(men_men_n1243_));
  NA3        u1215(.A(men_men_n1243_), .B(men_men_n1242_), .C(men_men_n160_), .Y(men_men_n1244_));
  NO2        u1216(.A(men_men_n246_), .B(men_men_n189_), .Y(men_men_n1245_));
  NA2        u1217(.A(men_men_n1245_), .B(men_men_n449_), .Y(men_men_n1246_));
  NA3        u1218(.A(men_men_n187_), .B(men_men_n115_), .C(g), .Y(men_men_n1247_));
  NA3        u1219(.A(men_men_n488_), .B(men_men_n40_), .C(f), .Y(men_men_n1248_));
  NOi31      u1220(.An(men_men_n923_), .B(men_men_n1248_), .C(men_men_n1247_), .Y(men_men_n1249_));
  NAi31      u1221(.An(men_men_n193_), .B(men_men_n910_), .C(men_men_n488_), .Y(men_men_n1250_));
  NAi31      u1222(.An(men_men_n1249_), .B(men_men_n1250_), .C(men_men_n1246_), .Y(men_men_n1251_));
  NO3        u1223(.A(men_men_n448_), .B(men_men_n880_), .C(n), .Y(men_men_n1252_));
  AOI210     u1224(.A0(men_men_n1252_), .A1(men_men_n1630_), .B0(men_men_n1137_), .Y(men_men_n1253_));
  NAi31      u1225(.An(men_men_n1106_), .B(men_men_n1253_), .C(men_men_n73_), .Y(men_men_n1254_));
  NO4        u1226(.A(men_men_n1254_), .B(men_men_n1251_), .C(men_men_n1244_), .D(men_men_n545_), .Y(men_men_n1255_));
  AN3        u1227(.A(men_men_n1255_), .B(men_men_n1241_), .C(men_men_n1231_), .Y(men_men_n1256_));
  NA2        u1228(.A(men_men_n563_), .B(men_men_n103_), .Y(men_men_n1257_));
  NA3        u1229(.A(men_men_n1169_), .B(men_men_n641_), .C(men_men_n487_), .Y(men_men_n1258_));
  NA4        u1230(.A(men_men_n1258_), .B(men_men_n590_), .C(men_men_n1257_), .D(men_men_n249_), .Y(men_men_n1259_));
  NA2        u1231(.A(men_men_n1162_), .B(men_men_n563_), .Y(men_men_n1260_));
  NA4        u1232(.A(d), .B(men_men_n212_), .C(men_men_n228_), .D(men_men_n169_), .Y(men_men_n1261_));
  NA3        u1233(.A(men_men_n1261_), .B(men_men_n1260_), .C(men_men_n309_), .Y(men_men_n1262_));
  OAI210     u1234(.A0(men_men_n486_), .A1(men_men_n123_), .B0(men_men_n916_), .Y(men_men_n1263_));
  AOI220     u1235(.A0(men_men_n1263_), .A1(men_men_n1203_), .B0(men_men_n589_), .B1(men_men_n430_), .Y(men_men_n1264_));
  OR4        u1236(.A(men_men_n1103_), .B(men_men_n282_), .C(men_men_n229_), .D(e), .Y(men_men_n1265_));
  AOI220     u1237(.A0(d), .A1(men_men_n284_), .B0(men_men_n897_), .B1(men_men_n222_), .Y(men_men_n1266_));
  OAI210     u1238(.A0(men_men_n375_), .A1(men_men_n326_), .B0(men_men_n469_), .Y(men_men_n1267_));
  NA4        u1239(.A(men_men_n1267_), .B(men_men_n1266_), .C(men_men_n1265_), .D(men_men_n1264_), .Y(men_men_n1268_));
  AOI210     u1240(.A0(d), .A1(men_men_n901_), .B0(men_men_n868_), .Y(men_men_n1269_));
  AOI220     u1241(.A0(men_men_n1009_), .A1(men_men_n606_), .B0(d), .B1(men_men_n252_), .Y(men_men_n1270_));
  NO2        u1242(.A(men_men_n67_), .B(h), .Y(men_men_n1271_));
  NO3        u1243(.A(men_men_n1103_), .B(men_men_n1101_), .C(men_men_n767_), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n1134_), .B(men_men_n136_), .Y(men_men_n1273_));
  AN2        u1245(.A(men_men_n1273_), .B(men_men_n1149_), .Y(men_men_n1274_));
  OAI210     u1246(.A0(men_men_n1274_), .A1(men_men_n1272_), .B0(men_men_n1271_), .Y(men_men_n1275_));
  NA4        u1247(.A(men_men_n1275_), .B(men_men_n1270_), .C(men_men_n1269_), .D(men_men_n918_), .Y(men_men_n1276_));
  NO4        u1248(.A(men_men_n1276_), .B(men_men_n1268_), .C(men_men_n1262_), .D(men_men_n1259_), .Y(men_men_n1277_));
  NA2        u1249(.A(men_men_n885_), .B(men_men_n800_), .Y(men_men_n1278_));
  NA4        u1250(.A(men_men_n1278_), .B(men_men_n1277_), .C(men_men_n1256_), .D(men_men_n1224_), .Y(men01));
  AN2        u1251(.A(men_men_n1082_), .B(men_men_n1080_), .Y(men_men_n1280_));
  NO4        u1252(.A(men_men_n849_), .B(men_men_n841_), .C(men_men_n502_), .D(men_men_n293_), .Y(men_men_n1281_));
  NO2        u1253(.A(men_men_n623_), .B(men_men_n302_), .Y(men_men_n1282_));
  OAI210     u1254(.A0(men_men_n1282_), .A1(men_men_n414_), .B0(i), .Y(men_men_n1283_));
  NA3        u1255(.A(men_men_n1283_), .B(men_men_n1281_), .C(men_men_n1280_), .Y(men_men_n1284_));
  NA2        u1256(.A(men_men_n619_), .B(men_men_n91_), .Y(men_men_n1285_));
  NA2        u1257(.A(men_men_n582_), .B(men_men_n281_), .Y(men_men_n1286_));
  NA2        u1258(.A(men_men_n1016_), .B(men_men_n1286_), .Y(men_men_n1287_));
  NA4        u1259(.A(men_men_n1287_), .B(men_men_n1285_), .C(men_men_n967_), .D(men_men_n349_), .Y(men_men_n1288_));
  NA2        u1260(.A(men_men_n45_), .B(f), .Y(men_men_n1289_));
  NA2        u1261(.A(men_men_n746_), .B(men_men_n98_), .Y(men_men_n1290_));
  OAI220     u1262(.A0(men_men_n1290_), .A1(men_men_n1289_), .B0(men_men_n371_), .B1(men_men_n297_), .Y(men_men_n1291_));
  OAI210     u1263(.A0(men_men_n827_), .A1(men_men_n636_), .B0(men_men_n1261_), .Y(men_men_n1292_));
  AOI210     u1264(.A0(men_men_n1291_), .A1(men_men_n671_), .B0(men_men_n1292_), .Y(men_men_n1293_));
  NA2        u1265(.A(men_men_n121_), .B(l), .Y(men_men_n1294_));
  OA220      u1266(.A0(men_men_n1294_), .A1(men_men_n616_), .B0(men_men_n697_), .B1(men_men_n389_), .Y(men_men_n1295_));
  NAi41      u1267(.An(men_men_n168_), .B(men_men_n1295_), .C(men_men_n1293_), .D(men_men_n951_), .Y(men_men_n1296_));
  NO3        u1268(.A(men_men_n828_), .B(men_men_n712_), .C(men_men_n538_), .Y(men_men_n1297_));
  NA4        u1269(.A(men_men_n746_), .B(men_men_n98_), .C(men_men_n45_), .D(men_men_n220_), .Y(men_men_n1298_));
  OA220      u1270(.A0(men_men_n1298_), .A1(men_men_n705_), .B0(men_men_n201_), .B1(men_men_n1626_), .Y(men_men_n1299_));
  NA3        u1271(.A(men_men_n1299_), .B(men_men_n1297_), .C(men_men_n142_), .Y(men_men_n1300_));
  NO4        u1272(.A(men_men_n1300_), .B(men_men_n1296_), .C(men_men_n1288_), .D(men_men_n1284_), .Y(men_men_n1301_));
  NA2        u1273(.A(men_men_n1233_), .B(men_men_n213_), .Y(men_men_n1302_));
  OAI210     u1274(.A0(men_men_n1302_), .A1(men_men_n315_), .B0(men_men_n558_), .Y(men_men_n1303_));
  NA2        u1275(.A(men_men_n566_), .B(men_men_n416_), .Y(men_men_n1304_));
  NA2        u1276(.A(men_men_n75_), .B(i), .Y(men_men_n1305_));
  AOI210     u1277(.A0(men_men_n622_), .A1(men_men_n616_), .B0(men_men_n1305_), .Y(men_men_n1306_));
  NOi21      u1278(.An(men_men_n591_), .B(men_men_n613_), .Y(men_men_n1307_));
  AOI210     u1279(.A0(men_men_n1307_), .A1(men_men_n1304_), .B0(men_men_n1306_), .Y(men_men_n1308_));
  AOI210     u1280(.A0(men_men_n210_), .A1(men_men_n90_), .B0(men_men_n220_), .Y(men_men_n1309_));
  OAI210     u1281(.A0(men_men_n855_), .A1(men_men_n449_), .B0(men_men_n1309_), .Y(men_men_n1310_));
  AN3        u1282(.A(m), .B(l), .C(k), .Y(men_men_n1311_));
  OAI210     u1283(.A0(men_men_n377_), .A1(men_men_n34_), .B0(men_men_n1311_), .Y(men_men_n1312_));
  NA2        u1284(.A(men_men_n209_), .B(men_men_n34_), .Y(men_men_n1313_));
  AO210      u1285(.A0(men_men_n1313_), .A1(men_men_n1312_), .B0(men_men_n348_), .Y(men_men_n1314_));
  NA4        u1286(.A(men_men_n1314_), .B(men_men_n1310_), .C(men_men_n1308_), .D(men_men_n1303_), .Y(men_men_n1315_));
  AOI210     u1287(.A0(men_men_n628_), .A1(men_men_n121_), .B0(men_men_n634_), .Y(men_men_n1316_));
  OAI210     u1288(.A0(men_men_n1294_), .A1(men_men_n625_), .B0(men_men_n1316_), .Y(men_men_n1317_));
  NA2        u1289(.A(men_men_n292_), .B(men_men_n201_), .Y(men_men_n1318_));
  OAI210     u1290(.A0(men_men_n1318_), .A1(men_men_n406_), .B0(men_men_n702_), .Y(men_men_n1319_));
  NO3        u1291(.A(men_men_n867_), .B(men_men_n210_), .C(men_men_n428_), .Y(men_men_n1320_));
  NO2        u1292(.A(men_men_n1320_), .B(men_men_n1013_), .Y(men_men_n1321_));
  OAI210     u1293(.A0(men_men_n1291_), .A1(men_men_n342_), .B0(men_men_n713_), .Y(men_men_n1322_));
  NA4        u1294(.A(men_men_n1322_), .B(men_men_n1321_), .C(men_men_n1319_), .D(men_men_n831_), .Y(men_men_n1323_));
  NO3        u1295(.A(men_men_n1323_), .B(men_men_n1317_), .C(men_men_n1315_), .Y(men_men_n1324_));
  NA3        u1296(.A(men_men_n637_), .B(men_men_n29_), .C(f), .Y(men_men_n1325_));
  NO2        u1297(.A(men_men_n1325_), .B(men_men_n210_), .Y(men_men_n1326_));
  AOI210     u1298(.A0(men_men_n530_), .A1(men_men_n58_), .B0(men_men_n1326_), .Y(men_men_n1327_));
  OR3        u1299(.A(men_men_n1290_), .B(men_men_n638_), .C(men_men_n1289_), .Y(men_men_n1328_));
  NA3        u1300(.A(men_men_n781_), .B(men_men_n75_), .C(i), .Y(men_men_n1329_));
  AOI210     u1301(.A0(men_men_n1329_), .A1(men_men_n1298_), .B0(men_men_n1034_), .Y(men_men_n1330_));
  NO2        u1302(.A(men_men_n213_), .B(men_men_n114_), .Y(men_men_n1331_));
  NO3        u1303(.A(men_men_n1331_), .B(men_men_n1330_), .C(men_men_n1229_), .Y(men_men_n1332_));
  NA4        u1304(.A(men_men_n1332_), .B(men_men_n1328_), .C(men_men_n1327_), .D(men_men_n799_), .Y(men_men_n1333_));
  NO2        u1305(.A(g), .B(men_men_n239_), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n1022_), .B(men_men_n584_), .Y(men_men_n1335_));
  OAI210     u1307(.A0(men_men_n1335_), .A1(men_men_n1334_), .B0(men_men_n357_), .Y(men_men_n1336_));
  NA2        u1308(.A(men_men_n601_), .B(men_men_n599_), .Y(men_men_n1337_));
  NO3        u1309(.A(men_men_n80_), .B(men_men_n313_), .C(men_men_n45_), .Y(men_men_n1338_));
  NA2        u1310(.A(men_men_n1338_), .B(men_men_n581_), .Y(men_men_n1339_));
  NA3        u1311(.A(men_men_n1339_), .B(men_men_n1337_), .C(men_men_n707_), .Y(men_men_n1340_));
  OR2        u1312(.A(men_men_n1233_), .B(men_men_n1226_), .Y(men_men_n1341_));
  NO2        u1313(.A(men_men_n389_), .B(men_men_n72_), .Y(men_men_n1342_));
  AOI210     u1314(.A0(men_men_n772_), .A1(men_men_n651_), .B0(men_men_n1342_), .Y(men_men_n1343_));
  NA2        u1315(.A(men_men_n1338_), .B(men_men_n858_), .Y(men_men_n1344_));
  NA4        u1316(.A(men_men_n1344_), .B(men_men_n1343_), .C(men_men_n1341_), .D(men_men_n407_), .Y(men_men_n1345_));
  NOi41      u1317(.An(men_men_n1336_), .B(men_men_n1345_), .C(men_men_n1340_), .D(men_men_n1333_), .Y(men_men_n1346_));
  NO2        u1318(.A(men_men_n135_), .B(men_men_n45_), .Y(men_men_n1347_));
  AO220      u1319(.A0(i), .A1(men_men_n657_), .B0(men_men_n1347_), .B1(men_men_n744_), .Y(men_men_n1348_));
  NA2        u1320(.A(men_men_n1348_), .B(men_men_n357_), .Y(men_men_n1349_));
  NA2        u1321(.A(men_men_n481_), .B(men_men_n139_), .Y(men_men_n1350_));
  NO3        u1322(.A(men_men_n1147_), .B(men_men_n184_), .C(men_men_n88_), .Y(men_men_n1351_));
  AOI220     u1323(.A0(men_men_n1351_), .A1(men_men_n1350_), .B0(men_men_n1338_), .B1(men_men_n1025_), .Y(men_men_n1352_));
  NA2        u1324(.A(men_men_n1352_), .B(men_men_n1349_), .Y(men_men_n1353_));
  NO2        u1325(.A(men_men_n648_), .B(f), .Y(men_men_n1354_));
  NO4        u1326(.A(men_men_n1147_), .B(men_men_n1354_), .C(men_men_n182_), .D(men_men_n88_), .Y(men_men_n1355_));
  NO3        u1327(.A(men_men_n1355_), .B(men_men_n1353_), .C(men_men_n675_), .Y(men_men_n1356_));
  NA4        u1328(.A(men_men_n1356_), .B(men_men_n1346_), .C(men_men_n1324_), .D(men_men_n1301_), .Y(men06));
  NO2        u1329(.A(men_men_n429_), .B(men_men_n588_), .Y(men_men_n1358_));
  NO2        u1330(.A(men_men_n774_), .B(i), .Y(men_men_n1359_));
  OAI210     u1331(.A0(men_men_n1359_), .A1(men_men_n277_), .B0(men_men_n1358_), .Y(men_men_n1360_));
  NO2        u1332(.A(men_men_n231_), .B(men_men_n105_), .Y(men_men_n1361_));
  OAI210     u1333(.A0(men_men_n1361_), .A1(men_men_n1351_), .B0(men_men_n403_), .Y(men_men_n1362_));
  NO3        u1334(.A(men_men_n632_), .B(men_men_n853_), .C(men_men_n635_), .Y(men_men_n1363_));
  OR2        u1335(.A(men_men_n1363_), .B(men_men_n938_), .Y(men_men_n1364_));
  NA4        u1336(.A(men_men_n1364_), .B(men_men_n1362_), .C(men_men_n1360_), .D(men_men_n1336_), .Y(men_men_n1365_));
  NO3        u1337(.A(men_men_n1365_), .B(men_men_n1340_), .C(men_men_n265_), .Y(men_men_n1366_));
  AOI210     u1338(.A0(i), .A1(men_men_n1026_), .B0(men_men_n1334_), .Y(men_men_n1367_));
  AOI210     u1339(.A0(i), .A1(men_men_n585_), .B0(men_men_n1348_), .Y(men_men_n1368_));
  AOI210     u1340(.A0(men_men_n1368_), .A1(men_men_n1367_), .B0(men_men_n354_), .Y(men_men_n1369_));
  OAI210     u1341(.A0(men_men_n90_), .A1(men_men_n40_), .B0(men_men_n711_), .Y(men_men_n1370_));
  NA2        u1342(.A(men_men_n1370_), .B(men_men_n380_), .Y(men_men_n1371_));
  NO2        u1343(.A(men_men_n541_), .B(men_men_n180_), .Y(men_men_n1372_));
  NOi21      u1344(.An(men_men_n141_), .B(men_men_n45_), .Y(men_men_n1373_));
  AOI210     u1345(.A0(men_men_n642_), .A1(men_men_n57_), .B0(men_men_n1170_), .Y(men_men_n1374_));
  OAI210     u1346(.A0(men_men_n481_), .A1(men_men_n256_), .B0(men_men_n961_), .Y(men_men_n1375_));
  NO4        u1347(.A(men_men_n1375_), .B(men_men_n1374_), .C(men_men_n1373_), .D(men_men_n1372_), .Y(men_men_n1376_));
  OR2        u1348(.A(men_men_n633_), .B(men_men_n631_), .Y(men_men_n1377_));
  NO2        u1349(.A(men_men_n388_), .B(men_men_n140_), .Y(men_men_n1378_));
  AOI210     u1350(.A0(men_men_n1378_), .A1(men_men_n619_), .B0(men_men_n1377_), .Y(men_men_n1379_));
  NA3        u1351(.A(men_men_n1379_), .B(men_men_n1376_), .C(men_men_n1371_), .Y(men_men_n1380_));
  NO2        u1352(.A(men_men_n790_), .B(men_men_n387_), .Y(men_men_n1381_));
  NO3        u1353(.A(men_men_n713_), .B(men_men_n801_), .C(men_men_n671_), .Y(men_men_n1382_));
  NOi21      u1354(.An(men_men_n1381_), .B(men_men_n1382_), .Y(men_men_n1383_));
  AN2        u1355(.A(men_men_n1009_), .B(men_men_n681_), .Y(men_men_n1384_));
  NO4        u1356(.A(men_men_n1384_), .B(men_men_n1383_), .C(men_men_n1380_), .D(men_men_n1369_), .Y(men_men_n1385_));
  NO2        u1357(.A(men_men_n848_), .B(men_men_n288_), .Y(men_men_n1386_));
  OAI220     u1358(.A0(men_men_n774_), .A1(men_men_n47_), .B0(men_men_n231_), .B1(men_men_n650_), .Y(men_men_n1387_));
  OAI210     u1359(.A0(men_men_n288_), .A1(c), .B0(men_men_n678_), .Y(men_men_n1388_));
  AOI220     u1360(.A0(men_men_n1388_), .A1(men_men_n1387_), .B0(men_men_n1386_), .B1(men_men_n277_), .Y(men_men_n1389_));
  NO3        u1361(.A(men_men_n251_), .B(men_men_n105_), .C(men_men_n295_), .Y(men_men_n1390_));
  OAI220     u1362(.A0(men_men_n736_), .A1(men_men_n256_), .B0(men_men_n537_), .B1(men_men_n541_), .Y(men_men_n1391_));
  OAI210     u1363(.A0(l), .A1(i), .B0(k), .Y(men_men_n1392_));
  NO3        u1364(.A(men_men_n1392_), .B(men_men_n630_), .C(j), .Y(men_men_n1393_));
  NOi21      u1365(.An(men_men_n1393_), .B(men_men_n705_), .Y(men_men_n1394_));
  NO4        u1366(.A(men_men_n1394_), .B(men_men_n1391_), .C(men_men_n1390_), .D(men_men_n1173_), .Y(men_men_n1395_));
  NA4        u1367(.A(men_men_n839_), .B(men_men_n838_), .C(men_men_n458_), .D(men_men_n930_), .Y(men_men_n1396_));
  NAi31      u1368(.An(men_men_n790_), .B(men_men_n1396_), .C(men_men_n209_), .Y(men_men_n1397_));
  NA4        u1369(.A(men_men_n1397_), .B(men_men_n1395_), .C(men_men_n1389_), .D(men_men_n1270_), .Y(men_men_n1398_));
  NOi31      u1370(.An(men_men_n1363_), .B(men_men_n485_), .C(men_men_n415_), .Y(men_men_n1399_));
  OR3        u1371(.A(men_men_n1399_), .B(men_men_n827_), .C(men_men_n569_), .Y(men_men_n1400_));
  OR3        u1372(.A(men_men_n391_), .B(men_men_n231_), .C(men_men_n650_), .Y(men_men_n1401_));
  AOI210     u1373(.A0(men_men_n601_), .A1(men_men_n469_), .B0(men_men_n393_), .Y(men_men_n1402_));
  NA2        u1374(.A(men_men_n1393_), .B(men_men_n835_), .Y(men_men_n1403_));
  NA4        u1375(.A(men_men_n1403_), .B(men_men_n1402_), .C(men_men_n1401_), .D(men_men_n1400_), .Y(men_men_n1404_));
  AOI220     u1376(.A0(men_men_n1381_), .A1(men_men_n800_), .B0(men_men_n1378_), .B1(men_men_n245_), .Y(men_men_n1405_));
  NO4        u1377(.A(men_men_n983_), .B(men_men_n928_), .C(men_men_n526_), .D(men_men_n505_), .Y(men_men_n1406_));
  NA3        u1378(.A(men_men_n1406_), .B(men_men_n1405_), .C(men_men_n1344_), .Y(men_men_n1407_));
  NAi21      u1379(.An(j), .B(i), .Y(men_men_n1408_));
  NO4        u1380(.A(men_men_n1354_), .B(men_men_n1408_), .C(men_men_n464_), .D(men_men_n242_), .Y(men_men_n1409_));
  NO4        u1381(.A(men_men_n1409_), .B(men_men_n1407_), .C(men_men_n1404_), .D(men_men_n1398_), .Y(men_men_n1410_));
  NA4        u1382(.A(men_men_n1410_), .B(men_men_n1385_), .C(men_men_n1366_), .D(men_men_n1356_), .Y(men07));
  NOi21      u1383(.An(j), .B(k), .Y(men_men_n1412_));
  NA4        u1384(.A(men_men_n187_), .B(men_men_n111_), .C(men_men_n1412_), .D(f), .Y(men_men_n1413_));
  NAi32      u1385(.An(m), .Bn(b), .C(n), .Y(men_men_n1414_));
  NO3        u1386(.A(men_men_n1414_), .B(g), .C(f), .Y(men_men_n1415_));
  OAI210     u1387(.A0(men_men_n336_), .A1(men_men_n507_), .B0(men_men_n1415_), .Y(men_men_n1416_));
  NAi21      u1388(.An(f), .B(c), .Y(men_men_n1417_));
  OR2        u1389(.A(e), .B(d), .Y(men_men_n1418_));
  NOi31      u1390(.An(n), .B(m), .C(b), .Y(men_men_n1419_));
  NO3        u1391(.A(men_men_n136_), .B(men_men_n471_), .C(h), .Y(men_men_n1420_));
  NA2        u1392(.A(men_men_n1416_), .B(men_men_n1413_), .Y(men_men_n1421_));
  NOi41      u1393(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1422_));
  NA3        u1394(.A(men_men_n1422_), .B(men_men_n920_), .C(men_men_n431_), .Y(men_men_n1423_));
  NOi21      u1395(.An(h), .B(k), .Y(men_men_n1424_));
  NO2        u1396(.A(men_men_n1423_), .B(men_men_n56_), .Y(men_men_n1425_));
  NO3        u1397(.A(men_men_n1109_), .B(men_men_n152_), .C(men_men_n221_), .Y(men_men_n1426_));
  OAI210     u1398(.A0(men_men_n1149_), .A1(men_men_n1426_), .B0(men_men_n228_), .Y(men_men_n1427_));
  NO2        u1399(.A(men_men_n1427_), .B(men_men_n60_), .Y(men_men_n1428_));
  NO2        u1400(.A(k), .B(i), .Y(men_men_n1429_));
  NA2        u1401(.A(men_men_n88_), .B(men_men_n45_), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n1109_), .B(men_men_n464_), .Y(men_men_n1431_));
  NA3        u1403(.A(men_men_n1431_), .B(men_men_n1430_), .C(men_men_n221_), .Y(men_men_n1432_));
  NO2        u1404(.A(men_men_n1119_), .B(men_men_n321_), .Y(men_men_n1433_));
  NA2        u1405(.A(men_men_n570_), .B(men_men_n81_), .Y(men_men_n1434_));
  NA2        u1406(.A(men_men_n1271_), .B(men_men_n303_), .Y(men_men_n1435_));
  NA3        u1407(.A(men_men_n1435_), .B(men_men_n1434_), .C(men_men_n1432_), .Y(men_men_n1436_));
  NO4        u1408(.A(men_men_n1436_), .B(men_men_n1428_), .C(men_men_n1425_), .D(men_men_n1421_), .Y(men_men_n1437_));
  NO3        u1409(.A(e), .B(d), .C(c), .Y(men_men_n1438_));
  AOI210     u1410(.A0(men_men_n1126_), .A1(men_men_n221_), .B0(men_men_n1438_), .Y(men_men_n1439_));
  OAI210     u1411(.A0(men_men_n136_), .A1(men_men_n221_), .B0(men_men_n639_), .Y(men_men_n1440_));
  NA2        u1412(.A(men_men_n1440_), .B(men_men_n1438_), .Y(men_men_n1441_));
  NO2        u1413(.A(men_men_n1441_), .B(men_men_n1439_), .Y(men_men_n1442_));
  OR2        u1414(.A(h), .B(f), .Y(men_men_n1443_));
  NO3        u1415(.A(n), .B(m), .C(i), .Y(men_men_n1444_));
  OAI210     u1416(.A0(men_men_n1171_), .A1(men_men_n163_), .B0(men_men_n1444_), .Y(men_men_n1445_));
  NO2        u1417(.A(i), .B(g), .Y(men_men_n1446_));
  OR3        u1418(.A(men_men_n1446_), .B(men_men_n1414_), .C(men_men_n71_), .Y(men_men_n1447_));
  OAI220     u1419(.A0(men_men_n1447_), .A1(men_men_n507_), .B0(men_men_n1445_), .B1(men_men_n1443_), .Y(men_men_n1448_));
  NA3        u1420(.A(men_men_n1419_), .B(men_men_n1116_), .C(men_men_n709_), .Y(men_men_n1449_));
  NO2        u1421(.A(men_men_n1449_), .B(men_men_n45_), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1444_), .B(men_men_n677_), .Y(men_men_n1451_));
  NO2        u1423(.A(l), .B(k), .Y(men_men_n1452_));
  NOi41      u1424(.An(men_men_n574_), .B(men_men_n1452_), .C(men_men_n500_), .D(men_men_n464_), .Y(men_men_n1453_));
  NO4        u1425(.A(men_men_n1453_), .B(men_men_n1450_), .C(men_men_n1448_), .D(men_men_n1442_), .Y(men_men_n1454_));
  NO2        u1426(.A(men_men_n153_), .B(h), .Y(men_men_n1455_));
  NO2        u1427(.A(g), .B(c), .Y(men_men_n1456_));
  NA3        u1428(.A(men_men_n1456_), .B(men_men_n147_), .C(men_men_n194_), .Y(men_men_n1457_));
  NO2        u1429(.A(men_men_n1457_), .B(men_men_n1621_), .Y(men_men_n1458_));
  NA2        u1430(.A(men_men_n1458_), .B(men_men_n187_), .Y(men_men_n1459_));
  OAI210     u1431(.A0(men_men_n1424_), .A1(men_men_n220_), .B0(men_men_n1129_), .Y(men_men_n1460_));
  NO2        u1432(.A(men_men_n474_), .B(a), .Y(men_men_n1461_));
  NA3        u1433(.A(men_men_n1461_), .B(men_men_n1460_), .C(men_men_n116_), .Y(men_men_n1462_));
  NO2        u1434(.A(i), .B(h), .Y(men_men_n1463_));
  NA2        u1435(.A(men_men_n1463_), .B(men_men_n228_), .Y(men_men_n1464_));
  AOI210     u1436(.A0(men_men_n266_), .A1(men_men_n119_), .B0(men_men_n558_), .Y(men_men_n1465_));
  NO2        u1437(.A(men_men_n1465_), .B(men_men_n1464_), .Y(men_men_n1466_));
  NO2        u1438(.A(men_men_n797_), .B(men_men_n195_), .Y(men_men_n1467_));
  NOi31      u1439(.An(m), .B(n), .C(b), .Y(men_men_n1468_));
  NOi31      u1440(.An(f), .B(d), .C(c), .Y(men_men_n1469_));
  NA2        u1441(.A(men_men_n1469_), .B(men_men_n1468_), .Y(men_men_n1470_));
  INV        u1442(.A(men_men_n1470_), .Y(men_men_n1471_));
  NO3        u1443(.A(men_men_n1471_), .B(men_men_n1467_), .C(men_men_n1466_), .Y(men_men_n1472_));
  NA2        u1444(.A(men_men_n1140_), .B(men_men_n488_), .Y(men_men_n1473_));
  NO4        u1445(.A(men_men_n1473_), .B(men_men_n1116_), .C(men_men_n464_), .D(men_men_n45_), .Y(men_men_n1474_));
  NO3        u1446(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1475_));
  INV        u1447(.A(men_men_n1474_), .Y(men_men_n1476_));
  AN4        u1448(.A(men_men_n1476_), .B(men_men_n1472_), .C(men_men_n1462_), .D(men_men_n1459_), .Y(men_men_n1477_));
  NA2        u1449(.A(men_men_n1419_), .B(men_men_n400_), .Y(men_men_n1478_));
  NO2        u1450(.A(men_men_n1478_), .B(men_men_n1100_), .Y(men_men_n1479_));
  NO2        u1451(.A(men_men_n195_), .B(b), .Y(men_men_n1480_));
  AOI220     u1452(.A0(men_men_n1227_), .A1(men_men_n1480_), .B0(men_men_n1148_), .B1(men_men_n1473_), .Y(men_men_n1481_));
  NO2        u1453(.A(i), .B(men_men_n220_), .Y(men_men_n1482_));
  NA4        u1454(.A(men_men_n1201_), .B(men_men_n1482_), .C(men_men_n106_), .D(m), .Y(men_men_n1483_));
  NAi31      u1455(.An(men_men_n1479_), .B(men_men_n1483_), .C(men_men_n1481_), .Y(men_men_n1484_));
  NO4        u1456(.A(men_men_n136_), .B(g), .C(f), .D(e), .Y(men_men_n1485_));
  NA3        u1457(.A(men_men_n1429_), .B(men_men_n304_), .C(h), .Y(men_men_n1486_));
  NA2        u1458(.A(men_men_n200_), .B(men_men_n100_), .Y(men_men_n1487_));
  OR2        u1459(.A(e), .B(a), .Y(men_men_n1488_));
  NOi41      u1460(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1489_));
  NA2        u1461(.A(men_men_n1489_), .B(men_men_n116_), .Y(men_men_n1490_));
  INV        u1462(.A(men_men_n1490_), .Y(men_men_n1491_));
  OR3        u1463(.A(men_men_n569_), .B(men_men_n568_), .C(men_men_n115_), .Y(men_men_n1492_));
  NA2        u1464(.A(men_men_n1169_), .B(men_men_n428_), .Y(men_men_n1493_));
  OAI220     u1465(.A0(men_men_n1493_), .A1(men_men_n457_), .B0(men_men_n1492_), .B1(men_men_n313_), .Y(men_men_n1494_));
  AO210      u1466(.A0(men_men_n1494_), .A1(men_men_n119_), .B0(men_men_n1491_), .Y(men_men_n1495_));
  NO2        u1467(.A(men_men_n1495_), .B(men_men_n1484_), .Y(men_men_n1496_));
  NA4        u1468(.A(men_men_n1496_), .B(men_men_n1477_), .C(men_men_n1454_), .D(men_men_n1437_), .Y(men_men_n1497_));
  NO2        u1469(.A(men_men_n1185_), .B(men_men_n113_), .Y(men_men_n1498_));
  NA2        u1470(.A(men_men_n400_), .B(men_men_n56_), .Y(men_men_n1499_));
  AOI210     u1471(.A0(men_men_n1499_), .A1(men_men_n1109_), .B0(men_men_n1451_), .Y(men_men_n1500_));
  NA2        u1472(.A(men_men_n222_), .B(men_men_n187_), .Y(men_men_n1501_));
  AOI210     u1473(.A0(men_men_n1501_), .A1(men_men_n1247_), .B0(men_men_n1499_), .Y(men_men_n1502_));
  NO2        u1474(.A(men_men_n1141_), .B(men_men_n1136_), .Y(men_men_n1503_));
  NO3        u1475(.A(men_men_n1503_), .B(men_men_n1502_), .C(men_men_n1500_), .Y(men_men_n1504_));
  NO2        u1476(.A(men_men_n411_), .B(j), .Y(men_men_n1505_));
  NA3        u1477(.A(men_men_n1475_), .B(men_men_n1418_), .C(men_men_n1169_), .Y(men_men_n1506_));
  NAi41      u1478(.An(men_men_n1463_), .B(men_men_n1127_), .C(men_men_n176_), .D(men_men_n156_), .Y(men_men_n1507_));
  NA2        u1479(.A(men_men_n1507_), .B(men_men_n1506_), .Y(men_men_n1508_));
  NA3        u1480(.A(g), .B(men_men_n1505_), .C(men_men_n165_), .Y(men_men_n1509_));
  INV        u1481(.A(men_men_n1509_), .Y(men_men_n1510_));
  NO2        u1482(.A(men_men_n1510_), .B(men_men_n1508_), .Y(men_men_n1511_));
  NO3        u1483(.A(men_men_n1136_), .B(men_men_n613_), .C(g), .Y(men_men_n1512_));
  NOi21      u1484(.An(men_men_n1501_), .B(men_men_n1512_), .Y(men_men_n1513_));
  AOI210     u1485(.A0(men_men_n1513_), .A1(men_men_n1487_), .B0(men_men_n1109_), .Y(men_men_n1514_));
  OAI220     u1486(.A0(men_men_n703_), .A1(g), .B0(men_men_n231_), .B1(c), .Y(men_men_n1515_));
  AOI210     u1487(.A0(men_men_n1480_), .A1(men_men_n41_), .B0(men_men_n1515_), .Y(men_men_n1516_));
  NO2        u1488(.A(men_men_n136_), .B(l), .Y(men_men_n1517_));
  NO2        u1489(.A(men_men_n231_), .B(k), .Y(men_men_n1518_));
  OAI210     u1490(.A0(men_men_n1518_), .A1(men_men_n1463_), .B0(men_men_n1517_), .Y(men_men_n1519_));
  OAI220     u1491(.A0(men_men_n1519_), .A1(men_men_n31_), .B0(men_men_n1516_), .B1(men_men_n184_), .Y(men_men_n1520_));
  NO3        u1492(.A(men_men_n1492_), .B(men_men_n488_), .C(men_men_n371_), .Y(men_men_n1521_));
  NO3        u1493(.A(men_men_n1521_), .B(men_men_n1520_), .C(men_men_n1514_), .Y(men_men_n1522_));
  NO2        u1494(.A(men_men_n49_), .B(men_men_n613_), .Y(men_men_n1523_));
  NO3        u1495(.A(men_men_n1151_), .B(men_men_n1418_), .C(men_men_n49_), .Y(men_men_n1524_));
  AOI220     u1496(.A0(men_men_n1524_), .A1(men_men_n221_), .B0(men_men_n1152_), .B1(men_men_n1523_), .Y(men_men_n1525_));
  NO2        u1497(.A(men_men_n1136_), .B(h), .Y(men_men_n1526_));
  NA3        u1498(.A(men_men_n1526_), .B(d), .C(men_men_n1101_), .Y(men_men_n1527_));
  OAI220     u1499(.A0(men_men_n1527_), .A1(c), .B0(men_men_n1525_), .B1(j), .Y(men_men_n1528_));
  NA3        u1500(.A(men_men_n1498_), .B(men_men_n488_), .C(f), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n187_), .B(men_men_n115_), .Y(men_men_n1530_));
  NO2        u1502(.A(men_men_n1412_), .B(men_men_n42_), .Y(men_men_n1531_));
  AOI210     u1503(.A0(men_men_n116_), .A1(men_men_n40_), .B0(men_men_n1531_), .Y(men_men_n1532_));
  NO2        u1504(.A(men_men_n1532_), .B(men_men_n1529_), .Y(men_men_n1533_));
  AOI210     u1505(.A0(men_men_n553_), .A1(h), .B0(men_men_n68_), .Y(men_men_n1534_));
  NA2        u1506(.A(men_men_n1534_), .B(men_men_n1461_), .Y(men_men_n1535_));
  NO2        u1507(.A(men_men_n1408_), .B(men_men_n182_), .Y(men_men_n1536_));
  NOi21      u1508(.An(d), .B(f), .Y(men_men_n1537_));
  NO3        u1509(.A(men_men_n1469_), .B(men_men_n1537_), .C(men_men_n40_), .Y(men_men_n1538_));
  NA2        u1510(.A(men_men_n1538_), .B(men_men_n1536_), .Y(men_men_n1539_));
  NO2        u1511(.A(men_men_n1418_), .B(f), .Y(men_men_n1540_));
  NA2        u1512(.A(men_men_n1461_), .B(men_men_n1531_), .Y(men_men_n1541_));
  NO2        u1513(.A(men_men_n313_), .B(c), .Y(men_men_n1542_));
  NA2        u1514(.A(men_men_n1542_), .B(men_men_n570_), .Y(men_men_n1543_));
  NA4        u1515(.A(men_men_n1543_), .B(men_men_n1541_), .C(men_men_n1539_), .D(men_men_n1535_), .Y(men_men_n1544_));
  NO3        u1516(.A(men_men_n1544_), .B(men_men_n1533_), .C(men_men_n1528_), .Y(men_men_n1545_));
  NA4        u1517(.A(men_men_n1545_), .B(men_men_n1522_), .C(men_men_n1511_), .D(men_men_n1504_), .Y(men_men_n1546_));
  NO3        u1518(.A(men_men_n1140_), .B(men_men_n1126_), .C(men_men_n40_), .Y(men_men_n1547_));
  OAI220     u1519(.A0(men_men_n488_), .A1(men_men_n313_), .B0(men_men_n135_), .B1(men_men_n59_), .Y(men_men_n1548_));
  OAI210     u1520(.A0(men_men_n1548_), .A1(men_men_n1547_), .B0(men_men_n1433_), .Y(men_men_n1549_));
  OAI210     u1521(.A0(men_men_n1485_), .A1(men_men_n1419_), .B0(men_men_n935_), .Y(men_men_n1550_));
  OAI220     u1522(.A0(men_men_n1098_), .A1(men_men_n136_), .B0(men_men_n703_), .B1(men_men_n182_), .Y(men_men_n1551_));
  NA2        u1523(.A(men_men_n1551_), .B(men_men_n656_), .Y(men_men_n1552_));
  NA3        u1524(.A(men_men_n1552_), .B(men_men_n1550_), .C(men_men_n1549_), .Y(men_men_n1553_));
  NA3        u1525(.A(men_men_n1149_), .B(men_men_n111_), .C(men_men_n228_), .Y(men_men_n1554_));
  OAI220     u1526(.A0(men_men_n157_), .A1(men_men_n189_), .B0(men_men_n471_), .B1(g), .Y(men_men_n1555_));
  OAI210     u1527(.A0(men_men_n1555_), .A1(men_men_n113_), .B0(men_men_n1468_), .Y(men_men_n1556_));
  NA2        u1528(.A(men_men_n1556_), .B(men_men_n1554_), .Y(men_men_n1557_));
  NO2        u1529(.A(men_men_n1557_), .B(men_men_n1553_), .Y(men_men_n1558_));
  NO2        u1530(.A(men_men_n1417_), .B(e), .Y(men_men_n1559_));
  NA2        u1531(.A(men_men_n1559_), .B(men_men_n426_), .Y(men_men_n1560_));
  OR3        u1532(.A(men_men_n1518_), .B(men_men_n1271_), .C(men_men_n136_), .Y(men_men_n1561_));
  NO2        u1533(.A(men_men_n1561_), .B(men_men_n1560_), .Y(men_men_n1562_));
  NO3        u1534(.A(men_men_n1492_), .B(men_men_n371_), .C(a), .Y(men_men_n1563_));
  NO2        u1535(.A(men_men_n1563_), .B(men_men_n1562_), .Y(men_men_n1564_));
  INV        u1536(.A(men_men_n1524_), .Y(men_men_n1565_));
  NO2        u1537(.A(men_men_n1488_), .B(f), .Y(men_men_n1566_));
  AOI210     u1538(.A0(men_men_n1180_), .A1(a), .B0(men_men_n1566_), .Y(men_men_n1567_));
  OAI220     u1539(.A0(men_men_n1567_), .A1(men_men_n68_), .B0(men_men_n1565_), .B1(men_men_n220_), .Y(men_men_n1568_));
  AOI210     u1540(.A0(men_men_n955_), .A1(men_men_n438_), .B0(men_men_n107_), .Y(men_men_n1569_));
  OR2        u1541(.A(men_men_n1569_), .B(men_men_n568_), .Y(men_men_n1570_));
  NA2        u1542(.A(men_men_n1566_), .B(men_men_n1430_), .Y(men_men_n1571_));
  OAI220     u1543(.A0(men_men_n1571_), .A1(men_men_n49_), .B0(men_men_n1570_), .B1(men_men_n182_), .Y(men_men_n1572_));
  NA4        u1544(.A(men_men_n1149_), .B(men_men_n1146_), .C(men_men_n228_), .D(men_men_n67_), .Y(men_men_n1573_));
  NA2        u1545(.A(men_men_n1420_), .B(men_men_n190_), .Y(men_men_n1574_));
  NO2        u1546(.A(men_men_n49_), .B(l), .Y(men_men_n1575_));
  OAI210     u1547(.A0(men_men_n1488_), .A1(men_men_n912_), .B0(men_men_n507_), .Y(men_men_n1576_));
  OAI210     u1548(.A0(men_men_n1576_), .A1(men_men_n1152_), .B0(men_men_n1575_), .Y(men_men_n1577_));
  NO2        u1549(.A(men_men_n261_), .B(g), .Y(men_men_n1578_));
  NO2        u1550(.A(m), .B(i), .Y(men_men_n1579_));
  AOI220     u1551(.A0(men_men_n1579_), .A1(men_men_n1455_), .B0(men_men_n1127_), .B1(men_men_n1578_), .Y(men_men_n1580_));
  NA4        u1552(.A(men_men_n1580_), .B(men_men_n1577_), .C(men_men_n1574_), .D(men_men_n1573_), .Y(men_men_n1581_));
  NO3        u1553(.A(men_men_n1581_), .B(men_men_n1572_), .C(men_men_n1568_), .Y(men_men_n1582_));
  NA3        u1554(.A(men_men_n1582_), .B(men_men_n1564_), .C(men_men_n1558_), .Y(men_men_n1583_));
  NA3        u1555(.A(men_men_n1015_), .B(men_men_n143_), .C(men_men_n46_), .Y(men_men_n1584_));
  AOI210     u1556(.A0(men_men_n154_), .A1(c), .B0(men_men_n1584_), .Y(men_men_n1585_));
  OAI210     u1557(.A0(men_men_n613_), .A1(g), .B0(men_men_n192_), .Y(men_men_n1586_));
  NA2        u1558(.A(men_men_n1586_), .B(men_men_n1526_), .Y(men_men_n1587_));
  AO210      u1559(.A0(men_men_n137_), .A1(l), .B0(men_men_n1478_), .Y(men_men_n1588_));
  NO2        u1560(.A(men_men_n71_), .B(c), .Y(men_men_n1589_));
  NO4        u1561(.A(men_men_n1443_), .B(men_men_n193_), .C(men_men_n471_), .D(men_men_n45_), .Y(men_men_n1590_));
  AOI210     u1562(.A0(men_men_n1536_), .A1(men_men_n1589_), .B0(men_men_n1590_), .Y(men_men_n1591_));
  NA3        u1563(.A(men_men_n1591_), .B(men_men_n1588_), .C(men_men_n1587_), .Y(men_men_n1592_));
  NO2        u1564(.A(men_men_n1592_), .B(men_men_n1585_), .Y(men_men_n1593_));
  NO4        u1565(.A(men_men_n231_), .B(men_men_n193_), .C(men_men_n266_), .D(k), .Y(men_men_n1594_));
  AOI210     u1566(.A0(men_men_n163_), .A1(men_men_n56_), .B0(men_men_n1559_), .Y(men_men_n1595_));
  NO2        u1567(.A(men_men_n1595_), .B(men_men_n1530_), .Y(men_men_n1596_));
  NO2        u1568(.A(men_men_n1584_), .B(men_men_n113_), .Y(men_men_n1597_));
  NOi21      u1569(.An(men_men_n1420_), .B(e), .Y(men_men_n1598_));
  NO4        u1570(.A(men_men_n1598_), .B(men_men_n1597_), .C(men_men_n1596_), .D(men_men_n1594_), .Y(men_men_n1599_));
  AO220      u1571(.A0(men_men_n1149_), .A1(men_men_n1134_), .B0(men_men_n1426_), .B1(men_men_n805_), .Y(men_men_n1600_));
  AOI220     u1572(.A0(men_men_n1579_), .A1(men_men_n677_), .B0(men_men_n1113_), .B1(men_men_n166_), .Y(men_men_n1601_));
  NOi31      u1573(.An(men_men_n30_), .B(men_men_n1601_), .C(n), .Y(men_men_n1602_));
  AOI210     u1574(.A0(men_men_n1600_), .A1(men_men_n1227_), .B0(men_men_n1602_), .Y(men_men_n1603_));
  NO2        u1575(.A(men_men_n1529_), .B(men_men_n68_), .Y(men_men_n1604_));
  NO2        u1576(.A(men_men_n1429_), .B(men_men_n121_), .Y(men_men_n1605_));
  NO2        u1577(.A(men_men_n1605_), .B(men_men_n1478_), .Y(men_men_n1606_));
  NO2        u1578(.A(men_men_n1606_), .B(men_men_n1604_), .Y(men_men_n1607_));
  NA4        u1579(.A(men_men_n1607_), .B(men_men_n1603_), .C(men_men_n1599_), .D(men_men_n1593_), .Y(men_men_n1608_));
  OR4        u1580(.A(men_men_n1608_), .B(men_men_n1583_), .C(men_men_n1546_), .D(men_men_n1497_), .Y(men04));
  NOi31      u1581(.An(men_men_n1485_), .B(men_men_n1486_), .C(men_men_n1103_), .Y(men_men_n1610_));
  NA2        u1582(.A(men_men_n1540_), .B(men_men_n872_), .Y(men_men_n1611_));
  NO4        u1583(.A(men_men_n1611_), .B(men_men_n1094_), .C(men_men_n508_), .D(j), .Y(men_men_n1612_));
  OR3        u1584(.A(men_men_n1612_), .B(men_men_n1610_), .C(men_men_n1117_), .Y(men_men_n1613_));
  NO3        u1585(.A(men_men_n1430_), .B(men_men_n92_), .C(k), .Y(men_men_n1614_));
  AOI210     u1586(.A0(men_men_n1614_), .A1(men_men_n1625_), .B0(men_men_n1249_), .Y(men_men_n1615_));
  NA2        u1587(.A(men_men_n1615_), .B(men_men_n1275_), .Y(men_men_n1616_));
  NO4        u1588(.A(men_men_n1616_), .B(men_men_n1613_), .C(men_men_n1125_), .D(men_men_n1108_), .Y(men_men_n1617_));
  NA4        u1589(.A(men_men_n1617_), .B(men_men_n1182_), .C(men_men_n1167_), .D(men_men_n1155_), .Y(men05));
  INV        u1590(.A(l), .Y(men_men_n1621_));
  INV        u1591(.A(f), .Y(men_men_n1622_));
  INV        u1592(.A(n), .Y(men_men_n1623_));
  INV        u1593(.A(m), .Y(men_men_n1624_));
  INV        u1594(.A(men_men_n321_), .Y(men_men_n1625_));
  INV        u1595(.A(f), .Y(men_men_n1626_));
  INV        u1596(.A(men_men_n322_), .Y(men_men_n1627_));
  INV        u1597(.A(men_men_n464_), .Y(men_men_n1628_));
  INV        u1598(.A(e), .Y(men_men_n1629_));
  INV        u1599(.A(g), .Y(men_men_n1630_));
  INV        u1600(.A(m), .Y(men_men_n1631_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule