//Benchmark atmr_9sym_175_0.125

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n133_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n119_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  INV        o002(.A(i_5_), .Y(ori_ori_n13_));
  NOi21      o003(.An(i_3_), .B(i_7_), .Y(ori_ori_n14_));
  INV        o004(.A(i_0_), .Y(ori_ori_n15_));
  NOi21      o005(.An(i_1_), .B(i_3_), .Y(ori_ori_n16_));
  INV        o006(.A(i_4_), .Y(ori_ori_n17_));
  NA2        o007(.A(i_0_), .B(ori_ori_n17_), .Y(ori_ori_n18_));
  NOi21      o008(.An(i_8_), .B(i_6_), .Y(ori_ori_n19_));
  AOI210     o009(.A0(ori_ori_n19_), .A1(i_5_), .B0(i_2_), .Y(ori_ori_n20_));
  NO2        o010(.A(ori_ori_n20_), .B(ori_ori_n18_), .Y(ori_ori_n21_));
  NA2        o011(.A(ori_ori_n21_), .B(ori_ori_n11_), .Y(ori_ori_n22_));
  NA2        o012(.A(ori_ori_n15_), .B(i_5_), .Y(ori_ori_n23_));
  INV        o013(.A(i_2_), .Y(ori_ori_n24_));
  NOi21      o014(.An(i_5_), .B(i_0_), .Y(ori_ori_n25_));
  NOi21      o015(.An(i_6_), .B(i_8_), .Y(ori_ori_n26_));
  NOi21      o016(.An(i_7_), .B(i_1_), .Y(ori_ori_n27_));
  NOi21      o017(.An(i_5_), .B(i_6_), .Y(ori_ori_n28_));
  AOI220     o018(.A0(ori_ori_n28_), .A1(ori_ori_n27_), .B0(ori_ori_n26_), .B1(ori_ori_n25_), .Y(ori_ori_n29_));
  NOi21      o019(.An(i_0_), .B(i_4_), .Y(ori_ori_n30_));
  XO2        o020(.A(i_1_), .B(i_3_), .Y(ori_ori_n31_));
  INV        o021(.A(i_1_), .Y(ori_ori_n32_));
  NOi21      o022(.An(i_3_), .B(i_0_), .Y(ori_ori_n33_));
  INV        o023(.A(i_8_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_4_), .B(i_0_), .Y(ori_ori_n35_));
  NO2        o025(.A(ori_ori_n19_), .B(ori_ori_n14_), .Y(ori_ori_n36_));
  NA2        o026(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n37_));
  NOi21      o027(.An(i_2_), .B(i_8_), .Y(ori_ori_n38_));
  NO2        o028(.A(ori_ori_n35_), .B(ori_ori_n30_), .Y(ori_ori_n39_));
  NO3        o029(.A(ori_ori_n39_), .B(ori_ori_n37_), .C(ori_ori_n36_), .Y(ori_ori_n40_));
  INV        o030(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NOi31      o031(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n42_));
  NOi21      o032(.An(i_4_), .B(i_3_), .Y(ori_ori_n43_));
  NOi21      o033(.An(i_1_), .B(i_4_), .Y(ori_ori_n44_));
  AN2        o034(.A(i_8_), .B(i_7_), .Y(ori_ori_n45_));
  NA2        o035(.A(ori_ori_n45_), .B(ori_ori_n12_), .Y(ori_ori_n46_));
  NOi21      o036(.An(i_8_), .B(i_7_), .Y(ori_ori_n47_));
  NO2        o037(.A(ori_ori_n46_), .B(ori_ori_n37_), .Y(ori_ori_n48_));
  INV        o038(.A(ori_ori_n48_), .Y(ori_ori_n49_));
  NA4        o039(.A(ori_ori_n49_), .B(ori_ori_n41_), .C(ori_ori_n29_), .D(ori_ori_n22_), .Y(ori_ori_n50_));
  INV        o040(.A(i_8_), .Y(ori_ori_n51_));
  AOI220     o041(.A0(ori_ori_n33_), .A1(i_1_), .B0(ori_ori_n31_), .B1(i_2_), .Y(ori_ori_n52_));
  NOi21      o042(.An(i_1_), .B(i_2_), .Y(ori_ori_n53_));
  NO2        o043(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n54_));
  NA2        o044(.A(ori_ori_n54_), .B(ori_ori_n13_), .Y(ori_ori_n55_));
  NA3        o045(.A(ori_ori_n47_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n56_));
  INV        o046(.A(ori_ori_n56_), .Y(ori_ori_n57_));
  NA3        o047(.A(ori_ori_n16_), .B(i_2_), .C(i_6_), .Y(ori_ori_n58_));
  INV        o048(.A(ori_ori_n58_), .Y(ori_ori_n59_));
  INV        o049(.A(i_0_), .Y(ori_ori_n60_));
  AOI220     o050(.A0(ori_ori_n60_), .A1(ori_ori_n59_), .B0(ori_ori_n57_), .B1(ori_ori_n43_), .Y(ori_ori_n61_));
  NA2        o051(.A(ori_ori_n61_), .B(ori_ori_n55_), .Y(ori_ori_n62_));
  NAi21      o052(.An(i_3_), .B(i_6_), .Y(ori_ori_n63_));
  NO2        o053(.A(ori_ori_n63_), .B(ori_ori_n34_), .Y(ori_ori_n64_));
  NOi21      o054(.An(i_7_), .B(i_8_), .Y(ori_ori_n65_));
  NOi31      o055(.An(i_6_), .B(i_5_), .C(i_7_), .Y(ori_ori_n66_));
  AOI210     o056(.A0(ori_ori_n65_), .A1(ori_ori_n12_), .B0(ori_ori_n66_), .Y(ori_ori_n67_));
  NO2        o057(.A(ori_ori_n67_), .B(ori_ori_n11_), .Y(ori_ori_n68_));
  OAI210     o058(.A0(ori_ori_n68_), .A1(ori_ori_n64_), .B0(ori_ori_n53_), .Y(ori_ori_n69_));
  NA3        o059(.A(ori_ori_n47_), .B(ori_ori_n24_), .C(i_3_), .Y(ori_ori_n70_));
  NA2        o060(.A(ori_ori_n32_), .B(i_6_), .Y(ori_ori_n71_));
  AOI210     o061(.A0(ori_ori_n71_), .A1(ori_ori_n18_), .B0(ori_ori_n70_), .Y(ori_ori_n72_));
  NA2        o062(.A(ori_ori_n53_), .B(ori_ori_n26_), .Y(ori_ori_n73_));
  INV        o063(.A(ori_ori_n72_), .Y(ori_ori_n74_));
  INV        o064(.A(i_1_), .Y(ori_ori_n75_));
  AOI220     o065(.A0(ori_ori_n75_), .A1(i_7_), .B0(ori_ori_n19_), .B1(i_5_), .Y(ori_ori_n76_));
  NOi31      o066(.An(ori_ori_n35_), .B(ori_ori_n76_), .C(i_2_), .Y(ori_ori_n77_));
  NA2        o067(.A(ori_ori_n47_), .B(ori_ori_n12_), .Y(ori_ori_n78_));
  NOi21      o068(.An(i_3_), .B(i_1_), .Y(ori_ori_n79_));
  NA2        o069(.A(ori_ori_n79_), .B(i_4_), .Y(ori_ori_n80_));
  NO2        o070(.A(ori_ori_n78_), .B(ori_ori_n80_), .Y(ori_ori_n81_));
  NO2        o071(.A(ori_ori_n81_), .B(ori_ori_n77_), .Y(ori_ori_n82_));
  NA3        o072(.A(ori_ori_n82_), .B(ori_ori_n74_), .C(ori_ori_n69_), .Y(ori_ori_n83_));
  NOi31      o073(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n84_));
  NA2        o074(.A(ori_ori_n84_), .B(i_7_), .Y(ori_ori_n85_));
  NA2        o075(.A(ori_ori_n85_), .B(ori_ori_n73_), .Y(ori_ori_n86_));
  NA2        o076(.A(ori_ori_n86_), .B(ori_ori_n30_), .Y(ori_ori_n87_));
  NO2        o077(.A(ori_ori_n56_), .B(ori_ori_n23_), .Y(ori_ori_n88_));
  NA3        o078(.A(ori_ori_n47_), .B(ori_ori_n42_), .C(i_6_), .Y(ori_ori_n89_));
  INV        o079(.A(ori_ori_n89_), .Y(ori_ori_n90_));
  NOi21      o080(.An(i_0_), .B(i_2_), .Y(ori_ori_n91_));
  NA2        o081(.A(ori_ori_n91_), .B(ori_ori_n43_), .Y(ori_ori_n92_));
  INV        o082(.A(ori_ori_n92_), .Y(ori_ori_n93_));
  NA3        o083(.A(ori_ori_n42_), .B(ori_ori_n13_), .C(i_7_), .Y(ori_ori_n94_));
  NA4        o084(.A(ori_ori_n44_), .B(ori_ori_n28_), .C(ori_ori_n15_), .D(i_8_), .Y(ori_ori_n95_));
  NA2        o085(.A(ori_ori_n95_), .B(ori_ori_n94_), .Y(ori_ori_n96_));
  NO4        o086(.A(ori_ori_n96_), .B(ori_ori_n93_), .C(ori_ori_n90_), .D(ori_ori_n88_), .Y(ori_ori_n97_));
  INV        o087(.A(ori_ori_n65_), .Y(ori_ori_n98_));
  NO2        o088(.A(ori_ori_n98_), .B(ori_ori_n71_), .Y(ori_ori_n99_));
  NO4        o089(.A(i_2_), .B(ori_ori_n17_), .C(ori_ori_n11_), .D(ori_ori_n13_), .Y(ori_ori_n100_));
  NA2        o090(.A(i_2_), .B(i_4_), .Y(ori_ori_n101_));
  INV        o091(.A(ori_ori_n101_), .Y(ori_ori_n102_));
  NO2        o092(.A(i_8_), .B(i_7_), .Y(ori_ori_n103_));
  OA210      o093(.A0(ori_ori_n102_), .A1(ori_ori_n100_), .B0(ori_ori_n103_), .Y(ori_ori_n104_));
  NA2        o094(.A(ori_ori_n79_), .B(i_0_), .Y(ori_ori_n105_));
  NO2        o095(.A(ori_ori_n105_), .B(i_4_), .Y(ori_ori_n106_));
  NO3        o096(.A(ori_ori_n106_), .B(ori_ori_n104_), .C(ori_ori_n99_), .Y(ori_ori_n107_));
  INV        o097(.A(ori_ori_n65_), .Y(ori_ori_n108_));
  NA2        o098(.A(i_2_), .B(ori_ori_n13_), .Y(ori_ori_n109_));
  INV        o099(.A(ori_ori_n35_), .Y(ori_ori_n110_));
  AOI210     o100(.A0(ori_ori_n110_), .A1(ori_ori_n109_), .B0(ori_ori_n108_), .Y(ori_ori_n111_));
  NO2        o101(.A(ori_ori_n70_), .B(ori_ori_n23_), .Y(ori_ori_n112_));
  NA3        o102(.A(ori_ori_n45_), .B(ori_ori_n32_), .C(ori_ori_n17_), .Y(ori_ori_n113_));
  NA2        o103(.A(ori_ori_n38_), .B(ori_ori_n14_), .Y(ori_ori_n114_));
  NA2        o104(.A(ori_ori_n114_), .B(ori_ori_n113_), .Y(ori_ori_n115_));
  NO3        o105(.A(ori_ori_n115_), .B(ori_ori_n112_), .C(ori_ori_n111_), .Y(ori_ori_n116_));
  NA4        o106(.A(ori_ori_n116_), .B(ori_ori_n107_), .C(ori_ori_n97_), .D(ori_ori_n87_), .Y(ori_ori_n117_));
  OR4        o107(.A(ori_ori_n117_), .B(ori_ori_n83_), .C(ori_ori_n62_), .D(ori_ori_n50_), .Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NA3        m013(.A(i_6_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n24_));
  NO2        m014(.A(mai_mai_n24_), .B(mai_mai_n22_), .Y(mai_mai_n25_));
  AOI210     m015(.A0(mai_mai_n25_), .A1(mai_mai_n11_), .B0(mai_mai_n20_), .Y(mai_mai_n26_));
  NA2        m016(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n27_));
  NA2        m017(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n28_));
  NO2        m018(.A(i_2_), .B(i_4_), .Y(mai_mai_n29_));
  NA3        m019(.A(mai_mai_n29_), .B(i_6_), .C(i_8_), .Y(mai_mai_n30_));
  AOI210     m020(.A0(mai_mai_n28_), .A1(mai_mai_n27_), .B0(mai_mai_n30_), .Y(mai_mai_n31_));
  INV        m021(.A(i_2_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_6_), .B(i_8_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_5_), .B(i_6_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_0_), .B(i_4_), .Y(mai_mai_n35_));
  XO2        m025(.A(i_1_), .B(i_3_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_7_), .B(i_5_), .Y(mai_mai_n37_));
  AN3        m027(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(mai_mai_n35_), .Y(mai_mai_n38_));
  INV        m028(.A(i_1_), .Y(mai_mai_n39_));
  NOi21      m029(.An(i_3_), .B(i_0_), .Y(mai_mai_n40_));
  NO2        m030(.A(mai_mai_n38_), .B(mai_mai_n31_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_4_), .B(i_0_), .Y(mai_mai_n42_));
  INV        m032(.A(mai_mai_n15_), .Y(mai_mai_n43_));
  NA2        m033(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n44_));
  NOi21      m034(.An(i_2_), .B(i_8_), .Y(mai_mai_n45_));
  NO3        m035(.A(mai_mai_n45_), .B(mai_mai_n42_), .C(mai_mai_n35_), .Y(mai_mai_n46_));
  NO3        m036(.A(mai_mai_n46_), .B(mai_mai_n44_), .C(mai_mai_n43_), .Y(mai_mai_n47_));
  INV        m037(.A(mai_mai_n47_), .Y(mai_mai_n48_));
  NOi31      m038(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n49_));
  NOi21      m039(.An(i_4_), .B(i_3_), .Y(mai_mai_n50_));
  NOi21      m040(.An(i_1_), .B(i_4_), .Y(mai_mai_n51_));
  AN2        m041(.A(i_8_), .B(i_7_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_8_), .B(i_7_), .Y(mai_mai_n53_));
  NA2        m043(.A(mai_mai_n45_), .B(mai_mai_n34_), .Y(mai_mai_n54_));
  NA4        m044(.A(mai_mai_n54_), .B(mai_mai_n48_), .C(mai_mai_n41_), .D(mai_mai_n26_), .Y(mai_mai_n55_));
  NA2        m045(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n56_));
  AOI220     m046(.A0(mai_mai_n40_), .A1(i_1_), .B0(mai_mai_n36_), .B1(i_2_), .Y(mai_mai_n57_));
  NOi21      m047(.An(i_1_), .B(i_2_), .Y(mai_mai_n58_));
  NO2        m048(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  INV        m049(.A(mai_mai_n59_), .Y(mai_mai_n60_));
  NOi32      m050(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n61_));
  NA2        m051(.A(mai_mai_n61_), .B(i_3_), .Y(mai_mai_n62_));
  NA3        m052(.A(mai_mai_n18_), .B(i_2_), .C(i_6_), .Y(mai_mai_n63_));
  NA2        m053(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n64_));
  NO2        m054(.A(i_0_), .B(i_4_), .Y(mai_mai_n65_));
  AOI220     m055(.A0(mai_mai_n65_), .A1(mai_mai_n64_), .B0(mai_mai_n53_), .B1(mai_mai_n50_), .Y(mai_mai_n66_));
  NA2        m056(.A(mai_mai_n66_), .B(mai_mai_n60_), .Y(mai_mai_n67_));
  NOi21      m057(.An(i_7_), .B(i_8_), .Y(mai_mai_n68_));
  AOI220     m058(.A0(mai_mai_n40_), .A1(mai_mai_n39_), .B0(mai_mai_n18_), .B1(mai_mai_n32_), .Y(mai_mai_n69_));
  NA3        m059(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n70_));
  NO2        m060(.A(mai_mai_n70_), .B(mai_mai_n69_), .Y(mai_mai_n71_));
  INV        m061(.A(mai_mai_n71_), .Y(mai_mai_n72_));
  NA3        m062(.A(mai_mai_n53_), .B(mai_mai_n32_), .C(i_3_), .Y(mai_mai_n73_));
  NA2        m063(.A(mai_mai_n39_), .B(i_6_), .Y(mai_mai_n74_));
  AOI210     m064(.A0(mai_mai_n74_), .A1(mai_mai_n22_), .B0(mai_mai_n73_), .Y(mai_mai_n75_));
  NOi21      m065(.An(i_2_), .B(i_1_), .Y(mai_mai_n76_));
  AN3        m066(.A(mai_mai_n68_), .B(mai_mai_n76_), .C(mai_mai_n42_), .Y(mai_mai_n77_));
  NAi21      m067(.An(i_6_), .B(i_0_), .Y(mai_mai_n78_));
  NA2        m068(.A(mai_mai_n51_), .B(mai_mai_n23_), .Y(mai_mai_n79_));
  NOi21      m069(.An(i_4_), .B(i_6_), .Y(mai_mai_n80_));
  NOi21      m070(.An(i_5_), .B(i_3_), .Y(mai_mai_n81_));
  NA3        m071(.A(mai_mai_n81_), .B(mai_mai_n58_), .C(mai_mai_n80_), .Y(mai_mai_n82_));
  OAI210     m072(.A0(mai_mai_n79_), .A1(mai_mai_n78_), .B0(mai_mai_n82_), .Y(mai_mai_n83_));
  NA2        m073(.A(mai_mai_n58_), .B(mai_mai_n33_), .Y(mai_mai_n84_));
  NOi21      m074(.An(mai_mai_n37_), .B(mai_mai_n84_), .Y(mai_mai_n85_));
  NO4        m075(.A(mai_mai_n85_), .B(mai_mai_n83_), .C(mai_mai_n77_), .D(mai_mai_n75_), .Y(mai_mai_n86_));
  NOi31      m076(.An(mai_mai_n42_), .B(mai_mai_n133_), .C(i_2_), .Y(mai_mai_n87_));
  NA2        m077(.A(mai_mai_n33_), .B(mai_mai_n14_), .Y(mai_mai_n88_));
  NOi21      m078(.An(i_3_), .B(i_1_), .Y(mai_mai_n89_));
  NA2        m079(.A(mai_mai_n89_), .B(i_4_), .Y(mai_mai_n90_));
  NO2        m080(.A(mai_mai_n88_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  NO2        m081(.A(mai_mai_n91_), .B(mai_mai_n87_), .Y(mai_mai_n92_));
  NA3        m082(.A(mai_mai_n92_), .B(mai_mai_n86_), .C(mai_mai_n72_), .Y(mai_mai_n93_));
  NA2        m083(.A(mai_mai_n45_), .B(mai_mai_n15_), .Y(mai_mai_n94_));
  NOi31      m084(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n95_));
  NA2        m085(.A(mai_mai_n95_), .B(i_7_), .Y(mai_mai_n96_));
  INV        m086(.A(mai_mai_n33_), .Y(mai_mai_n97_));
  NA3        m087(.A(mai_mai_n97_), .B(mai_mai_n96_), .C(mai_mai_n94_), .Y(mai_mai_n98_));
  NA2        m088(.A(mai_mai_n98_), .B(mai_mai_n35_), .Y(mai_mai_n99_));
  NA4        m089(.A(mai_mai_n52_), .B(mai_mai_n76_), .C(mai_mai_n17_), .D(mai_mai_n12_), .Y(mai_mai_n100_));
  NAi31      m090(.An(mai_mai_n78_), .B(mai_mai_n68_), .C(mai_mai_n76_), .Y(mai_mai_n101_));
  NA2        m091(.A(mai_mai_n101_), .B(mai_mai_n100_), .Y(mai_mai_n102_));
  NOi21      m092(.An(i_0_), .B(i_2_), .Y(mai_mai_n103_));
  NA3        m093(.A(mai_mai_n103_), .B(i_7_), .C(mai_mai_n80_), .Y(mai_mai_n104_));
  NA2        m094(.A(mai_mai_n50_), .B(mai_mai_n33_), .Y(mai_mai_n105_));
  NA2        m095(.A(mai_mai_n105_), .B(mai_mai_n104_), .Y(mai_mai_n106_));
  NA3        m096(.A(mai_mai_n49_), .B(i_6_), .C(i_7_), .Y(mai_mai_n107_));
  NA3        m097(.A(mai_mai_n51_), .B(mai_mai_n34_), .C(mai_mai_n17_), .Y(mai_mai_n108_));
  NA2        m098(.A(mai_mai_n108_), .B(mai_mai_n107_), .Y(mai_mai_n109_));
  NO3        m099(.A(mai_mai_n109_), .B(mai_mai_n106_), .C(mai_mai_n102_), .Y(mai_mai_n110_));
  NOi21      m100(.An(i_5_), .B(i_2_), .Y(mai_mai_n111_));
  AOI220     m101(.A0(mai_mai_n111_), .A1(mai_mai_n68_), .B0(mai_mai_n52_), .B1(mai_mai_n29_), .Y(mai_mai_n112_));
  AOI210     m102(.A0(mai_mai_n112_), .A1(mai_mai_n94_), .B0(mai_mai_n74_), .Y(mai_mai_n113_));
  NO3        m103(.A(i_2_), .B(mai_mai_n11_), .C(mai_mai_n14_), .Y(mai_mai_n114_));
  NO2        m104(.A(i_8_), .B(i_7_), .Y(mai_mai_n115_));
  AN2        m105(.A(mai_mai_n114_), .B(mai_mai_n115_), .Y(mai_mai_n116_));
  NO2        m106(.A(mai_mai_n116_), .B(mai_mai_n113_), .Y(mai_mai_n117_));
  NA2        m107(.A(mai_mai_n68_), .B(mai_mai_n12_), .Y(mai_mai_n118_));
  NA2        m108(.A(i_2_), .B(i_1_), .Y(mai_mai_n119_));
  NA2        m109(.A(mai_mai_n42_), .B(i_3_), .Y(mai_mai_n120_));
  AOI210     m110(.A0(mai_mai_n120_), .A1(mai_mai_n119_), .B0(mai_mai_n118_), .Y(mai_mai_n121_));
  NA3        m111(.A(mai_mai_n103_), .B(mai_mai_n53_), .C(mai_mai_n80_), .Y(mai_mai_n122_));
  INV        m112(.A(mai_mai_n122_), .Y(mai_mai_n123_));
  NA3        m113(.A(mai_mai_n81_), .B(mai_mai_n52_), .C(mai_mai_n39_), .Y(mai_mai_n124_));
  NOi31      m114(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n125_));
  NA2        m115(.A(mai_mai_n61_), .B(mai_mai_n125_), .Y(mai_mai_n126_));
  NA2        m116(.A(mai_mai_n126_), .B(mai_mai_n124_), .Y(mai_mai_n127_));
  NO3        m117(.A(mai_mai_n127_), .B(mai_mai_n123_), .C(mai_mai_n121_), .Y(mai_mai_n128_));
  NA4        m118(.A(mai_mai_n128_), .B(mai_mai_n117_), .C(mai_mai_n110_), .D(mai_mai_n99_), .Y(mai_mai_n129_));
  OR4        m119(.A(mai_mai_n129_), .B(mai_mai_n93_), .C(mai_mai_n67_), .D(mai_mai_n55_), .Y(mai00));
  INV        m120(.A(i_8_), .Y(mai_mai_n133_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  INV        u005(.A(i_0_), .Y(men_men_n16_));
  NOi21      u006(.An(i_1_), .B(i_3_), .Y(men_men_n17_));
  INV        u007(.A(i_4_), .Y(men_men_n18_));
  INV        u008(.A(i_7_), .Y(men_men_n19_));
  NOi21      u009(.An(i_8_), .B(i_6_), .Y(men_men_n20_));
  NOi21      u010(.An(i_1_), .B(i_8_), .Y(men_men_n21_));
  NA2        u011(.A(men_men_n21_), .B(i_2_), .Y(men_men_n22_));
  NO2        u012(.A(men_men_n22_), .B(i_4_), .Y(men_men_n23_));
  NA2        u013(.A(men_men_n23_), .B(men_men_n11_), .Y(men_men_n24_));
  NO2        u014(.A(i_2_), .B(i_4_), .Y(men_men_n25_));
  NA3        u015(.A(men_men_n25_), .B(i_6_), .C(i_8_), .Y(men_men_n26_));
  INV        u016(.A(men_men_n26_), .Y(men_men_n27_));
  INV        u017(.A(i_2_), .Y(men_men_n28_));
  NOi21      u018(.An(i_5_), .B(i_0_), .Y(men_men_n29_));
  NOi21      u019(.An(i_5_), .B(i_6_), .Y(men_men_n30_));
  AOI220     u020(.A0(men_men_n30_), .A1(i_7_), .B0(i_6_), .B1(men_men_n29_), .Y(men_men_n31_));
  NO3        u021(.A(men_men_n31_), .B(men_men_n28_), .C(i_4_), .Y(men_men_n32_));
  NOi21      u022(.An(i_0_), .B(i_4_), .Y(men_men_n33_));
  NOi21      u023(.An(i_7_), .B(i_5_), .Y(men_men_n34_));
  AN2        u024(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  INV        u025(.A(i_1_), .Y(men_men_n36_));
  NOi21      u026(.An(i_3_), .B(i_0_), .Y(men_men_n37_));
  NA2        u027(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u028(.A(men_men_n119_), .B(men_men_n38_), .Y(men_men_n39_));
  NO4        u029(.A(men_men_n39_), .B(men_men_n35_), .C(men_men_n32_), .D(men_men_n27_), .Y(men_men_n40_));
  NOi21      u030(.An(i_4_), .B(i_0_), .Y(men_men_n41_));
  INV        u031(.A(men_men_n15_), .Y(men_men_n42_));
  NA2        u032(.A(i_1_), .B(men_men_n14_), .Y(men_men_n43_));
  NOi21      u033(.An(i_2_), .B(i_8_), .Y(men_men_n44_));
  NO2        u034(.A(men_men_n43_), .B(men_men_n42_), .Y(men_men_n45_));
  INV        u035(.A(men_men_n45_), .Y(men_men_n46_));
  NOi21      u036(.An(i_4_), .B(i_3_), .Y(men_men_n47_));
  NOi21      u037(.An(i_1_), .B(i_4_), .Y(men_men_n48_));
  INV        u038(.A(i_8_), .Y(men_men_n49_));
  NOi21      u039(.An(i_8_), .B(i_7_), .Y(men_men_n50_));
  NA3        u040(.A(men_men_n50_), .B(men_men_n47_), .C(i_6_), .Y(men_men_n51_));
  OAI210     u041(.A0(men_men_n49_), .A1(men_men_n43_), .B0(men_men_n51_), .Y(men_men_n52_));
  AOI220     u042(.A0(men_men_n52_), .A1(men_men_n28_), .B0(men_men_n47_), .B1(men_men_n30_), .Y(men_men_n53_));
  NA4        u043(.A(men_men_n53_), .B(men_men_n46_), .C(men_men_n40_), .D(men_men_n24_), .Y(men_men_n54_));
  NA2        u044(.A(i_8_), .B(i_7_), .Y(men_men_n55_));
  NO3        u045(.A(men_men_n55_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n56_));
  NA2        u046(.A(i_8_), .B(men_men_n19_), .Y(men_men_n57_));
  INV        u047(.A(i_2_), .Y(men_men_n58_));
  NOi21      u048(.An(i_1_), .B(i_2_), .Y(men_men_n59_));
  NO2        u049(.A(men_men_n58_), .B(men_men_n57_), .Y(men_men_n60_));
  OAI210     u050(.A0(men_men_n60_), .A1(men_men_n56_), .B0(men_men_n14_), .Y(men_men_n61_));
  NA3        u051(.A(men_men_n50_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n62_));
  NA3        u052(.A(men_men_n21_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n63_));
  INV        u053(.A(men_men_n63_), .Y(men_men_n64_));
  NA2        u054(.A(i_7_), .B(i_3_), .Y(men_men_n65_));
  INV        u055(.A(men_men_n65_), .Y(men_men_n66_));
  NO2        u056(.A(i_0_), .B(i_4_), .Y(men_men_n67_));
  AOI220     u057(.A0(men_men_n67_), .A1(men_men_n66_), .B0(men_men_n64_), .B1(men_men_n47_), .Y(men_men_n68_));
  NA2        u058(.A(men_men_n68_), .B(men_men_n61_), .Y(men_men_n69_));
  NAi21      u059(.An(i_3_), .B(i_6_), .Y(men_men_n70_));
  NO2        u060(.A(men_men_n70_), .B(i_0_), .Y(men_men_n71_));
  NOi21      u061(.An(i_7_), .B(i_8_), .Y(men_men_n72_));
  OAI210     u062(.A0(men_men_n72_), .A1(men_men_n71_), .B0(men_men_n59_), .Y(men_men_n73_));
  NA3        u063(.A(men_men_n20_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n74_));
  NO2        u064(.A(i_3_), .B(men_men_n74_), .Y(men_men_n75_));
  NA2        u065(.A(i_4_), .B(i_5_), .Y(men_men_n76_));
  NA3        u066(.A(men_men_n55_), .B(men_men_n17_), .C(men_men_n16_), .Y(men_men_n77_));
  NO2        u067(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NO2        u068(.A(men_men_n78_), .B(men_men_n75_), .Y(men_men_n79_));
  NA3        u069(.A(men_men_n50_), .B(men_men_n28_), .C(i_3_), .Y(men_men_n80_));
  NOi21      u070(.An(i_2_), .B(i_1_), .Y(men_men_n81_));
  NAi21      u071(.An(i_6_), .B(i_0_), .Y(men_men_n82_));
  NOi21      u072(.An(i_4_), .B(i_6_), .Y(men_men_n83_));
  NOi21      u073(.An(i_6_), .B(i_1_), .Y(men_men_n84_));
  NA2        u074(.A(men_men_n84_), .B(i_7_), .Y(men_men_n85_));
  NOi21      u075(.An(men_men_n41_), .B(men_men_n85_), .Y(men_men_n86_));
  AOI210     u076(.A0(men_men_n72_), .A1(men_men_n14_), .B0(men_men_n83_), .Y(men_men_n87_));
  NOi21      u077(.An(men_men_n37_), .B(men_men_n87_), .Y(men_men_n88_));
  NO2        u078(.A(men_men_n88_), .B(men_men_n86_), .Y(men_men_n89_));
  NA4        u079(.A(men_men_n89_), .B(men_men_n80_), .C(men_men_n79_), .D(men_men_n73_), .Y(men_men_n90_));
  NOi31      u080(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n91_));
  INV        u081(.A(men_men_n62_), .Y(men_men_n92_));
  NAi31      u082(.An(men_men_n82_), .B(men_men_n72_), .C(men_men_n81_), .Y(men_men_n93_));
  INV        u083(.A(men_men_n93_), .Y(men_men_n94_));
  NA3        u084(.A(men_men_n41_), .B(men_men_n34_), .C(men_men_n17_), .Y(men_men_n95_));
  NOi32      u085(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n96_));
  NA2        u086(.A(men_men_n96_), .B(men_men_n91_), .Y(men_men_n97_));
  NA2        u087(.A(men_men_n97_), .B(men_men_n95_), .Y(men_men_n98_));
  NA4        u088(.A(men_men_n48_), .B(men_men_n37_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n99_));
  INV        u089(.A(men_men_n99_), .Y(men_men_n100_));
  NO4        u090(.A(men_men_n100_), .B(men_men_n98_), .C(men_men_n94_), .D(men_men_n92_), .Y(men_men_n101_));
  NO3        u091(.A(i_2_), .B(men_men_n18_), .C(men_men_n11_), .Y(men_men_n102_));
  NA2        u092(.A(i_2_), .B(i_4_), .Y(men_men_n103_));
  NO2        u093(.A(men_men_n82_), .B(men_men_n103_), .Y(men_men_n104_));
  INV        u094(.A(i_7_), .Y(men_men_n105_));
  OA210      u095(.A0(men_men_n104_), .A1(men_men_n102_), .B0(men_men_n105_), .Y(men_men_n106_));
  NA3        u096(.A(i_0_), .B(i_5_), .C(men_men_n19_), .Y(men_men_n107_));
  NO2        u097(.A(men_men_n107_), .B(i_4_), .Y(men_men_n108_));
  NO2        u098(.A(men_men_n108_), .B(men_men_n106_), .Y(men_men_n109_));
  NA3        u099(.A(men_men_n44_), .B(men_men_n29_), .C(men_men_n15_), .Y(men_men_n110_));
  NOi31      u100(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n111_));
  NA2        u101(.A(i_7_), .B(men_men_n111_), .Y(men_men_n112_));
  NA2        u102(.A(men_men_n112_), .B(men_men_n110_), .Y(men_men_n113_));
  INV        u103(.A(men_men_n113_), .Y(men_men_n114_));
  NA3        u104(.A(men_men_n114_), .B(men_men_n109_), .C(men_men_n101_), .Y(men_men_n115_));
  OR4        u105(.A(men_men_n115_), .B(men_men_n90_), .C(men_men_n69_), .D(men_men_n54_), .Y(men00));
  INV        u106(.A(i_6_), .Y(men_men_n119_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule