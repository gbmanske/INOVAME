// Benchmark "top" written by ABC on Fri Jun 21 17:49:26 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n133_, new_new_n134_, new_new_n135_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n731_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n955_,
    new_new_n956_, new_new_n957_, new_new_n958_, new_new_n959_,
    new_new_n960_, new_new_n961_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA3        g031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  OAI210     g034(.A0(new_new_n56_), .A1(new_new_n55_), .B0(new_new_n54_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_12_), .Y(new_new_n58_));
  NAi21      g036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g037(.A(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA3        g039(.A(new_new_n61_), .B(new_new_n59_), .C(new_new_n31_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_10_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NAi31      g042(.An(new_new_n64_), .B(new_new_n62_), .C(new_new_n58_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n50_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NA2        g055(.A(i_2_), .B(i_8_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_9_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_7_), .Y(new_new_n80_));
  NO3        g058(.A(new_new_n80_), .B(new_new_n79_), .C(new_new_n60_), .Y(new_new_n81_));
  INV        g059(.A(i_6_), .Y(new_new_n82_));
  NO2        g060(.A(i_2_), .B(i_7_), .Y(new_new_n83_));
  INV        g061(.A(new_new_n83_), .Y(new_new_n84_));
  NA2        g062(.A(new_new_n81_), .B(new_new_n84_), .Y(new_new_n85_));
  NAi21      g063(.An(i_6_), .B(i_10_), .Y(new_new_n86_));
  NA2        g064(.A(i_6_), .B(i_9_), .Y(new_new_n87_));
  AOI210     g065(.A0(new_new_n87_), .A1(new_new_n86_), .B0(new_new_n60_), .Y(new_new_n88_));
  NA2        g066(.A(i_2_), .B(i_6_), .Y(new_new_n89_));
  NO3        g067(.A(new_new_n89_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n90_));
  NO2        g068(.A(new_new_n90_), .B(new_new_n88_), .Y(new_new_n91_));
  AOI210     g069(.A0(new_new_n91_), .A1(new_new_n85_), .B0(new_new_n77_), .Y(new_new_n92_));
  AN3        g070(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n93_));
  NAi21      g071(.An(i_6_), .B(i_11_), .Y(new_new_n94_));
  NO2        g072(.A(i_5_), .B(i_8_), .Y(new_new_n95_));
  NOi21      g073(.An(new_new_n95_), .B(new_new_n94_), .Y(new_new_n96_));
  AOI220     g074(.A0(new_new_n96_), .A1(new_new_n59_), .B0(new_new_n93_), .B1(new_new_n32_), .Y(new_new_n97_));
  INV        g075(.A(i_7_), .Y(new_new_n98_));
  NA2        g076(.A(new_new_n46_), .B(new_new_n98_), .Y(new_new_n99_));
  NO2        g077(.A(i_0_), .B(i_5_), .Y(new_new_n100_));
  NO2        g078(.A(new_new_n100_), .B(new_new_n82_), .Y(new_new_n101_));
  NA2        g079(.A(i_12_), .B(i_3_), .Y(new_new_n102_));
  INV        g080(.A(new_new_n102_), .Y(new_new_n103_));
  NA3        g081(.A(new_new_n103_), .B(new_new_n101_), .C(new_new_n99_), .Y(new_new_n104_));
  NAi21      g082(.An(i_7_), .B(i_11_), .Y(new_new_n105_));
  NO3        g083(.A(new_new_n105_), .B(new_new_n86_), .C(new_new_n51_), .Y(new_new_n106_));
  AN2        g084(.A(i_2_), .B(i_10_), .Y(new_new_n107_));
  NO2        g085(.A(new_new_n107_), .B(i_7_), .Y(new_new_n108_));
  OR2        g086(.A(new_new_n77_), .B(new_new_n55_), .Y(new_new_n109_));
  NO2        g087(.A(i_8_), .B(new_new_n98_), .Y(new_new_n110_));
  NO3        g088(.A(new_new_n110_), .B(new_new_n109_), .C(new_new_n108_), .Y(new_new_n111_));
  NA2        g089(.A(i_12_), .B(i_7_), .Y(new_new_n112_));
  NA2        g090(.A(i_11_), .B(i_12_), .Y(new_new_n113_));
  INV        g091(.A(new_new_n113_), .Y(new_new_n114_));
  NO2        g092(.A(new_new_n114_), .B(new_new_n111_), .Y(new_new_n115_));
  NAi41      g093(.An(new_new_n106_), .B(new_new_n115_), .C(new_new_n104_), .D(new_new_n97_), .Y(new_new_n116_));
  NOi21      g094(.An(i_1_), .B(i_5_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(i_11_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n98_), .B(new_new_n37_), .Y(new_new_n119_));
  NA2        g097(.A(i_7_), .B(new_new_n25_), .Y(new_new_n120_));
  NA2        g098(.A(new_new_n120_), .B(new_new_n119_), .Y(new_new_n121_));
  NO2        g099(.A(new_new_n121_), .B(new_new_n46_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n87_), .B(new_new_n86_), .Y(new_new_n123_));
  NAi21      g101(.An(i_3_), .B(i_8_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(new_new_n59_), .Y(new_new_n125_));
  NOi31      g103(.An(new_new_n125_), .B(new_new_n123_), .C(new_new_n122_), .Y(new_new_n126_));
  NO2        g104(.A(i_1_), .B(new_new_n82_), .Y(new_new_n127_));
  NO2        g105(.A(i_6_), .B(i_5_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(i_3_), .Y(new_new_n129_));
  OAI220     g107(.A0(new_new_n129_), .A1(new_new_n105_), .B0(new_new_n126_), .B1(new_new_n118_), .Y(new_new_n130_));
  NO3        g108(.A(new_new_n130_), .B(new_new_n116_), .C(new_new_n92_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(new_new_n76_), .Y(mai2));
  NO2        g110(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n133_));
  NA2        g111(.A(i_6_), .B(new_new_n25_), .Y(new_new_n134_));
  NA2        g112(.A(new_new_n134_), .B(new_new_n133_), .Y(new_new_n135_));
  NA4        g113(.A(new_new_n135_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(mai0));
  AN2        g114(.A(i_8_), .B(i_7_), .Y(new_new_n137_));
  NA2        g115(.A(new_new_n137_), .B(i_6_), .Y(new_new_n138_));
  NO2        g116(.A(i_12_), .B(i_13_), .Y(new_new_n139_));
  NAi21      g117(.An(i_5_), .B(i_11_), .Y(new_new_n140_));
  NOi21      g118(.An(new_new_n139_), .B(new_new_n140_), .Y(new_new_n141_));
  NO2        g119(.A(i_0_), .B(i_1_), .Y(new_new_n142_));
  NA2        g120(.A(i_2_), .B(i_3_), .Y(new_new_n143_));
  NO2        g121(.A(new_new_n143_), .B(i_4_), .Y(new_new_n144_));
  NA3        g122(.A(new_new_n144_), .B(new_new_n142_), .C(new_new_n141_), .Y(new_new_n145_));
  AN2        g123(.A(new_new_n139_), .B(new_new_n79_), .Y(new_new_n146_));
  NA2        g124(.A(i_1_), .B(i_5_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n70_), .B(new_new_n46_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n36_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n149_), .B(new_new_n147_), .C(i_13_), .Y(new_new_n150_));
  OR2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NO3        g129(.A(new_new_n151_), .B(new_new_n77_), .C(i_13_), .Y(new_new_n152_));
  NAi32      g130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n153_));
  NAi21      g131(.An(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  NOi21      g132(.An(i_4_), .B(i_10_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n40_), .Y(new_new_n156_));
  NO3        g134(.A(new_new_n70_), .B(i_2_), .C(i_1_), .Y(new_new_n157_));
  INV        g135(.A(new_new_n157_), .Y(new_new_n158_));
  OAI210     g136(.A0(new_new_n158_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n159_));
  NO2        g137(.A(new_new_n159_), .B(new_new_n150_), .Y(new_new_n160_));
  AOI210     g138(.A0(new_new_n160_), .A1(new_new_n145_), .B0(new_new_n138_), .Y(new_new_n161_));
  INV        g139(.A(i_1_), .Y(new_new_n162_));
  NA2        g140(.A(i_3_), .B(new_new_n48_), .Y(new_new_n163_));
  NOi21      g141(.An(i_4_), .B(i_9_), .Y(new_new_n164_));
  NOi21      g142(.An(i_11_), .B(i_13_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OR2        g144(.A(new_new_n166_), .B(new_new_n163_), .Y(new_new_n167_));
  NO2        g145(.A(i_4_), .B(i_5_), .Y(new_new_n168_));
  NAi21      g146(.An(i_12_), .B(i_11_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n169_), .B(i_13_), .Y(new_new_n170_));
  NA3        g148(.A(new_new_n170_), .B(new_new_n168_), .C(new_new_n79_), .Y(new_new_n171_));
  AOI210     g149(.A0(new_new_n171_), .A1(new_new_n167_), .B0(new_new_n162_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n70_), .B(new_new_n60_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(new_new_n46_), .Y(new_new_n174_));
  NAi31      g152(.An(new_new_n959_), .B(new_new_n146_), .C(i_11_), .Y(new_new_n175_));
  NA2        g153(.A(i_3_), .B(i_5_), .Y(new_new_n176_));
  AOI210     g154(.A0(new_new_n166_), .A1(new_new_n175_), .B0(new_new_n174_), .Y(new_new_n177_));
  NO2        g155(.A(new_new_n70_), .B(i_5_), .Y(new_new_n178_));
  NO2        g156(.A(i_13_), .B(i_10_), .Y(new_new_n179_));
  NA3        g157(.A(new_new_n179_), .B(new_new_n178_), .C(new_new_n44_), .Y(new_new_n180_));
  NO2        g158(.A(i_2_), .B(i_1_), .Y(new_new_n181_));
  NA2        g159(.A(new_new_n181_), .B(i_3_), .Y(new_new_n182_));
  NAi21      g160(.An(i_4_), .B(i_12_), .Y(new_new_n183_));
  NO3        g161(.A(new_new_n183_), .B(new_new_n182_), .C(new_new_n180_), .Y(new_new_n184_));
  NO3        g162(.A(new_new_n184_), .B(new_new_n177_), .C(new_new_n172_), .Y(new_new_n185_));
  INV        g163(.A(i_8_), .Y(new_new_n186_));
  NA2        g164(.A(new_new_n961_), .B(i_6_), .Y(new_new_n187_));
  NO3        g165(.A(i_3_), .B(new_new_n82_), .C(new_new_n48_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n188_), .B(new_new_n110_), .Y(new_new_n189_));
  NO3        g167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n190_));
  NA3        g168(.A(new_new_n190_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n191_));
  NO3        g169(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n192_));
  OAI210     g170(.A0(new_new_n93_), .A1(i_12_), .B0(new_new_n192_), .Y(new_new_n193_));
  AOI210     g171(.A0(new_new_n193_), .A1(new_new_n191_), .B0(new_new_n189_), .Y(new_new_n194_));
  NO2        g172(.A(i_3_), .B(i_8_), .Y(new_new_n195_));
  NO3        g173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n196_));
  NO2        g174(.A(i_13_), .B(i_9_), .Y(new_new_n197_));
  NA3        g175(.A(new_new_n197_), .B(i_6_), .C(new_new_n186_), .Y(new_new_n198_));
  NAi21      g176(.An(i_12_), .B(i_3_), .Y(new_new_n199_));
  BUFFER     g177(.A(new_new_n198_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n44_), .B(i_5_), .Y(new_new_n201_));
  NO3        g179(.A(i_0_), .B(i_2_), .C(new_new_n60_), .Y(new_new_n202_));
  NA3        g180(.A(new_new_n202_), .B(new_new_n201_), .C(i_10_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n203_), .B(new_new_n200_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n204_), .B(new_new_n194_), .Y(new_new_n205_));
  OAI220     g183(.A0(new_new_n205_), .A1(i_4_), .B0(new_new_n187_), .B1(new_new_n185_), .Y(new_new_n206_));
  NAi21      g184(.An(i_12_), .B(i_7_), .Y(new_new_n207_));
  NA3        g185(.A(i_13_), .B(new_new_n186_), .C(i_10_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n208_), .B(new_new_n207_), .Y(new_new_n209_));
  NA2        g187(.A(i_0_), .B(i_5_), .Y(new_new_n210_));
  NA2        g188(.A(new_new_n210_), .B(new_new_n101_), .Y(new_new_n211_));
  OAI220     g189(.A0(new_new_n211_), .A1(new_new_n182_), .B0(new_new_n174_), .B1(new_new_n129_), .Y(new_new_n212_));
  NAi31      g190(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n36_), .B(i_13_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n70_), .B(new_new_n26_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n46_), .B(new_new_n60_), .Y(new_new_n216_));
  NA3        g194(.A(new_new_n216_), .B(new_new_n215_), .C(new_new_n214_), .Y(new_new_n217_));
  INV        g195(.A(i_13_), .Y(new_new_n218_));
  NO2        g196(.A(i_12_), .B(new_new_n218_), .Y(new_new_n219_));
  NA3        g197(.A(new_new_n219_), .B(new_new_n190_), .C(new_new_n188_), .Y(new_new_n220_));
  OAI210     g198(.A0(new_new_n217_), .A1(new_new_n213_), .B0(new_new_n220_), .Y(new_new_n221_));
  AOI220     g199(.A0(new_new_n221_), .A1(new_new_n137_), .B0(new_new_n212_), .B1(new_new_n209_), .Y(new_new_n222_));
  NO2        g200(.A(i_12_), .B(new_new_n37_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n176_), .B(i_4_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n225_));
  OR2        g203(.A(i_8_), .B(i_7_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n226_), .B(new_new_n82_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n51_), .B(i_1_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n229_));
  INV        g207(.A(i_12_), .Y(new_new_n230_));
  NO2        g208(.A(new_new_n44_), .B(new_new_n230_), .Y(new_new_n231_));
  NO3        g209(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n232_));
  NA2        g210(.A(i_2_), .B(i_1_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n229_), .B(new_new_n225_), .Y(new_new_n234_));
  NO3        g212(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n235_));
  NAi21      g213(.An(i_4_), .B(i_3_), .Y(new_new_n236_));
  INV        g214(.A(new_new_n72_), .Y(new_new_n237_));
  NO2        g215(.A(i_0_), .B(i_6_), .Y(new_new_n238_));
  NOi41      g216(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n239_));
  NA2        g217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  INV        g218(.A(new_new_n234_), .Y(new_new_n241_));
  NO2        g219(.A(i_11_), .B(new_new_n218_), .Y(new_new_n242_));
  NOi21      g220(.An(i_1_), .B(i_6_), .Y(new_new_n243_));
  NAi21      g221(.An(i_3_), .B(i_7_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n230_), .B(i_9_), .Y(new_new_n245_));
  OR4        g223(.A(new_new_n245_), .B(new_new_n244_), .C(new_new_n243_), .D(new_new_n178_), .Y(new_new_n246_));
  NO2        g224(.A(i_12_), .B(i_3_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n70_), .B(i_5_), .Y(new_new_n248_));
  NA2        g226(.A(i_3_), .B(i_9_), .Y(new_new_n249_));
  NAi21      g227(.An(i_7_), .B(i_10_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n250_), .B(new_new_n249_), .Y(new_new_n251_));
  NA3        g229(.A(new_new_n251_), .B(new_new_n248_), .C(new_new_n61_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n252_), .B(new_new_n246_), .Y(new_new_n253_));
  NA3        g231(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n254_));
  INV        g232(.A(new_new_n138_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n230_), .B(i_13_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n256_), .B(new_new_n72_), .Y(new_new_n257_));
  AOI220     g235(.A0(new_new_n257_), .A1(new_new_n255_), .B0(new_new_n253_), .B1(new_new_n242_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n226_), .B(new_new_n37_), .Y(new_new_n259_));
  NA2        g237(.A(i_12_), .B(i_6_), .Y(new_new_n260_));
  OR2        g238(.A(i_13_), .B(i_9_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n236_), .B(i_2_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n242_), .B(i_9_), .Y(new_new_n263_));
  NA2        g241(.A(new_new_n148_), .B(new_new_n60_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n244_), .B(i_8_), .Y(new_new_n265_));
  NO2        g243(.A(i_6_), .B(new_new_n48_), .Y(new_new_n266_));
  NA3        g244(.A(new_new_n266_), .B(new_new_n265_), .C(i_13_), .Y(new_new_n267_));
  NA3        g245(.A(i_6_), .B(new_new_n259_), .C(new_new_n219_), .Y(new_new_n268_));
  AOI210     g246(.A0(new_new_n268_), .A1(new_new_n267_), .B0(new_new_n264_), .Y(new_new_n269_));
  INV        g247(.A(new_new_n269_), .Y(new_new_n270_));
  NA4        g248(.A(new_new_n270_), .B(new_new_n258_), .C(new_new_n241_), .D(new_new_n222_), .Y(new_new_n271_));
  NO3        g249(.A(i_12_), .B(new_new_n218_), .C(new_new_n37_), .Y(new_new_n272_));
  INV        g250(.A(new_new_n272_), .Y(new_new_n273_));
  NA2        g251(.A(i_8_), .B(new_new_n98_), .Y(new_new_n274_));
  NO3        g252(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n275_));
  AOI220     g253(.A0(new_new_n275_), .A1(new_new_n188_), .B0(i_6_), .B1(new_new_n228_), .Y(new_new_n276_));
  NO2        g254(.A(new_new_n276_), .B(new_new_n274_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n233_), .B(i_0_), .Y(new_new_n278_));
  AOI220     g256(.A0(new_new_n278_), .A1(new_new_n961_), .B0(i_1_), .B1(new_new_n137_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n266_), .B(new_new_n26_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(new_new_n279_), .Y(new_new_n281_));
  NA2        g259(.A(i_0_), .B(i_1_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n282_), .B(i_2_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n56_), .B(i_6_), .Y(new_new_n284_));
  NA2        g262(.A(new_new_n284_), .B(new_new_n283_), .Y(new_new_n285_));
  OAI210     g263(.A0(new_new_n158_), .A1(new_new_n138_), .B0(new_new_n285_), .Y(new_new_n286_));
  NO3        g264(.A(new_new_n286_), .B(new_new_n281_), .C(new_new_n277_), .Y(new_new_n287_));
  NO2        g265(.A(i_3_), .B(i_10_), .Y(new_new_n288_));
  NA3        g266(.A(new_new_n288_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n289_));
  NO2        g267(.A(i_2_), .B(new_new_n98_), .Y(new_new_n290_));
  NA2        g268(.A(i_1_), .B(new_new_n36_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n291_), .B(i_8_), .Y(new_new_n292_));
  NA2        g270(.A(new_new_n292_), .B(new_new_n290_), .Y(new_new_n293_));
  AN2        g271(.A(i_3_), .B(i_10_), .Y(new_new_n294_));
  NA3        g272(.A(new_new_n294_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n295_));
  NO2        g273(.A(i_5_), .B(new_new_n37_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n297_));
  OR2        g275(.A(new_new_n293_), .B(new_new_n289_), .Y(new_new_n298_));
  OAI220     g276(.A0(new_new_n298_), .A1(i_6_), .B0(new_new_n287_), .B1(new_new_n273_), .Y(new_new_n299_));
  NO4        g277(.A(new_new_n299_), .B(new_new_n271_), .C(new_new_n206_), .D(new_new_n161_), .Y(new_new_n300_));
  NO3        g278(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n301_));
  NO3        g279(.A(i_6_), .B(new_new_n186_), .C(i_7_), .Y(new_new_n302_));
  AOI210     g280(.A0(new_new_n186_), .A1(new_new_n233_), .B0(new_new_n163_), .Y(new_new_n303_));
  NO2        g281(.A(i_2_), .B(i_3_), .Y(new_new_n304_));
  OR2        g282(.A(i_0_), .B(i_5_), .Y(new_new_n305_));
  NA2        g283(.A(new_new_n210_), .B(new_new_n305_), .Y(new_new_n306_));
  NA4        g284(.A(new_new_n306_), .B(new_new_n227_), .C(new_new_n304_), .D(i_1_), .Y(new_new_n307_));
  NA3        g285(.A(new_new_n278_), .B(i_6_), .C(new_new_n110_), .Y(new_new_n308_));
  NAi21      g286(.An(i_8_), .B(i_7_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n309_), .B(i_6_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n151_), .B(new_new_n46_), .Y(new_new_n311_));
  NA2        g289(.A(new_new_n311_), .B(new_new_n310_), .Y(new_new_n312_));
  NA3        g290(.A(new_new_n312_), .B(new_new_n308_), .C(new_new_n307_), .Y(new_new_n313_));
  OAI210     g291(.A0(new_new_n313_), .A1(new_new_n303_), .B0(i_4_), .Y(new_new_n314_));
  NO2        g292(.A(i_12_), .B(i_10_), .Y(new_new_n315_));
  NOi21      g293(.An(i_5_), .B(i_0_), .Y(new_new_n316_));
  NA4        g294(.A(new_new_n80_), .B(new_new_n36_), .C(new_new_n82_), .D(i_8_), .Y(new_new_n317_));
  NO2        g295(.A(i_6_), .B(i_8_), .Y(new_new_n318_));
  NOi21      g296(.An(i_0_), .B(i_2_), .Y(new_new_n319_));
  AN2        g297(.A(new_new_n319_), .B(new_new_n318_), .Y(new_new_n320_));
  NO2        g298(.A(i_1_), .B(i_7_), .Y(new_new_n321_));
  AO220      g299(.A0(new_new_n321_), .A1(new_new_n320_), .B0(new_new_n310_), .B1(new_new_n228_), .Y(new_new_n322_));
  NA3        g300(.A(new_new_n322_), .B(i_4_), .C(i_5_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n323_), .B(new_new_n314_), .Y(new_new_n324_));
  INV        g302(.A(i_6_), .Y(new_new_n325_));
  INV        g303(.A(new_new_n306_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n100_), .B(new_new_n120_), .Y(new_new_n327_));
  OAI210     g305(.A0(new_new_n327_), .A1(new_new_n326_), .B0(i_3_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n282_), .B(new_new_n78_), .Y(new_new_n329_));
  NA2        g307(.A(new_new_n329_), .B(new_new_n128_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n89_), .B(new_new_n186_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n331_), .B(new_new_n60_), .Y(new_new_n332_));
  AOI210     g310(.A0(new_new_n332_), .A1(new_new_n330_), .B0(i_7_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n186_), .B(i_9_), .Y(new_new_n334_));
  NO3        g312(.A(new_new_n334_), .B(new_new_n333_), .C(new_new_n281_), .Y(new_new_n335_));
  AOI210     g313(.A0(new_new_n335_), .A1(new_new_n328_), .B0(new_new_n156_), .Y(new_new_n336_));
  AOI210     g314(.A0(new_new_n324_), .A1(new_new_n301_), .B0(new_new_n336_), .Y(new_new_n337_));
  NOi32      g315(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n338_));
  INV        g316(.A(new_new_n338_), .Y(new_new_n339_));
  NAi21      g317(.An(i_0_), .B(i_6_), .Y(new_new_n340_));
  NAi21      g318(.An(i_1_), .B(i_5_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n341_), .B(new_new_n340_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n342_), .B(new_new_n25_), .Y(new_new_n343_));
  OAI210     g321(.A0(new_new_n343_), .A1(new_new_n153_), .B0(new_new_n240_), .Y(new_new_n344_));
  NAi41      g322(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n153_), .B(new_new_n151_), .Y(new_new_n346_));
  NOi32      g324(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n347_));
  NO2        g325(.A(i_1_), .B(new_new_n98_), .Y(new_new_n348_));
  NAi21      g326(.An(i_3_), .B(i_4_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(i_9_), .Y(new_new_n350_));
  AN2        g328(.A(i_6_), .B(i_7_), .Y(new_new_n351_));
  OAI210     g329(.A0(new_new_n351_), .A1(new_new_n348_), .B0(new_new_n350_), .Y(new_new_n352_));
  NA2        g330(.A(i_2_), .B(i_7_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n349_), .B(i_10_), .Y(new_new_n354_));
  NA3        g332(.A(new_new_n354_), .B(new_new_n353_), .C(new_new_n238_), .Y(new_new_n355_));
  AOI210     g333(.A0(new_new_n355_), .A1(new_new_n352_), .B0(new_new_n178_), .Y(new_new_n356_));
  AOI210     g334(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n357_));
  OAI210     g335(.A0(new_new_n357_), .A1(new_new_n181_), .B0(new_new_n354_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n358_), .B(i_5_), .Y(new_new_n359_));
  NO4        g337(.A(new_new_n359_), .B(new_new_n356_), .C(new_new_n346_), .D(new_new_n344_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n360_), .B(new_new_n339_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n56_), .B(new_new_n25_), .Y(new_new_n362_));
  AN2        g340(.A(i_12_), .B(i_5_), .Y(new_new_n363_));
  NO2        g341(.A(i_4_), .B(new_new_n26_), .Y(new_new_n364_));
  NA2        g342(.A(new_new_n364_), .B(new_new_n363_), .Y(new_new_n365_));
  NO2        g343(.A(i_11_), .B(i_6_), .Y(new_new_n366_));
  NA3        g344(.A(new_new_n366_), .B(new_new_n311_), .C(new_new_n218_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(new_new_n365_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n236_), .B(i_5_), .Y(new_new_n369_));
  NO2        g347(.A(i_5_), .B(i_10_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n139_), .B(new_new_n45_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n371_), .B(new_new_n236_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n372_), .B(new_new_n362_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n374_));
  INV        g352(.A(new_new_n368_), .Y(new_new_n375_));
  NO3        g353(.A(new_new_n82_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n376_));
  NO2        g354(.A(i_11_), .B(i_12_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n370_), .B(new_new_n230_), .Y(new_new_n378_));
  NA3        g356(.A(new_new_n110_), .B(i_4_), .C(i_11_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n213_), .Y(new_new_n380_));
  NAi21      g358(.An(i_13_), .B(i_0_), .Y(new_new_n381_));
  INV        g359(.A(new_new_n381_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n380_), .B(new_new_n382_), .Y(new_new_n383_));
  NA3        g361(.A(new_new_n383_), .B(new_new_n375_), .C(new_new_n373_), .Y(new_new_n384_));
  NO3        g362(.A(i_1_), .B(i_12_), .C(new_new_n82_), .Y(new_new_n385_));
  NO2        g363(.A(i_0_), .B(i_11_), .Y(new_new_n386_));
  INV        g364(.A(i_5_), .Y(new_new_n387_));
  AN2        g365(.A(i_1_), .B(i_6_), .Y(new_new_n388_));
  NOi21      g366(.An(i_2_), .B(i_12_), .Y(new_new_n389_));
  NA2        g367(.A(new_new_n389_), .B(new_new_n388_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n387_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n137_), .B(i_9_), .Y(new_new_n392_));
  NO2        g370(.A(new_new_n392_), .B(i_4_), .Y(new_new_n393_));
  NA2        g371(.A(new_new_n391_), .B(new_new_n393_), .Y(new_new_n394_));
  NAi21      g372(.An(i_9_), .B(i_4_), .Y(new_new_n395_));
  OR2        g373(.A(i_13_), .B(i_10_), .Y(new_new_n396_));
  NO3        g374(.A(new_new_n396_), .B(new_new_n113_), .C(new_new_n395_), .Y(new_new_n397_));
  OR2        g375(.A(new_new_n208_), .B(new_new_n207_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n98_), .B(new_new_n25_), .Y(new_new_n399_));
  NA2        g377(.A(new_new_n272_), .B(new_new_n399_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n266_), .B(new_new_n202_), .Y(new_new_n401_));
  OAI220     g379(.A0(new_new_n401_), .A1(new_new_n398_), .B0(new_new_n400_), .B1(new_new_n100_), .Y(new_new_n402_));
  INV        g380(.A(new_new_n402_), .Y(new_new_n403_));
  AOI210     g381(.A0(new_new_n403_), .A1(new_new_n394_), .B0(new_new_n26_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n308_), .B(new_new_n307_), .Y(new_new_n405_));
  AOI220     g383(.A0(new_new_n284_), .A1(new_new_n275_), .B0(new_new_n278_), .B1(i_6_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n406_), .B(new_new_n163_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n176_), .B(new_new_n82_), .Y(new_new_n408_));
  AOI220     g386(.A0(new_new_n408_), .A1(new_new_n283_), .B0(i_6_), .B1(new_new_n202_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n409_), .B(new_new_n274_), .Y(new_new_n410_));
  NO3        g388(.A(new_new_n410_), .B(new_new_n407_), .C(new_new_n405_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n188_), .B(new_new_n93_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n311_), .B(new_new_n82_), .Y(new_new_n413_));
  AOI210     g391(.A0(new_new_n413_), .A1(new_new_n412_), .B0(new_new_n309_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n186_), .B(i_10_), .Y(new_new_n415_));
  NA3        g393(.A(new_new_n248_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n284_), .B(new_new_n228_), .Y(new_new_n417_));
  OAI220     g395(.A0(new_new_n417_), .A1(new_new_n176_), .B0(new_new_n416_), .B1(new_new_n415_), .Y(new_new_n418_));
  NA3        g396(.A(new_new_n321_), .B(new_new_n320_), .C(i_5_), .Y(new_new_n419_));
  INV        g397(.A(new_new_n302_), .Y(new_new_n420_));
  OAI210     g398(.A0(new_new_n420_), .A1(new_new_n182_), .B0(new_new_n419_), .Y(new_new_n421_));
  NO3        g399(.A(new_new_n421_), .B(new_new_n418_), .C(new_new_n414_), .Y(new_new_n422_));
  AOI210     g400(.A0(new_new_n422_), .A1(new_new_n411_), .B0(new_new_n263_), .Y(new_new_n423_));
  NO4        g401(.A(new_new_n423_), .B(new_new_n404_), .C(new_new_n384_), .D(new_new_n361_), .Y(new_new_n424_));
  NO2        g402(.A(new_new_n60_), .B(i_4_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n70_), .B(i_13_), .Y(new_new_n426_));
  NO2        g404(.A(i_10_), .B(i_9_), .Y(new_new_n427_));
  NAi21      g405(.An(i_12_), .B(i_8_), .Y(new_new_n428_));
  NO2        g406(.A(new_new_n428_), .B(i_3_), .Y(new_new_n429_));
  INV        g407(.A(i_0_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n260_), .B(new_new_n94_), .Y(new_new_n431_));
  NA2        g409(.A(i_8_), .B(i_9_), .Y(new_new_n432_));
  NO3        g410(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n433_));
  NA3        g411(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n434_));
  OR2        g412(.A(new_new_n282_), .B(new_new_n198_), .Y(new_new_n435_));
  BUFFER     g413(.A(new_new_n285_), .Y(new_new_n436_));
  OA220      g414(.A0(new_new_n436_), .A1(new_new_n156_), .B0(new_new_n435_), .B1(new_new_n225_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n93_), .B(i_13_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n408_), .B(new_new_n362_), .Y(new_new_n439_));
  NO2        g417(.A(i_2_), .B(i_13_), .Y(new_new_n440_));
  NA3        g418(.A(new_new_n440_), .B(new_new_n155_), .C(new_new_n96_), .Y(new_new_n441_));
  OAI220     g419(.A0(new_new_n441_), .A1(new_new_n230_), .B0(new_new_n439_), .B1(new_new_n438_), .Y(new_new_n442_));
  NO3        g420(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n443_));
  NO2        g421(.A(i_6_), .B(i_7_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n444_), .B(new_new_n443_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n70_), .B(i_3_), .Y(new_new_n446_));
  NOi21      g424(.An(i_2_), .B(i_7_), .Y(new_new_n447_));
  NAi31      g425(.An(i_11_), .B(new_new_n447_), .C(new_new_n446_), .Y(new_new_n448_));
  INV        g426(.A(new_new_n396_), .Y(new_new_n449_));
  NA3        g427(.A(new_new_n449_), .B(new_new_n425_), .C(new_new_n72_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n450_), .B(new_new_n448_), .Y(new_new_n451_));
  NO2        g429(.A(i_6_), .B(i_10_), .Y(new_new_n452_));
  NA4        g430(.A(new_new_n452_), .B(new_new_n301_), .C(i_8_), .D(new_new_n230_), .Y(new_new_n453_));
  NO2        g431(.A(new_new_n453_), .B(new_new_n149_), .Y(new_new_n454_));
  NA3        g432(.A(new_new_n239_), .B(new_new_n165_), .C(new_new_n128_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n151_), .B(i_3_), .Y(new_new_n457_));
  NAi31      g435(.An(new_new_n456_), .B(new_new_n457_), .C(new_new_n219_), .Y(new_new_n458_));
  NA3        g436(.A(new_new_n374_), .B(new_new_n173_), .C(new_new_n144_), .Y(new_new_n459_));
  NA3        g437(.A(new_new_n459_), .B(new_new_n458_), .C(new_new_n455_), .Y(new_new_n460_));
  NO4        g438(.A(new_new_n460_), .B(new_new_n454_), .C(new_new_n451_), .D(new_new_n442_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n433_), .B(new_new_n370_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n462_), .B(new_new_n217_), .Y(new_new_n463_));
  NAi21      g441(.An(new_new_n208_), .B(new_new_n377_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n26_), .B(i_5_), .Y(new_new_n465_));
  NO2        g443(.A(i_0_), .B(new_new_n82_), .Y(new_new_n466_));
  NA3        g444(.A(new_new_n466_), .B(new_new_n465_), .C(new_new_n137_), .Y(new_new_n467_));
  OR3        g445(.A(new_new_n291_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n468_), .B(new_new_n467_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n27_), .B(i_10_), .Y(new_new_n470_));
  NA2        g448(.A(new_new_n301_), .B(new_new_n232_), .Y(new_new_n471_));
  OAI220     g449(.A0(new_new_n471_), .A1(new_new_n416_), .B0(new_new_n470_), .B1(new_new_n438_), .Y(new_new_n472_));
  NA4        g450(.A(new_new_n294_), .B(new_new_n216_), .C(new_new_n70_), .D(new_new_n230_), .Y(new_new_n473_));
  NO2        g451(.A(new_new_n473_), .B(new_new_n445_), .Y(new_new_n474_));
  NO4        g452(.A(new_new_n474_), .B(new_new_n472_), .C(new_new_n469_), .D(new_new_n463_), .Y(new_new_n475_));
  NA3        g453(.A(new_new_n475_), .B(new_new_n461_), .C(new_new_n437_), .Y(new_new_n476_));
  NA3        g454(.A(new_new_n294_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n477_));
  INV        g455(.A(new_new_n477_), .Y(new_new_n478_));
  BUFFER     g456(.A(new_new_n275_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n479_), .B(new_new_n478_), .Y(new_new_n480_));
  INV        g458(.A(new_new_n157_), .Y(new_new_n481_));
  OAI210     g459(.A0(new_new_n481_), .A1(new_new_n225_), .B0(new_new_n295_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n482_), .B(new_new_n310_), .Y(new_new_n483_));
  NA2        g461(.A(new_new_n363_), .B(new_new_n218_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n351_), .B(new_new_n347_), .Y(new_new_n485_));
  OR2        g463(.A(new_new_n484_), .B(new_new_n485_), .Y(new_new_n486_));
  NO2        g464(.A(new_new_n36_), .B(i_8_), .Y(new_new_n487_));
  AOI210     g465(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n397_), .Y(new_new_n488_));
  NA2        g466(.A(new_new_n488_), .B(new_new_n486_), .Y(new_new_n489_));
  INV        g467(.A(new_new_n489_), .Y(new_new_n490_));
  NO2        g468(.A(i_7_), .B(new_new_n191_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n176_), .B(new_new_n82_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n492_), .B(new_new_n491_), .Y(new_new_n493_));
  NA4        g471(.A(new_new_n493_), .B(new_new_n490_), .C(new_new_n483_), .D(new_new_n480_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n369_), .B(new_new_n283_), .Y(new_new_n495_));
  OAI210     g473(.A0(new_new_n365_), .A1(new_new_n162_), .B0(new_new_n495_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n958_), .B(new_new_n218_), .Y(new_new_n497_));
  NA2        g475(.A(new_new_n452_), .B(new_new_n27_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n498_), .B(new_new_n497_), .Y(new_new_n499_));
  NOi31      g477(.An(new_new_n302_), .B(new_new_n396_), .C(new_new_n38_), .Y(new_new_n500_));
  OAI210     g478(.A0(new_new_n500_), .A1(new_new_n499_), .B0(new_new_n496_), .Y(new_new_n501_));
  NO2        g479(.A(i_8_), .B(i_7_), .Y(new_new_n502_));
  OAI210     g480(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n503_), .B(new_new_n216_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n228_), .B(new_new_n197_), .Y(new_new_n505_));
  OAI220     g483(.A0(new_new_n505_), .A1(new_new_n176_), .B0(new_new_n504_), .B1(new_new_n236_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n44_), .B(i_10_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(i_6_), .Y(new_new_n508_));
  NA3        g486(.A(new_new_n508_), .B(new_new_n506_), .C(new_new_n502_), .Y(new_new_n509_));
  AOI220     g487(.A0(new_new_n408_), .A1(new_new_n311_), .B0(i_2_), .B1(new_new_n238_), .Y(new_new_n510_));
  OAI220     g488(.A0(new_new_n510_), .A1(new_new_n256_), .B0(new_new_n438_), .B1(new_new_n129_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n511_), .B(new_new_n259_), .Y(new_new_n512_));
  NOi31      g490(.An(new_new_n278_), .B(new_new_n289_), .C(new_new_n959_), .Y(new_new_n513_));
  NO2        g491(.A(new_new_n214_), .B(new_new_n44_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n151_), .B(i_5_), .Y(new_new_n515_));
  NA2        g493(.A(new_new_n515_), .B(new_new_n304_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n516_), .B(new_new_n514_), .Y(new_new_n517_));
  OAI210     g495(.A0(new_new_n517_), .A1(new_new_n513_), .B0(new_new_n433_), .Y(new_new_n518_));
  NA4        g496(.A(new_new_n518_), .B(new_new_n512_), .C(new_new_n509_), .D(new_new_n501_), .Y(new_new_n519_));
  NA3        g497(.A(new_new_n210_), .B(new_new_n68_), .C(new_new_n44_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n272_), .B(new_new_n80_), .Y(new_new_n521_));
  AOI210     g499(.A0(new_new_n520_), .A1(new_new_n330_), .B0(new_new_n521_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n56_), .B(new_new_n167_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n524_));
  NA2        g502(.A(new_new_n427_), .B(new_new_n214_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n524_), .B(new_new_n525_), .Y(new_new_n526_));
  NO3        g504(.A(new_new_n526_), .B(new_new_n523_), .C(new_new_n522_), .Y(new_new_n527_));
  NO4        g505(.A(new_new_n243_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n528_));
  NO3        g506(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n529_));
  NO2        g507(.A(new_new_n226_), .B(new_new_n36_), .Y(new_new_n530_));
  AN2        g508(.A(new_new_n530_), .B(new_new_n529_), .Y(new_new_n531_));
  OA210      g509(.A0(new_new_n531_), .A1(new_new_n528_), .B0(new_new_n338_), .Y(new_new_n532_));
  NO2        g510(.A(new_new_n396_), .B(i_1_), .Y(new_new_n533_));
  NOi31      g511(.An(new_new_n533_), .B(new_new_n431_), .C(new_new_n70_), .Y(new_new_n534_));
  AN3        g512(.A(new_new_n534_), .B(new_new_n393_), .C(i_2_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n406_), .B(new_new_n171_), .Y(new_new_n536_));
  NO3        g514(.A(new_new_n536_), .B(new_new_n535_), .C(new_new_n532_), .Y(new_new_n537_));
  NOi21      g515(.An(i_10_), .B(i_6_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n112_), .B(new_new_n23_), .Y(new_new_n539_));
  NA2        g517(.A(new_new_n302_), .B(new_new_n157_), .Y(new_new_n540_));
  AOI220     g518(.A0(new_new_n540_), .A1(new_new_n417_), .B0(new_new_n166_), .B1(new_new_n175_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n190_), .B(new_new_n37_), .Y(new_new_n542_));
  NOi31      g520(.An(new_new_n141_), .B(new_new_n542_), .C(new_new_n317_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n543_), .B(new_new_n541_), .Y(new_new_n544_));
  INV        g522(.A(new_new_n304_), .Y(new_new_n545_));
  NO2        g523(.A(i_12_), .B(new_new_n82_), .Y(new_new_n546_));
  NO3        g524(.A(i_4_), .B(new_new_n325_), .C(new_new_n289_), .Y(new_new_n547_));
  OR2        g525(.A(i_2_), .B(i_5_), .Y(new_new_n548_));
  OR2        g526(.A(new_new_n548_), .B(new_new_n388_), .Y(new_new_n549_));
  NA2        g527(.A(new_new_n353_), .B(new_new_n238_), .Y(new_new_n550_));
  AOI210     g528(.A0(new_new_n550_), .A1(new_new_n549_), .B0(new_new_n464_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n551_), .B(new_new_n547_), .Y(new_new_n552_));
  NA4        g530(.A(new_new_n552_), .B(new_new_n544_), .C(new_new_n537_), .D(new_new_n527_), .Y(new_new_n553_));
  NO4        g531(.A(new_new_n553_), .B(new_new_n519_), .C(new_new_n494_), .D(new_new_n476_), .Y(new_new_n554_));
  NA4        g532(.A(new_new_n554_), .B(new_new_n424_), .C(new_new_n337_), .D(new_new_n300_), .Y(mai7));
  NO2        g533(.A(new_new_n89_), .B(new_new_n52_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n452_), .B(new_new_n80_), .Y(new_new_n557_));
  NA2        g535(.A(i_11_), .B(new_new_n186_), .Y(new_new_n558_));
  NA3        g536(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n230_), .B(i_4_), .Y(new_new_n560_));
  NA2        g538(.A(new_new_n560_), .B(i_8_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n102_), .B(new_new_n559_), .Y(new_new_n562_));
  NA2        g540(.A(i_2_), .B(new_new_n82_), .Y(new_new_n563_));
  OAI210     g541(.A0(new_new_n83_), .A1(new_new_n195_), .B0(new_new_n196_), .Y(new_new_n564_));
  NO2        g542(.A(i_7_), .B(new_new_n37_), .Y(new_new_n565_));
  NA2        g543(.A(i_4_), .B(i_8_), .Y(new_new_n566_));
  AOI210     g544(.A0(new_new_n566_), .A1(new_new_n294_), .B0(new_new_n565_), .Y(new_new_n567_));
  OAI220     g545(.A0(new_new_n567_), .A1(new_new_n563_), .B0(new_new_n564_), .B1(i_13_), .Y(new_new_n568_));
  NO3        g546(.A(new_new_n568_), .B(new_new_n562_), .C(new_new_n556_), .Y(new_new_n569_));
  AOI210     g547(.A0(new_new_n124_), .A1(new_new_n59_), .B0(i_10_), .Y(new_new_n570_));
  AOI210     g548(.A0(new_new_n570_), .A1(new_new_n230_), .B0(new_new_n155_), .Y(new_new_n571_));
  OR2        g549(.A(i_6_), .B(i_10_), .Y(new_new_n572_));
  NO2        g550(.A(new_new_n572_), .B(new_new_n23_), .Y(new_new_n573_));
  OR3        g551(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n574_));
  NO3        g552(.A(new_new_n574_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n575_));
  INV        g553(.A(new_new_n192_), .Y(new_new_n576_));
  NO2        g554(.A(new_new_n575_), .B(new_new_n573_), .Y(new_new_n577_));
  OA220      g555(.A0(new_new_n577_), .A1(new_new_n545_), .B0(new_new_n571_), .B1(new_new_n261_), .Y(new_new_n578_));
  AOI210     g556(.A0(new_new_n578_), .A1(new_new_n569_), .B0(new_new_n60_), .Y(new_new_n579_));
  NOi21      g557(.An(i_11_), .B(i_7_), .Y(new_new_n580_));
  AO210      g558(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n581_), .B(new_new_n580_), .Y(new_new_n582_));
  NA3        g560(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n583_));
  NO3        g561(.A(new_new_n250_), .B(new_new_n199_), .C(new_new_n558_), .Y(new_new_n584_));
  OAI210     g562(.A0(new_new_n584_), .A1(new_new_n219_), .B0(new_new_n60_), .Y(new_new_n585_));
  NO2        g563(.A(new_new_n60_), .B(i_9_), .Y(new_new_n586_));
  NO2        g564(.A(i_1_), .B(i_12_), .Y(new_new_n587_));
  INV        g565(.A(new_new_n585_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n588_), .B(i_6_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n583_), .B(new_new_n105_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n590_), .B(new_new_n546_), .Y(new_new_n591_));
  NO2        g569(.A(i_6_), .B(i_11_), .Y(new_new_n592_));
  INV        g570(.A(new_new_n591_), .Y(new_new_n593_));
  NO4        g571(.A(new_new_n207_), .B(new_new_n124_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n594_));
  NA2        g572(.A(new_new_n594_), .B(new_new_n586_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n230_), .B(i_6_), .Y(new_new_n596_));
  NO3        g574(.A(new_new_n572_), .B(new_new_n226_), .C(new_new_n23_), .Y(new_new_n597_));
  AOI210     g575(.A0(i_1_), .A1(new_new_n251_), .B0(new_new_n597_), .Y(new_new_n598_));
  OAI210     g576(.A0(new_new_n598_), .A1(new_new_n44_), .B0(new_new_n595_), .Y(new_new_n599_));
  NA3        g577(.A(new_new_n502_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n133_), .B(i_9_), .Y(new_new_n601_));
  NA3        g579(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n46_), .B(i_1_), .Y(new_new_n603_));
  NA3        g581(.A(new_new_n603_), .B(new_new_n260_), .C(new_new_n44_), .Y(new_new_n604_));
  OAI220     g582(.A0(new_new_n604_), .A1(new_new_n602_), .B0(new_new_n601_), .B1(new_new_n956_), .Y(new_new_n605_));
  NA3        g583(.A(new_new_n586_), .B(new_new_n304_), .C(i_6_), .Y(new_new_n606_));
  NO2        g584(.A(new_new_n606_), .B(new_new_n23_), .Y(new_new_n607_));
  NAi21      g585(.An(new_new_n600_), .B(new_new_n88_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n603_), .B(new_new_n260_), .Y(new_new_n609_));
  NO2        g587(.A(i_11_), .B(new_new_n37_), .Y(new_new_n610_));
  NA2        g588(.A(new_new_n610_), .B(new_new_n24_), .Y(new_new_n611_));
  OAI210     g589(.A0(new_new_n611_), .A1(new_new_n609_), .B0(new_new_n608_), .Y(new_new_n612_));
  OR3        g590(.A(new_new_n612_), .B(new_new_n607_), .C(new_new_n605_), .Y(new_new_n613_));
  NO3        g591(.A(new_new_n613_), .B(new_new_n599_), .C(new_new_n593_), .Y(new_new_n614_));
  NO2        g592(.A(new_new_n230_), .B(new_new_n98_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n615_), .B(new_new_n580_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n616_), .B(i_1_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n617_), .B(new_new_n574_), .Y(new_new_n618_));
  NO2        g596(.A(new_new_n395_), .B(new_new_n82_), .Y(new_new_n619_));
  NA2        g597(.A(new_new_n618_), .B(new_new_n46_), .Y(new_new_n620_));
  NO2        g598(.A(i_8_), .B(new_new_n112_), .Y(new_new_n621_));
  AN2        g599(.A(new_new_n621_), .B(new_new_n508_), .Y(new_new_n622_));
  NO2        g600(.A(new_new_n226_), .B(new_new_n44_), .Y(new_new_n623_));
  NO3        g601(.A(new_new_n623_), .B(new_new_n297_), .C(new_new_n231_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n113_), .B(new_new_n37_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(i_6_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n82_), .B(i_9_), .Y(new_new_n627_));
  NO2        g605(.A(new_new_n627_), .B(new_new_n60_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n628_), .B(new_new_n587_), .Y(new_new_n629_));
  NO4        g607(.A(new_new_n629_), .B(new_new_n626_), .C(new_new_n624_), .D(i_4_), .Y(new_new_n630_));
  NA2        g608(.A(i_1_), .B(i_3_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n432_), .B(new_new_n89_), .Y(new_new_n632_));
  AOI210     g610(.A0(new_new_n623_), .A1(new_new_n538_), .B0(new_new_n632_), .Y(new_new_n633_));
  NO2        g611(.A(new_new_n633_), .B(new_new_n631_), .Y(new_new_n634_));
  NO3        g612(.A(new_new_n634_), .B(new_new_n630_), .C(new_new_n622_), .Y(new_new_n635_));
  NA4        g613(.A(new_new_n635_), .B(new_new_n620_), .C(new_new_n614_), .D(new_new_n589_), .Y(new_new_n636_));
  NO3        g614(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n637_));
  NOi21      g615(.An(new_new_n637_), .B(i_10_), .Y(new_new_n638_));
  OA210      g616(.A0(new_new_n638_), .A1(new_new_n239_), .B0(new_new_n82_), .Y(new_new_n639_));
  NA2        g617(.A(new_new_n351_), .B(new_new_n350_), .Y(new_new_n640_));
  NA3        g618(.A(new_new_n452_), .B(new_new_n487_), .C(new_new_n46_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n641_), .B(new_new_n640_), .Y(new_new_n642_));
  OAI210     g620(.A0(new_new_n642_), .A1(new_new_n639_), .B0(i_1_), .Y(new_new_n643_));
  AOI210     g621(.A0(new_new_n260_), .A1(new_new_n94_), .B0(i_1_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n349_), .B(i_2_), .Y(new_new_n645_));
  NA2        g623(.A(new_new_n645_), .B(new_new_n644_), .Y(new_new_n646_));
  OAI210     g624(.A0(new_new_n606_), .A1(new_new_n428_), .B0(new_new_n646_), .Y(new_new_n647_));
  INV        g625(.A(new_new_n647_), .Y(new_new_n648_));
  AOI210     g626(.A0(new_new_n648_), .A1(new_new_n643_), .B0(i_13_), .Y(new_new_n649_));
  OR2        g627(.A(i_11_), .B(i_7_), .Y(new_new_n650_));
  NO2        g628(.A(new_new_n52_), .B(i_12_), .Y(new_new_n651_));
  AOI220     g629(.A0(i_7_), .A1(new_new_n619_), .B0(new_new_n239_), .B1(new_new_n127_), .Y(new_new_n652_));
  OAI220     g630(.A0(new_new_n652_), .A1(new_new_n41_), .B0(new_new_n955_), .B1(new_new_n89_), .Y(new_new_n653_));
  INV        g631(.A(new_new_n653_), .Y(new_new_n654_));
  AOI210     g632(.A0(new_new_n428_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n655_));
  NOi31      g633(.An(new_new_n655_), .B(new_new_n557_), .C(new_new_n44_), .Y(new_new_n656_));
  NA2        g634(.A(new_new_n123_), .B(i_13_), .Y(new_new_n657_));
  NO2        g635(.A(new_new_n602_), .B(new_new_n112_), .Y(new_new_n658_));
  INV        g636(.A(new_new_n658_), .Y(new_new_n659_));
  OAI220     g637(.A0(new_new_n659_), .A1(new_new_n68_), .B0(new_new_n657_), .B1(new_new_n644_), .Y(new_new_n660_));
  NA2        g638(.A(new_new_n26_), .B(new_new_n186_), .Y(new_new_n661_));
  NA2        g639(.A(new_new_n661_), .B(i_7_), .Y(new_new_n662_));
  NO3        g640(.A(new_new_n447_), .B(new_new_n230_), .C(new_new_n82_), .Y(new_new_n663_));
  NA2        g641(.A(new_new_n663_), .B(new_new_n662_), .Y(new_new_n664_));
  AOI220     g642(.A0(new_new_n366_), .A1(new_new_n603_), .B0(new_new_n88_), .B1(new_new_n99_), .Y(new_new_n665_));
  OAI220     g643(.A0(new_new_n665_), .A1(new_new_n561_), .B0(new_new_n664_), .B1(new_new_n576_), .Y(new_new_n666_));
  NO3        g644(.A(new_new_n666_), .B(new_new_n660_), .C(new_new_n656_), .Y(new_new_n667_));
  OR2        g645(.A(i_11_), .B(i_6_), .Y(new_new_n668_));
  NA3        g646(.A(new_new_n560_), .B(new_new_n661_), .C(i_7_), .Y(new_new_n669_));
  AOI210     g647(.A0(new_new_n669_), .A1(new_new_n659_), .B0(new_new_n668_), .Y(new_new_n670_));
  NA3        g648(.A(new_new_n389_), .B(new_new_n565_), .C(new_new_n94_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n592_), .B(i_13_), .Y(new_new_n672_));
  NAi21      g650(.An(i_11_), .B(i_12_), .Y(new_new_n673_));
  NOi41      g651(.An(new_new_n108_), .B(new_new_n673_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n674_));
  INV        g652(.A(new_new_n674_), .Y(new_new_n675_));
  NA3        g653(.A(new_new_n675_), .B(new_new_n672_), .C(new_new_n671_), .Y(new_new_n676_));
  OAI210     g654(.A0(new_new_n676_), .A1(new_new_n670_), .B0(new_new_n60_), .Y(new_new_n677_));
  NO2        g655(.A(i_2_), .B(i_12_), .Y(new_new_n678_));
  NA2        g656(.A(new_new_n348_), .B(new_new_n678_), .Y(new_new_n679_));
  NO3        g657(.A(i_9_), .B(new_new_n364_), .C(new_new_n560_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n680_), .B(new_new_n348_), .Y(new_new_n681_));
  NO2        g659(.A(new_new_n124_), .B(i_2_), .Y(new_new_n682_));
  NA2        g660(.A(new_new_n682_), .B(new_new_n587_), .Y(new_new_n683_));
  NA3        g661(.A(new_new_n683_), .B(new_new_n681_), .C(new_new_n679_), .Y(new_new_n684_));
  NA3        g662(.A(new_new_n684_), .B(new_new_n45_), .C(new_new_n218_), .Y(new_new_n685_));
  NA4        g663(.A(new_new_n685_), .B(new_new_n677_), .C(new_new_n667_), .D(new_new_n654_), .Y(new_new_n686_));
  OR4        g664(.A(new_new_n686_), .B(new_new_n649_), .C(new_new_n636_), .D(new_new_n579_), .Y(mai5));
  NA2        g665(.A(new_new_n616_), .B(new_new_n262_), .Y(new_new_n688_));
  AN2        g666(.A(new_new_n24_), .B(i_10_), .Y(new_new_n689_));
  NA3        g667(.A(new_new_n689_), .B(new_new_n678_), .C(new_new_n105_), .Y(new_new_n690_));
  NO2        g668(.A(new_new_n561_), .B(i_11_), .Y(new_new_n691_));
  NA2        g669(.A(new_new_n83_), .B(new_new_n691_), .Y(new_new_n692_));
  NA3        g670(.A(new_new_n692_), .B(new_new_n690_), .C(new_new_n688_), .Y(new_new_n693_));
  NO3        g671(.A(i_11_), .B(new_new_n230_), .C(i_13_), .Y(new_new_n694_));
  NO2        g672(.A(new_new_n120_), .B(new_new_n23_), .Y(new_new_n695_));
  NA2        g673(.A(i_12_), .B(i_8_), .Y(new_new_n696_));
  INV        g674(.A(new_new_n427_), .Y(new_new_n697_));
  AOI220     g675(.A0(new_new_n304_), .A1(new_new_n539_), .B0(i_12_), .B1(new_new_n695_), .Y(new_new_n698_));
  INV        g676(.A(new_new_n698_), .Y(new_new_n699_));
  NO2        g677(.A(new_new_n699_), .B(new_new_n693_), .Y(new_new_n700_));
  INV        g678(.A(new_new_n165_), .Y(new_new_n701_));
  INV        g679(.A(new_new_n239_), .Y(new_new_n702_));
  OAI210     g680(.A0(new_new_n645_), .A1(new_new_n429_), .B0(new_new_n108_), .Y(new_new_n703_));
  AOI210     g681(.A0(new_new_n703_), .A1(new_new_n702_), .B0(new_new_n701_), .Y(new_new_n704_));
  INV        g682(.A(new_new_n399_), .Y(new_new_n705_));
  NA2        g683(.A(new_new_n705_), .B(i_2_), .Y(new_new_n706_));
  INV        g684(.A(new_new_n706_), .Y(new_new_n707_));
  AOI210     g685(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n396_), .Y(new_new_n708_));
  AOI210     g686(.A0(new_new_n708_), .A1(new_new_n707_), .B0(new_new_n704_), .Y(new_new_n709_));
  NO2        g687(.A(new_new_n183_), .B(new_new_n121_), .Y(new_new_n710_));
  OAI210     g688(.A0(new_new_n710_), .A1(new_new_n695_), .B0(i_2_), .Y(new_new_n711_));
  INV        g689(.A(new_new_n166_), .Y(new_new_n712_));
  NO3        g690(.A(new_new_n581_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n713_));
  AOI210     g691(.A0(new_new_n712_), .A1(new_new_n83_), .B0(new_new_n713_), .Y(new_new_n714_));
  AOI210     g692(.A0(new_new_n714_), .A1(new_new_n711_), .B0(new_new_n186_), .Y(new_new_n715_));
  OA210      g693(.A0(new_new_n582_), .A1(new_new_n122_), .B0(i_13_), .Y(new_new_n716_));
  INV        g694(.A(new_new_n146_), .Y(new_new_n717_));
  NO2        g695(.A(new_new_n717_), .B(new_new_n353_), .Y(new_new_n718_));
  AOI210     g696(.A0(new_new_n199_), .A1(new_new_n143_), .B0(new_new_n487_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n719_), .B(new_new_n399_), .Y(new_new_n720_));
  NO2        g698(.A(new_new_n99_), .B(new_new_n44_), .Y(new_new_n721_));
  INV        g699(.A(new_new_n290_), .Y(new_new_n722_));
  NA4        g700(.A(new_new_n722_), .B(new_new_n294_), .C(new_new_n120_), .D(new_new_n42_), .Y(new_new_n723_));
  OAI210     g701(.A0(new_new_n723_), .A1(new_new_n721_), .B0(new_new_n720_), .Y(new_new_n724_));
  NO4        g702(.A(new_new_n724_), .B(new_new_n718_), .C(new_new_n716_), .D(new_new_n715_), .Y(new_new_n725_));
  NO2        g703(.A(new_new_n59_), .B(i_12_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n726_), .B(new_new_n122_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n727_), .B(new_new_n558_), .Y(new_new_n728_));
  NA2        g706(.A(new_new_n728_), .B(new_new_n36_), .Y(new_new_n729_));
  NA4        g707(.A(new_new_n729_), .B(new_new_n725_), .C(new_new_n709_), .D(new_new_n700_), .Y(mai6));
  NO3        g708(.A(i_9_), .B(new_new_n296_), .C(i_1_), .Y(new_new_n731_));
  NO2        g709(.A(new_new_n178_), .B(new_new_n134_), .Y(new_new_n732_));
  OAI210     g710(.A0(new_new_n732_), .A1(new_new_n731_), .B0(new_new_n682_), .Y(new_new_n733_));
  NO2        g711(.A(new_new_n213_), .B(new_new_n456_), .Y(new_new_n734_));
  INV        g712(.A(new_new_n316_), .Y(new_new_n735_));
  AO210      g713(.A0(new_new_n735_), .A1(new_new_n733_), .B0(i_12_), .Y(new_new_n736_));
  NA2        g714(.A(new_new_n354_), .B(new_new_n321_), .Y(new_new_n737_));
  NA2        g715(.A(new_new_n546_), .B(new_new_n60_), .Y(new_new_n738_));
  NA2        g716(.A(new_new_n638_), .B(new_new_n68_), .Y(new_new_n739_));
  NA3        g717(.A(new_new_n739_), .B(new_new_n738_), .C(new_new_n737_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n740_), .B(new_new_n70_), .Y(new_new_n741_));
  INV        g719(.A(new_new_n315_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n72_), .B(new_new_n127_), .Y(new_new_n743_));
  INV        g721(.A(new_new_n120_), .Y(new_new_n744_));
  NA2        g722(.A(new_new_n744_), .B(new_new_n46_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n745_), .A1(new_new_n743_), .B0(new_new_n742_), .Y(new_new_n746_));
  NO2        g724(.A(new_new_n32_), .B(i_11_), .Y(new_new_n747_));
  NA3        g725(.A(new_new_n747_), .B(new_new_n444_), .C(new_new_n370_), .Y(new_new_n748_));
  OAI210     g726(.A0(new_new_n637_), .A1(new_new_n530_), .B0(new_new_n529_), .Y(new_new_n749_));
  NA2        g727(.A(new_new_n749_), .B(new_new_n748_), .Y(new_new_n750_));
  OR2        g728(.A(new_new_n750_), .B(new_new_n746_), .Y(new_new_n751_));
  NO2        g729(.A(new_new_n650_), .B(i_2_), .Y(new_new_n752_));
  NA2        g730(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n753_));
  NO2        g731(.A(new_new_n753_), .B(new_new_n388_), .Y(new_new_n754_));
  NA2        g732(.A(new_new_n754_), .B(new_new_n752_), .Y(new_new_n755_));
  AO210      g733(.A0(new_new_n342_), .A1(new_new_n334_), .B0(new_new_n376_), .Y(new_new_n756_));
  NA3        g734(.A(new_new_n756_), .B(new_new_n247_), .C(i_7_), .Y(new_new_n757_));
  OR2        g735(.A(new_new_n582_), .B(new_new_n429_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n758_), .B(new_new_n142_), .Y(new_new_n759_));
  AO210      g737(.A0(new_new_n462_), .A1(new_new_n697_), .B0(new_new_n36_), .Y(new_new_n760_));
  NA4        g738(.A(new_new_n760_), .B(new_new_n759_), .C(new_new_n757_), .D(new_new_n755_), .Y(new_new_n761_));
  NO2        g739(.A(i_6_), .B(i_11_), .Y(new_new_n762_));
  AOI220     g740(.A0(new_new_n762_), .A1(new_new_n529_), .B0(new_new_n734_), .B1(new_new_n662_), .Y(new_new_n763_));
  NA3        g741(.A(new_new_n353_), .B(new_new_n232_), .C(new_new_n142_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n376_), .B(new_new_n67_), .Y(new_new_n765_));
  NA4        g743(.A(new_new_n765_), .B(new_new_n764_), .C(new_new_n763_), .D(new_new_n564_), .Y(new_new_n766_));
  AOI210     g744(.A0(new_new_n429_), .A1(new_new_n427_), .B0(new_new_n528_), .Y(new_new_n767_));
  NO2        g745(.A(new_new_n572_), .B(new_new_n99_), .Y(new_new_n768_));
  OAI210     g746(.A0(new_new_n768_), .A1(new_new_n109_), .B0(new_new_n386_), .Y(new_new_n769_));
  INV        g747(.A(new_new_n549_), .Y(new_new_n770_));
  NA3        g748(.A(new_new_n770_), .B(new_new_n315_), .C(i_7_), .Y(new_new_n771_));
  NA3        g749(.A(new_new_n771_), .B(new_new_n769_), .C(new_new_n767_), .Y(new_new_n772_));
  NO4        g750(.A(new_new_n772_), .B(new_new_n766_), .C(new_new_n761_), .D(new_new_n751_), .Y(new_new_n773_));
  NA4        g751(.A(new_new_n773_), .B(new_new_n741_), .C(new_new_n736_), .D(new_new_n360_), .Y(mai3));
  NA2        g752(.A(i_6_), .B(i_7_), .Y(new_new_n775_));
  NO2        g753(.A(new_new_n775_), .B(i_0_), .Y(new_new_n776_));
  NO2        g754(.A(i_11_), .B(new_new_n230_), .Y(new_new_n777_));
  NA2        g755(.A(new_new_n278_), .B(new_new_n777_), .Y(new_new_n778_));
  NO2        g756(.A(new_new_n778_), .B(new_new_n186_), .Y(new_new_n779_));
  NO3        g757(.A(new_new_n430_), .B(new_new_n86_), .C(new_new_n44_), .Y(new_new_n780_));
  OA210      g758(.A0(new_new_n780_), .A1(new_new_n779_), .B0(new_new_n168_), .Y(new_new_n781_));
  NA2        g759(.A(new_new_n764_), .B(new_new_n352_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n782_), .B(new_new_n40_), .Y(new_new_n783_));
  AN2        g761(.A(new_new_n431_), .B(new_new_n53_), .Y(new_new_n784_));
  AOI210     g762(.A0(new_new_n957_), .A1(new_new_n783_), .B0(new_new_n48_), .Y(new_new_n785_));
  NO4        g763(.A(new_new_n357_), .B(new_new_n363_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n786_));
  INV        g764(.A(new_new_n786_), .Y(new_new_n787_));
  NA2        g765(.A(new_new_n655_), .B(new_new_n627_), .Y(new_new_n788_));
  NA2        g766(.A(new_new_n319_), .B(i_5_), .Y(new_new_n789_));
  OAI220     g767(.A0(new_new_n789_), .A1(new_new_n788_), .B0(new_new_n787_), .B1(new_new_n60_), .Y(new_new_n790_));
  NOi21      g768(.An(i_5_), .B(i_9_), .Y(new_new_n791_));
  NA2        g769(.A(new_new_n791_), .B(new_new_n426_), .Y(new_new_n792_));
  NO3        g770(.A(new_new_n392_), .B(new_new_n260_), .C(new_new_n70_), .Y(new_new_n793_));
  NO2        g771(.A(new_new_n169_), .B(new_new_n143_), .Y(new_new_n794_));
  AOI210     g772(.A0(new_new_n794_), .A1(new_new_n238_), .B0(new_new_n793_), .Y(new_new_n795_));
  NO2        g773(.A(new_new_n795_), .B(new_new_n959_), .Y(new_new_n796_));
  NO4        g774(.A(new_new_n796_), .B(new_new_n790_), .C(new_new_n785_), .D(new_new_n781_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n178_), .B(new_new_n24_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n301_), .B(new_new_n125_), .Y(new_new_n799_));
  NAi21      g777(.An(new_new_n156_), .B(i_5_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n799_), .B(new_new_n378_), .Y(new_new_n801_));
  INV        g779(.A(new_new_n801_), .Y(new_new_n802_));
  NO2        g780(.A(new_new_n370_), .B(new_new_n282_), .Y(new_new_n803_));
  NA2        g781(.A(new_new_n803_), .B(new_new_n658_), .Y(new_new_n804_));
  NO4        g782(.A(new_new_n548_), .B(new_new_n207_), .C(new_new_n396_), .D(new_new_n388_), .Y(new_new_n805_));
  AN2        g783(.A(new_new_n93_), .B(new_new_n237_), .Y(new_new_n806_));
  NA2        g784(.A(new_new_n694_), .B(new_new_n316_), .Y(new_new_n807_));
  AOI210     g785(.A0(new_new_n452_), .A1(new_new_n83_), .B0(new_new_n55_), .Y(new_new_n808_));
  OAI220     g786(.A0(new_new_n808_), .A1(new_new_n807_), .B0(new_new_n611_), .B1(new_new_n504_), .Y(new_new_n809_));
  NO2        g787(.A(new_new_n245_), .B(new_new_n147_), .Y(new_new_n810_));
  NA2        g788(.A(i_0_), .B(i_10_), .Y(new_new_n811_));
  AN2        g789(.A(new_new_n810_), .B(i_6_), .Y(new_new_n812_));
  AOI220     g790(.A0(new_new_n319_), .A1(new_new_n95_), .B0(new_new_n178_), .B1(new_new_n80_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n533_), .B(i_4_), .Y(new_new_n814_));
  NA2        g792(.A(new_new_n181_), .B(new_new_n195_), .Y(new_new_n815_));
  OAI220     g793(.A0(new_new_n815_), .A1(new_new_n807_), .B0(new_new_n814_), .B1(new_new_n813_), .Y(new_new_n816_));
  NO4        g794(.A(new_new_n816_), .B(new_new_n812_), .C(new_new_n809_), .D(new_new_n806_), .Y(new_new_n817_));
  NA3        g795(.A(new_new_n817_), .B(new_new_n804_), .C(new_new_n802_), .Y(new_new_n818_));
  NO2        g796(.A(new_new_n48_), .B(i_7_), .Y(new_new_n819_));
  NA2        g797(.A(new_new_n374_), .B(new_new_n173_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n820_), .B(new_new_n154_), .Y(new_new_n821_));
  NO2        g799(.A(new_new_n169_), .B(i_0_), .Y(new_new_n822_));
  INV        g800(.A(new_new_n822_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n444_), .B(new_new_n224_), .Y(new_new_n824_));
  INV        g802(.A(new_new_n385_), .Y(new_new_n825_));
  OAI220     g803(.A0(new_new_n825_), .A1(new_new_n792_), .B0(new_new_n824_), .B1(new_new_n823_), .Y(new_new_n826_));
  NO2        g804(.A(new_new_n826_), .B(new_new_n821_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n610_), .B(new_new_n117_), .Y(new_new_n828_));
  NO2        g806(.A(i_6_), .B(new_new_n828_), .Y(new_new_n829_));
  AOI210     g807(.A0(new_new_n428_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n165_), .B(new_new_n100_), .Y(new_new_n831_));
  NOi32      g809(.An(new_new_n830_), .Bn(new_new_n181_), .C(new_new_n831_), .Y(new_new_n832_));
  NO2        g810(.A(new_new_n832_), .B(new_new_n829_), .Y(new_new_n833_));
  NOi21      g811(.An(i_7_), .B(i_5_), .Y(new_new_n834_));
  NOi31      g812(.An(new_new_n834_), .B(i_0_), .C(new_new_n673_), .Y(new_new_n835_));
  NA3        g813(.A(new_new_n835_), .B(new_new_n364_), .C(i_6_), .Y(new_new_n836_));
  OA210      g814(.A0(new_new_n831_), .A1(new_new_n485_), .B0(new_new_n836_), .Y(new_new_n837_));
  NO3        g815(.A(new_new_n381_), .B(new_new_n345_), .C(new_new_n341_), .Y(new_new_n838_));
  NO2        g816(.A(new_new_n254_), .B(new_new_n305_), .Y(new_new_n839_));
  NO2        g817(.A(new_new_n673_), .B(new_new_n249_), .Y(new_new_n840_));
  AOI210     g818(.A0(new_new_n840_), .A1(new_new_n839_), .B0(new_new_n838_), .Y(new_new_n841_));
  NA4        g819(.A(new_new_n841_), .B(new_new_n837_), .C(new_new_n833_), .D(new_new_n827_), .Y(new_new_n842_));
  NO2        g820(.A(new_new_n798_), .B(new_new_n233_), .Y(new_new_n843_));
  AN2        g821(.A(new_new_n318_), .B(new_new_n316_), .Y(new_new_n844_));
  NA2        g822(.A(new_new_n843_), .B(i_10_), .Y(new_new_n845_));
  OA210      g823(.A0(new_new_n444_), .A1(new_new_n216_), .B0(new_new_n443_), .Y(new_new_n846_));
  NA3        g824(.A(new_new_n443_), .B(new_new_n389_), .C(new_new_n45_), .Y(new_new_n847_));
  OAI210     g825(.A0(new_new_n800_), .A1(i_6_), .B0(new_new_n847_), .Y(new_new_n848_));
  INV        g826(.A(new_new_n180_), .Y(new_new_n849_));
  AOI220     g827(.A0(new_new_n849_), .A1(new_new_n444_), .B0(new_new_n848_), .B1(new_new_n70_), .Y(new_new_n850_));
  NA2        g828(.A(new_new_n89_), .B(new_new_n44_), .Y(new_new_n851_));
  NO2        g829(.A(new_new_n72_), .B(new_new_n696_), .Y(new_new_n852_));
  NA2        g830(.A(new_new_n852_), .B(new_new_n851_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n853_), .B(new_new_n47_), .Y(new_new_n854_));
  NO2        g832(.A(new_new_n559_), .B(new_new_n102_), .Y(new_new_n855_));
  NA2        g833(.A(new_new_n855_), .B(i_0_), .Y(new_new_n856_));
  NO2        g834(.A(new_new_n856_), .B(new_new_n82_), .Y(new_new_n857_));
  NO3        g835(.A(new_new_n857_), .B(new_new_n854_), .C(new_new_n489_), .Y(new_new_n858_));
  NA3        g836(.A(new_new_n858_), .B(new_new_n850_), .C(new_new_n845_), .Y(new_new_n859_));
  NO3        g837(.A(new_new_n859_), .B(new_new_n842_), .C(new_new_n818_), .Y(new_new_n860_));
  NO2        g838(.A(i_0_), .B(new_new_n673_), .Y(new_new_n861_));
  NA2        g839(.A(new_new_n70_), .B(new_new_n44_), .Y(new_new_n862_));
  INV        g840(.A(new_new_n862_), .Y(new_new_n863_));
  NO3        g841(.A(new_new_n102_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n864_));
  AO220      g842(.A0(new_new_n864_), .A1(new_new_n863_), .B0(new_new_n861_), .B1(new_new_n168_), .Y(new_new_n865_));
  AOI210     g843(.A0(new_new_n738_), .A1(new_new_n640_), .B0(new_new_n831_), .Y(new_new_n866_));
  AOI210     g844(.A0(new_new_n865_), .A1(new_new_n331_), .B0(new_new_n866_), .Y(new_new_n867_));
  NA3        g845(.A(new_new_n141_), .B(new_new_n627_), .C(new_new_n70_), .Y(new_new_n868_));
  NO2        g846(.A(new_new_n749_), .B(new_new_n381_), .Y(new_new_n869_));
  NA3        g847(.A(new_new_n776_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n870_));
  NA2        g848(.A(new_new_n777_), .B(i_9_), .Y(new_new_n871_));
  AOI210     g849(.A0(new_new_n870_), .A1(new_new_n467_), .B0(new_new_n871_), .Y(new_new_n872_));
  NA2        g850(.A(new_new_n238_), .B(new_new_n223_), .Y(new_new_n873_));
  NO2        g851(.A(new_new_n873_), .B(new_new_n147_), .Y(new_new_n874_));
  NO3        g852(.A(new_new_n874_), .B(new_new_n872_), .C(new_new_n869_), .Y(new_new_n875_));
  NA3        g853(.A(new_new_n875_), .B(new_new_n868_), .C(new_new_n867_), .Y(new_new_n876_));
  NA2        g854(.A(new_new_n844_), .B(new_new_n353_), .Y(new_new_n877_));
  AOI210     g855(.A0(new_new_n289_), .A1(new_new_n156_), .B0(new_new_n877_), .Y(new_new_n878_));
  NA2        g856(.A(new_new_n40_), .B(new_new_n44_), .Y(new_new_n879_));
  NA2        g857(.A(new_new_n819_), .B(new_new_n457_), .Y(new_new_n880_));
  AOI210     g858(.A0(new_new_n879_), .A1(new_new_n156_), .B0(new_new_n880_), .Y(new_new_n881_));
  NO2        g859(.A(new_new_n881_), .B(new_new_n878_), .Y(new_new_n882_));
  NO3        g860(.A(new_new_n811_), .B(new_new_n791_), .C(new_new_n183_), .Y(new_new_n883_));
  AOI220     g861(.A0(new_new_n883_), .A1(i_11_), .B0(new_new_n534_), .B1(new_new_n72_), .Y(new_new_n884_));
  NO3        g862(.A(new_new_n201_), .B(new_new_n363_), .C(i_0_), .Y(new_new_n885_));
  OAI210     g863(.A0(new_new_n885_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n886_));
  INV        g864(.A(new_new_n210_), .Y(new_new_n887_));
  OAI220     g865(.A0(new_new_n497_), .A1(new_new_n134_), .B0(new_new_n596_), .B1(new_new_n576_), .Y(new_new_n888_));
  NA3        g866(.A(new_new_n888_), .B(i_7_), .C(new_new_n887_), .Y(new_new_n889_));
  NA4        g867(.A(new_new_n889_), .B(new_new_n886_), .C(new_new_n884_), .D(new_new_n882_), .Y(new_new_n890_));
  INV        g868(.A(new_new_n106_), .Y(new_new_n891_));
  NA2        g869(.A(new_new_n834_), .B(new_new_n457_), .Y(new_new_n892_));
  INV        g870(.A(new_new_n170_), .Y(new_new_n893_));
  OA220      g871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n891_), .B1(i_5_), .Y(new_new_n894_));
  AOI210     g872(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n169_), .Y(new_new_n895_));
  NA2        g873(.A(new_new_n895_), .B(new_new_n846_), .Y(new_new_n896_));
  NA3        g874(.A(new_new_n370_), .B(new_new_n320_), .C(new_new_n214_), .Y(new_new_n897_));
  INV        g875(.A(new_new_n897_), .Y(new_new_n898_));
  NOi31      g876(.An(new_new_n369_), .B(new_new_n862_), .C(new_new_n233_), .Y(new_new_n899_));
  NO2        g877(.A(new_new_n899_), .B(new_new_n898_), .Y(new_new_n900_));
  NA4        g878(.A(new_new_n900_), .B(new_new_n441_), .C(new_new_n896_), .D(new_new_n894_), .Y(new_new_n901_));
  NA3        g879(.A(new_new_n294_), .B(i_5_), .C(new_new_n186_), .Y(new_new_n902_));
  NAi31      g880(.An(new_new_n235_), .B(new_new_n902_), .C(new_new_n236_), .Y(new_new_n903_));
  NO4        g881(.A(new_new_n233_), .B(new_new_n201_), .C(i_0_), .D(i_12_), .Y(new_new_n904_));
  NA2        g882(.A(new_new_n904_), .B(new_new_n903_), .Y(new_new_n905_));
  AN2        g883(.A(new_new_n811_), .B(new_new_n147_), .Y(new_new_n906_));
  NO4        g884(.A(new_new_n906_), .B(i_12_), .C(new_new_n600_), .D(new_new_n127_), .Y(new_new_n907_));
  NA2        g885(.A(new_new_n907_), .B(new_new_n210_), .Y(new_new_n908_));
  NA3        g886(.A(new_new_n95_), .B(new_new_n538_), .C(i_11_), .Y(new_new_n909_));
  NA2        g887(.A(new_new_n834_), .B(new_new_n440_), .Y(new_new_n910_));
  NA2        g888(.A(new_new_n61_), .B(new_new_n98_), .Y(new_new_n911_));
  OAI220     g889(.A0(new_new_n911_), .A1(new_new_n902_), .B0(new_new_n910_), .B1(new_new_n628_), .Y(new_new_n912_));
  NA2        g890(.A(new_new_n912_), .B(new_new_n822_), .Y(new_new_n913_));
  NA3        g891(.A(new_new_n913_), .B(new_new_n908_), .C(new_new_n905_), .Y(new_new_n914_));
  NO4        g892(.A(new_new_n914_), .B(new_new_n901_), .C(new_new_n890_), .D(new_new_n876_), .Y(new_new_n915_));
  OAI210     g893(.A0(new_new_n752_), .A1(new_new_n747_), .B0(new_new_n37_), .Y(new_new_n916_));
  NA3        g894(.A(new_new_n830_), .B(new_new_n348_), .C(i_5_), .Y(new_new_n917_));
  NA3        g895(.A(new_new_n917_), .B(new_new_n916_), .C(new_new_n571_), .Y(new_new_n918_));
  NA2        g896(.A(new_new_n918_), .B(new_new_n197_), .Y(new_new_n919_));
  BUFFER     g897(.A(new_new_n349_), .Y(new_new_n920_));
  NA2        g898(.A(new_new_n179_), .B(new_new_n181_), .Y(new_new_n921_));
  AO210      g899(.A0(new_new_n920_), .A1(new_new_n33_), .B0(new_new_n921_), .Y(new_new_n922_));
  OAI210     g900(.A0(new_new_n575_), .A1(new_new_n573_), .B0(new_new_n304_), .Y(new_new_n923_));
  NAi31      g901(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n924_));
  NO2        g902(.A(new_new_n67_), .B(new_new_n924_), .Y(new_new_n925_));
  NO2        g903(.A(new_new_n925_), .B(new_new_n597_), .Y(new_new_n926_));
  NA3        g904(.A(new_new_n926_), .B(new_new_n923_), .C(new_new_n922_), .Y(new_new_n927_));
  NO2        g905(.A(new_new_n434_), .B(new_new_n260_), .Y(new_new_n928_));
  NO4        g906(.A(new_new_n226_), .B(new_new_n140_), .C(new_new_n631_), .D(new_new_n37_), .Y(new_new_n929_));
  NO3        g907(.A(new_new_n929_), .B(new_new_n928_), .C(new_new_n805_), .Y(new_new_n930_));
  OAI210     g908(.A0(new_new_n909_), .A1(new_new_n143_), .B0(new_new_n930_), .Y(new_new_n931_));
  AOI210     g909(.A0(new_new_n927_), .A1(new_new_n48_), .B0(new_new_n931_), .Y(new_new_n932_));
  AOI210     g910(.A0(new_new_n932_), .A1(new_new_n919_), .B0(new_new_n70_), .Y(new_new_n933_));
  NO2        g911(.A(new_new_n531_), .B(new_new_n359_), .Y(new_new_n934_));
  NO2        g912(.A(new_new_n934_), .B(new_new_n701_), .Y(new_new_n935_));
  OAI210     g913(.A0(new_new_n77_), .A1(new_new_n52_), .B0(new_new_n105_), .Y(new_new_n936_));
  NA2        g914(.A(new_new_n936_), .B(new_new_n73_), .Y(new_new_n937_));
  AOI210     g915(.A0(new_new_n895_), .A1(new_new_n819_), .B0(new_new_n835_), .Y(new_new_n938_));
  AOI210     g916(.A0(new_new_n938_), .A1(new_new_n937_), .B0(new_new_n631_), .Y(new_new_n939_));
  NA2        g917(.A(new_new_n254_), .B(new_new_n54_), .Y(new_new_n940_));
  NA2        g918(.A(new_new_n940_), .B(new_new_n73_), .Y(new_new_n941_));
  NO2        g919(.A(new_new_n941_), .B(new_new_n230_), .Y(new_new_n942_));
  NA3        g920(.A(new_new_n93_), .B(new_new_n296_), .C(new_new_n31_), .Y(new_new_n943_));
  INV        g921(.A(new_new_n943_), .Y(new_new_n944_));
  NO3        g922(.A(new_new_n944_), .B(new_new_n942_), .C(new_new_n939_), .Y(new_new_n945_));
  OAI210     g923(.A0(new_new_n960_), .A1(new_new_n830_), .B0(new_new_n197_), .Y(new_new_n946_));
  NA2        g924(.A(new_new_n157_), .B(i_5_), .Y(new_new_n947_));
  NO2        g925(.A(new_new_n946_), .B(new_new_n947_), .Y(new_new_n948_));
  INV        g926(.A(new_new_n948_), .Y(new_new_n949_));
  OAI210     g927(.A0(new_new_n945_), .A1(i_4_), .B0(new_new_n949_), .Y(new_new_n950_));
  NO3        g928(.A(new_new_n950_), .B(new_new_n935_), .C(new_new_n933_), .Y(new_new_n951_));
  NA4        g929(.A(new_new_n951_), .B(new_new_n915_), .C(new_new_n860_), .D(new_new_n797_), .Y(mai4));
  INV        g930(.A(new_new_n651_), .Y(new_new_n955_));
  INV        g931(.A(i_2_), .Y(new_new_n956_));
  INV        g932(.A(new_new_n784_), .Y(new_new_n957_));
  INV        g933(.A(i_12_), .Y(new_new_n958_));
  INV        g934(.A(i_5_), .Y(new_new_n959_));
  INV        g935(.A(i_12_), .Y(new_new_n960_));
  INV        g936(.A(i_7_), .Y(new_new_n961_));
endmodule


