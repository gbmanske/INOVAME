//Benchmark atmr_9sym_175_0.0625

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n154_, mai_mai_n155_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n156_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  NA2        o002(.A(i_4_), .B(ori_ori_n12_), .Y(ori_ori_n13_));
  INV        o003(.A(i_5_), .Y(ori_ori_n14_));
  NOi21      o004(.An(i_3_), .B(i_7_), .Y(ori_ori_n15_));
  INV        o005(.A(ori_ori_n15_), .Y(ori_ori_n16_));
  INV        o006(.A(i_0_), .Y(ori_ori_n17_));
  NOi21      o007(.An(i_1_), .B(i_3_), .Y(ori_ori_n18_));
  NO2        o008(.A(ori_ori_n16_), .B(ori_ori_n13_), .Y(ori_ori_n19_));
  INV        o009(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o010(.A(i_0_), .B(ori_ori_n20_), .Y(ori_ori_n21_));
  INV        o011(.A(i_7_), .Y(ori_ori_n22_));
  NA3        o012(.A(i_6_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n23_));
  NOi21      o013(.An(i_8_), .B(i_6_), .Y(ori_ori_n24_));
  NOi21      o014(.An(i_1_), .B(i_8_), .Y(ori_ori_n25_));
  AOI220     o015(.A0(ori_ori_n25_), .A1(i_2_), .B0(ori_ori_n24_), .B1(i_5_), .Y(ori_ori_n26_));
  AOI210     o016(.A0(ori_ori_n26_), .A1(ori_ori_n23_), .B0(ori_ori_n21_), .Y(ori_ori_n27_));
  AOI210     o017(.A0(ori_ori_n27_), .A1(ori_ori_n11_), .B0(ori_ori_n19_), .Y(ori_ori_n28_));
  INV        o018(.A(i_0_), .Y(ori_ori_n29_));
  NA2        o019(.A(ori_ori_n17_), .B(i_5_), .Y(ori_ori_n30_));
  NO2        o020(.A(i_2_), .B(i_4_), .Y(ori_ori_n31_));
  NA3        o021(.A(ori_ori_n31_), .B(i_6_), .C(i_8_), .Y(ori_ori_n32_));
  AOI210     o022(.A0(ori_ori_n30_), .A1(ori_ori_n29_), .B0(ori_ori_n32_), .Y(ori_ori_n33_));
  INV        o023(.A(i_2_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_5_), .B(i_0_), .Y(ori_ori_n35_));
  NOi21      o025(.An(i_6_), .B(i_8_), .Y(ori_ori_n36_));
  NOi21      o026(.An(i_5_), .B(i_6_), .Y(ori_ori_n37_));
  NA2        o027(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n38_));
  NO3        o028(.A(ori_ori_n38_), .B(ori_ori_n34_), .C(i_4_), .Y(ori_ori_n39_));
  NOi21      o029(.An(i_0_), .B(i_4_), .Y(ori_ori_n40_));
  XO2        o030(.A(i_1_), .B(i_3_), .Y(ori_ori_n41_));
  INV        o031(.A(i_1_), .Y(ori_ori_n42_));
  NOi21      o032(.An(i_3_), .B(i_0_), .Y(ori_ori_n43_));
  NA2        o033(.A(ori_ori_n43_), .B(ori_ori_n42_), .Y(ori_ori_n44_));
  NO2        o034(.A(ori_ori_n23_), .B(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o035(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n33_), .Y(ori_ori_n46_));
  NO2        o036(.A(ori_ori_n24_), .B(ori_ori_n15_), .Y(ori_ori_n47_));
  NA2        o037(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n48_));
  NOi21      o038(.An(i_2_), .B(i_8_), .Y(ori_ori_n49_));
  NO2        o039(.A(ori_ori_n49_), .B(ori_ori_n40_), .Y(ori_ori_n50_));
  NO3        o040(.A(ori_ori_n50_), .B(ori_ori_n48_), .C(ori_ori_n47_), .Y(ori_ori_n51_));
  INV        o041(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NOi31      o042(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n53_));
  NA2        o043(.A(ori_ori_n53_), .B(i_0_), .Y(ori_ori_n54_));
  NOi21      o044(.An(i_4_), .B(i_3_), .Y(ori_ori_n55_));
  NOi21      o045(.An(i_1_), .B(i_4_), .Y(ori_ori_n56_));
  NA2        o046(.A(ori_ori_n56_), .B(ori_ori_n49_), .Y(ori_ori_n57_));
  NA2        o047(.A(ori_ori_n57_), .B(ori_ori_n54_), .Y(ori_ori_n58_));
  AN2        o048(.A(i_8_), .B(i_7_), .Y(ori_ori_n59_));
  INV        o049(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  NOi21      o050(.An(i_8_), .B(i_7_), .Y(ori_ori_n61_));
  NA2        o051(.A(ori_ori_n61_), .B(ori_ori_n55_), .Y(ori_ori_n62_));
  OAI210     o052(.A0(ori_ori_n60_), .A1(ori_ori_n48_), .B0(ori_ori_n62_), .Y(ori_ori_n63_));
  AOI220     o053(.A0(ori_ori_n63_), .A1(ori_ori_n34_), .B0(ori_ori_n58_), .B1(ori_ori_n37_), .Y(ori_ori_n64_));
  NA4        o054(.A(ori_ori_n64_), .B(ori_ori_n52_), .C(ori_ori_n46_), .D(ori_ori_n28_), .Y(ori_ori_n65_));
  NA2        o055(.A(i_8_), .B(ori_ori_n22_), .Y(ori_ori_n66_));
  AOI220     o056(.A0(ori_ori_n43_), .A1(i_1_), .B0(ori_ori_n41_), .B1(i_2_), .Y(ori_ori_n67_));
  NOi21      o057(.An(i_1_), .B(i_2_), .Y(ori_ori_n68_));
  NO2        o058(.A(ori_ori_n67_), .B(ori_ori_n66_), .Y(ori_ori_n69_));
  NA2        o059(.A(ori_ori_n69_), .B(ori_ori_n14_), .Y(ori_ori_n70_));
  NA2        o060(.A(ori_ori_n61_), .B(ori_ori_n12_), .Y(ori_ori_n71_));
  NA2        o061(.A(ori_ori_n25_), .B(ori_ori_n14_), .Y(ori_ori_n72_));
  NA2        o062(.A(ori_ori_n72_), .B(ori_ori_n71_), .Y(ori_ori_n73_));
  AN2        o063(.A(i_8_), .B(i_7_), .Y(ori_ori_n74_));
  NA2        o064(.A(ori_ori_n18_), .B(i_6_), .Y(ori_ori_n75_));
  INV        o065(.A(ori_ori_n75_), .Y(ori_ori_n76_));
  INV        o066(.A(i_0_), .Y(ori_ori_n77_));
  AOI220     o067(.A0(ori_ori_n77_), .A1(ori_ori_n76_), .B0(ori_ori_n73_), .B1(ori_ori_n55_), .Y(ori_ori_n78_));
  NA2        o068(.A(ori_ori_n78_), .B(ori_ori_n70_), .Y(ori_ori_n79_));
  NAi21      o069(.An(i_3_), .B(i_6_), .Y(ori_ori_n80_));
  NA2        o070(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n81_));
  NOi21      o071(.An(i_7_), .B(i_8_), .Y(ori_ori_n82_));
  NOi21      o072(.An(i_6_), .B(i_5_), .Y(ori_ori_n83_));
  AOI210     o073(.A0(ori_ori_n82_), .A1(ori_ori_n12_), .B0(ori_ori_n83_), .Y(ori_ori_n84_));
  OAI210     o074(.A0(ori_ori_n84_), .A1(ori_ori_n11_), .B0(ori_ori_n81_), .Y(ori_ori_n85_));
  NA2        o075(.A(ori_ori_n85_), .B(ori_ori_n68_), .Y(ori_ori_n86_));
  NA3        o076(.A(ori_ori_n24_), .B(i_2_), .C(ori_ori_n14_), .Y(ori_ori_n87_));
  INV        o077(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  NA3        o078(.A(ori_ori_n20_), .B(i_5_), .C(i_7_), .Y(ori_ori_n89_));
  NO2        o079(.A(ori_ori_n89_), .B(i_2_), .Y(ori_ori_n90_));
  NO2        o080(.A(ori_ori_n90_), .B(ori_ori_n88_), .Y(ori_ori_n91_));
  NA3        o081(.A(ori_ori_n61_), .B(ori_ori_n34_), .C(i_3_), .Y(ori_ori_n92_));
  NA2        o082(.A(ori_ori_n42_), .B(i_6_), .Y(ori_ori_n93_));
  NO2        o083(.A(ori_ori_n93_), .B(ori_ori_n92_), .Y(ori_ori_n94_));
  NAi21      o084(.An(i_6_), .B(i_0_), .Y(ori_ori_n95_));
  NA3        o085(.A(ori_ori_n56_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n96_));
  BUFFER     o086(.A(i_4_), .Y(ori_ori_n97_));
  INV        o087(.A(i_3_), .Y(ori_ori_n98_));
  NA3        o088(.A(ori_ori_n98_), .B(ori_ori_n68_), .C(ori_ori_n97_), .Y(ori_ori_n99_));
  OAI210     o089(.A0(ori_ori_n96_), .A1(ori_ori_n95_), .B0(ori_ori_n99_), .Y(ori_ori_n100_));
  NO2        o090(.A(ori_ori_n100_), .B(ori_ori_n94_), .Y(ori_ori_n101_));
  NOi21      o091(.An(i_3_), .B(i_1_), .Y(ori_ori_n102_));
  NA2        o092(.A(ori_ori_n102_), .B(i_4_), .Y(ori_ori_n103_));
  NO2        o093(.A(i_8_), .B(ori_ori_n103_), .Y(ori_ori_n104_));
  NOi31      o094(.An(ori_ori_n43_), .B(i_5_), .C(ori_ori_n34_), .Y(ori_ori_n105_));
  NO2        o095(.A(ori_ori_n105_), .B(ori_ori_n104_), .Y(ori_ori_n106_));
  NA4        o096(.A(ori_ori_n106_), .B(ori_ori_n101_), .C(ori_ori_n91_), .D(ori_ori_n86_), .Y(ori_ori_n107_));
  NA2        o097(.A(ori_ori_n36_), .B(ori_ori_n40_), .Y(ori_ori_n108_));
  INV        o098(.A(ori_ori_n55_), .Y(ori_ori_n109_));
  NO2        o099(.A(ori_ori_n109_), .B(ori_ori_n30_), .Y(ori_ori_n110_));
  NA2        o100(.A(ori_ori_n61_), .B(ori_ori_n53_), .Y(ori_ori_n111_));
  INV        o101(.A(ori_ori_n111_), .Y(ori_ori_n112_));
  NA3        o102(.A(ori_ori_n53_), .B(ori_ori_n14_), .C(i_7_), .Y(ori_ori_n113_));
  NA3        o103(.A(ori_ori_n37_), .B(ori_ori_n17_), .C(i_8_), .Y(ori_ori_n114_));
  NA4        o104(.A(ori_ori_n56_), .B(ori_ori_n43_), .C(i_5_), .D(ori_ori_n22_), .Y(ori_ori_n115_));
  NA3        o105(.A(ori_ori_n115_), .B(ori_ori_n114_), .C(ori_ori_n113_), .Y(ori_ori_n116_));
  NO3        o106(.A(ori_ori_n116_), .B(ori_ori_n112_), .C(ori_ori_n110_), .Y(ori_ori_n117_));
  INV        o107(.A(ori_ori_n82_), .Y(ori_ori_n118_));
  NO2        o108(.A(ori_ori_n118_), .B(ori_ori_n93_), .Y(ori_ori_n119_));
  NO3        o109(.A(i_2_), .B(ori_ori_n20_), .C(ori_ori_n14_), .Y(ori_ori_n120_));
  NA2        o110(.A(i_2_), .B(i_4_), .Y(ori_ori_n121_));
  AOI210     o111(.A0(ori_ori_n95_), .A1(ori_ori_n80_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  NO2        o112(.A(i_8_), .B(i_7_), .Y(ori_ori_n123_));
  OA210      o113(.A0(ori_ori_n122_), .A1(ori_ori_n120_), .B0(ori_ori_n123_), .Y(ori_ori_n124_));
  NA2        o114(.A(ori_ori_n102_), .B(i_0_), .Y(ori_ori_n125_));
  NO2        o115(.A(ori_ori_n125_), .B(i_4_), .Y(ori_ori_n126_));
  NO3        o116(.A(ori_ori_n126_), .B(ori_ori_n124_), .C(ori_ori_n119_), .Y(ori_ori_n127_));
  NA2        o117(.A(ori_ori_n82_), .B(ori_ori_n12_), .Y(ori_ori_n128_));
  INV        o118(.A(i_2_), .Y(ori_ori_n129_));
  NO2        o119(.A(ori_ori_n129_), .B(ori_ori_n128_), .Y(ori_ori_n130_));
  NO2        o120(.A(ori_ori_n92_), .B(ori_ori_n30_), .Y(ori_ori_n131_));
  NA3        o121(.A(ori_ori_n59_), .B(ori_ori_n42_), .C(ori_ori_n20_), .Y(ori_ori_n132_));
  NA3        o122(.A(ori_ori_n49_), .B(ori_ori_n35_), .C(ori_ori_n15_), .Y(ori_ori_n133_));
  NO2        o123(.A(i_2_), .B(i_1_), .Y(ori_ori_n134_));
  NA2        o124(.A(ori_ori_n74_), .B(ori_ori_n134_), .Y(ori_ori_n135_));
  NA3        o125(.A(ori_ori_n135_), .B(ori_ori_n133_), .C(ori_ori_n132_), .Y(ori_ori_n136_));
  NO3        o126(.A(ori_ori_n136_), .B(ori_ori_n131_), .C(ori_ori_n130_), .Y(ori_ori_n137_));
  NA4        o127(.A(ori_ori_n137_), .B(ori_ori_n127_), .C(ori_ori_n117_), .D(ori_ori_n108_), .Y(ori_ori_n138_));
  OR4        o128(.A(ori_ori_n138_), .B(ori_ori_n107_), .C(ori_ori_n79_), .D(ori_ori_n65_), .Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NO2        m008(.A(mai_mai_n16_), .B(mai_mai_n13_), .Y(mai_mai_n19_));
  INV        m009(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m010(.A(i_0_), .B(mai_mai_n20_), .Y(mai_mai_n21_));
  INV        m011(.A(i_7_), .Y(mai_mai_n22_));
  NA3        m012(.A(i_6_), .B(i_5_), .C(mai_mai_n22_), .Y(mai_mai_n23_));
  NOi21      m013(.An(i_8_), .B(i_6_), .Y(mai_mai_n24_));
  AOI210     m014(.A0(mai_mai_n154_), .A1(mai_mai_n23_), .B0(mai_mai_n21_), .Y(mai_mai_n25_));
  AOI210     m015(.A0(mai_mai_n25_), .A1(mai_mai_n11_), .B0(mai_mai_n19_), .Y(mai_mai_n26_));
  NA2        m016(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n27_));
  NO2        m017(.A(i_2_), .B(i_4_), .Y(mai_mai_n28_));
  NA3        m018(.A(mai_mai_n28_), .B(i_6_), .C(i_8_), .Y(mai_mai_n29_));
  AOI210     m019(.A0(mai_mai_n27_), .A1(i_5_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  INV        m020(.A(i_2_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_5_), .B(i_0_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_6_), .B(i_8_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_7_), .B(i_1_), .Y(mai_mai_n34_));
  BUFFER     m024(.A(i_5_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_0_), .B(i_4_), .Y(mai_mai_n36_));
  XO2        m026(.A(i_1_), .B(i_3_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_7_), .B(i_5_), .Y(mai_mai_n38_));
  INV        m028(.A(i_1_), .Y(mai_mai_n39_));
  NOi21      m029(.An(i_3_), .B(i_0_), .Y(mai_mai_n40_));
  NA2        m030(.A(mai_mai_n40_), .B(mai_mai_n39_), .Y(mai_mai_n41_));
  NA3        m031(.A(i_6_), .B(mai_mai_n14_), .C(i_7_), .Y(mai_mai_n42_));
  AOI210     m032(.A0(mai_mai_n42_), .A1(mai_mai_n23_), .B0(mai_mai_n41_), .Y(mai_mai_n43_));
  NO2        m033(.A(mai_mai_n43_), .B(mai_mai_n30_), .Y(mai_mai_n44_));
  NOi21      m034(.An(i_4_), .B(i_0_), .Y(mai_mai_n45_));
  AOI210     m035(.A0(mai_mai_n45_), .A1(mai_mai_n24_), .B0(mai_mai_n15_), .Y(mai_mai_n46_));
  NA2        m036(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n47_));
  NOi21      m037(.An(i_2_), .B(i_8_), .Y(mai_mai_n48_));
  NO3        m038(.A(mai_mai_n48_), .B(mai_mai_n45_), .C(mai_mai_n36_), .Y(mai_mai_n49_));
  NO3        m039(.A(mai_mai_n49_), .B(mai_mai_n47_), .C(mai_mai_n46_), .Y(mai_mai_n50_));
  INV        m040(.A(mai_mai_n50_), .Y(mai_mai_n51_));
  NOi31      m041(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_4_), .B(i_3_), .Y(mai_mai_n53_));
  NOi21      m043(.An(i_1_), .B(i_4_), .Y(mai_mai_n54_));
  AN2        m044(.A(i_8_), .B(i_7_), .Y(mai_mai_n55_));
  NA2        m045(.A(mai_mai_n55_), .B(mai_mai_n12_), .Y(mai_mai_n56_));
  NOi21      m046(.An(i_8_), .B(i_7_), .Y(mai_mai_n57_));
  NA3        m047(.A(mai_mai_n57_), .B(mai_mai_n53_), .C(i_6_), .Y(mai_mai_n58_));
  OAI210     m048(.A0(mai_mai_n56_), .A1(mai_mai_n47_), .B0(mai_mai_n58_), .Y(mai_mai_n59_));
  AOI220     m049(.A0(mai_mai_n59_), .A1(mai_mai_n31_), .B0(mai_mai_n52_), .B1(mai_mai_n35_), .Y(mai_mai_n60_));
  NA4        m050(.A(mai_mai_n60_), .B(mai_mai_n51_), .C(mai_mai_n44_), .D(mai_mai_n26_), .Y(mai_mai_n61_));
  NA2        m051(.A(i_8_), .B(mai_mai_n22_), .Y(mai_mai_n62_));
  AOI220     m052(.A0(mai_mai_n40_), .A1(i_1_), .B0(mai_mai_n37_), .B1(i_2_), .Y(mai_mai_n63_));
  NOi21      m053(.An(i_1_), .B(i_2_), .Y(mai_mai_n64_));
  NO2        m054(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n65_));
  NA2        m055(.A(mai_mai_n65_), .B(mai_mai_n14_), .Y(mai_mai_n66_));
  NA3        m056(.A(mai_mai_n57_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n67_));
  NA3        m057(.A(i_1_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n68_));
  NA2        m058(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  NOi32      m059(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n70_));
  NA2        m060(.A(mai_mai_n70_), .B(i_3_), .Y(mai_mai_n71_));
  NA3        m061(.A(mai_mai_n18_), .B(i_2_), .C(i_6_), .Y(mai_mai_n72_));
  NA2        m062(.A(mai_mai_n72_), .B(mai_mai_n71_), .Y(mai_mai_n73_));
  NO2        m063(.A(i_0_), .B(i_4_), .Y(mai_mai_n74_));
  AOI220     m064(.A0(mai_mai_n74_), .A1(mai_mai_n73_), .B0(mai_mai_n69_), .B1(mai_mai_n53_), .Y(mai_mai_n75_));
  NA2        m065(.A(mai_mai_n75_), .B(mai_mai_n66_), .Y(mai_mai_n76_));
  NA2        m066(.A(mai_mai_n33_), .B(mai_mai_n32_), .Y(mai_mai_n77_));
  NOi21      m067(.An(i_7_), .B(i_8_), .Y(mai_mai_n78_));
  NOi31      m068(.An(i_6_), .B(i_5_), .C(i_7_), .Y(mai_mai_n79_));
  AOI210     m069(.A0(mai_mai_n78_), .A1(mai_mai_n12_), .B0(mai_mai_n79_), .Y(mai_mai_n80_));
  OAI210     m070(.A0(mai_mai_n80_), .A1(mai_mai_n11_), .B0(mai_mai_n77_), .Y(mai_mai_n81_));
  NA2        m071(.A(mai_mai_n81_), .B(mai_mai_n64_), .Y(mai_mai_n82_));
  AOI220     m072(.A0(mai_mai_n40_), .A1(mai_mai_n39_), .B0(mai_mai_n18_), .B1(mai_mai_n31_), .Y(mai_mai_n83_));
  NA3        m073(.A(mai_mai_n20_), .B(i_5_), .C(i_7_), .Y(mai_mai_n84_));
  NO2        m074(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n85_));
  INV        m075(.A(mai_mai_n85_), .Y(mai_mai_n86_));
  NA3        m076(.A(mai_mai_n57_), .B(mai_mai_n31_), .C(i_3_), .Y(mai_mai_n87_));
  NA2        m077(.A(mai_mai_n39_), .B(i_6_), .Y(mai_mai_n88_));
  AOI210     m078(.A0(mai_mai_n88_), .A1(mai_mai_n21_), .B0(mai_mai_n87_), .Y(mai_mai_n89_));
  NOi21      m079(.An(i_2_), .B(i_1_), .Y(mai_mai_n90_));
  NAi21      m080(.An(i_6_), .B(i_0_), .Y(mai_mai_n91_));
  NOi21      m081(.An(i_4_), .B(i_6_), .Y(mai_mai_n92_));
  NOi21      m082(.An(i_5_), .B(i_3_), .Y(mai_mai_n93_));
  NA3        m083(.A(mai_mai_n93_), .B(mai_mai_n64_), .C(mai_mai_n92_), .Y(mai_mai_n94_));
  INV        m084(.A(mai_mai_n94_), .Y(mai_mai_n95_));
  NA2        m085(.A(mai_mai_n64_), .B(mai_mai_n33_), .Y(mai_mai_n96_));
  NOi21      m086(.An(mai_mai_n38_), .B(mai_mai_n96_), .Y(mai_mai_n97_));
  NO3        m087(.A(mai_mai_n97_), .B(mai_mai_n95_), .C(mai_mai_n89_), .Y(mai_mai_n98_));
  NOi31      m088(.An(mai_mai_n45_), .B(mai_mai_n155_), .C(i_2_), .Y(mai_mai_n99_));
  NA2        m089(.A(mai_mai_n57_), .B(mai_mai_n12_), .Y(mai_mai_n100_));
  NA2        m090(.A(mai_mai_n33_), .B(mai_mai_n14_), .Y(mai_mai_n101_));
  NOi21      m091(.An(i_3_), .B(i_1_), .Y(mai_mai_n102_));
  NA2        m092(.A(mai_mai_n102_), .B(i_4_), .Y(mai_mai_n103_));
  AOI210     m093(.A0(mai_mai_n101_), .A1(mai_mai_n100_), .B0(mai_mai_n103_), .Y(mai_mai_n104_));
  AOI220     m094(.A0(mai_mai_n78_), .A1(mai_mai_n14_), .B0(mai_mai_n92_), .B1(mai_mai_n22_), .Y(mai_mai_n105_));
  NOi31      m095(.An(mai_mai_n40_), .B(mai_mai_n105_), .C(mai_mai_n31_), .Y(mai_mai_n106_));
  NO3        m096(.A(mai_mai_n106_), .B(mai_mai_n104_), .C(mai_mai_n99_), .Y(mai_mai_n107_));
  NA4        m097(.A(mai_mai_n107_), .B(mai_mai_n98_), .C(mai_mai_n86_), .D(mai_mai_n82_), .Y(mai_mai_n108_));
  NA2        m098(.A(mai_mai_n48_), .B(mai_mai_n15_), .Y(mai_mai_n109_));
  NOi31      m099(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n110_));
  NOi31      m100(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n111_));
  OAI210     m101(.A0(mai_mai_n111_), .A1(mai_mai_n110_), .B0(i_7_), .Y(mai_mai_n112_));
  NA3        m102(.A(mai_mai_n33_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n113_));
  NA4        m103(.A(mai_mai_n113_), .B(mai_mai_n112_), .C(mai_mai_n109_), .D(mai_mai_n96_), .Y(mai_mai_n114_));
  NA2        m104(.A(mai_mai_n114_), .B(mai_mai_n36_), .Y(mai_mai_n115_));
  NA3        m105(.A(mai_mai_n55_), .B(mai_mai_n90_), .C(mai_mai_n12_), .Y(mai_mai_n116_));
  NAi31      m106(.An(mai_mai_n91_), .B(mai_mai_n78_), .C(mai_mai_n90_), .Y(mai_mai_n117_));
  NA3        m107(.A(mai_mai_n57_), .B(mai_mai_n52_), .C(i_6_), .Y(mai_mai_n118_));
  NA3        m108(.A(mai_mai_n118_), .B(mai_mai_n117_), .C(mai_mai_n116_), .Y(mai_mai_n119_));
  NOi21      m109(.An(i_0_), .B(i_2_), .Y(mai_mai_n120_));
  NA3        m110(.A(mai_mai_n120_), .B(mai_mai_n34_), .C(mai_mai_n92_), .Y(mai_mai_n121_));
  NA3        m111(.A(mai_mai_n45_), .B(mai_mai_n38_), .C(mai_mai_n18_), .Y(mai_mai_n122_));
  NA3        m112(.A(mai_mai_n120_), .B(mai_mai_n53_), .C(mai_mai_n33_), .Y(mai_mai_n123_));
  NA3        m113(.A(mai_mai_n123_), .B(mai_mai_n122_), .C(mai_mai_n121_), .Y(mai_mai_n124_));
  NA4        m114(.A(mai_mai_n52_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n125_));
  NA4        m115(.A(mai_mai_n54_), .B(mai_mai_n35_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n126_));
  NA2        m116(.A(mai_mai_n126_), .B(mai_mai_n125_), .Y(mai_mai_n127_));
  NO3        m117(.A(mai_mai_n127_), .B(mai_mai_n124_), .C(mai_mai_n119_), .Y(mai_mai_n128_));
  NO2        m118(.A(mai_mai_n109_), .B(mai_mai_n88_), .Y(mai_mai_n129_));
  NO3        m119(.A(i_2_), .B(mai_mai_n11_), .C(mai_mai_n14_), .Y(mai_mai_n130_));
  NA2        m120(.A(i_2_), .B(i_4_), .Y(mai_mai_n131_));
  AOI210     m121(.A0(mai_mai_n91_), .A1(i_3_), .B0(mai_mai_n131_), .Y(mai_mai_n132_));
  NO2        m122(.A(i_8_), .B(i_7_), .Y(mai_mai_n133_));
  OA210      m123(.A0(mai_mai_n132_), .A1(mai_mai_n130_), .B0(mai_mai_n133_), .Y(mai_mai_n134_));
  NA3        m124(.A(mai_mai_n102_), .B(i_5_), .C(mai_mai_n22_), .Y(mai_mai_n135_));
  NO2        m125(.A(mai_mai_n135_), .B(i_4_), .Y(mai_mai_n136_));
  NO3        m126(.A(mai_mai_n136_), .B(mai_mai_n134_), .C(mai_mai_n129_), .Y(mai_mai_n137_));
  NA2        m127(.A(mai_mai_n78_), .B(mai_mai_n12_), .Y(mai_mai_n138_));
  NA3        m128(.A(i_2_), .B(i_1_), .C(mai_mai_n14_), .Y(mai_mai_n139_));
  INV        m129(.A(mai_mai_n45_), .Y(mai_mai_n140_));
  AOI210     m130(.A0(mai_mai_n140_), .A1(mai_mai_n139_), .B0(mai_mai_n138_), .Y(mai_mai_n141_));
  NA3        m131(.A(mai_mai_n120_), .B(mai_mai_n57_), .C(mai_mai_n92_), .Y(mai_mai_n142_));
  OAI210     m132(.A0(mai_mai_n87_), .A1(mai_mai_n27_), .B0(mai_mai_n142_), .Y(mai_mai_n143_));
  NA3        m133(.A(mai_mai_n93_), .B(mai_mai_n55_), .C(mai_mai_n39_), .Y(mai_mai_n144_));
  NA2        m134(.A(mai_mai_n48_), .B(mai_mai_n32_), .Y(mai_mai_n145_));
  NOi31      m135(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n146_));
  NA2        m136(.A(mai_mai_n70_), .B(mai_mai_n146_), .Y(mai_mai_n147_));
  NA3        m137(.A(mai_mai_n147_), .B(mai_mai_n145_), .C(mai_mai_n144_), .Y(mai_mai_n148_));
  NO3        m138(.A(mai_mai_n148_), .B(mai_mai_n143_), .C(mai_mai_n141_), .Y(mai_mai_n149_));
  NA4        m139(.A(mai_mai_n149_), .B(mai_mai_n137_), .C(mai_mai_n128_), .D(mai_mai_n115_), .Y(mai_mai_n150_));
  OR4        m140(.A(mai_mai_n150_), .B(mai_mai_n108_), .C(mai_mai_n76_), .D(mai_mai_n61_), .Y(mai00));
  INV        m141(.A(i_1_), .Y(mai_mai_n154_));
  INV        m142(.A(i_7_), .Y(mai_mai_n155_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  INV        u005(.A(i_0_), .Y(men_men_n16_));
  NOi21      u006(.An(i_1_), .B(i_3_), .Y(men_men_n17_));
  NA3        u007(.A(men_men_n17_), .B(men_men_n16_), .C(i_2_), .Y(men_men_n18_));
  NO2        u008(.A(men_men_n18_), .B(men_men_n13_), .Y(men_men_n19_));
  INV        u009(.A(i_4_), .Y(men_men_n20_));
  NA2        u010(.A(i_0_), .B(men_men_n20_), .Y(men_men_n21_));
  INV        u011(.A(i_7_), .Y(men_men_n22_));
  NA3        u012(.A(i_6_), .B(i_5_), .C(men_men_n22_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  NOi21      u014(.An(i_1_), .B(i_8_), .Y(men_men_n25_));
  AOI220     u015(.A0(men_men_n25_), .A1(i_2_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n26_));
  AOI210     u016(.A0(men_men_n26_), .A1(men_men_n23_), .B0(men_men_n21_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n11_), .B0(men_men_n19_), .Y(men_men_n28_));
  NA2        u018(.A(i_0_), .B(men_men_n14_), .Y(men_men_n29_));
  NA2        u019(.A(men_men_n16_), .B(i_5_), .Y(men_men_n30_));
  NO2        u020(.A(i_2_), .B(i_4_), .Y(men_men_n31_));
  NA3        u021(.A(men_men_n31_), .B(i_6_), .C(i_8_), .Y(men_men_n32_));
  AOI210     u022(.A0(men_men_n30_), .A1(men_men_n29_), .B0(men_men_n32_), .Y(men_men_n33_));
  INV        u023(.A(i_2_), .Y(men_men_n34_));
  NOi21      u024(.An(i_5_), .B(i_0_), .Y(men_men_n35_));
  NOi21      u025(.An(i_6_), .B(i_8_), .Y(men_men_n36_));
  NOi21      u026(.An(i_7_), .B(i_1_), .Y(men_men_n37_));
  NOi21      u027(.An(i_5_), .B(i_6_), .Y(men_men_n38_));
  AOI220     u028(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n36_), .B1(men_men_n35_), .Y(men_men_n39_));
  NO3        u029(.A(men_men_n39_), .B(men_men_n34_), .C(i_4_), .Y(men_men_n40_));
  NOi21      u030(.An(i_0_), .B(i_4_), .Y(men_men_n41_));
  XO2        u031(.A(i_1_), .B(i_3_), .Y(men_men_n42_));
  NOi21      u032(.An(i_7_), .B(i_5_), .Y(men_men_n43_));
  AN3        u033(.A(men_men_n43_), .B(men_men_n42_), .C(men_men_n41_), .Y(men_men_n44_));
  INV        u034(.A(i_1_), .Y(men_men_n45_));
  NOi21      u035(.An(i_3_), .B(i_0_), .Y(men_men_n46_));
  NA2        u036(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  AOI210     u037(.A0(men_men_n156_), .A1(men_men_n23_), .B0(men_men_n47_), .Y(men_men_n48_));
  NO4        u038(.A(men_men_n48_), .B(men_men_n44_), .C(men_men_n40_), .D(men_men_n33_), .Y(men_men_n49_));
  INV        u039(.A(i_8_), .Y(men_men_n50_));
  NA2        u040(.A(i_1_), .B(men_men_n11_), .Y(men_men_n51_));
  NOi21      u041(.An(i_4_), .B(i_0_), .Y(men_men_n52_));
  AOI210     u042(.A0(men_men_n52_), .A1(men_men_n24_), .B0(men_men_n15_), .Y(men_men_n53_));
  NA2        u043(.A(i_1_), .B(men_men_n14_), .Y(men_men_n54_));
  NOi21      u044(.An(i_2_), .B(i_8_), .Y(men_men_n55_));
  NO2        u045(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n56_));
  INV        u046(.A(men_men_n56_), .Y(men_men_n57_));
  NOi31      u047(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n58_), .B(i_0_), .Y(men_men_n59_));
  NOi21      u049(.An(i_4_), .B(i_3_), .Y(men_men_n60_));
  NOi21      u050(.An(i_1_), .B(i_4_), .Y(men_men_n61_));
  OAI210     u051(.A0(men_men_n61_), .A1(men_men_n60_), .B0(men_men_n55_), .Y(men_men_n62_));
  NA2        u052(.A(men_men_n62_), .B(men_men_n59_), .Y(men_men_n63_));
  AN2        u053(.A(i_8_), .B(i_7_), .Y(men_men_n64_));
  NOi21      u054(.An(i_8_), .B(i_7_), .Y(men_men_n65_));
  NA3        u055(.A(men_men_n65_), .B(men_men_n60_), .C(i_6_), .Y(men_men_n66_));
  INV        u056(.A(men_men_n66_), .Y(men_men_n67_));
  AOI220     u057(.A0(men_men_n67_), .A1(men_men_n34_), .B0(men_men_n63_), .B1(men_men_n38_), .Y(men_men_n68_));
  NA4        u058(.A(men_men_n68_), .B(men_men_n57_), .C(men_men_n49_), .D(men_men_n28_), .Y(men_men_n69_));
  NA2        u059(.A(i_8_), .B(i_7_), .Y(men_men_n70_));
  NO3        u060(.A(men_men_n70_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n71_));
  NA2        u061(.A(i_8_), .B(men_men_n22_), .Y(men_men_n72_));
  NA2        u062(.A(men_men_n42_), .B(i_2_), .Y(men_men_n73_));
  NOi21      u063(.An(i_1_), .B(i_2_), .Y(men_men_n74_));
  NA3        u064(.A(men_men_n74_), .B(men_men_n52_), .C(i_6_), .Y(men_men_n75_));
  OAI210     u065(.A0(men_men_n73_), .A1(men_men_n72_), .B0(men_men_n75_), .Y(men_men_n76_));
  OAI210     u066(.A0(men_men_n76_), .A1(men_men_n71_), .B0(men_men_n14_), .Y(men_men_n77_));
  NA3        u067(.A(men_men_n65_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n78_));
  INV        u068(.A(men_men_n78_), .Y(men_men_n79_));
  NOi32      u069(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n80_));
  NA2        u070(.A(men_men_n80_), .B(i_3_), .Y(men_men_n81_));
  NA3        u071(.A(men_men_n17_), .B(i_2_), .C(i_6_), .Y(men_men_n82_));
  NA2        u072(.A(men_men_n82_), .B(men_men_n81_), .Y(men_men_n83_));
  NO2        u073(.A(i_0_), .B(i_4_), .Y(men_men_n84_));
  AOI220     u074(.A0(men_men_n84_), .A1(men_men_n83_), .B0(men_men_n79_), .B1(men_men_n60_), .Y(men_men_n85_));
  NA2        u075(.A(men_men_n85_), .B(men_men_n77_), .Y(men_men_n86_));
  NAi21      u076(.An(i_3_), .B(i_6_), .Y(men_men_n87_));
  NO3        u077(.A(men_men_n87_), .B(i_0_), .C(men_men_n50_), .Y(men_men_n88_));
  NA2        u078(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n89_));
  NOi21      u079(.An(i_7_), .B(i_8_), .Y(men_men_n90_));
  NOi31      u080(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n91_));
  OAI210     u081(.A0(i_6_), .A1(men_men_n11_), .B0(men_men_n89_), .Y(men_men_n92_));
  OAI210     u082(.A0(men_men_n92_), .A1(men_men_n88_), .B0(men_men_n74_), .Y(men_men_n93_));
  NA3        u083(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n94_));
  AOI210     u084(.A0(men_men_n21_), .A1(men_men_n51_), .B0(men_men_n94_), .Y(men_men_n95_));
  OAI210     u085(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n96_));
  NA3        u086(.A(men_men_n70_), .B(men_men_n17_), .C(men_men_n16_), .Y(men_men_n97_));
  NO2        u087(.A(men_men_n97_), .B(men_men_n96_), .Y(men_men_n98_));
  NO2        u088(.A(men_men_n98_), .B(men_men_n95_), .Y(men_men_n99_));
  NA3        u089(.A(men_men_n65_), .B(men_men_n34_), .C(i_3_), .Y(men_men_n100_));
  NA2        u090(.A(men_men_n45_), .B(i_6_), .Y(men_men_n101_));
  NOi21      u091(.An(i_2_), .B(i_1_), .Y(men_men_n102_));
  NAi21      u092(.An(i_6_), .B(i_0_), .Y(men_men_n103_));
  NOi21      u093(.An(i_4_), .B(i_6_), .Y(men_men_n104_));
  NA2        u094(.A(men_men_n74_), .B(men_men_n36_), .Y(men_men_n105_));
  NA2        u095(.A(men_men_n24_), .B(i_5_), .Y(men_men_n106_));
  NOi31      u096(.An(men_men_n52_), .B(men_men_n106_), .C(i_2_), .Y(men_men_n107_));
  INV        u097(.A(men_men_n107_), .Y(men_men_n108_));
  NA4        u098(.A(men_men_n108_), .B(men_men_n100_), .C(men_men_n99_), .D(men_men_n93_), .Y(men_men_n109_));
  NA2        u099(.A(men_men_n55_), .B(men_men_n15_), .Y(men_men_n110_));
  NOi31      u100(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n111_));
  NOi31      u101(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n112_));
  OAI210     u102(.A0(men_men_n112_), .A1(men_men_n111_), .B0(i_7_), .Y(men_men_n113_));
  NA3        u103(.A(men_men_n113_), .B(men_men_n110_), .C(men_men_n105_), .Y(men_men_n114_));
  NA2        u104(.A(men_men_n114_), .B(men_men_n41_), .Y(men_men_n115_));
  NA2        u105(.A(men_men_n60_), .B(men_men_n37_), .Y(men_men_n116_));
  AOI210     u106(.A0(men_men_n116_), .A1(men_men_n78_), .B0(men_men_n30_), .Y(men_men_n117_));
  NAi31      u107(.An(men_men_n103_), .B(men_men_n90_), .C(men_men_n102_), .Y(men_men_n118_));
  NA3        u108(.A(men_men_n65_), .B(men_men_n58_), .C(i_6_), .Y(men_men_n119_));
  NA2        u109(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NOi21      u110(.An(i_0_), .B(i_2_), .Y(men_men_n121_));
  NOi32      u111(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n122_));
  NA2        u112(.A(men_men_n122_), .B(men_men_n111_), .Y(men_men_n123_));
  NA3        u113(.A(men_men_n121_), .B(men_men_n60_), .C(men_men_n36_), .Y(men_men_n124_));
  NA2        u114(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NA3        u115(.A(men_men_n58_), .B(i_6_), .C(men_men_n14_), .Y(men_men_n126_));
  NA4        u116(.A(men_men_n61_), .B(men_men_n38_), .C(men_men_n16_), .D(i_8_), .Y(men_men_n127_));
  NA2        u117(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n128_));
  NO4        u118(.A(men_men_n128_), .B(men_men_n125_), .C(men_men_n120_), .D(men_men_n117_), .Y(men_men_n129_));
  NOi21      u119(.An(i_5_), .B(i_2_), .Y(men_men_n130_));
  AOI220     u120(.A0(men_men_n130_), .A1(men_men_n90_), .B0(men_men_n64_), .B1(men_men_n31_), .Y(men_men_n131_));
  AOI210     u121(.A0(men_men_n131_), .A1(men_men_n110_), .B0(men_men_n101_), .Y(men_men_n132_));
  NO4        u122(.A(i_2_), .B(men_men_n20_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n133_));
  NA2        u123(.A(i_2_), .B(i_4_), .Y(men_men_n134_));
  AOI210     u124(.A0(men_men_n103_), .A1(men_men_n87_), .B0(men_men_n134_), .Y(men_men_n135_));
  NO2        u125(.A(i_8_), .B(i_7_), .Y(men_men_n136_));
  OA210      u126(.A0(men_men_n135_), .A1(men_men_n133_), .B0(men_men_n136_), .Y(men_men_n137_));
  NA4        u127(.A(i_3_), .B(i_0_), .C(i_5_), .D(men_men_n22_), .Y(men_men_n138_));
  NO2        u128(.A(men_men_n138_), .B(i_4_), .Y(men_men_n139_));
  NO3        u129(.A(men_men_n139_), .B(men_men_n137_), .C(men_men_n132_), .Y(men_men_n140_));
  INV        u130(.A(men_men_n90_), .Y(men_men_n141_));
  NA2        u131(.A(i_1_), .B(men_men_n14_), .Y(men_men_n142_));
  NO2        u132(.A(men_men_n142_), .B(men_men_n141_), .Y(men_men_n143_));
  NA2        u133(.A(men_men_n121_), .B(men_men_n104_), .Y(men_men_n144_));
  INV        u134(.A(men_men_n144_), .Y(men_men_n145_));
  NA2        u135(.A(men_men_n91_), .B(i_3_), .Y(men_men_n146_));
  NA3        u136(.A(men_men_n55_), .B(men_men_n35_), .C(men_men_n15_), .Y(men_men_n147_));
  NOi31      u137(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n148_));
  OAI210     u138(.A0(men_men_n122_), .A1(men_men_n80_), .B0(men_men_n148_), .Y(men_men_n149_));
  NA3        u139(.A(men_men_n149_), .B(men_men_n147_), .C(men_men_n146_), .Y(men_men_n150_));
  NO3        u140(.A(men_men_n150_), .B(men_men_n145_), .C(men_men_n143_), .Y(men_men_n151_));
  NA4        u141(.A(men_men_n151_), .B(men_men_n140_), .C(men_men_n129_), .D(men_men_n115_), .Y(men_men_n152_));
  OR4        u142(.A(men_men_n152_), .B(men_men_n109_), .C(men_men_n86_), .D(men_men_n69_), .Y(men00));
  INV        u143(.A(i_7_), .Y(men_men_n156_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule