//Benchmark atmr_intb_466_0.25

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n152_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n285_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n383_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n454_, men_men_n455_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  INV        o026(.A(x09), .Y(ori_ori_n49_));
  NO2        o027(.A(x10), .B(x02), .Y(ori_ori_n50_));
  NOi21      o028(.An(x01), .B(x09), .Y(ori_ori_n51_));
  INV        o029(.A(x00), .Y(ori_ori_n52_));
  NO2        o030(.A(ori_ori_n49_), .B(ori_ori_n52_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(ori_ori_n51_), .Y(ori_ori_n54_));
  NA2        o032(.A(x09), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  INV        o033(.A(x07), .Y(ori_ori_n56_));
  INV        o034(.A(ori_ori_n54_), .Y(ori_ori_n57_));
  NO2        o035(.A(x02), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n58_), .B(ori_ori_n31_), .Y(ori_ori_n59_));
  NO2        o037(.A(ori_ori_n59_), .B(x05), .Y(ori_ori_n60_));
  NO2        o038(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n61_));
  NO2        o039(.A(x08), .B(x01), .Y(ori_ori_n62_));
  OAI210     o040(.A0(ori_ori_n62_), .A1(ori_ori_n61_), .B0(ori_ori_n35_), .Y(ori_ori_n63_));
  NO2        o041(.A(ori_ori_n63_), .B(x02), .Y(ori_ori_n64_));
  AN2        o042(.A(ori_ori_n64_), .B(ori_ori_n170_), .Y(ori_ori_n65_));
  INV        o043(.A(ori_ori_n63_), .Y(ori_ori_n66_));
  NA2        o044(.A(x11), .B(x00), .Y(ori_ori_n67_));
  NO2        o045(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n68_));
  NOi21      o046(.An(ori_ori_n67_), .B(ori_ori_n68_), .Y(ori_ori_n69_));
  INV        o047(.A(ori_ori_n69_), .Y(ori_ori_n70_));
  NOi21      o048(.An(x01), .B(x10), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n29_), .B(ori_ori_n52_), .Y(ori_ori_n72_));
  NO3        o050(.A(ori_ori_n72_), .B(ori_ori_n71_), .C(x06), .Y(ori_ori_n73_));
  NA2        o051(.A(ori_ori_n73_), .B(ori_ori_n27_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n70_), .A1(x07), .B0(ori_ori_n74_), .Y(ori_ori_n75_));
  NO3        o053(.A(ori_ori_n75_), .B(ori_ori_n65_), .C(ori_ori_n60_), .Y(ori01));
  INV        o054(.A(x12), .Y(ori_ori_n77_));
  INV        o055(.A(x13), .Y(ori_ori_n78_));
  NA2        o056(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n79_));
  NA2        o057(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n80_));
  NO2        o058(.A(ori_ori_n80_), .B(x05), .Y(ori_ori_n81_));
  NA2        o059(.A(ori_ori_n35_), .B(ori_ori_n52_), .Y(ori_ori_n82_));
  NA2        o060(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n83_));
  NA2        o061(.A(x10), .B(ori_ori_n52_), .Y(ori_ori_n84_));
  NA2        o062(.A(ori_ori_n84_), .B(ori_ori_n83_), .Y(ori_ori_n85_));
  NA2        o063(.A(ori_ori_n49_), .B(x05), .Y(ori_ori_n86_));
  NO2        o064(.A(ori_ori_n55_), .B(x05), .Y(ori_ori_n87_));
  NO2        o065(.A(ori_ori_n49_), .B(ori_ori_n41_), .Y(ori_ori_n88_));
  NO2        o066(.A(x09), .B(x05), .Y(ori_ori_n89_));
  NA2        o067(.A(ori_ori_n89_), .B(ori_ori_n47_), .Y(ori_ori_n90_));
  NO2        o068(.A(x03), .B(x02), .Y(ori_ori_n91_));
  NA2        o069(.A(ori_ori_n63_), .B(ori_ori_n78_), .Y(ori_ori_n92_));
  NA2        o070(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n94_));
  NO2        o072(.A(x09), .B(x01), .Y(ori_ori_n95_));
  NA2        o073(.A(x01), .B(ori_ori_n84_), .Y(ori_ori_n96_));
  NA2        o074(.A(x06), .B(x05), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n97_), .B(ori_ori_n77_), .Y(ori_ori_n98_));
  AOI210     o076(.A0(x10), .A1(ori_ori_n53_), .B0(ori_ori_n98_), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n99_), .B(ori_ori_n96_), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n78_), .B(x12), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n102_));
  NO2        o080(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n103_), .B(x02), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n102_), .B(ori_ori_n100_), .Y(ori_ori_n105_));
  INV        o083(.A(ori_ori_n105_), .Y(ori_ori_n106_));
  AOI210     o084(.A0(ori_ori_n171_), .A1(ori_ori_n77_), .B0(ori_ori_n106_), .Y(ori_ori_n107_));
  NO2        o085(.A(ori_ori_n49_), .B(x03), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n109_));
  NA2        o087(.A(x13), .B(ori_ori_n77_), .Y(ori_ori_n110_));
  NA3        o088(.A(ori_ori_n110_), .B(ori_ori_n98_), .C(ori_ori_n69_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(x07), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n49_), .B(ori_ori_n41_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n113_), .B(x01), .Y(ori_ori_n114_));
  NO2        o092(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n115_));
  NA2        o093(.A(x06), .B(ori_ori_n115_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n109_), .B(ori_ori_n28_), .Y(ori_ori_n117_));
  OAI210     o095(.A0(ori_ori_n72_), .A1(x06), .B0(ori_ori_n117_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n118_), .B(ori_ori_n116_), .Y(ori_ori_n119_));
  NO2        o097(.A(ori_ori_n119_), .B(ori_ori_n112_), .Y(ori_ori_n120_));
  OAI210     o098(.A0(ori_ori_n107_), .A1(ori_ori_n56_), .B0(ori_ori_n120_), .Y(ori02));
  NA2        o099(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n88_), .B(x03), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n77_), .B(ori_ori_n41_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n124_), .B(ori_ori_n85_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n125_), .B(ori_ori_n48_), .Y(ori_ori_n126_));
  INV        o104(.A(ori_ori_n103_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n128_));
  OAI210     o106(.A0(ori_ori_n127_), .A1(ori_ori_n54_), .B0(ori_ori_n128_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n129_), .B(x02), .Y(ori_ori_n130_));
  NO3        o108(.A(ori_ori_n101_), .B(ori_ori_n94_), .C(ori_ori_n50_), .Y(ori_ori_n131_));
  OAI210     o109(.A0(x12), .A1(x01), .B0(ori_ori_n131_), .Y(ori_ori_n132_));
  NA3        o110(.A(ori_ori_n132_), .B(ori_ori_n130_), .C(x06), .Y(ori_ori_n133_));
  NA2        o111(.A(ori_ori_n133_), .B(ori_ori_n126_), .Y(ori_ori_n134_));
  OAI210     o112(.A0(ori_ori_n122_), .A1(x12), .B0(ori_ori_n134_), .Y(ori03));
  OR2        o113(.A(ori_ori_n42_), .B(ori_ori_n108_), .Y(ori_ori_n136_));
  AOI210     o114(.A0(ori_ori_n92_), .A1(ori_ori_n77_), .B0(ori_ori_n136_), .Y(ori_ori_n137_));
  NA2        o115(.A(ori_ori_n101_), .B(ori_ori_n91_), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n138_), .B(ori_ori_n104_), .Y(ori_ori_n139_));
  OAI210     o117(.A0(ori_ori_n139_), .A1(ori_ori_n137_), .B0(x05), .Y(ori_ori_n140_));
  INV        o118(.A(ori_ori_n81_), .Y(ori_ori_n141_));
  NO2        o119(.A(ori_ori_n141_), .B(ori_ori_n54_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n142_), .B(ori_ori_n77_), .Y(ori_ori_n143_));
  AOI210     o121(.A0(ori_ori_n90_), .A1(ori_ori_n55_), .B0(ori_ori_n38_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n95_), .B(ori_ori_n87_), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n145_), .B(ori_ori_n37_), .Y(ori_ori_n146_));
  OAI210     o124(.A0(ori_ori_n146_), .A1(ori_ori_n144_), .B0(x04), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n77_), .B(ori_ori_n90_), .Y(ori_ori_n148_));
  AN2        o126(.A(x12), .B(ori_ori_n87_), .Y(ori_ori_n149_));
  NO2        o127(.A(ori_ori_n149_), .B(ori_ori_n148_), .Y(ori_ori_n150_));
  NA4        o128(.A(ori_ori_n150_), .B(ori_ori_n147_), .C(ori_ori_n143_), .D(ori_ori_n140_), .Y(ori04));
  NO2        o129(.A(ori_ori_n66_), .B(ori_ori_n39_), .Y(ori_ori_n152_));
  XO2        o130(.A(ori_ori_n152_), .B(ori_ori_n110_), .Y(ori05));
  AOI210     o131(.A0(ori_ori_n172_), .A1(x12), .B0(ori_ori_n26_), .Y(ori_ori_n154_));
  NA2        o132(.A(x12), .B(ori_ori_n79_), .Y(ori_ori_n155_));
  NOi21      o133(.An(ori_ori_n123_), .B(ori_ori_n87_), .Y(ori_ori_n156_));
  NO3        o134(.A(x01), .B(ori_ori_n155_), .C(x08), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n86_), .B(ori_ori_n28_), .Y(ori_ori_n158_));
  NO2        o136(.A(ori_ori_n158_), .B(ori_ori_n114_), .Y(ori_ori_n159_));
  NA3        o137(.A(ori_ori_n127_), .B(ori_ori_n82_), .C(x12), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(x08), .Y(ori_ori_n161_));
  INV        o139(.A(ori_ori_n161_), .Y(ori_ori_n162_));
  NO2        o140(.A(ori_ori_n157_), .B(ori_ori_n162_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n159_), .B(ori_ori_n156_), .Y(ori_ori_n164_));
  NA2        o142(.A(x14), .B(ori_ori_n164_), .Y(ori_ori_n165_));
  OAI210     o143(.A0(x07), .A1(ori_ori_n67_), .B0(x12), .Y(ori_ori_n166_));
  NO4        o144(.A(ori_ori_n166_), .B(ori_ori_n165_), .C(ori_ori_n163_), .D(ori_ori_n154_), .Y(ori06));
  INV        o145(.A(x03), .Y(ori_ori_n170_));
  INV        o146(.A(ori_ori_n93_), .Y(ori_ori_n171_));
  INV        o147(.A(x07), .Y(ori_ori_n172_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NO3        m026(.A(x02), .B(x11), .C(x09), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  NA2        m029(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(x07), .Y(mai_mai_n53_));
  OAI210     m031(.A0(mai_mai_n53_), .A1(mai_mai_n49_), .B0(mai_mai_n47_), .Y(mai_mai_n54_));
  NOi21      m032(.An(x01), .B(x09), .Y(mai_mai_n55_));
  INV        m033(.A(x00), .Y(mai_mai_n56_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n56_), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n57_), .B(mai_mai_n55_), .Y(mai_mai_n58_));
  NA2        m036(.A(x09), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  INV        m037(.A(x07), .Y(mai_mai_n60_));
  AOI220     m038(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n60_), .Y(mai_mai_n61_));
  INV        m039(.A(mai_mai_n58_), .Y(mai_mai_n62_));
  OAI220     m040(.A0(mai_mai_n23_), .A1(mai_mai_n62_), .B0(mai_mai_n61_), .B1(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n60_), .B(mai_mai_n48_), .Y(mai_mai_n64_));
  OAI210     m042(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n64_), .Y(mai_mai_n65_));
  AOI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n58_), .B0(mai_mai_n63_), .B1(mai_mai_n31_), .Y(mai_mai_n66_));
  AOI210     m044(.A0(mai_mai_n66_), .A1(mai_mai_n54_), .B0(x05), .Y(mai_mai_n67_));
  NO2        m045(.A(mai_mai_n60_), .B(mai_mai_n23_), .Y(mai_mai_n68_));
  NA2        m046(.A(x09), .B(x05), .Y(mai_mai_n69_));
  NA2        m047(.A(x10), .B(x06), .Y(mai_mai_n70_));
  NA3        m048(.A(mai_mai_n70_), .B(mai_mai_n69_), .C(mai_mai_n28_), .Y(mai_mai_n71_));
  OAI210     m049(.A0(mai_mai_n71_), .A1(mai_mai_n68_), .B0(x03), .Y(mai_mai_n72_));
  NOi31      m050(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n73_));
  AOI210     m051(.A0(mai_mai_n312_), .A1(mai_mai_n73_), .B0(mai_mai_n24_), .Y(mai_mai_n74_));
  NO2        m052(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n76_));
  NO2        m054(.A(x08), .B(x01), .Y(mai_mai_n77_));
  OAI210     m055(.A0(mai_mai_n77_), .A1(mai_mai_n76_), .B0(mai_mai_n35_), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n78_), .B(mai_mai_n74_), .Y(mai_mai_n79_));
  AN2        m057(.A(mai_mai_n79_), .B(mai_mai_n72_), .Y(mai_mai_n80_));
  INV        m058(.A(mai_mai_n78_), .Y(mai_mai_n81_));
  NO2        m059(.A(x06), .B(x05), .Y(mai_mai_n82_));
  NA2        m060(.A(x11), .B(x00), .Y(mai_mai_n83_));
  NO2        m061(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n84_));
  NOi21      m062(.An(mai_mai_n83_), .B(mai_mai_n84_), .Y(mai_mai_n85_));
  AOI210     m063(.A0(mai_mai_n82_), .A1(mai_mai_n81_), .B0(mai_mai_n85_), .Y(mai_mai_n86_));
  NO2        m064(.A(mai_mai_n52_), .B(x11), .Y(mai_mai_n87_));
  NOi21      m065(.An(x01), .B(x10), .Y(mai_mai_n88_));
  NO2        m066(.A(mai_mai_n29_), .B(mai_mai_n56_), .Y(mai_mai_n89_));
  NO3        m067(.A(mai_mai_n89_), .B(mai_mai_n88_), .C(x06), .Y(mai_mai_n90_));
  AOI220     m068(.A0(mai_mai_n90_), .A1(mai_mai_n27_), .B0(mai_mai_n87_), .B1(mai_mai_n81_), .Y(mai_mai_n91_));
  OAI210     m069(.A0(mai_mai_n86_), .A1(x07), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NO3        m070(.A(mai_mai_n92_), .B(mai_mai_n80_), .C(mai_mai_n67_), .Y(mai01));
  INV        m071(.A(x12), .Y(mai_mai_n94_));
  INV        m072(.A(x13), .Y(mai_mai_n95_));
  NA2        m073(.A(x08), .B(x04), .Y(mai_mai_n96_));
  NA2        m074(.A(mai_mai_n88_), .B(mai_mai_n28_), .Y(mai_mai_n97_));
  NO2        m075(.A(x10), .B(x01), .Y(mai_mai_n98_));
  NO2        m076(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n99_));
  NA2        m077(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n100_));
  NO3        m078(.A(mai_mai_n100_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n55_), .B(x05), .Y(mai_mai_n102_));
  NOi21      m080(.An(mai_mai_n102_), .B(mai_mai_n57_), .Y(mai_mai_n103_));
  NA3        m081(.A(x08), .B(x04), .C(x06), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n104_), .B(mai_mai_n103_), .Y(mai_mai_n105_));
  NO2        m083(.A(x04), .B(x05), .Y(mai_mai_n106_));
  NA2        m084(.A(mai_mai_n35_), .B(mai_mai_n56_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n108_));
  NA2        m086(.A(x10), .B(mai_mai_n56_), .Y(mai_mai_n109_));
  NA2        m087(.A(mai_mai_n109_), .B(mai_mai_n108_), .Y(mai_mai_n110_));
  NA2        m088(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n59_), .B(x05), .Y(mai_mai_n112_));
  NO2        m090(.A(x06), .B(x03), .Y(mai_mai_n113_));
  NO4        m091(.A(mai_mai_n113_), .B(mai_mai_n313_), .C(mai_mai_n105_), .D(mai_mai_n101_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n115_));
  NA2        m093(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n116_));
  NO2        m094(.A(x09), .B(x05), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n117_), .B(mai_mai_n47_), .Y(mai_mai_n118_));
  NA2        m096(.A(x09), .B(x00), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n102_), .B(mai_mai_n119_), .Y(mai_mai_n120_));
  NO2        m098(.A(x03), .B(x02), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n78_), .B(mai_mai_n95_), .Y(mai_mai_n122_));
  INV        m100(.A(mai_mai_n121_), .Y(mai_mai_n123_));
  OA210      m101(.A0(x02), .A1(x11), .B0(mai_mai_n123_), .Y(mai_mai_n124_));
  OAI210     m102(.A0(mai_mai_n114_), .A1(mai_mai_n23_), .B0(mai_mai_n124_), .Y(mai_mai_n125_));
  NAi21      m103(.An(x06), .B(x10), .Y(mai_mai_n126_));
  NOi21      m104(.An(x01), .B(x13), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n128_));
  NO2        m106(.A(mai_mai_n31_), .B(mai_mai_n41_), .Y(mai_mai_n129_));
  NO2        m107(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n95_), .B(x01), .Y(mai_mai_n131_));
  NO2        m109(.A(mai_mai_n131_), .B(x08), .Y(mai_mai_n132_));
  OAI210     m110(.A0(x05), .A1(mai_mai_n132_), .B0(mai_mai_n50_), .Y(mai_mai_n133_));
  AOI210     m111(.A0(mai_mai_n133_), .A1(mai_mai_n130_), .B0(mai_mai_n48_), .Y(mai_mai_n134_));
  AOI210     m112(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n135_));
  OAI210     m113(.A0(mai_mai_n134_), .A1(mai_mai_n129_), .B0(mai_mai_n135_), .Y(mai_mai_n136_));
  NA2        m114(.A(x04), .B(x02), .Y(mai_mai_n137_));
  NA2        m115(.A(x10), .B(x05), .Y(mai_mai_n138_));
  NO2        m116(.A(mai_mai_n102_), .B(x08), .Y(mai_mai_n139_));
  NA3        m117(.A(mai_mai_n127_), .B(mai_mai_n126_), .C(mai_mai_n50_), .Y(mai_mai_n140_));
  INV        m118(.A(mai_mai_n140_), .Y(mai_mai_n141_));
  AOI210     m119(.A0(mai_mai_n139_), .A1(x06), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n142_), .B(x11), .Y(mai_mai_n143_));
  NAi21      m121(.An(mai_mai_n137_), .B(mai_mai_n143_), .Y(mai_mai_n144_));
  INV        m122(.A(mai_mai_n25_), .Y(mai_mai_n145_));
  NAi21      m123(.An(x13), .B(x00), .Y(mai_mai_n146_));
  AOI210     m124(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n146_), .Y(mai_mai_n147_));
  AOI220     m125(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n148_));
  OAI210     m126(.A0(mai_mai_n138_), .A1(mai_mai_n35_), .B0(mai_mai_n148_), .Y(mai_mai_n149_));
  AN2        m127(.A(mai_mai_n149_), .B(mai_mai_n147_), .Y(mai_mai_n150_));
  NO2        m128(.A(mai_mai_n146_), .B(mai_mai_n36_), .Y(mai_mai_n151_));
  INV        m129(.A(mai_mai_n151_), .Y(mai_mai_n152_));
  OAI210     m130(.A0(mai_mai_n151_), .A1(mai_mai_n150_), .B0(mai_mai_n145_), .Y(mai_mai_n153_));
  NA2        m131(.A(x10), .B(x08), .Y(mai_mai_n154_));
  NO2        m132(.A(mai_mai_n95_), .B(x12), .Y(mai_mai_n155_));
  AOI210     m133(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n155_), .Y(mai_mai_n156_));
  NA2        m134(.A(mai_mai_n88_), .B(mai_mai_n50_), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n156_), .B(x12), .Y(mai_mai_n159_));
  NA4        m137(.A(mai_mai_n159_), .B(mai_mai_n153_), .C(mai_mai_n144_), .D(mai_mai_n136_), .Y(mai_mai_n160_));
  AOI210     m138(.A0(mai_mai_n125_), .A1(mai_mai_n94_), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  AOI210     m139(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n162_));
  NO2        m140(.A(mai_mai_n108_), .B(x06), .Y(mai_mai_n163_));
  NO2        m141(.A(mai_mai_n162_), .B(mai_mai_n163_), .Y(mai_mai_n164_));
  AOI210     m142(.A0(mai_mai_n164_), .A1(mai_mai_n71_), .B0(x12), .Y(mai_mai_n165_));
  INV        m143(.A(mai_mai_n73_), .Y(mai_mai_n166_));
  AOI210     m144(.A0(mai_mai_n154_), .A1(x05), .B0(mai_mai_n50_), .Y(mai_mai_n167_));
  OAI210     m145(.A0(mai_mai_n167_), .A1(mai_mai_n128_), .B0(mai_mai_n56_), .Y(mai_mai_n168_));
  NA2        m146(.A(mai_mai_n168_), .B(mai_mai_n166_), .Y(mai_mai_n169_));
  AOI210     m147(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n50_), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n170_), .B(mai_mai_n41_), .Y(mai_mai_n171_));
  NA2        m149(.A(x09), .B(mai_mai_n116_), .Y(mai_mai_n172_));
  OAI210     m150(.A0(mai_mai_n172_), .A1(mai_mai_n171_), .B0(x02), .Y(mai_mai_n173_));
  AOI210     m151(.A0(mai_mai_n173_), .A1(mai_mai_n169_), .B0(mai_mai_n23_), .Y(mai_mai_n174_));
  OAI210     m152(.A0(mai_mai_n165_), .A1(mai_mai_n56_), .B0(mai_mai_n174_), .Y(mai_mai_n175_));
  NO2        m153(.A(mai_mai_n50_), .B(x03), .Y(mai_mai_n176_));
  NO2        m154(.A(mai_mai_n95_), .B(x03), .Y(mai_mai_n177_));
  INV        m155(.A(x05), .Y(mai_mai_n178_));
  INV        m156(.A(mai_mai_n84_), .Y(mai_mai_n179_));
  NO2        m157(.A(mai_mai_n179_), .B(x12), .Y(mai_mai_n180_));
  NA2        m158(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n181_));
  NO2        m159(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n182_));
  OAI210     m160(.A0(mai_mai_n182_), .A1(mai_mai_n149_), .B0(mai_mai_n147_), .Y(mai_mai_n183_));
  AOI210     m161(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n184_), .B(mai_mai_n41_), .Y(mai_mai_n185_));
  OAI210     m163(.A0(mai_mai_n96_), .A1(mai_mai_n119_), .B0(mai_mai_n70_), .Y(mai_mai_n186_));
  NO2        m164(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  NA2        m165(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n188_), .B(x03), .Y(mai_mai_n189_));
  OA210      m167(.A0(mai_mai_n189_), .A1(mai_mai_n187_), .B0(mai_mai_n183_), .Y(mai_mai_n190_));
  NA2        m168(.A(x13), .B(mai_mai_n94_), .Y(mai_mai_n191_));
  NA3        m169(.A(mai_mai_n191_), .B(x12), .C(mai_mai_n85_), .Y(mai_mai_n192_));
  OAI210     m170(.A0(mai_mai_n190_), .A1(mai_mai_n181_), .B0(mai_mai_n192_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n180_), .B(mai_mai_n193_), .Y(mai_mai_n194_));
  AOI210     m172(.A0(mai_mai_n194_), .A1(mai_mai_n175_), .B0(x07), .Y(mai_mai_n195_));
  NO2        m173(.A(x08), .B(x05), .Y(mai_mai_n196_));
  NO2        m174(.A(x12), .B(x02), .Y(mai_mai_n197_));
  INV        m175(.A(mai_mai_n197_), .Y(mai_mai_n198_));
  NO2        m176(.A(mai_mai_n198_), .B(mai_mai_n179_), .Y(mai_mai_n199_));
  NA2        m177(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n200_), .B(x01), .Y(mai_mai_n201_));
  NA2        m179(.A(mai_mai_n95_), .B(x04), .Y(mai_mai_n202_));
  NO3        m180(.A(mai_mai_n83_), .B(x12), .C(x03), .Y(mai_mai_n203_));
  INV        m181(.A(mai_mai_n203_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n157_), .B(mai_mai_n96_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n206_));
  OAI210     m184(.A0(mai_mai_n315_), .A1(mai_mai_n205_), .B0(mai_mai_n206_), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n57_), .B(x05), .Y(mai_mai_n208_));
  NA2        m186(.A(mai_mai_n207_), .B(mai_mai_n204_), .Y(mai_mai_n209_));
  NO3        m187(.A(mai_mai_n209_), .B(mai_mai_n199_), .C(mai_mai_n195_), .Y(mai_mai_n210_));
  OAI210     m188(.A0(mai_mai_n161_), .A1(mai_mai_n60_), .B0(mai_mai_n210_), .Y(mai02));
  INV        m189(.A(mai_mai_n111_), .Y(mai_mai_n212_));
  NA3        m190(.A(x04), .B(x08), .C(mai_mai_n55_), .Y(mai_mai_n213_));
  NA2        m191(.A(mai_mai_n32_), .B(mai_mai_n213_), .Y(mai_mai_n214_));
  OAI210     m192(.A0(mai_mai_n214_), .A1(mai_mai_n212_), .B0(mai_mai_n138_), .Y(mai_mai_n215_));
  INV        m193(.A(mai_mai_n138_), .Y(mai_mai_n216_));
  OAI210     m194(.A0(mai_mai_n78_), .A1(mai_mai_n50_), .B0(mai_mai_n95_), .Y(mai_mai_n217_));
  NA2        m195(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  AOI210     m196(.A0(mai_mai_n218_), .A1(mai_mai_n215_), .B0(mai_mai_n48_), .Y(mai_mai_n219_));
  AOI220     m197(.A0(mai_mai_n196_), .A1(mai_mai_n57_), .B0(mai_mai_n55_), .B1(mai_mai_n36_), .Y(mai_mai_n220_));
  NOi21      m198(.An(x04), .B(mai_mai_n220_), .Y(mai_mai_n221_));
  AOI210     m199(.A0(x13), .A1(mai_mai_n75_), .B0(mai_mai_n221_), .Y(mai_mai_n222_));
  AOI210     m200(.A0(mai_mai_n222_), .A1(x02), .B0(mai_mai_n116_), .Y(mai_mai_n223_));
  NAi21      m201(.An(mai_mai_n178_), .B(x03), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n188_), .B(mai_mai_n47_), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n226_));
  OAI210     m204(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n227_), .Y(mai_mai_n228_));
  OAI210     m206(.A0(mai_mai_n228_), .A1(mai_mai_n177_), .B0(mai_mai_n89_), .Y(mai_mai_n229_));
  NA3        m207(.A(mai_mai_n89_), .B(mai_mai_n77_), .C(mai_mai_n176_), .Y(mai_mai_n230_));
  NA3        m208(.A(mai_mai_n88_), .B(mai_mai_n76_), .C(mai_mai_n42_), .Y(mai_mai_n231_));
  AOI210     m209(.A0(mai_mai_n231_), .A1(mai_mai_n230_), .B0(x04), .Y(mai_mai_n232_));
  INV        m210(.A(mai_mai_n97_), .Y(mai_mai_n233_));
  AOI210     m211(.A0(mai_mai_n233_), .A1(x13), .B0(mai_mai_n232_), .Y(mai_mai_n234_));
  NA3        m212(.A(mai_mai_n234_), .B(mai_mai_n229_), .C(mai_mai_n226_), .Y(mai_mai_n235_));
  NO3        m213(.A(mai_mai_n235_), .B(mai_mai_n223_), .C(mai_mai_n219_), .Y(mai_mai_n236_));
  NA2        m214(.A(mai_mai_n115_), .B(x03), .Y(mai_mai_n237_));
  INV        m215(.A(mai_mai_n146_), .Y(mai_mai_n238_));
  OAI210     m216(.A0(mai_mai_n50_), .A1(mai_mai_n35_), .B0(mai_mai_n36_), .Y(mai_mai_n239_));
  AOI220     m217(.A0(mai_mai_n239_), .A1(mai_mai_n238_), .B0(mai_mai_n158_), .B1(x08), .Y(mai_mai_n240_));
  OAI210     m218(.A0(mai_mai_n240_), .A1(mai_mai_n208_), .B0(mai_mai_n237_), .Y(mai_mai_n241_));
  NA2        m219(.A(mai_mai_n241_), .B(mai_mai_n98_), .Y(mai_mai_n242_));
  NA2        m220(.A(mai_mai_n137_), .B(mai_mai_n131_), .Y(mai_mai_n243_));
  AN2        m221(.A(mai_mai_n243_), .B(mai_mai_n139_), .Y(mai_mai_n244_));
  OAI220     m222(.A0(mai_mai_n202_), .A1(x09), .B0(mai_mai_n111_), .B1(mai_mai_n28_), .Y(mai_mai_n245_));
  OAI210     m223(.A0(mai_mai_n245_), .A1(mai_mai_n244_), .B0(mai_mai_n99_), .Y(mai_mai_n246_));
  NA2        m224(.A(mai_mai_n202_), .B(mai_mai_n94_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n94_), .B(mai_mai_n41_), .Y(mai_mai_n248_));
  NA3        m226(.A(mai_mai_n248_), .B(mai_mai_n247_), .C(mai_mai_n110_), .Y(mai_mai_n249_));
  NA4        m227(.A(mai_mai_n249_), .B(mai_mai_n246_), .C(mai_mai_n242_), .D(mai_mai_n48_), .Y(mai_mai_n250_));
  INV        m228(.A(mai_mai_n158_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n155_), .B(x04), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n252_), .B(mai_mai_n50_), .Y(mai_mai_n253_));
  NO3        m231(.A(mai_mai_n148_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n254_));
  OAI210     m232(.A0(mai_mai_n254_), .A1(mai_mai_n253_), .B0(mai_mai_n89_), .Y(mai_mai_n255_));
  NO3        m233(.A(mai_mai_n155_), .B(mai_mai_n130_), .C(mai_mai_n51_), .Y(mai_mai_n256_));
  OAI210     m234(.A0(mai_mai_n119_), .A1(mai_mai_n36_), .B0(mai_mai_n94_), .Y(mai_mai_n257_));
  NA2        m235(.A(mai_mai_n257_), .B(mai_mai_n256_), .Y(mai_mai_n258_));
  NA3        m236(.A(mai_mai_n258_), .B(mai_mai_n255_), .C(x06), .Y(mai_mai_n259_));
  NO3        m237(.A(mai_mai_n208_), .B(mai_mai_n108_), .C(x08), .Y(mai_mai_n260_));
  INV        m238(.A(mai_mai_n260_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n262_));
  NO3        m240(.A(mai_mai_n102_), .B(mai_mai_n109_), .C(mai_mai_n38_), .Y(mai_mai_n263_));
  AOI210     m241(.A0(mai_mai_n256_), .A1(mai_mai_n262_), .B0(mai_mai_n263_), .Y(mai_mai_n264_));
  OAI210     m242(.A0(mai_mai_n261_), .A1(mai_mai_n28_), .B0(mai_mai_n264_), .Y(mai_mai_n265_));
  AN2        m243(.A(mai_mai_n265_), .B(x04), .Y(mai_mai_n266_));
  AOI210     m244(.A0(mai_mai_n259_), .A1(mai_mai_n250_), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  OAI210     m245(.A0(mai_mai_n236_), .A1(x12), .B0(mai_mai_n267_), .Y(mai03));
  OR2        m246(.A(mai_mai_n42_), .B(mai_mai_n176_), .Y(mai_mai_n269_));
  AOI210     m247(.A0(mai_mai_n122_), .A1(mai_mai_n94_), .B0(mai_mai_n269_), .Y(mai_mai_n270_));
  OAI210     m248(.A0(mai_mai_n314_), .A1(mai_mai_n270_), .B0(x05), .Y(mai_mai_n271_));
  NA2        m249(.A(mai_mai_n269_), .B(x05), .Y(mai_mai_n272_));
  AOI210     m250(.A0(x04), .A1(mai_mai_n166_), .B0(mai_mai_n272_), .Y(mai_mai_n273_));
  AOI210     m251(.A0(mai_mai_n177_), .A1(x08), .B0(mai_mai_n106_), .Y(mai_mai_n274_));
  OAI220     m252(.A0(mai_mai_n274_), .A1(mai_mai_n58_), .B0(x02), .B1(mai_mai_n220_), .Y(mai_mai_n275_));
  OAI210     m253(.A0(mai_mai_n275_), .A1(mai_mai_n273_), .B0(mai_mai_n94_), .Y(mai_mai_n276_));
  AOI210     m254(.A0(mai_mai_n118_), .A1(mai_mai_n59_), .B0(mai_mai_n38_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n120_), .B(x13), .Y(mai_mai_n278_));
  OAI210     m256(.A0(mai_mai_n278_), .A1(mai_mai_n277_), .B0(x04), .Y(mai_mai_n279_));
  NO3        m257(.A(mai_mai_n248_), .B(mai_mai_n78_), .C(mai_mai_n58_), .Y(mai_mai_n280_));
  AOI210     m258(.A0(mai_mai_n152_), .A1(mai_mai_n94_), .B0(mai_mai_n118_), .Y(mai_mai_n281_));
  OA210      m259(.A0(mai_mai_n132_), .A1(x12), .B0(mai_mai_n112_), .Y(mai_mai_n282_));
  NO3        m260(.A(mai_mai_n282_), .B(mai_mai_n281_), .C(mai_mai_n280_), .Y(mai_mai_n283_));
  NA4        m261(.A(mai_mai_n283_), .B(mai_mai_n279_), .C(mai_mai_n276_), .D(mai_mai_n271_), .Y(mai04));
  NO2        m262(.A(mai_mai_n81_), .B(mai_mai_n39_), .Y(mai_mai_n285_));
  XO2        m263(.A(mai_mai_n285_), .B(mai_mai_n191_), .Y(mai05));
  OAI210     m264(.A0(mai_mai_n26_), .A1(mai_mai_n94_), .B0(x07), .Y(mai_mai_n287_));
  INV        m265(.A(mai_mai_n287_), .Y(mai_mai_n288_));
  AOI210     m266(.A0(x12), .A1(mai_mai_n84_), .B0(x07), .Y(mai_mai_n289_));
  NO2        m267(.A(mai_mai_n288_), .B(mai_mai_n289_), .Y(mai_mai_n290_));
  AOI210     m268(.A0(mai_mai_n252_), .A1(mai_mai_n100_), .B0(mai_mai_n197_), .Y(mai_mai_n291_));
  NOi21      m269(.An(mai_mai_n237_), .B(mai_mai_n112_), .Y(mai_mai_n292_));
  OAI210     m270(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n293_));
  AOI210     m271(.A0(mai_mai_n191_), .A1(mai_mai_n47_), .B0(mai_mai_n293_), .Y(mai_mai_n294_));
  NO3        m272(.A(mai_mai_n294_), .B(mai_mai_n291_), .C(x08), .Y(mai_mai_n295_));
  NO2        m273(.A(mai_mai_n111_), .B(mai_mai_n28_), .Y(mai_mai_n296_));
  NO2        m274(.A(mai_mai_n296_), .B(mai_mai_n201_), .Y(mai_mai_n297_));
  NA3        m275(.A(mai_mai_n251_), .B(mai_mai_n107_), .C(x12), .Y(mai_mai_n298_));
  AO210      m276(.A0(mai_mai_n251_), .A1(mai_mai_n107_), .B0(mai_mai_n191_), .Y(mai_mai_n299_));
  NA3        m277(.A(mai_mai_n299_), .B(mai_mai_n298_), .C(x08), .Y(mai_mai_n300_));
  INV        m278(.A(mai_mai_n300_), .Y(mai_mai_n301_));
  NO2        m279(.A(mai_mai_n295_), .B(mai_mai_n301_), .Y(mai_mai_n302_));
  NA3        m280(.A(mai_mai_n297_), .B(mai_mai_n292_), .C(mai_mai_n247_), .Y(mai_mai_n303_));
  NA2        m281(.A(x14), .B(mai_mai_n303_), .Y(mai_mai_n304_));
  NOi21      m282(.An(mai_mai_n202_), .B(mai_mai_n120_), .Y(mai_mai_n305_));
  NO2        m283(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n306_));
  OAI210     m284(.A0(mai_mai_n306_), .A1(mai_mai_n305_), .B0(mai_mai_n94_), .Y(mai_mai_n307_));
  INV        m285(.A(mai_mai_n307_), .Y(mai_mai_n308_));
  NO4        m286(.A(mai_mai_n308_), .B(mai_mai_n304_), .C(mai_mai_n302_), .D(mai_mai_n290_), .Y(mai06));
  INV        m287(.A(x07), .Y(mai_mai_n312_));
  INV        m288(.A(mai_mai_n70_), .Y(mai_mai_n313_));
  INV        m289(.A(mai_mai_n252_), .Y(mai_mai_n314_));
  INV        m290(.A(mai_mai_n69_), .Y(mai_mai_n315_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  OAI210     u030(.A0(men_men_n52_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n53_));
  NOi21      u031(.An(x01), .B(x09), .Y(men_men_n54_));
  INV        u032(.A(x00), .Y(men_men_n55_));
  NO2        u033(.A(men_men_n51_), .B(men_men_n55_), .Y(men_men_n56_));
  NO2        u034(.A(men_men_n56_), .B(men_men_n54_), .Y(men_men_n57_));
  NA2        u035(.A(x09), .B(men_men_n55_), .Y(men_men_n58_));
  INV        u036(.A(x07), .Y(men_men_n59_));
  AOI220     u037(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n59_), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n29_), .B(x02), .Y(men_men_n61_));
  OAI220     u039(.A0(men_men_n29_), .A1(men_men_n56_), .B0(men_men_n60_), .B1(men_men_n58_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n59_), .B(men_men_n48_), .Y(men_men_n63_));
  OAI210     u041(.A0(men_men_n30_), .A1(x11), .B0(men_men_n63_), .Y(men_men_n64_));
  AOI220     u042(.A0(men_men_n64_), .A1(men_men_n57_), .B0(men_men_n62_), .B1(men_men_n31_), .Y(men_men_n65_));
  AOI210     u043(.A0(men_men_n65_), .A1(men_men_n53_), .B0(x05), .Y(men_men_n66_));
  NA2        u044(.A(x10), .B(x09), .Y(men_men_n67_));
  NA2        u045(.A(x09), .B(x05), .Y(men_men_n68_));
  NA2        u046(.A(x10), .B(x06), .Y(men_men_n69_));
  NA3        u047(.A(men_men_n69_), .B(men_men_n68_), .C(men_men_n28_), .Y(men_men_n70_));
  NO2        u048(.A(men_men_n59_), .B(men_men_n41_), .Y(men_men_n71_));
  NA2        u049(.A(men_men_n70_), .B(x03), .Y(men_men_n72_));
  NOi31      u050(.An(x08), .B(x04), .C(x00), .Y(men_men_n73_));
  NO2        u051(.A(x10), .B(x09), .Y(men_men_n74_));
  NO2        u052(.A(x09), .B(men_men_n41_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n75_), .B(men_men_n36_), .Y(men_men_n76_));
  OAI210     u054(.A0(men_men_n75_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n77_));
  AOI210     u055(.A0(men_men_n76_), .A1(men_men_n48_), .B0(men_men_n77_), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n36_), .B(x00), .Y(men_men_n79_));
  NO2        u057(.A(x08), .B(x01), .Y(men_men_n80_));
  OAI210     u058(.A0(men_men_n80_), .A1(men_men_n79_), .B0(men_men_n35_), .Y(men_men_n81_));
  NA2        u059(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n82_));
  NO2        u060(.A(men_men_n81_), .B(men_men_n78_), .Y(men_men_n83_));
  AN2        u061(.A(men_men_n83_), .B(men_men_n72_), .Y(men_men_n84_));
  INV        u062(.A(men_men_n81_), .Y(men_men_n85_));
  NO2        u063(.A(x06), .B(x05), .Y(men_men_n86_));
  NA2        u064(.A(x11), .B(x00), .Y(men_men_n87_));
  NO2        u065(.A(x11), .B(men_men_n47_), .Y(men_men_n88_));
  NOi21      u066(.An(men_men_n87_), .B(men_men_n88_), .Y(men_men_n89_));
  AOI210     u067(.A0(men_men_n86_), .A1(men_men_n85_), .B0(men_men_n89_), .Y(men_men_n90_));
  NOi21      u068(.An(x01), .B(x10), .Y(men_men_n91_));
  NO2        u069(.A(men_men_n29_), .B(men_men_n55_), .Y(men_men_n92_));
  NO3        u070(.A(men_men_n92_), .B(men_men_n91_), .C(x06), .Y(men_men_n93_));
  AOI220     u071(.A0(men_men_n93_), .A1(men_men_n27_), .B0(men_men_n52_), .B1(men_men_n85_), .Y(men_men_n94_));
  OAI210     u072(.A0(men_men_n90_), .A1(x07), .B0(men_men_n94_), .Y(men_men_n95_));
  NO3        u073(.A(men_men_n95_), .B(men_men_n84_), .C(men_men_n66_), .Y(men01));
  INV        u074(.A(x12), .Y(men_men_n97_));
  INV        u075(.A(x13), .Y(men_men_n98_));
  NA2        u076(.A(x08), .B(x04), .Y(men_men_n99_));
  NO2        u077(.A(men_men_n99_), .B(men_men_n55_), .Y(men_men_n100_));
  NA2        u078(.A(men_men_n100_), .B(men_men_n86_), .Y(men_men_n101_));
  NA2        u079(.A(men_men_n91_), .B(men_men_n28_), .Y(men_men_n102_));
  NO2        u080(.A(men_men_n102_), .B(men_men_n68_), .Y(men_men_n103_));
  NO2        u081(.A(x10), .B(x01), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n29_), .B(x00), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n105_), .B(men_men_n104_), .Y(men_men_n106_));
  NA2        u084(.A(x04), .B(men_men_n28_), .Y(men_men_n107_));
  NO3        u085(.A(men_men_n107_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n108_));
  AOI210     u086(.A0(men_men_n108_), .A1(men_men_n106_), .B0(men_men_n103_), .Y(men_men_n109_));
  AOI210     u087(.A0(men_men_n109_), .A1(men_men_n101_), .B0(men_men_n98_), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n54_), .B(x05), .Y(men_men_n111_));
  NOi21      u089(.An(men_men_n111_), .B(men_men_n56_), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n35_), .B(x02), .Y(men_men_n113_));
  NO2        u091(.A(men_men_n98_), .B(men_men_n36_), .Y(men_men_n114_));
  NA3        u092(.A(men_men_n114_), .B(men_men_n113_), .C(x06), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n115_), .B(men_men_n112_), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n80_), .B(x13), .Y(men_men_n117_));
  NA2        u095(.A(x09), .B(men_men_n35_), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n119_));
  NA2        u097(.A(x13), .B(men_men_n35_), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n120_), .B(x05), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n121_), .B(men_men_n119_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n35_), .B(men_men_n55_), .Y(men_men_n123_));
  NA2        u101(.A(men_men_n123_), .B(men_men_n98_), .Y(men_men_n124_));
  AOI210     u102(.A0(men_men_n124_), .A1(men_men_n76_), .B0(men_men_n112_), .Y(men_men_n125_));
  AOI210     u103(.A0(men_men_n125_), .A1(men_men_n122_), .B0(men_men_n69_), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n127_));
  NA2        u105(.A(x10), .B(men_men_n55_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n128_), .B(men_men_n127_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n51_), .B(x05), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n36_), .B(x04), .Y(men_men_n131_));
  NA3        u109(.A(men_men_n131_), .B(men_men_n130_), .C(x13), .Y(men_men_n132_));
  NO3        u110(.A(men_men_n123_), .B(men_men_n75_), .C(men_men_n36_), .Y(men_men_n133_));
  NO2        u111(.A(men_men_n58_), .B(x05), .Y(men_men_n134_));
  NOi41      u112(.An(men_men_n132_), .B(men_men_n134_), .C(men_men_n133_), .D(men_men_n129_), .Y(men_men_n135_));
  NO3        u113(.A(men_men_n135_), .B(x06), .C(x03), .Y(men_men_n136_));
  NO4        u114(.A(men_men_n136_), .B(men_men_n126_), .C(men_men_n116_), .D(men_men_n110_), .Y(men_men_n137_));
  NA2        u115(.A(x13), .B(men_men_n36_), .Y(men_men_n138_));
  OAI210     u116(.A0(men_men_n80_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NOi21      u118(.An(men_men_n86_), .B(men_men_n55_), .Y(men_men_n141_));
  NO2        u119(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n142_));
  OA210      u120(.A0(men_men_n141_), .A1(men_men_n74_), .B0(men_men_n142_), .Y(men_men_n143_));
  NO2        u121(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n144_));
  NA2        u122(.A(men_men_n29_), .B(x06), .Y(men_men_n145_));
  AOI210     u123(.A0(men_men_n145_), .A1(men_men_n49_), .B0(men_men_n144_), .Y(men_men_n146_));
  OA210      u124(.A0(men_men_n146_), .A1(men_men_n143_), .B0(men_men_n140_), .Y(men_men_n147_));
  NO2        u125(.A(x09), .B(x05), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n148_), .B(men_men_n47_), .Y(men_men_n149_));
  AOI210     u127(.A0(men_men_n149_), .A1(men_men_n106_), .B0(men_men_n49_), .Y(men_men_n150_));
  NA2        u128(.A(x09), .B(x00), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n111_), .B(men_men_n151_), .Y(men_men_n152_));
  NA2        u130(.A(men_men_n73_), .B(men_men_n51_), .Y(men_men_n153_));
  AOI210     u131(.A0(men_men_n153_), .A1(men_men_n152_), .B0(men_men_n145_), .Y(men_men_n154_));
  NO3        u132(.A(men_men_n154_), .B(men_men_n150_), .C(men_men_n147_), .Y(men_men_n155_));
  NO2        u133(.A(x03), .B(x02), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n81_), .B(men_men_n98_), .Y(men_men_n157_));
  OAI210     u135(.A0(men_men_n157_), .A1(men_men_n112_), .B0(men_men_n156_), .Y(men_men_n158_));
  OA210      u136(.A0(men_men_n155_), .A1(x11), .B0(men_men_n158_), .Y(men_men_n159_));
  OAI210     u137(.A0(men_men_n137_), .A1(men_men_n23_), .B0(men_men_n159_), .Y(men_men_n160_));
  NA2        u138(.A(men_men_n106_), .B(men_men_n40_), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n162_));
  NAi21      u140(.An(x06), .B(x10), .Y(men_men_n163_));
  NOi21      u141(.An(x01), .B(x13), .Y(men_men_n164_));
  NA2        u142(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  OR2        u143(.A(men_men_n165_), .B(men_men_n162_), .Y(men_men_n166_));
  AOI210     u144(.A0(men_men_n166_), .A1(men_men_n161_), .B0(men_men_n41_), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n29_), .B(x03), .Y(men_men_n168_));
  NA2        u146(.A(men_men_n98_), .B(x01), .Y(men_men_n169_));
  NO2        u147(.A(men_men_n169_), .B(x08), .Y(men_men_n170_));
  OAI210     u148(.A0(x05), .A1(men_men_n170_), .B0(men_men_n51_), .Y(men_men_n171_));
  AOI210     u149(.A0(men_men_n171_), .A1(men_men_n168_), .B0(men_men_n48_), .Y(men_men_n172_));
  AOI210     u150(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n173_));
  OAI210     u151(.A0(men_men_n172_), .A1(men_men_n167_), .B0(men_men_n173_), .Y(men_men_n174_));
  NA2        u152(.A(x04), .B(x02), .Y(men_men_n175_));
  NA2        u153(.A(x10), .B(x05), .Y(men_men_n176_));
  NA2        u154(.A(x09), .B(x06), .Y(men_men_n177_));
  AOI210     u155(.A0(men_men_n177_), .A1(men_men_n176_), .B0(men_men_n162_), .Y(men_men_n178_));
  NO2        u156(.A(x09), .B(x01), .Y(men_men_n179_));
  NO3        u157(.A(men_men_n179_), .B(men_men_n104_), .C(men_men_n31_), .Y(men_men_n180_));
  OAI210     u158(.A0(men_men_n180_), .A1(men_men_n178_), .B0(x00), .Y(men_men_n181_));
  NO2        u159(.A(men_men_n111_), .B(x08), .Y(men_men_n182_));
  NA3        u160(.A(men_men_n164_), .B(men_men_n163_), .C(men_men_n51_), .Y(men_men_n183_));
  NA2        u161(.A(men_men_n91_), .B(x05), .Y(men_men_n184_));
  OAI210     u162(.A0(men_men_n184_), .A1(men_men_n114_), .B0(men_men_n183_), .Y(men_men_n185_));
  AOI210     u163(.A0(men_men_n182_), .A1(x06), .B0(men_men_n185_), .Y(men_men_n186_));
  OAI210     u164(.A0(men_men_n186_), .A1(x11), .B0(men_men_n181_), .Y(men_men_n187_));
  NAi21      u165(.An(men_men_n175_), .B(men_men_n187_), .Y(men_men_n188_));
  INV        u166(.A(men_men_n25_), .Y(men_men_n189_));
  NAi21      u167(.An(x13), .B(x00), .Y(men_men_n190_));
  AOI210     u168(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n190_), .Y(men_men_n191_));
  AOI220     u169(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n192_));
  OAI210     u170(.A0(men_men_n176_), .A1(men_men_n35_), .B0(men_men_n192_), .Y(men_men_n193_));
  AN2        u171(.A(men_men_n193_), .B(men_men_n191_), .Y(men_men_n194_));
  NO2        u172(.A(men_men_n92_), .B(x06), .Y(men_men_n195_));
  NO2        u173(.A(men_men_n190_), .B(men_men_n36_), .Y(men_men_n196_));
  OAI220     u174(.A0(men_men_n190_), .A1(men_men_n177_), .B0(men_men_n195_), .B1(men_men_n68_), .Y(men_men_n197_));
  OAI210     u175(.A0(men_men_n197_), .A1(men_men_n194_), .B0(men_men_n189_), .Y(men_men_n198_));
  NOi21      u176(.An(x09), .B(x00), .Y(men_men_n199_));
  NO3        u177(.A(men_men_n79_), .B(men_men_n199_), .C(men_men_n47_), .Y(men_men_n200_));
  NA2        u178(.A(men_men_n200_), .B(men_men_n128_), .Y(men_men_n201_));
  NA2        u179(.A(x10), .B(x08), .Y(men_men_n202_));
  INV        u180(.A(men_men_n202_), .Y(men_men_n203_));
  NA2        u181(.A(x06), .B(x05), .Y(men_men_n204_));
  OAI210     u182(.A0(men_men_n204_), .A1(men_men_n35_), .B0(men_men_n97_), .Y(men_men_n205_));
  AOI210     u183(.A0(men_men_n203_), .A1(men_men_n56_), .B0(men_men_n205_), .Y(men_men_n206_));
  NA2        u184(.A(men_men_n206_), .B(men_men_n201_), .Y(men_men_n207_));
  NO2        u185(.A(men_men_n98_), .B(x12), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n208_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n91_), .B(men_men_n51_), .Y(men_men_n210_));
  NO2        u188(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n211_), .B(x02), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n212_), .B(men_men_n210_), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n209_), .A1(men_men_n207_), .B0(men_men_n213_), .Y(men_men_n214_));
  NA4        u192(.A(men_men_n214_), .B(men_men_n198_), .C(men_men_n188_), .D(men_men_n174_), .Y(men_men_n215_));
  AOI210     u193(.A0(men_men_n160_), .A1(men_men_n97_), .B0(men_men_n215_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n28_), .B(men_men_n140_), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n218_));
  NA2        u196(.A(men_men_n218_), .B(men_men_n139_), .Y(men_men_n219_));
  AOI210     u197(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n220_));
  NO2        u198(.A(men_men_n127_), .B(x06), .Y(men_men_n221_));
  AOI210     u199(.A0(men_men_n220_), .A1(men_men_n219_), .B0(men_men_n221_), .Y(men_men_n222_));
  AOI210     u200(.A0(men_men_n222_), .A1(men_men_n217_), .B0(x12), .Y(men_men_n223_));
  INV        u201(.A(men_men_n73_), .Y(men_men_n224_));
  AOI210     u202(.A0(men_men_n202_), .A1(x05), .B0(men_men_n51_), .Y(men_men_n225_));
  OAI210     u203(.A0(men_men_n225_), .A1(men_men_n165_), .B0(men_men_n55_), .Y(men_men_n226_));
  NA2        u204(.A(men_men_n226_), .B(men_men_n224_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n91_), .B(x06), .Y(men_men_n228_));
  AOI210     u206(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n229_));
  NO3        u207(.A(men_men_n229_), .B(men_men_n228_), .C(men_men_n41_), .Y(men_men_n230_));
  NA4        u208(.A(men_men_n163_), .B(men_men_n54_), .C(men_men_n36_), .D(x04), .Y(men_men_n231_));
  NA2        u209(.A(men_men_n231_), .B(men_men_n145_), .Y(men_men_n232_));
  OAI210     u210(.A0(men_men_n232_), .A1(men_men_n230_), .B0(x02), .Y(men_men_n233_));
  AOI210     u211(.A0(men_men_n233_), .A1(men_men_n227_), .B0(men_men_n23_), .Y(men_men_n234_));
  OAI210     u212(.A0(men_men_n223_), .A1(men_men_n55_), .B0(men_men_n234_), .Y(men_men_n235_));
  INV        u213(.A(men_men_n145_), .Y(men_men_n236_));
  NO2        u214(.A(men_men_n51_), .B(x03), .Y(men_men_n237_));
  OAI210     u215(.A0(men_men_n75_), .A1(men_men_n36_), .B0(men_men_n118_), .Y(men_men_n238_));
  NO2        u216(.A(men_men_n98_), .B(x03), .Y(men_men_n239_));
  AOI220     u217(.A0(men_men_n239_), .A1(men_men_n238_), .B0(men_men_n73_), .B1(men_men_n237_), .Y(men_men_n240_));
  NA2        u218(.A(men_men_n32_), .B(x06), .Y(men_men_n241_));
  INV        u219(.A(men_men_n163_), .Y(men_men_n242_));
  NOi21      u220(.An(x13), .B(x04), .Y(men_men_n243_));
  NO3        u221(.A(men_men_n243_), .B(men_men_n73_), .C(men_men_n199_), .Y(men_men_n244_));
  NO2        u222(.A(men_men_n244_), .B(x05), .Y(men_men_n245_));
  AOI220     u223(.A0(men_men_n245_), .A1(men_men_n241_), .B0(men_men_n242_), .B1(men_men_n55_), .Y(men_men_n246_));
  OAI210     u224(.A0(men_men_n240_), .A1(men_men_n236_), .B0(men_men_n246_), .Y(men_men_n247_));
  INV        u225(.A(men_men_n88_), .Y(men_men_n248_));
  NA2        u226(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n249_));
  NO2        u227(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n250_));
  OAI210     u228(.A0(men_men_n250_), .A1(men_men_n193_), .B0(men_men_n191_), .Y(men_men_n251_));
  AOI210     u229(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n252_));
  NO2        u230(.A(x06), .B(x00), .Y(men_men_n253_));
  NO3        u231(.A(men_men_n253_), .B(men_men_n252_), .C(men_men_n41_), .Y(men_men_n254_));
  OAI210     u232(.A0(men_men_n99_), .A1(men_men_n151_), .B0(men_men_n69_), .Y(men_men_n255_));
  NO2        u233(.A(men_men_n255_), .B(men_men_n254_), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n257_));
  INV        u235(.A(x03), .Y(men_men_n258_));
  OA210      u236(.A0(men_men_n258_), .A1(men_men_n256_), .B0(men_men_n251_), .Y(men_men_n259_));
  NA2        u237(.A(x13), .B(men_men_n97_), .Y(men_men_n260_));
  NA3        u238(.A(men_men_n260_), .B(men_men_n205_), .C(men_men_n89_), .Y(men_men_n261_));
  OAI210     u239(.A0(men_men_n259_), .A1(men_men_n249_), .B0(men_men_n261_), .Y(men_men_n262_));
  AOI210     u240(.A0(men_men_n88_), .A1(men_men_n247_), .B0(men_men_n262_), .Y(men_men_n263_));
  AOI210     u241(.A0(men_men_n263_), .A1(men_men_n235_), .B0(x07), .Y(men_men_n264_));
  NA2        u242(.A(men_men_n68_), .B(men_men_n29_), .Y(men_men_n265_));
  NOi31      u243(.An(men_men_n138_), .B(men_men_n243_), .C(men_men_n199_), .Y(men_men_n266_));
  AOI210     u244(.A0(men_men_n266_), .A1(men_men_n153_), .B0(men_men_n265_), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n98_), .B(x06), .Y(men_men_n268_));
  INV        u246(.A(men_men_n268_), .Y(men_men_n269_));
  NO2        u247(.A(x08), .B(x05), .Y(men_men_n270_));
  NO2        u248(.A(men_men_n270_), .B(men_men_n252_), .Y(men_men_n271_));
  OAI210     u249(.A0(men_men_n73_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n272_));
  OAI210     u250(.A0(men_men_n271_), .A1(men_men_n269_), .B0(men_men_n272_), .Y(men_men_n273_));
  NO2        u251(.A(x02), .B(men_men_n248_), .Y(men_men_n274_));
  OA210      u252(.A0(men_men_n273_), .A1(men_men_n267_), .B0(men_men_n274_), .Y(men_men_n275_));
  NA2        u253(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n276_));
  NO2        u254(.A(men_men_n276_), .B(x01), .Y(men_men_n277_));
  NOi21      u255(.An(men_men_n80_), .B(men_men_n118_), .Y(men_men_n278_));
  NO2        u256(.A(men_men_n278_), .B(men_men_n277_), .Y(men_men_n279_));
  AOI210     u257(.A0(men_men_n279_), .A1(men_men_n132_), .B0(men_men_n29_), .Y(men_men_n280_));
  NA2        u258(.A(men_men_n268_), .B(men_men_n238_), .Y(men_men_n281_));
  NA2        u259(.A(men_men_n98_), .B(x04), .Y(men_men_n282_));
  NA2        u260(.A(men_men_n282_), .B(men_men_n28_), .Y(men_men_n283_));
  OAI210     u261(.A0(men_men_n283_), .A1(men_men_n117_), .B0(men_men_n281_), .Y(men_men_n284_));
  NO3        u262(.A(men_men_n87_), .B(x12), .C(x03), .Y(men_men_n285_));
  OAI210     u263(.A0(men_men_n284_), .A1(men_men_n280_), .B0(men_men_n285_), .Y(men_men_n286_));
  AOI210     u264(.A0(men_men_n210_), .A1(men_men_n204_), .B0(men_men_n99_), .Y(men_men_n287_));
  NOi21      u265(.An(men_men_n265_), .B(men_men_n228_), .Y(men_men_n288_));
  NO2        u266(.A(men_men_n25_), .B(x00), .Y(men_men_n289_));
  OAI210     u267(.A0(men_men_n288_), .A1(men_men_n287_), .B0(men_men_n289_), .Y(men_men_n290_));
  NO2        u268(.A(men_men_n56_), .B(x05), .Y(men_men_n291_));
  NO3        u269(.A(men_men_n291_), .B(men_men_n229_), .C(men_men_n195_), .Y(men_men_n292_));
  NO2        u270(.A(men_men_n249_), .B(men_men_n28_), .Y(men_men_n293_));
  OAI210     u271(.A0(men_men_n292_), .A1(men_men_n236_), .B0(men_men_n293_), .Y(men_men_n294_));
  NA3        u272(.A(men_men_n294_), .B(men_men_n290_), .C(men_men_n286_), .Y(men_men_n295_));
  NO3        u273(.A(men_men_n295_), .B(men_men_n275_), .C(men_men_n264_), .Y(men_men_n296_));
  OAI210     u274(.A0(men_men_n216_), .A1(men_men_n59_), .B0(men_men_n296_), .Y(men02));
  AOI210     u275(.A0(men_men_n138_), .A1(men_men_n81_), .B0(men_men_n130_), .Y(men_men_n298_));
  NOi21      u276(.An(men_men_n244_), .B(men_men_n179_), .Y(men_men_n299_));
  NA3        u277(.A(x13), .B(men_men_n203_), .C(men_men_n54_), .Y(men_men_n300_));
  OAI210     u278(.A0(men_men_n299_), .A1(men_men_n32_), .B0(men_men_n300_), .Y(men_men_n301_));
  OAI210     u279(.A0(men_men_n301_), .A1(men_men_n298_), .B0(men_men_n176_), .Y(men_men_n302_));
  INV        u280(.A(men_men_n176_), .Y(men_men_n303_));
  AOI210     u281(.A0(men_men_n113_), .A1(men_men_n82_), .B0(men_men_n229_), .Y(men_men_n304_));
  OAI220     u282(.A0(men_men_n304_), .A1(men_men_n98_), .B0(men_men_n81_), .B1(men_men_n51_), .Y(men_men_n305_));
  AOI220     u283(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n157_), .B1(men_men_n156_), .Y(men_men_n306_));
  AOI210     u284(.A0(men_men_n306_), .A1(men_men_n302_), .B0(men_men_n48_), .Y(men_men_n307_));
  NO2        u285(.A(x05), .B(x02), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n219_), .A1(men_men_n199_), .B0(men_men_n308_), .Y(men_men_n309_));
  NOi21      u287(.An(x13), .B(men_men_n454_), .Y(men_men_n310_));
  AOI210     u288(.A0(men_men_n243_), .A1(men_men_n75_), .B0(men_men_n310_), .Y(men_men_n311_));
  AOI210     u289(.A0(men_men_n311_), .A1(men_men_n309_), .B0(men_men_n145_), .Y(men_men_n312_));
  NAi21      u290(.An(men_men_n245_), .B(men_men_n240_), .Y(men_men_n313_));
  NO2        u291(.A(men_men_n257_), .B(men_men_n47_), .Y(men_men_n314_));
  NA2        u292(.A(men_men_n314_), .B(men_men_n313_), .Y(men_men_n315_));
  AN2        u293(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n316_));
  OAI210     u294(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n317_));
  NA2        u295(.A(x13), .B(men_men_n28_), .Y(men_men_n318_));
  OA210      u296(.A0(men_men_n318_), .A1(x08), .B0(men_men_n149_), .Y(men_men_n319_));
  AOI210     u297(.A0(men_men_n319_), .A1(men_men_n139_), .B0(men_men_n317_), .Y(men_men_n320_));
  OAI210     u298(.A0(men_men_n320_), .A1(men_men_n316_), .B0(men_men_n92_), .Y(men_men_n321_));
  NA3        u299(.A(men_men_n92_), .B(men_men_n80_), .C(men_men_n237_), .Y(men_men_n322_));
  NA3        u300(.A(men_men_n91_), .B(men_men_n79_), .C(men_men_n42_), .Y(men_men_n323_));
  AOI210     u301(.A0(men_men_n323_), .A1(men_men_n322_), .B0(x04), .Y(men_men_n324_));
  NO2        u302(.A(men_men_n271_), .B(men_men_n102_), .Y(men_men_n325_));
  AOI210     u303(.A0(men_men_n325_), .A1(x13), .B0(men_men_n324_), .Y(men_men_n326_));
  NA3        u304(.A(men_men_n326_), .B(men_men_n321_), .C(men_men_n315_), .Y(men_men_n327_));
  NO3        u305(.A(men_men_n327_), .B(men_men_n312_), .C(men_men_n307_), .Y(men_men_n328_));
  NA2        u306(.A(men_men_n144_), .B(x03), .Y(men_men_n329_));
  INV        u307(.A(men_men_n190_), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n51_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n331_));
  AOI220     u309(.A0(men_men_n331_), .A1(men_men_n330_), .B0(men_men_n211_), .B1(x08), .Y(men_men_n332_));
  OAI210     u310(.A0(men_men_n332_), .A1(men_men_n291_), .B0(men_men_n329_), .Y(men_men_n333_));
  NA2        u311(.A(men_men_n333_), .B(men_men_n104_), .Y(men_men_n334_));
  NA2        u312(.A(men_men_n175_), .B(men_men_n169_), .Y(men_men_n335_));
  AN2        u313(.A(men_men_n335_), .B(men_men_n182_), .Y(men_men_n336_));
  INV        u314(.A(men_men_n54_), .Y(men_men_n337_));
  OAI220     u315(.A0(men_men_n282_), .A1(men_men_n337_), .B0(men_men_n130_), .B1(men_men_n28_), .Y(men_men_n338_));
  OAI210     u316(.A0(men_men_n338_), .A1(men_men_n336_), .B0(men_men_n105_), .Y(men_men_n339_));
  NA2        u317(.A(men_men_n97_), .B(men_men_n41_), .Y(men_men_n340_));
  NA3        u318(.A(men_men_n340_), .B(x12), .C(men_men_n129_), .Y(men_men_n341_));
  NA4        u319(.A(men_men_n341_), .B(men_men_n339_), .C(men_men_n334_), .D(men_men_n48_), .Y(men_men_n342_));
  INV        u320(.A(men_men_n211_), .Y(men_men_n343_));
  NO2        u321(.A(men_men_n170_), .B(men_men_n40_), .Y(men_men_n344_));
  NA2        u322(.A(men_men_n32_), .B(x05), .Y(men_men_n345_));
  OAI220     u323(.A0(men_men_n345_), .A1(men_men_n344_), .B0(men_men_n343_), .B1(men_men_n57_), .Y(men_men_n346_));
  NA2        u324(.A(men_men_n346_), .B(x02), .Y(men_men_n347_));
  INV        u325(.A(men_men_n250_), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n208_), .B(x04), .Y(men_men_n349_));
  NO2        u327(.A(men_men_n349_), .B(men_men_n348_), .Y(men_men_n350_));
  NO3        u328(.A(men_men_n192_), .B(x13), .C(men_men_n31_), .Y(men_men_n351_));
  OAI210     u329(.A0(men_men_n351_), .A1(men_men_n350_), .B0(men_men_n92_), .Y(men_men_n352_));
  NO3        u330(.A(men_men_n208_), .B(men_men_n168_), .C(men_men_n52_), .Y(men_men_n353_));
  OAI210     u331(.A0(men_men_n151_), .A1(men_men_n36_), .B0(men_men_n97_), .Y(men_men_n354_));
  OAI210     u332(.A0(men_men_n354_), .A1(men_men_n200_), .B0(men_men_n353_), .Y(men_men_n355_));
  NA4        u333(.A(men_men_n355_), .B(men_men_n352_), .C(men_men_n347_), .D(x06), .Y(men_men_n356_));
  NA2        u334(.A(x09), .B(x03), .Y(men_men_n357_));
  OAI220     u335(.A0(men_men_n357_), .A1(men_men_n128_), .B0(men_men_n218_), .B1(men_men_n61_), .Y(men_men_n358_));
  OAI220     u336(.A0(men_men_n169_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n359_));
  NO3        u337(.A(men_men_n291_), .B(men_men_n127_), .C(x08), .Y(men_men_n360_));
  AOI210     u338(.A0(men_men_n359_), .A1(men_men_n236_), .B0(men_men_n360_), .Y(men_men_n361_));
  NO2        u339(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n362_));
  NO3        u340(.A(men_men_n111_), .B(men_men_n128_), .C(men_men_n38_), .Y(men_men_n363_));
  AOI210     u341(.A0(men_men_n353_), .A1(men_men_n362_), .B0(men_men_n363_), .Y(men_men_n364_));
  OAI210     u342(.A0(men_men_n361_), .A1(men_men_n28_), .B0(men_men_n364_), .Y(men_men_n365_));
  AO220      u343(.A0(men_men_n365_), .A1(x04), .B0(men_men_n358_), .B1(x05), .Y(men_men_n366_));
  AOI210     u344(.A0(men_men_n356_), .A1(men_men_n342_), .B0(men_men_n366_), .Y(men_men_n367_));
  OAI210     u345(.A0(men_men_n328_), .A1(x12), .B0(men_men_n367_), .Y(men03));
  OR2        u346(.A(men_men_n42_), .B(men_men_n237_), .Y(men_men_n369_));
  AOI210     u347(.A0(men_men_n157_), .A1(men_men_n97_), .B0(men_men_n369_), .Y(men_men_n370_));
  AO210      u348(.A0(men_men_n348_), .A1(men_men_n82_), .B0(men_men_n349_), .Y(men_men_n371_));
  INV        u349(.A(men_men_n371_), .Y(men_men_n372_));
  OAI210     u350(.A0(men_men_n372_), .A1(men_men_n370_), .B0(x05), .Y(men_men_n373_));
  NA2        u351(.A(men_men_n369_), .B(x05), .Y(men_men_n374_));
  AOI210     u352(.A0(men_men_n139_), .A1(men_men_n224_), .B0(men_men_n374_), .Y(men_men_n375_));
  AOI210     u353(.A0(men_men_n239_), .A1(men_men_n76_), .B0(men_men_n121_), .Y(men_men_n376_));
  OAI220     u354(.A0(men_men_n376_), .A1(men_men_n57_), .B0(men_men_n318_), .B1(men_men_n454_), .Y(men_men_n377_));
  OAI210     u355(.A0(men_men_n377_), .A1(men_men_n375_), .B0(men_men_n97_), .Y(men_men_n378_));
  NO3        u356(.A(men_men_n340_), .B(men_men_n81_), .C(men_men_n57_), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n190_), .A1(men_men_n97_), .B0(men_men_n149_), .Y(men_men_n380_));
  NO3        u358(.A(men_men_n134_), .B(men_men_n380_), .C(men_men_n379_), .Y(men_men_n381_));
  NA4        u359(.A(men_men_n381_), .B(men_men_n152_), .C(men_men_n378_), .D(men_men_n373_), .Y(men04));
  NO2        u360(.A(men_men_n85_), .B(men_men_n39_), .Y(men_men_n383_));
  XO2        u361(.A(men_men_n383_), .B(men_men_n260_), .Y(men05));
  AOI210     u362(.A0(men_men_n68_), .A1(men_men_n52_), .B0(men_men_n221_), .Y(men_men_n385_));
  AOI210     u363(.A0(men_men_n385_), .A1(men_men_n317_), .B0(men_men_n25_), .Y(men_men_n386_));
  NAi41      u364(.An(men_men_n74_), .B(men_men_n145_), .C(men_men_n130_), .D(men_men_n31_), .Y(men_men_n387_));
  AOI210     u365(.A0(men_men_n242_), .A1(men_men_n55_), .B0(men_men_n86_), .Y(men_men_n388_));
  AOI210     u366(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n24_), .Y(men_men_n389_));
  OAI210     u367(.A0(men_men_n389_), .A1(men_men_n386_), .B0(men_men_n97_), .Y(men_men_n390_));
  NA2        u368(.A(x11), .B(men_men_n31_), .Y(men_men_n391_));
  NA2        u369(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n392_));
  NA2        u370(.A(men_men_n265_), .B(x03), .Y(men_men_n393_));
  OAI220     u371(.A0(men_men_n393_), .A1(men_men_n392_), .B0(men_men_n391_), .B1(men_men_n77_), .Y(men_men_n394_));
  AOI210     u372(.A0(men_men_n394_), .A1(x06), .B0(men_men_n455_), .Y(men_men_n395_));
  AOI220     u373(.A0(men_men_n77_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n396_));
  NO3        u374(.A(men_men_n396_), .B(men_men_n23_), .C(x00), .Y(men_men_n397_));
  NA2        u375(.A(men_men_n67_), .B(x02), .Y(men_men_n398_));
  AOI210     u376(.A0(men_men_n398_), .A1(men_men_n393_), .B0(men_men_n268_), .Y(men_men_n399_));
  OR2        u377(.A(men_men_n399_), .B(men_men_n249_), .Y(men_men_n400_));
  NA2        u378(.A(men_men_n164_), .B(x05), .Y(men_men_n401_));
  NA3        u379(.A(men_men_n401_), .B(men_men_n253_), .C(men_men_n248_), .Y(men_men_n402_));
  NO2        u380(.A(men_men_n23_), .B(x10), .Y(men_men_n403_));
  OAI210     u381(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n404_));
  OR3        u382(.A(men_men_n404_), .B(men_men_n403_), .C(men_men_n44_), .Y(men_men_n405_));
  NA3        u383(.A(men_men_n405_), .B(men_men_n402_), .C(men_men_n400_), .Y(men_men_n406_));
  OAI210     u384(.A0(men_men_n406_), .A1(men_men_n397_), .B0(men_men_n97_), .Y(men_men_n407_));
  NA2        u385(.A(men_men_n33_), .B(men_men_n97_), .Y(men_men_n408_));
  AOI210     u386(.A0(men_men_n408_), .A1(men_men_n88_), .B0(x07), .Y(men_men_n409_));
  AOI220     u387(.A0(men_men_n409_), .A1(men_men_n407_), .B0(men_men_n395_), .B1(men_men_n390_), .Y(men_men_n410_));
  NA3        u388(.A(men_men_n23_), .B(men_men_n59_), .C(men_men_n48_), .Y(men_men_n411_));
  AO210      u389(.A0(men_men_n411_), .A1(men_men_n276_), .B0(x02), .Y(men_men_n412_));
  AOI210     u390(.A0(men_men_n403_), .A1(men_men_n71_), .B0(men_men_n144_), .Y(men_men_n413_));
  OR2        u391(.A(men_men_n413_), .B(x03), .Y(men_men_n414_));
  NA2        u392(.A(men_men_n362_), .B(men_men_n59_), .Y(men_men_n415_));
  NO2        u393(.A(men_men_n415_), .B(x11), .Y(men_men_n416_));
  NO3        u394(.A(men_men_n416_), .B(men_men_n148_), .C(men_men_n28_), .Y(men_men_n417_));
  AOI220     u395(.A0(men_men_n417_), .A1(men_men_n414_), .B0(men_men_n412_), .B1(men_men_n47_), .Y(men_men_n418_));
  NO4        u396(.A(men_men_n340_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n419_));
  OAI210     u397(.A0(men_men_n419_), .A1(men_men_n418_), .B0(men_men_n98_), .Y(men_men_n420_));
  NOi21      u398(.An(men_men_n329_), .B(men_men_n134_), .Y(men_men_n421_));
  NO2        u399(.A(men_men_n421_), .B(x02), .Y(men_men_n422_));
  NO2        u400(.A(men_men_n422_), .B(x08), .Y(men_men_n423_));
  AOI210     u401(.A0(men_men_n403_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n424_));
  NA2        u402(.A(x09), .B(men_men_n41_), .Y(men_men_n425_));
  OAI220     u403(.A0(men_men_n425_), .A1(men_men_n424_), .B0(men_men_n391_), .B1(men_men_n63_), .Y(men_men_n426_));
  NO2        u404(.A(x13), .B(x12), .Y(men_men_n427_));
  NO2        u405(.A(men_men_n130_), .B(men_men_n28_), .Y(men_men_n428_));
  NO2        u406(.A(men_men_n428_), .B(men_men_n277_), .Y(men_men_n429_));
  OR3        u407(.A(men_men_n429_), .B(x12), .C(x03), .Y(men_men_n430_));
  NA2        u408(.A(men_men_n430_), .B(x08), .Y(men_men_n431_));
  AOI210     u409(.A0(men_men_n427_), .A1(men_men_n426_), .B0(men_men_n431_), .Y(men_men_n432_));
  AOI210     u410(.A0(men_men_n423_), .A1(men_men_n420_), .B0(men_men_n432_), .Y(men_men_n433_));
  OAI210     u411(.A0(men_men_n415_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n434_));
  NA2        u412(.A(men_men_n303_), .B(x07), .Y(men_men_n435_));
  OAI220     u413(.A0(men_men_n435_), .A1(men_men_n392_), .B0(men_men_n148_), .B1(men_men_n43_), .Y(men_men_n436_));
  OAI210     u414(.A0(men_men_n436_), .A1(men_men_n434_), .B0(men_men_n196_), .Y(men_men_n437_));
  NA3        u415(.A(men_men_n429_), .B(men_men_n421_), .C(x12), .Y(men_men_n438_));
  INV        u416(.A(x14), .Y(men_men_n439_));
  NO3        u417(.A(men_men_n329_), .B(men_men_n102_), .C(x11), .Y(men_men_n440_));
  NO3        u418(.A(men_men_n169_), .B(men_men_n71_), .C(men_men_n55_), .Y(men_men_n441_));
  NO3        u419(.A(men_men_n411_), .B(men_men_n340_), .C(men_men_n190_), .Y(men_men_n442_));
  NO4        u420(.A(men_men_n442_), .B(men_men_n441_), .C(men_men_n440_), .D(men_men_n439_), .Y(men_men_n443_));
  NA3        u421(.A(men_men_n443_), .B(men_men_n438_), .C(men_men_n437_), .Y(men_men_n444_));
  AOI220     u422(.A0(men_men_n408_), .A1(men_men_n59_), .B0(men_men_n428_), .B1(men_men_n168_), .Y(men_men_n445_));
  NO3        u423(.A(men_men_n127_), .B(men_men_n24_), .C(x06), .Y(men_men_n446_));
  AOI210     u424(.A0(men_men_n289_), .A1(men_men_n242_), .B0(men_men_n446_), .Y(men_men_n447_));
  INV        u425(.A(men_men_n447_), .Y(men_men_n448_));
  NA2        u426(.A(men_men_n448_), .B(men_men_n97_), .Y(men_men_n449_));
  OAI210     u427(.A0(men_men_n445_), .A1(men_men_n87_), .B0(men_men_n449_), .Y(men_men_n450_));
  NO4        u428(.A(men_men_n450_), .B(men_men_n444_), .C(men_men_n433_), .D(men_men_n410_), .Y(men06));
  INV        u429(.A(men_men_n270_), .Y(men_men_n454_));
  INV        u430(.A(x07), .Y(men_men_n455_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule