//Benchmark atmr_prom1_2672_0.5

module atmr_prom1(x0, x1, x2, x3, x4, x5, x6, x7, x8, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27, z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27, z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39;
 wire ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1375_, ori_ori_n1376_, ori_ori_n1377_, ori_ori_n1378_, ori_ori_n1379_, ori_ori_n1380_, ori_ori_n1381_, ori_ori_n1382_, ori_ori_n1383_, ori_ori_n1384_, ori_ori_n1385_, ori_ori_n1386_, ori_ori_n1387_, ori_ori_n1388_, ori_ori_n1389_, ori_ori_n1390_, ori_ori_n1391_, ori_ori_n1392_, ori_ori_n1393_, ori_ori_n1395_, ori_ori_n1396_, ori_ori_n1397_, ori_ori_n1398_, ori_ori_n1399_, ori_ori_n1400_, ori_ori_n1401_, ori_ori_n1402_, ori_ori_n1403_, ori_ori_n1404_, ori_ori_n1405_, ori_ori_n1406_, ori_ori_n1407_, ori_ori_n1408_, ori_ori_n1409_, ori_ori_n1410_, ori_ori_n1411_, ori_ori_n1412_, ori_ori_n1413_, ori_ori_n1414_, ori_ori_n1415_, ori_ori_n1416_, ori_ori_n1417_, ori_ori_n1418_, ori_ori_n1419_, ori_ori_n1420_, ori_ori_n1421_, ori_ori_n1422_, ori_ori_n1423_, ori_ori_n1424_, ori_ori_n1425_, ori_ori_n1426_, ori_ori_n1427_, ori_ori_n1428_, ori_ori_n1429_, ori_ori_n1430_, ori_ori_n1431_, ori_ori_n1432_, ori_ori_n1433_, ori_ori_n1434_, ori_ori_n1435_, ori_ori_n1436_, ori_ori_n1437_, ori_ori_n1438_, ori_ori_n1439_, ori_ori_n1440_, ori_ori_n1441_, ori_ori_n1442_, ori_ori_n1443_, ori_ori_n1444_, ori_ori_n1445_, ori_ori_n1446_, ori_ori_n1447_, ori_ori_n1448_, ori_ori_n1449_, ori_ori_n1450_, ori_ori_n1451_, ori_ori_n1452_, ori_ori_n1453_, ori_ori_n1454_, ori_ori_n1455_, ori_ori_n1456_, ori_ori_n1457_, ori_ori_n1458_, ori_ori_n1459_, ori_ori_n1460_, ori_ori_n1461_, ori_ori_n1462_, ori_ori_n1463_, ori_ori_n1465_, ori_ori_n1466_, ori_ori_n1467_, ori_ori_n1468_, ori_ori_n1469_, ori_ori_n1470_, ori_ori_n1471_, ori_ori_n1472_, ori_ori_n1473_, ori_ori_n1474_, ori_ori_n1475_, ori_ori_n1476_, ori_ori_n1477_, ori_ori_n1478_, ori_ori_n1479_, ori_ori_n1480_, ori_ori_n1481_, ori_ori_n1482_, ori_ori_n1483_, ori_ori_n1484_, ori_ori_n1485_, ori_ori_n1486_, ori_ori_n1487_, ori_ori_n1488_, ori_ori_n1489_, ori_ori_n1490_, ori_ori_n1491_, ori_ori_n1492_, ori_ori_n1493_, ori_ori_n1494_, ori_ori_n1495_, ori_ori_n1496_, ori_ori_n1497_, ori_ori_n1498_, ori_ori_n1499_, ori_ori_n1500_, ori_ori_n1501_, ori_ori_n1502_, ori_ori_n1503_, ori_ori_n1504_, ori_ori_n1505_, ori_ori_n1506_, ori_ori_n1507_, ori_ori_n1508_, ori_ori_n1509_, ori_ori_n1510_, ori_ori_n1512_, ori_ori_n1513_, ori_ori_n1514_, ori_ori_n1515_, ori_ori_n1516_, ori_ori_n1517_, ori_ori_n1518_, ori_ori_n1519_, ori_ori_n1520_, ori_ori_n1521_, ori_ori_n1522_, ori_ori_n1523_, ori_ori_n1524_, ori_ori_n1525_, ori_ori_n1526_, ori_ori_n1528_, ori_ori_n1529_, ori_ori_n1530_, ori_ori_n1531_, ori_ori_n1532_, ori_ori_n1533_, ori_ori_n1534_, ori_ori_n1535_, ori_ori_n1536_, ori_ori_n1537_, ori_ori_n1538_, ori_ori_n1540_, ori_ori_n1541_, ori_ori_n1542_, ori_ori_n1543_, ori_ori_n1544_, ori_ori_n1545_, ori_ori_n1546_, ori_ori_n1547_, ori_ori_n1548_, ori_ori_n1549_, ori_ori_n1551_, ori_ori_n1552_, ori_ori_n1553_, ori_ori_n1554_, ori_ori_n1555_, ori_ori_n1556_, ori_ori_n1557_, ori_ori_n1558_, ori_ori_n1559_, ori_ori_n1560_, ori_ori_n1561_, ori_ori_n1562_, ori_ori_n1563_, ori_ori_n1564_, ori_ori_n1565_, ori_ori_n1566_, ori_ori_n1567_, ori_ori_n1568_, ori_ori_n1569_, ori_ori_n1570_, ori_ori_n1571_, ori_ori_n1572_, ori_ori_n1573_, ori_ori_n1574_, ori_ori_n1575_, ori_ori_n1576_, ori_ori_n1577_, ori_ori_n1578_, ori_ori_n1579_, ori_ori_n1580_, ori_ori_n1581_, ori_ori_n1582_, ori_ori_n1583_, ori_ori_n1584_, ori_ori_n1585_, ori_ori_n1586_, ori_ori_n1587_, ori_ori_n1588_, ori_ori_n1589_, ori_ori_n1590_, ori_ori_n1591_, ori_ori_n1592_, ori_ori_n1593_, ori_ori_n1594_, ori_ori_n1596_, ori_ori_n1597_, ori_ori_n1598_, ori_ori_n1599_, ori_ori_n1600_, ori_ori_n1601_, ori_ori_n1602_, ori_ori_n1603_, ori_ori_n1604_, ori_ori_n1605_, ori_ori_n1606_, ori_ori_n1607_, ori_ori_n1608_, ori_ori_n1609_, ori_ori_n1611_, ori_ori_n1612_, ori_ori_n1613_, ori_ori_n1614_, ori_ori_n1615_, ori_ori_n1616_, ori_ori_n1617_, ori_ori_n1618_, ori_ori_n1619_, ori_ori_n1620_, ori_ori_n1621_, ori_ori_n1622_, ori_ori_n1623_, ori_ori_n1624_, ori_ori_n1625_, ori_ori_n1626_, ori_ori_n1627_, ori_ori_n1628_, ori_ori_n1629_, ori_ori_n1630_, ori_ori_n1631_, ori_ori_n1632_, ori_ori_n1633_, ori_ori_n1634_, ori_ori_n1635_, ori_ori_n1636_, ori_ori_n1637_, ori_ori_n1638_, ori_ori_n1639_, ori_ori_n1640_, ori_ori_n1641_, ori_ori_n1642_, ori_ori_n1643_, ori_ori_n1644_, ori_ori_n1645_, ori_ori_n1646_, ori_ori_n1647_, ori_ori_n1648_, ori_ori_n1649_, ori_ori_n1650_, ori_ori_n1651_, ori_ori_n1652_, ori_ori_n1653_, ori_ori_n1655_, ori_ori_n1656_, ori_ori_n1657_, ori_ori_n1658_, ori_ori_n1659_, ori_ori_n1660_, ori_ori_n1661_, ori_ori_n1662_, ori_ori_n1663_, ori_ori_n1664_, ori_ori_n1665_, ori_ori_n1666_, ori_ori_n1667_, ori_ori_n1668_, ori_ori_n1669_, ori_ori_n1670_, ori_ori_n1671_, ori_ori_n1672_, ori_ori_n1673_, ori_ori_n1674_, ori_ori_n1675_, ori_ori_n1676_, ori_ori_n1677_, ori_ori_n1678_, ori_ori_n1679_, ori_ori_n1680_, ori_ori_n1681_, ori_ori_n1682_, ori_ori_n1683_, ori_ori_n1684_, ori_ori_n1685_, ori_ori_n1686_, ori_ori_n1687_, ori_ori_n1688_, ori_ori_n1689_, ori_ori_n1690_, ori_ori_n1691_, ori_ori_n1692_, ori_ori_n1693_, ori_ori_n1694_, ori_ori_n1695_, ori_ori_n1696_, ori_ori_n1697_, ori_ori_n1698_, ori_ori_n1699_, ori_ori_n1700_, ori_ori_n1701_, ori_ori_n1702_, ori_ori_n1703_, ori_ori_n1704_, ori_ori_n1705_, ori_ori_n1706_, ori_ori_n1707_, ori_ori_n1708_, ori_ori_n1710_, ori_ori_n1711_, ori_ori_n1712_, ori_ori_n1713_, ori_ori_n1714_, ori_ori_n1715_, ori_ori_n1716_, ori_ori_n1717_, ori_ori_n1718_, ori_ori_n1719_, ori_ori_n1720_, ori_ori_n1721_, ori_ori_n1722_, ori_ori_n1723_, ori_ori_n1724_, ori_ori_n1725_, ori_ori_n1726_, ori_ori_n1727_, ori_ori_n1728_, ori_ori_n1729_, ori_ori_n1730_, ori_ori_n1731_, ori_ori_n1732_, ori_ori_n1733_, ori_ori_n1734_, ori_ori_n1735_, ori_ori_n1736_, ori_ori_n1737_, ori_ori_n1738_, ori_ori_n1739_, ori_ori_n1740_, ori_ori_n1741_, ori_ori_n1742_, ori_ori_n1743_, ori_ori_n1744_, ori_ori_n1745_, ori_ori_n1746_, ori_ori_n1747_, ori_ori_n1748_, ori_ori_n1749_, ori_ori_n1750_, ori_ori_n1751_, ori_ori_n1752_, ori_ori_n1753_, ori_ori_n1754_, ori_ori_n1755_, ori_ori_n1756_, ori_ori_n1757_, ori_ori_n1758_, ori_ori_n1759_, ori_ori_n1760_, ori_ori_n1761_, ori_ori_n1762_, ori_ori_n1763_, ori_ori_n1764_, ori_ori_n1765_, ori_ori_n1766_, ori_ori_n1767_, ori_ori_n1769_, ori_ori_n1770_, ori_ori_n1771_, ori_ori_n1772_, ori_ori_n1773_, ori_ori_n1774_, ori_ori_n1775_, ori_ori_n1776_, ori_ori_n1777_, ori_ori_n1778_, ori_ori_n1779_, ori_ori_n1780_, ori_ori_n1781_, ori_ori_n1782_, ori_ori_n1783_, ori_ori_n1784_, ori_ori_n1785_, ori_ori_n1786_, ori_ori_n1787_, ori_ori_n1788_, ori_ori_n1789_, ori_ori_n1790_, ori_ori_n1791_, ori_ori_n1792_, ori_ori_n1793_, ori_ori_n1794_, ori_ori_n1795_, ori_ori_n1796_, ori_ori_n1797_, ori_ori_n1798_, ori_ori_n1799_, ori_ori_n1800_, ori_ori_n1801_, ori_ori_n1802_, ori_ori_n1803_, ori_ori_n1804_, ori_ori_n1805_, ori_ori_n1806_, ori_ori_n1807_, ori_ori_n1808_, ori_ori_n1809_, ori_ori_n1810_, ori_ori_n1811_, ori_ori_n1812_, ori_ori_n1813_, ori_ori_n1814_, ori_ori_n1815_, ori_ori_n1816_, ori_ori_n1817_, ori_ori_n1818_, ori_ori_n1819_, ori_ori_n1820_, ori_ori_n1821_, ori_ori_n1822_, ori_ori_n1823_, ori_ori_n1824_, ori_ori_n1825_, ori_ori_n1827_, ori_ori_n1828_, ori_ori_n1829_, ori_ori_n1830_, ori_ori_n1831_, ori_ori_n1832_, ori_ori_n1833_, ori_ori_n1834_, ori_ori_n1835_, ori_ori_n1836_, ori_ori_n1837_, ori_ori_n1838_, ori_ori_n1839_, ori_ori_n1840_, ori_ori_n1841_, ori_ori_n1842_, ori_ori_n1843_, ori_ori_n1844_, ori_ori_n1845_, ori_ori_n1846_, ori_ori_n1847_, ori_ori_n1848_, ori_ori_n1849_, ori_ori_n1850_, ori_ori_n1851_, ori_ori_n1852_, ori_ori_n1853_, ori_ori_n1854_, ori_ori_n1855_, ori_ori_n1856_, ori_ori_n1857_, ori_ori_n1858_, ori_ori_n1859_, ori_ori_n1860_, ori_ori_n1861_, ori_ori_n1862_, ori_ori_n1863_, ori_ori_n1864_, ori_ori_n1865_, ori_ori_n1866_, ori_ori_n1867_, ori_ori_n1868_, ori_ori_n1869_, ori_ori_n1870_, ori_ori_n1871_, ori_ori_n1872_, ori_ori_n1873_, ori_ori_n1874_, ori_ori_n1875_, ori_ori_n1876_, ori_ori_n1877_, ori_ori_n1878_, ori_ori_n1879_, ori_ori_n1880_, ori_ori_n1881_, ori_ori_n1882_, ori_ori_n1883_, ori_ori_n1884_, ori_ori_n1885_, ori_ori_n1886_, ori_ori_n1887_, ori_ori_n1888_, ori_ori_n1889_, ori_ori_n1890_, ori_ori_n1891_, ori_ori_n1892_, ori_ori_n1894_, ori_ori_n1895_, ori_ori_n1896_, ori_ori_n1897_, ori_ori_n1898_, ori_ori_n1899_, ori_ori_n1900_, ori_ori_n1901_, ori_ori_n1902_, ori_ori_n1903_, ori_ori_n1904_, ori_ori_n1905_, ori_ori_n1906_, ori_ori_n1907_, ori_ori_n1908_, ori_ori_n1909_, ori_ori_n1910_, ori_ori_n1911_, ori_ori_n1912_, ori_ori_n1913_, ori_ori_n1914_, ori_ori_n1915_, ori_ori_n1916_, ori_ori_n1917_, ori_ori_n1918_, ori_ori_n1919_, ori_ori_n1920_, ori_ori_n1921_, ori_ori_n1922_, ori_ori_n1923_, ori_ori_n1924_, ori_ori_n1925_, ori_ori_n1926_, ori_ori_n1927_, ori_ori_n1928_, ori_ori_n1929_, ori_ori_n1930_, ori_ori_n1931_, ori_ori_n1932_, ori_ori_n1933_, ori_ori_n1934_, ori_ori_n1935_, ori_ori_n1936_, ori_ori_n1937_, ori_ori_n1938_, ori_ori_n1940_, ori_ori_n1941_, ori_ori_n1942_, ori_ori_n1943_, ori_ori_n1944_, ori_ori_n1945_, ori_ori_n1946_, ori_ori_n1947_, ori_ori_n1948_, ori_ori_n1949_, ori_ori_n1950_, ori_ori_n1951_, ori_ori_n1952_, ori_ori_n1953_, ori_ori_n1954_, ori_ori_n1955_, ori_ori_n1956_, ori_ori_n1957_, ori_ori_n1958_, ori_ori_n1959_, ori_ori_n1960_, ori_ori_n1961_, ori_ori_n1962_, ori_ori_n1963_, ori_ori_n1964_, ori_ori_n1965_, ori_ori_n1966_, ori_ori_n1967_, ori_ori_n1968_, ori_ori_n1969_, ori_ori_n1970_, ori_ori_n1971_, ori_ori_n1972_, ori_ori_n1973_, ori_ori_n1974_, ori_ori_n1975_, ori_ori_n1976_, ori_ori_n1977_, ori_ori_n1978_, ori_ori_n1979_, ori_ori_n1980_, ori_ori_n1981_, ori_ori_n1982_, ori_ori_n1983_, ori_ori_n1984_, ori_ori_n1985_, ori_ori_n1986_, ori_ori_n1987_, ori_ori_n1988_, ori_ori_n1989_, ori_ori_n1991_, ori_ori_n1992_, ori_ori_n1993_, ori_ori_n1994_, ori_ori_n1995_, ori_ori_n1996_, ori_ori_n1997_, ori_ori_n1998_, ori_ori_n1999_, ori_ori_n2000_, ori_ori_n2001_, ori_ori_n2002_, ori_ori_n2003_, ori_ori_n2004_, ori_ori_n2005_, ori_ori_n2006_, ori_ori_n2007_, ori_ori_n2008_, ori_ori_n2009_, ori_ori_n2010_, ori_ori_n2011_, ori_ori_n2012_, ori_ori_n2013_, ori_ori_n2014_, ori_ori_n2015_, ori_ori_n2016_, ori_ori_n2017_, ori_ori_n2018_, ori_ori_n2019_, ori_ori_n2020_, ori_ori_n2021_, ori_ori_n2022_, ori_ori_n2023_, ori_ori_n2024_, ori_ori_n2025_, ori_ori_n2026_, ori_ori_n2027_, ori_ori_n2028_, ori_ori_n2029_, ori_ori_n2030_, ori_ori_n2031_, ori_ori_n2032_, ori_ori_n2033_, ori_ori_n2034_, ori_ori_n2035_, ori_ori_n2036_, ori_ori_n2037_, ori_ori_n2038_, ori_ori_n2039_, ori_ori_n2040_, ori_ori_n2041_, ori_ori_n2042_, ori_ori_n2043_, ori_ori_n2045_, ori_ori_n2046_, ori_ori_n2047_, ori_ori_n2048_, ori_ori_n2049_, ori_ori_n2050_, ori_ori_n2051_, ori_ori_n2052_, ori_ori_n2053_, ori_ori_n2054_, ori_ori_n2055_, ori_ori_n2056_, ori_ori_n2057_, ori_ori_n2058_, ori_ori_n2059_, ori_ori_n2060_, ori_ori_n2061_, ori_ori_n2062_, ori_ori_n2063_, ori_ori_n2064_, ori_ori_n2065_, ori_ori_n2066_, ori_ori_n2067_, ori_ori_n2068_, ori_ori_n2069_, ori_ori_n2070_, ori_ori_n2071_, ori_ori_n2072_, ori_ori_n2073_, ori_ori_n2074_, ori_ori_n2075_, ori_ori_n2076_, ori_ori_n2077_, ori_ori_n2078_, ori_ori_n2080_, ori_ori_n2081_, ori_ori_n2082_, ori_ori_n2083_, ori_ori_n2084_, ori_ori_n2085_, ori_ori_n2086_, ori_ori_n2087_, ori_ori_n2088_, ori_ori_n2089_, ori_ori_n2090_, ori_ori_n2091_, ori_ori_n2092_, ori_ori_n2093_, ori_ori_n2094_, ori_ori_n2095_, ori_ori_n2096_, ori_ori_n2097_, ori_ori_n2098_, ori_ori_n2099_, ori_ori_n2100_, ori_ori_n2101_, ori_ori_n2102_, ori_ori_n2103_, ori_ori_n2104_, ori_ori_n2105_, ori_ori_n2106_, ori_ori_n2107_, ori_ori_n2108_, ori_ori_n2109_, ori_ori_n2110_, ori_ori_n2111_, ori_ori_n2112_, ori_ori_n2113_, ori_ori_n2114_, ori_ori_n2115_, ori_ori_n2116_, ori_ori_n2117_, ori_ori_n2118_, ori_ori_n2119_, ori_ori_n2120_, ori_ori_n2121_, ori_ori_n2122_, ori_ori_n2124_, ori_ori_n2125_, ori_ori_n2126_, ori_ori_n2127_, ori_ori_n2128_, ori_ori_n2129_, ori_ori_n2130_, ori_ori_n2131_, ori_ori_n2132_, ori_ori_n2133_, ori_ori_n2134_, ori_ori_n2135_, ori_ori_n2136_, ori_ori_n2137_, ori_ori_n2138_, ori_ori_n2139_, ori_ori_n2140_, ori_ori_n2141_, ori_ori_n2142_, ori_ori_n2143_, ori_ori_n2144_, ori_ori_n2145_, ori_ori_n2146_, ori_ori_n2147_, ori_ori_n2148_, ori_ori_n2149_, ori_ori_n2150_, ori_ori_n2151_, ori_ori_n2152_, ori_ori_n2153_, ori_ori_n2154_, ori_ori_n2155_, ori_ori_n2156_, ori_ori_n2157_, ori_ori_n2158_, ori_ori_n2159_, ori_ori_n2160_, ori_ori_n2164_, ori_ori_n2165_, ori_ori_n2166_, ori_ori_n2167_, ori_ori_n2168_, ori_ori_n2169_, ori_ori_n2170_, ori_ori_n2171_, ori_ori_n2172_, ori_ori_n2173_, ori_ori_n2174_, ori_ori_n2175_, ori_ori_n2176_, ori_ori_n2177_, ori_ori_n2178_, ori_ori_n2179_, ori_ori_n2180_, ori_ori_n2181_, ori_ori_n2182_, ori_ori_n2183_, ori_ori_n2184_, ori_ori_n2185_, ori_ori_n2186_, ori_ori_n2187_, ori_ori_n2188_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1533_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1543_, mai_mai_n1544_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1549_, mai_mai_n1550_, mai_mai_n1551_, mai_mai_n1552_, mai_mai_n1553_, mai_mai_n1554_, mai_mai_n1555_, mai_mai_n1556_, mai_mai_n1557_, mai_mai_n1558_, mai_mai_n1560_, mai_mai_n1561_, mai_mai_n1562_, mai_mai_n1563_, mai_mai_n1564_, mai_mai_n1565_, mai_mai_n1567_, mai_mai_n1568_, mai_mai_n1569_, mai_mai_n1570_, mai_mai_n1571_, mai_mai_n1572_, mai_mai_n1573_, mai_mai_n1574_, mai_mai_n1575_, mai_mai_n1576_, mai_mai_n1578_, mai_mai_n1579_, mai_mai_n1580_, mai_mai_n1581_, mai_mai_n1582_, mai_mai_n1583_, mai_mai_n1584_, mai_mai_n1585_, mai_mai_n1586_, mai_mai_n1587_, mai_mai_n1588_, mai_mai_n1589_, mai_mai_n1590_, mai_mai_n1591_, mai_mai_n1592_, mai_mai_n1593_, mai_mai_n1594_, mai_mai_n1595_, mai_mai_n1596_, mai_mai_n1597_, mai_mai_n1598_, mai_mai_n1599_, mai_mai_n1600_, mai_mai_n1601_, mai_mai_n1602_, mai_mai_n1603_, mai_mai_n1604_, mai_mai_n1605_, mai_mai_n1607_, mai_mai_n1608_, mai_mai_n1609_, mai_mai_n1610_, mai_mai_n1611_, mai_mai_n1612_, mai_mai_n1613_, mai_mai_n1614_, mai_mai_n1615_, mai_mai_n1616_, mai_mai_n1617_, mai_mai_n1618_, mai_mai_n1619_, mai_mai_n1621_, mai_mai_n1622_, mai_mai_n1623_, mai_mai_n1624_, mai_mai_n1625_, mai_mai_n1626_, mai_mai_n1627_, mai_mai_n1628_, mai_mai_n1629_, mai_mai_n1630_, mai_mai_n1631_, mai_mai_n1632_, mai_mai_n1633_, mai_mai_n1634_, mai_mai_n1635_, mai_mai_n1636_, mai_mai_n1637_, mai_mai_n1638_, mai_mai_n1639_, mai_mai_n1640_, mai_mai_n1641_, mai_mai_n1642_, mai_mai_n1643_, mai_mai_n1644_, mai_mai_n1645_, mai_mai_n1646_, mai_mai_n1647_, mai_mai_n1648_, mai_mai_n1649_, mai_mai_n1650_, mai_mai_n1651_, mai_mai_n1652_, mai_mai_n1654_, mai_mai_n1655_, mai_mai_n1656_, mai_mai_n1657_, mai_mai_n1658_, mai_mai_n1659_, mai_mai_n1660_, mai_mai_n1661_, mai_mai_n1662_, mai_mai_n1663_, mai_mai_n1664_, mai_mai_n1665_, mai_mai_n1666_, mai_mai_n1667_, mai_mai_n1668_, mai_mai_n1669_, mai_mai_n1670_, mai_mai_n1671_, mai_mai_n1672_, mai_mai_n1673_, mai_mai_n1674_, mai_mai_n1675_, mai_mai_n1676_, mai_mai_n1677_, mai_mai_n1678_, mai_mai_n1679_, mai_mai_n1680_, mai_mai_n1681_, mai_mai_n1682_, mai_mai_n1683_, mai_mai_n1684_, mai_mai_n1685_, mai_mai_n1686_, mai_mai_n1687_, mai_mai_n1688_, mai_mai_n1689_, mai_mai_n1690_, mai_mai_n1691_, mai_mai_n1692_, mai_mai_n1693_, mai_mai_n1694_, mai_mai_n1695_, mai_mai_n1696_, mai_mai_n1697_, mai_mai_n1698_, mai_mai_n1699_, mai_mai_n1700_, mai_mai_n1701_, mai_mai_n1702_, mai_mai_n1703_, mai_mai_n1704_, mai_mai_n1706_, mai_mai_n1707_, mai_mai_n1708_, mai_mai_n1709_, mai_mai_n1710_, mai_mai_n1711_, mai_mai_n1712_, mai_mai_n1713_, mai_mai_n1714_, mai_mai_n1715_, mai_mai_n1716_, mai_mai_n1717_, mai_mai_n1718_, mai_mai_n1719_, mai_mai_n1720_, mai_mai_n1721_, mai_mai_n1722_, mai_mai_n1723_, mai_mai_n1724_, mai_mai_n1725_, mai_mai_n1726_, mai_mai_n1727_, mai_mai_n1728_, mai_mai_n1729_, mai_mai_n1730_, mai_mai_n1731_, mai_mai_n1732_, mai_mai_n1733_, mai_mai_n1734_, mai_mai_n1735_, mai_mai_n1736_, mai_mai_n1737_, mai_mai_n1738_, mai_mai_n1739_, mai_mai_n1740_, mai_mai_n1741_, mai_mai_n1742_, mai_mai_n1743_, mai_mai_n1744_, mai_mai_n1745_, mai_mai_n1746_, mai_mai_n1747_, mai_mai_n1748_, mai_mai_n1749_, mai_mai_n1750_, mai_mai_n1751_, mai_mai_n1752_, mai_mai_n1753_, mai_mai_n1754_, mai_mai_n1755_, mai_mai_n1756_, mai_mai_n1757_, mai_mai_n1758_, mai_mai_n1759_, mai_mai_n1760_, mai_mai_n1761_, mai_mai_n1762_, mai_mai_n1763_, mai_mai_n1764_, mai_mai_n1765_, mai_mai_n1766_, mai_mai_n1767_, mai_mai_n1768_, mai_mai_n1769_, mai_mai_n1770_, mai_mai_n1771_, mai_mai_n1772_, mai_mai_n1773_, mai_mai_n1775_, mai_mai_n1776_, mai_mai_n1777_, mai_mai_n1778_, mai_mai_n1779_, mai_mai_n1780_, mai_mai_n1781_, mai_mai_n1782_, mai_mai_n1783_, mai_mai_n1784_, mai_mai_n1785_, mai_mai_n1786_, mai_mai_n1787_, mai_mai_n1788_, mai_mai_n1789_, mai_mai_n1790_, mai_mai_n1791_, mai_mai_n1792_, mai_mai_n1793_, mai_mai_n1794_, mai_mai_n1795_, mai_mai_n1796_, mai_mai_n1797_, mai_mai_n1798_, mai_mai_n1799_, mai_mai_n1800_, mai_mai_n1801_, mai_mai_n1802_, mai_mai_n1803_, mai_mai_n1804_, mai_mai_n1805_, mai_mai_n1806_, mai_mai_n1807_, mai_mai_n1808_, mai_mai_n1809_, mai_mai_n1810_, mai_mai_n1811_, mai_mai_n1812_, mai_mai_n1813_, mai_mai_n1814_, mai_mai_n1815_, mai_mai_n1816_, mai_mai_n1817_, mai_mai_n1818_, mai_mai_n1819_, mai_mai_n1820_, mai_mai_n1821_, mai_mai_n1822_, mai_mai_n1823_, mai_mai_n1824_, mai_mai_n1825_, mai_mai_n1826_, mai_mai_n1827_, mai_mai_n1828_, mai_mai_n1829_, mai_mai_n1830_, mai_mai_n1831_, mai_mai_n1832_, mai_mai_n1833_, mai_mai_n1834_, mai_mai_n1836_, mai_mai_n1837_, mai_mai_n1838_, mai_mai_n1839_, mai_mai_n1840_, mai_mai_n1841_, mai_mai_n1842_, mai_mai_n1843_, mai_mai_n1844_, mai_mai_n1845_, mai_mai_n1846_, mai_mai_n1847_, mai_mai_n1848_, mai_mai_n1849_, mai_mai_n1850_, mai_mai_n1851_, mai_mai_n1852_, mai_mai_n1853_, mai_mai_n1854_, mai_mai_n1855_, mai_mai_n1856_, mai_mai_n1857_, mai_mai_n1858_, mai_mai_n1859_, mai_mai_n1860_, mai_mai_n1861_, mai_mai_n1862_, mai_mai_n1863_, mai_mai_n1864_, mai_mai_n1865_, mai_mai_n1866_, mai_mai_n1867_, mai_mai_n1868_, mai_mai_n1869_, mai_mai_n1870_, mai_mai_n1871_, mai_mai_n1872_, mai_mai_n1873_, mai_mai_n1874_, mai_mai_n1875_, mai_mai_n1876_, mai_mai_n1877_, mai_mai_n1878_, mai_mai_n1879_, mai_mai_n1880_, mai_mai_n1881_, mai_mai_n1882_, mai_mai_n1883_, mai_mai_n1884_, mai_mai_n1885_, mai_mai_n1886_, mai_mai_n1887_, mai_mai_n1888_, mai_mai_n1889_, mai_mai_n1890_, mai_mai_n1891_, mai_mai_n1892_, mai_mai_n1893_, mai_mai_n1894_, mai_mai_n1896_, mai_mai_n1897_, mai_mai_n1898_, mai_mai_n1899_, mai_mai_n1900_, mai_mai_n1901_, mai_mai_n1902_, mai_mai_n1903_, mai_mai_n1904_, mai_mai_n1905_, mai_mai_n1906_, mai_mai_n1907_, mai_mai_n1908_, mai_mai_n1909_, mai_mai_n1910_, mai_mai_n1911_, mai_mai_n1912_, mai_mai_n1913_, mai_mai_n1914_, mai_mai_n1915_, mai_mai_n1916_, mai_mai_n1917_, mai_mai_n1918_, mai_mai_n1919_, mai_mai_n1920_, mai_mai_n1921_, mai_mai_n1922_, mai_mai_n1923_, mai_mai_n1924_, mai_mai_n1925_, mai_mai_n1926_, mai_mai_n1927_, mai_mai_n1928_, mai_mai_n1929_, mai_mai_n1930_, mai_mai_n1931_, mai_mai_n1932_, mai_mai_n1933_, mai_mai_n1934_, mai_mai_n1935_, mai_mai_n1936_, mai_mai_n1937_, mai_mai_n1938_, mai_mai_n1939_, mai_mai_n1940_, mai_mai_n1941_, mai_mai_n1942_, mai_mai_n1943_, mai_mai_n1944_, mai_mai_n1945_, mai_mai_n1946_, mai_mai_n1948_, mai_mai_n1949_, mai_mai_n1950_, mai_mai_n1951_, mai_mai_n1952_, mai_mai_n1953_, mai_mai_n1954_, mai_mai_n1955_, mai_mai_n1956_, mai_mai_n1957_, mai_mai_n1958_, mai_mai_n1959_, mai_mai_n1960_, mai_mai_n1961_, mai_mai_n1962_, mai_mai_n1963_, mai_mai_n1964_, mai_mai_n1965_, mai_mai_n1966_, mai_mai_n1967_, mai_mai_n1968_, mai_mai_n1969_, mai_mai_n1970_, mai_mai_n1971_, mai_mai_n1972_, mai_mai_n1973_, mai_mai_n1974_, mai_mai_n1975_, mai_mai_n1976_, mai_mai_n1977_, mai_mai_n1978_, mai_mai_n1979_, mai_mai_n1980_, mai_mai_n1981_, mai_mai_n1982_, mai_mai_n1983_, mai_mai_n1984_, mai_mai_n1985_, mai_mai_n1986_, mai_mai_n1987_, mai_mai_n1988_, mai_mai_n1989_, mai_mai_n1990_, mai_mai_n1991_, mai_mai_n1992_, mai_mai_n1993_, mai_mai_n1994_, mai_mai_n1996_, mai_mai_n1997_, mai_mai_n1998_, mai_mai_n1999_, mai_mai_n2000_, mai_mai_n2001_, mai_mai_n2002_, mai_mai_n2003_, mai_mai_n2004_, mai_mai_n2005_, mai_mai_n2006_, mai_mai_n2007_, mai_mai_n2008_, mai_mai_n2009_, mai_mai_n2010_, mai_mai_n2011_, mai_mai_n2012_, mai_mai_n2013_, mai_mai_n2014_, mai_mai_n2015_, mai_mai_n2016_, mai_mai_n2017_, mai_mai_n2018_, mai_mai_n2019_, mai_mai_n2020_, mai_mai_n2021_, mai_mai_n2022_, mai_mai_n2023_, mai_mai_n2024_, mai_mai_n2025_, mai_mai_n2026_, mai_mai_n2027_, mai_mai_n2028_, mai_mai_n2029_, mai_mai_n2030_, mai_mai_n2031_, mai_mai_n2032_, mai_mai_n2033_, mai_mai_n2034_, mai_mai_n2035_, mai_mai_n2036_, mai_mai_n2037_, mai_mai_n2038_, mai_mai_n2039_, mai_mai_n2040_, mai_mai_n2041_, mai_mai_n2042_, mai_mai_n2043_, mai_mai_n2044_, mai_mai_n2045_, mai_mai_n2046_, mai_mai_n2047_, mai_mai_n2048_, mai_mai_n2049_, mai_mai_n2050_, mai_mai_n2051_, mai_mai_n2052_, mai_mai_n2053_, mai_mai_n2054_, mai_mai_n2056_, mai_mai_n2057_, mai_mai_n2058_, mai_mai_n2059_, mai_mai_n2060_, mai_mai_n2061_, mai_mai_n2062_, mai_mai_n2063_, mai_mai_n2064_, mai_mai_n2065_, mai_mai_n2066_, mai_mai_n2067_, mai_mai_n2068_, mai_mai_n2069_, mai_mai_n2070_, mai_mai_n2071_, mai_mai_n2072_, mai_mai_n2073_, mai_mai_n2074_, mai_mai_n2075_, mai_mai_n2076_, mai_mai_n2077_, mai_mai_n2078_, mai_mai_n2079_, mai_mai_n2080_, mai_mai_n2081_, mai_mai_n2082_, mai_mai_n2083_, mai_mai_n2084_, mai_mai_n2085_, mai_mai_n2086_, mai_mai_n2087_, mai_mai_n2088_, mai_mai_n2089_, mai_mai_n2090_, mai_mai_n2091_, mai_mai_n2092_, mai_mai_n2093_, mai_mai_n2094_, mai_mai_n2095_, mai_mai_n2096_, mai_mai_n2097_, mai_mai_n2098_, mai_mai_n2099_, mai_mai_n2100_, mai_mai_n2101_, mai_mai_n2102_, mai_mai_n2103_, mai_mai_n2104_, mai_mai_n2105_, mai_mai_n2107_, mai_mai_n2108_, mai_mai_n2109_, mai_mai_n2110_, mai_mai_n2111_, mai_mai_n2112_, mai_mai_n2113_, mai_mai_n2114_, mai_mai_n2115_, mai_mai_n2116_, mai_mai_n2117_, mai_mai_n2118_, mai_mai_n2119_, mai_mai_n2120_, mai_mai_n2121_, mai_mai_n2122_, mai_mai_n2123_, mai_mai_n2124_, mai_mai_n2125_, mai_mai_n2126_, mai_mai_n2127_, mai_mai_n2128_, mai_mai_n2129_, mai_mai_n2130_, mai_mai_n2131_, mai_mai_n2132_, mai_mai_n2133_, mai_mai_n2134_, mai_mai_n2135_, mai_mai_n2136_, mai_mai_n2137_, mai_mai_n2138_, mai_mai_n2139_, mai_mai_n2140_, mai_mai_n2141_, mai_mai_n2142_, mai_mai_n2143_, mai_mai_n2144_, mai_mai_n2145_, mai_mai_n2146_, mai_mai_n2147_, mai_mai_n2148_, mai_mai_n2149_, mai_mai_n2150_, mai_mai_n2151_, mai_mai_n2152_, mai_mai_n2153_, mai_mai_n2154_, mai_mai_n2155_, mai_mai_n2156_, mai_mai_n2158_, mai_mai_n2159_, mai_mai_n2160_, mai_mai_n2161_, mai_mai_n2162_, mai_mai_n2163_, mai_mai_n2164_, mai_mai_n2165_, mai_mai_n2166_, mai_mai_n2167_, mai_mai_n2168_, mai_mai_n2169_, mai_mai_n2170_, mai_mai_n2171_, mai_mai_n2172_, mai_mai_n2173_, mai_mai_n2174_, mai_mai_n2175_, mai_mai_n2176_, mai_mai_n2177_, mai_mai_n2178_, mai_mai_n2179_, mai_mai_n2180_, mai_mai_n2181_, mai_mai_n2182_, mai_mai_n2183_, mai_mai_n2184_, mai_mai_n2185_, mai_mai_n2186_, mai_mai_n2187_, mai_mai_n2188_, mai_mai_n2189_, mai_mai_n2190_, mai_mai_n2191_, mai_mai_n2192_, mai_mai_n2193_, mai_mai_n2194_, mai_mai_n2195_, mai_mai_n2196_, mai_mai_n2197_, mai_mai_n2198_, mai_mai_n2199_, mai_mai_n2200_, mai_mai_n2201_, mai_mai_n2202_, mai_mai_n2203_, mai_mai_n2204_, mai_mai_n2205_, mai_mai_n2206_, mai_mai_n2207_, mai_mai_n2208_, mai_mai_n2209_, mai_mai_n2210_, mai_mai_n2211_, mai_mai_n2212_, mai_mai_n2216_, mai_mai_n2217_, mai_mai_n2218_, mai_mai_n2219_, mai_mai_n2220_, mai_mai_n2221_, mai_mai_n2222_, mai_mai_n2223_, mai_mai_n2224_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1606_, men_men_n1607_, men_men_n1608_, men_men_n1609_, men_men_n1610_, men_men_n1611_, men_men_n1612_, men_men_n1613_, men_men_n1615_, men_men_n1616_, men_men_n1617_, men_men_n1618_, men_men_n1619_, men_men_n1620_, men_men_n1621_, men_men_n1622_, men_men_n1623_, men_men_n1624_, men_men_n1625_, men_men_n1626_, men_men_n1627_, men_men_n1628_, men_men_n1629_, men_men_n1630_, men_men_n1631_, men_men_n1632_, men_men_n1633_, men_men_n1634_, men_men_n1635_, men_men_n1636_, men_men_n1637_, men_men_n1638_, men_men_n1639_, men_men_n1640_, men_men_n1641_, men_men_n1642_, men_men_n1643_, men_men_n1644_, men_men_n1645_, men_men_n1646_, men_men_n1647_, men_men_n1648_, men_men_n1649_, men_men_n1650_, men_men_n1651_, men_men_n1652_, men_men_n1653_, men_men_n1654_, men_men_n1655_, men_men_n1657_, men_men_n1658_, men_men_n1659_, men_men_n1660_, men_men_n1661_, men_men_n1662_, men_men_n1663_, men_men_n1664_, men_men_n1665_, men_men_n1666_, men_men_n1667_, men_men_n1669_, men_men_n1670_, men_men_n1671_, men_men_n1672_, men_men_n1673_, men_men_n1674_, men_men_n1675_, men_men_n1676_, men_men_n1677_, men_men_n1678_, men_men_n1679_, men_men_n1680_, men_men_n1681_, men_men_n1682_, men_men_n1683_, men_men_n1684_, men_men_n1685_, men_men_n1686_, men_men_n1687_, men_men_n1688_, men_men_n1689_, men_men_n1690_, men_men_n1691_, men_men_n1692_, men_men_n1693_, men_men_n1694_, men_men_n1695_, men_men_n1696_, men_men_n1697_, men_men_n1698_, men_men_n1699_, men_men_n1700_, men_men_n1701_, men_men_n1702_, men_men_n1703_, men_men_n1704_, men_men_n1705_, men_men_n1706_, men_men_n1707_, men_men_n1708_, men_men_n1709_, men_men_n1710_, men_men_n1711_, men_men_n1712_, men_men_n1713_, men_men_n1714_, men_men_n1715_, men_men_n1716_, men_men_n1718_, men_men_n1719_, men_men_n1720_, men_men_n1721_, men_men_n1722_, men_men_n1723_, men_men_n1724_, men_men_n1725_, men_men_n1726_, men_men_n1727_, men_men_n1728_, men_men_n1729_, men_men_n1730_, men_men_n1731_, men_men_n1732_, men_men_n1733_, men_men_n1734_, men_men_n1735_, men_men_n1736_, men_men_n1737_, men_men_n1738_, men_men_n1739_, men_men_n1740_, men_men_n1741_, men_men_n1742_, men_men_n1743_, men_men_n1744_, men_men_n1745_, men_men_n1746_, men_men_n1747_, men_men_n1748_, men_men_n1749_, men_men_n1750_, men_men_n1751_, men_men_n1752_, men_men_n1753_, men_men_n1754_, men_men_n1755_, men_men_n1756_, men_men_n1757_, men_men_n1758_, men_men_n1759_, men_men_n1760_, men_men_n1761_, men_men_n1762_, men_men_n1763_, men_men_n1764_, men_men_n1765_, men_men_n1766_, men_men_n1767_, men_men_n1768_, men_men_n1769_, men_men_n1770_, men_men_n1772_, men_men_n1773_, men_men_n1774_, men_men_n1775_, men_men_n1776_, men_men_n1777_, men_men_n1778_, men_men_n1779_, men_men_n1780_, men_men_n1781_, men_men_n1782_, men_men_n1783_, men_men_n1784_, men_men_n1785_, men_men_n1786_, men_men_n1787_, men_men_n1788_, men_men_n1789_, men_men_n1790_, men_men_n1791_, men_men_n1792_, men_men_n1793_, men_men_n1794_, men_men_n1795_, men_men_n1796_, men_men_n1797_, men_men_n1798_, men_men_n1799_, men_men_n1800_, men_men_n1801_, men_men_n1802_, men_men_n1803_, men_men_n1804_, men_men_n1805_, men_men_n1806_, men_men_n1807_, men_men_n1808_, men_men_n1809_, men_men_n1810_, men_men_n1811_, men_men_n1812_, men_men_n1813_, men_men_n1814_, men_men_n1815_, men_men_n1816_, men_men_n1817_, men_men_n1818_, men_men_n1819_, men_men_n1820_, men_men_n1821_, men_men_n1822_, men_men_n1823_, men_men_n1824_, men_men_n1825_, men_men_n1826_, men_men_n1827_, men_men_n1828_, men_men_n1829_, men_men_n1831_, men_men_n1832_, men_men_n1833_, men_men_n1834_, men_men_n1835_, men_men_n1836_, men_men_n1837_, men_men_n1838_, men_men_n1839_, men_men_n1840_, men_men_n1841_, men_men_n1842_, men_men_n1843_, men_men_n1844_, men_men_n1845_, men_men_n1846_, men_men_n1847_, men_men_n1848_, men_men_n1849_, men_men_n1850_, men_men_n1851_, men_men_n1852_, men_men_n1853_, men_men_n1854_, men_men_n1855_, men_men_n1856_, men_men_n1857_, men_men_n1858_, men_men_n1859_, men_men_n1860_, men_men_n1861_, men_men_n1862_, men_men_n1863_, men_men_n1864_, men_men_n1865_, men_men_n1866_, men_men_n1867_, men_men_n1868_, men_men_n1869_, men_men_n1870_, men_men_n1871_, men_men_n1872_, men_men_n1873_, men_men_n1874_, men_men_n1875_, men_men_n1876_, men_men_n1877_, men_men_n1878_, men_men_n1879_, men_men_n1880_, men_men_n1881_, men_men_n1882_, men_men_n1883_, men_men_n1884_, men_men_n1885_, men_men_n1886_, men_men_n1887_, men_men_n1888_, men_men_n1890_, men_men_n1891_, men_men_n1892_, men_men_n1893_, men_men_n1894_, men_men_n1895_, men_men_n1896_, men_men_n1897_, men_men_n1898_, men_men_n1899_, men_men_n1900_, men_men_n1901_, men_men_n1902_, men_men_n1903_, men_men_n1904_, men_men_n1905_, men_men_n1906_, men_men_n1907_, men_men_n1908_, men_men_n1909_, men_men_n1910_, men_men_n1911_, men_men_n1912_, men_men_n1913_, men_men_n1914_, men_men_n1915_, men_men_n1916_, men_men_n1917_, men_men_n1918_, men_men_n1919_, men_men_n1920_, men_men_n1921_, men_men_n1922_, men_men_n1923_, men_men_n1924_, men_men_n1925_, men_men_n1926_, men_men_n1927_, men_men_n1928_, men_men_n1929_, men_men_n1930_, men_men_n1931_, men_men_n1932_, men_men_n1933_, men_men_n1934_, men_men_n1935_, men_men_n1936_, men_men_n1937_, men_men_n1938_, men_men_n1939_, men_men_n1940_, men_men_n1941_, men_men_n1942_, men_men_n1943_, men_men_n1944_, men_men_n1945_, men_men_n1946_, men_men_n1947_, men_men_n1948_, men_men_n1949_, men_men_n1950_, men_men_n1951_, men_men_n1952_, men_men_n1954_, men_men_n1955_, men_men_n1956_, men_men_n1957_, men_men_n1958_, men_men_n1959_, men_men_n1960_, men_men_n1961_, men_men_n1962_, men_men_n1963_, men_men_n1964_, men_men_n1965_, men_men_n1966_, men_men_n1967_, men_men_n1968_, men_men_n1969_, men_men_n1970_, men_men_n1971_, men_men_n1972_, men_men_n1973_, men_men_n1974_, men_men_n1975_, men_men_n1976_, men_men_n1977_, men_men_n1978_, men_men_n1979_, men_men_n1980_, men_men_n1981_, men_men_n1982_, men_men_n1983_, men_men_n1984_, men_men_n1985_, men_men_n1986_, men_men_n1987_, men_men_n1988_, men_men_n1989_, men_men_n1990_, men_men_n1991_, men_men_n1992_, men_men_n1993_, men_men_n1994_, men_men_n1995_, men_men_n1996_, men_men_n1997_, men_men_n1998_, men_men_n1999_, men_men_n2000_, men_men_n2001_, men_men_n2002_, men_men_n2003_, men_men_n2004_, men_men_n2005_, men_men_n2006_, men_men_n2007_, men_men_n2008_, men_men_n2009_, men_men_n2010_, men_men_n2011_, men_men_n2012_, men_men_n2013_, men_men_n2015_, men_men_n2016_, men_men_n2017_, men_men_n2018_, men_men_n2019_, men_men_n2020_, men_men_n2021_, men_men_n2022_, men_men_n2023_, men_men_n2024_, men_men_n2025_, men_men_n2026_, men_men_n2027_, men_men_n2028_, men_men_n2029_, men_men_n2030_, men_men_n2031_, men_men_n2032_, men_men_n2033_, men_men_n2034_, men_men_n2035_, men_men_n2036_, men_men_n2037_, men_men_n2038_, men_men_n2039_, men_men_n2040_, men_men_n2041_, men_men_n2042_, men_men_n2043_, men_men_n2044_, men_men_n2045_, men_men_n2046_, men_men_n2047_, men_men_n2048_, men_men_n2049_, men_men_n2050_, men_men_n2051_, men_men_n2052_, men_men_n2053_, men_men_n2054_, men_men_n2055_, men_men_n2056_, men_men_n2057_, men_men_n2058_, men_men_n2059_, men_men_n2060_, men_men_n2061_, men_men_n2062_, men_men_n2063_, men_men_n2064_, men_men_n2065_, men_men_n2067_, men_men_n2068_, men_men_n2069_, men_men_n2070_, men_men_n2071_, men_men_n2072_, men_men_n2073_, men_men_n2074_, men_men_n2075_, men_men_n2076_, men_men_n2077_, men_men_n2078_, men_men_n2079_, men_men_n2080_, men_men_n2081_, men_men_n2082_, men_men_n2083_, men_men_n2084_, men_men_n2085_, men_men_n2086_, men_men_n2087_, men_men_n2088_, men_men_n2089_, men_men_n2090_, men_men_n2091_, men_men_n2092_, men_men_n2093_, men_men_n2094_, men_men_n2095_, men_men_n2096_, men_men_n2097_, men_men_n2098_, men_men_n2099_, men_men_n2100_, men_men_n2101_, men_men_n2102_, men_men_n2103_, men_men_n2104_, men_men_n2105_, men_men_n2106_, men_men_n2107_, men_men_n2108_, men_men_n2109_, men_men_n2110_, men_men_n2111_, men_men_n2112_, men_men_n2113_, men_men_n2114_, men_men_n2115_, men_men_n2116_, men_men_n2117_, men_men_n2118_, men_men_n2119_, men_men_n2120_, men_men_n2121_, men_men_n2122_, men_men_n2123_, men_men_n2124_, men_men_n2125_, men_men_n2126_, men_men_n2127_, men_men_n2129_, men_men_n2130_, men_men_n2131_, men_men_n2132_, men_men_n2133_, men_men_n2134_, men_men_n2135_, men_men_n2136_, men_men_n2137_, men_men_n2138_, men_men_n2139_, men_men_n2140_, men_men_n2141_, men_men_n2142_, men_men_n2143_, men_men_n2144_, men_men_n2145_, men_men_n2146_, men_men_n2147_, men_men_n2148_, men_men_n2149_, men_men_n2150_, men_men_n2151_, men_men_n2152_, men_men_n2153_, men_men_n2154_, men_men_n2155_, men_men_n2156_, men_men_n2157_, men_men_n2158_, men_men_n2159_, men_men_n2160_, men_men_n2161_, men_men_n2162_, men_men_n2163_, men_men_n2164_, men_men_n2165_, men_men_n2166_, men_men_n2167_, men_men_n2168_, men_men_n2169_, men_men_n2170_, men_men_n2171_, men_men_n2172_, men_men_n2173_, men_men_n2174_, men_men_n2175_, men_men_n2176_, men_men_n2177_, men_men_n2178_, men_men_n2179_, men_men_n2180_, men_men_n2181_, men_men_n2182_, men_men_n2183_, men_men_n2184_, men_men_n2185_, men_men_n2187_, men_men_n2188_, men_men_n2189_, men_men_n2190_, men_men_n2191_, men_men_n2192_, men_men_n2193_, men_men_n2194_, men_men_n2195_, men_men_n2196_, men_men_n2197_, men_men_n2198_, men_men_n2199_, men_men_n2200_, men_men_n2201_, men_men_n2202_, men_men_n2203_, men_men_n2204_, men_men_n2205_, men_men_n2206_, men_men_n2207_, men_men_n2208_, men_men_n2209_, men_men_n2210_, men_men_n2211_, men_men_n2212_, men_men_n2213_, men_men_n2214_, men_men_n2215_, men_men_n2216_, men_men_n2217_, men_men_n2218_, men_men_n2219_, men_men_n2220_, men_men_n2221_, men_men_n2222_, men_men_n2223_, men_men_n2224_, men_men_n2225_, men_men_n2226_, men_men_n2227_, men_men_n2228_, men_men_n2229_, men_men_n2230_, men_men_n2231_, men_men_n2232_, men_men_n2233_, men_men_n2234_, men_men_n2235_, men_men_n2236_, men_men_n2237_, men_men_n2238_, men_men_n2239_, men_men_n2240_, men_men_n2241_, men_men_n2242_, men_men_n2243_, men_men_n2244_, men_men_n2245_, men_men_n2247_, men_men_n2248_, men_men_n2249_, men_men_n2250_, men_men_n2251_, men_men_n2252_, men_men_n2253_, men_men_n2254_, men_men_n2255_, men_men_n2256_, men_men_n2257_, men_men_n2258_, men_men_n2259_, men_men_n2260_, men_men_n2261_, men_men_n2262_, men_men_n2263_, men_men_n2264_, men_men_n2265_, men_men_n2266_, men_men_n2267_, men_men_n2268_, men_men_n2269_, men_men_n2270_, men_men_n2271_, men_men_n2272_, men_men_n2273_, men_men_n2274_, men_men_n2275_, men_men_n2276_, men_men_n2277_, men_men_n2278_, men_men_n2279_, men_men_n2280_, men_men_n2281_, men_men_n2282_, men_men_n2283_, men_men_n2284_, men_men_n2285_, men_men_n2286_, men_men_n2287_, men_men_n2288_, men_men_n2289_, men_men_n2290_, men_men_n2291_, men_men_n2292_, men_men_n2293_, men_men_n2294_, men_men_n2295_, men_men_n2296_, men_men_n2297_, men_men_n2298_, men_men_n2299_, men_men_n2300_, men_men_n2301_, men_men_n2302_, men_men_n2303_, men_men_n2304_, men_men_n2308_, men_men_n2309_, men_men_n2310_, men_men_n2311_, men_men_n2312_, men_men_n2313_, men_men_n2314_, men_men_n2315_, men_men_n2316_, men_men_n2317_, men_men_n2318_, men_men_n2319_, men_men_n2320_, men_men_n2321_, men_men_n2322_, men_men_n2323_, men_men_n2324_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13, ori14, mai14, men14, ori15, mai15, men15, ori16, mai16, men16, ori17, mai17, men17, ori18, mai18, men18, ori19, mai19, men19, ori20, mai20, men20, ori21, mai21, men21, ori22, mai22, men22, ori23, mai23, men23, ori24, mai24, men24, ori25, mai25, men25, ori26, mai26, men26, ori27, mai27, men27, ori28, mai28, men28, ori29, mai29, men29, ori30, mai30, men30, ori31, mai31, men31, ori32, mai32, men32, ori33, mai33, men33, ori34, mai34, men34, ori35, mai35, men35, ori36, mai36, men36, ori37, mai37, men37, ori38, mai38, men38, ori39, mai39, men39;
  INV        o0000(.A(x3), .Y(ori_ori_n50_));
  NA2        o0001(.A(ori_ori_n50_), .B(x2), .Y(ori_ori_n51_));
  NA2        o0002(.A(x7), .B(x0), .Y(ori_ori_n52_));
  INV        o0003(.A(x1), .Y(ori_ori_n53_));
  NA2        o0004(.A(x5), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  INV        o0005(.A(x8), .Y(ori_ori_n55_));
  INV        o0006(.A(x4), .Y(ori_ori_n56_));
  INV        o0007(.A(x0), .Y(ori_ori_n57_));
  NA2        o0008(.A(x4), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NA3        o0009(.A(ori_ori_n58_), .B(ori_ori_n55_), .C(x6), .Y(ori_ori_n59_));
  NA2        o0010(.A(ori_ori_n56_), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  NO2        o0011(.A(ori_ori_n55_), .B(x6), .Y(ori_ori_n61_));
  NA2        o0012(.A(ori_ori_n61_), .B(ori_ori_n60_), .Y(ori_ori_n62_));
  AOI210     o0013(.A0(ori_ori_n62_), .A1(ori_ori_n59_), .B0(ori_ori_n54_), .Y(ori_ori_n63_));
  INV        o0014(.A(x8), .Y(ori_ori_n64_));
  NO2        o0015(.A(x7), .B(ori_ori_n57_), .Y(ori_ori_n65_));
  NO2        o0016(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  NAi21      o0017(.An(x5), .B(x1), .Y(ori_ori_n67_));
  INV        o0018(.A(x6), .Y(ori_ori_n68_));
  NA2        o0019(.A(ori_ori_n68_), .B(x4), .Y(ori_ori_n69_));
  NO3        o0020(.A(ori_ori_n69_), .B(ori_ori_n67_), .C(ori_ori_n66_), .Y(ori_ori_n70_));
  OAI210     o0021(.A0(ori_ori_n70_), .A1(ori_ori_n63_), .B0(ori_ori_n52_), .Y(ori_ori_n71_));
  NA2        o0022(.A(x7), .B(x4), .Y(ori_ori_n72_));
  NO2        o0023(.A(ori_ori_n72_), .B(x1), .Y(ori_ori_n73_));
  NO2        o0024(.A(ori_ori_n68_), .B(x5), .Y(ori_ori_n74_));
  NO2        o0025(.A(x8), .B(ori_ori_n57_), .Y(ori_ori_n75_));
  NA3        o0026(.A(ori_ori_n75_), .B(ori_ori_n74_), .C(ori_ori_n73_), .Y(ori_ori_n76_));
  AOI210     o0027(.A0(ori_ori_n76_), .A1(ori_ori_n71_), .B0(ori_ori_n51_), .Y(ori_ori_n77_));
  NA2        o0028(.A(x5), .B(x3), .Y(ori_ori_n78_));
  NO2        o0029(.A(x6), .B(x0), .Y(ori_ori_n79_));
  NO2        o0030(.A(ori_ori_n79_), .B(x4), .Y(ori_ori_n80_));
  NO2        o0031(.A(x4), .B(x2), .Y(ori_ori_n81_));
  NO2        o0032(.A(ori_ori_n68_), .B(ori_ori_n57_), .Y(ori_ori_n82_));
  NA2        o0033(.A(x8), .B(x1), .Y(ori_ori_n83_));
  NO2        o0034(.A(x8), .B(x6), .Y(ori_ori_n84_));
  NO2        o0035(.A(x1), .B(ori_ori_n57_), .Y(ori_ori_n85_));
  NO2        o0036(.A(ori_ori_n56_), .B(x2), .Y(ori_ori_n86_));
  XO2        o0037(.A(x7), .B(x1), .Y(ori_ori_n87_));
  INV        o0038(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  NO2        o0039(.A(ori_ori_n88_), .B(x6), .Y(ori_ori_n89_));
  NO2        o0040(.A(ori_ori_n50_), .B(x0), .Y(ori_ori_n90_));
  NA2        o0041(.A(ori_ori_n90_), .B(ori_ori_n55_), .Y(ori_ori_n91_));
  NO2        o0042(.A(x6), .B(x5), .Y(ori_ori_n92_));
  INV        o0043(.A(x5), .Y(ori_ori_n93_));
  NA2        o0044(.A(x6), .B(x1), .Y(ori_ori_n94_));
  NA2        o0045(.A(ori_ori_n94_), .B(ori_ori_n81_), .Y(ori_ori_n95_));
  NO4        o0046(.A(ori_ori_n95_), .B(x5), .C(ori_ori_n91_), .D(ori_ori_n89_), .Y(ori_ori_n96_));
  NA2        o0047(.A(x3), .B(x0), .Y(ori_ori_n97_));
  INV        o0048(.A(x5), .Y(ori_ori_n98_));
  NA2        o0049(.A(ori_ori_n68_), .B(ori_ori_n98_), .Y(ori_ori_n99_));
  INV        o0050(.A(x2), .Y(ori_ori_n100_));
  NO2        o0051(.A(ori_ori_n56_), .B(ori_ori_n100_), .Y(ori_ori_n101_));
  NA2        o0052(.A(ori_ori_n101_), .B(ori_ori_n99_), .Y(ori_ori_n102_));
  NO3        o0053(.A(ori_ori_n102_), .B(ori_ori_n97_), .C(ori_ori_n53_), .Y(ori_ori_n103_));
  NO3        o0054(.A(ori_ori_n103_), .B(ori_ori_n96_), .C(ori_ori_n77_), .Y(ori00));
  NO2        o0055(.A(x7), .B(x6), .Y(ori_ori_n105_));
  INV        o0056(.A(ori_ori_n105_), .Y(ori_ori_n106_));
  NO2        o0057(.A(ori_ori_n55_), .B(ori_ori_n53_), .Y(ori_ori_n107_));
  NA2        o0058(.A(ori_ori_n107_), .B(ori_ori_n56_), .Y(ori_ori_n108_));
  XN2        o0059(.A(x6), .B(x1), .Y(ori_ori_n109_));
  INV        o0060(.A(ori_ori_n109_), .Y(ori_ori_n110_));
  NO2        o0061(.A(x6), .B(x4), .Y(ori_ori_n111_));
  NA2        o0062(.A(x6), .B(x4), .Y(ori_ori_n112_));
  NAi21      o0063(.An(ori_ori_n111_), .B(ori_ori_n112_), .Y(ori_ori_n113_));
  XN2        o0064(.A(x7), .B(x6), .Y(ori_ori_n114_));
  NO4        o0065(.A(ori_ori_n114_), .B(ori_ori_n113_), .C(ori_ori_n110_), .D(x8), .Y(ori_ori_n115_));
  NO2        o0066(.A(x3), .B(ori_ori_n100_), .Y(ori_ori_n116_));
  NA2        o0067(.A(ori_ori_n116_), .B(ori_ori_n98_), .Y(ori_ori_n117_));
  NO2        o0068(.A(ori_ori_n117_), .B(ori_ori_n57_), .Y(ori_ori_n118_));
  OAI210     o0069(.A0(ori_ori_n115_), .A1(ori_ori_n105_), .B0(ori_ori_n118_), .Y(ori_ori_n119_));
  NA2        o0070(.A(x3), .B(ori_ori_n100_), .Y(ori_ori_n120_));
  NA2        o0071(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n121_));
  INV        o0072(.A(x2), .Y(ori_ori_n122_));
  NA2        o0073(.A(x8), .B(x3), .Y(ori_ori_n123_));
  NA2        o0074(.A(ori_ori_n123_), .B(ori_ori_n72_), .Y(ori_ori_n124_));
  OAI220     o0075(.A0(ori_ori_n124_), .A1(ori_ori_n122_), .B0(ori_ori_n121_), .B1(ori_ori_n120_), .Y(ori_ori_n125_));
  NO2        o0076(.A(x5), .B(x0), .Y(ori_ori_n126_));
  NO2        o0077(.A(x6), .B(x1), .Y(ori_ori_n127_));
  NA3        o0078(.A(ori_ori_n127_), .B(ori_ori_n126_), .C(ori_ori_n125_), .Y(ori_ori_n128_));
  NA2        o0079(.A(x8), .B(ori_ori_n98_), .Y(ori_ori_n129_));
  NA2        o0080(.A(x4), .B(ori_ori_n50_), .Y(ori_ori_n130_));
  NO3        o0081(.A(ori_ori_n130_), .B(ori_ori_n129_), .C(ori_ori_n94_), .Y(ori_ori_n131_));
  NAi21      o0082(.An(x7), .B(x2), .Y(ori_ori_n132_));
  XO2        o0083(.A(x8), .B(x7), .Y(ori_ori_n133_));
  NA2        o0084(.A(ori_ori_n133_), .B(ori_ori_n100_), .Y(ori_ori_n134_));
  NA2        o0085(.A(x6), .B(x5), .Y(ori_ori_n135_));
  NO2        o0086(.A(ori_ori_n56_), .B(x0), .Y(ori_ori_n136_));
  NO2        o0087(.A(ori_ori_n50_), .B(x1), .Y(ori_ori_n137_));
  NA2        o0088(.A(ori_ori_n137_), .B(ori_ori_n136_), .Y(ori_ori_n138_));
  NO3        o0089(.A(ori_ori_n138_), .B(ori_ori_n135_), .C(ori_ori_n134_), .Y(ori_ori_n139_));
  AOI210     o0090(.A0(ori_ori_n2181_), .A1(ori_ori_n131_), .B0(ori_ori_n139_), .Y(ori_ori_n140_));
  NA3        o0091(.A(ori_ori_n140_), .B(ori_ori_n128_), .C(ori_ori_n119_), .Y(ori01));
  NO2        o0092(.A(x2), .B(x1), .Y(ori_ori_n142_));
  NA2        o0093(.A(x2), .B(x1), .Y(ori_ori_n143_));
  NOi21      o0094(.An(ori_ori_n143_), .B(ori_ori_n142_), .Y(ori_ori_n144_));
  NA2        o0095(.A(ori_ori_n98_), .B(ori_ori_n53_), .Y(ori_ori_n145_));
  NAi21      o0096(.An(x8), .B(x1), .Y(ori_ori_n146_));
  NO2        o0097(.A(ori_ori_n146_), .B(x3), .Y(ori_ori_n147_));
  NO2        o0098(.A(x5), .B(ori_ori_n50_), .Y(ori_ori_n148_));
  NO2        o0099(.A(ori_ori_n100_), .B(x1), .Y(ori_ori_n149_));
  NA2        o0100(.A(ori_ori_n149_), .B(ori_ori_n148_), .Y(ori_ori_n150_));
  NAi21      o0101(.An(x7), .B(x0), .Y(ori_ori_n151_));
  NO2        o0102(.A(ori_ori_n55_), .B(x2), .Y(ori_ori_n152_));
  NO2        o0103(.A(ori_ori_n78_), .B(x1), .Y(ori_ori_n153_));
  NA2        o0104(.A(x5), .B(ori_ori_n50_), .Y(ori_ori_n154_));
  NO2        o0105(.A(ori_ori_n154_), .B(ori_ori_n146_), .Y(ori_ori_n155_));
  NA2        o0106(.A(x8), .B(x5), .Y(ori_ori_n156_));
  NO3        o0107(.A(x3), .B(ori_ori_n100_), .C(ori_ori_n53_), .Y(ori_ori_n157_));
  INV        o0108(.A(ori_ori_n151_), .Y(ori_ori_n158_));
  INV        o0109(.A(x3), .Y(ori_ori_n159_));
  NO2        o0110(.A(ori_ori_n55_), .B(x0), .Y(ori_ori_n160_));
  NA3        o0111(.A(ori_ori_n98_), .B(ori_ori_n100_), .C(x1), .Y(ori_ori_n161_));
  NO2        o0112(.A(ori_ori_n161_), .B(ori_ori_n160_), .Y(ori_ori_n162_));
  NO2        o0113(.A(ori_ori_n83_), .B(ori_ori_n50_), .Y(ori_ori_n163_));
  NA2        o0114(.A(ori_ori_n98_), .B(x0), .Y(ori_ori_n164_));
  NA2        o0115(.A(ori_ori_n162_), .B(ori_ori_n159_), .Y(ori_ori_n165_));
  NA2        o0116(.A(x7), .B(ori_ori_n100_), .Y(ori_ori_n166_));
  NA2        o0117(.A(ori_ori_n148_), .B(x8), .Y(ori_ori_n167_));
  NA4        o0118(.A(x5), .B(x3), .C(x1), .D(x0), .Y(ori_ori_n168_));
  AO210      o0119(.A0(ori_ori_n168_), .A1(ori_ori_n167_), .B0(ori_ori_n166_), .Y(ori_ori_n169_));
  NO2        o0120(.A(ori_ori_n143_), .B(ori_ori_n50_), .Y(ori_ori_n170_));
  NAi21      o0121(.An(x1), .B(x2), .Y(ori_ori_n171_));
  NO2        o0122(.A(ori_ori_n154_), .B(ori_ori_n171_), .Y(ori_ori_n172_));
  NA2        o0123(.A(x8), .B(x7), .Y(ori_ori_n173_));
  NO2        o0124(.A(ori_ori_n173_), .B(x0), .Y(ori_ori_n174_));
  OAI210     o0125(.A0(ori_ori_n172_), .A1(ori_ori_n170_), .B0(ori_ori_n174_), .Y(ori_ori_n175_));
  NA3        o0126(.A(ori_ori_n175_), .B(ori_ori_n169_), .C(ori_ori_n165_), .Y(ori_ori_n176_));
  NO2        o0127(.A(ori_ori_n176_), .B(ori_ori_n158_), .Y(ori_ori_n177_));
  NA2        o0128(.A(x3), .B(x1), .Y(ori_ori_n178_));
  NA2        o0129(.A(ori_ori_n50_), .B(ori_ori_n100_), .Y(ori_ori_n179_));
  NO2        o0130(.A(ori_ori_n179_), .B(ori_ori_n67_), .Y(ori_ori_n180_));
  OAI210     o0131(.A0(ori_ori_n180_), .A1(ori_ori_n172_), .B0(ori_ori_n64_), .Y(ori_ori_n181_));
  NA2        o0132(.A(x8), .B(ori_ori_n100_), .Y(ori_ori_n182_));
  OAI210     o0133(.A0(ori_ori_n182_), .A1(ori_ori_n178_), .B0(ori_ori_n181_), .Y(ori_ori_n183_));
  XO2        o0134(.A(x5), .B(x3), .Y(ori_ori_n184_));
  NA2        o0135(.A(ori_ori_n184_), .B(x8), .Y(ori_ori_n185_));
  NA2        o0136(.A(x8), .B(ori_ori_n57_), .Y(ori_ori_n186_));
  NA2        o0137(.A(ori_ori_n186_), .B(ori_ori_n123_), .Y(ori_ori_n187_));
  NA2        o0138(.A(x7), .B(ori_ori_n68_), .Y(ori_ori_n188_));
  NO2        o0139(.A(ori_ori_n171_), .B(ori_ori_n188_), .Y(ori_ori_n189_));
  OA210      o0140(.A0(ori_ori_n187_), .A1(ori_ori_n184_), .B0(ori_ori_n189_), .Y(ori_ori_n190_));
  AOI220     o0141(.A0(ori_ori_n190_), .A1(ori_ori_n185_), .B0(ori_ori_n183_), .B1(x0), .Y(ori_ori_n191_));
  OAI210     o0142(.A0(ori_ori_n177_), .A1(ori_ori_n68_), .B0(ori_ori_n191_), .Y(ori_ori_n192_));
  NA4        o0143(.A(ori_ori_n55_), .B(x5), .C(x3), .D(x2), .Y(ori_ori_n193_));
  NA2        o0144(.A(x8), .B(ori_ori_n50_), .Y(ori_ori_n194_));
  NA2        o0145(.A(ori_ori_n194_), .B(x2), .Y(ori_ori_n195_));
  NA2        o0146(.A(ori_ori_n55_), .B(x3), .Y(ori_ori_n196_));
  NA4        o0147(.A(ori_ori_n196_), .B(ori_ori_n195_), .C(ori_ori_n184_), .D(ori_ori_n79_), .Y(ori_ori_n197_));
  AOI210     o0148(.A0(ori_ori_n197_), .A1(ori_ori_n193_), .B0(ori_ori_n53_), .Y(ori_ori_n198_));
  NO2        o0149(.A(ori_ori_n100_), .B(ori_ori_n57_), .Y(ori_ori_n199_));
  NA2        o0150(.A(x5), .B(x1), .Y(ori_ori_n200_));
  NO2        o0151(.A(ori_ori_n200_), .B(x6), .Y(ori_ori_n201_));
  NO2        o0152(.A(x3), .B(x1), .Y(ori_ori_n202_));
  AOI210     o0153(.A0(ori_ori_n202_), .A1(ori_ori_n74_), .B0(ori_ori_n201_), .Y(ori_ori_n203_));
  NO2        o0154(.A(ori_ori_n78_), .B(ori_ori_n55_), .Y(ori_ori_n204_));
  NO2        o0155(.A(ori_ori_n94_), .B(ori_ori_n50_), .Y(ori_ori_n205_));
  NO2        o0156(.A(ori_ori_n205_), .B(ori_ori_n204_), .Y(ori_ori_n206_));
  OAI210     o0157(.A0(ori_ori_n203_), .A1(x8), .B0(ori_ori_n206_), .Y(ori_ori_n207_));
  NO2        o0158(.A(ori_ori_n55_), .B(x5), .Y(ori_ori_n208_));
  NA2        o0159(.A(ori_ori_n208_), .B(ori_ori_n68_), .Y(ori_ori_n209_));
  NAi21      o0160(.An(x2), .B(x5), .Y(ori_ori_n210_));
  NA2        o0161(.A(x8), .B(x6), .Y(ori_ori_n211_));
  OAI210     o0162(.A0(ori_ori_n211_), .A1(ori_ori_n210_), .B0(ori_ori_n209_), .Y(ori_ori_n212_));
  NA2        o0163(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n213_));
  NO2        o0164(.A(ori_ori_n213_), .B(ori_ori_n57_), .Y(ori_ori_n214_));
  AO220      o0165(.A0(ori_ori_n214_), .A1(ori_ori_n212_), .B0(ori_ori_n207_), .B1(ori_ori_n199_), .Y(ori_ori_n215_));
  OAI210     o0166(.A0(ori_ori_n215_), .A1(ori_ori_n198_), .B0(x4), .Y(ori_ori_n216_));
  NA2        o0167(.A(ori_ori_n68_), .B(ori_ori_n56_), .Y(ori_ori_n217_));
  NO2        o0168(.A(ori_ori_n217_), .B(x7), .Y(ori_ori_n218_));
  NO2        o0169(.A(ori_ori_n98_), .B(ori_ori_n53_), .Y(ori_ori_n219_));
  NA2        o0170(.A(ori_ori_n219_), .B(ori_ori_n100_), .Y(ori_ori_n220_));
  NA2        o0171(.A(x3), .B(ori_ori_n57_), .Y(ori_ori_n221_));
  NO2        o0172(.A(ori_ori_n161_), .B(ori_ori_n221_), .Y(ori_ori_n222_));
  NO2        o0173(.A(x1), .B(x0), .Y(ori_ori_n223_));
  NA2        o0174(.A(ori_ori_n223_), .B(ori_ori_n100_), .Y(ori_ori_n224_));
  NA2        o0175(.A(ori_ori_n98_), .B(ori_ori_n50_), .Y(ori_ori_n225_));
  XN2        o0176(.A(x3), .B(x2), .Y(ori_ori_n226_));
  NO2        o0177(.A(ori_ori_n98_), .B(x0), .Y(ori_ori_n227_));
  NA2        o0178(.A(x8), .B(ori_ori_n53_), .Y(ori_ori_n228_));
  OAI210     o0179(.A0(ori_ori_n226_), .A1(x8), .B0(ori_ori_n218_), .Y(ori_ori_n229_));
  NO2        o0180(.A(x7), .B(x1), .Y(ori_ori_n230_));
  NOi21      o0181(.An(x8), .B(x3), .Y(ori_ori_n231_));
  NA2        o0182(.A(ori_ori_n231_), .B(ori_ori_n57_), .Y(ori_ori_n232_));
  NA2        o0183(.A(x5), .B(x0), .Y(ori_ori_n233_));
  NAi21      o0184(.An(ori_ori_n126_), .B(ori_ori_n233_), .Y(ori_ori_n234_));
  NA2        o0185(.A(ori_ori_n68_), .B(ori_ori_n50_), .Y(ori_ori_n235_));
  NA2        o0186(.A(ori_ori_n129_), .B(ori_ori_n230_), .Y(ori_ori_n236_));
  NO2        o0187(.A(ori_ori_n137_), .B(ori_ori_n68_), .Y(ori_ori_n237_));
  NA2        o0188(.A(x1), .B(x0), .Y(ori_ori_n238_));
  NA2        o0189(.A(ori_ori_n50_), .B(ori_ori_n57_), .Y(ori_ori_n239_));
  NA2        o0190(.A(ori_ori_n236_), .B(ori_ori_n168_), .Y(ori_ori_n240_));
  NO2        o0191(.A(ori_ori_n98_), .B(x3), .Y(ori_ori_n241_));
  NO2        o0192(.A(ori_ori_n100_), .B(x0), .Y(ori_ori_n242_));
  NA2        o0193(.A(ori_ori_n242_), .B(ori_ori_n241_), .Y(ori_ori_n243_));
  NO2        o0194(.A(ori_ori_n55_), .B(x7), .Y(ori_ori_n244_));
  NO3        o0195(.A(x8), .B(ori_ori_n50_), .C(x0), .Y(ori_ori_n245_));
  NAi21      o0196(.An(x8), .B(x0), .Y(ori_ori_n246_));
  NAi21      o0197(.An(x1), .B(x3), .Y(ori_ori_n247_));
  NO2        o0198(.A(ori_ori_n247_), .B(ori_ori_n246_), .Y(ori_ori_n248_));
  NO2        o0199(.A(x2), .B(ori_ori_n53_), .Y(ori_ori_n249_));
  AOI210     o0200(.A0(ori_ori_n249_), .A1(ori_ori_n245_), .B0(ori_ori_n248_), .Y(ori_ori_n250_));
  NOi21      o0201(.An(x5), .B(x6), .Y(ori_ori_n251_));
  INV        o0202(.A(x4), .Y(ori_ori_n252_));
  NA2        o0203(.A(ori_ori_n252_), .B(ori_ori_n251_), .Y(ori_ori_n253_));
  NO2        o0204(.A(ori_ori_n253_), .B(ori_ori_n250_), .Y(ori_ori_n254_));
  AOI210     o0205(.A0(ori_ori_n240_), .A1(ori_ori_n101_), .B0(ori_ori_n254_), .Y(ori_ori_n255_));
  NA3        o0206(.A(ori_ori_n255_), .B(ori_ori_n229_), .C(ori_ori_n216_), .Y(ori_ori_n256_));
  AOI210     o0207(.A0(ori_ori_n192_), .A1(ori_ori_n56_), .B0(ori_ori_n256_), .Y(ori02));
  NO2        o0208(.A(x8), .B(ori_ori_n98_), .Y(ori_ori_n258_));
  XN2        o0209(.A(x7), .B(x3), .Y(ori_ori_n259_));
  INV        o0210(.A(ori_ori_n259_), .Y(ori_ori_n260_));
  NO2        o0211(.A(x2), .B(x0), .Y(ori_ori_n261_));
  NA2        o0212(.A(ori_ori_n261_), .B(ori_ori_n68_), .Y(ori_ori_n262_));
  INV        o0213(.A(x1), .Y(ori_ori_n263_));
  NO3        o0214(.A(ori_ori_n263_), .B(ori_ori_n262_), .C(ori_ori_n260_), .Y(ori_ori_n264_));
  NA2        o0215(.A(ori_ori_n53_), .B(x0), .Y(ori_ori_n265_));
  NO2        o0216(.A(ori_ori_n247_), .B(x6), .Y(ori_ori_n266_));
  XO2        o0217(.A(x7), .B(x0), .Y(ori_ori_n267_));
  NO2        o0218(.A(ori_ori_n267_), .B(ori_ori_n261_), .Y(ori_ori_n268_));
  NA2        o0219(.A(ori_ori_n268_), .B(ori_ori_n266_), .Y(ori_ori_n269_));
  AN2        o0220(.A(x7), .B(x2), .Y(ori_ori_n270_));
  NA2        o0221(.A(ori_ori_n270_), .B(ori_ori_n50_), .Y(ori_ori_n271_));
  OAI210     o0222(.A0(ori_ori_n271_), .A1(ori_ori_n265_), .B0(ori_ori_n269_), .Y(ori_ori_n272_));
  OAI210     o0223(.A0(ori_ori_n272_), .A1(ori_ori_n264_), .B0(ori_ori_n258_), .Y(ori_ori_n273_));
  NAi21      o0224(.An(x8), .B(x6), .Y(ori_ori_n274_));
  NO2        o0225(.A(ori_ori_n98_), .B(ori_ori_n57_), .Y(ori_ori_n275_));
  NA2        o0226(.A(x7), .B(x3), .Y(ori_ori_n276_));
  NO2        o0227(.A(ori_ori_n276_), .B(x2), .Y(ori_ori_n277_));
  NA2        o0228(.A(x2), .B(x0), .Y(ori_ori_n278_));
  NA2        o0229(.A(ori_ori_n100_), .B(ori_ori_n57_), .Y(ori_ori_n279_));
  NAi21      o0230(.An(x7), .B(x1), .Y(ori_ori_n280_));
  AOI220     o0231(.A0(ori_ori_n2186_), .A1(x0), .B0(ori_ori_n277_), .B1(ori_ori_n275_), .Y(ori_ori_n281_));
  NA2        o0232(.A(ori_ori_n249_), .B(ori_ori_n50_), .Y(ori_ori_n282_));
  NA3        o0233(.A(x7), .B(ori_ori_n98_), .C(x0), .Y(ori_ori_n283_));
  OR2        o0234(.A(ori_ori_n283_), .B(ori_ori_n282_), .Y(ori_ori_n284_));
  AOI210     o0235(.A0(ori_ori_n284_), .A1(ori_ori_n281_), .B0(ori_ori_n274_), .Y(ori_ori_n285_));
  INV        o0236(.A(ori_ori_n267_), .Y(ori_ori_n286_));
  NO2        o0237(.A(x7), .B(ori_ori_n68_), .Y(ori_ori_n287_));
  NA2        o0238(.A(ori_ori_n98_), .B(x3), .Y(ori_ori_n288_));
  INV        o0239(.A(ori_ori_n288_), .Y(ori_ori_n289_));
  NA2        o0240(.A(ori_ori_n289_), .B(ori_ori_n286_), .Y(ori_ori_n290_));
  NA2        o0241(.A(ori_ori_n50_), .B(x0), .Y(ori_ori_n291_));
  NA2        o0242(.A(ori_ori_n152_), .B(x1), .Y(ori_ori_n292_));
  AOI210     o0243(.A0(x7), .A1(ori_ori_n290_), .B0(ori_ori_n292_), .Y(ori_ori_n293_));
  NO2        o0244(.A(ori_ori_n55_), .B(ori_ori_n100_), .Y(ori_ori_n294_));
  NA3        o0245(.A(ori_ori_n294_), .B(x3), .C(ori_ori_n57_), .Y(ori_ori_n295_));
  NO2        o0246(.A(ori_ori_n145_), .B(x6), .Y(ori_ori_n296_));
  NO2        o0247(.A(ori_ori_n94_), .B(ori_ori_n98_), .Y(ori_ori_n297_));
  NO2        o0248(.A(ori_ori_n295_), .B(ori_ori_n94_), .Y(ori_ori_n298_));
  NO3        o0249(.A(ori_ori_n298_), .B(ori_ori_n293_), .C(ori_ori_n285_), .Y(ori_ori_n299_));
  AOI210     o0250(.A0(ori_ori_n299_), .A1(ori_ori_n273_), .B0(x4), .Y(ori_ori_n300_));
  NA2        o0251(.A(x8), .B(ori_ori_n68_), .Y(ori_ori_n301_));
  NO2        o0252(.A(x3), .B(ori_ori_n57_), .Y(ori_ori_n302_));
  NA3        o0253(.A(ori_ori_n302_), .B(ori_ori_n98_), .C(ori_ori_n53_), .Y(ori_ori_n303_));
  NO2        o0254(.A(x3), .B(x0), .Y(ori_ori_n304_));
  NAi21      o0255(.An(ori_ori_n304_), .B(ori_ori_n97_), .Y(ori_ori_n305_));
  NA2        o0256(.A(x5), .B(x2), .Y(ori_ori_n306_));
  NO2        o0257(.A(ori_ori_n306_), .B(ori_ori_n202_), .Y(ori_ori_n307_));
  AOI210     o0258(.A0(ori_ori_n307_), .A1(ori_ori_n305_), .B0(ori_ori_n222_), .Y(ori_ori_n308_));
  AO210      o0259(.A0(ori_ori_n308_), .A1(ori_ori_n303_), .B0(ori_ori_n301_), .Y(ori_ori_n309_));
  NO2        o0260(.A(ori_ori_n100_), .B(ori_ori_n53_), .Y(ori_ori_n310_));
  NA2        o0261(.A(ori_ori_n310_), .B(x3), .Y(ori_ori_n311_));
  NO2        o0262(.A(ori_ori_n55_), .B(x1), .Y(ori_ori_n312_));
  NA2        o0263(.A(ori_ori_n312_), .B(ori_ori_n100_), .Y(ori_ori_n313_));
  OAI210     o0264(.A0(ori_ori_n313_), .A1(ori_ori_n154_), .B0(ori_ori_n311_), .Y(ori_ori_n314_));
  NAi32      o0265(.An(x3), .Bn(x0), .C(x2), .Y(ori_ori_n315_));
  NO2        o0266(.A(ori_ori_n50_), .B(x2), .Y(ori_ori_n316_));
  NAi21      o0267(.An(x6), .B(x5), .Y(ori_ori_n317_));
  NO2        o0268(.A(x2), .B(ori_ori_n57_), .Y(ori_ori_n318_));
  NO4        o0269(.A(ori_ori_n318_), .B(ori_ori_n317_), .C(ori_ori_n146_), .D(ori_ori_n316_), .Y(ori_ori_n319_));
  AOI220     o0270(.A0(ori_ori_n319_), .A1(ori_ori_n315_), .B0(ori_ori_n314_), .B1(ori_ori_n82_), .Y(ori_ori_n320_));
  AOI210     o0271(.A0(ori_ori_n320_), .A1(ori_ori_n309_), .B0(ori_ori_n72_), .Y(ori_ori_n321_));
  NA2        o0272(.A(ori_ori_n312_), .B(ori_ori_n56_), .Y(ori_ori_n322_));
  NO2        o0273(.A(ori_ori_n98_), .B(ori_ori_n50_), .Y(ori_ori_n323_));
  NO2        o0274(.A(ori_ori_n261_), .B(ori_ori_n199_), .Y(ori_ori_n324_));
  XO2        o0275(.A(x7), .B(x2), .Y(ori_ori_n325_));
  INV        o0276(.A(ori_ori_n325_), .Y(ori_ori_n326_));
  XO2        o0277(.A(x6), .B(x2), .Y(ori_ori_n327_));
  NA4        o0278(.A(ori_ori_n327_), .B(ori_ori_n326_), .C(ori_ori_n324_), .D(ori_ori_n323_), .Y(ori_ori_n328_));
  NAi21      o0279(.An(x0), .B(x6), .Y(ori_ori_n329_));
  AOI210     o0280(.A0(ori_ori_n329_), .A1(ori_ori_n132_), .B0(ori_ori_n242_), .Y(ori_ori_n330_));
  XN2        o0281(.A(x7), .B(x5), .Y(ori_ori_n331_));
  NA2        o0282(.A(ori_ori_n331_), .B(ori_ori_n68_), .Y(ori_ori_n332_));
  NA2        o0283(.A(x7), .B(x5), .Y(ori_ori_n333_));
  AOI210     o0284(.A0(ori_ori_n333_), .A1(x6), .B0(ori_ori_n315_), .Y(ori_ori_n334_));
  AOI220     o0285(.A0(ori_ori_n334_), .A1(ori_ori_n332_), .B0(ori_ori_n330_), .B1(ori_ori_n289_), .Y(ori_ori_n335_));
  AOI210     o0286(.A0(ori_ori_n335_), .A1(ori_ori_n328_), .B0(ori_ori_n322_), .Y(ori_ori_n336_));
  NO2        o0287(.A(x8), .B(x6), .Y(ori_ori_n337_));
  NAi21      o0288(.An(ori_ori_n337_), .B(ori_ori_n211_), .Y(ori_ori_n338_));
  NA2        o0289(.A(ori_ori_n98_), .B(x2), .Y(ori_ori_n339_));
  NA2        o0290(.A(x1), .B(ori_ori_n57_), .Y(ori_ori_n340_));
  NA2        o0291(.A(x4), .B(x2), .Y(ori_ori_n341_));
  NO2        o0292(.A(ori_ori_n341_), .B(ori_ori_n98_), .Y(ori_ori_n342_));
  NAi21      o0293(.An(x1), .B(x6), .Y(ori_ori_n343_));
  NA2        o0294(.A(ori_ori_n304_), .B(ori_ori_n244_), .Y(ori_ori_n344_));
  NA2        o0295(.A(x8), .B(x2), .Y(ori_ori_n345_));
  NO2        o0296(.A(ori_ori_n345_), .B(ori_ori_n50_), .Y(ori_ori_n346_));
  INV        o0297(.A(ori_ori_n201_), .Y(ori_ori_n347_));
  NO2        o0298(.A(ori_ori_n347_), .B(ori_ori_n52_), .Y(ori_ori_n348_));
  AOI220     o0299(.A0(ori_ori_n348_), .A1(ori_ori_n346_), .B0(ori_ori_n2166_), .B1(ori_ori_n342_), .Y(ori_ori_n349_));
  INV        o0300(.A(ori_ori_n349_), .Y(ori_ori_n350_));
  NO4        o0301(.A(ori_ori_n350_), .B(ori_ori_n336_), .C(ori_ori_n321_), .D(ori_ori_n300_), .Y(ori03));
  NAi21      o0302(.An(x2), .B(x0), .Y(ori_ori_n352_));
  NO3        o0303(.A(x8), .B(x6), .C(x4), .Y(ori_ori_n353_));
  INV        o0304(.A(ori_ori_n353_), .Y(ori_ori_n354_));
  NO2        o0305(.A(ori_ori_n354_), .B(ori_ori_n352_), .Y(ori_ori_n355_));
  NA2        o0306(.A(ori_ori_n101_), .B(ori_ori_n57_), .Y(ori_ori_n356_));
  NO2        o0307(.A(ori_ori_n356_), .B(ori_ori_n55_), .Y(ori_ori_n357_));
  OAI210     o0308(.A0(ori_ori_n357_), .A1(ori_ori_n355_), .B0(ori_ori_n148_), .Y(ori_ori_n358_));
  NA2        o0309(.A(x3), .B(x2), .Y(ori_ori_n359_));
  NO2        o0310(.A(ori_ori_n146_), .B(x0), .Y(ori_ori_n360_));
  NA2        o0311(.A(x8), .B(x0), .Y(ori_ori_n361_));
  NO2        o0312(.A(ori_ori_n361_), .B(x6), .Y(ori_ori_n362_));
  NO2        o0313(.A(x5), .B(ori_ori_n57_), .Y(ori_ori_n363_));
  NO2        o0314(.A(x3), .B(x2), .Y(ori_ori_n364_));
  NA2        o0315(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n365_));
  NO2        o0316(.A(ori_ori_n53_), .B(x0), .Y(ori_ori_n366_));
  NA2        o0317(.A(ori_ori_n366_), .B(x5), .Y(ori_ori_n367_));
  NO2        o0318(.A(ori_ori_n50_), .B(ori_ori_n57_), .Y(ori_ori_n368_));
  NO2        o0319(.A(ori_ori_n68_), .B(x0), .Y(ori_ori_n369_));
  OAI210     o0320(.A0(x5), .A1(ori_ori_n360_), .B0(x4), .Y(ori_ori_n370_));
  NO2        o0321(.A(x4), .B(ori_ori_n53_), .Y(ori_ori_n371_));
  NA2        o0322(.A(ori_ori_n371_), .B(ori_ori_n57_), .Y(ori_ori_n372_));
  NO3        o0323(.A(ori_ori_n372_), .B(ori_ori_n211_), .C(x5), .Y(ori_ori_n373_));
  NA2        o0324(.A(x7), .B(ori_ori_n98_), .Y(ori_ori_n374_));
  NO3        o0325(.A(x5), .B(ori_ori_n53_), .C(x0), .Y(ori_ori_n375_));
  INV        o0326(.A(ori_ori_n375_), .Y(ori_ori_n376_));
  NO2        o0327(.A(x6), .B(ori_ori_n56_), .Y(ori_ori_n377_));
  NO2        o0328(.A(x8), .B(ori_ori_n50_), .Y(ori_ori_n378_));
  NA2        o0329(.A(ori_ori_n378_), .B(ori_ori_n377_), .Y(ori_ori_n379_));
  AOI210     o0330(.A0(ori_ori_n373_), .A1(x2), .B0(x7), .Y(ori_ori_n380_));
  AOI220     o0331(.A0(ori_ori_n380_), .A1(ori_ori_n370_), .B0(ori_ori_n358_), .B1(x7), .Y(ori_ori_n381_));
  NO2        o0332(.A(ori_ori_n231_), .B(ori_ori_n100_), .Y(ori_ori_n382_));
  NO2        o0333(.A(ori_ori_n55_), .B(ori_ori_n57_), .Y(ori_ori_n383_));
  NO3        o0334(.A(ori_ori_n383_), .B(ori_ori_n382_), .C(ori_ori_n135_), .Y(ori_ori_n384_));
  AOI210     o0335(.A0(ori_ori_n187_), .A1(ori_ori_n92_), .B0(ori_ori_n384_), .Y(ori_ori_n385_));
  NO2        o0336(.A(x5), .B(x2), .Y(ori_ori_n386_));
  NO2        o0337(.A(x8), .B(x3), .Y(ori_ori_n387_));
  NA2        o0338(.A(ori_ori_n186_), .B(x2), .Y(ori_ori_n388_));
  NO3        o0339(.A(ori_ori_n387_), .B(ori_ori_n305_), .C(ori_ori_n317_), .Y(ori_ori_n389_));
  NA2        o0340(.A(ori_ori_n389_), .B(ori_ori_n388_), .Y(ori_ori_n390_));
  OAI210     o0341(.A0(ori_ori_n385_), .A1(ori_ori_n261_), .B0(ori_ori_n390_), .Y(ori_ori_n391_));
  NA2        o0342(.A(ori_ori_n391_), .B(x4), .Y(ori_ori_n392_));
  NA2        o0343(.A(ori_ori_n55_), .B(ori_ori_n57_), .Y(ori_ori_n393_));
  NO2        o0344(.A(ori_ori_n393_), .B(x5), .Y(ori_ori_n394_));
  NAi21      o0345(.An(x4), .B(x6), .Y(ori_ori_n395_));
  NO2        o0346(.A(ori_ori_n395_), .B(ori_ori_n51_), .Y(ori_ori_n396_));
  NO2        o0347(.A(ori_ori_n55_), .B(ori_ori_n68_), .Y(ori_ori_n397_));
  NO2        o0348(.A(ori_ori_n50_), .B(ori_ori_n100_), .Y(ori_ori_n398_));
  NO2        o0349(.A(ori_ori_n211_), .B(x0), .Y(ori_ori_n399_));
  NO2        o0350(.A(ori_ori_n317_), .B(x8), .Y(ori_ori_n400_));
  OAI210     o0351(.A0(ori_ori_n400_), .A1(ori_ori_n399_), .B0(ori_ori_n398_), .Y(ori_ori_n401_));
  OAI210     o0352(.A0(ori_ori_n365_), .A1(ori_ori_n397_), .B0(ori_ori_n401_), .Y(ori_ori_n402_));
  AOI220     o0353(.A0(ori_ori_n402_), .A1(ori_ori_n56_), .B0(ori_ori_n396_), .B1(ori_ori_n394_), .Y(ori_ori_n403_));
  AOI210     o0354(.A0(ori_ori_n403_), .A1(ori_ori_n392_), .B0(x1), .Y(ori_ori_n404_));
  NO2        o0355(.A(ori_ori_n68_), .B(ori_ori_n56_), .Y(ori_ori_n405_));
  NA2        o0356(.A(ori_ori_n316_), .B(ori_ori_n57_), .Y(ori_ori_n406_));
  NO2        o0357(.A(x8), .B(x5), .Y(ori_ori_n407_));
  NAi21      o0358(.An(ori_ori_n407_), .B(ori_ori_n156_), .Y(ori_ori_n408_));
  NA2        o0359(.A(ori_ori_n324_), .B(ori_ori_n74_), .Y(ori_ori_n409_));
  NOi21      o0360(.An(x3), .B(x4), .Y(ori_ori_n410_));
  NA2        o0361(.A(ori_ori_n55_), .B(ori_ori_n100_), .Y(ori_ori_n411_));
  NO2        o0362(.A(ori_ori_n135_), .B(ori_ori_n55_), .Y(ori_ori_n412_));
  NO3        o0363(.A(ori_ori_n56_), .B(x2), .C(x0), .Y(ori_ori_n413_));
  NA2        o0364(.A(x7), .B(x1), .Y(ori_ori_n414_));
  NO3        o0365(.A(x5), .B(x4), .C(x2), .Y(ori_ori_n415_));
  AN2        o0366(.A(ori_ori_n415_), .B(ori_ori_n337_), .Y(ori_ori_n416_));
  NO3        o0367(.A(ori_ori_n416_), .B(ori_ori_n412_), .C(ori_ori_n342_), .Y(ori_ori_n417_));
  OAI210     o0368(.A0(ori_ori_n337_), .A1(ori_ori_n81_), .B0(ori_ori_n304_), .Y(ori_ori_n418_));
  NO2        o0369(.A(ori_ori_n418_), .B(ori_ori_n417_), .Y(ori_ori_n419_));
  NO2        o0370(.A(x4), .B(ori_ori_n100_), .Y(ori_ori_n420_));
  NA2        o0371(.A(ori_ori_n420_), .B(x6), .Y(ori_ori_n421_));
  NA3        o0372(.A(ori_ori_n98_), .B(x4), .C(ori_ori_n100_), .Y(ori_ori_n422_));
  AOI210     o0373(.A0(ori_ori_n422_), .A1(ori_ori_n421_), .B0(ori_ori_n91_), .Y(ori_ori_n423_));
  NA2        o0374(.A(ori_ori_n410_), .B(ori_ori_n68_), .Y(ori_ori_n424_));
  NA2        o0375(.A(ori_ori_n152_), .B(ori_ori_n57_), .Y(ori_ori_n425_));
  NO2        o0376(.A(ori_ori_n425_), .B(ori_ori_n424_), .Y(ori_ori_n426_));
  NA2        o0377(.A(ori_ori_n398_), .B(x4), .Y(ori_ori_n427_));
  NO3        o0378(.A(ori_ori_n427_), .B(ori_ori_n337_), .C(ori_ori_n369_), .Y(ori_ori_n428_));
  NO4        o0379(.A(ori_ori_n428_), .B(ori_ori_n426_), .C(ori_ori_n423_), .D(ori_ori_n419_), .Y(ori_ori_n429_));
  NA2        o0380(.A(x5), .B(x4), .Y(ori_ori_n430_));
  NO2        o0381(.A(ori_ori_n68_), .B(ori_ori_n53_), .Y(ori_ori_n431_));
  NO3        o0382(.A(x8), .B(x3), .C(x2), .Y(ori_ori_n432_));
  NA3        o0383(.A(ori_ori_n432_), .B(ori_ori_n431_), .C(ori_ori_n57_), .Y(ori_ori_n433_));
  NO3        o0384(.A(x6), .B(x5), .C(x2), .Y(ori_ori_n434_));
  NA3        o0385(.A(ori_ori_n434_), .B(ori_ori_n263_), .C(ori_ori_n75_), .Y(ori_ori_n435_));
  OAI210     o0386(.A0(ori_ori_n433_), .A1(ori_ori_n430_), .B0(ori_ori_n435_), .Y(ori_ori_n436_));
  NA2        o0387(.A(ori_ori_n68_), .B(x2), .Y(ori_ori_n437_));
  NO3        o0388(.A(x4), .B(x3), .C(ori_ori_n57_), .Y(ori_ori_n438_));
  NA2        o0389(.A(ori_ori_n438_), .B(ori_ori_n208_), .Y(ori_ori_n439_));
  NO3        o0390(.A(ori_ori_n439_), .B(ori_ori_n437_), .C(ori_ori_n87_), .Y(ori_ori_n440_));
  XO2        o0391(.A(x4), .B(x0), .Y(ori_ori_n441_));
  NA2        o0392(.A(ori_ori_n239_), .B(x5), .Y(ori_ori_n442_));
  NO2        o0393(.A(ori_ori_n56_), .B(ori_ori_n50_), .Y(ori_ori_n443_));
  NO2        o0394(.A(ori_ori_n443_), .B(ori_ori_n61_), .Y(ori_ori_n444_));
  NO4        o0395(.A(ori_ori_n444_), .B(ori_ori_n442_), .C(ori_ori_n441_), .D(ori_ori_n143_), .Y(ori_ori_n445_));
  NO3        o0396(.A(ori_ori_n445_), .B(ori_ori_n440_), .C(ori_ori_n436_), .Y(ori_ori_n446_));
  OAI210     o0397(.A0(ori_ori_n429_), .A1(ori_ori_n414_), .B0(ori_ori_n446_), .Y(ori_ori_n447_));
  NO3        o0398(.A(ori_ori_n447_), .B(ori_ori_n404_), .C(ori_ori_n381_), .Y(ori04));
  NO2        o0399(.A(x7), .B(x2), .Y(ori_ori_n449_));
  NO2        o0400(.A(x3), .B(ori_ori_n53_), .Y(ori_ori_n450_));
  NO2        o0401(.A(ori_ori_n450_), .B(ori_ori_n137_), .Y(ori_ori_n451_));
  XN2        o0402(.A(x8), .B(x1), .Y(ori_ori_n452_));
  NO2        o0403(.A(ori_ori_n452_), .B(ori_ori_n135_), .Y(ori_ori_n453_));
  NA2        o0404(.A(ori_ori_n453_), .B(ori_ori_n451_), .Y(ori_ori_n454_));
  NA2        o0405(.A(x6), .B(x3), .Y(ori_ori_n455_));
  NA2        o0406(.A(ori_ori_n68_), .B(x1), .Y(ori_ori_n456_));
  NO2        o0407(.A(ori_ori_n407_), .B(ori_ori_n231_), .Y(ori_ori_n457_));
  NOi21      o0408(.An(ori_ori_n156_), .B(ori_ori_n407_), .Y(ori_ori_n458_));
  NA2        o0409(.A(ori_ori_n99_), .B(x1), .Y(ori_ori_n459_));
  NA2        o0410(.A(ori_ori_n123_), .B(ori_ori_n221_), .Y(ori_ori_n460_));
  OR4        o0411(.A(ori_ori_n460_), .B(ori_ori_n338_), .C(ori_ori_n79_), .D(ori_ori_n54_), .Y(ori_ori_n461_));
  OR2        o0412(.A(x6), .B(x0), .Y(ori_ori_n462_));
  NO3        o0413(.A(ori_ori_n462_), .B(x3), .C(x1), .Y(ori_ori_n463_));
  AOI220     o0414(.A0(ori_ori_n463_), .A1(ori_ori_n98_), .B0(ori_ori_n251_), .B1(ori_ori_n245_), .Y(ori_ori_n464_));
  AOI210     o0415(.A0(ori_ori_n464_), .A1(ori_ori_n461_), .B0(ori_ori_n166_), .Y(ori_ori_n465_));
  NA2        o0416(.A(x7), .B(x2), .Y(ori_ori_n466_));
  INV        o0417(.A(ori_ori_n123_), .Y(ori_ori_n467_));
  OAI210     o0418(.A0(ori_ori_n155_), .A1(ori_ori_n467_), .B0(ori_ori_n79_), .Y(ori_ori_n468_));
  NO2        o0419(.A(ori_ori_n288_), .B(ori_ori_n55_), .Y(ori_ori_n469_));
  NO3        o0420(.A(x3), .B(x1), .C(x0), .Y(ori_ori_n470_));
  OR2        o0421(.A(x6), .B(x1), .Y(ori_ori_n471_));
  NA2        o0422(.A(ori_ori_n471_), .B(x0), .Y(ori_ori_n472_));
  AOI220     o0423(.A0(ori_ori_n472_), .A1(ori_ori_n469_), .B0(ori_ori_n470_), .B1(ori_ori_n412_), .Y(ori_ori_n473_));
  AOI210     o0424(.A0(ori_ori_n473_), .A1(ori_ori_n468_), .B0(ori_ori_n466_), .Y(ori_ori_n474_));
  NA2        o0425(.A(ori_ori_n68_), .B(x0), .Y(ori_ori_n475_));
  NO3        o0426(.A(ori_ori_n474_), .B(ori_ori_n465_), .C(ori_ori_n56_), .Y(ori_ori_n476_));
  INV        o0427(.A(ori_ori_n476_), .Y(ori_ori_n477_));
  NA3        o0428(.A(x8), .B(x7), .C(x0), .Y(ori_ori_n478_));
  INV        o0429(.A(ori_ori_n478_), .Y(ori_ori_n479_));
  AOI210     o0430(.A0(ori_ori_n244_), .A1(ori_ori_n90_), .B0(ori_ori_n479_), .Y(ori_ori_n480_));
  NO2        o0431(.A(ori_ori_n480_), .B(ori_ori_n143_), .Y(ori_ori_n481_));
  NO2        o0432(.A(x8), .B(x0), .Y(ori_ori_n482_));
  NA2        o0433(.A(ori_ori_n482_), .B(ori_ori_n326_), .Y(ori_ori_n483_));
  NO2        o0434(.A(ori_ori_n483_), .B(ori_ori_n247_), .Y(ori_ori_n484_));
  OAI210     o0435(.A0(ori_ori_n484_), .A1(ori_ori_n481_), .B0(ori_ori_n251_), .Y(ori_ori_n485_));
  NO2        o0436(.A(ori_ori_n68_), .B(ori_ori_n100_), .Y(ori_ori_n486_));
  NO2        o0437(.A(ori_ori_n333_), .B(x8), .Y(ori_ori_n487_));
  INV        o0438(.A(ori_ori_n487_), .Y(ori_ori_n488_));
  NO3        o0439(.A(ori_ori_n488_), .B(ori_ori_n340_), .C(ori_ori_n241_), .Y(ori_ori_n489_));
  NO2        o0440(.A(ori_ori_n260_), .B(x8), .Y(ori_ori_n490_));
  OAI210     o0441(.A0(ori_ori_n407_), .A1(x3), .B0(ori_ori_n223_), .Y(ori_ori_n491_));
  NA2        o0442(.A(ori_ori_n312_), .B(ori_ori_n159_), .Y(ori_ori_n492_));
  OAI220     o0443(.A0(ori_ori_n492_), .A1(ori_ori_n57_), .B0(ori_ori_n491_), .B1(ori_ori_n490_), .Y(ori_ori_n493_));
  OAI210     o0444(.A0(ori_ori_n493_), .A1(ori_ori_n489_), .B0(ori_ori_n486_), .Y(ori_ori_n494_));
  NO2        o0445(.A(x8), .B(x2), .Y(ori_ori_n495_));
  INV        o0446(.A(ori_ori_n202_), .Y(ori_ori_n496_));
  NA3        o0447(.A(ori_ori_n496_), .B(ori_ori_n495_), .C(ori_ori_n305_), .Y(ori_ori_n497_));
  NO2        o0448(.A(ori_ori_n224_), .B(ori_ori_n123_), .Y(ori_ori_n498_));
  AOI210     o0449(.A0(ori_ori_n2179_), .A1(ori_ori_n149_), .B0(ori_ori_n498_), .Y(ori_ori_n499_));
  AOI210     o0450(.A0(ori_ori_n499_), .A1(ori_ori_n497_), .B0(ori_ori_n99_), .Y(ori_ori_n500_));
  NA2        o0451(.A(ori_ori_n302_), .B(x2), .Y(ori_ori_n501_));
  NA2        o0452(.A(x1), .B(ori_ori_n61_), .Y(ori_ori_n502_));
  AOI210     o0453(.A0(ori_ori_n501_), .A1(ori_ori_n406_), .B0(ori_ori_n502_), .Y(ori_ori_n503_));
  NA2        o0454(.A(ori_ori_n100_), .B(ori_ori_n53_), .Y(ori_ori_n504_));
  NO2        o0455(.A(ori_ori_n504_), .B(x8), .Y(ori_ori_n505_));
  NA2        o0456(.A(x7), .B(ori_ori_n50_), .Y(ori_ori_n506_));
  NO2        o0457(.A(ori_ori_n164_), .B(ori_ori_n506_), .Y(ori_ori_n507_));
  AN2        o0458(.A(ori_ori_n507_), .B(ori_ori_n505_), .Y(ori_ori_n508_));
  NA2        o0459(.A(ori_ori_n363_), .B(ori_ori_n137_), .Y(ori_ori_n509_));
  NO2        o0460(.A(ori_ori_n68_), .B(x2), .Y(ori_ori_n510_));
  NA2        o0461(.A(ori_ori_n510_), .B(ori_ori_n244_), .Y(ori_ori_n511_));
  OAI210     o0462(.A0(ori_ori_n511_), .A1(ori_ori_n509_), .B0(ori_ori_n56_), .Y(ori_ori_n512_));
  NO4        o0463(.A(ori_ori_n512_), .B(ori_ori_n508_), .C(ori_ori_n503_), .D(ori_ori_n500_), .Y(ori_ori_n513_));
  NA3        o0464(.A(ori_ori_n513_), .B(ori_ori_n494_), .C(ori_ori_n485_), .Y(ori_ori_n514_));
  NA2        o0465(.A(ori_ori_n53_), .B(ori_ori_n57_), .Y(ori_ori_n515_));
  NOi21      o0466(.An(x2), .B(x7), .Y(ori_ori_n516_));
  NO2        o0467(.A(x6), .B(x3), .Y(ori_ori_n517_));
  NA2        o0468(.A(ori_ori_n517_), .B(ori_ori_n516_), .Y(ori_ori_n518_));
  NO2        o0469(.A(x6), .B(ori_ori_n57_), .Y(ori_ori_n519_));
  NO2        o0470(.A(x2), .B(x1), .Y(ori_ori_n520_));
  NO2        o0471(.A(x2), .B(x0), .Y(ori_ori_n521_));
  AOI220     o0472(.A0(ori_ori_n521_), .A1(ori_ori_n205_), .B0(ori_ori_n520_), .B1(ori_ori_n519_), .Y(ori_ori_n522_));
  OAI210     o0473(.A0(ori_ori_n518_), .A1(ori_ori_n515_), .B0(ori_ori_n522_), .Y(ori_ori_n523_));
  NO2        o0474(.A(ori_ori_n92_), .B(ori_ori_n53_), .Y(ori_ori_n524_));
  NO2        o0475(.A(ori_ori_n524_), .B(ori_ori_n400_), .Y(ori_ori_n525_));
  NO3        o0476(.A(ori_ori_n525_), .B(ori_ori_n427_), .C(ori_ori_n57_), .Y(ori_ori_n526_));
  AO210      o0477(.A0(ori_ori_n523_), .A1(ori_ori_n407_), .B0(ori_ori_n526_), .Y(ori_ori_n527_));
  AOI210     o0478(.A0(ori_ori_n514_), .A1(ori_ori_n477_), .B0(ori_ori_n527_), .Y(ori05));
  AOI210     o0479(.A0(ori_ori_n148_), .A1(ori_ori_n55_), .B0(ori_ori_n443_), .Y(ori_ori_n529_));
  NO2        o0480(.A(x7), .B(ori_ori_n98_), .Y(ori_ori_n530_));
  NO2        o0481(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n531_));
  NA2        o0482(.A(x5), .B(ori_ori_n56_), .Y(ori_ori_n532_));
  NO2        o0483(.A(ori_ori_n532_), .B(ori_ori_n506_), .Y(ori_ori_n533_));
  AOI210     o0484(.A0(ori_ori_n531_), .A1(ori_ori_n530_), .B0(ori_ori_n533_), .Y(ori_ori_n534_));
  AOI210     o0485(.A0(ori_ori_n534_), .A1(ori_ori_n529_), .B0(ori_ori_n100_), .Y(ori_ori_n535_));
  NO2        o0486(.A(x7), .B(x4), .Y(ori_ori_n536_));
  NO2        o0487(.A(ori_ori_n179_), .B(x5), .Y(ori_ori_n537_));
  NA2        o0488(.A(ori_ori_n98_), .B(ori_ori_n100_), .Y(ori_ori_n538_));
  NO2        o0489(.A(ori_ori_n538_), .B(ori_ori_n196_), .Y(ori_ori_n539_));
  AN2        o0490(.A(ori_ori_n539_), .B(ori_ori_n536_), .Y(ori_ori_n540_));
  OAI210     o0491(.A0(ori_ori_n540_), .A1(ori_ori_n535_), .B0(ori_ori_n431_), .Y(ori_ori_n541_));
  NO2        o0492(.A(x6), .B(ori_ori_n50_), .Y(ori_ori_n542_));
  NA2        o0493(.A(ori_ori_n55_), .B(x4), .Y(ori_ori_n543_));
  NO2        o0494(.A(ori_ori_n98_), .B(ori_ori_n100_), .Y(ori_ori_n544_));
  NA2        o0495(.A(ori_ori_n544_), .B(x7), .Y(ori_ori_n545_));
  NA2        o0496(.A(ori_ori_n386_), .B(ori_ori_n230_), .Y(ori_ori_n546_));
  AOI210     o0497(.A0(ori_ori_n546_), .A1(ori_ori_n545_), .B0(ori_ori_n543_), .Y(ori_ori_n547_));
  NA2        o0498(.A(ori_ori_n98_), .B(x4), .Y(ori_ori_n548_));
  XO2        o0499(.A(x7), .B(x5), .Y(ori_ori_n549_));
  NO2        o0500(.A(ori_ori_n549_), .B(ori_ori_n53_), .Y(ori_ori_n550_));
  NA2        o0501(.A(ori_ori_n550_), .B(ori_ori_n294_), .Y(ori_ori_n551_));
  NO2        o0502(.A(ori_ori_n98_), .B(x2), .Y(ori_ori_n552_));
  NO2        o0503(.A(ori_ori_n72_), .B(ori_ori_n55_), .Y(ori_ori_n553_));
  NA2        o0504(.A(ori_ori_n553_), .B(ori_ori_n552_), .Y(ori_ori_n554_));
  NA2        o0505(.A(ori_ori_n554_), .B(ori_ori_n551_), .Y(ori_ori_n555_));
  OAI210     o0506(.A0(ori_ori_n555_), .A1(ori_ori_n547_), .B0(ori_ori_n542_), .Y(ori_ori_n556_));
  NO2        o0507(.A(ori_ori_n68_), .B(ori_ori_n50_), .Y(ori_ori_n557_));
  NO2        o0508(.A(ori_ori_n173_), .B(x4), .Y(ori_ori_n558_));
  NO2        o0509(.A(x5), .B(ori_ori_n56_), .Y(ori_ori_n559_));
  XO2        o0510(.A(x5), .B(x2), .Y(ori_ori_n560_));
  NO3        o0511(.A(x8), .B(x7), .C(ori_ori_n100_), .Y(ori_ori_n561_));
  AO220      o0512(.A0(ori_ori_n561_), .A1(ori_ori_n559_), .B0(ori_ori_n560_), .B1(ori_ori_n558_), .Y(ori_ori_n562_));
  NA3        o0513(.A(ori_ori_n562_), .B(ori_ori_n557_), .C(ori_ori_n53_), .Y(ori_ori_n563_));
  NA2        o0514(.A(ori_ori_n241_), .B(ori_ori_n516_), .Y(ori_ori_n564_));
  NOi21      o0515(.An(x4), .B(x1), .Y(ori_ori_n565_));
  NA2        o0516(.A(ori_ori_n565_), .B(ori_ori_n61_), .Y(ori_ori_n566_));
  NA2        o0517(.A(x4), .B(x1), .Y(ori_ori_n567_));
  NO2        o0518(.A(ori_ori_n567_), .B(ori_ori_n50_), .Y(ori_ori_n568_));
  AOI210     o0519(.A0(ori_ori_n568_), .A1(ori_ori_n544_), .B0(ori_ori_n57_), .Y(ori_ori_n569_));
  OA210      o0520(.A0(ori_ori_n566_), .A1(ori_ori_n564_), .B0(ori_ori_n569_), .Y(ori_ori_n570_));
  NA4        o0521(.A(ori_ori_n570_), .B(ori_ori_n563_), .C(ori_ori_n556_), .D(ori_ori_n541_), .Y(ori_ori_n571_));
  NA2        o0522(.A(ori_ori_n557_), .B(ori_ori_n56_), .Y(ori_ori_n572_));
  OAI210     o0523(.A0(x7), .A1(ori_ori_n150_), .B0(ori_ori_n57_), .Y(ori_ori_n573_));
  INV        o0524(.A(x3), .Y(ori_ori_n574_));
  NA2        o0525(.A(ori_ori_n559_), .B(ori_ori_n142_), .Y(ori_ori_n575_));
  NO3        o0526(.A(ori_ori_n575_), .B(ori_ori_n574_), .C(ori_ori_n378_), .Y(ori_ori_n576_));
  NA2        o0527(.A(ori_ori_n252_), .B(ori_ori_n68_), .Y(ori_ori_n577_));
  NO2        o0528(.A(ori_ori_n345_), .B(x3), .Y(ori_ori_n578_));
  NA2        o0529(.A(ori_ori_n578_), .B(ori_ori_n219_), .Y(ori_ori_n579_));
  NO2        o0530(.A(ori_ori_n378_), .B(ori_ori_n558_), .Y(ori_ori_n580_));
  NO2        o0531(.A(ori_ori_n410_), .B(ori_ori_n98_), .Y(ori_ori_n581_));
  NO2        o0532(.A(ori_ori_n504_), .B(x6), .Y(ori_ori_n582_));
  NA2        o0533(.A(ori_ori_n582_), .B(ori_ori_n581_), .Y(ori_ori_n583_));
  OAI220     o0534(.A0(ori_ori_n583_), .A1(ori_ori_n580_), .B0(ori_ori_n579_), .B1(ori_ori_n577_), .Y(ori_ori_n584_));
  NO3        o0535(.A(ori_ori_n584_), .B(ori_ori_n576_), .C(ori_ori_n573_), .Y(ori_ori_n585_));
  NA2        o0536(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n586_));
  NO2        o0537(.A(ori_ori_n586_), .B(ori_ori_n120_), .Y(ori_ori_n587_));
  NA2        o0538(.A(x8), .B(x4), .Y(ori_ori_n588_));
  NO2        o0539(.A(x8), .B(x4), .Y(ori_ori_n589_));
  NAi21      o0540(.An(ori_ori_n589_), .B(ori_ori_n588_), .Y(ori_ori_n590_));
  NAi21      o0541(.An(ori_ori_n495_), .B(ori_ori_n345_), .Y(ori_ori_n591_));
  NO3        o0542(.A(x8), .B(ori_ori_n98_), .C(x4), .Y(ori_ori_n592_));
  INV        o0543(.A(ori_ori_n592_), .Y(ori_ori_n593_));
  NO2        o0544(.A(x5), .B(x4), .Y(ori_ori_n594_));
  NO2        o0545(.A(x6), .B(ori_ori_n100_), .Y(ori_ori_n595_));
  NA2        o0546(.A(ori_ori_n586_), .B(ori_ori_n595_), .Y(ori_ori_n596_));
  NA2        o0547(.A(ori_ori_n2173_), .B(ori_ori_n2186_), .Y(ori_ori_n597_));
  NA2        o0548(.A(ori_ori_n597_), .B(ori_ori_n585_), .Y(ori_ori_n598_));
  OR2        o0549(.A(x4), .B(x1), .Y(ori_ori_n599_));
  NO2        o0550(.A(ori_ori_n599_), .B(x3), .Y(ori_ori_n600_));
  NA2        o0551(.A(ori_ori_n55_), .B(x2), .Y(ori_ori_n601_));
  NO3        o0552(.A(ori_ori_n331_), .B(ori_ori_n601_), .C(x6), .Y(ori_ori_n602_));
  AOI220     o0553(.A0(ori_ori_n602_), .A1(ori_ori_n600_), .B0(ori_ori_n598_), .B1(ori_ori_n571_), .Y(ori06));
  NA2        o0554(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n604_));
  NA2        o0555(.A(x6), .B(ori_ori_n100_), .Y(ori_ori_n605_));
  NA2        o0556(.A(x5), .B(ori_ori_n57_), .Y(ori_ori_n606_));
  NA2        o0557(.A(ori_ori_n301_), .B(x2), .Y(ori_ori_n607_));
  NOi21      o0558(.An(x6), .B(x8), .Y(ori_ori_n608_));
  NA2        o0559(.A(ori_ori_n56_), .B(ori_ori_n50_), .Y(ori_ori_n609_));
  NO2        o0560(.A(ori_ori_n68_), .B(ori_ori_n98_), .Y(ori_ori_n610_));
  NO2        o0561(.A(ori_ori_n53_), .B(ori_ori_n57_), .Y(ori_ori_n611_));
  NO2        o0562(.A(ori_ori_n54_), .B(x0), .Y(ori_ori_n612_));
  NA2        o0563(.A(x4), .B(x3), .Y(ori_ori_n613_));
  NO2        o0564(.A(ori_ori_n94_), .B(ori_ori_n56_), .Y(ori_ori_n614_));
  NO2        o0565(.A(ori_ori_n366_), .B(x8), .Y(ori_ori_n615_));
  NO2        o0566(.A(x5), .B(x3), .Y(ori_ori_n616_));
  NA2        o0567(.A(x7), .B(ori_ori_n56_), .Y(ori_ori_n617_));
  NO2        o0568(.A(ori_ori_n544_), .B(ori_ori_n57_), .Y(ori_ori_n618_));
  NA2        o0569(.A(ori_ori_n618_), .B(ori_ori_n557_), .Y(ori_ori_n619_));
  NO2        o0570(.A(ori_ori_n154_), .B(x6), .Y(ori_ori_n620_));
  NA2        o0571(.A(ori_ori_n620_), .B(ori_ori_n261_), .Y(ori_ori_n621_));
  AOI210     o0572(.A0(ori_ori_n621_), .A1(ori_ori_n619_), .B0(ori_ori_n617_), .Y(ori_ori_n622_));
  AN2        o0573(.A(ori_ori_n413_), .B(ori_ori_n289_), .Y(ori_ori_n623_));
  OAI210     o0574(.A0(ori_ori_n623_), .A1(ori_ori_n622_), .B0(ori_ori_n312_), .Y(ori_ori_n624_));
  NO2        o0575(.A(ori_ori_n278_), .B(ori_ori_n98_), .Y(ori_ori_n625_));
  NO2        o0576(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n626_));
  NA2        o0577(.A(ori_ori_n626_), .B(ori_ori_n68_), .Y(ori_ori_n627_));
  NO2        o0578(.A(ori_ori_n627_), .B(ori_ori_n228_), .Y(ori_ori_n628_));
  NO2        o0579(.A(ori_ori_n68_), .B(x3), .Y(ori_ori_n629_));
  NA3        o0580(.A(ori_ori_n629_), .B(x1), .C(ori_ori_n56_), .Y(ori_ori_n630_));
  INV        o0581(.A(x6), .Y(ori_ori_n631_));
  NA2        o0582(.A(ori_ori_n163_), .B(ori_ori_n631_), .Y(ori_ori_n632_));
  NA3        o0583(.A(ori_ori_n531_), .B(x3), .C(ori_ori_n68_), .Y(ori_ori_n633_));
  NA3        o0584(.A(ori_ori_n633_), .B(ori_ori_n632_), .C(ori_ori_n630_), .Y(ori_ori_n634_));
  OR3        o0585(.A(ori_ori_n634_), .B(ori_ori_n628_), .C(ori_ori_n568_), .Y(ori_ori_n635_));
  NA2        o0586(.A(ori_ori_n635_), .B(ori_ori_n625_), .Y(ori_ori_n636_));
  NA2        o0587(.A(ori_ori_n612_), .B(ori_ori_n557_), .Y(ori_ori_n637_));
  NA4        o0588(.A(ori_ori_n238_), .B(ori_ori_n517_), .C(ori_ori_n200_), .D(ori_ori_n233_), .Y(ori_ori_n638_));
  NA2        o0589(.A(ori_ori_n420_), .B(ori_ori_n64_), .Y(ori_ori_n639_));
  AOI210     o0590(.A0(ori_ori_n638_), .A1(ori_ori_n637_), .B0(ori_ori_n639_), .Y(ori_ori_n640_));
  NA2        o0591(.A(x7), .B(x6), .Y(ori_ori_n641_));
  NA3        o0592(.A(x2), .B(x1), .C(x0), .Y(ori_ori_n642_));
  NO3        o0593(.A(ori_ori_n642_), .B(ori_ori_n641_), .C(ori_ori_n529_), .Y(ori_ori_n643_));
  NO2        o0594(.A(x5), .B(x1), .Y(ori_ori_n644_));
  NA2        o0595(.A(ori_ori_n644_), .B(ori_ori_n631_), .Y(ori_ori_n645_));
  NA2        o0596(.A(x4), .B(x0), .Y(ori_ori_n646_));
  NO2        o0597(.A(x6), .B(x2), .Y(ori_ori_n647_));
  NA2        o0598(.A(ori_ori_n647_), .B(ori_ori_n204_), .Y(ori_ori_n648_));
  NO2        o0599(.A(ori_ori_n648_), .B(ori_ori_n646_), .Y(ori_ori_n649_));
  NO3        o0600(.A(ori_ori_n649_), .B(ori_ori_n643_), .C(ori_ori_n640_), .Y(ori_ori_n650_));
  NA3        o0601(.A(ori_ori_n650_), .B(ori_ori_n636_), .C(ori_ori_n624_), .Y(ori_ori_n651_));
  INV        o0602(.A(ori_ori_n651_), .Y(ori07));
  NA2        o0603(.A(ori_ori_n98_), .B(ori_ori_n57_), .Y(ori_ori_n653_));
  NOi21      o0604(.An(ori_ori_n641_), .B(ori_ori_n105_), .Y(ori_ori_n654_));
  NO4        o0605(.A(ori_ori_n654_), .B(ori_ori_n557_), .C(ori_ori_n228_), .D(ori_ori_n653_), .Y(ori_ori_n655_));
  NO2        o0606(.A(x5), .B(x1), .Y(ori_ori_n656_));
  NA2        o0607(.A(ori_ori_n656_), .B(ori_ori_n337_), .Y(ori_ori_n657_));
  NA2        o0608(.A(x6), .B(ori_ori_n85_), .Y(ori_ori_n658_));
  OAI220     o0609(.A0(ori_ori_n658_), .A1(ori_ori_n123_), .B0(ori_ori_n657_), .B1(ori_ori_n291_), .Y(ori_ori_n659_));
  OAI210     o0610(.A0(ori_ori_n659_), .A1(ori_ori_n655_), .B0(x2), .Y(ori_ori_n660_));
  NAi21      o0611(.An(ori_ori_n142_), .B(ori_ori_n143_), .Y(ori_ori_n661_));
  NA3        o0612(.A(ori_ori_n661_), .B(ori_ori_n84_), .C(x3), .Y(ori_ori_n662_));
  INV        o0613(.A(ori_ori_n662_), .Y(ori_ori_n663_));
  NO2        o0614(.A(x8), .B(ori_ori_n53_), .Y(ori_ori_n664_));
  NA2        o0615(.A(ori_ori_n664_), .B(ori_ori_n57_), .Y(ori_ori_n665_));
  NO2        o0616(.A(x7), .B(x3), .Y(ori_ori_n666_));
  NA2        o0617(.A(ori_ori_n666_), .B(ori_ori_n92_), .Y(ori_ori_n667_));
  INV        o0618(.A(ori_ori_n667_), .Y(ori_ori_n668_));
  AOI210     o0619(.A0(ori_ori_n663_), .A1(ori_ori_n227_), .B0(ori_ori_n668_), .Y(ori_ori_n669_));
  AOI210     o0620(.A0(ori_ori_n669_), .A1(ori_ori_n660_), .B0(x4), .Y(ori_ori_n670_));
  NA3        o0621(.A(ori_ori_n644_), .B(ori_ori_n287_), .C(ori_ori_n55_), .Y(ori_ori_n671_));
  AOI210     o0622(.A0(ori_ori_n671_), .A1(ori_ori_n525_), .B0(ori_ori_n100_), .Y(ori_ori_n672_));
  XO2        o0623(.A(x5), .B(x1), .Y(ori_ori_n673_));
  NO4        o0624(.A(ori_ori_n673_), .B(ori_ori_n149_), .C(ori_ori_n188_), .D(ori_ori_n55_), .Y(ori_ori_n674_));
  OAI210     o0625(.A0(ori_ori_n674_), .A1(ori_ori_n672_), .B0(ori_ori_n368_), .Y(ori_ori_n675_));
  NO3        o0626(.A(ori_ori_n50_), .B(x2), .C(x0), .Y(ori_ori_n676_));
  NA2        o0627(.A(x6), .B(x0), .Y(ori_ori_n677_));
  NO2        o0628(.A(ori_ori_n601_), .B(ori_ori_n677_), .Y(ori_ori_n678_));
  INV        o0629(.A(ori_ori_n657_), .Y(ori_ori_n679_));
  NA2        o0630(.A(ori_ori_n679_), .B(ori_ori_n676_), .Y(ori_ori_n680_));
  AOI210     o0631(.A0(ori_ori_n680_), .A1(ori_ori_n675_), .B0(ori_ori_n56_), .Y(ori_ori_n681_));
  NOi21      o0632(.An(ori_ori_n211_), .B(ori_ori_n337_), .Y(ori_ori_n682_));
  NO3        o0633(.A(ori_ori_n682_), .B(ori_ori_n220_), .C(ori_ori_n64_), .Y(ori_ori_n683_));
  NO2        o0634(.A(ori_ori_n171_), .B(ori_ori_n68_), .Y(ori_ori_n684_));
  NO2        o0635(.A(ori_ori_n280_), .B(x6), .Y(ori_ori_n685_));
  AO220      o0636(.A0(ori_ori_n685_), .A1(ori_ori_n294_), .B0(ori_ori_n684_), .B1(ori_ori_n487_), .Y(ori_ori_n686_));
  OAI210     o0637(.A0(ori_ori_n686_), .A1(ori_ori_n683_), .B0(ori_ori_n57_), .Y(ori_ori_n687_));
  NA2        o0638(.A(ori_ori_n85_), .B(ori_ori_n68_), .Y(ori_ori_n688_));
  NAi21      o0639(.An(x8), .B(x7), .Y(ori_ori_n689_));
  NA2        o0640(.A(ori_ori_n682_), .B(ori_ori_n689_), .Y(ori_ori_n690_));
  NA2        o0641(.A(ori_ori_n363_), .B(ori_ori_n100_), .Y(ori_ori_n691_));
  NO2        o0642(.A(ori_ori_n608_), .B(x1), .Y(ori_ori_n692_));
  NO3        o0643(.A(ori_ori_n692_), .B(ori_ori_n691_), .C(x1), .Y(ori_ori_n693_));
  AOI210     o0644(.A0(ori_ori_n693_), .A1(ori_ori_n690_), .B0(ori_ori_n530_), .Y(ori_ori_n694_));
  AOI210     o0645(.A0(ori_ori_n694_), .A1(ori_ori_n687_), .B0(ori_ori_n130_), .Y(ori_ori_n695_));
  NO2        o0646(.A(x8), .B(x7), .Y(ori_ori_n696_));
  INV        o0647(.A(x3), .Y(ori_ori_n697_));
  NA3        o0648(.A(ori_ori_n697_), .B(ori_ori_n326_), .C(x1), .Y(ori_ori_n698_));
  NO2        o0649(.A(x8), .B(ori_ori_n100_), .Y(ori_ori_n699_));
  NA2        o0650(.A(x3), .B(ori_ori_n312_), .Y(ori_ori_n700_));
  NO2        o0651(.A(ori_ori_n68_), .B(x4), .Y(ori_ori_n701_));
  NA2        o0652(.A(ori_ori_n701_), .B(ori_ori_n275_), .Y(ori_ori_n702_));
  AOI210     o0653(.A0(ori_ori_n700_), .A1(ori_ori_n698_), .B0(ori_ori_n702_), .Y(ori_ori_n703_));
  NO4        o0654(.A(ori_ori_n703_), .B(ori_ori_n695_), .C(ori_ori_n681_), .D(ori_ori_n670_), .Y(ori08));
  NA2        o0655(.A(ori_ori_n50_), .B(x1), .Y(ori_ori_n705_));
  XN2        o0656(.A(x5), .B(x4), .Y(ori_ori_n706_));
  INV        o0657(.A(ori_ori_n706_), .Y(ori_ori_n707_));
  NO2        o0658(.A(ori_ori_n221_), .B(ori_ori_n98_), .Y(ori_ori_n708_));
  INV        o0659(.A(ori_ori_n244_), .Y(ori_ori_n709_));
  AOI210     o0660(.A0(ori_ori_n243_), .A1(ori_ori_n691_), .B0(ori_ori_n543_), .Y(ori_ori_n710_));
  NA2        o0661(.A(ori_ori_n538_), .B(ori_ori_n154_), .Y(ori_ori_n711_));
  OAI220     o0662(.A0(ori_ori_n711_), .A1(ori_ori_n586_), .B0(ori_ori_n422_), .B1(ori_ori_n50_), .Y(ori_ori_n712_));
  AO210      o0663(.A0(ori_ori_n712_), .A1(ori_ori_n305_), .B0(ori_ori_n710_), .Y(ori_ori_n713_));
  NA2        o0664(.A(ori_ori_n249_), .B(ori_ori_n136_), .Y(ori_ori_n714_));
  NA2        o0665(.A(ori_ori_n130_), .B(x7), .Y(ori_ori_n715_));
  OR3        o0666(.A(ori_ori_n642_), .B(ori_ori_n410_), .C(ori_ori_n616_), .Y(ori_ori_n716_));
  OAI220     o0667(.A0(ori_ori_n716_), .A1(ori_ori_n715_), .B0(ori_ori_n714_), .B1(ori_ori_n185_), .Y(ori_ori_n717_));
  AOI210     o0668(.A0(ori_ori_n713_), .A1(ori_ori_n263_), .B0(ori_ori_n717_), .Y(ori_ori_n718_));
  AOI210     o0669(.A0(ori_ori_n718_), .A1(ori_ori_n709_), .B0(ori_ori_n68_), .Y(ori_ori_n719_));
  NO2        o0670(.A(ori_ori_n696_), .B(ori_ori_n100_), .Y(ori_ori_n720_));
  NA2        o0671(.A(ori_ori_n720_), .B(ori_ori_n173_), .Y(ori_ori_n721_));
  OAI210     o0672(.A0(ori_ori_n366_), .A1(ori_ori_n275_), .B0(ori_ori_n305_), .Y(ori_ori_n722_));
  NA2        o0673(.A(ori_ori_n615_), .B(ori_ori_n97_), .Y(ori_ori_n723_));
  OAI220     o0674(.A0(ori_ori_n723_), .A1(ori_ori_n2178_), .B0(ori_ori_n722_), .B1(ori_ori_n721_), .Y(ori_ori_n724_));
  NA2        o0675(.A(ori_ori_n724_), .B(ori_ori_n259_), .Y(ori_ori_n725_));
  NO3        o0676(.A(ori_ori_n366_), .B(ori_ori_n123_), .C(ori_ori_n65_), .Y(ori_ori_n726_));
  NO2        o0677(.A(ori_ori_n611_), .B(ori_ori_n223_), .Y(ori_ori_n727_));
  NO3        o0678(.A(ori_ori_n496_), .B(ori_ori_n411_), .C(ori_ori_n90_), .Y(ori_ori_n728_));
  AO220      o0679(.A0(ori_ori_n728_), .A1(ori_ori_n727_), .B0(ori_ori_n726_), .B1(x1), .Y(ori_ori_n729_));
  NA2        o0680(.A(x7), .B(ori_ori_n57_), .Y(ori_ori_n730_));
  NO3        o0681(.A(ori_ori_n282_), .B(ori_ori_n730_), .C(ori_ori_n258_), .Y(ori_ori_n731_));
  AOI210     o0682(.A0(ori_ori_n729_), .A1(x5), .B0(ori_ori_n731_), .Y(ori_ori_n732_));
  AOI210     o0683(.A0(ori_ori_n732_), .A1(ori_ori_n725_), .B0(ori_ori_n69_), .Y(ori_ori_n733_));
  NO2        o0684(.A(ori_ori_n67_), .B(x3), .Y(ori_ori_n734_));
  NA2        o0685(.A(ori_ori_n734_), .B(ori_ori_n134_), .Y(ori_ori_n735_));
  MUX2       o0686(.S(x3), .A(ori_ori_n149_), .B(ori_ori_n661_), .Y(ori_ori_n736_));
  NA2        o0687(.A(ori_ori_n736_), .B(ori_ori_n487_), .Y(ori_ori_n737_));
  NO3        o0688(.A(x6), .B(x4), .C(x0), .Y(ori_ori_n738_));
  INV        o0689(.A(ori_ori_n738_), .Y(ori_ori_n739_));
  AOI210     o0690(.A0(ori_ori_n737_), .A1(ori_ori_n735_), .B0(ori_ori_n739_), .Y(ori_ori_n740_));
  NO3        o0691(.A(x5), .B(x3), .C(ori_ori_n100_), .Y(ori_ori_n741_));
  OR2        o0692(.A(x8), .B(x1), .Y(ori_ori_n742_));
  NO2        o0693(.A(ori_ori_n742_), .B(ori_ori_n626_), .Y(ori_ori_n743_));
  NAi21      o0694(.An(x4), .B(x1), .Y(ori_ori_n744_));
  NO2        o0695(.A(ori_ori_n744_), .B(x0), .Y(ori_ori_n745_));
  NA2        o0696(.A(ori_ori_n537_), .B(ori_ori_n745_), .Y(ori_ori_n746_));
  NA3        o0697(.A(ori_ori_n55_), .B(x1), .C(x0), .Y(ori_ori_n747_));
  OAI210     o0698(.A0(ori_ori_n747_), .A1(ori_ori_n341_), .B0(ori_ori_n746_), .Y(ori_ori_n748_));
  OAI210     o0699(.A0(ori_ori_n748_), .A1(ori_ori_n743_), .B0(ori_ori_n287_), .Y(ori_ori_n749_));
  NA2        o0700(.A(ori_ori_n98_), .B(ori_ori_n56_), .Y(ori_ori_n750_));
  NO2        o0701(.A(ori_ori_n750_), .B(ori_ori_n235_), .Y(ori_ori_n751_));
  INV        o0702(.A(x2), .Y(ori_ori_n752_));
  NO4        o0703(.A(ori_ori_n294_), .B(ori_ori_n752_), .C(ori_ori_n696_), .D(ori_ori_n265_), .Y(ori_ori_n753_));
  AOI220     o0704(.A0(ori_ori_n753_), .A1(ori_ori_n751_), .B0(ori_ori_n625_), .B1(ori_ori_n568_), .Y(ori_ori_n754_));
  NA2        o0705(.A(ori_ori_n754_), .B(ori_ori_n749_), .Y(ori_ori_n755_));
  NO4        o0706(.A(ori_ori_n755_), .B(ori_ori_n740_), .C(ori_ori_n733_), .D(ori_ori_n719_), .Y(ori09));
  NO3        o0707(.A(ori_ori_n673_), .B(ori_ori_n109_), .C(ori_ori_n87_), .Y(ori_ori_n757_));
  AOI220     o0708(.A0(ori_ori_n270_), .A1(ori_ori_n67_), .B0(ori_ori_n516_), .B1(ori_ori_n471_), .Y(ori_ori_n758_));
  OAI210     o0709(.A0(ori_ori_n757_), .A1(x2), .B0(ori_ori_n758_), .Y(ori_ori_n759_));
  AOI210     o0710(.A0(ori_ori_n759_), .A1(ori_ori_n645_), .B0(ori_ori_n393_), .Y(ori_ori_n760_));
  NO2        o0711(.A(ori_ori_n644_), .B(ori_ori_n301_), .Y(ori_ori_n761_));
  NO3        o0712(.A(ori_ori_n530_), .B(ori_ori_n93_), .C(ori_ori_n100_), .Y(ori_ori_n762_));
  AN2        o0713(.A(ori_ori_n762_), .B(ori_ori_n761_), .Y(ori_ori_n763_));
  OAI210     o0714(.A0(ori_ori_n763_), .A1(ori_ori_n760_), .B0(x4), .Y(ori_ori_n764_));
  OAI220     o0715(.A0(ori_ori_n329_), .A1(ori_ori_n132_), .B0(ori_ori_n352_), .B1(ori_ori_n251_), .Y(ori_ori_n765_));
  NO2        o0716(.A(ori_ori_n171_), .B(ori_ori_n98_), .Y(ori_ori_n766_));
  AOI220     o0717(.A0(ori_ori_n766_), .A1(ori_ori_n114_), .B0(ori_ori_n765_), .B1(ori_ori_n550_), .Y(ori_ori_n767_));
  NO2        o0718(.A(ori_ori_n673_), .B(ori_ori_n87_), .Y(ori_ori_n768_));
  NAi21      o0719(.An(x0), .B(x2), .Y(ori_ori_n769_));
  NO2        o0720(.A(ori_ori_n274_), .B(ori_ori_n769_), .Y(ori_ori_n770_));
  OAI210     o0721(.A0(ori_ori_n414_), .A1(ori_ori_n246_), .B0(ori_ori_n171_), .Y(ori_ori_n771_));
  AOI210     o0722(.A0(ori_ori_n151_), .A1(ori_ori_n689_), .B0(ori_ori_n317_), .Y(ori_ori_n772_));
  AOI220     o0723(.A0(ori_ori_n772_), .A1(ori_ori_n771_), .B0(ori_ori_n770_), .B1(ori_ori_n768_), .Y(ori_ori_n773_));
  OAI210     o0724(.A0(ori_ori_n767_), .A1(ori_ori_n55_), .B0(ori_ori_n773_), .Y(ori_ori_n774_));
  NA2        o0725(.A(ori_ori_n774_), .B(ori_ori_n56_), .Y(ori_ori_n775_));
  NO2        o0726(.A(ori_ori_n56_), .B(ori_ori_n57_), .Y(ori_ori_n776_));
  INV        o0727(.A(ori_ori_n114_), .Y(ori_ori_n777_));
  NA2        o0728(.A(ori_ori_n644_), .B(ori_ori_n55_), .Y(ori_ori_n778_));
  AOI210     o0729(.A0(x6), .A1(x1), .B0(x5), .Y(ori_ori_n779_));
  OAI210     o0730(.A0(ori_ori_n779_), .A1(ori_ori_n297_), .B0(x2), .Y(ori_ori_n780_));
  AOI210     o0731(.A0(ori_ori_n780_), .A1(ori_ori_n778_), .B0(ori_ori_n777_), .Y(ori_ori_n781_));
  NA2        o0732(.A(ori_ori_n486_), .B(ori_ori_n55_), .Y(ori_ori_n782_));
  NO2        o0733(.A(ori_ori_n210_), .B(ori_ori_n343_), .Y(ori_ori_n783_));
  NO2        o0734(.A(ori_ori_n280_), .B(ori_ori_n135_), .Y(ori_ori_n784_));
  NO2        o0735(.A(ori_ori_n784_), .B(ori_ori_n783_), .Y(ori_ori_n785_));
  NO2        o0736(.A(ori_ori_n785_), .B(ori_ori_n55_), .Y(ori_ori_n786_));
  OAI210     o0737(.A0(ori_ori_n786_), .A1(ori_ori_n781_), .B0(ori_ori_n776_), .Y(ori_ori_n787_));
  NO2        o0738(.A(ori_ori_n361_), .B(ori_ori_n98_), .Y(ori_ori_n788_));
  NA2        o0739(.A(ori_ori_n189_), .B(ori_ori_n208_), .Y(ori_ori_n789_));
  NA4        o0740(.A(ori_ori_n789_), .B(ori_ori_n787_), .C(ori_ori_n775_), .D(ori_ori_n764_), .Y(ori_ori_n790_));
  NA2        o0741(.A(ori_ori_n790_), .B(ori_ori_n50_), .Y(ori_ori_n791_));
  NO2        o0742(.A(ori_ori_n339_), .B(ori_ori_n146_), .Y(ori_ori_n792_));
  OAI210     o0743(.A0(x1), .A1(ori_ori_n699_), .B0(ori_ori_n2176_), .Y(ori_ori_n793_));
  OAI210     o0744(.A0(ori_ori_n793_), .A1(ori_ori_n792_), .B0(x0), .Y(ori_ori_n794_));
  NO3        o0745(.A(x8), .B(x7), .C(x2), .Y(ori_ori_n795_));
  NO2        o0746(.A(x5), .B(x2), .Y(ori_ori_n796_));
  OAI210     o0747(.A0(ori_ori_n796_), .A1(ori_ori_n795_), .B0(ori_ori_n452_), .Y(ori_ori_n797_));
  AOI210     o0748(.A0(ori_ori_n797_), .A1(ori_ori_n794_), .B0(x4), .Y(ori_ori_n798_));
  NO2        o0749(.A(ori_ori_n376_), .B(ori_ori_n134_), .Y(ori_ori_n799_));
  NO2        o0750(.A(ori_ori_n52_), .B(x2), .Y(ori_ori_n800_));
  NO2        o0751(.A(ori_ori_n98_), .B(ori_ori_n56_), .Y(ori_ori_n801_));
  NA2        o0752(.A(ori_ori_n801_), .B(x8), .Y(ori_ori_n802_));
  NA2        o0753(.A(ori_ori_n802_), .B(ori_ori_n778_), .Y(ori_ori_n803_));
  AO210      o0754(.A0(ori_ori_n803_), .A1(ori_ori_n800_), .B0(ori_ori_n799_), .Y(ori_ori_n804_));
  OAI210     o0755(.A0(ori_ori_n804_), .A1(ori_ori_n798_), .B0(ori_ori_n542_), .Y(ori_ori_n805_));
  NO2        o0756(.A(ori_ori_n234_), .B(ori_ori_n108_), .Y(ori_ori_n806_));
  OAI210     o0757(.A0(x4), .A1(x2), .B0(x0), .Y(ori_ori_n807_));
  NA3        o0758(.A(ori_ori_n532_), .B(ori_ori_n543_), .C(ori_ori_n306_), .Y(ori_ori_n808_));
  OAI210     o0759(.A0(ori_ori_n807_), .A1(ori_ori_n258_), .B0(ori_ori_n53_), .Y(ori_ori_n809_));
  AOI210     o0760(.A0(ori_ori_n808_), .A1(ori_ori_n807_), .B0(ori_ori_n809_), .Y(ori_ori_n810_));
  OAI210     o0761(.A0(ori_ori_n810_), .A1(ori_ori_n806_), .B0(x3), .Y(ori_ori_n811_));
  NA2        o0762(.A(ori_ori_n363_), .B(ori_ori_n661_), .Y(ori_ori_n812_));
  NA2        o0763(.A(ori_ori_n227_), .B(ori_ori_n149_), .Y(ori_ori_n813_));
  AO210      o0764(.A0(ori_ori_n813_), .A1(ori_ori_n812_), .B0(ori_ori_n121_), .Y(ori_ori_n814_));
  NO2        o0765(.A(ori_ori_n387_), .B(x2), .Y(ori_ori_n815_));
  NO2        o0766(.A(x7), .B(ori_ori_n53_), .Y(ori_ori_n816_));
  NA2        o0767(.A(ori_ori_n589_), .B(ori_ori_n222_), .Y(ori_ori_n817_));
  NA3        o0768(.A(ori_ori_n817_), .B(ori_ori_n814_), .C(ori_ori_n811_), .Y(ori_ori_n818_));
  AOI220     o0769(.A0(ori_ori_n531_), .A1(ori_ori_n530_), .B0(ori_ori_n252_), .B1(x5), .Y(ori_ori_n819_));
  NO2        o0770(.A(ori_ori_n594_), .B(ori_ori_n171_), .Y(ori_ori_n820_));
  NA3        o0771(.A(ori_ori_n820_), .B(ori_ori_n590_), .C(x7), .Y(ori_ori_n821_));
  OAI210     o0772(.A0(ori_ori_n819_), .A1(ori_ori_n311_), .B0(ori_ori_n821_), .Y(ori_ori_n822_));
  NA2        o0773(.A(ori_ori_n822_), .B(ori_ori_n79_), .Y(ori_ori_n823_));
  NO2        o0774(.A(x5), .B(ori_ori_n53_), .Y(ori_ori_n824_));
  NAi21      o0775(.An(x1), .B(x4), .Y(ori_ori_n825_));
  NA2        o0776(.A(ori_ori_n825_), .B(ori_ori_n744_), .Y(ori_ori_n826_));
  NO3        o0777(.A(ori_ori_n826_), .B(ori_ori_n182_), .C(ori_ori_n824_), .Y(ori_ori_n827_));
  NA2        o0778(.A(ori_ori_n827_), .B(ori_ori_n368_), .Y(ori_ori_n828_));
  NA2        o0779(.A(ori_ori_n828_), .B(ori_ori_n823_), .Y(ori_ori_n829_));
  AOI210     o0780(.A0(ori_ori_n818_), .A1(x6), .B0(ori_ori_n829_), .Y(ori_ori_n830_));
  NA3        o0781(.A(ori_ori_n830_), .B(ori_ori_n805_), .C(ori_ori_n791_), .Y(ori10));
  NO2        o0782(.A(x4), .B(x1), .Y(ori_ori_n832_));
  NO2        o0783(.A(ori_ori_n832_), .B(ori_ori_n136_), .Y(ori_ori_n833_));
  NA3        o0784(.A(x5), .B(x4), .C(x0), .Y(ori_ori_n834_));
  OAI220     o0785(.A0(ori_ori_n834_), .A1(ori_ori_n247_), .B0(ori_ori_n611_), .B1(ori_ori_n225_), .Y(ori_ori_n835_));
  NA2        o0786(.A(ori_ori_n835_), .B(ori_ori_n833_), .Y(ori_ori_n836_));
  NO3        o0787(.A(ori_ori_n318_), .B(ori_ori_n288_), .C(ori_ori_n85_), .Y(ori_ori_n837_));
  NA3        o0788(.A(ori_ori_n837_), .B(ori_ori_n341_), .C(ori_ori_n60_), .Y(ori_ori_n838_));
  AOI210     o0789(.A0(ori_ori_n838_), .A1(ori_ori_n836_), .B0(ori_ori_n274_), .Y(ori_ori_n839_));
  NOi21      o0790(.An(ori_ori_n233_), .B(ori_ori_n126_), .Y(ori_ori_n840_));
  AOI210     o0791(.A0(ori_ori_n438_), .A1(ori_ori_n544_), .B0(ori_ori_n294_), .Y(ori_ori_n841_));
  NO2        o0792(.A(ori_ori_n776_), .B(ori_ori_n304_), .Y(ori_ori_n842_));
  NOi31      o0793(.An(ori_ori_n842_), .B(ori_ori_n841_), .C(ori_ori_n840_), .Y(ori_ori_n843_));
  NA2        o0794(.A(x4), .B(ori_ori_n100_), .Y(ori_ori_n844_));
  NO2        o0795(.A(ori_ori_n291_), .B(ori_ori_n844_), .Y(ori_ori_n845_));
  NA2        o0796(.A(ori_ori_n90_), .B(x5), .Y(ori_ori_n846_));
  NO3        o0797(.A(ori_ori_n846_), .B(ori_ori_n101_), .C(ori_ori_n55_), .Y(ori_ori_n847_));
  NO3        o0798(.A(ori_ori_n847_), .B(ori_ori_n845_), .C(ori_ori_n843_), .Y(ori_ori_n848_));
  NA2        o0799(.A(ori_ori_n824_), .B(ori_ori_n50_), .Y(ori_ori_n849_));
  NA2        o0800(.A(ori_ori_n531_), .B(ori_ori_n242_), .Y(ori_ori_n850_));
  NO2        o0801(.A(ori_ori_n850_), .B(ori_ori_n849_), .Y(ori_ori_n851_));
  OAI220     o0802(.A0(ori_ori_n802_), .A1(ori_ori_n97_), .B0(ori_ori_n750_), .B1(ori_ori_n393_), .Y(ori_ori_n852_));
  AOI210     o0803(.A0(ori_ori_n852_), .A1(ori_ori_n249_), .B0(ori_ori_n851_), .Y(ori_ori_n853_));
  OAI210     o0804(.A0(ori_ori_n848_), .A1(ori_ori_n343_), .B0(ori_ori_n853_), .Y(ori_ori_n854_));
  OAI210     o0805(.A0(ori_ori_n854_), .A1(ori_ori_n839_), .B0(x7), .Y(ori_ori_n855_));
  NA2        o0806(.A(ori_ori_n55_), .B(ori_ori_n68_), .Y(ori_ori_n856_));
  NO3        o0807(.A(ori_ori_n395_), .B(ori_ori_n769_), .C(x5), .Y(ori_ori_n857_));
  NO2        o0808(.A(ori_ori_n318_), .B(ori_ori_n129_), .Y(ori_ori_n858_));
  NO2        o0809(.A(x5), .B(ori_ori_n100_), .Y(ori_ori_n859_));
  NA3        o0810(.A(ori_ori_n407_), .B(ori_ori_n120_), .C(ori_ori_n377_), .Y(ori_ori_n860_));
  OAI210     o0811(.A0(ori_ori_n395_), .A1(ori_ori_n193_), .B0(ori_ori_n860_), .Y(ori_ori_n861_));
  NO2        o0812(.A(ori_ori_n231_), .B(ori_ori_n861_), .Y(ori_ori_n862_));
  NO2        o0813(.A(ori_ori_n862_), .B(ori_ori_n57_), .Y(ori_ori_n863_));
  OAI210     o0814(.A0(ori_ori_n863_), .A1(ori_ori_n857_), .B0(ori_ori_n816_), .Y(ori_ori_n864_));
  NO2        o0815(.A(x4), .B(x3), .Y(ori_ori_n865_));
  NO3        o0816(.A(ori_ori_n865_), .B(ori_ori_n305_), .C(ori_ori_n83_), .Y(ori_ori_n866_));
  OAI210     o0817(.A0(ori_ori_n866_), .A1(ori_ori_n248_), .B0(ori_ori_n386_), .Y(ori_ori_n867_));
  AOI210     o0818(.A0(ori_ori_n356_), .A1(ori_ori_n117_), .B0(ori_ori_n228_), .Y(ori_ori_n868_));
  NA2        o0819(.A(ori_ori_n832_), .B(ori_ori_n55_), .Y(ori_ori_n869_));
  NO2        o0820(.A(ori_ori_n869_), .B(ori_ori_n846_), .Y(ori_ori_n870_));
  NO2        o0821(.A(ori_ori_n458_), .B(ori_ori_n323_), .Y(ori_ori_n871_));
  NO3        o0822(.A(x4), .B(ori_ori_n100_), .C(ori_ori_n57_), .Y(ori_ori_n872_));
  NO2        o0823(.A(ori_ori_n387_), .B(x1), .Y(ori_ori_n873_));
  NOi31      o0824(.An(ori_ori_n872_), .B(ori_ori_n873_), .C(ori_ori_n871_), .Y(ori_ori_n874_));
  NA2        o0825(.A(ori_ori_n55_), .B(x5), .Y(ori_ori_n875_));
  NO4        o0826(.A(ori_ori_n833_), .B(ori_ori_n451_), .C(ori_ori_n875_), .D(x2), .Y(ori_ori_n876_));
  NO4        o0827(.A(ori_ori_n876_), .B(ori_ori_n874_), .C(ori_ori_n870_), .D(ori_ori_n868_), .Y(ori_ori_n877_));
  AOI210     o0828(.A0(ori_ori_n877_), .A1(ori_ori_n867_), .B0(ori_ori_n188_), .Y(ori_ori_n878_));
  NO2        o0829(.A(x6), .B(x2), .Y(ori_ori_n879_));
  NO2        o0830(.A(ori_ori_n750_), .B(ori_ori_n393_), .Y(ori_ori_n880_));
  NA3        o0831(.A(x4), .B(x3), .C(ori_ori_n100_), .Y(ori_ori_n881_));
  NO2        o0832(.A(ori_ori_n55_), .B(ori_ori_n56_), .Y(ori_ori_n882_));
  NOi21      o0833(.An(ori_ori_n112_), .B(ori_ori_n111_), .Y(ori_ori_n883_));
  NO3        o0834(.A(ori_ori_n306_), .B(ori_ori_n291_), .C(ori_ori_n883_), .Y(ori_ori_n884_));
  NA2        o0835(.A(ori_ori_n884_), .B(ori_ori_n230_), .Y(ori_ori_n885_));
  NO2        o0836(.A(ori_ori_n885_), .B(ori_ori_n882_), .Y(ori_ori_n886_));
  NA2        o0837(.A(ori_ori_n455_), .B(ori_ori_n235_), .Y(ori_ori_n887_));
  NO2        o0838(.A(ori_ori_n422_), .B(ori_ori_n515_), .Y(ori_ori_n888_));
  NO2        o0839(.A(ori_ori_n164_), .B(ori_ori_n100_), .Y(ori_ori_n889_));
  NA3        o0840(.A(ori_ori_n889_), .B(ori_ori_n163_), .C(ori_ori_n111_), .Y(ori_ori_n890_));
  INV        o0841(.A(ori_ori_n890_), .Y(ori_ori_n891_));
  NO3        o0842(.A(ori_ori_n891_), .B(ori_ori_n886_), .C(ori_ori_n878_), .Y(ori_ori_n892_));
  NA3        o0843(.A(ori_ori_n892_), .B(ori_ori_n864_), .C(ori_ori_n855_), .Y(ori11));
  NO2        o0844(.A(ori_ori_n661_), .B(x5), .Y(ori_ori_n894_));
  NO2        o0845(.A(ori_ori_n302_), .B(ori_ori_n378_), .Y(ori_ori_n895_));
  NO2        o0846(.A(ori_ori_n55_), .B(ori_ori_n98_), .Y(ori_ori_n896_));
  NO2        o0847(.A(ori_ori_n68_), .B(x1), .Y(ori_ori_n897_));
  NA2        o0848(.A(ori_ori_n897_), .B(ori_ori_n75_), .Y(ori_ori_n898_));
  NO2        o0849(.A(ori_ori_n386_), .B(x3), .Y(ori_ori_n899_));
  NA2        o0850(.A(ori_ori_n100_), .B(x1), .Y(ori_ori_n900_));
  NO2        o0851(.A(ori_ori_n544_), .B(ori_ori_n199_), .Y(ori_ori_n901_));
  NA3        o0852(.A(x6), .B(x5), .C(ori_ori_n100_), .Y(ori_ori_n902_));
  NO2        o0853(.A(ori_ori_n902_), .B(ori_ori_n247_), .Y(ori_ori_n903_));
  NO2        o0854(.A(ori_ori_n395_), .B(x0), .Y(ori_ori_n904_));
  NA2        o0855(.A(ori_ori_n742_), .B(ori_ori_n83_), .Y(ori_ori_n905_));
  NO3        o0856(.A(ori_ori_n408_), .B(ori_ori_n664_), .C(ori_ori_n112_), .Y(ori_ori_n906_));
  AOI210     o0857(.A0(ori_ori_n905_), .A1(ori_ori_n92_), .B0(ori_ori_n906_), .Y(ori_ori_n907_));
  NO2        o0858(.A(x8), .B(x1), .Y(ori_ori_n908_));
  NO3        o0859(.A(ori_ori_n908_), .B(ori_ori_n604_), .C(ori_ori_n397_), .Y(ori_ori_n909_));
  OAI210     o0860(.A0(ori_ori_n74_), .A1(ori_ori_n53_), .B0(ori_ori_n909_), .Y(ori_ori_n910_));
  OAI210     o0861(.A0(ori_ori_n907_), .A1(x3), .B0(ori_ori_n910_), .Y(ori_ori_n911_));
  NO2        o0862(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n912_));
  OAI210     o0863(.A0(ori_ori_n912_), .A1(x2), .B0(ori_ori_n213_), .Y(ori_ori_n913_));
  NO2        o0864(.A(ori_ori_n532_), .B(ori_ori_n211_), .Y(ori_ori_n914_));
  NA2        o0865(.A(ori_ori_n914_), .B(ori_ori_n913_), .Y(ori_ori_n915_));
  NO2        o0866(.A(ori_ori_n455_), .B(x4), .Y(ori_ori_n916_));
  NO3        o0867(.A(ori_ori_n55_), .B(x6), .C(x1), .Y(ori_ori_n917_));
  NOi21      o0868(.An(ori_ori_n917_), .B(ori_ori_n422_), .Y(ori_ori_n918_));
  AOI210     o0869(.A0(ori_ori_n916_), .A1(ori_ori_n505_), .B0(ori_ori_n918_), .Y(ori_ori_n919_));
  NA2        o0870(.A(ori_ori_n919_), .B(ori_ori_n915_), .Y(ori_ori_n920_));
  AOI210     o0871(.A0(ori_ori_n911_), .A1(x2), .B0(ori_ori_n920_), .Y(ori_ori_n921_));
  NO2        o0872(.A(ori_ori_n211_), .B(x2), .Y(ori_ori_n922_));
  NA2        o0873(.A(ori_ori_n922_), .B(ori_ori_n865_), .Y(ori_ori_n923_));
  NOi21      o0874(.An(ori_ori_n345_), .B(ori_ori_n495_), .Y(ori_ori_n924_));
  NO3        o0875(.A(ori_ori_n924_), .B(ori_ori_n531_), .C(ori_ori_n291_), .Y(ori_ori_n925_));
  NA2        o0876(.A(x8), .B(ori_ori_n100_), .Y(ori_ori_n926_));
  OAI220     o0877(.A0(ori_ori_n613_), .A1(ori_ori_n926_), .B0(ori_ori_n291_), .B1(ori_ori_n341_), .Y(ori_ori_n927_));
  OAI210     o0878(.A0(ori_ori_n927_), .A1(ori_ori_n925_), .B0(ori_ori_n68_), .Y(ori_ori_n928_));
  NO2        o0879(.A(ori_ori_n98_), .B(x1), .Y(ori_ori_n929_));
  NA2        o0880(.A(ori_ori_n929_), .B(x7), .Y(ori_ori_n930_));
  AOI210     o0881(.A0(ori_ori_n928_), .A1(ori_ori_n923_), .B0(ori_ori_n930_), .Y(ori_ori_n931_));
  NA2        o0882(.A(ori_ori_n81_), .B(ori_ori_n68_), .Y(ori_ori_n932_));
  INV        o0883(.A(ori_ori_n226_), .Y(ori_ori_n933_));
  NA2        o0884(.A(ori_ori_n933_), .B(ori_ori_n136_), .Y(ori_ori_n934_));
  OAI220     o0885(.A0(ori_ori_n934_), .A1(ori_ori_n327_), .B0(ori_ori_n932_), .B1(ori_ori_n291_), .Y(ori_ori_n935_));
  NO2        o0886(.A(ori_ori_n145_), .B(ori_ori_n55_), .Y(ori_ori_n936_));
  AOI210     o0887(.A0(ori_ori_n936_), .A1(ori_ori_n935_), .B0(ori_ori_n931_), .Y(ori_ori_n937_));
  OAI210     o0888(.A0(ori_ori_n921_), .A1(ori_ori_n730_), .B0(ori_ori_n937_), .Y(ori12));
  NA2        o0889(.A(ori_ori_n2187_), .B(ori_ori_n248_), .Y(ori_ori_n939_));
  INV        o0890(.A(ori_ori_n939_), .Y(ori_ori_n940_));
  NOi21      o0891(.An(ori_ori_n361_), .B(ori_ori_n482_), .Y(ori_ori_n941_));
  NO2        o0892(.A(x7), .B(ori_ori_n50_), .Y(ori_ori_n942_));
  INV        o0893(.A(ori_ori_n532_), .Y(ori_ori_n943_));
  NA2        o0894(.A(ori_ori_n943_), .B(ori_ori_n873_), .Y(ori_ori_n944_));
  NA2        o0895(.A(ori_ori_n896_), .B(ori_ori_n56_), .Y(ori_ori_n945_));
  OAI220     o0896(.A0(ori_ori_n945_), .A1(ori_ori_n506_), .B0(ori_ori_n944_), .B1(ori_ori_n941_), .Y(ori_ori_n946_));
  OAI210     o0897(.A0(ori_ori_n946_), .A1(ori_ori_n940_), .B0(ori_ori_n510_), .Y(ori_ori_n947_));
  NA2        o0898(.A(ori_ori_n83_), .B(x5), .Y(ori_ori_n948_));
  NA2        o0899(.A(ori_ori_n258_), .B(ori_ori_n50_), .Y(ori_ori_n949_));
  NO2        o0900(.A(ori_ori_n905_), .B(ori_ori_n450_), .Y(ori_ori_n950_));
  NO3        o0901(.A(ori_ori_n219_), .B(ori_ori_n241_), .C(ori_ori_n58_), .Y(ori_ori_n951_));
  AOI220     o0902(.A0(ori_ori_n951_), .A1(ori_ori_n950_), .B0(ori_ori_n530_), .B1(ori_ori_n56_), .Y(ori_ori_n952_));
  INV        o0903(.A(ori_ori_n952_), .Y(ori_ori_n953_));
  INV        o0904(.A(x0), .Y(ori_ori_n954_));
  NO2        o0905(.A(ori_ori_n586_), .B(ori_ori_n288_), .Y(ori_ori_n955_));
  NO2        o0906(.A(ori_ori_n646_), .B(x3), .Y(ori_ori_n956_));
  NA2        o0907(.A(ori_ori_n955_), .B(ori_ori_n954_), .Y(ori_ori_n957_));
  NO3        o0908(.A(ori_ori_n2170_), .B(ori_ori_n533_), .C(x8), .Y(ori_ori_n958_));
  NA4        o0909(.A(ori_ori_n588_), .B(ori_ori_n582_), .C(ori_ori_n185_), .D(x0), .Y(ori_ori_n959_));
  OAI220     o0910(.A0(ori_ori_n959_), .A1(ori_ori_n958_), .B0(ori_ori_n957_), .B1(ori_ori_n504_), .Y(ori_ori_n960_));
  AOI210     o0911(.A0(ori_ori_n953_), .A1(ori_ori_n879_), .B0(ori_ori_n960_), .Y(ori_ori_n961_));
  NO2        o0912(.A(ori_ori_n225_), .B(ori_ori_n55_), .Y(ori_ori_n962_));
  NOi32      o0913(.An(ori_ori_n2182_), .Bn(ori_ori_n184_), .C(ori_ori_n496_), .Y(ori_ori_n963_));
  NO2        o0914(.A(ori_ori_n2164_), .B(ori_ori_n58_), .Y(ori_ori_n964_));
  OAI210     o0915(.A0(ori_ori_n963_), .A1(ori_ori_n962_), .B0(ori_ori_n964_), .Y(ori_ori_n965_));
  NO2        o0916(.A(ori_ori_n816_), .B(ori_ori_n91_), .Y(ori_ori_n966_));
  NO2        o0917(.A(ori_ori_n151_), .B(ori_ori_n53_), .Y(ori_ori_n967_));
  AOI210     o0918(.A0(ori_ori_n302_), .A1(x8), .B0(ori_ori_n967_), .Y(ori_ori_n968_));
  AOI210     o0919(.A0(ori_ori_n196_), .A1(ori_ori_n87_), .B0(ori_ori_n968_), .Y(ori_ori_n969_));
  OAI210     o0920(.A0(ori_ori_n969_), .A1(ori_ori_n966_), .B0(ori_ori_n594_), .Y(ori_ori_n970_));
  NO2        o0921(.A(x7), .B(x0), .Y(ori_ori_n971_));
  NO3        o0922(.A(ori_ori_n145_), .B(ori_ori_n971_), .C(ori_ori_n133_), .Y(ori_ori_n972_));
  XN2        o0923(.A(x8), .B(x7), .Y(ori_ori_n973_));
  NO3        o0924(.A(ori_ori_n908_), .B(ori_ori_n233_), .C(ori_ori_n973_), .Y(ori_ori_n974_));
  OAI210     o0925(.A0(ori_ori_n974_), .A1(ori_ori_n972_), .B0(ori_ori_n626_), .Y(ori_ori_n975_));
  NO2        o0926(.A(ori_ori_n98_), .B(x4), .Y(ori_ori_n976_));
  NA2        o0927(.A(ori_ori_n248_), .B(ori_ori_n976_), .Y(ori_ori_n977_));
  NA4        o0928(.A(ori_ori_n977_), .B(ori_ori_n975_), .C(ori_ori_n970_), .D(ori_ori_n965_), .Y(ori_ori_n978_));
  NA2        o0929(.A(ori_ori_n978_), .B(ori_ori_n486_), .Y(ori_ori_n979_));
  NO2        o0930(.A(ori_ori_n55_), .B(x4), .Y(ori_ori_n980_));
  NA2        o0931(.A(ori_ori_n980_), .B(ori_ori_n148_), .Y(ori_ori_n981_));
  NO2        o0932(.A(ori_ori_n590_), .B(ori_ori_n233_), .Y(ori_ori_n982_));
  OAI210     o0933(.A0(ori_ori_n982_), .A1(ori_ori_n880_), .B0(ori_ori_n50_), .Y(ori_ori_n983_));
  AOI210     o0934(.A0(ori_ori_n983_), .A1(ori_ori_n981_), .B0(x1), .Y(ori_ori_n984_));
  NO2        o0935(.A(ori_ori_n260_), .B(ori_ori_n246_), .Y(ori_ori_n985_));
  NA3        o0936(.A(ori_ori_n985_), .B(ori_ori_n594_), .C(x1), .Y(ori_ori_n986_));
  OAI210     o0937(.A0(x8), .A1(x0), .B0(x4), .Y(ori_ori_n987_));
  NO2        o0938(.A(x7), .B(ori_ori_n56_), .Y(ori_ori_n988_));
  NOi21      o0939(.An(ori_ori_n987_), .B(x7), .Y(ori_ori_n989_));
  NO2        o0940(.A(ori_ori_n588_), .B(ori_ori_n291_), .Y(ori_ori_n990_));
  INV        o0941(.A(ori_ori_n200_), .Y(ori_ori_n991_));
  OAI210     o0942(.A0(ori_ori_n990_), .A1(ori_ori_n989_), .B0(ori_ori_n991_), .Y(ori_ori_n992_));
  NO2        o0943(.A(ori_ori_n705_), .B(ori_ori_n374_), .Y(ori_ori_n993_));
  NA2        o0944(.A(x3), .B(ori_ori_n57_), .Y(ori_ori_n994_));
  NO2        o0945(.A(ori_ori_n945_), .B(ori_ori_n994_), .Y(ori_ori_n995_));
  AOI210     o0946(.A0(ori_ori_n993_), .A1(ori_ori_n160_), .B0(ori_ori_n995_), .Y(ori_ori_n996_));
  NA3        o0947(.A(ori_ori_n996_), .B(ori_ori_n992_), .C(ori_ori_n986_), .Y(ori_ori_n997_));
  OAI210     o0948(.A0(ori_ori_n997_), .A1(ori_ori_n984_), .B0(ori_ori_n595_), .Y(ori_ori_n998_));
  NA4        o0949(.A(ori_ori_n998_), .B(ori_ori_n979_), .C(ori_ori_n961_), .D(ori_ori_n947_), .Y(ori13));
  NO2        o0950(.A(ori_ori_n407_), .B(ori_ori_n312_), .Y(ori_ori_n1000_));
  NOi41      o0951(.An(ori_ori_n1000_), .B(ori_ori_n594_), .C(ori_ori_n262_), .D(ori_ori_n219_), .Y(ori_ori_n1001_));
  NO2        o0952(.A(ori_ori_n744_), .B(ori_ori_n164_), .Y(ori_ori_n1002_));
  NO2        o0953(.A(ori_ori_n144_), .B(ori_ori_n68_), .Y(ori_ori_n1003_));
  XN2        o0954(.A(x4), .B(x0), .Y(ori_ori_n1004_));
  NO3        o0955(.A(ori_ori_n1004_), .B(ori_ori_n101_), .C(ori_ori_n374_), .Y(ori_ori_n1005_));
  AN2        o0956(.A(ori_ori_n1005_), .B(ori_ori_n1003_), .Y(ori_ori_n1006_));
  OAI210     o0957(.A0(ori_ori_n1006_), .A1(ori_ori_n1001_), .B0(x3), .Y(ori_ori_n1007_));
  NO2        o0958(.A(ori_ori_n744_), .B(x6), .Y(ori_ori_n1008_));
  NO2        o0959(.A(ori_ori_n949_), .B(ori_ori_n352_), .Y(ori_ori_n1009_));
  NO3        o0960(.A(x8), .B(x5), .C(ori_ori_n100_), .Y(ori_ori_n1010_));
  NO2        o0961(.A(ori_ori_n532_), .B(ori_ori_n179_), .Y(ori_ori_n1011_));
  NA2        o0962(.A(ori_ori_n56_), .B(ori_ori_n100_), .Y(ori_ori_n1012_));
  NA2        o0963(.A(ori_ori_n1012_), .B(x1), .Y(ori_ori_n1013_));
  NO2        o0964(.A(ori_ori_n288_), .B(x6), .Y(ori_ori_n1014_));
  NO2        o0965(.A(ori_ori_n2177_), .B(ori_ori_n1014_), .Y(ori_ori_n1015_));
  NA2        o0966(.A(ori_ori_n1015_), .B(ori_ori_n532_), .Y(ori_ori_n1016_));
  AOI220     o0967(.A0(ori_ori_n1016_), .A1(ori_ori_n65_), .B0(ori_ori_n1009_), .B1(ori_ori_n1008_), .Y(ori_ori_n1017_));
  NA2        o0968(.A(ori_ori_n68_), .B(x3), .Y(ori_ori_n1018_));
  NA2        o0969(.A(ori_ori_n544_), .B(ori_ori_n55_), .Y(ori_ori_n1019_));
  NA2        o0970(.A(x6), .B(ori_ori_n50_), .Y(ori_ori_n1020_));
  NA2        o0971(.A(ori_ori_n1020_), .B(ori_ori_n471_), .Y(ori_ori_n1021_));
  OAI210     o0972(.A0(ori_ori_n544_), .A1(ori_ori_n644_), .B0(ori_ori_n971_), .Y(ori_ori_n1022_));
  NAi21      o0973(.An(ori_ori_n81_), .B(ori_ori_n341_), .Y(ori_ori_n1023_));
  NO2        o0974(.A(ori_ori_n1023_), .B(ori_ori_n68_), .Y(ori_ori_n1024_));
  AOI210     o0975(.A0(ori_ori_n148_), .A1(x4), .B0(ori_ori_n157_), .Y(ori_ori_n1025_));
  NO2        o0976(.A(ori_ori_n1025_), .B(x0), .Y(ori_ori_n1026_));
  NO2        o0977(.A(ori_ori_n154_), .B(ori_ori_n265_), .Y(ori_ori_n1027_));
  OAI210     o0978(.A0(ori_ori_n1027_), .A1(ori_ori_n1026_), .B0(ori_ori_n1024_), .Y(ori_ori_n1028_));
  NA3        o0979(.A(ori_ori_n976_), .B(ori_ori_n170_), .C(ori_ori_n68_), .Y(ori_ori_n1029_));
  NO2        o0980(.A(x4), .B(x0), .Y(ori_ori_n1030_));
  NO3        o0981(.A(ori_ori_n859_), .B(ori_ori_n226_), .C(ori_ori_n471_), .Y(ori_ori_n1031_));
  OAI210     o0982(.A0(ori_ori_n1031_), .A1(ori_ori_n180_), .B0(ori_ori_n1030_), .Y(ori_ori_n1032_));
  NA3        o0983(.A(ori_ori_n1032_), .B(ori_ori_n1029_), .C(ori_ori_n1028_), .Y(ori_ori_n1033_));
  NA2        o0984(.A(ori_ori_n227_), .B(ori_ori_n626_), .Y(ori_ori_n1034_));
  NO2        o0985(.A(ori_ori_n1034_), .B(ori_ori_n456_), .Y(ori_ori_n1035_));
  NA2        o0986(.A(ori_ori_n56_), .B(x0), .Y(ori_ori_n1036_));
  NO3        o0987(.A(ori_ori_n1036_), .B(ori_ori_n431_), .C(ori_ori_n78_), .Y(ori_ori_n1037_));
  OAI210     o0988(.A0(ori_ori_n1037_), .A1(ori_ori_n1035_), .B0(x2), .Y(ori_ori_n1038_));
  NO2        o0989(.A(ori_ori_n291_), .B(ori_ori_n341_), .Y(ori_ori_n1039_));
  NO2        o0990(.A(ori_ori_n604_), .B(x0), .Y(ori_ori_n1040_));
  OAI210     o0991(.A0(ori_ori_n1040_), .A1(ori_ori_n1039_), .B0(ori_ori_n297_), .Y(ori_ori_n1041_));
  NO2        o0992(.A(ori_ori_n677_), .B(x1), .Y(ori_ori_n1042_));
  AOI220     o0993(.A0(ori_ori_n1042_), .A1(ori_ori_n537_), .B0(ori_ori_n415_), .B1(ori_ori_n266_), .Y(ori_ori_n1043_));
  NA2        o0994(.A(ori_ori_n437_), .B(ori_ori_n50_), .Y(ori_ori_n1044_));
  AOI220     o0995(.A0(ori_ori_n1044_), .A1(ori_ori_n1002_), .B0(ori_ori_n845_), .B1(ori_ori_n92_), .Y(ori_ori_n1045_));
  NA4        o0996(.A(ori_ori_n1045_), .B(ori_ori_n1043_), .C(ori_ori_n1041_), .D(ori_ori_n1038_), .Y(ori_ori_n1046_));
  AOI220     o0997(.A0(ori_ori_n1046_), .A1(x8), .B0(ori_ori_n1033_), .B1(ori_ori_n64_), .Y(ori_ori_n1047_));
  NA4        o0998(.A(ori_ori_n1047_), .B(ori_ori_n1022_), .C(ori_ori_n1017_), .D(ori_ori_n1007_), .Y(ori14));
  NO2        o0999(.A(ori_ori_n333_), .B(ori_ori_n68_), .Y(ori_ori_n1049_));
  NO3        o1000(.A(x7), .B(x6), .C(x0), .Y(ori_ori_n1050_));
  NA2        o1001(.A(ori_ori_n1049_), .B(x8), .Y(ori_ori_n1051_));
  NO2        o1002(.A(ori_ori_n1051_), .B(ori_ori_n143_), .Y(ori_ori_n1052_));
  AOI220     o1003(.A0(ori_ori_n337_), .A1(ori_ori_n730_), .B0(ori_ori_n397_), .B1(ori_ori_n374_), .Y(ori_ori_n1053_));
  NA2        o1004(.A(ori_ori_n249_), .B(ori_ori_n840_), .Y(ori_ori_n1054_));
  OAI220     o1005(.A0(ori_ori_n1054_), .A1(ori_ori_n1053_), .B0(ori_ori_n409_), .B1(ori_ori_n689_), .Y(ori_ori_n1055_));
  OA210      o1006(.A0(ori_ori_n1055_), .A1(ori_ori_n1052_), .B0(x4), .Y(ori_ori_n1056_));
  NO2        o1007(.A(ori_ori_n129_), .B(ori_ori_n536_), .Y(ori_ori_n1057_));
  NA2        o1008(.A(x6), .B(x2), .Y(ori_ori_n1058_));
  NO2        o1009(.A(ori_ori_n553_), .B(ori_ori_n1058_), .Y(ori_ori_n1059_));
  OA210      o1010(.A0(ori_ori_n1057_), .A1(x4), .B0(ori_ori_n1059_), .Y(ori_ori_n1060_));
  NO4        o1011(.A(ori_ori_n532_), .B(ori_ori_n338_), .C(ori_ori_n270_), .D(ori_ori_n105_), .Y(ori_ori_n1061_));
  OAI210     o1012(.A0(ori_ori_n1061_), .A1(ori_ori_n1060_), .B0(ori_ori_n57_), .Y(ori_ori_n1062_));
  NA2        o1013(.A(x6), .B(ori_ori_n98_), .Y(ori_ori_n1063_));
  NO2        o1014(.A(ori_ori_n586_), .B(ori_ori_n1063_), .Y(ori_ori_n1064_));
  NA2        o1015(.A(ori_ori_n1064_), .B(ori_ori_n800_), .Y(ori_ori_n1065_));
  INV        o1016(.A(x1), .Y(ori_ori_n1066_));
  NO2        o1017(.A(ori_ori_n466_), .B(x5), .Y(ori_ori_n1067_));
  NA3        o1018(.A(ori_ori_n1067_), .B(ori_ori_n111_), .C(x0), .Y(ori_ori_n1068_));
  AN4        o1019(.A(ori_ori_n2167_), .B(ori_ori_n1068_), .C(ori_ori_n1066_), .D(ori_ori_n1065_), .Y(ori_ori_n1069_));
  AO210      o1020(.A0(ori_ori_n1049_), .A1(ori_ori_n872_), .B0(ori_ori_n53_), .Y(ori_ori_n1070_));
  INV        o1021(.A(ori_ori_n1070_), .Y(ori_ori_n1071_));
  AOI210     o1022(.A0(ori_ori_n1069_), .A1(ori_ori_n1062_), .B0(ori_ori_n1071_), .Y(ori_ori_n1072_));
  NO2        o1023(.A(x6), .B(ori_ori_n151_), .Y(ori_ori_n1073_));
  NO3        o1024(.A(ori_ori_n1073_), .B(ori_ori_n1072_), .C(ori_ori_n1056_), .Y(ori_ori_n1074_));
  NO2        o1025(.A(ori_ori_n288_), .B(x2), .Y(ori_ori_n1075_));
  XN2        o1026(.A(x4), .B(x1), .Y(ori_ori_n1076_));
  NO2        o1027(.A(ori_ori_n1076_), .B(ori_ori_n274_), .Y(ori_ori_n1077_));
  BUFFER     o1028(.A(ori_ori_n1077_), .Y(ori_ori_n1078_));
  NO2        o1029(.A(ori_ori_n301_), .B(ori_ori_n58_), .Y(ori_ori_n1079_));
  OAI210     o1030(.A0(ori_ori_n1079_), .A1(ori_ori_n1078_), .B0(ori_ori_n1075_), .Y(ori_ori_n1080_));
  OAI220     o1031(.A0(x4), .A1(ori_ori_n144_), .B0(ori_ori_n171_), .B1(ori_ori_n68_), .Y(ori_ori_n1081_));
  AOI220     o1032(.A0(ori_ori_n126_), .A1(ori_ori_n56_), .B0(ori_ori_n86_), .B1(x5), .Y(ori_ori_n1082_));
  NO2        o1033(.A(x6), .B(ori_ori_n1082_), .Y(ori_ori_n1083_));
  AOI210     o1034(.A0(x5), .A1(ori_ori_n1081_), .B0(ori_ori_n1083_), .Y(ori_ori_n1084_));
  AOI210     o1035(.A0(ori_ori_n1084_), .A1(ori_ori_n1080_), .B0(x7), .Y(ori_ori_n1085_));
  NO2        o1036(.A(ori_ori_n430_), .B(x6), .Y(ori_ori_n1086_));
  AOI210     o1037(.A0(ori_ori_n701_), .A1(ori_ori_n824_), .B0(ori_ori_n1086_), .Y(ori_ori_n1087_));
  OAI220     o1038(.A0(ori_ori_n1087_), .A1(ori_ori_n55_), .B0(ori_ori_n430_), .B1(ori_ori_n94_), .Y(ori_ori_n1088_));
  NA2        o1039(.A(ori_ori_n1088_), .B(ori_ori_n318_), .Y(ori_ori_n1089_));
  NA3        o1040(.A(ori_ori_n538_), .B(ori_ori_n900_), .C(ori_ori_n67_), .Y(ori_ori_n1090_));
  NO4        o1041(.A(ori_ori_n1090_), .B(ori_ori_n1036_), .C(ori_ori_n109_), .D(ori_ori_n55_), .Y(ori_ori_n1091_));
  NO3        o1042(.A(ori_ori_n898_), .B(ori_ori_n707_), .C(ori_ori_n420_), .Y(ori_ori_n1092_));
  NO3        o1043(.A(ori_ori_n646_), .B(ori_ori_n437_), .C(ori_ori_n54_), .Y(ori_ori_n1093_));
  NO4        o1044(.A(ori_ori_n1093_), .B(ori_ori_n1092_), .C(ori_ori_n1091_), .D(ori_ori_n888_), .Y(ori_ori_n1094_));
  AOI210     o1045(.A0(ori_ori_n1094_), .A1(ori_ori_n1089_), .B0(ori_ori_n276_), .Y(ori_ori_n1095_));
  NA2        o1046(.A(ori_ori_n776_), .B(ori_ori_n53_), .Y(ori_ori_n1096_));
  OAI210     o1047(.A0(ori_ori_n223_), .A1(ori_ori_n107_), .B0(x2), .Y(ori_ori_n1097_));
  NA2        o1048(.A(ori_ori_n56_), .B(x2), .Y(ori_ori_n1098_));
  NO2        o1049(.A(ori_ori_n1098_), .B(ori_ori_n178_), .Y(ori_ori_n1099_));
  NA4        o1050(.A(ori_ori_n1099_), .B(ori_ori_n329_), .C(ori_ori_n233_), .D(ori_ori_n64_), .Y(ori_ori_n1100_));
  INV        o1051(.A(ori_ori_n1100_), .Y(ori_ori_n1101_));
  NO3        o1052(.A(ori_ori_n1101_), .B(ori_ori_n1095_), .C(ori_ori_n1085_), .Y(ori_ori_n1102_));
  OAI210     o1053(.A0(ori_ori_n1074_), .A1(x3), .B0(ori_ori_n1102_), .Y(ori15));
  NAi41      o1054(.An(x2), .B(x7), .C(x6), .D(x0), .Y(ori_ori_n1104_));
  NO2        o1055(.A(ori_ori_n1104_), .B(ori_ori_n53_), .Y(ori_ori_n1105_));
  NA2        o1056(.A(ori_ori_n1105_), .B(ori_ori_n976_), .Y(ori_ori_n1106_));
  NA4        o1057(.A(x2), .B(ori_ori_n565_), .C(x0), .D(x6), .Y(ori_ori_n1107_));
  AOI210     o1058(.A0(ori_ori_n625_), .A1(ori_ori_n73_), .B0(x3), .Y(ori_ori_n1108_));
  NA3        o1059(.A(ori_ori_n1108_), .B(ori_ori_n1107_), .C(ori_ori_n1106_), .Y(ori_ori_n1109_));
  AOI210     o1060(.A0(ori_ori_n904_), .A1(ori_ori_n520_), .B0(ori_ori_n50_), .Y(ori_ori_n1110_));
  NO2        o1061(.A(ori_ori_n265_), .B(ori_ori_n100_), .Y(ori_ori_n1111_));
  NO2        o1062(.A(ori_ori_n217_), .B(x5), .Y(ori_ori_n1112_));
  NA2        o1063(.A(ori_ori_n1112_), .B(ori_ori_n1111_), .Y(ori_ori_n1113_));
  NA3        o1064(.A(ori_ori_n1113_), .B(ori_ori_n1110_), .C(ori_ori_n1068_), .Y(ori_ori_n1114_));
  INV        o1065(.A(ori_ori_n304_), .Y(ori_ori_n1115_));
  NO2        o1066(.A(ori_ori_n1013_), .B(ori_ori_n1115_), .Y(ori_ori_n1116_));
  NA4        o1067(.A(ori_ori_n1013_), .B(ori_ori_n609_), .C(ori_ori_n954_), .D(ori_ori_n341_), .Y(ori_ori_n1117_));
  NA2        o1068(.A(ori_ori_n520_), .B(ori_ori_n410_), .Y(ori_ori_n1118_));
  NO2        o1069(.A(ori_ori_n646_), .B(ori_ori_n53_), .Y(ori_ori_n1119_));
  NA2        o1070(.A(ori_ori_n2180_), .B(ori_ori_n1119_), .Y(ori_ori_n1120_));
  NA3        o1071(.A(ori_ori_n1120_), .B(ori_ori_n1118_), .C(ori_ori_n1117_), .Y(ori_ori_n1121_));
  OAI210     o1072(.A0(ori_ori_n1121_), .A1(ori_ori_n1116_), .B0(ori_ori_n74_), .Y(ori_ori_n1122_));
  NA2        o1073(.A(ori_ori_n331_), .B(ori_ori_n611_), .Y(ori_ori_n1123_));
  NA2        o1074(.A(x1), .B(ori_ori_n56_), .Y(ori_ori_n1124_));
  NA2        o1075(.A(ori_ori_n1124_), .B(ori_ori_n304_), .Y(ori_ori_n1125_));
  AOI210     o1076(.A0(ori_ori_n1125_), .A1(ori_ori_n1123_), .B0(ori_ori_n437_), .Y(ori_ori_n1126_));
  NO3        o1077(.A(ori_ori_n688_), .B(ori_ori_n549_), .C(ori_ori_n179_), .Y(ori_ori_n1127_));
  OAI210     o1078(.A0(ori_ori_n1127_), .A1(ori_ori_n1126_), .B0(ori_ori_n430_), .Y(ori_ori_n1128_));
  NO2        o1079(.A(ori_ori_n750_), .B(ori_ori_n50_), .Y(ori_ori_n1129_));
  AN2        o1080(.A(ori_ori_n1129_), .B(ori_ori_n366_), .Y(ori_ori_n1130_));
  NO2        o1081(.A(ori_ori_n846_), .B(ori_ori_n599_), .Y(ori_ori_n1131_));
  OAI210     o1082(.A0(ori_ori_n1131_), .A1(ori_ori_n1130_), .B0(ori_ori_n879_), .Y(ori_ori_n1132_));
  NO2        o1083(.A(ori_ori_n1058_), .B(x0), .Y(ori_ori_n1133_));
  AOI210     o1084(.A0(ori_ori_n1133_), .A1(ori_ori_n533_), .B0(x8), .Y(ori_ori_n1134_));
  NO2        o1085(.A(x1), .B(ori_ori_n78_), .Y(ori_ori_n1135_));
  NO2        o1086(.A(ori_ori_n807_), .B(ori_ori_n68_), .Y(ori_ori_n1136_));
  NA2        o1087(.A(ori_ori_n1136_), .B(ori_ori_n1135_), .Y(ori_ori_n1137_));
  NO2        o1088(.A(ori_ori_n844_), .B(x6), .Y(ori_ori_n1138_));
  NA3        o1089(.A(ori_ori_n1138_), .B(ori_ori_n145_), .C(ori_ori_n368_), .Y(ori_ori_n1139_));
  AN3        o1090(.A(ori_ori_n1139_), .B(ori_ori_n1137_), .C(ori_ori_n1134_), .Y(ori_ori_n1140_));
  NA4        o1091(.A(ori_ori_n1140_), .B(ori_ori_n1132_), .C(ori_ori_n1128_), .D(ori_ori_n1122_), .Y(ori_ori_n1141_));
  NA2        o1092(.A(ori_ori_n149_), .B(ori_ori_n631_), .Y(ori_ori_n1142_));
  OAI210     o1093(.A0(ori_ori_n65_), .A1(ori_ori_n53_), .B0(ori_ori_n132_), .Y(ori_ori_n1143_));
  NA2        o1094(.A(ori_ori_n82_), .B(ori_ori_n1143_), .Y(ori_ori_n1144_));
  AOI210     o1095(.A0(ori_ori_n1144_), .A1(ori_ori_n1142_), .B0(ori_ori_n288_), .Y(ori_ori_n1145_));
  NA3        o1096(.A(ori_ori_n68_), .B(x5), .C(x2), .Y(ori_ori_n1146_));
  NA4        o1097(.A(x7), .B(x3), .C(ori_ori_n53_), .D(x0), .Y(ori_ori_n1147_));
  NO2        o1098(.A(ori_ori_n1147_), .B(x6), .Y(ori_ori_n1148_));
  INV        o1099(.A(ori_ori_n1148_), .Y(ori_ori_n1149_));
  NAi21      o1100(.An(ori_ori_n105_), .B(ori_ori_n641_), .Y(ori_ori_n1150_));
  NA4        o1101(.A(ori_ori_n1150_), .B(ori_ori_n286_), .C(ori_ori_n260_), .D(ori_ori_n552_), .Y(ori_ori_n1151_));
  OAI220     o1102(.A0(ori_ori_n291_), .A1(x7), .B0(ori_ori_n120_), .B1(ori_ori_n68_), .Y(ori_ori_n1152_));
  NA3        o1103(.A(ori_ori_n1152_), .B(ori_ori_n677_), .C(ori_ori_n929_), .Y(ori_ori_n1153_));
  NA2        o1104(.A(ori_ori_n79_), .B(ori_ori_n50_), .Y(ori_ori_n1154_));
  AO210      o1105(.A0(ori_ori_n1154_), .A1(ori_ori_n283_), .B0(ori_ori_n143_), .Y(ori_ori_n1155_));
  NA4        o1106(.A(ori_ori_n1155_), .B(ori_ori_n1153_), .C(ori_ori_n1151_), .D(ori_ori_n1149_), .Y(ori_ori_n1156_));
  OAI210     o1107(.A0(ori_ori_n1156_), .A1(ori_ori_n1145_), .B0(ori_ori_n56_), .Y(ori_ori_n1157_));
  AOI210     o1108(.A0(ori_ori_n606_), .A1(x4), .B0(ori_ori_n824_), .Y(ori_ori_n1158_));
  NO2        o1109(.A(ori_ori_n1158_), .B(ori_ori_n271_), .Y(ori_ori_n1159_));
  NA2        o1110(.A(ori_ori_n715_), .B(ori_ori_n363_), .Y(ori_ori_n1160_));
  NA2        o1111(.A(ori_ori_n1135_), .B(ori_ori_n261_), .Y(ori_ori_n1161_));
  OAI210     o1112(.A0(ori_ori_n1160_), .A1(x1), .B0(ori_ori_n1161_), .Y(ori_ori_n1162_));
  OAI210     o1113(.A0(ori_ori_n1162_), .A1(ori_ori_n1159_), .B0(x6), .Y(ori_ori_n1163_));
  NA2        o1114(.A(ori_ori_n734_), .B(x0), .Y(ori_ori_n1164_));
  NA2        o1115(.A(ori_ori_n656_), .B(ori_ori_n261_), .Y(ori_ori_n1165_));
  NA3        o1116(.A(ori_ori_n544_), .B(ori_ori_n263_), .C(ori_ori_n221_), .Y(ori_ori_n1166_));
  NA3        o1117(.A(ori_ori_n1166_), .B(ori_ori_n1165_), .C(ori_ori_n1164_), .Y(ori_ori_n1167_));
  NA2        o1118(.A(ori_ori_n1167_), .B(ori_ori_n377_), .Y(ori_ori_n1168_));
  NA4        o1119(.A(x8), .B(ori_ori_n1168_), .C(ori_ori_n1163_), .D(ori_ori_n1157_), .Y(ori_ori_n1169_));
  AO220      o1120(.A0(ori_ori_n1169_), .A1(ori_ori_n1141_), .B0(ori_ori_n1114_), .B1(ori_ori_n1109_), .Y(ori16));
  NO2        o1121(.A(x4), .B(ori_ori_n57_), .Y(ori_ori_n1171_));
  NA3        o1122(.A(ori_ori_n211_), .B(ori_ori_n382_), .C(ori_ori_n824_), .Y(ori_ori_n1172_));
  INV        o1123(.A(ori_ori_n188_), .Y(ori_ori_n1173_));
  NO2        o1124(.A(ori_ori_n1172_), .B(ori_ori_n1173_), .Y(ori_ori_n1174_));
  NO3        o1125(.A(x8), .B(x6), .C(ori_ori_n50_), .Y(ori_ori_n1175_));
  NO2        o1126(.A(ori_ori_n629_), .B(ori_ori_n166_), .Y(ori_ori_n1176_));
  OAI210     o1127(.A0(ori_ori_n1175_), .A1(ori_ori_n219_), .B0(ori_ori_n1176_), .Y(ori_ori_n1177_));
  NA3        o1128(.A(ori_ori_n510_), .B(ori_ori_n469_), .C(ori_ori_n414_), .Y(ori_ori_n1178_));
  NA2        o1129(.A(ori_ori_n1178_), .B(ori_ori_n1177_), .Y(ori_ori_n1179_));
  OAI210     o1130(.A0(ori_ori_n1179_), .A1(ori_ori_n1174_), .B0(ori_ori_n1171_), .Y(ori_ori_n1180_));
  OAI210     o1131(.A0(ori_ori_n1075_), .A1(ori_ori_n800_), .B0(ori_ori_n374_), .Y(ori_ori_n1181_));
  NO2        o1132(.A(ori_ori_n1181_), .B(ori_ori_n566_), .Y(ori_ori_n1182_));
  NA2        o1133(.A(ori_ori_n908_), .B(ori_ori_n179_), .Y(ori_ori_n1183_));
  NA2        o1134(.A(ori_ori_n55_), .B(ori_ori_n98_), .Y(ori_ori_n1184_));
  NA2        o1135(.A(ori_ori_n1184_), .B(ori_ori_n601_), .Y(ori_ori_n1185_));
  NA2        o1136(.A(ori_ori_n339_), .B(ori_ori_n912_), .Y(ori_ori_n1186_));
  OA220      o1137(.A0(ori_ori_n1186_), .A1(ori_ori_n1185_), .B0(ori_ori_n1183_), .B1(ori_ori_n560_), .Y(ori_ori_n1187_));
  OAI210     o1138(.A0(ori_ori_n1187_), .A1(ori_ori_n577_), .B0(ori_ori_n435_), .Y(ori_ori_n1188_));
  INV        o1139(.A(ori_ori_n879_), .Y(ori_ori_n1189_));
  NO2        o1140(.A(ori_ori_n1189_), .B(ori_ori_n60_), .Y(ori_ori_n1190_));
  AOI220     o1141(.A0(ori_ori_n1190_), .A1(ori_ori_n241_), .B0(ori_ori_n1064_), .B1(ori_ori_n116_), .Y(ori_ori_n1191_));
  AOI210     o1142(.A0(ori_ori_n565_), .A1(ori_ori_n325_), .B0(ori_ori_n552_), .Y(ori_ori_n1192_));
  NA3        o1143(.A(ori_ori_n408_), .B(ori_ori_n517_), .C(ori_ori_n173_), .Y(ori_ori_n1193_));
  OAI220     o1144(.A0(ori_ori_n1193_), .A1(ori_ori_n1192_), .B0(ori_ori_n1191_), .B1(ori_ori_n280_), .Y(ori_ori_n1194_));
  NO3        o1145(.A(ori_ori_n1194_), .B(ori_ori_n1188_), .C(ori_ori_n1182_), .Y(ori_ori_n1195_));
  NO3        o1146(.A(x6), .B(x4), .C(x3), .Y(ori_ori_n1196_));
  NA2        o1147(.A(ori_ori_n1196_), .B(ori_ori_n466_), .Y(ori_ori_n1197_));
  NA3        o1148(.A(ori_ori_n613_), .B(ori_ori_n166_), .C(x6), .Y(ori_ori_n1198_));
  AOI210     o1149(.A0(ori_ori_n1198_), .A1(ori_ori_n1197_), .B0(ori_ori_n54_), .Y(ori_ori_n1199_));
  NO2        o1150(.A(ori_ori_n617_), .B(x3), .Y(ori_ori_n1200_));
  NO2        o1151(.A(ori_ori_n135_), .B(ori_ori_n900_), .Y(ori_ori_n1201_));
  OA210      o1152(.A0(ori_ori_n1200_), .A1(ori_ori_n377_), .B0(ori_ori_n1201_), .Y(ori_ori_n1202_));
  NO3        o1153(.A(ori_ori_n437_), .B(ori_ori_n200_), .C(ori_ori_n72_), .Y(ori_ori_n1203_));
  NO2        o1154(.A(ori_ori_n656_), .B(ori_ori_n449_), .Y(ori_ori_n1204_));
  NO3        o1155(.A(ori_ori_n1204_), .B(ori_ori_n235_), .C(ori_ori_n142_), .Y(ori_ori_n1205_));
  NO4        o1156(.A(ori_ori_n1205_), .B(ori_ori_n1203_), .C(ori_ori_n1202_), .D(ori_ori_n1199_), .Y(ori_ori_n1206_));
  NA2        o1157(.A(ori_ori_n364_), .B(ori_ori_n824_), .Y(ori_ori_n1207_));
  NA4        o1158(.A(ori_ori_n420_), .B(ori_ori_n333_), .C(ori_ori_n202_), .D(x6), .Y(ori_ori_n1208_));
  OAI210     o1159(.A0(ori_ori_n617_), .A1(ori_ori_n1207_), .B0(ori_ori_n1208_), .Y(ori_ori_n1209_));
  NA2        o1160(.A(ori_ori_n626_), .B(x7), .Y(ori_ori_n1210_));
  NO2        o1161(.A(ori_ori_n1210_), .B(ori_ori_n347_), .Y(ori_ori_n1211_));
  NA2        o1162(.A(ori_ori_n247_), .B(x2), .Y(ori_ori_n1212_));
  AOI210     o1163(.A0(ori_ori_n510_), .A1(ori_ori_n50_), .B0(ori_ori_n520_), .Y(ori_ori_n1213_));
  OAI210     o1164(.A0(ori_ori_n801_), .A1(ori_ori_n816_), .B0(ori_ori_n343_), .Y(ori_ori_n1214_));
  NO2        o1165(.A(ori_ori_n1214_), .B(ori_ori_n1213_), .Y(ori_ori_n1215_));
  NO3        o1166(.A(ori_ori_n1215_), .B(ori_ori_n1211_), .C(ori_ori_n1209_), .Y(ori_ori_n1216_));
  OA220      o1167(.A0(ori_ori_n1216_), .A1(ori_ori_n393_), .B0(ori_ori_n1206_), .B1(ori_ori_n186_), .Y(ori_ori_n1217_));
  NO2        o1168(.A(ori_ori_n796_), .B(ori_ori_n55_), .Y(ori_ori_n1218_));
  NA2        o1169(.A(ori_ori_n371_), .B(ori_ori_n689_), .Y(ori_ori_n1219_));
  NO2        o1170(.A(ori_ori_n1219_), .B(ori_ori_n1218_), .Y(ori_ori_n1220_));
  NA2        o1171(.A(ori_ori_n1220_), .B(x6), .Y(ori_ori_n1221_));
  NO2        o1172(.A(ori_ori_n924_), .B(ori_ori_n897_), .Y(ori_ori_n1222_));
  NA2        o1173(.A(ori_ori_n171_), .B(x7), .Y(ori_ori_n1223_));
  OAI220     o1174(.A0(ori_ori_n1223_), .A1(ori_ori_n1222_), .B0(x6), .B1(ori_ori_n83_), .Y(ori_ori_n1224_));
  NA2        o1175(.A(ori_ori_n1224_), .B(ori_ori_n801_), .Y(ori_ori_n1225_));
  NA2        o1176(.A(ori_ori_n752_), .B(ori_ori_n68_), .Y(ori_ori_n1226_));
  INV        o1177(.A(ori_ori_n869_), .Y(ori_ori_n1227_));
  INV        o1178(.A(ori_ori_n560_), .Y(ori_ori_n1228_));
  NA3        o1179(.A(ori_ori_n208_), .B(ori_ori_n73_), .C(ori_ori_n68_), .Y(ori_ori_n1229_));
  OAI210     o1180(.A0(ori_ori_n2176_), .A1(ori_ori_n211_), .B0(ori_ori_n1229_), .Y(ori_ori_n1230_));
  AOI210     o1181(.A0(ori_ori_n1228_), .A1(ori_ori_n1227_), .B0(ori_ori_n1230_), .Y(ori_ori_n1231_));
  NA3        o1182(.A(ori_ori_n1231_), .B(ori_ori_n1225_), .C(ori_ori_n1221_), .Y(ori_ori_n1232_));
  NO2        o1183(.A(ori_ori_n567_), .B(x6), .Y(ori_ori_n1233_));
  OAI210     o1184(.A0(ori_ori_n343_), .A1(ori_ori_n81_), .B0(ori_ori_n341_), .Y(ori_ori_n1234_));
  OA210      o1185(.A0(ori_ori_n1234_), .A1(ori_ori_n1233_), .B0(x8), .Y(ori_ori_n1235_));
  NO3        o1186(.A(ori_ori_n395_), .B(ori_ori_n345_), .C(x7), .Y(ori_ori_n1236_));
  NO3        o1187(.A(ori_ori_n146_), .B(ori_ori_n72_), .C(x2), .Y(ori_ori_n1237_));
  NO3        o1188(.A(ori_ori_n1237_), .B(ori_ori_n1236_), .C(ori_ori_n1235_), .Y(ori_ori_n1238_));
  NA2        o1189(.A(ori_ori_n917_), .B(x5), .Y(ori_ori_n1239_));
  NO2        o1190(.A(ori_ori_n1239_), .B(ori_ori_n56_), .Y(ori_ori_n1240_));
  NA2        o1191(.A(x6), .B(ori_ori_n664_), .Y(ori_ori_n1241_));
  NO2        o1192(.A(ori_ori_n1241_), .B(ori_ori_n1098_), .Y(ori_ori_n1242_));
  NO3        o1193(.A(ori_ori_n466_), .B(ori_ori_n156_), .C(ori_ori_n897_), .Y(ori_ori_n1243_));
  NO3        o1194(.A(ori_ori_n1243_), .B(ori_ori_n1242_), .C(ori_ori_n1240_), .Y(ori_ori_n1244_));
  OAI210     o1195(.A0(ori_ori_n1238_), .A1(x5), .B0(ori_ori_n1244_), .Y(ori_ori_n1245_));
  AOI220     o1196(.A0(ori_ori_n1245_), .A1(ori_ori_n90_), .B0(ori_ori_n1232_), .B1(ori_ori_n302_), .Y(ori_ori_n1246_));
  NA4        o1197(.A(ori_ori_n1246_), .B(ori_ori_n1217_), .C(ori_ori_n1195_), .D(ori_ori_n1180_), .Y(ori17));
  NO4        o1198(.A(ori_ori_n530_), .B(ori_ori_n610_), .C(ori_ori_n93_), .D(ori_ori_n92_), .Y(ori_ori_n1248_));
  AOI220     o1199(.A0(ori_ori_n2175_), .A1(ori_ori_n616_), .B0(ori_ori_n1248_), .B1(ori_ori_n443_), .Y(ori_ori_n1249_));
  NA2        o1200(.A(ori_ori_n149_), .B(ori_ori_n75_), .Y(ori_ori_n1250_));
  NOi21      o1201(.An(ori_ori_n341_), .B(ori_ori_n81_), .Y(ori_ori_n1251_));
  OAI210     o1202(.A0(ori_ori_n613_), .A1(x8), .B0(ori_ori_n1098_), .Y(ori_ori_n1252_));
  NA3        o1203(.A(ori_ori_n1252_), .B(ori_ori_n1049_), .C(ori_ori_n359_), .Y(ori_ori_n1253_));
  NA2        o1204(.A(ori_ori_n241_), .B(ori_ori_n516_), .Y(ori_ori_n1254_));
  NA3        o1205(.A(ori_ori_n648_), .B(ori_ori_n1254_), .C(ori_ori_n1253_), .Y(ori_ori_n1255_));
  NA3        o1206(.A(ori_ori_n148_), .B(ori_ori_n558_), .C(ori_ori_n897_), .Y(ori_ori_n1256_));
  AOI210     o1207(.A0(ori_ori_n914_), .A1(ori_ori_n277_), .B0(ori_ori_n57_), .Y(ori_ori_n1257_));
  NA2        o1208(.A(ori_ori_n1257_), .B(ori_ori_n1256_), .Y(ori_ori_n1258_));
  AOI210     o1209(.A0(ori_ori_n1255_), .A1(x1), .B0(ori_ori_n1258_), .Y(ori_ori_n1259_));
  OAI210     o1210(.A0(ori_ori_n68_), .A1(ori_ori_n903_), .B0(ori_ori_n536_), .Y(ori_ori_n1260_));
  NO3        o1211(.A(ori_ori_n560_), .B(ori_ori_n486_), .C(ori_ori_n459_), .Y(ori_ori_n1261_));
  OAI210     o1212(.A0(ori_ori_n1261_), .A1(ori_ori_n783_), .B0(ori_ori_n1200_), .Y(ori_ori_n1262_));
  AOI210     o1213(.A0(ori_ori_n1262_), .A1(ori_ori_n1260_), .B0(x8), .Y(ori_ori_n1263_));
  NA3        o1214(.A(ori_ori_n560_), .B(ori_ori_n244_), .C(ori_ori_n111_), .Y(ori_ori_n1264_));
  NO2        o1215(.A(ori_ori_n132_), .B(ori_ori_n130_), .Y(ori_ori_n1265_));
  NO2        o1216(.A(ori_ori_n1265_), .B(x0), .Y(ori_ori_n1266_));
  NA2        o1217(.A(ori_ori_n1264_), .B(ori_ori_n1266_), .Y(ori_ori_n1267_));
  NO2        o1218(.A(ori_ori_n1267_), .B(ori_ori_n1263_), .Y(ori_ori_n1268_));
  OAI220     o1219(.A0(ori_ori_n1268_), .A1(ori_ori_n1259_), .B0(ori_ori_n1250_), .B1(ori_ori_n1249_), .Y(ori18));
  AOI210     o1220(.A0(x8), .A1(x0), .B0(x5), .Y(ori_ori_n1270_));
  NOi31      o1221(.An(ori_ori_n277_), .B(ori_ori_n1270_), .C(ori_ori_n896_), .Y(ori_ori_n1271_));
  NO2        o1222(.A(ori_ori_n545_), .B(ori_ori_n665_), .Y(ori_ori_n1272_));
  NO2        o1223(.A(ori_ori_n1272_), .B(ori_ori_n1271_), .Y(ori_ori_n1273_));
  NA3        o1224(.A(ori_ori_n457_), .B(ori_ori_n196_), .C(x0), .Y(ori_ori_n1274_));
  NAi21      o1225(.An(ori_ori_n346_), .B(ori_ori_n1274_), .Y(ori_ori_n1275_));
  NO2        o1226(.A(ori_ori_n769_), .B(x5), .Y(ori_ori_n1276_));
  AOI210     o1227(.A0(ori_ori_n967_), .A1(x5), .B0(ori_ori_n1276_), .Y(ori_ori_n1277_));
  OR2        o1228(.A(ori_ori_n359_), .B(x5), .Y(ori_ori_n1278_));
  OAI220     o1229(.A0(ori_ori_n1278_), .A1(ori_ori_n265_), .B0(ori_ori_n1277_), .B1(ori_ori_n194_), .Y(ori_ori_n1279_));
  AOI210     o1230(.A0(ori_ori_n1275_), .A1(ori_ori_n263_), .B0(ori_ori_n1279_), .Y(ori_ori_n1280_));
  AOI210     o1231(.A0(ori_ori_n1280_), .A1(ori_ori_n1273_), .B0(x6), .Y(ori_ori_n1281_));
  NA3        o1232(.A(ori_ori_n458_), .B(ori_ori_n374_), .C(x2), .Y(ori_ori_n1282_));
  NO2        o1233(.A(ori_ori_n1282_), .B(ori_ori_n677_), .Y(ori_ori_n1283_));
  AOI210     o1234(.A0(ori_ori_n378_), .A1(ori_ori_n126_), .B0(ori_ori_n676_), .Y(ori_ori_n1284_));
  NA2        o1235(.A(ori_ori_n241_), .B(x6), .Y(ori_ori_n1285_));
  OAI210     o1236(.A0(ori_ori_n160_), .A1(ori_ori_n100_), .B0(ori_ori_n973_), .Y(ori_ori_n1286_));
  OAI220     o1237(.A0(ori_ori_n1286_), .A1(ori_ori_n1285_), .B0(ori_ori_n1284_), .B1(ori_ori_n641_), .Y(ori_ori_n1287_));
  OAI210     o1238(.A0(ori_ori_n1287_), .A1(ori_ori_n1283_), .B0(ori_ori_n53_), .Y(ori_ori_n1288_));
  NO2        o1239(.A(ori_ori_n238_), .B(x3), .Y(ori_ori_n1289_));
  NO3        o1240(.A(ori_ori_n386_), .B(ori_ori_n530_), .C(ori_ori_n720_), .Y(ori_ori_n1290_));
  NA2        o1241(.A(ori_ori_n1290_), .B(ori_ori_n1289_), .Y(ori_ori_n1291_));
  INV        o1242(.A(x4), .Y(ori_ori_n1292_));
  OAI210     o1243(.A0(ori_ori_n486_), .A1(ori_ori_n530_), .B0(ori_ori_n57_), .Y(ori_ori_n1293_));
  INV        o1244(.A(ori_ori_n1293_), .Y(ori_ori_n1294_));
  AO220      o1245(.A0(ori_ori_n1067_), .A1(ori_ori_n629_), .B0(ori_ori_n487_), .B1(ori_ori_n318_), .Y(ori_ori_n1295_));
  AOI220     o1246(.A0(ori_ori_n1295_), .A1(x1), .B0(ori_ori_n1294_), .B1(ori_ori_n147_), .Y(ori_ori_n1296_));
  NA4        o1247(.A(ori_ori_n1296_), .B(ori_ori_n1292_), .C(ori_ori_n1291_), .D(ori_ori_n1288_), .Y(ori_ori_n1297_));
  NO3        o1248(.A(ori_ori_n905_), .B(x8), .C(ori_ori_n120_), .Y(ori_ori_n1298_));
  OAI210     o1249(.A0(ori_ori_n1298_), .A1(ori_ori_n578_), .B0(ori_ori_n98_), .Y(ori_ori_n1299_));
  AOI210     o1250(.A0(ori_ori_n1299_), .A1(ori_ori_n492_), .B0(ori_ori_n677_), .Y(ori_ori_n1300_));
  NA3        o1251(.A(ori_ori_n1019_), .B(ori_ori_n171_), .C(ori_ori_n129_), .Y(ori_ori_n1301_));
  NA3        o1252(.A(ori_ori_n908_), .B(ori_ori_n666_), .C(ori_ori_n306_), .Y(ori_ori_n1302_));
  NA2        o1253(.A(ori_ori_n154_), .B(ori_ori_n664_), .Y(ori_ori_n1303_));
  OAI210     o1254(.A0(ori_ori_n1303_), .A1(x2), .B0(ori_ori_n1302_), .Y(ori_ori_n1304_));
  AOI210     o1255(.A0(ori_ori_n1301_), .A1(ori_ori_n159_), .B0(ori_ori_n1304_), .Y(ori_ori_n1305_));
  OAI210     o1256(.A0(ori_ori_n1305_), .A1(ori_ori_n475_), .B0(x4), .Y(ori_ori_n1306_));
  OAI220     o1257(.A0(ori_ori_n1306_), .A1(ori_ori_n1300_), .B0(ori_ori_n1297_), .B1(ori_ori_n1281_), .Y(ori_ori_n1307_));
  NO2        o1258(.A(ori_ori_n134_), .B(ori_ori_n112_), .Y(ori_ori_n1308_));
  NO2        o1259(.A(ori_ori_n171_), .B(ori_ori_n689_), .Y(ori_ori_n1309_));
  AOI210     o1260(.A0(ori_ori_n531_), .A1(ori_ori_n449_), .B0(ori_ori_n1309_), .Y(ori_ori_n1310_));
  NO2        o1261(.A(ori_ori_n1310_), .B(x6), .Y(ori_ori_n1311_));
  NO2        o1262(.A(ori_ori_n345_), .B(ori_ori_n230_), .Y(ori_ori_n1312_));
  NO2        o1263(.A(ori_ori_n825_), .B(ori_ori_n516_), .Y(ori_ori_n1313_));
  AO220      o1264(.A0(ori_ori_n1313_), .A1(ori_ori_n55_), .B0(ori_ori_n1312_), .B1(ori_ori_n114_), .Y(ori_ori_n1314_));
  NO3        o1265(.A(ori_ori_n1314_), .B(ori_ori_n1311_), .C(ori_ori_n1308_), .Y(ori_ori_n1315_));
  NA2        o1266(.A(ori_ori_n905_), .B(x3), .Y(ori_ori_n1316_));
  INV        o1267(.A(ori_ori_n1138_), .Y(ori_ori_n1317_));
  OAI220     o1268(.A0(ori_ori_n1317_), .A1(ori_ori_n1316_), .B0(ori_ori_n1315_), .B1(x3), .Y(ori_ori_n1318_));
  NO3        o1269(.A(ori_ori_n865_), .B(ori_ori_n605_), .C(x3), .Y(ori_ori_n1319_));
  AO210      o1270(.A0(ori_ori_n887_), .A1(ori_ori_n270_), .B0(ori_ori_n1319_), .Y(ori_ori_n1320_));
  AOI220     o1271(.A0(ori_ori_n1320_), .A1(x8), .B0(ori_ori_n1138_), .B1(ori_ori_n387_), .Y(ori_ori_n1321_));
  NA2        o1272(.A(ori_ori_n644_), .B(ori_ori_n287_), .Y(ori_ori_n1322_));
  NO4        o1273(.A(ori_ori_n331_), .B(ori_ori_n184_), .C(ori_ori_n301_), .D(x2), .Y(ori_ori_n1323_));
  NA2        o1274(.A(ori_ori_n1184_), .B(ori_ori_n100_), .Y(ori_ori_n1324_));
  NO3        o1275(.A(ori_ori_n1020_), .B(ori_ori_n859_), .C(ori_ori_n973_), .Y(ori_ori_n1325_));
  AOI210     o1276(.A0(ori_ori_n1325_), .A1(ori_ori_n1324_), .B0(ori_ori_n1323_), .Y(ori_ori_n1326_));
  OA220      o1277(.A0(ori_ori_n1326_), .A1(ori_ori_n825_), .B0(ori_ori_n1322_), .B1(ori_ori_n501_), .Y(ori_ori_n1327_));
  OAI210     o1278(.A0(ori_ori_n1321_), .A1(ori_ori_n367_), .B0(ori_ori_n1327_), .Y(ori_ori_n1328_));
  AOI210     o1279(.A0(ori_ori_n1318_), .A1(ori_ori_n126_), .B0(ori_ori_n1328_), .Y(ori_ori_n1329_));
  NA2        o1280(.A(ori_ori_n1329_), .B(ori_ori_n1307_), .Y(ori19));
  NO2        o1281(.A(ori_ori_n1226_), .B(ori_ori_n234_), .Y(ori_ori_n1331_));
  INV        o1282(.A(x3), .Y(ori_ori_n1332_));
  NO2        o1283(.A(ori_ori_n1104_), .B(ori_ori_n154_), .Y(ori_ori_n1333_));
  INV        o1284(.A(ori_ori_n1333_), .Y(ori_ori_n1334_));
  NO2        o1285(.A(ori_ori_n1334_), .B(ori_ori_n56_), .Y(ori_ori_n1335_));
  NO2        o1286(.A(ori_ori_n742_), .B(ori_ori_n1030_), .Y(ori_ori_n1336_));
  OAI210     o1287(.A0(ori_ori_n1335_), .A1(ori_ori_n1331_), .B0(ori_ori_n1336_), .Y(ori_ori_n1337_));
  NOi21      o1288(.An(ori_ori_n539_), .B(ori_ori_n577_), .Y(ori_ori_n1338_));
  AOI210     o1289(.A0(ori_ori_n316_), .A1(x6), .B0(ori_ori_n111_), .Y(ori_ori_n1339_));
  NO3        o1290(.A(ori_ori_n1339_), .B(ori_ori_n653_), .C(ori_ori_n116_), .Y(ori_ori_n1340_));
  NA2        o1291(.A(ori_ori_n1018_), .B(ori_ori_n112_), .Y(ori_ori_n1341_));
  NO4        o1292(.A(ori_ori_n1341_), .B(ori_ori_n865_), .C(ori_ori_n769_), .D(ori_ori_n74_), .Y(ori_ori_n1342_));
  NO3        o1293(.A(ori_ori_n1342_), .B(ori_ori_n1340_), .C(ori_ori_n884_), .Y(ori_ori_n1343_));
  NO2        o1294(.A(ori_ori_n475_), .B(ori_ori_n548_), .Y(ori_ori_n1344_));
  NA2        o1295(.A(ori_ori_n1344_), .B(ori_ori_n666_), .Y(ori_ori_n1345_));
  NA2        o1296(.A(ori_ori_n1343_), .B(ori_ori_n1345_), .Y(ori_ori_n1346_));
  AOI210     o1297(.A0(ori_ori_n1346_), .A1(ori_ori_n664_), .B0(ori_ori_n1338_), .Y(ori_ori_n1347_));
  NA2        o1298(.A(ori_ori_n708_), .B(ori_ori_n631_), .Y(ori_ori_n1348_));
  NO2        o1299(.A(ori_ori_n1348_), .B(x4), .Y(ori_ori_n1349_));
  NA3        o1300(.A(ori_ori_n629_), .B(ori_ori_n233_), .C(x7), .Y(ori_ori_n1350_));
  NA2        o1301(.A(ori_ori_n610_), .B(ori_ori_n988_), .Y(ori_ori_n1351_));
  AOI210     o1302(.A0(ori_ori_n1351_), .A1(ori_ori_n1350_), .B0(ori_ori_n441_), .Y(ori_ori_n1352_));
  OAI210     o1303(.A0(ori_ori_n1352_), .A1(ori_ori_n1349_), .B0(ori_ori_n699_), .Y(ori_ori_n1353_));
  NO2        o1304(.A(ori_ori_n641_), .B(ori_ori_n291_), .Y(ori_ori_n1354_));
  NA2        o1305(.A(ori_ori_n1354_), .B(ori_ori_n415_), .Y(ori_ori_n1355_));
  AO210      o1306(.A0(ori_ori_n1355_), .A1(ori_ori_n1353_), .B0(x1), .Y(ori_ori_n1356_));
  NA2        o1307(.A(ori_ori_n560_), .B(ori_ori_n897_), .Y(ori_ori_n1357_));
  NA2        o1308(.A(ori_ori_n135_), .B(ori_ori_n101_), .Y(ori_ori_n1358_));
  NOi21      o1309(.An(x1), .B(x6), .Y(ori_ori_n1359_));
  NA2        o1310(.A(ori_ori_n1359_), .B(ori_ori_n81_), .Y(ori_ori_n1360_));
  NA3        o1311(.A(ori_ori_n1360_), .B(ori_ori_n1358_), .C(ori_ori_n1357_), .Y(ori_ori_n1361_));
  AOI220     o1312(.A0(ori_ori_n1361_), .A1(x3), .B0(ori_ori_n1021_), .B1(ori_ori_n342_), .Y(ori_ori_n1362_));
  AOI220     o1313(.A0(ori_ori_n1067_), .A1(ori_ori_n111_), .B0(ori_ori_n796_), .B1(ori_ori_n701_), .Y(ori_ori_n1363_));
  AOI210     o1314(.A0(ori_ori_n1363_), .A1(x7), .B0(ori_ori_n291_), .Y(ori_ori_n1364_));
  NA3        o1315(.A(ori_ori_n1018_), .B(ori_ori_n343_), .C(ori_ori_n100_), .Y(ori_ori_n1365_));
  NO2        o1316(.A(ori_ori_n1365_), .B(ori_ori_n834_), .Y(ori_ori_n1366_));
  NO3        o1317(.A(ori_ori_n230_), .B(ori_ori_n1366_), .C(ori_ori_n1364_), .Y(ori_ori_n1367_));
  OAI210     o1318(.A0(ori_ori_n1362_), .A1(ori_ori_n730_), .B0(ori_ori_n1367_), .Y(ori_ori_n1368_));
  NO2        o1319(.A(ori_ori_n486_), .B(ori_ori_n65_), .Y(ori_ori_n1369_));
  OAI220     o1320(.A0(ori_ori_n1369_), .A1(ori_ori_n1332_), .B0(ori_ori_n278_), .B1(ori_ori_n777_), .Y(ori_ori_n1370_));
  NA2        o1321(.A(ori_ori_n1370_), .B(ori_ori_n56_), .Y(ori_ori_n1371_));
  NO2        o1322(.A(ori_ori_n1371_), .B(ori_ori_n54_), .Y(ori_ori_n1372_));
  OAI210     o1323(.A0(ori_ori_n1372_), .A1(ori_ori_n1368_), .B0(x8), .Y(ori_ori_n1373_));
  NA4        o1324(.A(ori_ori_n1373_), .B(ori_ori_n1356_), .C(ori_ori_n1347_), .D(ori_ori_n1337_), .Y(ori20));
  NA4        o1325(.A(ori_ori_n352_), .B(ori_ori_n251_), .C(ori_ori_n341_), .D(ori_ori_n60_), .Y(ori_ori_n1375_));
  NO2        o1326(.A(ori_ori_n1375_), .B(ori_ori_n83_), .Y(ori_ori_n1376_));
  OAI210     o1327(.A0(x5), .A1(ori_ori_n601_), .B0(x4), .Y(ori_ori_n1377_));
  OAI210     o1328(.A0(ori_ori_n1377_), .A1(ori_ori_n1376_), .B0(ori_ori_n942_), .Y(ori_ori_n1378_));
  NAi21      o1329(.An(ori_ori_n482_), .B(ori_ori_n361_), .Y(ori_ori_n1379_));
  NA3        o1330(.A(ori_ori_n1379_), .B(ori_ori_n856_), .C(ori_ori_n824_), .Y(ori_ori_n1380_));
  NA3        o1331(.A(ori_ori_n941_), .B(ori_ori_n251_), .C(ori_ori_n515_), .Y(ori_ori_n1381_));
  AOI210     o1332(.A0(ori_ori_n1381_), .A1(ori_ori_n1380_), .B0(ori_ori_n1098_), .Y(ori_ori_n1382_));
  NO2        o1333(.A(ori_ori_n644_), .B(ori_ori_n844_), .Y(ori_ori_n1383_));
  NOi31      o1334(.An(ori_ori_n1383_), .B(ori_ori_n1000_), .C(ori_ori_n462_), .Y(ori_ori_n1384_));
  OAI210     o1335(.A0(ori_ori_n1384_), .A1(ori_ori_n1382_), .B0(x3), .Y(ori_ori_n1385_));
  NA2        o1336(.A(ori_ori_n287_), .B(ori_ori_n86_), .Y(ori_ori_n1386_));
  NA2        o1337(.A(ori_ori_n294_), .B(ori_ori_n98_), .Y(ori_ori_n1387_));
  NO2        o1338(.A(ori_ori_n590_), .B(ori_ori_n536_), .Y(ori_ori_n1388_));
  NA2        o1339(.A(ori_ori_n825_), .B(ori_ori_n50_), .Y(ori_ori_n1389_));
  NO3        o1340(.A(ori_ori_n1389_), .B(ori_ori_n329_), .C(ori_ori_n210_), .Y(ori_ori_n1390_));
  NA3        o1341(.A(ori_ori_n302_), .B(ori_ori_n219_), .C(ori_ori_n689_), .Y(ori_ori_n1391_));
  NO2        o1342(.A(ori_ori_n1391_), .B(ori_ori_n596_), .Y(ori_ori_n1392_));
  AOI210     o1343(.A0(ori_ori_n1390_), .A1(ori_ori_n1388_), .B0(ori_ori_n1392_), .Y(ori_ori_n1393_));
  NA3        o1344(.A(ori_ori_n1393_), .B(ori_ori_n1385_), .C(ori_ori_n1378_), .Y(ori21));
  OAI210     o1345(.A0(ori_ori_n364_), .A1(ori_ori_n54_), .B0(x7), .Y(ori_ori_n1395_));
  OAI220     o1346(.A0(ori_ori_n1395_), .A1(ori_ori_n1090_), .B0(ori_ori_n899_), .B1(ori_ori_n87_), .Y(ori_ori_n1396_));
  NA2        o1347(.A(ori_ori_n1396_), .B(ori_ori_n75_), .Y(ori_ori_n1397_));
  NA2        o1348(.A(ori_ori_n263_), .B(ori_ori_n741_), .Y(ori_ori_n1398_));
  AOI220     o1349(.A0(ori_ori_n1398_), .A1(ori_ori_n280_), .B0(ori_ori_n501_), .B1(ori_ori_n57_), .Y(ori_ori_n1399_));
  NA2        o1350(.A(ori_ori_n470_), .B(ori_ori_n407_), .Y(ori_ori_n1400_));
  NA3        o1351(.A(ori_ori_n1400_), .B(ori_ori_n1165_), .C(ori_ori_n56_), .Y(ori_ori_n1401_));
  NO2        o1352(.A(ori_ori_n666_), .B(ori_ori_n386_), .Y(ori_ori_n1402_));
  NO3        o1353(.A(ori_ori_n1402_), .B(ori_ori_n618_), .C(ori_ori_n228_), .Y(ori_ori_n1403_));
  NOi31      o1354(.An(ori_ori_n174_), .B(ori_ori_n560_), .C(ori_ori_n929_), .Y(ori_ori_n1404_));
  NO4        o1355(.A(ori_ori_n1404_), .B(ori_ori_n1403_), .C(ori_ori_n1401_), .D(ori_ori_n1399_), .Y(ori_ori_n1405_));
  NO3        o1356(.A(ori_ori_n386_), .B(ori_ori_n249_), .C(ori_ori_n52_), .Y(ori_ori_n1406_));
  OA210      o1357(.A0(ori_ori_n1406_), .A1(ori_ori_n766_), .B0(x3), .Y(ori_ori_n1407_));
  OAI210     o1358(.A0(ori_ori_n2188_), .A1(ori_ori_n520_), .B0(ori_ori_n304_), .Y(ori_ori_n1408_));
  NO2        o1359(.A(ori_ori_n67_), .B(x2), .Y(ori_ori_n1409_));
  OAI210     o1360(.A0(ori_ori_n159_), .A1(x0), .B0(ori_ori_n1409_), .Y(ori_ori_n1410_));
  NA3        o1361(.A(ori_ori_n132_), .B(ori_ori_n1410_), .C(ori_ori_n1408_), .Y(ori_ori_n1411_));
  OAI210     o1362(.A0(ori_ori_n1411_), .A1(ori_ori_n1407_), .B0(x8), .Y(ori_ori_n1412_));
  NO3        o1363(.A(ori_ori_n665_), .B(ori_ori_n549_), .C(ori_ori_n516_), .Y(ori_ori_n1413_));
  NA2        o1364(.A(ori_ori_n55_), .B(ori_ori_n50_), .Y(ori_ori_n1414_));
  BUFFER     o1365(.A(ori_ori_n1414_), .Y(ori_ori_n1415_));
  NO2        o1366(.A(ori_ori_n220_), .B(ori_ori_n1415_), .Y(ori_ori_n1416_));
  INV        o1367(.A(x4), .Y(ori_ori_n1417_));
  NO3        o1368(.A(ori_ori_n1417_), .B(ori_ori_n1416_), .C(ori_ori_n1413_), .Y(ori_ori_n1418_));
  AO220      o1369(.A0(ori_ori_n1418_), .A1(ori_ori_n1412_), .B0(ori_ori_n1405_), .B1(ori_ori_n1397_), .Y(ori_ori_n1419_));
  AO220      o1370(.A0(ori_ori_n561_), .A1(ori_ori_n291_), .B0(ori_ori_n521_), .B1(x8), .Y(ori_ori_n1420_));
  NO2        o1371(.A(ori_ori_n742_), .B(x0), .Y(ori_ori_n1421_));
  NO3        o1372(.A(ori_ori_n1421_), .B(ori_ori_n479_), .C(ori_ori_n2164_), .Y(ori_ori_n1422_));
  NO2        o1373(.A(ori_ori_n146_), .B(x2), .Y(ori_ori_n1423_));
  NO3        o1374(.A(ori_ori_n340_), .B(ori_ori_n231_), .C(ori_ori_n166_), .Y(ori_ori_n1424_));
  INV        o1375(.A(ori_ori_n1424_), .Y(ori_ori_n1425_));
  OAI210     o1376(.A0(ori_ori_n1422_), .A1(ori_ori_n359_), .B0(ori_ori_n1425_), .Y(ori_ori_n1426_));
  AOI220     o1377(.A0(ori_ori_n1426_), .A1(x5), .B0(ori_ori_n1420_), .B1(ori_ori_n644_), .Y(ori_ori_n1427_));
  AOI210     o1378(.A0(ori_ori_n1427_), .A1(ori_ori_n1419_), .B0(ori_ori_n68_), .Y(ori_ori_n1428_));
  NO2        o1379(.A(ori_ori_n788_), .B(ori_ori_n153_), .Y(ori_ori_n1429_));
  NOi41      o1380(.An(ori_ori_n1212_), .B(ori_ori_n1270_), .C(ori_ori_n987_), .D(ori_ori_n734_), .Y(ori_ori_n1430_));
  NA2        o1381(.A(ori_ori_n1430_), .B(ori_ori_n1429_), .Y(ori_ori_n1431_));
  NO2        o1382(.A(ori_ori_n75_), .B(x4), .Y(ori_ori_n1432_));
  OAI210     o1383(.A0(ori_ori_n261_), .A1(ori_ori_n145_), .B0(ori_ori_n1432_), .Y(ori_ori_n1433_));
  OAI210     o1384(.A0(ori_ori_n366_), .A1(ori_ori_n378_), .B0(ori_ori_n210_), .Y(ori_ori_n1434_));
  NO2        o1385(.A(ori_ori_n233_), .B(ori_ori_n50_), .Y(ori_ori_n1435_));
  INV        o1386(.A(ori_ori_n1435_), .Y(ori_ori_n1436_));
  NA2        o1387(.A(ori_ori_n1436_), .B(ori_ori_n1434_), .Y(ori_ori_n1437_));
  AOI210     o1388(.A0(ori_ori_n1433_), .A1(ori_ori_n1431_), .B0(ori_ori_n1437_), .Y(ori_ori_n1438_));
  NA2        o1389(.A(ori_ori_n656_), .B(ori_ori_n482_), .Y(ori_ori_n1439_));
  AO210      o1390(.A0(ori_ori_n1439_), .A1(ori_ori_n834_), .B0(ori_ori_n50_), .Y(ori_ori_n1440_));
  NO2        o1391(.A(ori_ori_n1379_), .B(ori_ori_n1030_), .Y(ori_ori_n1441_));
  AOI220     o1392(.A0(ori_ori_n1441_), .A1(ori_ori_n993_), .B0(ori_ori_n1119_), .B1(ori_ori_n896_), .Y(ori_ori_n1442_));
  AOI210     o1393(.A0(ori_ori_n1442_), .A1(ori_ori_n1440_), .B0(ori_ori_n100_), .Y(ori_ori_n1443_));
  NA2        o1394(.A(ori_ori_n270_), .B(ori_ori_n98_), .Y(ori_ori_n1444_));
  NA2        o1395(.A(ori_ori_n776_), .B(ori_ori_n55_), .Y(ori_ori_n1445_));
  NO2        o1396(.A(ori_ori_n1445_), .B(ori_ori_n1444_), .Y(ori_ori_n1446_));
  NO2        o1397(.A(ori_ori_n593_), .B(ori_ori_n900_), .Y(ori_ori_n1447_));
  NO4        o1398(.A(ori_ori_n1447_), .B(ori_ori_n1446_), .C(ori_ori_n1443_), .D(ori_ori_n1438_), .Y(ori_ori_n1448_));
  NO2        o1399(.A(ori_ori_n1448_), .B(x6), .Y(ori_ori_n1449_));
  OA220      o1400(.A0(x1), .A1(ori_ori_n388_), .B0(ori_ori_n411_), .B1(ori_ori_n644_), .Y(ori_ori_n1450_));
  NA3        o1401(.A(ori_ori_n55_), .B(x2), .C(x0), .Y(ori_ori_n1451_));
  NA2        o1402(.A(ori_ori_n1450_), .B(ori_ori_n56_), .Y(ori_ori_n1452_));
  NA2        o1403(.A(ori_ori_n1452_), .B(ori_ori_n105_), .Y(ori_ori_n1453_));
  NO2        o1404(.A(ori_ori_n543_), .B(ori_ori_n276_), .Y(ori_ori_n1454_));
  INV        o1405(.A(ori_ori_n1454_), .Y(ori_ori_n1455_));
  NO2        o1406(.A(ori_ori_n1455_), .B(ori_ori_n100_), .Y(ori_ori_n1456_));
  NA2        o1407(.A(ori_ori_n613_), .B(ori_ori_n78_), .Y(ori_ori_n1457_));
  NO2        o1408(.A(ori_ori_n1445_), .B(ori_ori_n1444_), .Y(ori_ori_n1458_));
  OAI210     o1409(.A0(ori_ori_n1458_), .A1(ori_ori_n1456_), .B0(x1), .Y(ori_ori_n1459_));
  NO2        o1410(.A(ori_ori_n58_), .B(ori_ori_n98_), .Y(ori_ori_n1460_));
  NO4        o1411(.A(ori_ori_n1444_), .B(ori_ori_n832_), .C(ori_ori_n590_), .D(ori_ori_n50_), .Y(ori_ori_n1461_));
  AOI210     o1412(.A0(ori_ori_n1460_), .A1(ori_ori_n1309_), .B0(ori_ori_n1461_), .Y(ori_ori_n1462_));
  NA3        o1413(.A(ori_ori_n1462_), .B(ori_ori_n1459_), .C(ori_ori_n1453_), .Y(ori_ori_n1463_));
  NO3        o1414(.A(ori_ori_n1463_), .B(ori_ori_n1449_), .C(ori_ori_n1428_), .Y(ori22));
  NO2        o1415(.A(ori_ori_n486_), .B(ori_ori_n610_), .Y(ori_ori_n1465_));
  AOI210     o1416(.A0(x5), .A1(x2), .B0(x8), .Y(ori_ori_n1466_));
  OAI220     o1417(.A0(x0), .A1(ori_ori_n1465_), .B0(x5), .B1(ori_ori_n359_), .Y(ori_ori_n1467_));
  NA2        o1418(.A(ori_ori_n515_), .B(ori_ori_n83_), .Y(ori_ori_n1468_));
  NA2        o1419(.A(ori_ori_n246_), .B(ori_ori_n74_), .Y(ori_ori_n1469_));
  OA220      o1420(.A0(ori_ori_n1469_), .A1(ori_ori_n1468_), .B0(ori_ori_n727_), .B1(ori_ori_n875_), .Y(ori_ori_n1470_));
  NO3        o1421(.A(ori_ori_n1058_), .B(ori_ori_n83_), .C(x0), .Y(ori_ori_n1471_));
  NO2        o1422(.A(ori_ori_n2168_), .B(ori_ori_n1471_), .Y(ori_ori_n1472_));
  OAI210     o1423(.A0(ori_ori_n1470_), .A1(ori_ori_n179_), .B0(ori_ori_n1472_), .Y(ori_ori_n1473_));
  AOI210     o1424(.A0(ori_ori_n1467_), .A1(ori_ori_n53_), .B0(ori_ori_n1473_), .Y(ori_ori_n1474_));
  NA2        o1425(.A(ori_ori_n510_), .B(ori_ori_n223_), .Y(ori_ori_n1475_));
  NO3        o1426(.A(ori_ori_n437_), .B(ori_ori_n238_), .C(ori_ori_n194_), .Y(ori_ori_n1476_));
  NO2        o1427(.A(ori_ori_n411_), .B(ori_ori_n235_), .Y(ori_ori_n1477_));
  NA3        o1428(.A(ori_ori_n55_), .B(ori_ori_n68_), .C(x0), .Y(ori_ori_n1478_));
  OAI220     o1429(.A0(ori_ori_n1478_), .A1(ori_ori_n900_), .B0(ori_ori_n329_), .B1(ori_ori_n193_), .Y(ori_ori_n1479_));
  NO2        o1430(.A(ori_ori_n1479_), .B(x4), .Y(ori_ori_n1480_));
  NA2        o1431(.A(ori_ori_n233_), .B(ori_ori_n1480_), .Y(ori_ori_n1481_));
  AOI210     o1432(.A0(x8), .A1(ori_ori_n98_), .B0(ori_ori_n1481_), .Y(ori_ori_n1482_));
  OAI210     o1433(.A0(ori_ori_n691_), .A1(ori_ori_n146_), .B0(ori_ori_n813_), .Y(ori_ori_n1483_));
  OAI210     o1434(.A0(ori_ori_n1483_), .A1(ori_ori_n56_), .B0(ori_ori_n542_), .Y(ori_ori_n1484_));
  OA210      o1435(.A0(ori_ori_n1482_), .A1(ori_ori_n1474_), .B0(ori_ori_n1484_), .Y(ori_ori_n1485_));
  OAI210     o1436(.A0(ori_ori_n1002_), .A1(ori_ori_n612_), .B0(ori_ori_n608_), .Y(ori_ori_n1486_));
  NO2        o1437(.A(ori_ori_n317_), .B(x0), .Y(ori_ori_n1487_));
  NA3        o1438(.A(ori_ori_n1487_), .B(ori_ori_n312_), .C(ori_ori_n56_), .Y(ori_ori_n1488_));
  AOI210     o1439(.A0(ori_ori_n1488_), .A1(ori_ori_n1486_), .B0(ori_ori_n359_), .Y(ori_ori_n1489_));
  NO3        o1440(.A(ori_ori_n154_), .B(ori_ori_n146_), .C(ori_ori_n60_), .Y(ori_ori_n1490_));
  OAI210     o1441(.A0(ori_ori_n1490_), .A1(ori_ori_n373_), .B0(ori_ori_n100_), .Y(ori_ori_n1491_));
  NA2        o1442(.A(ori_ori_n129_), .B(ori_ori_n677_), .Y(ori_ori_n1492_));
  NA2        o1443(.A(ori_ori_n371_), .B(x3), .Y(ori_ori_n1493_));
  NAi31      o1444(.An(ori_ori_n1493_), .B(ori_ori_n1492_), .C(ori_ori_n1324_), .Y(ori_ori_n1494_));
  NO3        o1445(.A(ori_ori_n742_), .B(ori_ori_n410_), .C(ori_ori_n100_), .Y(ori_ori_n1495_));
  NO2        o1446(.A(ori_ori_n926_), .B(ori_ori_n130_), .Y(ori_ori_n1496_));
  NO3        o1447(.A(ori_ori_n779_), .B(ori_ori_n369_), .C(ori_ori_n275_), .Y(ori_ori_n1497_));
  AOI220     o1448(.A0(ori_ori_n1497_), .A1(ori_ori_n1496_), .B0(ori_ori_n1495_), .B1(ori_ori_n1487_), .Y(ori_ori_n1498_));
  NA3        o1449(.A(ori_ori_n369_), .B(ori_ori_n86_), .C(ori_ori_n78_), .Y(ori_ori_n1499_));
  AOI210     o1450(.A0(ori_ori_n538_), .A1(ori_ori_n405_), .B0(ori_ori_n434_), .Y(ori_ori_n1500_));
  NA2        o1451(.A(ori_ori_n1004_), .B(x3), .Y(ori_ori_n1501_));
  OAI210     o1452(.A0(ori_ori_n1501_), .A1(ori_ori_n1500_), .B0(ori_ori_n1499_), .Y(ori_ori_n1502_));
  NA3        o1453(.A(ori_ori_n56_), .B(ori_ori_n50_), .C(x0), .Y(ori_ori_n1503_));
  NOi21      o1454(.An(ori_ori_n80_), .B(ori_ori_n629_), .Y(ori_ori_n1504_));
  NA3        o1455(.A(x6), .B(x4), .C(ori_ori_n50_), .Y(ori_ori_n1505_));
  NA3        o1456(.A(ori_ori_n1505_), .B(ori_ori_n859_), .C(ori_ori_n239_), .Y(ori_ori_n1506_));
  OAI220     o1457(.A0(ori_ori_n1506_), .A1(ori_ori_n1504_), .B0(ori_ori_n902_), .B1(ori_ori_n1503_), .Y(ori_ori_n1507_));
  AOI220     o1458(.A0(ori_ori_n1507_), .A1(ori_ori_n908_), .B0(ori_ori_n1502_), .B1(ori_ori_n312_), .Y(ori_ori_n1508_));
  NA4        o1459(.A(ori_ori_n1508_), .B(ori_ori_n1498_), .C(ori_ori_n1494_), .D(ori_ori_n1491_), .Y(ori_ori_n1509_));
  AOI210     o1460(.A0(ori_ori_n1509_), .A1(x7), .B0(ori_ori_n1489_), .Y(ori_ori_n1510_));
  OAI210     o1461(.A0(ori_ori_n1485_), .A1(x7), .B0(ori_ori_n1510_), .Y(ori23));
  NO3        o1462(.A(ori_ori_n727_), .B(ori_ori_n524_), .C(ori_ori_n427_), .Y(ori_ori_n1512_));
  NO3        o1463(.A(ori_ori_n826_), .B(ori_ori_n137_), .C(ori_ori_n106_), .Y(ori_ori_n1513_));
  AOI210     o1464(.A0(ori_ori_n1513_), .A1(ori_ori_n889_), .B0(ori_ori_n1512_), .Y(ori_ori_n1514_));
  INV        o1465(.A(ori_ori_n1514_), .Y(ori_ori_n1515_));
  NA2        o1466(.A(ori_ori_n1515_), .B(ori_ori_n55_), .Y(ori_ori_n1516_));
  NO2        o1467(.A(ori_ori_n832_), .B(ori_ori_n454_), .Y(ori_ori_n1517_));
  AO220      o1468(.A0(ori_ori_n1086_), .A1(ori_ori_n163_), .B0(ori_ori_n865_), .B1(ori_ori_n644_), .Y(ori_ori_n1518_));
  OAI210     o1469(.A0(ori_ori_n1518_), .A1(ori_ori_n1517_), .B0(ori_ori_n521_), .Y(ori_ori_n1519_));
  NA2        o1470(.A(ori_ori_n160_), .B(ori_ori_n153_), .Y(ori_ori_n1520_));
  NA2        o1471(.A(ori_ori_n363_), .B(ori_ori_n147_), .Y(ori_ori_n1521_));
  AOI210     o1472(.A0(ori_ori_n1521_), .A1(ori_ori_n1520_), .B0(ori_ori_n217_), .Y(ori_ori_n1522_));
  NA3        o1473(.A(ori_ori_n750_), .B(ori_ori_n378_), .C(ori_ori_n233_), .Y(ori_ori_n1523_));
  AOI210     o1474(.A0(ori_ori_n1523_), .A1(ori_ori_n439_), .B0(ori_ori_n343_), .Y(ori_ori_n1524_));
  OAI210     o1475(.A0(ori_ori_n1524_), .A1(ori_ori_n1522_), .B0(ori_ori_n270_), .Y(ori_ori_n1525_));
  NA2        o1476(.A(ori_ori_n800_), .B(ori_ori_n131_), .Y(ori_ori_n1526_));
  NA4        o1477(.A(ori_ori_n1526_), .B(ori_ori_n1525_), .C(ori_ori_n1519_), .D(ori_ori_n1516_), .Y(ori24));
  NO2        o1478(.A(ori_ori_n221_), .B(x1), .Y(ori_ori_n1528_));
  NA2        o1479(.A(ori_ori_n302_), .B(ori_ori_n431_), .Y(ori_ori_n1529_));
  NAi21      o1480(.An(ori_ori_n1528_), .B(ori_ori_n1529_), .Y(ori_ori_n1530_));
  NO3        o1481(.A(ori_ori_n475_), .B(ori_ori_n604_), .C(ori_ori_n143_), .Y(ori_ori_n1531_));
  AOI210     o1482(.A0(ori_ori_n1530_), .A1(ori_ori_n86_), .B0(ori_ori_n1531_), .Y(ori_ori_n1532_));
  NA2        o1483(.A(ori_ori_n93_), .B(x8), .Y(ori_ori_n1533_));
  AN2        o1484(.A(ori_ori_n1077_), .B(x3), .Y(ori_ori_n1534_));
  NA2        o1485(.A(ori_ori_n405_), .B(x8), .Y(ori_ori_n1535_));
  NA2        o1486(.A(ori_ori_n591_), .B(ori_ori_n114_), .Y(ori_ori_n1536_));
  OAI220     o1487(.A0(ori_ori_n1536_), .A1(ori_ori_n1219_), .B0(ori_ori_n1535_), .B1(x1), .Y(ori_ori_n1537_));
  AOI220     o1488(.A0(ori_ori_n1537_), .A1(ori_ori_n1435_), .B0(ori_ori_n1534_), .B1(ori_ori_n889_), .Y(ori_ori_n1538_));
  OAI210     o1489(.A0(ori_ori_n1533_), .A1(ori_ori_n1532_), .B0(ori_ori_n1538_), .Y(ori25));
  NA2        o1490(.A(ori_ori_n1354_), .B(ori_ori_n1010_), .Y(ori_ori_n1540_));
  AOI210     o1491(.A0(ori_ori_n1540_), .A1(x7), .B0(ori_ori_n599_), .Y(ori_ori_n1541_));
  NO3        o1492(.A(ori_ori_n895_), .B(ori_ori_n132_), .C(ori_ori_n75_), .Y(ori_ori_n1542_));
  OAI210     o1493(.A0(ori_ori_n179_), .A1(ori_ori_n246_), .B0(ori_ori_n295_), .Y(ori_ori_n1543_));
  OAI210     o1494(.A0(ori_ori_n1543_), .A1(ori_ori_n1542_), .B0(ori_ori_n1008_), .Y(ori_ori_n1544_));
  NO2        o1495(.A(ori_ori_n1175_), .B(ori_ori_n399_), .Y(ori_ori_n1545_));
  NO3        o1496(.A(ori_ori_n1545_), .B(ori_ori_n466_), .C(ori_ori_n90_), .Y(ori_ori_n1546_));
  OAI210     o1497(.A0(ori_ori_n516_), .A1(ori_ori_n1546_), .B0(ori_ori_n565_), .Y(ori_ori_n1547_));
  AOI210     o1498(.A0(ori_ori_n1477_), .A1(ori_ori_n967_), .B0(ori_ori_n1265_), .Y(ori_ori_n1548_));
  NA3        o1499(.A(ori_ori_n1548_), .B(ori_ori_n1547_), .C(ori_ori_n1544_), .Y(ori_ori_n1549_));
  AO210      o1500(.A0(ori_ori_n1549_), .A1(ori_ori_n98_), .B0(ori_ori_n1541_), .Y(ori26));
  NA2        o1501(.A(ori_ori_n664_), .B(ori_ori_n50_), .Y(ori_ori_n1551_));
  OAI220     o1502(.A0(ori_ori_n276_), .A1(ori_ori_n228_), .B0(ori_ori_n1551_), .B1(x7), .Y(ori_ori_n1552_));
  AOI220     o1503(.A0(ori_ori_n1552_), .A1(ori_ori_n86_), .B0(ori_ori_n1099_), .B1(ori_ori_n973_), .Y(ori_ori_n1553_));
  NA2        o1504(.A(ori_ori_n553_), .B(ori_ori_n510_), .Y(ori_ori_n1554_));
  OAI210     o1505(.A0(ori_ori_n561_), .A1(ori_ori_n553_), .B0(ori_ori_n644_), .Y(ori_ori_n1555_));
  AOI210     o1506(.A0(ori_ori_n1554_), .A1(ori_ori_n1020_), .B0(ori_ori_n1555_), .Y(ori_ori_n1556_));
  NA2        o1507(.A(ori_ori_n882_), .B(ori_ori_n516_), .Y(ori_ori_n1557_));
  NO2        o1508(.A(ori_ori_n1557_), .B(ori_ori_n1063_), .Y(ori_ori_n1558_));
  AOI210     o1509(.A0(ori_ori_n1496_), .A1(x5), .B0(ori_ori_n1558_), .Y(ori_ori_n1559_));
  NO2        o1510(.A(ori_ori_n926_), .B(ori_ori_n72_), .Y(ori_ori_n1560_));
  NA2        o1511(.A(ori_ori_n699_), .B(ori_ori_n159_), .Y(ori_ori_n1561_));
  NO2        o1512(.A(ori_ori_n1561_), .B(ori_ori_n471_), .Y(ori_ori_n1562_));
  AOI210     o1513(.A0(ori_ori_n1560_), .A1(ori_ori_n517_), .B0(ori_ori_n1562_), .Y(ori_ori_n1563_));
  OAI220     o1514(.A0(ori_ori_n1563_), .A1(ori_ori_n98_), .B0(ori_ori_n1559_), .B1(ori_ori_n53_), .Y(ori_ori_n1564_));
  NO2        o1515(.A(ori_ori_n122_), .B(x8), .Y(ori_ori_n1565_));
  NA2        o1516(.A(ori_ori_n1565_), .B(ori_ori_n111_), .Y(ori_ori_n1566_));
  NA2        o1517(.A(ori_ori_n644_), .B(x3), .Y(ori_ori_n1567_));
  NO2        o1518(.A(ori_ori_n1566_), .B(ori_ori_n1567_), .Y(ori_ori_n1568_));
  NO2        o1519(.A(ori_ori_n875_), .B(x3), .Y(ori_ori_n1569_));
  AOI210     o1520(.A0(ori_ori_n397_), .A1(ori_ori_n98_), .B0(ori_ori_n1569_), .Y(ori_ori_n1570_));
  NA3        o1521(.A(x1), .B(ori_ori_n51_), .C(ori_ori_n56_), .Y(ori_ori_n1571_));
  AOI210     o1522(.A0(ori_ori_n1388_), .A1(ori_ori_n903_), .B0(x0), .Y(ori_ori_n1572_));
  OAI210     o1523(.A0(ori_ori_n1571_), .A1(ori_ori_n1570_), .B0(ori_ori_n1572_), .Y(ori_ori_n1573_));
  NO4        o1524(.A(ori_ori_n1573_), .B(ori_ori_n1568_), .C(ori_ori_n1564_), .D(ori_ori_n1556_), .Y(ori_ori_n1574_));
  AOI210     o1525(.A0(x8), .A1(x6), .B0(x5), .Y(ori_ori_n1575_));
  AO220      o1526(.A0(ori_ori_n1575_), .A1(ori_ori_n133_), .B0(ori_ori_n524_), .B1(ori_ori_n129_), .Y(ori_ori_n1576_));
  NA2        o1527(.A(ori_ori_n1576_), .B(ori_ori_n398_), .Y(ori_ori_n1577_));
  NO2        o1528(.A(ori_ori_n654_), .B(ori_ori_n133_), .Y(ori_ori_n1578_));
  NA3        o1529(.A(ori_ori_n1578_), .B(ori_ori_n1409_), .C(ori_ori_n123_), .Y(ori_ori_n1579_));
  INV        o1530(.A(ori_ori_n359_), .Y(ori_ori_n1580_));
  OAI210     o1531(.A0(ori_ori_n1580_), .A1(ori_ori_n1135_), .B0(ori_ori_n397_), .Y(ori_ori_n1581_));
  NA4        o1532(.A(ori_ori_n2174_), .B(ori_ori_n1581_), .C(ori_ori_n1579_), .D(ori_ori_n1577_), .Y(ori_ori_n1582_));
  NO2        o1533(.A(ori_ori_n2172_), .B(ori_ori_n106_), .Y(ori_ori_n1583_));
  NA3        o1534(.A(ori_ori_n701_), .B(ori_ori_n875_), .C(x7), .Y(ori_ori_n1584_));
  AOI210     o1535(.A0(ori_ori_n306_), .A1(ori_ori_n196_), .B0(ori_ori_n1584_), .Y(ori_ori_n1585_));
  NO2        o1536(.A(ori_ori_n782_), .B(ori_ori_n276_), .Y(ori_ori_n1586_));
  NO3        o1537(.A(ori_ori_n1586_), .B(ori_ori_n1585_), .C(ori_ori_n1583_), .Y(ori_ori_n1587_));
  NA3        o1538(.A(ori_ori_n591_), .B(ori_ori_n173_), .C(ori_ori_n824_), .Y(ori_ori_n1588_));
  NA2        o1539(.A(ori_ori_n1588_), .B(x7), .Y(ori_ori_n1589_));
  INV        o1540(.A(ori_ori_n129_), .Y(ori_ori_n1590_));
  OAI210     o1541(.A0(ori_ori_n1590_), .A1(ori_ori_n1208_), .B0(x0), .Y(ori_ori_n1591_));
  AOI210     o1542(.A0(ori_ori_n1589_), .A1(ori_ori_n1196_), .B0(ori_ori_n1591_), .Y(ori_ori_n1592_));
  OAI210     o1543(.A0(ori_ori_n1587_), .A1(ori_ori_n53_), .B0(ori_ori_n1592_), .Y(ori_ori_n1593_));
  AOI210     o1544(.A0(ori_ori_n1582_), .A1(x4), .B0(ori_ori_n1593_), .Y(ori_ori_n1594_));
  OA220      o1545(.A0(ori_ori_n1594_), .A1(ori_ori_n1574_), .B0(ori_ori_n1553_), .B1(ori_ori_n99_), .Y(ori27));
  NA2        o1546(.A(ori_ori_n976_), .B(ori_ori_n397_), .Y(ori_ori_n1596_));
  NO2        o1547(.A(ori_ori_n1596_), .B(ori_ori_n271_), .Y(ori_ori_n1597_));
  NA2        o1548(.A(ori_ori_n796_), .B(ori_ori_n701_), .Y(ori_ori_n1598_));
  NA3        o1549(.A(ori_ori_n707_), .B(ori_ori_n326_), .C(ori_ori_n883_), .Y(ori_ori_n1599_));
  AOI210     o1550(.A0(ori_ori_n1599_), .A1(ori_ori_n1598_), .B0(ori_ori_n196_), .Y(ori_ori_n1600_));
  OAI210     o1551(.A0(ori_ori_n1600_), .A1(ori_ori_n1597_), .B0(ori_ori_n611_), .Y(ori_ori_n1601_));
  XO2        o1552(.A(x8), .B(x4), .Y(ori_ori_n1602_));
  NO3        o1553(.A(ori_ori_n1602_), .B(ori_ori_n397_), .C(ori_ori_n154_), .Y(ori_ori_n1603_));
  OA210      o1554(.A0(ori_ori_n1603_), .A1(ori_ori_n1064_), .B0(ori_ori_n249_), .Y(ori_ori_n1604_));
  NO2        o1555(.A(ori_ori_n354_), .B(ori_ori_n150_), .Y(ori_ori_n1605_));
  OAI210     o1556(.A0(ori_ori_n1605_), .A1(ori_ori_n1604_), .B0(ori_ori_n954_), .Y(ori_ori_n1606_));
  AOI210     o1557(.A0(ori_ori_n561_), .A1(ori_ori_n56_), .B0(ori_ori_n1560_), .Y(ori_ori_n1607_));
  OAI220     o1558(.A0(ori_ori_n1607_), .A1(ori_ori_n1063_), .B0(ori_ori_n1019_), .B1(ori_ori_n188_), .Y(ori_ori_n1608_));
  NA2        o1559(.A(ori_ori_n1608_), .B(ori_ori_n470_), .Y(ori_ori_n1609_));
  NA3        o1560(.A(ori_ori_n1609_), .B(ori_ori_n1606_), .C(ori_ori_n1601_), .Y(ori28));
  OAI210     o1561(.A0(ori_ori_n57_), .A1(ori_ori_n1079_), .B0(ori_ori_n516_), .Y(ori_ori_n1611_));
  NA3        o1562(.A(ori_ori_n1010_), .B(ori_ori_n776_), .C(x7), .Y(ori_ori_n1612_));
  NA3        o1563(.A(ori_ori_n434_), .B(ori_ori_n75_), .C(ori_ori_n536_), .Y(ori_ori_n1613_));
  NA3        o1564(.A(ori_ori_n1613_), .B(ori_ori_n1612_), .C(ori_ori_n1611_), .Y(ori_ori_n1614_));
  NA2        o1565(.A(ori_ori_n1058_), .B(ori_ori_n395_), .Y(ori_ori_n1615_));
  NA3        o1566(.A(ori_ori_n1615_), .B(ori_ori_n1185_), .C(ori_ori_n368_), .Y(ori_ori_n1616_));
  NO2        o1567(.A(ori_ori_n279_), .B(x4), .Y(ori_ori_n1617_));
  AOI220     o1568(.A0(ori_ori_n1617_), .A1(ori_ori_n1569_), .B0(ori_ori_n955_), .B1(ori_ori_n595_), .Y(ori_ori_n1618_));
  NA2        o1569(.A(ori_ori_n1618_), .B(ori_ori_n1616_), .Y(ori_ori_n1619_));
  NO2        o1570(.A(ori_ori_n1058_), .B(ori_ori_n1036_), .Y(ori_ori_n1620_));
  NO4        o1571(.A(x6), .B(ori_ori_n56_), .C(x2), .D(x0), .Y(ori_ori_n1621_));
  OAI210     o1572(.A0(ori_ori_n1621_), .A1(ori_ori_n1620_), .B0(ori_ori_n896_), .Y(ori_ori_n1622_));
  NA2        o1573(.A(ori_ori_n1004_), .B(ori_ori_n98_), .Y(ori_ori_n1623_));
  NA2        o1574(.A(ori_ori_n922_), .B(ori_ori_n97_), .Y(ori_ori_n1624_));
  OAI210     o1575(.A0(ori_ori_n1624_), .A1(ori_ori_n1623_), .B0(ori_ori_n1622_), .Y(ori_ori_n1625_));
  OAI210     o1576(.A0(ori_ori_n1625_), .A1(ori_ori_n1619_), .B0(x7), .Y(ori_ori_n1626_));
  NO2        o1577(.A(ori_ori_n345_), .B(x7), .Y(ori_ori_n1627_));
  NO3        o1578(.A(ori_ori_n359_), .B(ori_ori_n244_), .C(ori_ori_n112_), .Y(ori_ori_n1628_));
  OAI210     o1579(.A0(ori_ori_n750_), .A1(ori_ori_n235_), .B0(ori_ori_n78_), .Y(ori_ori_n1629_));
  OAI220     o1580(.A0(ori_ori_n1629_), .A1(ori_ori_n1628_), .B0(ori_ori_n1627_), .B1(ori_ori_n101_), .Y(ori_ori_n1630_));
  AOI210     o1581(.A0(ori_ori_n416_), .A1(ori_ori_n50_), .B0(ori_ori_n449_), .Y(ori_ori_n1631_));
  AOI210     o1582(.A0(ori_ori_n1631_), .A1(ori_ori_n1630_), .B0(ori_ori_n57_), .Y(ori_ori_n1632_));
  AOI210     o1583(.A0(ori_ori_n1175_), .A1(ori_ori_n594_), .B0(ori_ori_n405_), .Y(ori_ori_n1633_));
  OAI210     o1584(.A0(ori_ori_n1633_), .A1(ori_ori_n132_), .B0(x1), .Y(ori_ori_n1634_));
  NO2        o1585(.A(ori_ori_n1634_), .B(ori_ori_n1632_), .Y(ori_ori_n1635_));
  AOI210     o1586(.A0(ori_ori_n1341_), .A1(ori_ori_n359_), .B0(ori_ori_n589_), .Y(ori_ori_n1636_));
  NO2        o1587(.A(ori_ori_n359_), .B(x5), .Y(ori_ori_n1637_));
  NO2        o1588(.A(ori_ori_n1637_), .B(ori_ori_n208_), .Y(ori_ori_n1638_));
  NO2        o1589(.A(ori_ori_n1638_), .B(ori_ori_n1636_), .Y(ori_ori_n1639_));
  NOi21      o1590(.An(ori_ori_n613_), .B(ori_ori_n865_), .Y(ori_ori_n1640_));
  NA3        o1591(.A(ori_ori_n1640_), .B(ori_ori_n922_), .C(ori_ori_n750_), .Y(ori_ori_n1641_));
  OAI210     o1592(.A0(ori_ori_n1146_), .A1(ori_ori_n1414_), .B0(ori_ori_n1641_), .Y(ori_ori_n1642_));
  OAI210     o1593(.A0(ori_ori_n1642_), .A1(ori_ori_n1639_), .B0(ori_ori_n954_), .Y(ori_ori_n1643_));
  NO2        o1594(.A(ori_ori_n601_), .B(x6), .Y(ori_ori_n1644_));
  NO2        o1595(.A(ori_ori_n274_), .B(x4), .Y(ori_ori_n1645_));
  AOI220     o1596(.A0(ori_ori_n1645_), .A1(ori_ori_n326_), .B0(ori_ori_n1644_), .B1(x4), .Y(ori_ori_n1646_));
  NO3        o1597(.A(ori_ori_n1646_), .B(ori_ori_n291_), .C(x5), .Y(ori_ori_n1647_));
  INV        o1598(.A(ori_ori_n613_), .Y(ori_ori_n1648_));
  NA2        o1599(.A(ori_ori_n1648_), .B(ori_ori_n397_), .Y(ori_ori_n1649_));
  AOI220     o1600(.A0(ori_ori_n587_), .A1(ori_ori_n631_), .B0(ori_ori_n432_), .B1(ori_ori_n218_), .Y(ori_ori_n1650_));
  AOI210     o1601(.A0(ori_ori_n1650_), .A1(ori_ori_n1649_), .B0(ori_ori_n233_), .Y(ori_ori_n1651_));
  NO3        o1602(.A(ori_ori_n1651_), .B(ori_ori_n1647_), .C(x1), .Y(ori_ori_n1652_));
  AOI220     o1603(.A0(ori_ori_n1652_), .A1(ori_ori_n1643_), .B0(ori_ori_n1635_), .B1(ori_ori_n1626_), .Y(ori_ori_n1653_));
  AOI210     o1604(.A0(ori_ori_n1614_), .A1(x3), .B0(ori_ori_n1653_), .Y(ori29));
  NA2        o1605(.A(ori_ori_n487_), .B(ori_ori_n626_), .Y(ori_ori_n1655_));
  INV        o1606(.A(ori_ori_n896_), .Y(ori_ori_n1656_));
  OR2        o1607(.A(ori_ori_n994_), .B(ori_ori_n1656_), .Y(ori_ori_n1657_));
  AOI210     o1608(.A0(ori_ori_n164_), .A1(ori_ori_n151_), .B0(ori_ori_n613_), .Y(ori_ori_n1658_));
  AOI210     o1609(.A0(ori_ori_n1200_), .A1(ori_ori_n75_), .B0(ori_ori_n1658_), .Y(ori_ori_n1659_));
  NA3        o1610(.A(ori_ori_n1659_), .B(ori_ori_n1657_), .C(ori_ori_n1655_), .Y(ori_ori_n1660_));
  NO3        o1611(.A(ori_ori_n589_), .B(ori_ori_n973_), .C(ori_ori_n50_), .Y(ori_ori_n1661_));
  NO3        o1612(.A(ori_ori_n1661_), .B(ori_ori_n1057_), .C(ori_ori_n487_), .Y(ori_ori_n1662_));
  NA2        o1613(.A(ori_ori_n592_), .B(x0), .Y(ori_ori_n1663_));
  OAI210     o1614(.A0(ori_ori_n1662_), .A1(ori_ori_n475_), .B0(ori_ori_n1663_), .Y(ori_ori_n1664_));
  AOI210     o1615(.A0(ori_ori_n1660_), .A1(x6), .B0(ori_ori_n1664_), .Y(ori_ori_n1665_));
  OAI210     o1616(.A0(x8), .A1(x4), .B0(x5), .Y(ori_ori_n1666_));
  INV        o1617(.A(ori_ori_n1666_), .Y(ori_ori_n1667_));
  NA2        o1618(.A(ori_ori_n274_), .B(ori_ori_n135_), .Y(ori_ori_n1668_));
  NA3        o1619(.A(ori_ori_n1668_), .B(ori_ori_n1667_), .C(ori_ori_n588_), .Y(ori_ori_n1669_));
  AOI210     o1620(.A0(ori_ori_n1112_), .A1(ori_ori_n244_), .B0(ori_ori_n1454_), .Y(ori_ori_n1670_));
  AOI210     o1621(.A0(ori_ori_n1670_), .A1(ori_ori_n1669_), .B0(ori_ori_n769_), .Y(ori_ori_n1671_));
  NA4        o1622(.A(ori_ori_n589_), .B(ori_ori_n279_), .C(ori_ori_n164_), .D(ori_ori_n151_), .Y(ori_ori_n1672_));
  NA3        o1623(.A(ori_ori_n559_), .B(ori_ori_n267_), .C(ori_ori_n689_), .Y(ori_ori_n1673_));
  AOI210     o1624(.A0(ori_ori_n1673_), .A1(ori_ori_n1672_), .B0(ori_ori_n1020_), .Y(ori_ori_n1674_));
  OAI210     o1625(.A0(ori_ori_n776_), .A1(x8), .B0(x7), .Y(ori_ori_n1675_));
  NO2        o1626(.A(ori_ori_n1675_), .B(ori_ori_n117_), .Y(ori_ori_n1676_));
  OR2        o1627(.A(ori_ori_n750_), .B(ori_ori_n246_), .Y(ori_ori_n1677_));
  NO2        o1628(.A(ori_ori_n1677_), .B(ori_ori_n518_), .Y(ori_ori_n1678_));
  NO4        o1629(.A(ori_ori_n1678_), .B(ori_ori_n1676_), .C(ori_ori_n1674_), .D(ori_ori_n1671_), .Y(ori_ori_n1679_));
  OAI210     o1630(.A0(ori_ori_n1665_), .A1(x2), .B0(ori_ori_n1679_), .Y(ori_ori_n1680_));
  NO3        o1631(.A(x5), .B(ori_ori_n327_), .C(ori_ori_n130_), .Y(ori_ori_n1681_));
  AOI210     o1632(.A0(ori_ori_n625_), .A1(ori_ori_n542_), .B0(ori_ori_n1681_), .Y(ori_ori_n1682_));
  NA2        o1633(.A(x7), .B(ori_ori_n1682_), .Y(ori_ori_n1683_));
  NA3        o1634(.A(ori_ori_n1637_), .B(ori_ori_n211_), .C(ori_ori_n80_), .Y(ori_ori_n1684_));
  NA2        o1635(.A(ori_ori_n1684_), .B(x7), .Y(ori_ori_n1685_));
  AOI210     o1636(.A0(ori_ori_n1683_), .A1(x8), .B0(ori_ori_n1685_), .Y(ori_ori_n1686_));
  OAI210     o1637(.A0(ori_ori_n393_), .A1(ori_ori_n225_), .B0(ori_ori_n834_), .Y(ori_ori_n1687_));
  OAI210     o1638(.A0(ori_ori_n1687_), .A1(ori_ori_n955_), .B0(ori_ori_n595_), .Y(ori_ori_n1688_));
  NO3        o1639(.A(ori_ori_n882_), .B(ori_ori_n317_), .C(ori_ori_n136_), .Y(ori_ori_n1689_));
  NA3        o1640(.A(ori_ori_n1689_), .B(ori_ori_n1098_), .C(ori_ori_n50_), .Y(ori_ori_n1690_));
  NO2        o1641(.A(ori_ori_n123_), .B(ori_ori_n86_), .Y(ori_ori_n1691_));
  AOI220     o1642(.A0(ori_ori_n1691_), .A1(ori_ori_n519_), .B0(ori_ori_n1620_), .B1(ori_ori_n323_), .Y(ori_ori_n1692_));
  NOi31      o1643(.An(ori_ori_n956_), .B(ori_ori_n1575_), .C(ori_ori_n552_), .Y(ori_ori_n1693_));
  NA2        o1644(.A(ori_ori_n156_), .B(x4), .Y(ori_ori_n1694_));
  NO3        o1645(.A(ori_ori_n1251_), .B(ori_ori_n221_), .C(ori_ori_n68_), .Y(ori_ori_n1695_));
  AOI210     o1646(.A0(ori_ori_n1695_), .A1(ori_ori_n1694_), .B0(ori_ori_n1693_), .Y(ori_ori_n1696_));
  NA4        o1647(.A(ori_ori_n1696_), .B(ori_ori_n1692_), .C(ori_ori_n1690_), .D(ori_ori_n1688_), .Y(ori_ori_n1697_));
  NO4        o1648(.A(ori_ori_n1036_), .B(ori_ori_n154_), .C(ori_ori_n55_), .D(ori_ori_n68_), .Y(ori_ori_n1698_));
  NO4        o1649(.A(ori_ori_n1018_), .B(ori_ori_n441_), .C(x0), .D(ori_ori_n98_), .Y(ori_ori_n1699_));
  OAI210     o1650(.A0(ori_ori_n1699_), .A1(ori_ori_n1698_), .B0(ori_ori_n100_), .Y(ori_ori_n1700_));
  AOI210     o1651(.A0(ori_ori_n278_), .A1(x4), .B0(ori_ori_n173_), .Y(ori_ori_n1701_));
  NA2        o1652(.A(ori_ori_n1701_), .B(ori_ori_n620_), .Y(ori_ori_n1702_));
  OR3        o1653(.A(ori_ori_n1469_), .B(ori_ori_n1210_), .C(ori_ori_n924_), .Y(ori_ori_n1703_));
  NA2        o1654(.A(ori_ori_n1621_), .B(ori_ori_n696_), .Y(ori_ori_n1704_));
  OA220      o1655(.A0(ori_ori_n1704_), .A1(ori_ori_n225_), .B0(ori_ori_n511_), .B1(ori_ori_n1503_), .Y(ori_ori_n1705_));
  NA4        o1656(.A(ori_ori_n1705_), .B(ori_ori_n1703_), .C(ori_ori_n1702_), .D(ori_ori_n1700_), .Y(ori_ori_n1706_));
  AOI210     o1657(.A0(ori_ori_n1697_), .A1(ori_ori_n263_), .B0(ori_ori_n1706_), .Y(ori_ori_n1707_));
  OAI210     o1658(.A0(ori_ori_n1686_), .A1(x1), .B0(ori_ori_n1707_), .Y(ori_ori_n1708_));
  AO210      o1659(.A0(ori_ori_n1680_), .A1(x1), .B0(ori_ori_n1708_), .Y(ori30));
  NO3        o1660(.A(ori_ori_n1487_), .B(ori_ori_n507_), .C(ori_ori_n90_), .Y(ori_ori_n1710_));
  NO3        o1661(.A(ori_ori_n971_), .B(ori_ori_n126_), .C(ori_ori_n343_), .Y(ori_ori_n1711_));
  AOI210     o1662(.A0(ori_ori_n620_), .A1(ori_ori_n230_), .B0(ori_ori_n1711_), .Y(ori_ori_n1712_));
  AOI210     o1663(.A0(ori_ori_n1712_), .A1(ori_ori_n1710_), .B0(ori_ori_n56_), .Y(ori_ori_n1713_));
  NA2        o1664(.A(ori_ori_n701_), .B(ori_ori_n304_), .Y(ori_ori_n1714_));
  NA2        o1665(.A(ori_ori_n1714_), .B(ori_ori_n1147_), .Y(ori_ori_n1715_));
  OAI210     o1666(.A0(ori_ori_n1715_), .A1(ori_ori_n1713_), .B0(ori_ori_n100_), .Y(ori_ori_n1716_));
  OAI210     o1667(.A0(ori_ori_n865_), .A1(x1), .B0(ori_ori_n595_), .Y(ori_ori_n1717_));
  AOI220     o1668(.A0(ori_ori_n398_), .A1(ori_ori_n816_), .B0(x3), .B1(ori_ori_n405_), .Y(ori_ori_n1718_));
  AOI210     o1669(.A0(ori_ori_n1718_), .A1(ori_ori_n1717_), .B0(ori_ori_n233_), .Y(ori_ori_n1719_));
  NO3        o1670(.A(ori_ori_n252_), .B(ori_ori_n113_), .C(x0), .Y(ori_ori_n1720_));
  AOI210     o1671(.A0(ori_ori_n443_), .A1(x6), .B0(ori_ori_n1720_), .Y(ori_ori_n1721_));
  AOI220     o1672(.A0(ori_ori_n967_), .A1(ori_ori_n377_), .B0(x6), .B1(ori_ori_n85_), .Y(ori_ori_n1722_));
  OAI220     o1673(.A0(ori_ori_n1722_), .A1(ori_ori_n225_), .B0(ori_ori_n1721_), .B1(ori_ori_n54_), .Y(ori_ori_n1723_));
  AO210      o1674(.A0(ori_ori_n501_), .A1(ori_ori_n456_), .B0(x5), .Y(ori_ori_n1724_));
  NO2        o1675(.A(ori_ori_n617_), .B(ori_ori_n1724_), .Y(ori_ori_n1725_));
  AOI210     o1676(.A0(ori_ori_n1359_), .A1(ori_ori_n50_), .B0(ori_ori_n405_), .Y(ori_ori_n1726_));
  NA2        o1677(.A(ori_ori_n178_), .B(x2), .Y(ori_ori_n1727_));
  OA220      o1678(.A0(ori_ori_n1727_), .A1(ori_ori_n1726_), .B0(ori_ori_n247_), .B1(x6), .Y(ori_ori_n1728_));
  NO3        o1679(.A(ori_ori_n1150_), .B(ori_ori_n306_), .C(ori_ori_n883_), .Y(ori_ori_n1729_));
  NO2        o1680(.A(ori_ori_n455_), .B(ori_ori_n744_), .Y(ori_ori_n1730_));
  NOi21      o1681(.An(ori_ori_n1730_), .B(ori_ori_n730_), .Y(ori_ori_n1731_));
  NO2        o1682(.A(ori_ori_n1731_), .B(ori_ori_n1729_), .Y(ori_ori_n1732_));
  OAI210     o1683(.A0(ori_ori_n1728_), .A1(ori_ori_n653_), .B0(ori_ori_n1732_), .Y(ori_ori_n1733_));
  NO4        o1684(.A(ori_ori_n1733_), .B(ori_ori_n1725_), .C(ori_ori_n1723_), .D(ori_ori_n1719_), .Y(ori_ori_n1734_));
  AOI210     o1685(.A0(ori_ori_n1734_), .A1(ori_ori_n1716_), .B0(x8), .Y(ori_ori_n1735_));
  NO3        o1686(.A(ori_ori_n430_), .B(ori_ori_n676_), .C(ori_ori_n53_), .Y(ori_ori_n1736_));
  OAI220     o1687(.A0(ori_ori_n1503_), .A1(ori_ori_n306_), .B0(ori_ori_n422_), .B1(ori_ori_n515_), .Y(ori_ori_n1737_));
  OAI210     o1688(.A0(ori_ori_n1737_), .A1(ori_ori_n1736_), .B0(x6), .Y(ori_ori_n1738_));
  OAI210     o1689(.A0(ori_ori_n894_), .A1(ori_ori_n470_), .B0(ori_ori_n701_), .Y(ori_ori_n1739_));
  OAI210     o1690(.A0(ori_ori_n1460_), .A1(ori_ori_n296_), .B0(ori_ori_n116_), .Y(ori_ori_n1740_));
  AOI210     o1691(.A0(ori_ori_n340_), .A1(ori_ori_n210_), .B0(ori_ori_n69_), .Y(ori_ori_n1741_));
  AOI210     o1692(.A0(ori_ori_n865_), .A1(ori_ori_n644_), .B0(ori_ori_n1741_), .Y(ori_ori_n1742_));
  NA4        o1693(.A(ori_ori_n1742_), .B(ori_ori_n1740_), .C(ori_ori_n1739_), .D(ori_ori_n1738_), .Y(ori_ori_n1743_));
  NA2        o1694(.A(ori_ori_n929_), .B(ori_ori_n57_), .Y(ori_ori_n1744_));
  AOI210     o1695(.A0(ori_ori_n801_), .A1(ori_ori_n431_), .B0(ori_ori_n600_), .Y(ori_ori_n1745_));
  OAI220     o1696(.A0(ori_ori_n1745_), .A1(ori_ori_n278_), .B0(ori_ori_n1744_), .B1(ori_ori_n421_), .Y(ori_ori_n1746_));
  AOI210     o1697(.A0(ori_ori_n1743_), .A1(x8), .B0(ori_ori_n1746_), .Y(ori_ori_n1747_));
  INV        o1698(.A(ori_ori_n1747_), .Y(ori_ori_n1748_));
  INV        o1699(.A(ori_ori_n800_), .Y(ori_ori_n1749_));
  NO2        o1700(.A(ori_ori_n1749_), .B(ori_ori_n395_), .Y(ori_ori_n1750_));
  NO2        o1701(.A(ori_ori_n565_), .B(ori_ori_n366_), .Y(ori_ori_n1751_));
  NO3        o1702(.A(ori_ori_n1751_), .B(ori_ori_n1063_), .C(x0), .Y(ori_ori_n1752_));
  AOI210     o1703(.A0(ori_ori_n275_), .A1(x1), .B0(ori_ori_n136_), .Y(ori_ori_n1753_));
  NO2        o1704(.A(ori_ori_n2184_), .B(ori_ori_n738_), .Y(ori_ori_n1754_));
  OAI220     o1705(.A0(ori_ori_n1754_), .A1(ori_ori_n901_), .B0(ori_ori_n1753_), .B1(ori_ori_n188_), .Y(ori_ori_n1755_));
  NO3        o1706(.A(ori_ori_n1755_), .B(ori_ori_n1752_), .C(ori_ori_n1750_), .Y(ori_ori_n1756_));
  NO2        o1707(.A(ori_ori_n275_), .B(ori_ori_n112_), .Y(ori_ori_n1757_));
  NA2        o1708(.A(ori_ori_n1757_), .B(ori_ori_n142_), .Y(ori_ori_n1758_));
  NA2        o1709(.A(ori_ori_n1119_), .B(x2), .Y(ori_ori_n1759_));
  AOI210     o1710(.A0(ori_ori_n1759_), .A1(ori_ori_n1758_), .B0(ori_ori_n50_), .Y(ori_ori_n1760_));
  NA3        o1711(.A(ori_ori_n2175_), .B(ori_ori_n2182_), .C(ori_ori_n414_), .Y(ori_ori_n1761_));
  NO2        o1712(.A(ori_ori_n1761_), .B(ori_ori_n538_), .Y(ori_ori_n1762_));
  AOI210     o1713(.A0(ori_ori_n883_), .A1(x1), .B0(ori_ori_n1112_), .Y(ori_ori_n1763_));
  NA2        o1714(.A(ori_ori_n990_), .B(ori_ori_n552_), .Y(ori_ori_n1764_));
  OAI210     o1715(.A0(ori_ori_n1763_), .A1(ori_ori_n425_), .B0(ori_ori_n1764_), .Y(ori_ori_n1765_));
  NO3        o1716(.A(ori_ori_n1765_), .B(ori_ori_n1762_), .C(ori_ori_n1760_), .Y(ori_ori_n1766_));
  OAI210     o1717(.A0(ori_ori_n1756_), .A1(ori_ori_n123_), .B0(ori_ori_n1766_), .Y(ori_ori_n1767_));
  NO3        o1718(.A(ori_ori_n1767_), .B(ori_ori_n1748_), .C(ori_ori_n1735_), .Y(ori31));
  NO2        o1719(.A(ori_ori_n677_), .B(ori_ori_n56_), .Y(ori_ori_n1769_));
  AOI220     o1720(.A0(ori_ori_n1769_), .A1(x2), .B0(ori_ori_n84_), .B1(x0), .Y(ori_ori_n1770_));
  NA3        o1721(.A(ori_ori_n1770_), .B(ori_ori_n1704_), .C(ori_ori_n1554_), .Y(ori_ori_n1771_));
  NA2        o1722(.A(ori_ori_n1771_), .B(ori_ori_n53_), .Y(ori_ori_n1772_));
  INV        o1723(.A(ori_ori_n595_), .Y(ori_ori_n1773_));
  NO3        o1724(.A(ori_ori_n1645_), .B(ori_ori_n1621_), .C(ori_ori_n770_), .Y(ori_ori_n1774_));
  OA220      o1725(.A0(ori_ori_n1774_), .A1(ori_ori_n414_), .B0(ori_ori_n1773_), .B1(x7), .Y(ori_ori_n1775_));
  AOI210     o1726(.A0(ori_ori_n1775_), .A1(ori_ori_n1772_), .B0(ori_ori_n98_), .Y(ori_ori_n1776_));
  NO2        o1727(.A(ori_ori_n437_), .B(ori_ori_n72_), .Y(ori_ori_n1777_));
  NA2        o1728(.A(ori_ori_n1777_), .B(ori_ori_n664_), .Y(ori_ori_n1778_));
  NO4        o1729(.A(ori_ori_n987_), .B(ori_ori_n327_), .C(ori_ori_n1359_), .D(ori_ori_n64_), .Y(ori_ori_n1779_));
  AOI210     o1730(.A0(ori_ori_n1386_), .A1(ori_ori_n1142_), .B0(ori_ori_n393_), .Y(ori_ori_n1780_));
  OAI220     o1731(.A0(ori_ori_n1104_), .A1(ori_ori_n825_), .B0(x2), .B1(ori_ori_n106_), .Y(ori_ori_n1781_));
  NO3        o1732(.A(ori_ori_n1781_), .B(ori_ori_n1780_), .C(ori_ori_n1779_), .Y(ori_ori_n1782_));
  AOI210     o1733(.A0(ori_ori_n1782_), .A1(ori_ori_n1778_), .B0(x5), .Y(ori_ori_n1783_));
  AOI220     o1734(.A0(ori_ori_n397_), .A1(ori_ori_n552_), .B0(x1), .B1(ori_ori_n61_), .Y(ori_ori_n1784_));
  AOI210     o1735(.A0(ori_ori_n1784_), .A1(ori_ori_n511_), .B0(ori_ori_n1036_), .Y(ori_ori_n1785_));
  NA2        o1736(.A(ori_ori_n833_), .B(ori_ori_n631_), .Y(ori_ori_n1786_));
  OAI220     o1737(.A0(ori_ori_n1786_), .A1(ori_ori_n345_), .B0(ori_ori_n421_), .B1(ori_ori_n665_), .Y(ori_ori_n1787_));
  NO4        o1738(.A(ori_ori_n1787_), .B(ori_ori_n1785_), .C(ori_ori_n1783_), .D(ori_ori_n1776_), .Y(ori_ori_n1788_));
  NA2        o1739(.A(ori_ori_n431_), .B(ori_ori_n57_), .Y(ori_ori_n1789_));
  AOI210     o1740(.A0(ori_ori_n475_), .A1(ori_ori_n1789_), .B0(ori_ori_n129_), .Y(ori_ori_n1790_));
  OAI210     o1741(.A0(ori_ori_n94_), .A1(ori_ori_n246_), .B0(ori_ori_n1744_), .Y(ori_ori_n1791_));
  OAI210     o1742(.A0(ori_ori_n1791_), .A1(ori_ori_n1790_), .B0(x7), .Y(ori_ori_n1792_));
  OA210      o1743(.A0(ori_ori_n2169_), .A1(ori_ori_n1111_), .B0(ori_ori_n92_), .Y(ori_ori_n1793_));
  NO2        o1744(.A(ori_ori_n782_), .B(ori_ori_n57_), .Y(ori_ori_n1794_));
  NA2        o1745(.A(ori_ori_n1312_), .B(x6), .Y(ori_ori_n1795_));
  AOI210     o1746(.A0(ori_ori_n1795_), .A1(ori_ori_n262_), .B0(ori_ori_n98_), .Y(ori_ori_n1796_));
  NO3        o1747(.A(ori_ori_n1796_), .B(ori_ori_n1794_), .C(ori_ori_n1793_), .Y(ori_ori_n1797_));
  AOI210     o1748(.A0(ori_ori_n1797_), .A1(ori_ori_n1792_), .B0(ori_ori_n604_), .Y(ori_ori_n1798_));
  NOi21      o1749(.An(ori_ori_n1478_), .B(ori_ori_n904_), .Y(ori_ori_n1799_));
  OAI220     o1750(.A0(ori_ori_n1799_), .A1(ori_ori_n1623_), .B0(ori_ori_n802_), .B1(ori_ori_n1789_), .Y(ori_ori_n1800_));
  NA2        o1751(.A(ori_ori_n1800_), .B(x3), .Y(ori_ori_n1801_));
  AOI220     o1752(.A0(ori_ori_n1171_), .A1(x8), .B0(ori_ori_n58_), .B1(x1), .Y(ori_ori_n1802_));
  NO3        o1753(.A(ori_ori_n1802_), .B(ori_ori_n948_), .C(x6), .Y(ori_ori_n1803_));
  AOI220     o1754(.A0(ori_ori_n542_), .A1(ori_ori_n366_), .B0(ori_ori_n431_), .B1(ori_ori_n75_), .Y(ori_ori_n1804_));
  NA2        o1755(.A(ori_ori_n107_), .B(ori_ori_n462_), .Y(ori_ori_n1805_));
  OAI220     o1756(.A0(ori_ori_n1805_), .A1(ori_ori_n1623_), .B0(ori_ori_n1804_), .B1(x4), .Y(ori_ori_n1806_));
  NO2        o1757(.A(ori_ori_n1806_), .B(ori_ori_n1803_), .Y(ori_ori_n1807_));
  AOI210     o1758(.A0(ori_ori_n1807_), .A1(ori_ori_n1801_), .B0(ori_ori_n166_), .Y(ori_ori_n1808_));
  NO4        o1759(.A(ori_ori_n543_), .B(ori_ori_n519_), .C(ori_ori_n611_), .D(ori_ori_n610_), .Y(ori_ori_n1809_));
  OAI210     o1760(.A0(ori_ori_n1809_), .A1(ori_ori_n917_), .B0(x3), .Y(ori_ori_n1810_));
  NO4        o1761(.A(ori_ori_n692_), .B(ori_ori_n1036_), .C(ori_ori_n664_), .D(x5), .Y(ori_ori_n1811_));
  NO3        o1762(.A(x6), .B(ori_ori_n56_), .C(x1), .Y(ori_ori_n1812_));
  NA2        o1763(.A(ori_ori_n1812_), .B(ori_ori_n258_), .Y(ori_ori_n1813_));
  OAI210     o1764(.A0(ori_ori_n1596_), .A1(ori_ori_n340_), .B0(ori_ori_n1813_), .Y(ori_ori_n1814_));
  NA4        o1765(.A(ori_ori_n565_), .B(ori_ori_n160_), .C(x6), .D(ori_ori_n98_), .Y(ori_ori_n1815_));
  NO2        o1766(.A(ori_ori_n739_), .B(ori_ori_n228_), .Y(ori_ori_n1816_));
  NOi41      o1767(.An(ori_ori_n1815_), .B(ori_ori_n1816_), .C(ori_ori_n1814_), .D(ori_ori_n1811_), .Y(ori_ori_n1817_));
  AOI210     o1768(.A0(ori_ori_n1817_), .A1(ori_ori_n1810_), .B0(ori_ori_n466_), .Y(ori_ori_n1818_));
  NO3        o1769(.A(ori_ori_n337_), .B(ori_ori_n74_), .C(ori_ori_n53_), .Y(ori_ori_n1819_));
  NA2        o1770(.A(ori_ori_n1819_), .B(ori_ori_n988_), .Y(ori_ori_n1820_));
  NO2        o1771(.A(ori_ori_n1820_), .B(ori_ori_n352_), .Y(ori_ori_n1821_));
  AOI220     o1772(.A0(ori_ori_n1341_), .A1(ori_ori_n788_), .B0(ori_ori_n245_), .B1(x4), .Y(ori_ori_n1822_));
  NO2        o1773(.A(ori_ori_n1822_), .B(ori_ori_n171_), .Y(ori_ori_n1823_));
  OR2        o1774(.A(ori_ori_n1823_), .B(ori_ori_n1821_), .Y(ori_ori_n1824_));
  NO4        o1775(.A(ori_ori_n1824_), .B(ori_ori_n1818_), .C(ori_ori_n1808_), .D(ori_ori_n1798_), .Y(ori_ori_n1825_));
  OAI210     o1776(.A0(ori_ori_n1788_), .A1(x3), .B0(ori_ori_n1825_), .Y(ori32));
  OAI210     o1777(.A0(ori_ori_n495_), .A1(ori_ori_n53_), .B0(ori_ori_n369_), .Y(ori_ori_n1827_));
  NA2        o1778(.A(ori_ori_n452_), .B(x2), .Y(ori_ori_n1828_));
  NA2        o1779(.A(ori_ori_n1828_), .B(ori_ori_n1827_), .Y(ori_ori_n1829_));
  OAI210     o1780(.A0(ori_ori_n1829_), .A1(ori_ori_n678_), .B0(ori_ori_n56_), .Y(ori_ori_n1830_));
  OAI210     o1781(.A0(ori_ori_n1445_), .A1(ori_ori_n1226_), .B0(ori_ori_n1250_), .Y(ori_ori_n1831_));
  AOI210     o1782(.A0(ori_ori_n1769_), .A1(ori_ori_n249_), .B0(ori_ori_n1831_), .Y(ori_ori_n1832_));
  AOI210     o1783(.A0(ori_ori_n1832_), .A1(ori_ori_n1830_), .B0(ori_ori_n50_), .Y(ori_ori_n1833_));
  NA3        o1784(.A(ori_ori_n55_), .B(ori_ori_n690_), .C(ori_ori_n261_), .Y(ori_ori_n1834_));
  NA2        o1785(.A(ori_ori_n642_), .B(ori_ori_n478_), .Y(ori_ori_n1835_));
  OAI220     o1786(.A0(ori_ori_n900_), .A1(ori_ori_n211_), .B0(ori_ori_n601_), .B1(ori_ori_n188_), .Y(ori_ori_n1836_));
  NO2        o1787(.A(ori_ori_n338_), .B(ori_ori_n504_), .Y(ori_ori_n1837_));
  NO3        o1788(.A(ori_ori_n1150_), .B(ori_ori_n515_), .C(ori_ori_n244_), .Y(ori_ori_n1838_));
  NO4        o1789(.A(ori_ori_n1838_), .B(ori_ori_n1837_), .C(ori_ori_n1836_), .D(ori_ori_n1835_), .Y(ori_ori_n1839_));
  AOI210     o1790(.A0(ori_ori_n1839_), .A1(ori_ori_n1834_), .B0(ori_ori_n130_), .Y(ori_ori_n1840_));
  OAI220     o1791(.A0(ori_ori_n361_), .A1(x7), .B0(ori_ori_n274_), .B1(ori_ori_n267_), .Y(ori_ori_n1841_));
  NA2        o1792(.A(ori_ori_n1841_), .B(ori_ori_n832_), .Y(ori_ori_n1842_));
  NO2        o1793(.A(ori_ori_n482_), .B(ori_ori_n744_), .Y(ori_ori_n1843_));
  AOI220     o1794(.A0(ori_ori_n1843_), .A1(ori_ori_n1578_), .B0(ori_ori_n463_), .B1(x8), .Y(ori_ori_n1844_));
  AOI210     o1795(.A0(ori_ori_n1844_), .A1(ori_ori_n1842_), .B0(ori_ori_n100_), .Y(ori_ori_n1845_));
  NA3        o1796(.A(ori_ori_n1111_), .B(ori_ori_n973_), .C(ori_ori_n106_), .Y(ori_ori_n1846_));
  INV        o1797(.A(ori_ori_n1050_), .Y(ori_ori_n1847_));
  AOI210     o1798(.A0(ori_ori_n1847_), .A1(ori_ori_n1846_), .B0(ori_ori_n56_), .Y(ori_ori_n1848_));
  NA2        o1799(.A(ori_ori_n879_), .B(ori_ori_n228_), .Y(ori_ori_n1849_));
  NO3        o1800(.A(ori_ori_n1849_), .B(ori_ori_n55_), .C(ori_ori_n57_), .Y(ori_ori_n1850_));
  OR4        o1801(.A(ori_ori_n1850_), .B(ori_ori_n1848_), .C(ori_ori_n1845_), .D(ori_ori_n1840_), .Y(ori_ori_n1851_));
  OAI210     o1802(.A0(ori_ori_n1851_), .A1(ori_ori_n1833_), .B0(ori_ori_n98_), .Y(ori_ori_n1852_));
  NO3        o1803(.A(ori_ori_n1036_), .B(ori_ori_n133_), .C(ori_ori_n114_), .Y(ori_ori_n1853_));
  NO2        o1804(.A(ori_ori_n341_), .B(ori_ori_n55_), .Y(ori_ori_n1854_));
  NA2        o1805(.A(ori_ori_n1854_), .B(ori_ori_n105_), .Y(ori_ori_n1855_));
  OAI210     o1806(.A0(ori_ori_n561_), .A1(ori_ori_n521_), .B0(ori_ori_n701_), .Y(ori_ori_n1856_));
  NA2        o1807(.A(ori_ori_n1856_), .B(ori_ori_n1855_), .Y(ori_ori_n1857_));
  OAI210     o1808(.A0(ori_ori_n1857_), .A1(ori_ori_n1853_), .B0(x3), .Y(ori_ori_n1858_));
  OAI210     o1809(.A0(ori_ori_n776_), .A1(ori_ori_n244_), .B0(ori_ori_n50_), .Y(ori_ori_n1859_));
  AOI210     o1810(.A0(ori_ori_n60_), .A1(ori_ori_n100_), .B0(ori_ori_n1859_), .Y(ori_ori_n1860_));
  OAI210     o1811(.A0(ori_ori_n1860_), .A1(ori_ori_n1560_), .B0(ori_ori_n610_), .Y(ori_ori_n1861_));
  NO3        o1812(.A(ori_ori_n276_), .B(ori_ori_n156_), .C(ori_ori_n112_), .Y(ori_ori_n1862_));
  NO3        o1813(.A(ori_ori_n690_), .B(ori_ori_n325_), .C(ori_ori_n130_), .Y(ori_ori_n1863_));
  OAI210     o1814(.A0(ori_ori_n1863_), .A1(ori_ori_n1862_), .B0(ori_ori_n57_), .Y(ori_ori_n1864_));
  NA2        o1815(.A(ori_ori_n976_), .B(ori_ori_n68_), .Y(ori_ori_n1865_));
  AOI210     o1816(.A0(ori_ori_n2183_), .A1(ori_ori_n1561_), .B0(ori_ori_n1865_), .Y(ori_ori_n1866_));
  INV        o1817(.A(ori_ori_n246_), .Y(ori_ori_n1867_));
  NOi31      o1818(.An(ori_ori_n620_), .B(ori_ori_n246_), .C(ori_ori_n252_), .Y(ori_ori_n1868_));
  NO3        o1819(.A(ori_ori_n1868_), .B(ori_ori_n1866_), .C(x1), .Y(ori_ori_n1869_));
  NA4        o1820(.A(ori_ori_n1869_), .B(ori_ori_n1864_), .C(ori_ori_n1861_), .D(ori_ori_n1858_), .Y(ori_ori_n1870_));
  AO210      o1821(.A0(ori_ori_n932_), .A1(ori_ori_n356_), .B0(ori_ori_n875_), .Y(ori_ori_n1871_));
  NA3        o1822(.A(ori_ori_n1602_), .B(ori_ori_n486_), .C(ori_ori_n246_), .Y(ori_ori_n1872_));
  AOI210     o1823(.A0(ori_ori_n1872_), .A1(ori_ori_n1871_), .B0(ori_ori_n276_), .Y(ori_ori_n1873_));
  NO3        o1824(.A(ori_ori_n1210_), .B(ori_ori_n875_), .C(x2), .Y(ori_ori_n1874_));
  NO2        o1825(.A(ori_ori_n1058_), .B(ori_ori_n344_), .Y(ori_ori_n1875_));
  NO3        o1826(.A(ori_ori_n1875_), .B(ori_ori_n1874_), .C(ori_ori_n53_), .Y(ori_ori_n1876_));
  OAI220     o1827(.A0(ori_ori_n604_), .A1(ori_ori_n156_), .B0(ori_ori_n317_), .B1(ori_ori_n130_), .Y(ori_ori_n1877_));
  NA2        o1828(.A(ori_ori_n1877_), .B(ori_ori_n65_), .Y(ori_ori_n1878_));
  NO2        o1829(.A(ori_ori_n1666_), .B(ori_ori_n329_), .Y(ori_ori_n1879_));
  NA2        o1830(.A(ori_ori_n1565_), .B(ori_ori_n1879_), .Y(ori_ori_n1880_));
  NA3        o1831(.A(ori_ori_n1880_), .B(ori_ori_n1878_), .C(ori_ori_n1876_), .Y(ori_ori_n1881_));
  OAI210     o1832(.A0(ori_ori_n1881_), .A1(ori_ori_n1873_), .B0(ori_ori_n1870_), .Y(ori_ori_n1882_));
  NO3        o1833(.A(ori_ori_n1023_), .B(ori_ori_n97_), .C(ori_ori_n68_), .Y(ori_ori_n1883_));
  NO2        o1834(.A(ori_ori_n495_), .B(ori_ori_n333_), .Y(ori_ori_n1884_));
  OAI210     o1835(.A0(ori_ori_n1883_), .A1(ori_ori_n1190_), .B0(ori_ori_n1884_), .Y(ori_ori_n1885_));
  NO3        o1836(.A(x8), .B(ori_ori_n68_), .C(x2), .Y(ori_ori_n1886_));
  OAI220     o1837(.A0(ori_ori_n1886_), .A1(ori_ori_n552_), .B0(ori_ori_n1200_), .B1(ori_ori_n84_), .Y(ori_ori_n1887_));
  AOI220     o1838(.A0(ori_ori_n487_), .A1(ori_ori_n701_), .B0(ori_ori_n595_), .B1(ori_ori_n231_), .Y(ori_ori_n1888_));
  AOI210     o1839(.A0(ori_ori_n1888_), .A1(ori_ori_n1887_), .B0(ori_ori_n238_), .Y(ori_ori_n1889_));
  NO2        o1840(.A(ori_ori_n400_), .B(ori_ori_n383_), .Y(ori_ori_n1890_));
  NOi31      o1841(.An(ori_ori_n1265_), .B(ori_ori_n1890_), .C(ori_ori_n519_), .Y(ori_ori_n1891_));
  NO2        o1842(.A(ori_ori_n1891_), .B(ori_ori_n1889_), .Y(ori_ori_n1892_));
  NA4        o1843(.A(ori_ori_n1892_), .B(ori_ori_n1885_), .C(ori_ori_n1882_), .D(ori_ori_n1852_), .Y(ori33));
  OAI210     o1844(.A0(ori_ori_n2184_), .A1(ori_ori_n159_), .B0(ori_ori_n294_), .Y(ori_ori_n1894_));
  OAI210     o1845(.A0(ori_ori_n912_), .A1(ori_ori_n696_), .B0(ori_ori_n316_), .Y(ori_ori_n1895_));
  NA3        o1846(.A(ori_ori_n1895_), .B(ori_ori_n1894_), .C(ori_ori_n564_), .Y(ori_ori_n1896_));
  AOI210     o1847(.A0(ori_ori_n100_), .A1(x5), .B0(ori_ori_n1896_), .Y(ori_ori_n1897_));
  NA2        o1848(.A(ori_ori_n210_), .B(ori_ori_n73_), .Y(ori_ori_n1898_));
  NA4        o1849(.A(ori_ori_n1466_), .B(ori_ori_n496_), .C(ori_ori_n225_), .D(x4), .Y(ori_ori_n1899_));
  AOI210     o1850(.A0(ori_ori_n1899_), .A1(ori_ori_n1898_), .B0(ori_ori_n316_), .Y(ori_ori_n1900_));
  NA2        o1851(.A(ori_ori_n1398_), .B(ori_ori_n68_), .Y(ori_ori_n1901_));
  NO2        o1852(.A(ori_ori_n1901_), .B(ori_ori_n1900_), .Y(ori_ori_n1902_));
  OAI210     o1853(.A0(ori_ori_n1897_), .A1(x4), .B0(ori_ori_n1902_), .Y(ori_ori_n1903_));
  OAI210     o1854(.A0(ori_ori_n132_), .A1(x5), .B0(ori_ori_n220_), .Y(ori_ori_n1904_));
  NA2        o1855(.A(ori_ori_n166_), .B(x4), .Y(ori_ori_n1905_));
  NA2        o1856(.A(ori_ori_n280_), .B(ori_ori_n258_), .Y(ori_ori_n1906_));
  NO2        o1857(.A(ori_ori_n832_), .B(ori_ori_n208_), .Y(ori_ori_n1907_));
  NA2        o1858(.A(ori_ori_n567_), .B(x7), .Y(ori_ori_n1908_));
  OAI220     o1859(.A0(ori_ori_n1908_), .A1(ori_ori_n1907_), .B0(ori_ori_n1906_), .B1(ori_ori_n1905_), .Y(ori_ori_n1909_));
  AOI210     o1860(.A0(ori_ori_n1904_), .A1(ori_ori_n882_), .B0(ori_ori_n1909_), .Y(ori_ori_n1910_));
  NA2        o1861(.A(x4), .B(ori_ori_n824_), .Y(ori_ori_n1911_));
  NO2        o1862(.A(ori_ori_n1911_), .B(ori_ori_n194_), .Y(ori_ori_n1912_));
  OAI210     o1863(.A0(ori_ori_n744_), .A1(ori_ori_n51_), .B0(x6), .Y(ori_ori_n1913_));
  NA3        o1864(.A(ori_ori_n796_), .B(ori_ori_n626_), .C(ori_ori_n55_), .Y(ori_ori_n1914_));
  OAI210     o1865(.A0(ori_ori_n546_), .A1(ori_ori_n443_), .B0(ori_ori_n1914_), .Y(ori_ori_n1915_));
  NO3        o1866(.A(ori_ori_n1915_), .B(ori_ori_n1913_), .C(ori_ori_n1912_), .Y(ori_ori_n1916_));
  OAI210     o1867(.A0(ori_ori_n1910_), .A1(ori_ori_n50_), .B0(ori_ori_n1916_), .Y(ori_ori_n1917_));
  NA3        o1868(.A(ori_ori_n1917_), .B(ori_ori_n1903_), .C(ori_ori_n57_), .Y(ori_ori_n1918_));
  NO2        o1869(.A(ori_ori_n130_), .B(ori_ori_n301_), .Y(ori_ori_n1919_));
  NAi21      o1870(.An(ori_ori_n1011_), .B(ori_ori_n427_), .Y(ori_ori_n1920_));
  NA4        o1871(.A(ori_ori_n567_), .B(ori_ori_n1098_), .C(ori_ori_n412_), .D(ori_ori_n50_), .Y(ori_ori_n1921_));
  OAI210     o1872(.A0(ori_ori_n1919_), .A1(ori_ori_n1730_), .B0(x2), .Y(ori_ori_n1922_));
  NA4        o1873(.A(ori_ori_n258_), .B(ori_ori_n143_), .C(ori_ori_n247_), .D(ori_ori_n111_), .Y(ori_ori_n1923_));
  NA3        o1874(.A(ori_ori_n1923_), .B(ori_ori_n1922_), .C(ori_ori_n1921_), .Y(ori_ori_n1924_));
  AO220      o1875(.A0(ori_ori_n1924_), .A1(x0), .B0(ori_ori_n1920_), .B1(ori_ori_n127_), .Y(ori_ori_n1925_));
  NA3        o1876(.A(ori_ori_n664_), .B(ori_ori_n316_), .C(ori_ori_n58_), .Y(ori_ori_n1926_));
  NO2        o1877(.A(ori_ori_n1886_), .B(ori_ori_n368_), .Y(ori_ori_n1927_));
  NA2        o1878(.A(ori_ori_n565_), .B(ori_ori_n455_), .Y(ori_ori_n1928_));
  OAI220     o1879(.A0(ori_ori_n1928_), .A1(ori_ori_n1927_), .B0(ori_ori_n1926_), .B1(ori_ori_n68_), .Y(ori_ori_n1929_));
  OAI210     o1880(.A0(ori_ori_n1289_), .A1(ori_ori_n312_), .B0(ori_ori_n101_), .Y(ori_ori_n1930_));
  AOI210     o1881(.A0(ori_ori_n519_), .A1(ori_ori_n410_), .B0(ori_ori_n127_), .Y(ori_ori_n1931_));
  OAI210     o1882(.A0(ori_ori_n1931_), .A1(ori_ori_n345_), .B0(ori_ori_n1930_), .Y(ori_ori_n1932_));
  OAI210     o1883(.A0(ori_ori_n1932_), .A1(ori_ori_n1929_), .B0(ori_ori_n93_), .Y(ori_ori_n1933_));
  NA3        o1884(.A(ori_ori_n1019_), .B(ori_ori_n121_), .C(ori_ori_n341_), .Y(ori_ori_n1934_));
  NA2        o1885(.A(ori_ori_n1934_), .B(ori_ori_n1528_), .Y(ori_ori_n1935_));
  NA2        o1886(.A(ori_ori_n1009_), .B(ori_ori_n614_), .Y(ori_ori_n1936_));
  NA3        o1887(.A(ori_ori_n1936_), .B(ori_ori_n1935_), .C(ori_ori_n1933_), .Y(ori_ori_n1937_));
  AOI210     o1888(.A0(ori_ori_n1925_), .A1(x7), .B0(ori_ori_n1937_), .Y(ori_ori_n1938_));
  NA2        o1889(.A(ori_ori_n1938_), .B(ori_ori_n1918_), .Y(ori34));
  NA2        o1890(.A(ori_ori_n383_), .B(x4), .Y(ori_ori_n1940_));
  NO2        o1891(.A(ori_ori_n1645_), .B(ori_ori_n738_), .Y(ori_ori_n1941_));
  AOI210     o1892(.A0(ori_ori_n1941_), .A1(ori_ori_n1940_), .B0(ori_ori_n288_), .Y(ori_ori_n1942_));
  NA2        o1893(.A(ori_ori_n258_), .B(ori_ori_n112_), .Y(ori_ori_n1943_));
  NO2        o1894(.A(ori_ori_n842_), .B(ori_ori_n1943_), .Y(ori_ori_n1944_));
  AOI210     o1895(.A0(ori_ori_n1714_), .A1(ori_ori_n475_), .B0(ori_ori_n129_), .Y(ori_ori_n1945_));
  NA2        o1896(.A(ori_ori_n1645_), .B(x0), .Y(ori_ori_n1946_));
  OAI210     o1897(.A0(ori_ori_n1535_), .A1(ori_ori_n846_), .B0(ori_ori_n1946_), .Y(ori_ori_n1947_));
  NO4        o1898(.A(ori_ori_n1947_), .B(ori_ori_n1945_), .C(ori_ori_n1944_), .D(ori_ori_n1942_), .Y(ori_ori_n1948_));
  NO2        o1899(.A(ori_ori_n1948_), .B(ori_ori_n414_), .Y(ori_ori_n1949_));
  NA2        o1900(.A(ori_ori_n629_), .B(x8), .Y(ori_ori_n1950_));
  OAI210     o1901(.A0(ori_ori_n111_), .A1(ori_ori_n897_), .B0(x5), .Y(ori_ori_n1951_));
  INV        o1902(.A(ori_ori_n1951_), .Y(ori_ori_n1952_));
  NA3        o1903(.A(ori_ori_n1952_), .B(ori_ori_n302_), .C(x8), .Y(ori_ori_n1953_));
  NA2        o1904(.A(ori_ori_n1344_), .B(x3), .Y(ori_ori_n1954_));
  NA3        o1905(.A(ori_ori_n2165_), .B(ori_ori_n1954_), .C(ori_ori_n1953_), .Y(ori_ori_n1955_));
  NA2        o1906(.A(ori_ori_n941_), .B(ori_ori_n644_), .Y(ori_ori_n1956_));
  NA3        o1907(.A(ori_ori_n973_), .B(ori_ori_n151_), .C(ori_ori_n929_), .Y(ori_ori_n1957_));
  AOI210     o1908(.A0(ori_ori_n1957_), .A1(ori_ori_n1956_), .B0(ori_ori_n654_), .Y(ori_ori_n1958_));
  AOI210     o1909(.A0(ori_ori_n1487_), .A1(x8), .B0(ori_ori_n1958_), .Y(ori_ori_n1959_));
  NO2        o1910(.A(ori_ori_n487_), .B(ori_ori_n230_), .Y(ori_ori_n1960_));
  OAI220     o1911(.A0(ori_ori_n1960_), .A1(ori_ori_n57_), .B0(x7), .B1(ori_ori_n55_), .Y(ori_ori_n1961_));
  NA3        o1912(.A(ori_ori_n1961_), .B(ori_ori_n629_), .C(ori_ori_n56_), .Y(ori_ori_n1962_));
  OAI210     o1913(.A0(ori_ori_n1959_), .A1(ori_ori_n130_), .B0(ori_ori_n1962_), .Y(ori_ori_n1963_));
  NO3        o1914(.A(ori_ori_n1963_), .B(ori_ori_n1955_), .C(ori_ori_n1949_), .Y(ori_ori_n1964_));
  NO2        o1915(.A(ori_ori_n2186_), .B(ori_ori_n824_), .Y(ori_ori_n1965_));
  NO3        o1916(.A(ori_ori_n1965_), .B(ori_ori_n393_), .C(x3), .Y(ori_ori_n1966_));
  NA2        o1917(.A(ori_ori_n673_), .B(ori_ori_n146_), .Y(ori_ori_n1967_));
  NO3        o1918(.A(ori_ori_n1867_), .B(ori_ori_n275_), .C(ori_ori_n929_), .Y(ori_ori_n1968_));
  OAI220     o1919(.A0(ori_ori_n1968_), .A1(ori_ori_n1316_), .B0(ori_ori_n1967_), .B1(ori_ori_n994_), .Y(ori_ori_n1969_));
  OAI210     o1920(.A0(ori_ori_n1969_), .A1(ori_ori_n1966_), .B0(x2), .Y(ori_ori_n1970_));
  OAI210     o1921(.A0(ori_ori_n747_), .A1(ori_ori_n333_), .B0(ori_ori_n1970_), .Y(ori_ori_n1971_));
  NA2        o1922(.A(ori_ori_n283_), .B(x4), .Y(ori_ori_n1972_));
  OAI220     o1923(.A0(ori_ori_n641_), .A1(ori_ori_n55_), .B0(ori_ori_n251_), .B1(ori_ori_n97_), .Y(ori_ori_n1973_));
  NO2        o1924(.A(ori_ori_n941_), .B(ori_ori_n259_), .Y(ori_ori_n1974_));
  NO3        o1925(.A(ori_ori_n1974_), .B(ori_ori_n1973_), .C(ori_ori_n1972_), .Y(ori_ori_n1975_));
  NA3        o1926(.A(ori_ori_n1175_), .B(ori_ori_n233_), .C(x7), .Y(ori_ori_n1976_));
  INV        o1927(.A(ori_ori_n1976_), .Y(ori_ori_n1977_));
  OAI210     o1928(.A0(ori_ori_n1977_), .A1(ori_ori_n1975_), .B0(ori_ori_n149_), .Y(ori_ori_n1978_));
  NA3        o1929(.A(ori_ori_n742_), .B(ori_ori_n83_), .C(x0), .Y(ori_ori_n1979_));
  NA4        o1930(.A(ori_ori_n1979_), .B(ori_ori_n976_), .C(ori_ori_n268_), .D(ori_ori_n517_), .Y(ori_ori_n1980_));
  NA2        o1931(.A(ori_ori_n980_), .B(ori_ori_n595_), .Y(ori_ori_n1981_));
  OAI210     o1932(.A0(ori_ori_n1981_), .A1(ori_ori_n239_), .B0(ori_ori_n1815_), .Y(ori_ori_n1982_));
  NA2        o1933(.A(ori_ori_n1982_), .B(x7), .Y(ori_ori_n1983_));
  INV        o1934(.A(ori_ori_n633_), .Y(ori_ori_n1984_));
  AOI210     o1935(.A0(ori_ori_n242_), .A1(ori_ori_n53_), .B0(ori_ori_n578_), .Y(ori_ori_n1985_));
  NO2        o1936(.A(ori_ori_n1985_), .B(ori_ori_n88_), .Y(ori_ori_n1986_));
  AOI220     o1937(.A0(ori_ori_n1986_), .A1(ori_ori_n1112_), .B0(ori_ori_n1984_), .B1(ori_ori_n1276_), .Y(ori_ori_n1987_));
  NA4        o1938(.A(ori_ori_n1987_), .B(ori_ori_n1983_), .C(ori_ori_n1980_), .D(ori_ori_n1978_), .Y(ori_ori_n1988_));
  AOI210     o1939(.A0(ori_ori_n1971_), .A1(ori_ori_n701_), .B0(ori_ori_n1988_), .Y(ori_ori_n1989_));
  OAI210     o1940(.A0(ori_ori_n1964_), .A1(x2), .B0(ori_ori_n1989_), .Y(ori35));
  NAi21      o1941(.An(ori_ori_n1423_), .B(ori_ori_n1097_), .Y(ori_ori_n1991_));
  NA2        o1942(.A(ori_ori_n194_), .B(ori_ori_n504_), .Y(ori_ori_n1992_));
  NO2        o1943(.A(ori_ori_n383_), .B(ori_ori_n378_), .Y(ori_ori_n1993_));
  AOI220     o1944(.A0(ori_ori_n1993_), .A1(ori_ori_n1992_), .B0(ori_ori_n1991_), .B1(ori_ori_n56_), .Y(ori_ori_n1994_));
  NA2        o1945(.A(x6), .B(ori_ori_n609_), .Y(ori_ori_n1995_));
  NO3        o1946(.A(ori_ori_n599_), .B(ori_ori_n55_), .C(x6), .Y(ori_ori_n1996_));
  OAI210     o1947(.A0(ori_ori_n1996_), .A1(ori_ori_n614_), .B0(ori_ori_n199_), .Y(ori_ori_n1997_));
  NA2        o1948(.A(ori_ori_n1119_), .B(ori_ori_n61_), .Y(ori_ori_n1998_));
  NA2        o1949(.A(x6), .B(ori_ori_n413_), .Y(ori_ori_n1999_));
  NA3        o1950(.A(ori_ori_n1999_), .B(ori_ori_n1998_), .C(ori_ori_n1997_), .Y(ori_ori_n2000_));
  NA3        o1951(.A(ori_ori_n1076_), .B(ori_ori_n646_), .C(x3), .Y(ori_ori_n2001_));
  NO3        o1952(.A(ori_ori_n2001_), .B(ori_ori_n601_), .C(ori_ori_n188_), .Y(ori_ori_n2002_));
  AOI210     o1953(.A0(ori_ori_n2000_), .A1(ori_ori_n50_), .B0(ori_ori_n2002_), .Y(ori_ori_n2003_));
  OAI210     o1954(.A0(ori_ori_n1995_), .A1(ori_ori_n1994_), .B0(ori_ori_n2003_), .Y(ori_ori_n2004_));
  INV        o1955(.A(ori_ori_n2004_), .Y(ori_ori_n2005_));
  NA2        o1956(.A(ori_ori_n832_), .B(ori_ori_n61_), .Y(ori_ori_n2006_));
  NO3        o1957(.A(ori_ori_n908_), .B(ori_ori_n495_), .C(ori_ori_n112_), .Y(ori_ori_n2007_));
  OAI210     o1958(.A0(ori_ori_n144_), .A1(ori_ori_n64_), .B0(ori_ori_n2007_), .Y(ori_ori_n2008_));
  AOI210     o1959(.A0(ori_ori_n2008_), .A1(ori_ori_n2006_), .B0(ori_ori_n50_), .Y(ori_ori_n2009_));
  NA3        o1960(.A(ori_ori_n410_), .B(ori_ori_n752_), .C(ori_ori_n94_), .Y(ori_ori_n2010_));
  OAI210     o1961(.A0(ori_ori_n832_), .A1(ori_ori_n231_), .B0(ori_ori_n647_), .Y(ori_ori_n2011_));
  OAI210     o1962(.A0(ori_ori_n231_), .A1(ori_ori_n516_), .B0(ori_ori_n1812_), .Y(ori_ori_n2012_));
  NA3        o1963(.A(ori_ori_n2012_), .B(ori_ori_n2011_), .C(ori_ori_n2010_), .Y(ori_ori_n2013_));
  OAI210     o1964(.A0(ori_ori_n2013_), .A1(ori_ori_n2009_), .B0(ori_ori_n57_), .Y(ori_ori_n2014_));
  AOI210     o1965(.A0(ori_ori_n742_), .A1(ori_ori_n466_), .B0(ori_ori_n1602_), .Y(ori_ori_n2015_));
  INV        o1966(.A(ori_ori_n2015_), .Y(ori_ori_n2016_));
  NO4        o1967(.A(ori_ori_n825_), .B(ori_ori_n495_), .C(ori_ori_n325_), .D(ori_ori_n364_), .Y(ori_ori_n2017_));
  XN2        o1968(.A(x4), .B(x3), .Y(ori_ori_n2018_));
  NO3        o1969(.A(ori_ori_n2018_), .B(ori_ori_n589_), .C(ori_ori_n280_), .Y(ori_ori_n2019_));
  NO3        o1970(.A(ori_ori_n2019_), .B(ori_ori_n2017_), .C(ori_ori_n1237_), .Y(ori_ori_n2020_));
  OAI210     o1971(.A0(ori_ori_n2016_), .A1(x3), .B0(ori_ori_n2020_), .Y(ori_ori_n2021_));
  NO3        o1972(.A(ori_ori_n641_), .B(ori_ori_n744_), .C(ori_ori_n246_), .Y(ori_ori_n2022_));
  OAI210     o1973(.A0(ori_ori_n2022_), .A1(ori_ori_n1237_), .B0(ori_ori_n50_), .Y(ori_ori_n2023_));
  NA2        o1974(.A(ori_ori_n2171_), .B(ori_ori_n2023_), .Y(ori_ori_n2024_));
  AOI210     o1975(.A0(ori_ori_n2021_), .A1(ori_ori_n519_), .B0(ori_ori_n2024_), .Y(ori_ori_n2025_));
  AOI210     o1976(.A0(ori_ori_n1210_), .A1(ori_ori_n572_), .B0(ori_ori_n601_), .Y(ori_ori_n2026_));
  OAI210     o1977(.A0(ori_ori_n1648_), .A1(ori_ori_n536_), .B0(ori_ori_n1886_), .Y(ori_ori_n2027_));
  OAI210     o1978(.A0(ori_ori_n1950_), .A1(x2), .B0(ori_ori_n2027_), .Y(ori_ori_n2028_));
  OAI210     o1979(.A0(ori_ori_n2028_), .A1(ori_ori_n2026_), .B0(ori_ori_n85_), .Y(ori_ori_n2029_));
  NO2        o1980(.A(ori_ori_n736_), .B(ori_ori_n586_), .Y(ori_ori_n2030_));
  NO2        o1981(.A(ori_ori_n259_), .B(x6), .Y(ori_ori_n2031_));
  OAI210     o1982(.A0(ori_ori_n2030_), .A1(ori_ori_n1495_), .B0(ori_ori_n2031_), .Y(ori_ori_n2032_));
  NA4        o1983(.A(ori_ori_n2032_), .B(ori_ori_n2029_), .C(ori_ori_n2025_), .D(ori_ori_n2014_), .Y(ori_ori_n2033_));
  NA4        o1984(.A(ori_ori_n543_), .B(ori_ori_n604_), .C(ori_ori_n382_), .D(x6), .Y(ori_ori_n2034_));
  AOI210     o1985(.A0(ori_ori_n2034_), .A1(ori_ori_n379_), .B0(x1), .Y(ori_ori_n2035_));
  NO2        o1986(.A(ori_ori_n627_), .B(ori_ori_n601_), .Y(ori_ori_n2036_));
  OAI210     o1987(.A0(ori_ori_n410_), .A1(ori_ori_n152_), .B0(ori_ori_n682_), .Y(ori_ori_n2037_));
  AOI210     o1988(.A0(ori_ori_n2037_), .A1(ori_ori_n881_), .B0(ori_ori_n53_), .Y(ori_ori_n2038_));
  NO3        o1989(.A(ori_ori_n2038_), .B(ori_ori_n2036_), .C(ori_ori_n2035_), .Y(ori_ori_n2039_));
  OAI220     o1990(.A0(ori_ori_n1104_), .A1(x8), .B0(ori_ori_n337_), .B1(ori_ori_n315_), .Y(ori_ori_n2040_));
  AOI210     o1991(.A0(ori_ori_n2040_), .A1(ori_ori_n371_), .B0(ori_ori_n795_), .Y(ori_ori_n2041_));
  OAI210     o1992(.A0(ori_ori_n2039_), .A1(ori_ori_n283_), .B0(ori_ori_n2041_), .Y(ori_ori_n2042_));
  AOI210     o1993(.A0(ori_ori_n2033_), .A1(x5), .B0(ori_ori_n2042_), .Y(ori_ori_n2043_));
  OAI210     o1994(.A0(ori_ori_n2005_), .A1(x5), .B0(ori_ori_n2043_), .Y(ori36));
  NO2        o1995(.A(ori_ori_n744_), .B(ori_ori_n274_), .Y(ori_ori_n2045_));
  NO3        o1996(.A(ori_ori_n111_), .B(ori_ori_n897_), .C(ori_ori_n55_), .Y(ori_ori_n2046_));
  NO3        o1997(.A(ori_ori_n2046_), .B(ori_ori_n1666_), .C(ori_ori_n908_), .Y(ori_ori_n2047_));
  OAI210     o1998(.A0(ori_ori_n2047_), .A1(ori_ori_n2045_), .B0(ori_ori_n100_), .Y(ori_ori_n2048_));
  OR4        o1999(.A(ori_ori_n826_), .B(ori_ori_n692_), .C(ori_ori_n339_), .D(ori_ori_n431_), .Y(ori_ori_n2049_));
  INV        o2000(.A(ori_ori_n869_), .Y(ori_ori_n2050_));
  OAI210     o2001(.A0(ori_ori_n1854_), .A1(ori_ori_n2050_), .B0(ori_ori_n251_), .Y(ori_ori_n2051_));
  NA3        o2002(.A(ori_ori_n395_), .B(ori_ori_n208_), .C(ori_ori_n110_), .Y(ori_ori_n2052_));
  NA4        o2003(.A(ori_ori_n2052_), .B(ori_ori_n2051_), .C(ori_ori_n2049_), .D(ori_ori_n2048_), .Y(ori_ori_n2053_));
  NO2        o2004(.A(ori_ori_n859_), .B(x8), .Y(ori_ori_n2054_));
  NO3        o2005(.A(ori_ori_n2054_), .B(ori_ori_n858_), .C(ori_ori_n471_), .Y(ori_ori_n2055_));
  AOI220     o2006(.A0(ori_ori_n275_), .A1(x1), .B0(ori_ori_n126_), .B1(x6), .Y(ori_ori_n2056_));
  AOI210     o2007(.A0(ori_ori_n929_), .A1(x6), .B0(ori_ori_n375_), .Y(ori_ori_n2057_));
  OAI220     o2008(.A0(ori_ori_n2057_), .A1(ori_ori_n324_), .B0(ori_ori_n2056_), .B1(ori_ori_n411_), .Y(ori_ori_n2058_));
  OAI210     o2009(.A0(ori_ori_n2058_), .A1(ori_ori_n2055_), .B0(ori_ori_n410_), .Y(ori_ori_n2059_));
  NA2        o2010(.A(ori_ori_n592_), .B(ori_ori_n431_), .Y(ori_ori_n2060_));
  AOI210     o2011(.A0(ori_ori_n2060_), .A1(ori_ori_n575_), .B0(ori_ori_n239_), .Y(ori_ori_n2061_));
  NO3        o2012(.A(ori_ori_n1575_), .B(ori_ori_n1358_), .C(ori_ori_n247_), .Y(ori_ori_n2062_));
  NO2        o2013(.A(ori_ori_n2006_), .B(ori_ori_n210_), .Y(ori_ori_n2063_));
  NO4        o2014(.A(ori_ori_n2063_), .B(ori_ori_n2062_), .C(ori_ori_n2061_), .D(ori_ori_n373_), .Y(ori_ori_n2064_));
  OAI210     o2015(.A0(ori_ori_n567_), .A1(ori_ori_n691_), .B0(ori_ori_n850_), .Y(ori_ori_n2065_));
  OAI220     o2016(.A0(ori_ori_n1389_), .A1(ori_ori_n1387_), .B0(ori_ori_n850_), .B1(ori_ori_n929_), .Y(ori_ori_n2066_));
  AOI220     o2017(.A0(ori_ori_n2066_), .A1(ori_ori_n109_), .B0(ori_ori_n2065_), .B1(ori_ori_n557_), .Y(ori_ori_n2067_));
  NA3        o2018(.A(ori_ori_n2067_), .B(ori_ori_n2064_), .C(ori_ori_n2059_), .Y(ori_ori_n2068_));
  AOI210     o2019(.A0(ori_ori_n2053_), .A1(ori_ori_n302_), .B0(ori_ori_n2068_), .Y(ori_ori_n2069_));
  NO3        o2020(.A(ori_ori_n2018_), .B(ori_ori_n782_), .C(ori_ori_n442_), .Y(ori_ori_n2070_));
  AOI210     o2021(.A0(ori_ori_n1079_), .A1(ori_ori_n241_), .B0(ori_ori_n2070_), .Y(ori_ori_n2071_));
  OAI210     o2022(.A0(ori_ori_n750_), .A1(ori_ori_n246_), .B0(ori_ori_n356_), .Y(ori_ori_n2072_));
  NO2        o2023(.A(ori_ori_n542_), .B(ori_ori_n100_), .Y(ori_ori_n2073_));
  AO210      o2024(.A0(ori_ori_n2073_), .A1(ori_ori_n2185_), .B0(ori_ori_n1477_), .Y(ori_ori_n2074_));
  NO2        o2025(.A(ori_ori_n407_), .B(ori_ori_n372_), .Y(ori_ori_n2075_));
  AOI220     o2026(.A0(ori_ori_n2075_), .A1(ori_ori_n2074_), .B0(ori_ori_n2072_), .B1(ori_ori_n266_), .Y(ori_ori_n2076_));
  OAI210     o2027(.A0(ori_ori_n2071_), .A1(x1), .B0(ori_ori_n2076_), .Y(ori_ori_n2077_));
  INV        o2028(.A(ori_ori_n2077_), .Y(ori_ori_n2078_));
  NA2        o2029(.A(ori_ori_n2069_), .B(ori_ori_n2078_), .Y(ori37));
  NO2        o2030(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n2080_));
  AOI220     o2031(.A0(ori_ori_n531_), .A1(ori_ori_n644_), .B0(ori_ori_n410_), .B1(ori_ori_n896_), .Y(ori_ori_n2081_));
  NO2        o2032(.A(ori_ori_n2081_), .B(ori_ori_n100_), .Y(ori_ori_n2082_));
  OAI210     o2033(.A0(ori_ori_n2082_), .A1(ori_ori_n2080_), .B0(ori_ori_n68_), .Y(ori_ori_n2083_));
  NA3        o2034(.A(ori_ori_n154_), .B(ori_ori_n2083_), .C(ori_ori_n605_), .Y(ori_ori_n2084_));
  NA2        o2035(.A(ori_ori_n378_), .B(ori_ori_n126_), .Y(ori_ori_n2085_));
  NO2        o2036(.A(ori_ori_n1445_), .B(ori_ori_n99_), .Y(ori_ori_n2086_));
  AOI210     o2037(.A0(ori_ori_n1668_), .A1(ori_ori_n745_), .B0(ori_ori_n2086_), .Y(ori_ori_n2087_));
  OAI220     o2038(.A0(ori_ori_n2087_), .A1(ori_ori_n51_), .B0(ori_ori_n1360_), .B1(ori_ori_n2085_), .Y(ori_ori_n2088_));
  AOI210     o2039(.A0(ori_ori_n2084_), .A1(ori_ori_n65_), .B0(ori_ori_n2088_), .Y(ori_ori_n2089_));
  OAI210     o2040(.A0(ori_ori_n242_), .A1(ori_ori_n933_), .B0(ori_ori_n425_), .Y(ori_ori_n2090_));
  NA3        o2041(.A(ori_ori_n2090_), .B(ori_ori_n239_), .C(ori_ori_n897_), .Y(ori_ori_n2091_));
  OAI210     o2042(.A0(ori_ori_n211_), .A1(ori_ori_n199_), .B0(ori_ori_n1451_), .Y(ori_ori_n2092_));
  NA2        o2043(.A(ori_ori_n310_), .B(ori_ori_n245_), .Y(ori_ori_n2093_));
  NA3        o2044(.A(ori_ori_n362_), .B(ori_ori_n705_), .C(ori_ori_n100_), .Y(ori_ori_n2094_));
  NO2        o2045(.A(ori_ori_n463_), .B(ori_ori_n56_), .Y(ori_ori_n2095_));
  NA3        o2046(.A(ori_ori_n2095_), .B(ori_ori_n2094_), .C(ori_ori_n2093_), .Y(ori_ori_n2096_));
  AOI210     o2047(.A0(ori_ori_n2092_), .A1(ori_ori_n450_), .B0(ori_ori_n2096_), .Y(ori_ori_n2097_));
  NO2        o2048(.A(ori_ori_n1003_), .B(ori_ori_n246_), .Y(ori_ori_n2098_));
  OAI210     o2049(.A0(ori_ori_n266_), .A1(ori_ori_n237_), .B0(ori_ori_n2098_), .Y(ori_ori_n2099_));
  OAI210     o2050(.A0(ori_ori_n591_), .A1(ori_ori_n127_), .B0(x3), .Y(ori_ori_n2100_));
  AOI210     o2051(.A0(ori_ori_n591_), .A1(ori_ori_n329_), .B0(ori_ori_n2100_), .Y(ori_ori_n2101_));
  AOI210     o2052(.A0(ori_ori_n1359_), .A1(ori_ori_n50_), .B0(ori_ori_n310_), .Y(ori_ori_n2102_));
  OAI210     o2053(.A0(ori_ori_n2102_), .A1(ori_ori_n361_), .B0(ori_ori_n56_), .Y(ori_ori_n2103_));
  NO2        o2054(.A(ori_ori_n2103_), .B(ori_ori_n2101_), .Y(ori_ori_n2104_));
  AOI220     o2055(.A0(ori_ori_n2104_), .A1(ori_ori_n2099_), .B0(ori_ori_n2097_), .B1(ori_ori_n2091_), .Y(ori_ori_n2105_));
  OAI210     o2056(.A0(ori_ori_n2105_), .A1(ori_ori_n1476_), .B0(ori_ori_n93_), .Y(ori_ori_n2106_));
  NO3        o2057(.A(ori_ori_n228_), .B(ori_ori_n316_), .C(ori_ori_n81_), .Y(ori_ori_n2107_));
  NO2        o2058(.A(ori_ori_n249_), .B(ori_ori_n664_), .Y(ori_ori_n2108_));
  NO3        o2059(.A(ori_ori_n2108_), .B(ori_ori_n1020_), .C(ori_ori_n1036_), .Y(ori_ori_n2109_));
  OAI220     o2060(.A0(ori_ori_n2109_), .A1(ori_ori_n2107_), .B0(ori_ori_n410_), .B1(ori_ori_n82_), .Y(ori_ori_n2110_));
  OR2        o2061(.A(ori_ori_n815_), .B(ori_ori_n646_), .Y(ori_ori_n2111_));
  NA2        o2062(.A(ori_ori_n1030_), .B(ori_ori_n55_), .Y(ori_ori_n2112_));
  NOi21      o2063(.An(ori_ori_n2112_), .B(ori_ori_n346_), .Y(ori_ori_n2113_));
  AOI210     o2064(.A0(ori_ori_n2113_), .A1(ori_ori_n2111_), .B0(x1), .Y(ori_ori_n2114_));
  NA2        o2065(.A(ori_ori_n238_), .B(ori_ori_n81_), .Y(ori_ori_n2115_));
  AOI210     o2066(.A0(ori_ori_n1316_), .A1(ori_ori_n361_), .B0(ori_ori_n2115_), .Y(ori_ori_n2116_));
  NA2        o2067(.A(ori_ori_n941_), .B(ori_ori_n60_), .Y(ori_ori_n2117_));
  NA2        o2068(.A(ori_ori_n980_), .B(ori_ori_n157_), .Y(ori_ori_n2118_));
  OAI210     o2069(.A0(ori_ori_n2117_), .A1(ori_ori_n282_), .B0(ori_ori_n2118_), .Y(ori_ori_n2119_));
  NO3        o2070(.A(ori_ori_n2119_), .B(ori_ori_n2116_), .C(ori_ori_n2114_), .Y(ori_ori_n2120_));
  OAI210     o2071(.A0(ori_ori_n2120_), .A1(x6), .B0(ori_ori_n2110_), .Y(ori_ori_n2121_));
  NA2        o2072(.A(ori_ori_n2121_), .B(x5), .Y(ori_ori_n2122_));
  NA3        o2073(.A(ori_ori_n2122_), .B(ori_ori_n2106_), .C(ori_ori_n2089_), .Y(ori38));
  NO2        o2074(.A(ori_ori_n168_), .B(ori_ori_n844_), .Y(ori_ori_n2124_));
  AOI210     o2075(.A0(ori_ori_n1034_), .A1(ori_ori_n509_), .B0(ori_ori_n926_), .Y(ori_ori_n2125_));
  AOI210     o2076(.A0(ori_ori_n2112_), .A1(ori_ori_n1551_), .B0(ori_ori_n210_), .Y(ori_ori_n2126_));
  NO3        o2077(.A(ori_ori_n1096_), .B(ori_ori_n288_), .C(x8), .Y(ori_ori_n2127_));
  NO4        o2078(.A(ori_ori_n2127_), .B(ori_ori_n2126_), .C(ori_ori_n2125_), .D(ori_ori_n2124_), .Y(ori_ori_n2128_));
  NO2        o2079(.A(ori_ori_n2128_), .B(x6), .Y(ori_ori_n2129_));
  NA4        o2080(.A(ori_ori_n340_), .B(ori_ori_n233_), .C(ori_ori_n171_), .D(x8), .Y(ori_ori_n2130_));
  NA2        o2081(.A(ori_ori_n360_), .B(ori_ori_n98_), .Y(ori_ori_n2131_));
  AOI210     o2082(.A0(ori_ori_n2131_), .A1(ori_ori_n2130_), .B0(ori_ori_n130_), .Y(ori_ori_n2132_));
  AOI210     o2083(.A0(ori_ori_n387_), .A1(ori_ori_n363_), .B0(ori_ori_n1457_), .Y(ori_ori_n2133_));
  NO2        o2084(.A(ori_ori_n699_), .B(ori_ori_n85_), .Y(ori_ori_n2134_));
  OAI210     o2085(.A0(ori_ori_n882_), .A1(ori_ori_n136_), .B0(ori_ori_n323_), .Y(ori_ori_n2135_));
  OAI220     o2086(.A0(ori_ori_n2135_), .A1(ori_ori_n2134_), .B0(ori_ori_n2133_), .B1(ori_ori_n171_), .Y(ori_ori_n2136_));
  OAI210     o2087(.A0(ori_ori_n2136_), .A1(ori_ori_n2132_), .B0(x6), .Y(ori_ori_n2137_));
  NO2        o2088(.A(ori_ori_n226_), .B(ori_ori_n664_), .Y(ori_ori_n2138_));
  NO3        o2089(.A(ori_ori_n2138_), .B(ori_ori_n1423_), .C(ori_ori_n233_), .Y(ori_ori_n2139_));
  NO3        o2090(.A(x3), .B(ori_ori_n53_), .C(x0), .Y(ori_ori_n2140_));
  OAI210     o2091(.A0(ori_ori_n458_), .A1(x2), .B0(ori_ori_n2140_), .Y(ori_ori_n2141_));
  NA3        o2092(.A(ori_ori_n386_), .B(ori_ori_n378_), .C(ori_ori_n265_), .Y(ori_ori_n2142_));
  NA2        o2093(.A(ori_ori_n2142_), .B(ori_ori_n2141_), .Y(ori_ori_n2143_));
  OAI210     o2094(.A0(ori_ori_n2143_), .A1(ori_ori_n2139_), .B0(ori_ori_n701_), .Y(ori_ori_n2144_));
  NO2        o2095(.A(ori_ori_n532_), .B(ori_ori_n247_), .Y(ori_ori_n2145_));
  AN3        o2096(.A(ori_ori_n706_), .B(ori_ori_n673_), .C(x0), .Y(ori_ori_n2146_));
  OAI210     o2097(.A0(ori_ori_n2146_), .A1(ori_ori_n2145_), .B0(ori_ori_n294_), .Y(ori_ori_n2147_));
  OAI220     o2098(.A0(ori_ori_n532_), .A1(ori_ori_n247_), .B0(ori_ori_n705_), .B1(ori_ori_n86_), .Y(ori_ori_n2148_));
  OAI210     o2099(.A0(ori_ori_n604_), .A1(x0), .B0(ori_ori_n51_), .Y(ori_ori_n2149_));
  AOI210     o2100(.A0(ori_ori_n515_), .A1(x4), .B0(ori_ori_n209_), .Y(ori_ori_n2150_));
  AOI220     o2101(.A0(ori_ori_n2150_), .A1(ori_ori_n2149_), .B0(ori_ori_n2148_), .B1(ori_ori_n362_), .Y(ori_ori_n2151_));
  NA4        o2102(.A(ori_ori_n2151_), .B(ori_ori_n2147_), .C(ori_ori_n2144_), .D(ori_ori_n2137_), .Y(ori_ori_n2152_));
  OAI210     o2103(.A0(ori_ori_n2152_), .A1(ori_ori_n2129_), .B0(x7), .Y(ori_ori_n2153_));
  AOI210     o2104(.A0(ori_ori_n1529_), .A1(ori_ori_n247_), .B0(ori_ori_n601_), .Y(ori_ori_n2154_));
  OAI210     o2105(.A0(ori_ori_n1475_), .A1(ori_ori_n194_), .B0(ori_ori_n433_), .Y(ori_ori_n2155_));
  OAI210     o2106(.A0(ori_ori_n2155_), .A1(ori_ori_n2154_), .B0(ori_ori_n559_), .Y(ori_ori_n2156_));
  OAI220     o2107(.A0(ori_ori_n1478_), .A1(ori_ori_n247_), .B0(ori_ori_n232_), .B1(ori_ori_n94_), .Y(ori_ori_n2157_));
  NA2        o2108(.A(ori_ori_n1569_), .B(ori_ori_n318_), .Y(ori_ori_n2158_));
  OAI220     o2109(.A0(ori_ori_n2158_), .A1(ori_ori_n567_), .B0(ori_ori_n607_), .B1(ori_ori_n138_), .Y(ori_ori_n2159_));
  AOI210     o2110(.A0(ori_ori_n2157_), .A1(ori_ori_n859_), .B0(ori_ori_n2159_), .Y(ori_ori_n2160_));
  NA3        o2111(.A(ori_ori_n2160_), .B(ori_ori_n2156_), .C(ori_ori_n2153_), .Y(ori39));
  INV        o2112(.A(x7), .Y(ori_ori_n2164_));
  INV        o2113(.A(ori_ori_n685_), .Y(ori_ori_n2165_));
  INV        o2114(.A(x7), .Y(ori_ori_n2166_));
  INV        o2115(.A(ori_ori_n65_), .Y(ori_ori_n2167_));
  INV        o2116(.A(x4), .Y(ori_ori_n2168_));
  INV        o2117(.A(x7), .Y(ori_ori_n2169_));
  INV        o2118(.A(x7), .Y(ori_ori_n2170_));
  INV        o2119(.A(ori_ori_n230_), .Y(ori_ori_n2171_));
  INV        o2120(.A(x5), .Y(ori_ori_n2172_));
  INV        o2121(.A(x6), .Y(ori_ori_n2173_));
  INV        o2122(.A(ori_ori_n230_), .Y(ori_ori_n2174_));
  INV        o2123(.A(x6), .Y(ori_ori_n2175_));
  INV        o2124(.A(ori_ori_n516_), .Y(ori_ori_n2176_));
  INV        o2125(.A(x2), .Y(ori_ori_n2177_));
  INV        o2126(.A(ori_ori_n386_), .Y(ori_ori_n2178_));
  INV        o2127(.A(x7), .Y(ori_ori_n2179_));
  INV        o2128(.A(x2), .Y(ori_ori_n2180_));
  INV        o2129(.A(x7), .Y(ori_ori_n2181_));
  INV        o2130(.A(x8), .Y(ori_ori_n2182_));
  INV        o2131(.A(ori_ori_n521_), .Y(ori_ori_n2183_));
  INV        o2132(.A(x7), .Y(ori_ori_n2184_));
  INV        o2133(.A(ori_ori_n156_), .Y(ori_ori_n2185_));
  INV        o2134(.A(x7), .Y(ori_ori_n2186_));
  INV        o2135(.A(x7), .Y(ori_ori_n2187_));
  INV        o2136(.A(x7), .Y(ori_ori_n2188_));
  INV        m0000(.A(x3), .Y(mai_mai_n50_));
  NA2        m0001(.A(mai_mai_n50_), .B(x2), .Y(mai_mai_n51_));
  NA2        m0002(.A(x7), .B(x0), .Y(mai_mai_n52_));
  INV        m0003(.A(x1), .Y(mai_mai_n53_));
  NA2        m0004(.A(x5), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  INV        m0005(.A(x8), .Y(mai_mai_n55_));
  INV        m0006(.A(x4), .Y(mai_mai_n56_));
  INV        m0007(.A(x7), .Y(mai_mai_n57_));
  NA2        m0008(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0009(.A(x0), .Y(mai_mai_n59_));
  NA2        m0010(.A(x4), .B(mai_mai_n59_), .Y(mai_mai_n60_));
  NA4        m0011(.A(mai_mai_n60_), .B(mai_mai_n58_), .C(mai_mai_n55_), .D(x6), .Y(mai_mai_n61_));
  NA2        m0012(.A(mai_mai_n56_), .B(mai_mai_n59_), .Y(mai_mai_n62_));
  NO2        m0013(.A(mai_mai_n55_), .B(x6), .Y(mai_mai_n63_));
  NA2        m0014(.A(mai_mai_n57_), .B(x4), .Y(mai_mai_n64_));
  NA3        m0015(.A(mai_mai_n64_), .B(mai_mai_n63_), .C(mai_mai_n62_), .Y(mai_mai_n65_));
  AOI210     m0016(.A0(mai_mai_n65_), .A1(mai_mai_n61_), .B0(mai_mai_n54_), .Y(mai_mai_n66_));
  NO2        m0017(.A(x8), .B(mai_mai_n57_), .Y(mai_mai_n67_));
  NO2        m0018(.A(x7), .B(mai_mai_n59_), .Y(mai_mai_n68_));
  NO2        m0019(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  NAi21      m0020(.An(x5), .B(x1), .Y(mai_mai_n70_));
  INV        m0021(.A(x6), .Y(mai_mai_n71_));
  NA2        m0022(.A(mai_mai_n71_), .B(x4), .Y(mai_mai_n72_));
  NO3        m0023(.A(mai_mai_n72_), .B(mai_mai_n70_), .C(mai_mai_n69_), .Y(mai_mai_n73_));
  NO2        m0024(.A(mai_mai_n73_), .B(mai_mai_n66_), .Y(mai_mai_n74_));
  NA2        m0025(.A(x7), .B(x4), .Y(mai_mai_n75_));
  NO2        m0026(.A(mai_mai_n75_), .B(x1), .Y(mai_mai_n76_));
  NO2        m0027(.A(mai_mai_n71_), .B(x5), .Y(mai_mai_n77_));
  NO2        m0028(.A(x8), .B(mai_mai_n59_), .Y(mai_mai_n78_));
  NA2        m0029(.A(mai_mai_n78_), .B(mai_mai_n76_), .Y(mai_mai_n79_));
  AOI210     m0030(.A0(mai_mai_n79_), .A1(mai_mai_n74_), .B0(mai_mai_n51_), .Y(mai_mai_n80_));
  NA2        m0031(.A(x5), .B(x3), .Y(mai_mai_n81_));
  NO2        m0032(.A(x6), .B(x0), .Y(mai_mai_n82_));
  NO2        m0033(.A(mai_mai_n82_), .B(x4), .Y(mai_mai_n83_));
  NO2        m0034(.A(x4), .B(x2), .Y(mai_mai_n84_));
  NO2        m0035(.A(mai_mai_n71_), .B(mai_mai_n59_), .Y(mai_mai_n85_));
  NO2        m0036(.A(mai_mai_n85_), .B(mai_mai_n84_), .Y(mai_mai_n86_));
  NA2        m0037(.A(x8), .B(x1), .Y(mai_mai_n87_));
  NO2        m0038(.A(mai_mai_n87_), .B(x7), .Y(mai_mai_n88_));
  INV        m0039(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  OR3        m0040(.A(mai_mai_n89_), .B(mai_mai_n86_), .C(mai_mai_n83_), .Y(mai_mai_n90_));
  NO3        m0041(.A(x8), .B(mai_mai_n57_), .C(x6), .Y(mai_mai_n91_));
  NO2        m0042(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n92_));
  NO2        m0043(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n93_));
  NA3        m0044(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(mai_mai_n91_), .Y(mai_mai_n94_));
  AOI210     m0045(.A0(mai_mai_n94_), .A1(mai_mai_n90_), .B0(mai_mai_n81_), .Y(mai_mai_n95_));
  XO2        m0046(.A(x7), .B(x1), .Y(mai_mai_n96_));
  INV        m0047(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NO2        m0048(.A(mai_mai_n50_), .B(x0), .Y(mai_mai_n98_));
  NO2        m0049(.A(x6), .B(x5), .Y(mai_mai_n99_));
  NO2        m0050(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n100_));
  NA2        m0051(.A(x6), .B(x1), .Y(mai_mai_n101_));
  NA2        m0052(.A(x3), .B(x0), .Y(mai_mai_n102_));
  INV        m0053(.A(x5), .Y(mai_mai_n103_));
  NA2        m0054(.A(mai_mai_n71_), .B(mai_mai_n103_), .Y(mai_mai_n104_));
  INV        m0055(.A(x2), .Y(mai_mai_n105_));
  NO2        m0056(.A(mai_mai_n56_), .B(mai_mai_n105_), .Y(mai_mai_n106_));
  NA2        m0057(.A(mai_mai_n57_), .B(mai_mai_n103_), .Y(mai_mai_n107_));
  NA3        m0058(.A(mai_mai_n107_), .B(mai_mai_n106_), .C(mai_mai_n104_), .Y(mai_mai_n108_));
  NO3        m0059(.A(mai_mai_n108_), .B(mai_mai_n102_), .C(mai_mai_n53_), .Y(mai_mai_n109_));
  NO3        m0060(.A(mai_mai_n109_), .B(mai_mai_n95_), .C(mai_mai_n80_), .Y(mai00));
  NO2        m0061(.A(x7), .B(x6), .Y(mai_mai_n111_));
  INV        m0062(.A(mai_mai_n111_), .Y(mai_mai_n112_));
  NO2        m0063(.A(mai_mai_n55_), .B(mai_mai_n53_), .Y(mai_mai_n113_));
  NA2        m0064(.A(mai_mai_n113_), .B(mai_mai_n56_), .Y(mai_mai_n114_));
  XN2        m0065(.A(x6), .B(x1), .Y(mai_mai_n115_));
  INV        m0066(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  NO2        m0067(.A(x6), .B(x4), .Y(mai_mai_n117_));
  NA2        m0068(.A(x6), .B(x4), .Y(mai_mai_n118_));
  NAi21      m0069(.An(mai_mai_n117_), .B(mai_mai_n118_), .Y(mai_mai_n119_));
  XN2        m0070(.A(x7), .B(x6), .Y(mai_mai_n120_));
  NO2        m0071(.A(x3), .B(mai_mai_n105_), .Y(mai_mai_n121_));
  NA2        m0072(.A(mai_mai_n121_), .B(mai_mai_n103_), .Y(mai_mai_n122_));
  NA2        m0073(.A(x3), .B(mai_mai_n105_), .Y(mai_mai_n123_));
  NO2        m0074(.A(mai_mai_n55_), .B(mai_mai_n57_), .Y(mai_mai_n124_));
  NA2        m0075(.A(mai_mai_n55_), .B(mai_mai_n57_), .Y(mai_mai_n125_));
  NA2        m0076(.A(mai_mai_n125_), .B(x2), .Y(mai_mai_n126_));
  NA2        m0077(.A(x8), .B(x3), .Y(mai_mai_n127_));
  NA2        m0078(.A(mai_mai_n127_), .B(mai_mai_n75_), .Y(mai_mai_n128_));
  NO2        m0079(.A(mai_mai_n128_), .B(mai_mai_n126_), .Y(mai_mai_n129_));
  NO2        m0080(.A(x5), .B(x0), .Y(mai_mai_n130_));
  NO2        m0081(.A(x6), .B(x1), .Y(mai_mai_n131_));
  NA3        m0082(.A(mai_mai_n131_), .B(mai_mai_n130_), .C(mai_mai_n129_), .Y(mai_mai_n132_));
  NA2        m0083(.A(x8), .B(mai_mai_n103_), .Y(mai_mai_n133_));
  NA2        m0084(.A(x4), .B(mai_mai_n50_), .Y(mai_mai_n134_));
  NAi21      m0085(.An(x7), .B(x2), .Y(mai_mai_n135_));
  XO2        m0086(.A(x8), .B(x7), .Y(mai_mai_n136_));
  NA2        m0087(.A(mai_mai_n136_), .B(mai_mai_n105_), .Y(mai_mai_n137_));
  NA2        m0088(.A(x6), .B(x5), .Y(mai_mai_n138_));
  NO2        m0089(.A(mai_mai_n56_), .B(x0), .Y(mai_mai_n139_));
  NO2        m0090(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n140_));
  NA2        m0091(.A(mai_mai_n140_), .B(mai_mai_n139_), .Y(mai_mai_n141_));
  INV        m0092(.A(mai_mai_n132_), .Y(mai01));
  NA2        m0093(.A(mai_mai_n57_), .B(mai_mai_n59_), .Y(mai_mai_n143_));
  NO2        m0094(.A(x2), .B(x1), .Y(mai_mai_n144_));
  NA2        m0095(.A(x2), .B(x1), .Y(mai_mai_n145_));
  NOi21      m0096(.An(mai_mai_n145_), .B(mai_mai_n144_), .Y(mai_mai_n146_));
  NA2        m0097(.A(mai_mai_n103_), .B(mai_mai_n53_), .Y(mai_mai_n147_));
  NO2        m0098(.A(mai_mai_n147_), .B(x8), .Y(mai_mai_n148_));
  NAi21      m0099(.An(x8), .B(x1), .Y(mai_mai_n149_));
  NO2        m0100(.A(mai_mai_n149_), .B(x3), .Y(mai_mai_n150_));
  OAI210     m0101(.A0(mai_mai_n150_), .A1(mai_mai_n148_), .B0(mai_mai_n146_), .Y(mai_mai_n151_));
  NO2        m0102(.A(x5), .B(mai_mai_n50_), .Y(mai_mai_n152_));
  NO2        m0103(.A(mai_mai_n105_), .B(x1), .Y(mai_mai_n153_));
  NA2        m0104(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  AOI210     m0105(.A0(mai_mai_n154_), .A1(mai_mai_n151_), .B0(mai_mai_n143_), .Y(mai_mai_n155_));
  NAi21      m0106(.An(x7), .B(x0), .Y(mai_mai_n156_));
  NO2        m0107(.A(mai_mai_n55_), .B(x2), .Y(mai_mai_n157_));
  NO2        m0108(.A(mai_mai_n81_), .B(x1), .Y(mai_mai_n158_));
  NA2        m0109(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NA2        m0110(.A(x5), .B(mai_mai_n50_), .Y(mai_mai_n160_));
  NO2        m0111(.A(mai_mai_n160_), .B(mai_mai_n149_), .Y(mai_mai_n161_));
  NA2        m0112(.A(x8), .B(x5), .Y(mai_mai_n162_));
  NO2        m0113(.A(mai_mai_n162_), .B(mai_mai_n51_), .Y(mai_mai_n163_));
  NO3        m0114(.A(x3), .B(mai_mai_n105_), .C(mai_mai_n53_), .Y(mai_mai_n164_));
  NO2        m0115(.A(mai_mai_n163_), .B(mai_mai_n161_), .Y(mai_mai_n165_));
  AOI210     m0116(.A0(mai_mai_n165_), .A1(mai_mai_n159_), .B0(mai_mai_n156_), .Y(mai_mai_n166_));
  NO2        m0117(.A(mai_mai_n57_), .B(x3), .Y(mai_mai_n167_));
  NO2        m0118(.A(mai_mai_n55_), .B(x0), .Y(mai_mai_n168_));
  NA3        m0119(.A(mai_mai_n103_), .B(mai_mai_n105_), .C(x1), .Y(mai_mai_n169_));
  NO2        m0120(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  NO2        m0121(.A(mai_mai_n87_), .B(mai_mai_n50_), .Y(mai_mai_n171_));
  NA2        m0122(.A(mai_mai_n103_), .B(x0), .Y(mai_mai_n172_));
  NA2        m0123(.A(mai_mai_n170_), .B(mai_mai_n167_), .Y(mai_mai_n173_));
  NA2        m0124(.A(x7), .B(mai_mai_n105_), .Y(mai_mai_n174_));
  NA4        m0125(.A(x5), .B(x3), .C(x1), .D(x0), .Y(mai_mai_n175_));
  NAi21      m0126(.An(x1), .B(x2), .Y(mai_mai_n176_));
  NO2        m0127(.A(mai_mai_n160_), .B(mai_mai_n176_), .Y(mai_mai_n177_));
  NA2        m0128(.A(x8), .B(x7), .Y(mai_mai_n178_));
  NO2        m0129(.A(mai_mai_n178_), .B(x0), .Y(mai_mai_n179_));
  OAI210     m0130(.A0(mai_mai_n177_), .A1(x2), .B0(mai_mai_n179_), .Y(mai_mai_n180_));
  NA2        m0131(.A(mai_mai_n180_), .B(mai_mai_n173_), .Y(mai_mai_n181_));
  NO3        m0132(.A(mai_mai_n181_), .B(mai_mai_n166_), .C(mai_mai_n155_), .Y(mai_mai_n182_));
  NA2        m0133(.A(x3), .B(x1), .Y(mai_mai_n183_));
  NA2        m0134(.A(mai_mai_n50_), .B(mai_mai_n105_), .Y(mai_mai_n184_));
  NA2        m0135(.A(mai_mai_n124_), .B(mai_mai_n105_), .Y(mai_mai_n185_));
  XO2        m0136(.A(x5), .B(x3), .Y(mai_mai_n186_));
  NA2        m0137(.A(mai_mai_n186_), .B(x8), .Y(mai_mai_n187_));
  NA2        m0138(.A(x8), .B(mai_mai_n59_), .Y(mai_mai_n188_));
  NA2        m0139(.A(mai_mai_n188_), .B(mai_mai_n127_), .Y(mai_mai_n189_));
  NA2        m0140(.A(x7), .B(mai_mai_n71_), .Y(mai_mai_n190_));
  NO2        m0141(.A(mai_mai_n176_), .B(mai_mai_n190_), .Y(mai_mai_n191_));
  OA210      m0142(.A0(mai_mai_n189_), .A1(mai_mai_n186_), .B0(mai_mai_n191_), .Y(mai_mai_n192_));
  NA2        m0143(.A(mai_mai_n192_), .B(mai_mai_n187_), .Y(mai_mai_n193_));
  OAI210     m0144(.A0(mai_mai_n182_), .A1(mai_mai_n71_), .B0(mai_mai_n193_), .Y(mai_mai_n194_));
  NO2        m0145(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n195_));
  NA4        m0146(.A(mai_mai_n55_), .B(x5), .C(x3), .D(x2), .Y(mai_mai_n196_));
  NA2        m0147(.A(x8), .B(mai_mai_n50_), .Y(mai_mai_n197_));
  NA2        m0148(.A(mai_mai_n197_), .B(x2), .Y(mai_mai_n198_));
  NA2        m0149(.A(mai_mai_n55_), .B(x3), .Y(mai_mai_n199_));
  NA3        m0150(.A(mai_mai_n198_), .B(mai_mai_n186_), .C(mai_mai_n82_), .Y(mai_mai_n200_));
  AOI210     m0151(.A0(mai_mai_n200_), .A1(mai_mai_n196_), .B0(mai_mai_n53_), .Y(mai_mai_n201_));
  NO2        m0152(.A(mai_mai_n105_), .B(mai_mai_n59_), .Y(mai_mai_n202_));
  NA2        m0153(.A(x5), .B(x1), .Y(mai_mai_n203_));
  NO2        m0154(.A(x3), .B(x1), .Y(mai_mai_n204_));
  NO2        m0155(.A(mai_mai_n81_), .B(mai_mai_n55_), .Y(mai_mai_n205_));
  NO2        m0156(.A(x3), .B(x8), .Y(mai_mai_n206_));
  NO2        m0157(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n207_));
  NA2        m0158(.A(mai_mai_n207_), .B(mai_mai_n71_), .Y(mai_mai_n208_));
  NAi21      m0159(.An(x2), .B(x5), .Y(mai_mai_n209_));
  NA2        m0160(.A(x8), .B(x6), .Y(mai_mai_n210_));
  OAI210     m0161(.A0(mai_mai_n210_), .A1(mai_mai_n209_), .B0(mai_mai_n208_), .Y(mai_mai_n211_));
  NA2        m0162(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n212_));
  NO2        m0163(.A(mai_mai_n212_), .B(mai_mai_n59_), .Y(mai_mai_n213_));
  AO220      m0164(.A0(mai_mai_n213_), .A1(mai_mai_n211_), .B0(mai_mai_n206_), .B1(mai_mai_n202_), .Y(mai_mai_n214_));
  OAI210     m0165(.A0(mai_mai_n214_), .A1(mai_mai_n201_), .B0(mai_mai_n195_), .Y(mai_mai_n215_));
  NA2        m0166(.A(mai_mai_n71_), .B(mai_mai_n56_), .Y(mai_mai_n216_));
  NO2        m0167(.A(mai_mai_n216_), .B(x7), .Y(mai_mai_n217_));
  NO2        m0168(.A(mai_mai_n103_), .B(mai_mai_n53_), .Y(mai_mai_n218_));
  NA2        m0169(.A(mai_mai_n218_), .B(mai_mai_n105_), .Y(mai_mai_n219_));
  AOI210     m0170(.A0(mai_mai_n219_), .A1(mai_mai_n154_), .B0(mai_mai_n59_), .Y(mai_mai_n220_));
  NA2        m0171(.A(x3), .B(mai_mai_n59_), .Y(mai_mai_n221_));
  NO2        m0172(.A(mai_mai_n169_), .B(mai_mai_n221_), .Y(mai_mai_n222_));
  OA210      m0173(.A0(mai_mai_n222_), .A1(mai_mai_n220_), .B0(x8), .Y(mai_mai_n223_));
  NO2        m0174(.A(x1), .B(x0), .Y(mai_mai_n224_));
  NA2        m0175(.A(mai_mai_n224_), .B(mai_mai_n105_), .Y(mai_mai_n225_));
  NA2        m0176(.A(mai_mai_n103_), .B(mai_mai_n50_), .Y(mai_mai_n226_));
  NO2        m0177(.A(mai_mai_n103_), .B(x0), .Y(mai_mai_n227_));
  NA2        m0178(.A(x8), .B(mai_mai_n53_), .Y(mai_mai_n228_));
  NO2        m0179(.A(mai_mai_n226_), .B(mai_mai_n225_), .Y(mai_mai_n229_));
  OAI210     m0180(.A0(mai_mai_n229_), .A1(mai_mai_n223_), .B0(mai_mai_n217_), .Y(mai_mai_n230_));
  NO2        m0181(.A(x7), .B(x1), .Y(mai_mai_n231_));
  NOi21      m0182(.An(x8), .B(x3), .Y(mai_mai_n232_));
  NA2        m0183(.A(mai_mai_n232_), .B(mai_mai_n59_), .Y(mai_mai_n233_));
  NA2        m0184(.A(x5), .B(x0), .Y(mai_mai_n234_));
  NAi21      m0185(.An(mai_mai_n130_), .B(mai_mai_n234_), .Y(mai_mai_n235_));
  NA2        m0186(.A(mai_mai_n71_), .B(mai_mai_n50_), .Y(mai_mai_n236_));
  OAI210     m0187(.A0(mai_mai_n236_), .A1(mai_mai_n235_), .B0(mai_mai_n233_), .Y(mai_mai_n237_));
  NA3        m0188(.A(mai_mai_n237_), .B(mai_mai_n133_), .C(mai_mai_n231_), .Y(mai_mai_n238_));
  NA2        m0189(.A(x8), .B(mai_mai_n57_), .Y(mai_mai_n239_));
  NO2        m0190(.A(mai_mai_n239_), .B(x5), .Y(mai_mai_n240_));
  NO2        m0191(.A(mai_mai_n140_), .B(mai_mai_n71_), .Y(mai_mai_n241_));
  NA2        m0192(.A(x1), .B(x0), .Y(mai_mai_n242_));
  NA2        m0193(.A(mai_mai_n50_), .B(mai_mai_n59_), .Y(mai_mai_n243_));
  NA3        m0194(.A(mai_mai_n242_), .B(mai_mai_n241_), .C(mai_mai_n240_), .Y(mai_mai_n244_));
  NA3        m0195(.A(mai_mai_n244_), .B(mai_mai_n238_), .C(mai_mai_n175_), .Y(mai_mai_n245_));
  NO2        m0196(.A(mai_mai_n103_), .B(x3), .Y(mai_mai_n246_));
  NO2        m0197(.A(mai_mai_n105_), .B(x0), .Y(mai_mai_n247_));
  NO2        m0198(.A(mai_mai_n55_), .B(x7), .Y(mai_mai_n248_));
  NO3        m0199(.A(x8), .B(mai_mai_n50_), .C(x0), .Y(mai_mai_n249_));
  NAi21      m0200(.An(x8), .B(x0), .Y(mai_mai_n250_));
  NAi21      m0201(.An(x1), .B(x3), .Y(mai_mai_n251_));
  NO2        m0202(.A(mai_mai_n251_), .B(mai_mai_n250_), .Y(mai_mai_n252_));
  NO2        m0203(.A(x2), .B(mai_mai_n53_), .Y(mai_mai_n253_));
  AOI210     m0204(.A0(mai_mai_n253_), .A1(mai_mai_n249_), .B0(mai_mai_n252_), .Y(mai_mai_n254_));
  NOi21      m0205(.An(x5), .B(x6), .Y(mai_mai_n255_));
  NO2        m0206(.A(mai_mai_n57_), .B(x4), .Y(mai_mai_n256_));
  NA2        m0207(.A(mai_mai_n256_), .B(mai_mai_n255_), .Y(mai_mai_n257_));
  NO2        m0208(.A(mai_mai_n257_), .B(mai_mai_n254_), .Y(mai_mai_n258_));
  AOI210     m0209(.A0(mai_mai_n245_), .A1(mai_mai_n106_), .B0(mai_mai_n258_), .Y(mai_mai_n259_));
  NA3        m0210(.A(mai_mai_n259_), .B(mai_mai_n230_), .C(mai_mai_n215_), .Y(mai_mai_n260_));
  AOI210     m0211(.A0(mai_mai_n194_), .A1(mai_mai_n56_), .B0(mai_mai_n260_), .Y(mai02));
  NO2        m0212(.A(x8), .B(mai_mai_n103_), .Y(mai_mai_n262_));
  XN2        m0213(.A(x7), .B(x3), .Y(mai_mai_n263_));
  NO2        m0214(.A(x2), .B(x0), .Y(mai_mai_n264_));
  NA2        m0215(.A(mai_mai_n264_), .B(mai_mai_n71_), .Y(mai_mai_n265_));
  NO2        m0216(.A(mai_mai_n57_), .B(x1), .Y(mai_mai_n266_));
  NO3        m0217(.A(mai_mai_n266_), .B(mai_mai_n265_), .C(x3), .Y(mai_mai_n267_));
  NA2        m0218(.A(mai_mai_n53_), .B(x0), .Y(mai_mai_n268_));
  NO2        m0219(.A(mai_mai_n251_), .B(x6), .Y(mai_mai_n269_));
  XO2        m0220(.A(x7), .B(x0), .Y(mai_mai_n270_));
  NO2        m0221(.A(mai_mai_n270_), .B(mai_mai_n264_), .Y(mai_mai_n271_));
  AN2        m0222(.A(x7), .B(x2), .Y(mai_mai_n272_));
  NA2        m0223(.A(mai_mai_n272_), .B(mai_mai_n50_), .Y(mai_mai_n273_));
  NA2        m0224(.A(mai_mai_n267_), .B(mai_mai_n262_), .Y(mai_mai_n274_));
  NAi21      m0225(.An(x8), .B(x6), .Y(mai_mai_n275_));
  NO2        m0226(.A(mai_mai_n103_), .B(mai_mai_n59_), .Y(mai_mai_n276_));
  NA2        m0227(.A(x7), .B(x3), .Y(mai_mai_n277_));
  NO2        m0228(.A(mai_mai_n277_), .B(x2), .Y(mai_mai_n278_));
  NA2        m0229(.A(x2), .B(x0), .Y(mai_mai_n279_));
  NA2        m0230(.A(mai_mai_n105_), .B(mai_mai_n59_), .Y(mai_mai_n280_));
  NA2        m0231(.A(mai_mai_n280_), .B(mai_mai_n279_), .Y(mai_mai_n281_));
  NAi21      m0232(.An(x7), .B(x1), .Y(mai_mai_n282_));
  NO2        m0233(.A(mai_mai_n282_), .B(x3), .Y(mai_mai_n283_));
  AOI220     m0234(.A0(mai_mai_n283_), .A1(mai_mai_n281_), .B0(mai_mai_n278_), .B1(mai_mai_n276_), .Y(mai_mai_n284_));
  NA2        m0235(.A(mai_mai_n253_), .B(mai_mai_n50_), .Y(mai_mai_n285_));
  NA3        m0236(.A(x7), .B(mai_mai_n103_), .C(x0), .Y(mai_mai_n286_));
  NA2        m0237(.A(mai_mai_n247_), .B(mai_mai_n53_), .Y(mai_mai_n287_));
  NA2        m0238(.A(mai_mai_n152_), .B(mai_mai_n57_), .Y(mai_mai_n288_));
  OR2        m0239(.A(mai_mai_n288_), .B(mai_mai_n287_), .Y(mai_mai_n289_));
  AOI210     m0240(.A0(mai_mai_n289_), .A1(mai_mai_n284_), .B0(mai_mai_n275_), .Y(mai_mai_n290_));
  INV        m0241(.A(mai_mai_n270_), .Y(mai_mai_n291_));
  NO2        m0242(.A(x7), .B(mai_mai_n71_), .Y(mai_mai_n292_));
  NA2        m0243(.A(mai_mai_n103_), .B(x3), .Y(mai_mai_n293_));
  NO2        m0244(.A(mai_mai_n293_), .B(mai_mai_n292_), .Y(mai_mai_n294_));
  NA2        m0245(.A(mai_mai_n294_), .B(mai_mai_n291_), .Y(mai_mai_n295_));
  NA2        m0246(.A(mai_mai_n50_), .B(x0), .Y(mai_mai_n296_));
  NO2        m0247(.A(mai_mai_n296_), .B(x7), .Y(mai_mai_n297_));
  NA2        m0248(.A(mai_mai_n297_), .B(mai_mai_n255_), .Y(mai_mai_n298_));
  NA2        m0249(.A(mai_mai_n157_), .B(x1), .Y(mai_mai_n299_));
  AOI210     m0250(.A0(mai_mai_n298_), .A1(mai_mai_n295_), .B0(mai_mai_n299_), .Y(mai_mai_n300_));
  NO2        m0251(.A(mai_mai_n57_), .B(mai_mai_n50_), .Y(mai_mai_n301_));
  NO2        m0252(.A(mai_mai_n55_), .B(mai_mai_n105_), .Y(mai_mai_n302_));
  NA3        m0253(.A(mai_mai_n302_), .B(mai_mai_n301_), .C(mai_mai_n59_), .Y(mai_mai_n303_));
  NO2        m0254(.A(mai_mai_n147_), .B(x6), .Y(mai_mai_n304_));
  NO2        m0255(.A(mai_mai_n101_), .B(mai_mai_n103_), .Y(mai_mai_n305_));
  NA2        m0256(.A(mai_mai_n57_), .B(mai_mai_n105_), .Y(mai_mai_n306_));
  NO2        m0257(.A(mai_mai_n306_), .B(mai_mai_n243_), .Y(mai_mai_n307_));
  OAI210     m0258(.A0(mai_mai_n305_), .A1(mai_mai_n304_), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  OAI210     m0259(.A0(mai_mai_n303_), .A1(mai_mai_n101_), .B0(mai_mai_n308_), .Y(mai_mai_n309_));
  NO3        m0260(.A(mai_mai_n309_), .B(mai_mai_n300_), .C(mai_mai_n290_), .Y(mai_mai_n310_));
  AOI210     m0261(.A0(mai_mai_n310_), .A1(mai_mai_n274_), .B0(x4), .Y(mai_mai_n311_));
  NA2        m0262(.A(x8), .B(mai_mai_n71_), .Y(mai_mai_n312_));
  NO2        m0263(.A(x3), .B(mai_mai_n59_), .Y(mai_mai_n313_));
  NA3        m0264(.A(mai_mai_n313_), .B(mai_mai_n103_), .C(mai_mai_n53_), .Y(mai_mai_n314_));
  NO2        m0265(.A(x3), .B(x0), .Y(mai_mai_n315_));
  NAi21      m0266(.An(mai_mai_n315_), .B(mai_mai_n102_), .Y(mai_mai_n316_));
  NA2        m0267(.A(x5), .B(x2), .Y(mai_mai_n317_));
  NO2        m0268(.A(mai_mai_n317_), .B(mai_mai_n204_), .Y(mai_mai_n318_));
  AOI210     m0269(.A0(mai_mai_n318_), .A1(mai_mai_n316_), .B0(mai_mai_n222_), .Y(mai_mai_n319_));
  AO210      m0270(.A0(mai_mai_n319_), .A1(mai_mai_n314_), .B0(mai_mai_n312_), .Y(mai_mai_n320_));
  NO2        m0271(.A(mai_mai_n105_), .B(mai_mai_n53_), .Y(mai_mai_n321_));
  NA2        m0272(.A(mai_mai_n321_), .B(x3), .Y(mai_mai_n322_));
  NO2        m0273(.A(mai_mai_n55_), .B(x1), .Y(mai_mai_n323_));
  NA2        m0274(.A(mai_mai_n323_), .B(mai_mai_n105_), .Y(mai_mai_n324_));
  INV        m0275(.A(mai_mai_n324_), .Y(mai_mai_n325_));
  NAi32      m0276(.An(x3), .Bn(x0), .C(x2), .Y(mai_mai_n326_));
  NO2        m0277(.A(mai_mai_n50_), .B(x2), .Y(mai_mai_n327_));
  NAi21      m0278(.An(x6), .B(x5), .Y(mai_mai_n328_));
  NO2        m0279(.A(x2), .B(mai_mai_n59_), .Y(mai_mai_n329_));
  NO3        m0280(.A(mai_mai_n328_), .B(mai_mai_n149_), .C(mai_mai_n327_), .Y(mai_mai_n330_));
  AOI220     m0281(.A0(mai_mai_n330_), .A1(mai_mai_n326_), .B0(mai_mai_n325_), .B1(mai_mai_n85_), .Y(mai_mai_n331_));
  AOI210     m0282(.A0(mai_mai_n331_), .A1(mai_mai_n320_), .B0(mai_mai_n75_), .Y(mai_mai_n332_));
  NA2        m0283(.A(mai_mai_n323_), .B(mai_mai_n56_), .Y(mai_mai_n333_));
  NO2        m0284(.A(mai_mai_n103_), .B(mai_mai_n50_), .Y(mai_mai_n334_));
  NO2        m0285(.A(mai_mai_n264_), .B(mai_mai_n202_), .Y(mai_mai_n335_));
  XO2        m0286(.A(x7), .B(x2), .Y(mai_mai_n336_));
  INV        m0287(.A(mai_mai_n336_), .Y(mai_mai_n337_));
  XO2        m0288(.A(x6), .B(x2), .Y(mai_mai_n338_));
  NA3        m0289(.A(mai_mai_n337_), .B(mai_mai_n335_), .C(mai_mai_n334_), .Y(mai_mai_n339_));
  NAi21      m0290(.An(x0), .B(x6), .Y(mai_mai_n340_));
  NA2        m0291(.A(mai_mai_n340_), .B(mai_mai_n135_), .Y(mai_mai_n341_));
  XN2        m0292(.A(x7), .B(x5), .Y(mai_mai_n342_));
  NA2        m0293(.A(mai_mai_n342_), .B(mai_mai_n71_), .Y(mai_mai_n343_));
  NA2        m0294(.A(x7), .B(x5), .Y(mai_mai_n344_));
  AOI210     m0295(.A0(mai_mai_n344_), .A1(x6), .B0(mai_mai_n326_), .Y(mai_mai_n345_));
  AOI220     m0296(.A0(mai_mai_n345_), .A1(mai_mai_n343_), .B0(mai_mai_n341_), .B1(mai_mai_n294_), .Y(mai_mai_n346_));
  AOI210     m0297(.A0(mai_mai_n346_), .A1(mai_mai_n339_), .B0(mai_mai_n333_), .Y(mai_mai_n347_));
  NO2        m0298(.A(x8), .B(x6), .Y(mai_mai_n348_));
  NAi21      m0299(.An(mai_mai_n348_), .B(mai_mai_n210_), .Y(mai_mai_n349_));
  AOI210     m0300(.A0(mai_mai_n349_), .A1(mai_mai_n92_), .B0(x3), .Y(mai_mai_n350_));
  NA2        m0301(.A(mai_mai_n103_), .B(x2), .Y(mai_mai_n351_));
  NO2        m0302(.A(mai_mai_n351_), .B(mai_mai_n64_), .Y(mai_mai_n352_));
  NA2        m0303(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n353_));
  NO2        m0304(.A(mai_mai_n353_), .B(mai_mai_n210_), .Y(mai_mai_n354_));
  OAI210     m0305(.A0(mai_mai_n354_), .A1(mai_mai_n50_), .B0(mai_mai_n352_), .Y(mai_mai_n355_));
  NA2        m0306(.A(x4), .B(x2), .Y(mai_mai_n356_));
  NO2        m0307(.A(mai_mai_n356_), .B(mai_mai_n103_), .Y(mai_mai_n357_));
  NAi21      m0308(.An(x1), .B(x6), .Y(mai_mai_n358_));
  NA2        m0309(.A(mai_mai_n315_), .B(mai_mai_n248_), .Y(mai_mai_n359_));
  OAI220     m0310(.A0(mai_mai_n359_), .A1(mai_mai_n358_), .B0(mai_mai_n102_), .B1(mai_mai_n53_), .Y(mai_mai_n360_));
  NA2        m0311(.A(x8), .B(x2), .Y(mai_mai_n361_));
  NO2        m0312(.A(mai_mai_n361_), .B(mai_mai_n50_), .Y(mai_mai_n362_));
  NA2        m0313(.A(mai_mai_n360_), .B(mai_mai_n357_), .Y(mai_mai_n363_));
  OAI210     m0314(.A0(mai_mai_n355_), .A1(mai_mai_n350_), .B0(mai_mai_n363_), .Y(mai_mai_n364_));
  NO4        m0315(.A(mai_mai_n364_), .B(mai_mai_n347_), .C(mai_mai_n332_), .D(mai_mai_n311_), .Y(mai03));
  NAi21      m0316(.An(x2), .B(x0), .Y(mai_mai_n366_));
  NO3        m0317(.A(x8), .B(x6), .C(x4), .Y(mai_mai_n367_));
  INV        m0318(.A(mai_mai_n367_), .Y(mai_mai_n368_));
  NO2        m0319(.A(mai_mai_n368_), .B(mai_mai_n366_), .Y(mai_mai_n369_));
  NA2        m0320(.A(mai_mai_n106_), .B(mai_mai_n59_), .Y(mai_mai_n370_));
  NO2        m0321(.A(mai_mai_n370_), .B(mai_mai_n55_), .Y(mai_mai_n371_));
  NA2        m0322(.A(mai_mai_n371_), .B(mai_mai_n152_), .Y(mai_mai_n372_));
  NA2        m0323(.A(x3), .B(x2), .Y(mai_mai_n373_));
  NO2        m0324(.A(mai_mai_n149_), .B(x0), .Y(mai_mai_n374_));
  NA2        m0325(.A(x8), .B(x0), .Y(mai_mai_n375_));
  NO2        m0326(.A(mai_mai_n375_), .B(x6), .Y(mai_mai_n376_));
  AOI210     m0327(.A0(mai_mai_n376_), .A1(x5), .B0(mai_mai_n374_), .Y(mai_mai_n377_));
  NO2        m0328(.A(mai_mai_n377_), .B(mai_mai_n373_), .Y(mai_mai_n378_));
  NO2        m0329(.A(x5), .B(mai_mai_n59_), .Y(mai_mai_n379_));
  NO2        m0330(.A(x3), .B(x2), .Y(mai_mai_n380_));
  NA2        m0331(.A(mai_mai_n380_), .B(mai_mai_n379_), .Y(mai_mai_n381_));
  NO2        m0332(.A(mai_mai_n53_), .B(x0), .Y(mai_mai_n382_));
  NA2        m0333(.A(mai_mai_n382_), .B(x5), .Y(mai_mai_n383_));
  AOI210     m0334(.A0(mai_mai_n383_), .A1(mai_mai_n381_), .B0(mai_mai_n275_), .Y(mai_mai_n384_));
  NA2        m0335(.A(mai_mai_n233_), .B(mai_mai_n162_), .Y(mai_mai_n385_));
  NO2        m0336(.A(mai_mai_n50_), .B(mai_mai_n59_), .Y(mai_mai_n386_));
  NO2        m0337(.A(mai_mai_n71_), .B(x0), .Y(mai_mai_n387_));
  NO4        m0338(.A(mai_mai_n387_), .B(mai_mai_n386_), .C(x2), .D(mai_mai_n53_), .Y(mai_mai_n388_));
  AO210      m0339(.A0(mai_mai_n388_), .A1(mai_mai_n385_), .B0(mai_mai_n384_), .Y(mai_mai_n389_));
  OAI210     m0340(.A0(mai_mai_n389_), .A1(mai_mai_n378_), .B0(x4), .Y(mai_mai_n390_));
  NO2        m0341(.A(x4), .B(mai_mai_n53_), .Y(mai_mai_n391_));
  NA2        m0342(.A(mai_mai_n391_), .B(mai_mai_n59_), .Y(mai_mai_n392_));
  NA2        m0343(.A(x7), .B(mai_mai_n103_), .Y(mai_mai_n393_));
  NO3        m0344(.A(x5), .B(mai_mai_n53_), .C(x0), .Y(mai_mai_n394_));
  NO2        m0345(.A(x6), .B(mai_mai_n56_), .Y(mai_mai_n395_));
  NO2        m0346(.A(x8), .B(mai_mai_n50_), .Y(mai_mai_n396_));
  AOI220     m0347(.A0(mai_mai_n393_), .A1(mai_mai_n390_), .B0(mai_mai_n372_), .B1(x7), .Y(mai_mai_n397_));
  NA2        m0348(.A(x7), .B(mai_mai_n53_), .Y(mai_mai_n398_));
  NO2        m0349(.A(mai_mai_n232_), .B(mai_mai_n105_), .Y(mai_mai_n399_));
  NO2        m0350(.A(mai_mai_n55_), .B(mai_mai_n59_), .Y(mai_mai_n400_));
  NA2        m0351(.A(mai_mai_n189_), .B(mai_mai_n99_), .Y(mai_mai_n401_));
  NO2        m0352(.A(x5), .B(x2), .Y(mai_mai_n402_));
  NO2        m0353(.A(x8), .B(x3), .Y(mai_mai_n403_));
  NA2        m0354(.A(mai_mai_n403_), .B(mai_mai_n402_), .Y(mai_mai_n404_));
  NO2        m0355(.A(mai_mai_n404_), .B(x6), .Y(mai_mai_n405_));
  NA2        m0356(.A(mai_mai_n188_), .B(x2), .Y(mai_mai_n406_));
  NO3        m0357(.A(mai_mai_n403_), .B(mai_mai_n316_), .C(mai_mai_n328_), .Y(mai_mai_n407_));
  AOI210     m0358(.A0(mai_mai_n407_), .A1(mai_mai_n406_), .B0(mai_mai_n405_), .Y(mai_mai_n408_));
  NA2        m0359(.A(mai_mai_n401_), .B(mai_mai_n408_), .Y(mai_mai_n409_));
  NA2        m0360(.A(mai_mai_n409_), .B(x4), .Y(mai_mai_n410_));
  NA2        m0361(.A(mai_mai_n55_), .B(mai_mai_n59_), .Y(mai_mai_n411_));
  NO2        m0362(.A(mai_mai_n411_), .B(x5), .Y(mai_mai_n412_));
  NAi21      m0363(.An(x4), .B(x6), .Y(mai_mai_n413_));
  NO2        m0364(.A(mai_mai_n55_), .B(mai_mai_n71_), .Y(mai_mai_n414_));
  NO2        m0365(.A(mai_mai_n50_), .B(mai_mai_n105_), .Y(mai_mai_n415_));
  NO2        m0366(.A(mai_mai_n210_), .B(x0), .Y(mai_mai_n416_));
  NO2        m0367(.A(mai_mai_n328_), .B(x8), .Y(mai_mai_n417_));
  OAI210     m0368(.A0(mai_mai_n417_), .A1(mai_mai_n416_), .B0(mai_mai_n415_), .Y(mai_mai_n418_));
  NA2        m0369(.A(mai_mai_n381_), .B(mai_mai_n418_), .Y(mai_mai_n419_));
  NA2        m0370(.A(mai_mai_n419_), .B(mai_mai_n56_), .Y(mai_mai_n420_));
  AOI210     m0371(.A0(mai_mai_n420_), .A1(mai_mai_n410_), .B0(mai_mai_n398_), .Y(mai_mai_n421_));
  NA2        m0372(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n422_));
  NO2        m0373(.A(mai_mai_n71_), .B(mai_mai_n56_), .Y(mai_mai_n423_));
  NA2        m0374(.A(mai_mai_n327_), .B(mai_mai_n59_), .Y(mai_mai_n424_));
  OAI220     m0375(.A0(mai_mai_n424_), .A1(mai_mai_n55_), .B0(mai_mai_n184_), .B1(mai_mai_n250_), .Y(mai_mai_n425_));
  NA2        m0376(.A(mai_mai_n425_), .B(mai_mai_n423_), .Y(mai_mai_n426_));
  NO3        m0377(.A(x6), .B(x4), .C(mai_mai_n50_), .Y(mai_mai_n427_));
  NA2        m0378(.A(mai_mai_n400_), .B(x5), .Y(mai_mai_n428_));
  NO2        m0379(.A(x8), .B(x5), .Y(mai_mai_n429_));
  NAi21      m0380(.An(mai_mai_n429_), .B(mai_mai_n162_), .Y(mai_mai_n430_));
  NA2        m0381(.A(mai_mai_n280_), .B(mai_mai_n428_), .Y(mai_mai_n431_));
  NA2        m0382(.A(mai_mai_n335_), .B(mai_mai_n77_), .Y(mai_mai_n432_));
  NOi21      m0383(.An(x3), .B(x4), .Y(mai_mai_n433_));
  NA2        m0384(.A(mai_mai_n55_), .B(mai_mai_n105_), .Y(mai_mai_n434_));
  NA2        m0385(.A(mai_mai_n434_), .B(mai_mai_n433_), .Y(mai_mai_n435_));
  NO2        m0386(.A(mai_mai_n51_), .B(x6), .Y(mai_mai_n436_));
  NO2        m0387(.A(mai_mai_n138_), .B(mai_mai_n55_), .Y(mai_mai_n437_));
  NO3        m0388(.A(mai_mai_n56_), .B(x2), .C(x0), .Y(mai_mai_n438_));
  AOI220     m0389(.A0(mai_mai_n438_), .A1(mai_mai_n437_), .B0(mai_mai_n436_), .B1(mai_mai_n412_), .Y(mai_mai_n439_));
  OAI210     m0390(.A0(mai_mai_n435_), .A1(mai_mai_n432_), .B0(mai_mai_n439_), .Y(mai_mai_n440_));
  AOI210     m0391(.A0(mai_mai_n431_), .A1(mai_mai_n427_), .B0(mai_mai_n440_), .Y(mai_mai_n441_));
  AOI210     m0392(.A0(mai_mai_n441_), .A1(mai_mai_n426_), .B0(mai_mai_n422_), .Y(mai_mai_n442_));
  NA2        m0393(.A(x7), .B(x1), .Y(mai_mai_n443_));
  NO3        m0394(.A(x5), .B(x4), .C(x2), .Y(mai_mai_n444_));
  NO2        m0395(.A(x4), .B(mai_mai_n105_), .Y(mai_mai_n445_));
  NA3        m0396(.A(mai_mai_n103_), .B(x4), .C(mai_mai_n105_), .Y(mai_mai_n446_));
  NA2        m0397(.A(mai_mai_n433_), .B(mai_mai_n71_), .Y(mai_mai_n447_));
  NA2        m0398(.A(mai_mai_n157_), .B(mai_mai_n59_), .Y(mai_mai_n448_));
  NO2        m0399(.A(mai_mai_n448_), .B(mai_mai_n447_), .Y(mai_mai_n449_));
  NA2        m0400(.A(mai_mai_n415_), .B(x4), .Y(mai_mai_n450_));
  NO3        m0401(.A(mai_mai_n450_), .B(mai_mai_n348_), .C(mai_mai_n387_), .Y(mai_mai_n451_));
  NO2        m0402(.A(mai_mai_n451_), .B(mai_mai_n449_), .Y(mai_mai_n452_));
  NA2        m0403(.A(x5), .B(x4), .Y(mai_mai_n453_));
  NO2        m0404(.A(mai_mai_n71_), .B(mai_mai_n53_), .Y(mai_mai_n454_));
  NO3        m0405(.A(x8), .B(x3), .C(x2), .Y(mai_mai_n455_));
  NA3        m0406(.A(mai_mai_n455_), .B(mai_mai_n454_), .C(mai_mai_n59_), .Y(mai_mai_n456_));
  NO3        m0407(.A(x6), .B(x5), .C(x2), .Y(mai_mai_n457_));
  NO2        m0408(.A(mai_mai_n456_), .B(mai_mai_n453_), .Y(mai_mai_n458_));
  NA2        m0409(.A(mai_mai_n71_), .B(x2), .Y(mai_mai_n459_));
  NO3        m0410(.A(x4), .B(x3), .C(mai_mai_n59_), .Y(mai_mai_n460_));
  NA2        m0411(.A(mai_mai_n460_), .B(mai_mai_n207_), .Y(mai_mai_n461_));
  NO3        m0412(.A(mai_mai_n461_), .B(mai_mai_n459_), .C(mai_mai_n96_), .Y(mai_mai_n462_));
  XO2        m0413(.A(x4), .B(x0), .Y(mai_mai_n463_));
  NA2        m0414(.A(mai_mai_n243_), .B(x5), .Y(mai_mai_n464_));
  NO2        m0415(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n465_));
  NO2        m0416(.A(mai_mai_n465_), .B(mai_mai_n63_), .Y(mai_mai_n466_));
  NO4        m0417(.A(mai_mai_n466_), .B(mai_mai_n464_), .C(mai_mai_n463_), .D(mai_mai_n145_), .Y(mai_mai_n467_));
  NO3        m0418(.A(mai_mai_n467_), .B(mai_mai_n462_), .C(mai_mai_n458_), .Y(mai_mai_n468_));
  OAI210     m0419(.A0(mai_mai_n452_), .A1(mai_mai_n443_), .B0(mai_mai_n468_), .Y(mai_mai_n469_));
  NO4        m0420(.A(mai_mai_n469_), .B(mai_mai_n442_), .C(mai_mai_n421_), .D(mai_mai_n397_), .Y(mai04));
  NO2        m0421(.A(x7), .B(x2), .Y(mai_mai_n471_));
  NO2        m0422(.A(x3), .B(mai_mai_n53_), .Y(mai_mai_n472_));
  NO2        m0423(.A(mai_mai_n472_), .B(mai_mai_n140_), .Y(mai_mai_n473_));
  XN2        m0424(.A(x8), .B(x1), .Y(mai_mai_n474_));
  NO2        m0425(.A(mai_mai_n474_), .B(mai_mai_n138_), .Y(mai_mai_n475_));
  NA2        m0426(.A(mai_mai_n475_), .B(mai_mai_n473_), .Y(mai_mai_n476_));
  NA2        m0427(.A(x6), .B(x3), .Y(mai_mai_n477_));
  NO2        m0428(.A(mai_mai_n477_), .B(x5), .Y(mai_mai_n478_));
  NA2        m0429(.A(mai_mai_n71_), .B(x1), .Y(mai_mai_n479_));
  NO2        m0430(.A(mai_mai_n429_), .B(mai_mai_n232_), .Y(mai_mai_n480_));
  NO3        m0431(.A(mai_mai_n480_), .B(mai_mai_n403_), .C(mai_mai_n479_), .Y(mai_mai_n481_));
  AOI210     m0432(.A0(mai_mai_n478_), .A1(mai_mai_n323_), .B0(mai_mai_n481_), .Y(mai_mai_n482_));
  AOI210     m0433(.A0(mai_mai_n482_), .A1(mai_mai_n476_), .B0(x0), .Y(mai_mai_n483_));
  NOi21      m0434(.An(mai_mai_n162_), .B(mai_mai_n429_), .Y(mai_mai_n484_));
  NO3        m0435(.A(mai_mai_n2222_), .B(mai_mai_n484_), .C(mai_mai_n296_), .Y(mai_mai_n485_));
  OAI210     m0436(.A0(mai_mai_n485_), .A1(mai_mai_n483_), .B0(mai_mai_n471_), .Y(mai_mai_n486_));
  NA2        m0437(.A(mai_mai_n127_), .B(mai_mai_n221_), .Y(mai_mai_n487_));
  OR3        m0438(.A(mai_mai_n349_), .B(mai_mai_n82_), .C(mai_mai_n54_), .Y(mai_mai_n488_));
  OR2        m0439(.A(x6), .B(x0), .Y(mai_mai_n489_));
  NO3        m0440(.A(mai_mai_n489_), .B(x3), .C(x1), .Y(mai_mai_n490_));
  AOI220     m0441(.A0(mai_mai_n490_), .A1(mai_mai_n103_), .B0(mai_mai_n255_), .B1(mai_mai_n249_), .Y(mai_mai_n491_));
  AOI210     m0442(.A0(mai_mai_n491_), .A1(mai_mai_n488_), .B0(mai_mai_n174_), .Y(mai_mai_n492_));
  NA2        m0443(.A(x7), .B(x2), .Y(mai_mai_n493_));
  INV        m0444(.A(mai_mai_n127_), .Y(mai_mai_n494_));
  NA2        m0445(.A(mai_mai_n494_), .B(mai_mai_n82_), .Y(mai_mai_n495_));
  NO2        m0446(.A(mai_mai_n293_), .B(mai_mai_n55_), .Y(mai_mai_n496_));
  NO3        m0447(.A(x3), .B(x1), .C(x0), .Y(mai_mai_n497_));
  OR2        m0448(.A(x6), .B(x1), .Y(mai_mai_n498_));
  NA2        m0449(.A(mai_mai_n498_), .B(x0), .Y(mai_mai_n499_));
  AOI220     m0450(.A0(mai_mai_n499_), .A1(mai_mai_n496_), .B0(mai_mai_n497_), .B1(mai_mai_n437_), .Y(mai_mai_n500_));
  AOI210     m0451(.A0(mai_mai_n500_), .A1(mai_mai_n495_), .B0(mai_mai_n493_), .Y(mai_mai_n501_));
  NA2        m0452(.A(mai_mai_n71_), .B(x0), .Y(mai_mai_n502_));
  NOi31      m0453(.An(mai_mai_n318_), .B(mai_mai_n502_), .C(mai_mai_n239_), .Y(mai_mai_n503_));
  NO4        m0454(.A(mai_mai_n503_), .B(mai_mai_n501_), .C(mai_mai_n492_), .D(mai_mai_n56_), .Y(mai_mai_n504_));
  NA2        m0455(.A(mai_mai_n504_), .B(mai_mai_n486_), .Y(mai_mai_n505_));
  NA3        m0456(.A(x8), .B(x7), .C(x0), .Y(mai_mai_n506_));
  INV        m0457(.A(mai_mai_n506_), .Y(mai_mai_n507_));
  NA2        m0458(.A(mai_mai_n400_), .B(mai_mai_n57_), .Y(mai_mai_n508_));
  NO2        m0459(.A(x8), .B(x0), .Y(mai_mai_n509_));
  NA2        m0460(.A(mai_mai_n509_), .B(mai_mai_n337_), .Y(mai_mai_n510_));
  AOI210     m0461(.A0(mai_mai_n510_), .A1(mai_mai_n508_), .B0(mai_mai_n251_), .Y(mai_mai_n511_));
  NA2        m0462(.A(mai_mai_n511_), .B(mai_mai_n255_), .Y(mai_mai_n512_));
  NO2        m0463(.A(mai_mai_n71_), .B(mai_mai_n105_), .Y(mai_mai_n513_));
  NO2        m0464(.A(mai_mai_n344_), .B(x8), .Y(mai_mai_n514_));
  INV        m0465(.A(mai_mai_n240_), .Y(mai_mai_n515_));
  NO2        m0466(.A(mai_mai_n515_), .B(mai_mai_n353_), .Y(mai_mai_n516_));
  NO2        m0467(.A(mai_mai_n57_), .B(mai_mai_n59_), .Y(mai_mai_n517_));
  OAI210     m0468(.A0(mai_mai_n517_), .A1(mai_mai_n516_), .B0(mai_mai_n513_), .Y(mai_mai_n518_));
  NO2        m0469(.A(x8), .B(x2), .Y(mai_mai_n519_));
  NO2        m0470(.A(mai_mai_n204_), .B(mai_mai_n57_), .Y(mai_mai_n520_));
  NO2        m0471(.A(mai_mai_n225_), .B(mai_mai_n127_), .Y(mai_mai_n521_));
  AOI210     m0472(.A0(mai_mai_n297_), .A1(mai_mai_n153_), .B0(mai_mai_n521_), .Y(mai_mai_n522_));
  NO2        m0473(.A(mai_mai_n522_), .B(mai_mai_n104_), .Y(mai_mai_n523_));
  NA2        m0474(.A(mai_mai_n313_), .B(x2), .Y(mai_mai_n524_));
  NO2        m0475(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n525_));
  NA2        m0476(.A(mai_mai_n525_), .B(mai_mai_n63_), .Y(mai_mai_n526_));
  AOI210     m0477(.A0(mai_mai_n524_), .A1(mai_mai_n424_), .B0(mai_mai_n526_), .Y(mai_mai_n527_));
  NA2        m0478(.A(mai_mai_n105_), .B(mai_mai_n53_), .Y(mai_mai_n528_));
  NA2        m0479(.A(x7), .B(mai_mai_n50_), .Y(mai_mai_n529_));
  NO2        m0480(.A(mai_mai_n172_), .B(mai_mai_n529_), .Y(mai_mai_n530_));
  NA2        m0481(.A(mai_mai_n379_), .B(mai_mai_n140_), .Y(mai_mai_n531_));
  NO2        m0482(.A(mai_mai_n71_), .B(x2), .Y(mai_mai_n532_));
  NA2        m0483(.A(mai_mai_n532_), .B(mai_mai_n248_), .Y(mai_mai_n533_));
  OAI210     m0484(.A0(mai_mai_n533_), .A1(mai_mai_n531_), .B0(mai_mai_n56_), .Y(mai_mai_n534_));
  NO3        m0485(.A(mai_mai_n534_), .B(mai_mai_n527_), .C(mai_mai_n523_), .Y(mai_mai_n535_));
  NA3        m0486(.A(mai_mai_n535_), .B(mai_mai_n518_), .C(mai_mai_n512_), .Y(mai_mai_n536_));
  NA2        m0487(.A(mai_mai_n53_), .B(mai_mai_n59_), .Y(mai_mai_n537_));
  NOi21      m0488(.An(x2), .B(x7), .Y(mai_mai_n538_));
  NO2        m0489(.A(x6), .B(x3), .Y(mai_mai_n539_));
  NA2        m0490(.A(mai_mai_n539_), .B(mai_mai_n538_), .Y(mai_mai_n540_));
  NO2        m0491(.A(x6), .B(mai_mai_n59_), .Y(mai_mai_n541_));
  NO3        m0492(.A(mai_mai_n57_), .B(x2), .C(x1), .Y(mai_mai_n542_));
  NO3        m0493(.A(mai_mai_n57_), .B(x2), .C(x0), .Y(mai_mai_n543_));
  NA2        m0494(.A(mai_mai_n542_), .B(mai_mai_n541_), .Y(mai_mai_n544_));
  OAI210     m0495(.A0(mai_mai_n540_), .A1(mai_mai_n537_), .B0(mai_mai_n544_), .Y(mai_mai_n545_));
  NO2        m0496(.A(mai_mai_n99_), .B(mai_mai_n53_), .Y(mai_mai_n546_));
  NA2        m0497(.A(mai_mai_n203_), .B(mai_mai_n57_), .Y(mai_mai_n547_));
  OAI210     m0498(.A0(mai_mai_n546_), .A1(mai_mai_n417_), .B0(mai_mai_n547_), .Y(mai_mai_n548_));
  NO3        m0499(.A(mai_mai_n548_), .B(mai_mai_n450_), .C(mai_mai_n59_), .Y(mai_mai_n549_));
  AO210      m0500(.A0(mai_mai_n545_), .A1(mai_mai_n429_), .B0(mai_mai_n549_), .Y(mai_mai_n550_));
  AOI210     m0501(.A0(mai_mai_n536_), .A1(mai_mai_n505_), .B0(mai_mai_n550_), .Y(mai05));
  NO2        m0502(.A(x7), .B(mai_mai_n103_), .Y(mai_mai_n552_));
  NO2        m0503(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n553_));
  NA2        m0504(.A(x5), .B(mai_mai_n56_), .Y(mai_mai_n554_));
  NO2        m0505(.A(mai_mai_n554_), .B(mai_mai_n529_), .Y(mai_mai_n555_));
  AOI210     m0506(.A0(mai_mai_n553_), .A1(mai_mai_n552_), .B0(mai_mai_n555_), .Y(mai_mai_n556_));
  NO2        m0507(.A(mai_mai_n556_), .B(mai_mai_n105_), .Y(mai_mai_n557_));
  NO2        m0508(.A(x7), .B(x4), .Y(mai_mai_n558_));
  NO2        m0509(.A(mai_mai_n64_), .B(mai_mai_n55_), .Y(mai_mai_n559_));
  NO2        m0510(.A(mai_mai_n184_), .B(x5), .Y(mai_mai_n560_));
  NA2        m0511(.A(mai_mai_n103_), .B(mai_mai_n105_), .Y(mai_mai_n561_));
  AN2        m0512(.A(mai_mai_n560_), .B(mai_mai_n559_), .Y(mai_mai_n562_));
  OAI210     m0513(.A0(mai_mai_n562_), .A1(mai_mai_n557_), .B0(mai_mai_n454_), .Y(mai_mai_n563_));
  NO2        m0514(.A(x6), .B(mai_mai_n50_), .Y(mai_mai_n564_));
  NA2        m0515(.A(mai_mai_n55_), .B(x4), .Y(mai_mai_n565_));
  NO2        m0516(.A(mai_mai_n103_), .B(mai_mai_n105_), .Y(mai_mai_n566_));
  NA2        m0517(.A(mai_mai_n566_), .B(x7), .Y(mai_mai_n567_));
  NA2        m0518(.A(mai_mai_n402_), .B(mai_mai_n231_), .Y(mai_mai_n568_));
  NA2        m0519(.A(mai_mai_n568_), .B(mai_mai_n567_), .Y(mai_mai_n569_));
  NA2        m0520(.A(mai_mai_n103_), .B(x4), .Y(mai_mai_n570_));
  XO2        m0521(.A(x7), .B(x5), .Y(mai_mai_n571_));
  NO2        m0522(.A(mai_mai_n103_), .B(x2), .Y(mai_mai_n572_));
  NO2        m0523(.A(mai_mai_n75_), .B(mai_mai_n55_), .Y(mai_mai_n573_));
  NA2        m0524(.A(mai_mai_n569_), .B(mai_mai_n564_), .Y(mai_mai_n574_));
  NO2        m0525(.A(mai_mai_n71_), .B(mai_mai_n50_), .Y(mai_mai_n575_));
  NO2        m0526(.A(mai_mai_n178_), .B(x4), .Y(mai_mai_n576_));
  NO2        m0527(.A(x5), .B(mai_mai_n56_), .Y(mai_mai_n577_));
  NO3        m0528(.A(x8), .B(x7), .C(mai_mai_n105_), .Y(mai_mai_n578_));
  AN2        m0529(.A(mai_mai_n578_), .B(mai_mai_n577_), .Y(mai_mai_n579_));
  NA3        m0530(.A(mai_mai_n579_), .B(mai_mai_n575_), .C(mai_mai_n53_), .Y(mai_mai_n580_));
  NA2        m0531(.A(mai_mai_n246_), .B(mai_mai_n538_), .Y(mai_mai_n581_));
  NOi21      m0532(.An(x4), .B(x1), .Y(mai_mai_n582_));
  NA2        m0533(.A(mai_mai_n582_), .B(mai_mai_n63_), .Y(mai_mai_n583_));
  NA2        m0534(.A(x4), .B(x1), .Y(mai_mai_n584_));
  NO2        m0535(.A(mai_mai_n584_), .B(mai_mai_n50_), .Y(mai_mai_n585_));
  AOI210     m0536(.A0(mai_mai_n585_), .A1(mai_mai_n566_), .B0(mai_mai_n59_), .Y(mai_mai_n586_));
  OA210      m0537(.A0(mai_mai_n583_), .A1(mai_mai_n581_), .B0(mai_mai_n586_), .Y(mai_mai_n587_));
  NA4        m0538(.A(mai_mai_n587_), .B(mai_mai_n580_), .C(mai_mai_n574_), .D(mai_mai_n563_), .Y(mai_mai_n588_));
  NA2        m0539(.A(mai_mai_n575_), .B(mai_mai_n56_), .Y(mai_mai_n589_));
  NA2        m0540(.A(mai_mai_n519_), .B(mai_mai_n552_), .Y(mai_mai_n590_));
  NO2        m0541(.A(mai_mai_n590_), .B(mai_mai_n589_), .Y(mai_mai_n591_));
  NA2        m0542(.A(mai_mai_n248_), .B(mai_mai_n117_), .Y(mai_mai_n592_));
  NA2        m0543(.A(mai_mai_n57_), .B(x6), .Y(mai_mai_n593_));
  AOI210     m0544(.A0(mai_mai_n593_), .A1(x3), .B0(mai_mai_n91_), .Y(mai_mai_n594_));
  NA2        m0545(.A(mai_mai_n577_), .B(mai_mai_n144_), .Y(mai_mai_n595_));
  NO3        m0546(.A(mai_mai_n595_), .B(mai_mai_n594_), .C(mai_mai_n396_), .Y(mai_mai_n596_));
  NA2        m0547(.A(mai_mai_n256_), .B(mai_mai_n71_), .Y(mai_mai_n597_));
  NO2        m0548(.A(mai_mai_n361_), .B(x3), .Y(mai_mai_n598_));
  NA2        m0549(.A(mai_mai_n598_), .B(mai_mai_n218_), .Y(mai_mai_n599_));
  NO2        m0550(.A(mai_mai_n396_), .B(mai_mai_n576_), .Y(mai_mai_n600_));
  NO2        m0551(.A(mai_mai_n433_), .B(mai_mai_n103_), .Y(mai_mai_n601_));
  NO2        m0552(.A(mai_mai_n528_), .B(x6), .Y(mai_mai_n602_));
  NA2        m0553(.A(mai_mai_n602_), .B(mai_mai_n601_), .Y(mai_mai_n603_));
  OAI220     m0554(.A0(mai_mai_n603_), .A1(mai_mai_n600_), .B0(mai_mai_n599_), .B1(mai_mai_n597_), .Y(mai_mai_n604_));
  NO4        m0555(.A(mai_mai_n604_), .B(mai_mai_n596_), .C(x0), .D(mai_mai_n591_), .Y(mai_mai_n605_));
  NA2        m0556(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n606_));
  NO2        m0557(.A(mai_mai_n606_), .B(x1), .Y(mai_mai_n607_));
  NA2        m0558(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n608_));
  NO2        m0559(.A(mai_mai_n608_), .B(mai_mai_n123_), .Y(mai_mai_n609_));
  NA2        m0560(.A(x8), .B(x4), .Y(mai_mai_n610_));
  NO2        m0561(.A(x8), .B(x4), .Y(mai_mai_n611_));
  NAi21      m0562(.An(mai_mai_n611_), .B(mai_mai_n610_), .Y(mai_mai_n612_));
  NAi21      m0563(.An(mai_mai_n519_), .B(mai_mai_n361_), .Y(mai_mai_n613_));
  NO4        m0564(.A(mai_mai_n613_), .B(mai_mai_n612_), .C(mai_mai_n396_), .D(mai_mai_n71_), .Y(mai_mai_n614_));
  OAI210     m0565(.A0(mai_mai_n614_), .A1(mai_mai_n609_), .B0(mai_mai_n607_), .Y(mai_mai_n615_));
  NO3        m0566(.A(x8), .B(mai_mai_n103_), .C(x4), .Y(mai_mai_n616_));
  INV        m0567(.A(mai_mai_n616_), .Y(mai_mai_n617_));
  NO2        m0568(.A(mai_mai_n617_), .B(mai_mai_n105_), .Y(mai_mai_n618_));
  NO2        m0569(.A(x5), .B(x4), .Y(mai_mai_n619_));
  NO2        m0570(.A(x6), .B(mai_mai_n105_), .Y(mai_mai_n620_));
  NA2        m0571(.A(mai_mai_n608_), .B(mai_mai_n620_), .Y(mai_mai_n621_));
  NO2        m0572(.A(mai_mai_n621_), .B(mai_mai_n484_), .Y(mai_mai_n622_));
  OAI210     m0573(.A0(mai_mai_n622_), .A1(mai_mai_n618_), .B0(mai_mai_n283_), .Y(mai_mai_n623_));
  NA3        m0574(.A(mai_mai_n623_), .B(mai_mai_n615_), .C(mai_mai_n605_), .Y(mai_mai_n624_));
  OR2        m0575(.A(x4), .B(x1), .Y(mai_mai_n625_));
  NO2        m0576(.A(mai_mai_n625_), .B(x3), .Y(mai_mai_n626_));
  NA2        m0577(.A(mai_mai_n55_), .B(x2), .Y(mai_mai_n627_));
  NO3        m0578(.A(mai_mai_n342_), .B(mai_mai_n627_), .C(x6), .Y(mai_mai_n628_));
  AOI220     m0579(.A0(mai_mai_n628_), .A1(mai_mai_n626_), .B0(mai_mai_n624_), .B1(mai_mai_n588_), .Y(mai06));
  NA2        m0580(.A(mai_mai_n56_), .B(x3), .Y(mai_mai_n630_));
  NA2        m0581(.A(x6), .B(mai_mai_n105_), .Y(mai_mai_n631_));
  NA2        m0582(.A(mai_mai_n631_), .B(mai_mai_n55_), .Y(mai_mai_n632_));
  NA2        m0583(.A(x5), .B(mai_mai_n59_), .Y(mai_mai_n633_));
  NO2        m0584(.A(mai_mai_n633_), .B(mai_mai_n113_), .Y(mai_mai_n634_));
  NA3        m0585(.A(mai_mai_n634_), .B(mai_mai_n632_), .C(mai_mai_n459_), .Y(mai_mai_n635_));
  NO2        m0586(.A(mai_mai_n361_), .B(x0), .Y(mai_mai_n636_));
  NA2        m0587(.A(mai_mai_n312_), .B(x2), .Y(mai_mai_n637_));
  NOi21      m0588(.An(x6), .B(x8), .Y(mai_mai_n638_));
  NO2        m0589(.A(mai_mai_n638_), .B(x2), .Y(mai_mai_n639_));
  NO3        m0590(.A(mai_mai_n639_), .B(mai_mai_n70_), .C(mai_mai_n59_), .Y(mai_mai_n640_));
  AOI220     m0591(.A0(mai_mai_n640_), .A1(mai_mai_n637_), .B0(mai_mai_n636_), .B1(mai_mai_n304_), .Y(mai_mai_n641_));
  AOI210     m0592(.A0(mai_mai_n641_), .A1(mai_mai_n635_), .B0(mai_mai_n630_), .Y(mai_mai_n642_));
  NA2        m0593(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n643_));
  NA2        m0594(.A(mai_mai_n340_), .B(mai_mai_n328_), .Y(mai_mai_n644_));
  NO2        m0595(.A(mai_mai_n71_), .B(mai_mai_n103_), .Y(mai_mai_n645_));
  NO2        m0596(.A(mai_mai_n53_), .B(mai_mai_n59_), .Y(mai_mai_n646_));
  NO4        m0597(.A(mai_mai_n646_), .B(mai_mai_n627_), .C(mai_mai_n645_), .D(mai_mai_n454_), .Y(mai_mai_n647_));
  AOI220     m0598(.A0(mai_mai_n647_), .A1(mai_mai_n644_), .B0(mai_mai_n394_), .B1(mai_mai_n63_), .Y(mai_mai_n648_));
  NO2        m0599(.A(mai_mai_n648_), .B(mai_mai_n643_), .Y(mai_mai_n649_));
  NO2        m0600(.A(mai_mai_n54_), .B(x0), .Y(mai_mai_n650_));
  NA2        m0601(.A(x4), .B(x3), .Y(mai_mai_n651_));
  OAI210     m0602(.A0(mai_mai_n651_), .A1(x8), .B0(mai_mai_n477_), .Y(mai_mai_n652_));
  NA2        m0603(.A(mai_mai_n652_), .B(mai_mai_n650_), .Y(mai_mai_n653_));
  NO2        m0604(.A(mai_mai_n101_), .B(mai_mai_n56_), .Y(mai_mai_n654_));
  NA3        m0605(.A(mai_mai_n654_), .B(mai_mai_n232_), .C(mai_mai_n379_), .Y(mai_mai_n655_));
  AOI210     m0606(.A0(mai_mai_n655_), .A1(mai_mai_n653_), .B0(x2), .Y(mai_mai_n656_));
  INV        m0607(.A(mai_mai_n357_), .Y(mai_mai_n657_));
  NO2        m0608(.A(mai_mai_n382_), .B(x8), .Y(mai_mai_n658_));
  NO2        m0609(.A(mai_mai_n233_), .B(mai_mai_n479_), .Y(mai_mai_n659_));
  AOI210     m0610(.A0(mai_mai_n658_), .A1(mai_mai_n241_), .B0(mai_mai_n659_), .Y(mai_mai_n660_));
  NO2        m0611(.A(x5), .B(x3), .Y(mai_mai_n661_));
  NA3        m0612(.A(mai_mai_n509_), .B(mai_mai_n661_), .C(x1), .Y(mai_mai_n662_));
  NA2        m0613(.A(mai_mai_n553_), .B(mai_mai_n513_), .Y(mai_mai_n663_));
  OA220      m0614(.A0(mai_mai_n663_), .A1(mai_mai_n531_), .B0(mai_mai_n662_), .B1(mai_mai_n459_), .Y(mai_mai_n664_));
  OAI210     m0615(.A0(mai_mai_n660_), .A1(mai_mai_n657_), .B0(mai_mai_n664_), .Y(mai_mai_n665_));
  OR4        m0616(.A(mai_mai_n665_), .B(mai_mai_n656_), .C(mai_mai_n649_), .D(mai_mai_n642_), .Y(mai_mai_n666_));
  NA2        m0617(.A(x7), .B(mai_mai_n56_), .Y(mai_mai_n667_));
  NO2        m0618(.A(mai_mai_n566_), .B(mai_mai_n59_), .Y(mai_mai_n668_));
  NO2        m0619(.A(mai_mai_n160_), .B(x6), .Y(mai_mai_n669_));
  NA2        m0620(.A(mai_mai_n669_), .B(mai_mai_n264_), .Y(mai_mai_n670_));
  NO2        m0621(.A(mai_mai_n670_), .B(mai_mai_n667_), .Y(mai_mai_n671_));
  NA2        m0622(.A(mai_mai_n671_), .B(mai_mai_n323_), .Y(mai_mai_n672_));
  NO2        m0623(.A(mai_mai_n279_), .B(mai_mai_n103_), .Y(mai_mai_n673_));
  NO2        m0624(.A(mai_mai_n56_), .B(x3), .Y(mai_mai_n674_));
  NA2        m0625(.A(mai_mai_n674_), .B(mai_mai_n71_), .Y(mai_mai_n675_));
  NO2        m0626(.A(mai_mai_n675_), .B(mai_mai_n228_), .Y(mai_mai_n676_));
  NO2        m0627(.A(mai_mai_n71_), .B(x3), .Y(mai_mai_n677_));
  NA3        m0628(.A(mai_mai_n677_), .B(mai_mai_n525_), .C(mai_mai_n56_), .Y(mai_mai_n678_));
  NO2        m0629(.A(mai_mai_n57_), .B(x6), .Y(mai_mai_n679_));
  NA3        m0630(.A(mai_mai_n553_), .B(mai_mai_n301_), .C(mai_mai_n71_), .Y(mai_mai_n680_));
  NA2        m0631(.A(mai_mai_n680_), .B(mai_mai_n678_), .Y(mai_mai_n681_));
  OR3        m0632(.A(mai_mai_n681_), .B(mai_mai_n676_), .C(mai_mai_n585_), .Y(mai_mai_n682_));
  NA2        m0633(.A(mai_mai_n682_), .B(mai_mai_n673_), .Y(mai_mai_n683_));
  NA3        m0634(.A(mai_mai_n242_), .B(mai_mai_n539_), .C(mai_mai_n234_), .Y(mai_mai_n684_));
  NA2        m0635(.A(mai_mai_n445_), .B(mai_mai_n67_), .Y(mai_mai_n685_));
  AOI210     m0636(.A0(mai_mai_n684_), .A1(mai_mai_n71_), .B0(mai_mai_n685_), .Y(mai_mai_n686_));
  NA2        m0637(.A(x7), .B(x6), .Y(mai_mai_n687_));
  NA3        m0638(.A(x2), .B(x1), .C(x0), .Y(mai_mai_n688_));
  NA2        m0639(.A(mai_mai_n455_), .B(mai_mai_n139_), .Y(mai_mai_n689_));
  NO2        m0640(.A(x5), .B(x1), .Y(mai_mai_n690_));
  NA2        m0641(.A(mai_mai_n690_), .B(mai_mai_n679_), .Y(mai_mai_n691_));
  NA2        m0642(.A(x4), .B(x0), .Y(mai_mai_n692_));
  NO3        m0643(.A(mai_mai_n57_), .B(x6), .C(x2), .Y(mai_mai_n693_));
  NO2        m0644(.A(mai_mai_n691_), .B(mai_mai_n689_), .Y(mai_mai_n694_));
  NO2        m0645(.A(mai_mai_n694_), .B(mai_mai_n686_), .Y(mai_mai_n695_));
  NA3        m0646(.A(mai_mai_n695_), .B(mai_mai_n683_), .C(mai_mai_n672_), .Y(mai_mai_n696_));
  AOI210     m0647(.A0(mai_mai_n666_), .A1(mai_mai_n57_), .B0(mai_mai_n696_), .Y(mai07));
  NA2        m0648(.A(mai_mai_n103_), .B(mai_mai_n59_), .Y(mai_mai_n698_));
  NOi21      m0649(.An(mai_mai_n687_), .B(mai_mai_n111_), .Y(mai_mai_n699_));
  NO3        m0650(.A(mai_mai_n57_), .B(x5), .C(x1), .Y(mai_mai_n700_));
  NA2        m0651(.A(mai_mai_n700_), .B(mai_mai_n348_), .Y(mai_mai_n701_));
  NO2        m0652(.A(mai_mai_n57_), .B(mai_mai_n71_), .Y(mai_mai_n702_));
  NO2        m0653(.A(mai_mai_n143_), .B(mai_mai_n104_), .Y(mai_mai_n703_));
  AOI210     m0654(.A0(mai_mai_n702_), .A1(mai_mai_n92_), .B0(mai_mai_n703_), .Y(mai_mai_n704_));
  OAI220     m0655(.A0(mai_mai_n704_), .A1(mai_mai_n127_), .B0(mai_mai_n701_), .B1(mai_mai_n296_), .Y(mai_mai_n705_));
  NA2        m0656(.A(mai_mai_n705_), .B(x2), .Y(mai_mai_n706_));
  NAi21      m0657(.An(mai_mai_n144_), .B(mai_mai_n145_), .Y(mai_mai_n707_));
  NA2        m0658(.A(mai_mai_n91_), .B(x3), .Y(mai_mai_n708_));
  NO3        m0659(.A(mai_mai_n55_), .B(x3), .C(x1), .Y(mai_mai_n709_));
  NO2        m0660(.A(mai_mai_n472_), .B(x2), .Y(mai_mai_n710_));
  AOI210     m0661(.A0(mai_mai_n710_), .A1(mai_mai_n474_), .B0(mai_mai_n709_), .Y(mai_mai_n711_));
  OAI210     m0662(.A0(mai_mai_n711_), .A1(mai_mai_n593_), .B0(mai_mai_n708_), .Y(mai_mai_n712_));
  NO2        m0663(.A(x8), .B(mai_mai_n53_), .Y(mai_mai_n713_));
  NA2        m0664(.A(mai_mai_n713_), .B(mai_mai_n59_), .Y(mai_mai_n714_));
  NO2        m0665(.A(x7), .B(x3), .Y(mai_mai_n715_));
  NA2        m0666(.A(mai_mai_n715_), .B(mai_mai_n99_), .Y(mai_mai_n716_));
  NO2        m0667(.A(mai_mai_n714_), .B(mai_mai_n716_), .Y(mai_mai_n717_));
  AOI210     m0668(.A0(mai_mai_n712_), .A1(mai_mai_n227_), .B0(mai_mai_n717_), .Y(mai_mai_n718_));
  AOI210     m0669(.A0(mai_mai_n718_), .A1(mai_mai_n706_), .B0(x4), .Y(mai_mai_n719_));
  NA3        m0670(.A(mai_mai_n690_), .B(mai_mai_n292_), .C(mai_mai_n55_), .Y(mai_mai_n720_));
  AOI210     m0671(.A0(mai_mai_n720_), .A1(mai_mai_n548_), .B0(mai_mai_n105_), .Y(mai_mai_n721_));
  XO2        m0672(.A(x5), .B(x1), .Y(mai_mai_n722_));
  NA2        m0673(.A(mai_mai_n721_), .B(mai_mai_n386_), .Y(mai_mai_n723_));
  NO3        m0674(.A(mai_mai_n50_), .B(x2), .C(x0), .Y(mai_mai_n724_));
  NO2        m0675(.A(mai_mai_n282_), .B(mai_mai_n103_), .Y(mai_mai_n725_));
  NA2        m0676(.A(x6), .B(x0), .Y(mai_mai_n726_));
  NO2        m0677(.A(mai_mai_n627_), .B(mai_mai_n726_), .Y(mai_mai_n727_));
  NO2        m0678(.A(mai_mai_n722_), .B(mai_mai_n638_), .Y(mai_mai_n728_));
  OAI210     m0679(.A0(mai_mai_n690_), .A1(mai_mai_n63_), .B0(mai_mai_n57_), .Y(mai_mai_n729_));
  OAI210     m0680(.A0(mai_mai_n729_), .A1(mai_mai_n728_), .B0(mai_mai_n701_), .Y(mai_mai_n730_));
  AOI220     m0681(.A0(mai_mai_n730_), .A1(mai_mai_n724_), .B0(mai_mai_n727_), .B1(mai_mai_n725_), .Y(mai_mai_n731_));
  AOI210     m0682(.A0(mai_mai_n731_), .A1(mai_mai_n723_), .B0(mai_mai_n56_), .Y(mai_mai_n732_));
  NOi21      m0683(.An(mai_mai_n210_), .B(mai_mai_n348_), .Y(mai_mai_n733_));
  NO3        m0684(.A(mai_mai_n733_), .B(mai_mai_n219_), .C(mai_mai_n67_), .Y(mai_mai_n734_));
  NO2        m0685(.A(mai_mai_n282_), .B(x6), .Y(mai_mai_n735_));
  AN2        m0686(.A(mai_mai_n735_), .B(mai_mai_n302_), .Y(mai_mai_n736_));
  OAI210     m0687(.A0(mai_mai_n736_), .A1(mai_mai_n734_), .B0(mai_mai_n59_), .Y(mai_mai_n737_));
  NA2        m0688(.A(mai_mai_n92_), .B(mai_mai_n71_), .Y(mai_mai_n738_));
  NO2        m0689(.A(mai_mai_n738_), .B(mai_mai_n590_), .Y(mai_mai_n739_));
  NAi21      m0690(.An(x8), .B(x7), .Y(mai_mai_n740_));
  NA2        m0691(.A(mai_mai_n733_), .B(mai_mai_n740_), .Y(mai_mai_n741_));
  NA2        m0692(.A(mai_mai_n379_), .B(mai_mai_n105_), .Y(mai_mai_n742_));
  NO3        m0693(.A(mai_mai_n2216_), .B(mai_mai_n742_), .C(mai_mai_n525_), .Y(mai_mai_n743_));
  AOI210     m0694(.A0(mai_mai_n743_), .A1(mai_mai_n741_), .B0(mai_mai_n739_), .Y(mai_mai_n744_));
  AOI210     m0695(.A0(mai_mai_n744_), .A1(mai_mai_n737_), .B0(mai_mai_n134_), .Y(mai_mai_n745_));
  NO2        m0696(.A(x8), .B(x7), .Y(mai_mai_n746_));
  NO2        m0697(.A(mai_mai_n746_), .B(x3), .Y(mai_mai_n747_));
  NA3        m0698(.A(mai_mai_n747_), .B(mai_mai_n337_), .C(x1), .Y(mai_mai_n748_));
  NO2        m0699(.A(x8), .B(mai_mai_n105_), .Y(mai_mai_n749_));
  NA2        m0700(.A(mai_mai_n749_), .B(mai_mai_n231_), .Y(mai_mai_n750_));
  NO2        m0701(.A(mai_mai_n71_), .B(x4), .Y(mai_mai_n751_));
  NA2        m0702(.A(mai_mai_n751_), .B(mai_mai_n276_), .Y(mai_mai_n752_));
  AOI210     m0703(.A0(mai_mai_n750_), .A1(mai_mai_n748_), .B0(mai_mai_n752_), .Y(mai_mai_n753_));
  NO4        m0704(.A(mai_mai_n753_), .B(mai_mai_n745_), .C(mai_mai_n732_), .D(mai_mai_n719_), .Y(mai08));
  NA2        m0705(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n755_));
  XN2        m0706(.A(x5), .B(x4), .Y(mai_mai_n756_));
  INV        m0707(.A(mai_mai_n756_), .Y(mai_mai_n757_));
  NO2        m0708(.A(mai_mai_n221_), .B(mai_mai_n103_), .Y(mai_mai_n758_));
  NA2        m0709(.A(mai_mai_n253_), .B(mai_mai_n139_), .Y(mai_mai_n759_));
  NO2        m0710(.A(mai_mai_n759_), .B(mai_mai_n187_), .Y(mai_mai_n760_));
  INV        m0711(.A(mai_mai_n760_), .Y(mai_mai_n761_));
  NO2        m0712(.A(mai_mai_n761_), .B(mai_mai_n71_), .Y(mai_mai_n762_));
  NO2        m0713(.A(mai_mai_n746_), .B(mai_mai_n105_), .Y(mai_mai_n763_));
  NA2        m0714(.A(mai_mai_n763_), .B(mai_mai_n178_), .Y(mai_mai_n764_));
  OAI210     m0715(.A0(mai_mai_n382_), .A1(mai_mai_n276_), .B0(mai_mai_n316_), .Y(mai_mai_n765_));
  NA2        m0716(.A(mai_mai_n402_), .B(mai_mai_n212_), .Y(mai_mai_n766_));
  OAI220     m0717(.A0(x8), .A1(mai_mai_n766_), .B0(mai_mai_n765_), .B1(mai_mai_n764_), .Y(mai_mai_n767_));
  NA2        m0718(.A(mai_mai_n767_), .B(mai_mai_n263_), .Y(mai_mai_n768_));
  NA2        m0719(.A(mai_mai_n306_), .B(mai_mai_n53_), .Y(mai_mai_n769_));
  NO3        m0720(.A(mai_mai_n382_), .B(mai_mai_n127_), .C(mai_mai_n68_), .Y(mai_mai_n770_));
  NO2        m0721(.A(mai_mai_n646_), .B(mai_mai_n224_), .Y(mai_mai_n771_));
  NO3        m0722(.A(mai_mai_n520_), .B(mai_mai_n434_), .C(mai_mai_n98_), .Y(mai_mai_n772_));
  AO220      m0723(.A0(mai_mai_n772_), .A1(mai_mai_n771_), .B0(mai_mai_n770_), .B1(mai_mai_n769_), .Y(mai_mai_n773_));
  NA2        m0724(.A(x7), .B(mai_mai_n59_), .Y(mai_mai_n774_));
  NO3        m0725(.A(mai_mai_n285_), .B(mai_mai_n774_), .C(mai_mai_n262_), .Y(mai_mai_n775_));
  AOI210     m0726(.A0(mai_mai_n773_), .A1(x5), .B0(mai_mai_n775_), .Y(mai_mai_n776_));
  AOI210     m0727(.A0(mai_mai_n776_), .A1(mai_mai_n768_), .B0(mai_mai_n72_), .Y(mai_mai_n777_));
  NO2        m0728(.A(mai_mai_n70_), .B(x3), .Y(mai_mai_n778_));
  OAI210     m0729(.A0(mai_mai_n778_), .A1(mai_mai_n240_), .B0(mai_mai_n137_), .Y(mai_mai_n779_));
  INV        m0730(.A(mai_mai_n514_), .Y(mai_mai_n780_));
  NO3        m0731(.A(x6), .B(x4), .C(x0), .Y(mai_mai_n781_));
  INV        m0732(.A(mai_mai_n781_), .Y(mai_mai_n782_));
  AOI210     m0733(.A0(mai_mai_n780_), .A1(mai_mai_n779_), .B0(mai_mai_n782_), .Y(mai_mai_n783_));
  NO3        m0734(.A(x5), .B(x3), .C(mai_mai_n105_), .Y(mai_mai_n784_));
  AOI220     m0735(.A0(mai_mai_n757_), .A1(mai_mai_n281_), .B0(mai_mai_n784_), .B1(mai_mai_n59_), .Y(mai_mai_n785_));
  OR2        m0736(.A(x8), .B(x1), .Y(mai_mai_n786_));
  NO3        m0737(.A(mai_mai_n786_), .B(mai_mai_n785_), .C(mai_mai_n674_), .Y(mai_mai_n787_));
  NAi21      m0738(.An(x4), .B(x1), .Y(mai_mai_n788_));
  NO2        m0739(.A(mai_mai_n788_), .B(x0), .Y(mai_mai_n789_));
  NA2        m0740(.A(mai_mai_n560_), .B(mai_mai_n789_), .Y(mai_mai_n790_));
  NA3        m0741(.A(mai_mai_n55_), .B(x1), .C(x0), .Y(mai_mai_n791_));
  OAI210     m0742(.A0(mai_mai_n791_), .A1(mai_mai_n657_), .B0(mai_mai_n790_), .Y(mai_mai_n792_));
  OAI210     m0743(.A0(mai_mai_n792_), .A1(mai_mai_n787_), .B0(mai_mai_n292_), .Y(mai_mai_n793_));
  AO210      m0744(.A0(mai_mai_n264_), .A1(mai_mai_n240_), .B0(mai_mai_n673_), .Y(mai_mai_n794_));
  NA2        m0745(.A(mai_mai_n103_), .B(mai_mai_n56_), .Y(mai_mai_n795_));
  NO2        m0746(.A(mai_mai_n795_), .B(mai_mai_n236_), .Y(mai_mai_n796_));
  NO2        m0747(.A(mai_mai_n57_), .B(x2), .Y(mai_mai_n797_));
  NO4        m0748(.A(mai_mai_n302_), .B(mai_mai_n797_), .C(mai_mai_n746_), .D(mai_mai_n268_), .Y(mai_mai_n798_));
  AOI220     m0749(.A0(mai_mai_n798_), .A1(mai_mai_n796_), .B0(mai_mai_n794_), .B1(mai_mai_n585_), .Y(mai_mai_n799_));
  NA2        m0750(.A(mai_mai_n799_), .B(mai_mai_n793_), .Y(mai_mai_n800_));
  NO4        m0751(.A(mai_mai_n800_), .B(mai_mai_n783_), .C(mai_mai_n777_), .D(mai_mai_n762_), .Y(mai09));
  NO3        m0752(.A(mai_mai_n722_), .B(mai_mai_n115_), .C(mai_mai_n96_), .Y(mai_mai_n802_));
  AOI220     m0753(.A0(mai_mai_n272_), .A1(mai_mai_n70_), .B0(mai_mai_n538_), .B1(mai_mai_n498_), .Y(mai_mai_n803_));
  OAI210     m0754(.A0(mai_mai_n802_), .A1(x2), .B0(mai_mai_n803_), .Y(mai_mai_n804_));
  AOI210     m0755(.A0(mai_mai_n804_), .A1(mai_mai_n691_), .B0(mai_mai_n411_), .Y(mai_mai_n805_));
  NO2        m0756(.A(mai_mai_n537_), .B(mai_mai_n239_), .Y(mai_mai_n806_));
  NO2        m0757(.A(mai_mai_n690_), .B(mai_mai_n312_), .Y(mai_mai_n807_));
  NO3        m0758(.A(mai_mai_n552_), .B(mai_mai_n100_), .C(mai_mai_n105_), .Y(mai_mai_n808_));
  AO220      m0759(.A0(mai_mai_n808_), .A1(mai_mai_n807_), .B0(mai_mai_n806_), .B1(mai_mai_n566_), .Y(mai_mai_n809_));
  OAI210     m0760(.A0(mai_mai_n809_), .A1(mai_mai_n805_), .B0(x4), .Y(mai_mai_n810_));
  NAi21      m0761(.An(x0), .B(x2), .Y(mai_mai_n811_));
  NO2        m0762(.A(mai_mai_n275_), .B(mai_mai_n811_), .Y(mai_mai_n812_));
  NA2        m0763(.A(mai_mai_n812_), .B(mai_mai_n56_), .Y(mai_mai_n813_));
  NO2        m0764(.A(mai_mai_n56_), .B(mai_mai_n59_), .Y(mai_mai_n814_));
  INV        m0765(.A(mai_mai_n120_), .Y(mai_mai_n815_));
  NA2        m0766(.A(mai_mai_n690_), .B(mai_mai_n55_), .Y(mai_mai_n816_));
  AOI210     m0767(.A0(x6), .A1(x1), .B0(x5), .Y(mai_mai_n817_));
  OAI210     m0768(.A0(mai_mai_n817_), .A1(mai_mai_n305_), .B0(x2), .Y(mai_mai_n818_));
  AOI210     m0769(.A0(mai_mai_n818_), .A1(mai_mai_n816_), .B0(mai_mai_n815_), .Y(mai_mai_n819_));
  NA2        m0770(.A(mai_mai_n513_), .B(mai_mai_n55_), .Y(mai_mai_n820_));
  NO4        m0771(.A(mai_mai_n57_), .B(x6), .C(x5), .D(x1), .Y(mai_mai_n821_));
  NO2        m0772(.A(mai_mai_n209_), .B(mai_mai_n358_), .Y(mai_mai_n822_));
  NO2        m0773(.A(mai_mai_n282_), .B(mai_mai_n138_), .Y(mai_mai_n823_));
  NO3        m0774(.A(mai_mai_n823_), .B(mai_mai_n822_), .C(mai_mai_n821_), .Y(mai_mai_n824_));
  OAI220     m0775(.A0(mai_mai_n824_), .A1(mai_mai_n55_), .B0(mai_mai_n820_), .B1(mai_mai_n422_), .Y(mai_mai_n825_));
  OAI210     m0776(.A0(mai_mai_n825_), .A1(mai_mai_n819_), .B0(mai_mai_n814_), .Y(mai_mai_n826_));
  NO2        m0777(.A(mai_mai_n375_), .B(mai_mai_n103_), .Y(mai_mai_n827_));
  NO2        m0778(.A(mai_mai_n306_), .B(mai_mai_n454_), .Y(mai_mai_n828_));
  AOI220     m0779(.A0(mai_mai_n828_), .A1(mai_mai_n827_), .B0(mai_mai_n191_), .B1(mai_mai_n207_), .Y(mai_mai_n829_));
  NA4        m0780(.A(mai_mai_n829_), .B(mai_mai_n826_), .C(mai_mai_n813_), .D(mai_mai_n810_), .Y(mai_mai_n830_));
  NA2        m0781(.A(mai_mai_n830_), .B(mai_mai_n50_), .Y(mai_mai_n831_));
  NO2        m0782(.A(mai_mai_n351_), .B(mai_mai_n149_), .Y(mai_mai_n832_));
  NA2        m0783(.A(mai_mai_n218_), .B(mai_mai_n538_), .Y(mai_mai_n833_));
  OAI210     m0784(.A0(mai_mai_n398_), .A1(mai_mai_n749_), .B0(mai_mai_n833_), .Y(mai_mai_n834_));
  OAI210     m0785(.A0(mai_mai_n834_), .A1(mai_mai_n832_), .B0(x0), .Y(mai_mai_n835_));
  NO3        m0786(.A(x8), .B(x7), .C(x2), .Y(mai_mai_n836_));
  NO3        m0787(.A(mai_mai_n57_), .B(x5), .C(x2), .Y(mai_mai_n837_));
  OAI210     m0788(.A0(mai_mai_n837_), .A1(mai_mai_n836_), .B0(mai_mai_n474_), .Y(mai_mai_n838_));
  AOI210     m0789(.A0(mai_mai_n838_), .A1(mai_mai_n835_), .B0(x4), .Y(mai_mai_n839_));
  NO2        m0790(.A(mai_mai_n103_), .B(mai_mai_n56_), .Y(mai_mai_n840_));
  NA2        m0791(.A(mai_mai_n839_), .B(mai_mai_n564_), .Y(mai_mai_n841_));
  NA2        m0792(.A(mai_mai_n565_), .B(mai_mai_n317_), .Y(mai_mai_n842_));
  NA2        m0793(.A(mai_mai_n56_), .B(mai_mai_n301_), .Y(mai_mai_n843_));
  AOI220     m0794(.A0(mai_mai_n610_), .A1(mai_mai_n321_), .B0(mai_mai_n323_), .B1(mai_mai_n93_), .Y(mai_mai_n844_));
  NA2        m0795(.A(mai_mai_n93_), .B(x5), .Y(mai_mai_n845_));
  OAI220     m0796(.A0(mai_mai_n845_), .A1(mai_mai_n786_), .B0(mai_mai_n844_), .B1(mai_mai_n293_), .Y(mai_mai_n846_));
  NA2        m0797(.A(mai_mai_n846_), .B(mai_mai_n68_), .Y(mai_mai_n847_));
  NA2        m0798(.A(mai_mai_n227_), .B(mai_mai_n153_), .Y(mai_mai_n848_));
  NO2        m0799(.A(mai_mai_n403_), .B(x2), .Y(mai_mai_n849_));
  NO2        m0800(.A(x7), .B(mai_mai_n53_), .Y(mai_mai_n850_));
  NA2        m0801(.A(mai_mai_n850_), .B(x5), .Y(mai_mai_n851_));
  NO2        m0802(.A(mai_mai_n851_), .B(mai_mai_n60_), .Y(mai_mai_n852_));
  AOI220     m0803(.A0(mai_mai_n852_), .A1(mai_mai_n849_), .B0(mai_mai_n611_), .B1(mai_mai_n222_), .Y(mai_mai_n853_));
  NA3        m0804(.A(mai_mai_n853_), .B(mai_mai_n847_), .C(mai_mai_n843_), .Y(mai_mai_n854_));
  NO4        m0805(.A(mai_mai_n842_), .B(mai_mai_n577_), .C(mai_mai_n422_), .D(mai_mai_n50_), .Y(mai_mai_n855_));
  AOI220     m0806(.A0(mai_mai_n553_), .A1(mai_mai_n552_), .B0(mai_mai_n256_), .B1(x5), .Y(mai_mai_n856_));
  NO2        m0807(.A(mai_mai_n619_), .B(mai_mai_n176_), .Y(mai_mai_n857_));
  NO2        m0808(.A(mai_mai_n856_), .B(mai_mai_n322_), .Y(mai_mai_n858_));
  OAI210     m0809(.A0(mai_mai_n858_), .A1(mai_mai_n855_), .B0(mai_mai_n82_), .Y(mai_mai_n859_));
  NA2        m0810(.A(mai_mai_n713_), .B(x2), .Y(mai_mai_n860_));
  NO2        m0811(.A(mai_mai_n860_), .B(mai_mai_n58_), .Y(mai_mai_n861_));
  NO2        m0812(.A(x5), .B(mai_mai_n53_), .Y(mai_mai_n862_));
  NAi21      m0813(.An(x1), .B(x4), .Y(mai_mai_n863_));
  INV        m0814(.A(mai_mai_n863_), .Y(mai_mai_n864_));
  NA2        m0815(.A(mai_mai_n861_), .B(mai_mai_n386_), .Y(mai_mai_n865_));
  NA3        m0816(.A(mai_mai_n369_), .B(mai_mai_n690_), .C(mai_mai_n57_), .Y(mai_mai_n866_));
  NA3        m0817(.A(mai_mai_n866_), .B(mai_mai_n865_), .C(mai_mai_n859_), .Y(mai_mai_n867_));
  AOI210     m0818(.A0(mai_mai_n854_), .A1(x6), .B0(mai_mai_n867_), .Y(mai_mai_n868_));
  NA3        m0819(.A(mai_mai_n868_), .B(mai_mai_n841_), .C(mai_mai_n831_), .Y(mai10));
  NO2        m0820(.A(x4), .B(x1), .Y(mai_mai_n870_));
  NO2        m0821(.A(mai_mai_n870_), .B(mai_mai_n139_), .Y(mai_mai_n871_));
  NA3        m0822(.A(x5), .B(x4), .C(x0), .Y(mai_mai_n872_));
  NOi21      m0823(.An(mai_mai_n234_), .B(mai_mai_n130_), .Y(mai_mai_n873_));
  NA2        m0824(.A(x4), .B(mai_mai_n105_), .Y(mai_mai_n874_));
  NO2        m0825(.A(mai_mai_n296_), .B(mai_mai_n874_), .Y(mai_mai_n875_));
  NA2        m0826(.A(mai_mai_n862_), .B(mai_mai_n50_), .Y(mai_mai_n876_));
  NA2        m0827(.A(mai_mai_n553_), .B(mai_mai_n247_), .Y(mai_mai_n877_));
  NO2        m0828(.A(mai_mai_n877_), .B(mai_mai_n876_), .Y(mai_mai_n878_));
  NA2        m0829(.A(mai_mai_n878_), .B(x7), .Y(mai_mai_n879_));
  NA2        m0830(.A(mai_mai_n55_), .B(mai_mai_n71_), .Y(mai_mai_n880_));
  AOI210     m0831(.A0(mai_mai_n411_), .A1(mai_mai_n328_), .B0(mai_mai_n874_), .Y(mai_mai_n881_));
  NA2        m0832(.A(mai_mai_n881_), .B(mai_mai_n880_), .Y(mai_mai_n882_));
  NO2        m0833(.A(mai_mai_n329_), .B(mai_mai_n133_), .Y(mai_mai_n883_));
  NA2        m0834(.A(mai_mai_n883_), .B(mai_mai_n395_), .Y(mai_mai_n884_));
  AOI210     m0835(.A0(mai_mai_n884_), .A1(mai_mai_n882_), .B0(x3), .Y(mai_mai_n885_));
  NA2        m0836(.A(mai_mai_n638_), .B(mai_mai_n227_), .Y(mai_mai_n886_));
  NO2        m0837(.A(x5), .B(mai_mai_n105_), .Y(mai_mai_n887_));
  OAI210     m0838(.A0(mai_mai_n887_), .A1(mai_mai_n216_), .B0(mai_mai_n845_), .Y(mai_mai_n888_));
  NA3        m0839(.A(mai_mai_n429_), .B(mai_mai_n123_), .C(mai_mai_n395_), .Y(mai_mai_n889_));
  OAI210     m0840(.A0(mai_mai_n413_), .A1(mai_mai_n196_), .B0(mai_mai_n889_), .Y(mai_mai_n890_));
  AOI210     m0841(.A0(mai_mai_n888_), .A1(mai_mai_n232_), .B0(mai_mai_n890_), .Y(mai_mai_n891_));
  OAI220     m0842(.A0(mai_mai_n891_), .A1(mai_mai_n59_), .B0(mai_mai_n886_), .B1(mai_mai_n651_), .Y(mai_mai_n892_));
  OAI210     m0843(.A0(mai_mai_n892_), .A1(mai_mai_n885_), .B0(mai_mai_n850_), .Y(mai_mai_n893_));
  NO2        m0844(.A(x4), .B(x3), .Y(mai_mai_n894_));
  NO3        m0845(.A(mai_mai_n894_), .B(mai_mai_n316_), .C(mai_mai_n87_), .Y(mai_mai_n895_));
  NA2        m0846(.A(mai_mai_n895_), .B(mai_mai_n402_), .Y(mai_mai_n896_));
  AOI210     m0847(.A0(mai_mai_n370_), .A1(mai_mai_n122_), .B0(mai_mai_n228_), .Y(mai_mai_n897_));
  NA2        m0848(.A(mai_mai_n870_), .B(mai_mai_n55_), .Y(mai_mai_n898_));
  NO2        m0849(.A(mai_mai_n898_), .B(mai_mai_n50_), .Y(mai_mai_n899_));
  NO3        m0850(.A(x4), .B(mai_mai_n105_), .C(mai_mai_n59_), .Y(mai_mai_n900_));
  NA2        m0851(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n901_));
  NO3        m0852(.A(mai_mai_n473_), .B(mai_mai_n901_), .C(x2), .Y(mai_mai_n902_));
  NO3        m0853(.A(mai_mai_n902_), .B(mai_mai_n899_), .C(mai_mai_n897_), .Y(mai_mai_n903_));
  AOI210     m0854(.A0(mai_mai_n903_), .A1(mai_mai_n896_), .B0(mai_mai_n190_), .Y(mai_mai_n904_));
  NO2        m0855(.A(mai_mai_n608_), .B(mai_mai_n459_), .Y(mai_mai_n905_));
  NO2        m0856(.A(x6), .B(x2), .Y(mai_mai_n906_));
  NO3        m0857(.A(mai_mai_n906_), .B(mai_mai_n638_), .C(mai_mai_n60_), .Y(mai_mai_n907_));
  OAI210     m0858(.A0(mai_mai_n907_), .A1(mai_mai_n905_), .B0(mai_mai_n246_), .Y(mai_mai_n908_));
  NO2        m0859(.A(mai_mai_n795_), .B(mai_mai_n411_), .Y(mai_mai_n909_));
  NA3        m0860(.A(x4), .B(x3), .C(mai_mai_n105_), .Y(mai_mai_n910_));
  NO3        m0861(.A(mai_mai_n910_), .B(mai_mai_n644_), .C(mai_mai_n429_), .Y(mai_mai_n911_));
  AOI210     m0862(.A0(mai_mai_n909_), .A1(mai_mai_n436_), .B0(mai_mai_n911_), .Y(mai_mai_n912_));
  AOI210     m0863(.A0(mai_mai_n912_), .A1(mai_mai_n908_), .B0(mai_mai_n422_), .Y(mai_mai_n913_));
  NO2        m0864(.A(mai_mai_n55_), .B(mai_mai_n56_), .Y(mai_mai_n914_));
  OAI220     m0865(.A0(mai_mai_n757_), .A1(mai_mai_n424_), .B0(mai_mai_n692_), .B1(mai_mai_n122_), .Y(mai_mai_n915_));
  NOi21      m0866(.An(mai_mai_n118_), .B(mai_mai_n117_), .Y(mai_mai_n916_));
  NO3        m0867(.A(mai_mai_n317_), .B(mai_mai_n296_), .C(mai_mai_n916_), .Y(mai_mai_n917_));
  AOI220     m0868(.A0(mai_mai_n917_), .A1(mai_mai_n231_), .B0(mai_mai_n915_), .B1(mai_mai_n111_), .Y(mai_mai_n918_));
  NO2        m0869(.A(mai_mai_n918_), .B(mai_mai_n914_), .Y(mai_mai_n919_));
  NA2        m0870(.A(mai_mai_n477_), .B(mai_mai_n236_), .Y(mai_mai_n920_));
  NO2        m0871(.A(mai_mai_n446_), .B(mai_mai_n537_), .Y(mai_mai_n921_));
  NA3        m0872(.A(mai_mai_n921_), .B(mai_mai_n920_), .C(mai_mai_n55_), .Y(mai_mai_n922_));
  NO2        m0873(.A(mai_mai_n172_), .B(mai_mai_n105_), .Y(mai_mai_n923_));
  INV        m0874(.A(mai_mai_n922_), .Y(mai_mai_n924_));
  NO4        m0875(.A(mai_mai_n924_), .B(mai_mai_n919_), .C(mai_mai_n913_), .D(mai_mai_n904_), .Y(mai_mai_n925_));
  NA3        m0876(.A(mai_mai_n925_), .B(mai_mai_n893_), .C(mai_mai_n879_), .Y(mai11));
  NA2        m0877(.A(mai_mai_n349_), .B(mai_mai_n92_), .Y(mai_mai_n927_));
  INV        m0878(.A(mai_mai_n812_), .Y(mai_mai_n928_));
  OAI220     m0879(.A0(mai_mai_n928_), .A1(mai_mai_n53_), .B0(mai_mai_n927_), .B1(mai_mai_n338_), .Y(mai_mai_n929_));
  NO2        m0880(.A(mai_mai_n707_), .B(x5), .Y(mai_mai_n930_));
  NO2        m0881(.A(mai_mai_n157_), .B(mai_mai_n489_), .Y(mai_mai_n931_));
  AOI220     m0882(.A0(mai_mai_n931_), .A1(mai_mai_n930_), .B0(mai_mai_n929_), .B1(x5), .Y(mai_mai_n932_));
  OAI220     m0883(.A0(mai_mai_n873_), .A1(mai_mai_n199_), .B0(mai_mai_n197_), .B1(mai_mai_n172_), .Y(mai_mai_n933_));
  NO2        m0884(.A(mai_mai_n313_), .B(mai_mai_n396_), .Y(mai_mai_n934_));
  AOI220     m0885(.A0(mai_mai_n934_), .A1(mai_mai_n170_), .B0(mai_mai_n933_), .B1(mai_mai_n153_), .Y(mai_mai_n935_));
  NO2        m0886(.A(mai_mai_n935_), .B(mai_mai_n413_), .Y(mai_mai_n936_));
  NO2        m0887(.A(mai_mai_n228_), .B(x2), .Y(mai_mai_n937_));
  OAI210     m0888(.A0(mai_mai_n832_), .A1(mai_mai_n937_), .B0(mai_mai_n387_), .Y(mai_mai_n938_));
  NO2        m0889(.A(mai_mai_n55_), .B(mai_mai_n103_), .Y(mai_mai_n939_));
  NA2        m0890(.A(mai_mai_n253_), .B(mai_mai_n939_), .Y(mai_mai_n940_));
  NO2        m0891(.A(mai_mai_n71_), .B(x1), .Y(mai_mai_n941_));
  NA2        m0892(.A(mai_mai_n941_), .B(mai_mai_n78_), .Y(mai_mai_n942_));
  OA220      m0893(.A0(mai_mai_n942_), .A1(mai_mai_n561_), .B0(mai_mai_n940_), .B1(mai_mai_n489_), .Y(mai_mai_n943_));
  AOI210     m0894(.A0(mai_mai_n943_), .A1(mai_mai_n938_), .B0(mai_mai_n651_), .Y(mai_mai_n944_));
  NO2        m0895(.A(mai_mai_n276_), .B(mai_mai_n53_), .Y(mai_mai_n945_));
  NO2        m0896(.A(mai_mai_n402_), .B(x3), .Y(mai_mai_n946_));
  NA3        m0897(.A(mai_mai_n946_), .B(mai_mai_n945_), .C(mai_mai_n811_), .Y(mai_mai_n947_));
  AOI210     m0898(.A0(mai_mai_n947_), .A1(mai_mai_n848_), .B0(mai_mai_n368_), .Y(mai_mai_n948_));
  NA2        m0899(.A(mai_mai_n105_), .B(x1), .Y(mai_mai_n949_));
  NO2        m0900(.A(mai_mai_n566_), .B(mai_mai_n202_), .Y(mai_mai_n950_));
  NA4        m0901(.A(mai_mai_n950_), .B(mai_mai_n807_), .C(mai_mai_n433_), .D(mai_mai_n949_), .Y(mai_mai_n951_));
  NA3        m0902(.A(x6), .B(x5), .C(mai_mai_n105_), .Y(mai_mai_n952_));
  NO2        m0903(.A(mai_mai_n952_), .B(mai_mai_n251_), .Y(mai_mai_n953_));
  NO2        m0904(.A(mai_mai_n413_), .B(x0), .Y(mai_mai_n954_));
  NOi31      m0905(.An(mai_mai_n954_), .B(mai_mai_n162_), .C(mai_mai_n51_), .Y(mai_mai_n955_));
  AOI210     m0906(.A0(mai_mai_n953_), .A1(mai_mai_n168_), .B0(mai_mai_n955_), .Y(mai_mai_n956_));
  NA2        m0907(.A(mai_mai_n956_), .B(mai_mai_n951_), .Y(mai_mai_n957_));
  NO4        m0908(.A(mai_mai_n957_), .B(mai_mai_n948_), .C(mai_mai_n944_), .D(mai_mai_n936_), .Y(mai_mai_n958_));
  OAI210     m0909(.A0(mai_mai_n932_), .A1(mai_mai_n134_), .B0(mai_mai_n958_), .Y(mai_mai_n959_));
  NA2        m0910(.A(mai_mai_n786_), .B(mai_mai_n87_), .Y(mai_mai_n960_));
  NA2        m0911(.A(mai_mai_n960_), .B(mai_mai_n99_), .Y(mai_mai_n961_));
  NO2        m0912(.A(x8), .B(x1), .Y(mai_mai_n962_));
  NO2        m0913(.A(mai_mai_n630_), .B(mai_mai_n414_), .Y(mai_mai_n963_));
  NA2        m0914(.A(mai_mai_n53_), .B(mai_mai_n963_), .Y(mai_mai_n964_));
  OAI210     m0915(.A0(mai_mai_n961_), .A1(x3), .B0(mai_mai_n964_), .Y(mai_mai_n965_));
  NO2        m0916(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n966_));
  OAI210     m0917(.A0(mai_mai_n966_), .A1(x2), .B0(mai_mai_n212_), .Y(mai_mai_n967_));
  NO3        m0918(.A(mai_mai_n55_), .B(x6), .C(x1), .Y(mai_mai_n968_));
  NOi21      m0919(.An(mai_mai_n968_), .B(mai_mai_n446_), .Y(mai_mai_n969_));
  AOI210     m0920(.A0(mai_mai_n965_), .A1(x2), .B0(mai_mai_n969_), .Y(mai_mai_n970_));
  NO2        m0921(.A(mai_mai_n210_), .B(x2), .Y(mai_mai_n971_));
  NOi21      m0922(.An(mai_mai_n361_), .B(mai_mai_n519_), .Y(mai_mai_n972_));
  NA2        m0923(.A(x8), .B(mai_mai_n105_), .Y(mai_mai_n973_));
  NO2        m0924(.A(mai_mai_n103_), .B(x1), .Y(mai_mai_n974_));
  NA2        m0925(.A(mai_mai_n84_), .B(mai_mai_n71_), .Y(mai_mai_n975_));
  NO2        m0926(.A(mai_mai_n970_), .B(mai_mai_n774_), .Y(mai_mai_n976_));
  AO210      m0927(.A0(mai_mai_n959_), .A1(mai_mai_n57_), .B0(mai_mai_n976_), .Y(mai12));
  NA2        m0928(.A(mai_mai_n806_), .B(mai_mai_n226_), .Y(mai_mai_n978_));
  NO2        m0929(.A(mai_mai_n570_), .B(x7), .Y(mai_mai_n979_));
  NA2        m0930(.A(mai_mai_n979_), .B(mai_mai_n252_), .Y(mai_mai_n980_));
  INV        m0931(.A(mai_mai_n795_), .Y(mai_mai_n981_));
  AOI210     m0932(.A0(mai_mai_n980_), .A1(mai_mai_n978_), .B0(mai_mai_n981_), .Y(mai_mai_n982_));
  NOi21      m0933(.An(mai_mai_n375_), .B(mai_mai_n509_), .Y(mai_mai_n983_));
  NO2        m0934(.A(x7), .B(mai_mai_n50_), .Y(mai_mai_n984_));
  NO3        m0935(.A(mai_mai_n788_), .B(mai_mai_n107_), .C(mai_mai_n98_), .Y(mai_mai_n985_));
  INV        m0936(.A(mai_mai_n985_), .Y(mai_mai_n986_));
  NA2        m0937(.A(mai_mai_n939_), .B(mai_mai_n56_), .Y(mai_mai_n987_));
  NO2        m0938(.A(mai_mai_n986_), .B(mai_mai_n983_), .Y(mai_mai_n988_));
  OAI210     m0939(.A0(mai_mai_n988_), .A1(mai_mai_n982_), .B0(mai_mai_n532_), .Y(mai_mai_n989_));
  NA2        m0940(.A(mai_mai_n87_), .B(x5), .Y(mai_mai_n990_));
  OAI210     m0941(.A0(mai_mai_n990_), .A1(mai_mai_n296_), .B0(mai_mai_n662_), .Y(mai_mai_n991_));
  AOI210     m0942(.A0(mai_mai_n758_), .A1(mai_mai_n113_), .B0(mai_mai_n991_), .Y(mai_mai_n992_));
  NO2        m0943(.A(mai_mai_n992_), .B(mai_mai_n64_), .Y(mai_mai_n993_));
  NO2        m0944(.A(mai_mai_n608_), .B(mai_mai_n293_), .Y(mai_mai_n994_));
  NO2        m0945(.A(mai_mai_n692_), .B(x3), .Y(mai_mai_n995_));
  NO2        m0946(.A(mai_mai_n606_), .B(x8), .Y(mai_mai_n996_));
  NA2        m0947(.A(mai_mai_n996_), .B(mai_mai_n995_), .Y(mai_mai_n997_));
  AOI210     m0948(.A0(mai_mai_n630_), .A1(mai_mai_n226_), .B0(x7), .Y(mai_mai_n998_));
  NO2        m0949(.A(mai_mai_n998_), .B(x8), .Y(mai_mai_n999_));
  NA4        m0950(.A(mai_mai_n610_), .B(mai_mai_n602_), .C(mai_mai_n187_), .D(x0), .Y(mai_mai_n1000_));
  OAI220     m0951(.A0(mai_mai_n1000_), .A1(mai_mai_n999_), .B0(mai_mai_n997_), .B1(mai_mai_n528_), .Y(mai_mai_n1001_));
  AOI210     m0952(.A0(mai_mai_n993_), .A1(mai_mai_n906_), .B0(mai_mai_n1001_), .Y(mai_mai_n1002_));
  NO2        m0953(.A(mai_mai_n226_), .B(mai_mai_n55_), .Y(mai_mai_n1003_));
  NO2        m0954(.A(mai_mai_n231_), .B(x8), .Y(mai_mai_n1004_));
  NOi32      m0955(.An(mai_mai_n1004_), .Bn(mai_mai_n186_), .C(mai_mai_n520_), .Y(mai_mai_n1005_));
  INV        m0956(.A(mai_mai_n60_), .Y(mai_mai_n1006_));
  OAI210     m0957(.A0(mai_mai_n1005_), .A1(mai_mai_n1003_), .B0(mai_mai_n1006_), .Y(mai_mai_n1007_));
  NO2        m0958(.A(x7), .B(x0), .Y(mai_mai_n1008_));
  NO3        m0959(.A(mai_mai_n147_), .B(mai_mai_n1008_), .C(mai_mai_n136_), .Y(mai_mai_n1009_));
  XN2        m0960(.A(x8), .B(x7), .Y(mai_mai_n1010_));
  NO2        m0961(.A(mai_mai_n234_), .B(mai_mai_n1010_), .Y(mai_mai_n1011_));
  OAI210     m0962(.A0(mai_mai_n1011_), .A1(mai_mai_n1009_), .B0(mai_mai_n674_), .Y(mai_mai_n1012_));
  NO2        m0963(.A(mai_mai_n243_), .B(mai_mai_n239_), .Y(mai_mai_n1013_));
  NO2        m0964(.A(mai_mai_n103_), .B(x4), .Y(mai_mai_n1014_));
  OAI210     m0965(.A0(mai_mai_n1013_), .A1(mai_mai_n252_), .B0(mai_mai_n1014_), .Y(mai_mai_n1015_));
  NA3        m0966(.A(mai_mai_n1015_), .B(mai_mai_n1012_), .C(mai_mai_n1007_), .Y(mai_mai_n1016_));
  NA2        m0967(.A(mai_mai_n1016_), .B(mai_mai_n513_), .Y(mai_mai_n1017_));
  NO2        m0968(.A(mai_mai_n55_), .B(x4), .Y(mai_mai_n1018_));
  NA2        m0969(.A(mai_mai_n1018_), .B(mai_mai_n152_), .Y(mai_mai_n1019_));
  NA2        m0970(.A(mai_mai_n909_), .B(mai_mai_n50_), .Y(mai_mai_n1020_));
  AOI210     m0971(.A0(mai_mai_n1020_), .A1(mai_mai_n1019_), .B0(mai_mai_n398_), .Y(mai_mai_n1021_));
  NA3        m0972(.A(x3), .B(mai_mai_n619_), .C(x1), .Y(mai_mai_n1022_));
  OAI210     m0973(.A0(x8), .A1(x0), .B0(x4), .Y(mai_mai_n1023_));
  NO2        m0974(.A(x7), .B(mai_mai_n56_), .Y(mai_mai_n1024_));
  NO2        m0975(.A(mai_mai_n68_), .B(mai_mai_n1024_), .Y(mai_mai_n1025_));
  NOi21      m0976(.An(mai_mai_n1023_), .B(mai_mai_n1025_), .Y(mai_mai_n1026_));
  NO2        m0977(.A(mai_mai_n610_), .B(mai_mai_n296_), .Y(mai_mai_n1027_));
  NO2        m0978(.A(mai_mai_n715_), .B(mai_mai_n203_), .Y(mai_mai_n1028_));
  OAI210     m0979(.A0(mai_mai_n1027_), .A1(mai_mai_n1026_), .B0(mai_mai_n1028_), .Y(mai_mai_n1029_));
  NO2        m0980(.A(mai_mai_n134_), .B(mai_mai_n133_), .Y(mai_mai_n1030_));
  NO2        m0981(.A(mai_mai_n554_), .B(mai_mai_n411_), .Y(mai_mai_n1031_));
  OAI210     m0982(.A0(mai_mai_n1031_), .A1(mai_mai_n1030_), .B0(mai_mai_n231_), .Y(mai_mai_n1032_));
  NO2        m0983(.A(mai_mai_n755_), .B(mai_mai_n393_), .Y(mai_mai_n1033_));
  NA2        m0984(.A(mai_mai_n301_), .B(mai_mai_n59_), .Y(mai_mai_n1034_));
  NO2        m0985(.A(mai_mai_n987_), .B(mai_mai_n1034_), .Y(mai_mai_n1035_));
  AOI210     m0986(.A0(mai_mai_n1033_), .A1(mai_mai_n168_), .B0(mai_mai_n1035_), .Y(mai_mai_n1036_));
  NA4        m0987(.A(mai_mai_n1036_), .B(mai_mai_n1032_), .C(mai_mai_n1029_), .D(mai_mai_n1022_), .Y(mai_mai_n1037_));
  OAI210     m0988(.A0(mai_mai_n1037_), .A1(mai_mai_n1021_), .B0(mai_mai_n620_), .Y(mai_mai_n1038_));
  NA4        m0989(.A(mai_mai_n1038_), .B(mai_mai_n1017_), .C(mai_mai_n1002_), .D(mai_mai_n989_), .Y(mai13));
  NO2        m0990(.A(mai_mai_n429_), .B(mai_mai_n323_), .Y(mai_mai_n1040_));
  NOi41      m0991(.An(mai_mai_n1040_), .B(mai_mai_n619_), .C(mai_mai_n265_), .D(mai_mai_n218_), .Y(mai_mai_n1041_));
  NO2        m0992(.A(mai_mai_n788_), .B(mai_mai_n172_), .Y(mai_mai_n1042_));
  NA2        m0993(.A(mai_mai_n1041_), .B(x3), .Y(mai_mai_n1043_));
  NO2        m0994(.A(mai_mai_n788_), .B(x6), .Y(mai_mai_n1044_));
  NO3        m0995(.A(x8), .B(x5), .C(mai_mai_n105_), .Y(mai_mai_n1045_));
  NA2        m0996(.A(mai_mai_n1045_), .B(mai_mai_n585_), .Y(mai_mai_n1046_));
  NO2        m0997(.A(mai_mai_n554_), .B(mai_mai_n184_), .Y(mai_mai_n1047_));
  NA2        m0998(.A(mai_mai_n1047_), .B(mai_mai_n968_), .Y(mai_mai_n1048_));
  NA2        m0999(.A(mai_mai_n414_), .B(mai_mai_n53_), .Y(mai_mai_n1049_));
  NO2        m1000(.A(mai_mai_n1049_), .B(mai_mai_n845_), .Y(mai_mai_n1050_));
  NA2        m1001(.A(mai_mai_n987_), .B(mai_mai_n434_), .Y(mai_mai_n1051_));
  NA2        m1002(.A(mai_mai_n56_), .B(mai_mai_n105_), .Y(mai_mai_n1052_));
  NA2        m1003(.A(mai_mai_n1052_), .B(x1), .Y(mai_mai_n1053_));
  NO2        m1004(.A(mai_mai_n1053_), .B(mai_mai_n236_), .Y(mai_mai_n1054_));
  NA2        m1005(.A(mai_mai_n1054_), .B(mai_mai_n1051_), .Y(mai_mai_n1055_));
  NAi41      m1006(.An(mai_mai_n1050_), .B(mai_mai_n1055_), .C(mai_mai_n1048_), .D(mai_mai_n1046_), .Y(mai_mai_n1056_));
  NA2        m1007(.A(mai_mai_n1056_), .B(mai_mai_n68_), .Y(mai_mai_n1057_));
  NA2        m1008(.A(mai_mai_n71_), .B(x3), .Y(mai_mai_n1058_));
  NA2        m1009(.A(mai_mai_n1058_), .B(mai_mai_n816_), .Y(mai_mai_n1059_));
  OAI220     m1010(.A0(mai_mai_n275_), .A1(mai_mai_n755_), .B0(mai_mai_n87_), .B1(mai_mai_n77_), .Y(mai_mai_n1060_));
  AOI210     m1011(.A0(mai_mai_n990_), .A1(mai_mai_n564_), .B0(mai_mai_n874_), .Y(mai_mai_n1061_));
  OA210      m1012(.A0(mai_mai_n1060_), .A1(mai_mai_n1059_), .B0(mai_mai_n1061_), .Y(mai_mai_n1062_));
  NA2        m1013(.A(mai_mai_n566_), .B(mai_mai_n55_), .Y(mai_mai_n1063_));
  NA2        m1014(.A(x6), .B(mai_mai_n50_), .Y(mai_mai_n1064_));
  NA2        m1015(.A(mai_mai_n1064_), .B(mai_mai_n498_), .Y(mai_mai_n1065_));
  NO2        m1016(.A(mai_mai_n149_), .B(mai_mai_n123_), .Y(mai_mai_n1066_));
  AOI210     m1017(.A0(mai_mai_n1065_), .A1(mai_mai_n399_), .B0(mai_mai_n1066_), .Y(mai_mai_n1067_));
  NO2        m1018(.A(mai_mai_n1067_), .B(mai_mai_n795_), .Y(mai_mai_n1068_));
  OAI210     m1019(.A0(mai_mai_n1068_), .A1(mai_mai_n1062_), .B0(mai_mai_n1008_), .Y(mai_mai_n1069_));
  NAi21      m1020(.An(mai_mai_n84_), .B(mai_mai_n356_), .Y(mai_mai_n1070_));
  NO2        m1021(.A(x4), .B(x0), .Y(mai_mai_n1071_));
  NA2        m1022(.A(mai_mai_n227_), .B(mai_mai_n674_), .Y(mai_mai_n1072_));
  NA2        m1023(.A(mai_mai_n56_), .B(x0), .Y(mai_mai_n1073_));
  NO2        m1024(.A(mai_mai_n296_), .B(mai_mai_n356_), .Y(mai_mai_n1074_));
  OAI210     m1025(.A0(mai_mai_n56_), .A1(mai_mai_n1074_), .B0(mai_mai_n305_), .Y(mai_mai_n1075_));
  NO2        m1026(.A(mai_mai_n726_), .B(x1), .Y(mai_mai_n1076_));
  NA2        m1027(.A(mai_mai_n459_), .B(mai_mai_n50_), .Y(mai_mai_n1077_));
  AOI220     m1028(.A0(mai_mai_n1077_), .A1(mai_mai_n1042_), .B0(mai_mai_n875_), .B1(mai_mai_n99_), .Y(mai_mai_n1078_));
  NA2        m1029(.A(mai_mai_n1078_), .B(mai_mai_n1075_), .Y(mai_mai_n1079_));
  AOI220     m1030(.A0(mai_mai_n1079_), .A1(mai_mai_n124_), .B0(mai_mai_n1014_), .B1(mai_mai_n67_), .Y(mai_mai_n1080_));
  NA4        m1031(.A(mai_mai_n1080_), .B(mai_mai_n1069_), .C(mai_mai_n1057_), .D(mai_mai_n1043_), .Y(mai14));
  NO2        m1032(.A(mai_mai_n344_), .B(mai_mai_n71_), .Y(mai_mai_n1082_));
  NO3        m1033(.A(x7), .B(x6), .C(x0), .Y(mai_mai_n1083_));
  OAI210     m1034(.A0(mai_mai_n1083_), .A1(mai_mai_n1082_), .B0(x8), .Y(mai_mai_n1084_));
  NA2        m1035(.A(mai_mai_n996_), .B(mai_mai_n85_), .Y(mai_mai_n1085_));
  AOI210     m1036(.A0(mai_mai_n1085_), .A1(mai_mai_n1084_), .B0(mai_mai_n145_), .Y(mai_mai_n1086_));
  AOI210     m1037(.A0(mai_mai_n348_), .A1(mai_mai_n774_), .B0(mai_mai_n414_), .Y(mai_mai_n1087_));
  NA2        m1038(.A(mai_mai_n253_), .B(mai_mai_n873_), .Y(mai_mai_n1088_));
  OAI220     m1039(.A0(mai_mai_n1088_), .A1(mai_mai_n1087_), .B0(mai_mai_n432_), .B1(mai_mai_n740_), .Y(mai_mai_n1089_));
  OA210      m1040(.A0(mai_mai_n1089_), .A1(mai_mai_n1086_), .B0(x4), .Y(mai_mai_n1090_));
  NA2        m1041(.A(x6), .B(x2), .Y(mai_mai_n1091_));
  NO4        m1042(.A(mai_mai_n554_), .B(mai_mai_n349_), .C(mai_mai_n272_), .D(mai_mai_n111_), .Y(mai_mai_n1092_));
  NA2        m1043(.A(mai_mai_n1092_), .B(mai_mai_n59_), .Y(mai_mai_n1093_));
  NA2        m1044(.A(x6), .B(mai_mai_n103_), .Y(mai_mai_n1094_));
  AOI210     m1045(.A0(mai_mai_n996_), .A1(mai_mai_n900_), .B0(x1), .Y(mai_mai_n1095_));
  NO2        m1046(.A(mai_mai_n493_), .B(x5), .Y(mai_mai_n1096_));
  NA3        m1047(.A(mai_mai_n1096_), .B(mai_mai_n117_), .C(x0), .Y(mai_mai_n1097_));
  NA4        m1048(.A(mai_mai_n637_), .B(mai_mai_n840_), .C(mai_mai_n275_), .D(mai_mai_n68_), .Y(mai_mai_n1098_));
  AN3        m1049(.A(mai_mai_n1098_), .B(mai_mai_n1097_), .C(mai_mai_n1095_), .Y(mai_mai_n1099_));
  NO2        m1050(.A(mai_mai_n644_), .B(mai_mai_n973_), .Y(mai_mai_n1100_));
  NO2        m1051(.A(mai_mai_n77_), .B(mai_mai_n58_), .Y(mai_mai_n1101_));
  OAI210     m1052(.A0(mai_mai_n1100_), .A1(mai_mai_n412_), .B0(mai_mai_n1101_), .Y(mai_mai_n1102_));
  AO210      m1053(.A0(mai_mai_n1082_), .A1(mai_mai_n900_), .B0(mai_mai_n53_), .Y(mai_mai_n1103_));
  AOI210     m1054(.A0(mai_mai_n703_), .A1(mai_mai_n749_), .B0(mai_mai_n1103_), .Y(mai_mai_n1104_));
  AOI220     m1055(.A0(mai_mai_n1104_), .A1(mai_mai_n1102_), .B0(mai_mai_n1099_), .B1(mai_mai_n1093_), .Y(mai_mai_n1105_));
  NO2        m1056(.A(mai_mai_n1105_), .B(mai_mai_n1090_), .Y(mai_mai_n1106_));
  NO2        m1057(.A(mai_mai_n293_), .B(x2), .Y(mai_mai_n1107_));
  XN2        m1058(.A(x4), .B(x1), .Y(mai_mai_n1108_));
  NO2        m1059(.A(mai_mai_n1108_), .B(mai_mai_n275_), .Y(mai_mai_n1109_));
  NO2        m1060(.A(mai_mai_n312_), .B(mai_mai_n60_), .Y(mai_mai_n1110_));
  NA2        m1061(.A(mai_mai_n631_), .B(mai_mai_n56_), .Y(mai_mai_n1111_));
  OAI220     m1062(.A0(mai_mai_n1111_), .A1(mai_mai_n146_), .B0(mai_mai_n176_), .B1(mai_mai_n71_), .Y(mai_mai_n1112_));
  NO2        m1063(.A(mai_mai_n199_), .B(mai_mai_n234_), .Y(mai_mai_n1113_));
  NA2        m1064(.A(mai_mai_n227_), .B(mai_mai_n327_), .Y(mai_mai_n1114_));
  NA2        m1065(.A(mai_mai_n584_), .B(mai_mai_n916_), .Y(mai_mai_n1115_));
  NO2        m1066(.A(mai_mai_n1115_), .B(mai_mai_n1114_), .Y(mai_mai_n1116_));
  AOI210     m1067(.A0(mai_mai_n1113_), .A1(mai_mai_n1112_), .B0(mai_mai_n1116_), .Y(mai_mai_n1117_));
  NO2        m1068(.A(mai_mai_n1117_), .B(x7), .Y(mai_mai_n1118_));
  NO2        m1069(.A(mai_mai_n453_), .B(x6), .Y(mai_mai_n1119_));
  NO3        m1070(.A(mai_mai_n692_), .B(mai_mai_n459_), .C(mai_mai_n54_), .Y(mai_mai_n1120_));
  INV        m1071(.A(mai_mai_n1120_), .Y(mai_mai_n1121_));
  NO2        m1072(.A(mai_mai_n1121_), .B(mai_mai_n277_), .Y(mai_mai_n1122_));
  NA2        m1073(.A(mai_mai_n814_), .B(mai_mai_n53_), .Y(mai_mai_n1123_));
  OAI210     m1074(.A0(mai_mai_n224_), .A1(mai_mai_n113_), .B0(x2), .Y(mai_mai_n1124_));
  OA220      m1075(.A0(x4), .A1(mai_mai_n1124_), .B0(mai_mai_n1123_), .B1(mai_mai_n348_), .Y(mai_mai_n1125_));
  NA3        m1076(.A(mai_mai_n921_), .B(mai_mai_n679_), .C(mai_mai_n55_), .Y(mai_mai_n1126_));
  NA2        m1077(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n1127_));
  NO2        m1078(.A(mai_mai_n1127_), .B(mai_mai_n183_), .Y(mai_mai_n1128_));
  NA4        m1079(.A(mai_mai_n1128_), .B(mai_mai_n340_), .C(mai_mai_n234_), .D(mai_mai_n67_), .Y(mai_mai_n1129_));
  NA3        m1080(.A(mai_mai_n1076_), .B(mai_mai_n566_), .C(mai_mai_n576_), .Y(mai_mai_n1130_));
  AN3        m1081(.A(mai_mai_n1130_), .B(mai_mai_n1129_), .C(mai_mai_n1126_), .Y(mai_mai_n1131_));
  OAI210     m1082(.A0(mai_mai_n1125_), .A1(mai_mai_n288_), .B0(mai_mai_n1131_), .Y(mai_mai_n1132_));
  NO3        m1083(.A(mai_mai_n1132_), .B(mai_mai_n1122_), .C(mai_mai_n1118_), .Y(mai_mai_n1133_));
  OAI210     m1084(.A0(mai_mai_n1106_), .A1(x3), .B0(mai_mai_n1133_), .Y(mai15));
  NA2        m1085(.A(mai_mai_n538_), .B(mai_mai_n59_), .Y(mai_mai_n1135_));
  INV        m1086(.A(mai_mai_n1135_), .Y(mai_mai_n1136_));
  NA3        m1087(.A(mai_mai_n57_), .B(x6), .C(mai_mai_n105_), .Y(mai_mai_n1137_));
  NO2        m1088(.A(mai_mai_n1137_), .B(mai_mai_n268_), .Y(mai_mai_n1138_));
  OAI210     m1089(.A0(mai_mai_n1138_), .A1(mai_mai_n1136_), .B0(mai_mai_n1014_), .Y(mai_mai_n1139_));
  NA2        m1090(.A(mai_mai_n107_), .B(mai_mai_n105_), .Y(mai_mai_n1140_));
  NA4        m1091(.A(mai_mai_n1140_), .B(mai_mai_n582_), .C(mai_mai_n281_), .D(x6), .Y(mai_mai_n1141_));
  INV        m1092(.A(x3), .Y(mai_mai_n1142_));
  NA3        m1093(.A(mai_mai_n1142_), .B(mai_mai_n1141_), .C(mai_mai_n1139_), .Y(mai_mai_n1143_));
  NO2        m1094(.A(mai_mai_n268_), .B(mai_mai_n105_), .Y(mai_mai_n1144_));
  NO2        m1095(.A(mai_mai_n216_), .B(x5), .Y(mai_mai_n1145_));
  NA2        m1096(.A(mai_mai_n1145_), .B(mai_mai_n1144_), .Y(mai_mai_n1146_));
  NA3        m1097(.A(mai_mai_n1076_), .B(mai_mai_n572_), .C(mai_mai_n1024_), .Y(mai_mai_n1147_));
  NA4        m1098(.A(mai_mai_n1147_), .B(mai_mai_n1146_), .C(x3), .D(mai_mai_n1097_), .Y(mai_mai_n1148_));
  NA2        m1099(.A(mai_mai_n306_), .B(mai_mai_n315_), .Y(mai_mai_n1149_));
  AOI210     m1100(.A0(mai_mai_n1053_), .A1(mai_mai_n58_), .B0(mai_mai_n1149_), .Y(mai_mai_n1150_));
  NA3        m1101(.A(mai_mai_n643_), .B(x7), .C(mai_mai_n356_), .Y(mai_mai_n1151_));
  NO2        m1102(.A(mai_mai_n692_), .B(mai_mai_n53_), .Y(mai_mai_n1152_));
  NA2        m1103(.A(x3), .B(mai_mai_n1152_), .Y(mai_mai_n1153_));
  NA2        m1104(.A(mai_mai_n1153_), .B(mai_mai_n1151_), .Y(mai_mai_n1154_));
  OAI210     m1105(.A0(mai_mai_n1154_), .A1(mai_mai_n1150_), .B0(mai_mai_n77_), .Y(mai_mai_n1155_));
  NA2        m1106(.A(mai_mai_n342_), .B(mai_mai_n646_), .Y(mai_mai_n1156_));
  NA2        m1107(.A(mai_mai_n525_), .B(mai_mai_n56_), .Y(mai_mai_n1157_));
  NA3        m1108(.A(mai_mai_n1157_), .B(mai_mai_n315_), .C(mai_mai_n107_), .Y(mai_mai_n1158_));
  AOI210     m1109(.A0(mai_mai_n1158_), .A1(mai_mai_n1156_), .B0(mai_mai_n459_), .Y(mai_mai_n1159_));
  NO3        m1110(.A(mai_mai_n738_), .B(mai_mai_n571_), .C(mai_mai_n184_), .Y(mai_mai_n1160_));
  OAI210     m1111(.A0(mai_mai_n1160_), .A1(mai_mai_n1159_), .B0(mai_mai_n453_), .Y(mai_mai_n1161_));
  NO2        m1112(.A(mai_mai_n226_), .B(mai_mai_n64_), .Y(mai_mai_n1162_));
  AN2        m1113(.A(mai_mai_n1162_), .B(mai_mai_n382_), .Y(mai_mai_n1163_));
  NA2        m1114(.A(mai_mai_n57_), .B(x3), .Y(mai_mai_n1164_));
  NO2        m1115(.A(mai_mai_n50_), .B(mai_mai_n625_), .Y(mai_mai_n1165_));
  OAI210     m1116(.A0(mai_mai_n1165_), .A1(mai_mai_n1163_), .B0(mai_mai_n906_), .Y(mai_mai_n1166_));
  NA2        m1117(.A(mai_mai_n1128_), .B(mai_mai_n68_), .Y(mai_mai_n1167_));
  AOI210     m1118(.A0(x2), .A1(mai_mai_n555_), .B0(x8), .Y(mai_mai_n1168_));
  NO2        m1119(.A(mai_mai_n874_), .B(x6), .Y(mai_mai_n1169_));
  AN2        m1120(.A(mai_mai_n1168_), .B(mai_mai_n1167_), .Y(mai_mai_n1170_));
  NA4        m1121(.A(mai_mai_n1170_), .B(mai_mai_n1166_), .C(mai_mai_n1161_), .D(mai_mai_n1155_), .Y(mai_mai_n1171_));
  NA2        m1122(.A(mai_mai_n153_), .B(mai_mai_n679_), .Y(mai_mai_n1172_));
  NO2        m1123(.A(mai_mai_n593_), .B(x2), .Y(mai_mai_n1173_));
  NA2        m1124(.A(mai_mai_n1173_), .B(x1), .Y(mai_mai_n1174_));
  AOI210     m1125(.A0(mai_mai_n1174_), .A1(mai_mai_n1172_), .B0(mai_mai_n293_), .Y(mai_mai_n1175_));
  NO3        m1126(.A(mai_mai_n1137_), .B(mai_mai_n242_), .C(mai_mai_n226_), .Y(mai_mai_n1176_));
  NA3        m1127(.A(mai_mai_n57_), .B(x1), .C(x0), .Y(mai_mai_n1177_));
  NA3        m1128(.A(mai_mai_n71_), .B(x5), .C(x2), .Y(mai_mai_n1178_));
  NO2        m1129(.A(mai_mai_n1178_), .B(mai_mai_n1177_), .Y(mai_mai_n1179_));
  NO2        m1130(.A(mai_mai_n1179_), .B(mai_mai_n1176_), .Y(mai_mai_n1180_));
  NAi21      m1131(.An(mai_mai_n111_), .B(mai_mai_n687_), .Y(mai_mai_n1181_));
  OAI220     m1132(.A0(mai_mai_n296_), .A1(x7), .B0(mai_mai_n123_), .B1(mai_mai_n71_), .Y(mai_mai_n1182_));
  NA3        m1133(.A(mai_mai_n1182_), .B(mai_mai_n726_), .C(mai_mai_n974_), .Y(mai_mai_n1183_));
  NA2        m1134(.A(mai_mai_n82_), .B(mai_mai_n50_), .Y(mai_mai_n1184_));
  AO210      m1135(.A0(mai_mai_n1184_), .A1(mai_mai_n286_), .B0(mai_mai_n145_), .Y(mai_mai_n1185_));
  NA3        m1136(.A(mai_mai_n1185_), .B(mai_mai_n1183_), .C(mai_mai_n1180_), .Y(mai_mai_n1186_));
  OAI210     m1137(.A0(mai_mai_n1186_), .A1(mai_mai_n1175_), .B0(mai_mai_n56_), .Y(mai_mai_n1187_));
  NA2        m1138(.A(mai_mai_n633_), .B(x4), .Y(mai_mai_n1188_));
  OAI220     m1139(.A0(mai_mai_n1188_), .A1(mai_mai_n273_), .B0(mai_mai_n910_), .B1(mai_mai_n851_), .Y(mai_mai_n1189_));
  NA2        m1140(.A(x3), .B(mai_mai_n379_), .Y(mai_mai_n1190_));
  NA2        m1141(.A(mai_mai_n1162_), .B(mai_mai_n264_), .Y(mai_mai_n1191_));
  OAI210     m1142(.A0(mai_mai_n1190_), .A1(mai_mai_n769_), .B0(mai_mai_n1191_), .Y(mai_mai_n1192_));
  OAI210     m1143(.A0(mai_mai_n1192_), .A1(mai_mai_n1189_), .B0(x6), .Y(mai_mai_n1193_));
  NO2        m1144(.A(x7), .B(x5), .Y(mai_mai_n1194_));
  NA2        m1145(.A(mai_mai_n497_), .B(mai_mai_n1194_), .Y(mai_mai_n1195_));
  NA2        m1146(.A(mai_mai_n700_), .B(mai_mai_n264_), .Y(mai_mai_n1196_));
  NA3        m1147(.A(mai_mai_n566_), .B(mai_mai_n266_), .C(mai_mai_n221_), .Y(mai_mai_n1197_));
  NA2        m1148(.A(mai_mai_n1197_), .B(mai_mai_n1195_), .Y(mai_mai_n1198_));
  NA2        m1149(.A(mai_mai_n1198_), .B(mai_mai_n395_), .Y(mai_mai_n1199_));
  AOI210     m1150(.A0(mai_mai_n352_), .A1(mai_mai_n313_), .B0(mai_mai_n55_), .Y(mai_mai_n1200_));
  NA4        m1151(.A(mai_mai_n1200_), .B(mai_mai_n1199_), .C(mai_mai_n1193_), .D(mai_mai_n1187_), .Y(mai_mai_n1201_));
  AO220      m1152(.A0(mai_mai_n1201_), .A1(mai_mai_n1171_), .B0(mai_mai_n1148_), .B1(mai_mai_n1143_), .Y(mai16));
  NO2        m1153(.A(x4), .B(mai_mai_n59_), .Y(mai_mai_n1203_));
  NA2        m1154(.A(mai_mai_n607_), .B(mai_mai_n494_), .Y(mai_mai_n1204_));
  INV        m1155(.A(mai_mai_n1204_), .Y(mai_mai_n1205_));
  NO3        m1156(.A(x8), .B(x6), .C(mai_mai_n50_), .Y(mai_mai_n1206_));
  NO2        m1157(.A(mai_mai_n149_), .B(x5), .Y(mai_mai_n1207_));
  NA2        m1158(.A(mai_mai_n1207_), .B(mai_mai_n1173_), .Y(mai_mai_n1208_));
  NA2        m1159(.A(mai_mai_n532_), .B(mai_mai_n496_), .Y(mai_mai_n1209_));
  NA2        m1160(.A(mai_mai_n1209_), .B(mai_mai_n1208_), .Y(mai_mai_n1210_));
  OAI210     m1161(.A0(mai_mai_n1210_), .A1(mai_mai_n1205_), .B0(mai_mai_n1203_), .Y(mai_mai_n1211_));
  NO2        m1162(.A(mai_mai_n293_), .B(x7), .Y(mai_mai_n1212_));
  NA2        m1163(.A(mai_mai_n1212_), .B(x0), .Y(mai_mai_n1213_));
  NO2        m1164(.A(mai_mai_n1213_), .B(mai_mai_n583_), .Y(mai_mai_n1214_));
  NA2        m1165(.A(mai_mai_n962_), .B(mai_mai_n184_), .Y(mai_mai_n1215_));
  NA2        m1166(.A(mai_mai_n55_), .B(mai_mai_n103_), .Y(mai_mai_n1216_));
  INV        m1167(.A(mai_mai_n906_), .Y(mai_mai_n1217_));
  NO2        m1168(.A(mai_mai_n1217_), .B(mai_mai_n62_), .Y(mai_mai_n1218_));
  AOI220     m1169(.A0(mai_mai_n582_), .A1(mai_mai_n336_), .B0(mai_mai_n572_), .B1(mai_mai_n88_), .Y(mai_mai_n1219_));
  NA3        m1170(.A(mai_mai_n430_), .B(mai_mai_n539_), .C(mai_mai_n178_), .Y(mai_mai_n1220_));
  NO2        m1171(.A(mai_mai_n1220_), .B(mai_mai_n1219_), .Y(mai_mai_n1221_));
  NO2        m1172(.A(mai_mai_n1221_), .B(mai_mai_n1214_), .Y(mai_mai_n1222_));
  NO3        m1173(.A(x6), .B(x4), .C(x3), .Y(mai_mai_n1223_));
  NA2        m1174(.A(mai_mai_n1223_), .B(mai_mai_n493_), .Y(mai_mai_n1224_));
  NA4        m1175(.A(mai_mai_n651_), .B(mai_mai_n174_), .C(mai_mai_n58_), .D(x6), .Y(mai_mai_n1225_));
  AOI210     m1176(.A0(mai_mai_n1225_), .A1(mai_mai_n1224_), .B0(mai_mai_n54_), .Y(mai_mai_n1226_));
  NO2        m1177(.A(mai_mai_n606_), .B(mai_mai_n949_), .Y(mai_mai_n1227_));
  AN2        m1178(.A(mai_mai_n395_), .B(mai_mai_n1227_), .Y(mai_mai_n1228_));
  NO2        m1179(.A(mai_mai_n700_), .B(mai_mai_n471_), .Y(mai_mai_n1229_));
  NO3        m1180(.A(mai_mai_n1229_), .B(mai_mai_n236_), .C(mai_mai_n144_), .Y(mai_mai_n1230_));
  NO3        m1181(.A(mai_mai_n1230_), .B(mai_mai_n1228_), .C(mai_mai_n1226_), .Y(mai_mai_n1231_));
  NA2        m1182(.A(mai_mai_n380_), .B(mai_mai_n862_), .Y(mai_mai_n1232_));
  NA2        m1183(.A(mai_mai_n823_), .B(mai_mai_n1127_), .Y(mai_mai_n1233_));
  NA2        m1184(.A(mai_mai_n674_), .B(x7), .Y(mai_mai_n1234_));
  INV        m1185(.A(mai_mai_n1233_), .Y(mai_mai_n1235_));
  NA2        m1186(.A(mai_mai_n251_), .B(x2), .Y(mai_mai_n1236_));
  NO3        m1187(.A(mai_mai_n1236_), .B(mai_mai_n547_), .C(mai_mai_n72_), .Y(mai_mai_n1237_));
  OA210      m1188(.A0(mai_mai_n1094_), .A1(mai_mai_n58_), .B0(mai_mai_n716_), .Y(mai_mai_n1238_));
  AOI210     m1189(.A0(mai_mai_n532_), .A1(mai_mai_n50_), .B0(mai_mai_n542_), .Y(mai_mai_n1239_));
  OAI210     m1190(.A0(mai_mai_n840_), .A1(mai_mai_n850_), .B0(mai_mai_n358_), .Y(mai_mai_n1240_));
  OAI220     m1191(.A0(mai_mai_n1240_), .A1(mai_mai_n1239_), .B0(mai_mai_n1238_), .B1(mai_mai_n176_), .Y(mai_mai_n1241_));
  NO3        m1192(.A(mai_mai_n1241_), .B(mai_mai_n1237_), .C(mai_mai_n1235_), .Y(mai_mai_n1242_));
  OA220      m1193(.A0(mai_mai_n1242_), .A1(mai_mai_n411_), .B0(mai_mai_n1231_), .B1(mai_mai_n188_), .Y(mai_mai_n1243_));
  NO2        m1194(.A(mai_mai_n837_), .B(mai_mai_n55_), .Y(mai_mai_n1244_));
  NA2        m1195(.A(mai_mai_n391_), .B(mai_mai_n740_), .Y(mai_mai_n1245_));
  NO2        m1196(.A(mai_mai_n1245_), .B(mai_mai_n1244_), .Y(mai_mai_n1246_));
  NO3        m1197(.A(mai_mai_n863_), .B(mai_mai_n306_), .C(x8), .Y(mai_mai_n1247_));
  OAI210     m1198(.A0(mai_mai_n1247_), .A1(mai_mai_n1246_), .B0(x6), .Y(mai_mai_n1248_));
  INV        m1199(.A(mai_mai_n972_), .Y(mai_mai_n1249_));
  OAI220     m1200(.A0(mai_mai_n2220_), .A1(mai_mai_n1249_), .B0(mai_mai_n702_), .B1(mai_mai_n87_), .Y(mai_mai_n1250_));
  NA2        m1201(.A(mai_mai_n1250_), .B(mai_mai_n840_), .Y(mai_mai_n1251_));
  NA2        m1202(.A(mai_mai_n797_), .B(mai_mai_n71_), .Y(mai_mai_n1252_));
  AOI210     m1203(.A0(mai_mai_n459_), .A1(mai_mai_n57_), .B0(x2), .Y(mai_mai_n1253_));
  NA3        m1204(.A(mai_mai_n207_), .B(mai_mai_n76_), .C(mai_mai_n71_), .Y(mai_mai_n1254_));
  OAI210     m1205(.A0(mai_mai_n833_), .A1(mai_mai_n210_), .B0(mai_mai_n1254_), .Y(mai_mai_n1255_));
  AOI210     m1206(.A0(mai_mai_n1253_), .A1(mai_mai_n53_), .B0(mai_mai_n1255_), .Y(mai_mai_n1256_));
  NA3        m1207(.A(mai_mai_n1256_), .B(mai_mai_n1251_), .C(mai_mai_n1248_), .Y(mai_mai_n1257_));
  NO2        m1208(.A(mai_mai_n584_), .B(x6), .Y(mai_mai_n1258_));
  INV        m1209(.A(mai_mai_n356_), .Y(mai_mai_n1259_));
  OA210      m1210(.A0(mai_mai_n1259_), .A1(mai_mai_n1258_), .B0(mai_mai_n124_), .Y(mai_mai_n1260_));
  NO3        m1211(.A(mai_mai_n149_), .B(mai_mai_n75_), .C(x2), .Y(mai_mai_n1261_));
  INV        m1212(.A(mai_mai_n1260_), .Y(mai_mai_n1262_));
  NO2        m1213(.A(mai_mai_n210_), .B(x1), .Y(mai_mai_n1263_));
  OAI210     m1214(.A0(mai_mai_n1263_), .A1(mai_mai_n417_), .B0(mai_mai_n471_), .Y(mai_mai_n1264_));
  NO2        m1215(.A(mai_mai_n57_), .B(mai_mai_n103_), .Y(mai_mai_n1265_));
  NO2        m1216(.A(mai_mai_n1264_), .B(mai_mai_n56_), .Y(mai_mai_n1266_));
  NO2        m1217(.A(mai_mai_n493_), .B(mai_mai_n162_), .Y(mai_mai_n1267_));
  NA2        m1218(.A(mai_mai_n850_), .B(x4), .Y(mai_mai_n1268_));
  OAI220     m1219(.A0(mai_mai_n1268_), .A1(mai_mai_n632_), .B0(mai_mai_n592_), .B1(mai_mai_n561_), .Y(mai_mai_n1269_));
  NO3        m1220(.A(mai_mai_n1269_), .B(mai_mai_n1267_), .C(mai_mai_n1266_), .Y(mai_mai_n1270_));
  OAI210     m1221(.A0(mai_mai_n1262_), .A1(x5), .B0(mai_mai_n1270_), .Y(mai_mai_n1271_));
  AOI220     m1222(.A0(mai_mai_n1271_), .A1(mai_mai_n98_), .B0(mai_mai_n1257_), .B1(mai_mai_n313_), .Y(mai_mai_n1272_));
  NA4        m1223(.A(mai_mai_n1272_), .B(mai_mai_n1243_), .C(mai_mai_n1222_), .D(mai_mai_n1211_), .Y(mai17));
  NO3        m1224(.A(mai_mai_n552_), .B(mai_mai_n645_), .C(mai_mai_n99_), .Y(mai_mai_n1274_));
  NO2        m1225(.A(mai_mai_n120_), .B(mai_mai_n1024_), .Y(mai_mai_n1275_));
  AOI220     m1226(.A0(mai_mai_n1275_), .A1(mai_mai_n661_), .B0(mai_mai_n1274_), .B1(mai_mai_n465_), .Y(mai_mai_n1276_));
  NA2        m1227(.A(mai_mai_n153_), .B(mai_mai_n78_), .Y(mai_mai_n1277_));
  NOi21      m1228(.An(mai_mai_n356_), .B(mai_mai_n84_), .Y(mai_mai_n1278_));
  OAI210     m1229(.A0(mai_mai_n572_), .A1(mai_mai_n55_), .B0(mai_mai_n1278_), .Y(mai_mai_n1279_));
  NA2        m1230(.A(mai_mai_n1070_), .B(mai_mai_n901_), .Y(mai_mai_n1280_));
  NA4        m1231(.A(mai_mai_n1280_), .B(mai_mai_n1279_), .C(mai_mai_n677_), .D(mai_mai_n57_), .Y(mai_mai_n1281_));
  NA2        m1232(.A(x8), .B(mai_mai_n1127_), .Y(mai_mai_n1282_));
  NA3        m1233(.A(mai_mai_n1282_), .B(mai_mai_n1082_), .C(mai_mai_n373_), .Y(mai_mai_n1283_));
  NA3        m1234(.A(mai_mai_n367_), .B(mai_mai_n246_), .C(mai_mai_n538_), .Y(mai_mai_n1284_));
  OR2        m1235(.A(mai_mai_n1137_), .B(mai_mai_n1019_), .Y(mai_mai_n1285_));
  NA4        m1236(.A(mai_mai_n1285_), .B(mai_mai_n1284_), .C(mai_mai_n1283_), .D(mai_mai_n1281_), .Y(mai_mai_n1286_));
  AOI210     m1237(.A0(mai_mai_n1286_), .A1(x1), .B0(mai_mai_n59_), .Y(mai_mai_n1287_));
  NO2        m1238(.A(mai_mai_n876_), .B(mai_mai_n459_), .Y(mai_mai_n1288_));
  OAI210     m1239(.A0(mai_mai_n1288_), .A1(mai_mai_n953_), .B0(mai_mai_n558_), .Y(mai_mai_n1289_));
  NO2        m1240(.A(mai_mai_n1289_), .B(x8), .Y(mai_mai_n1290_));
  NO2        m1241(.A(mai_mai_n135_), .B(mai_mai_n134_), .Y(mai_mai_n1291_));
  NO3        m1242(.A(mai_mai_n817_), .B(mai_mai_n713_), .C(mai_mai_n645_), .Y(mai_mai_n1292_));
  AOI210     m1243(.A0(mai_mai_n1292_), .A1(mai_mai_n1291_), .B0(x0), .Y(mai_mai_n1293_));
  INV        m1244(.A(mai_mai_n1293_), .Y(mai_mai_n1294_));
  NO2        m1245(.A(mai_mai_n1294_), .B(mai_mai_n1290_), .Y(mai_mai_n1295_));
  OAI220     m1246(.A0(mai_mai_n1295_), .A1(mai_mai_n1287_), .B0(mai_mai_n1277_), .B1(mai_mai_n1276_), .Y(mai18));
  AOI210     m1247(.A0(x8), .A1(x0), .B0(x5), .Y(mai_mai_n1297_));
  NOi21      m1248(.An(mai_mai_n278_), .B(mai_mai_n939_), .Y(mai_mai_n1298_));
  NA2        m1249(.A(mai_mai_n552_), .B(mai_mai_n59_), .Y(mai_mai_n1299_));
  AOI210     m1250(.A0(mai_mai_n1215_), .A1(mai_mai_n324_), .B0(mai_mai_n1299_), .Y(mai_mai_n1300_));
  NO2        m1251(.A(mai_mai_n567_), .B(mai_mai_n714_), .Y(mai_mai_n1301_));
  NO3        m1252(.A(mai_mai_n749_), .B(mai_mai_n143_), .C(mai_mai_n70_), .Y(mai_mai_n1302_));
  NO4        m1253(.A(mai_mai_n1302_), .B(mai_mai_n1301_), .C(mai_mai_n1300_), .D(mai_mai_n1298_), .Y(mai_mai_n1303_));
  NO2        m1254(.A(mai_mai_n811_), .B(x5), .Y(mai_mai_n1304_));
  AOI210     m1255(.A0(mai_mai_n2223_), .A1(x5), .B0(mai_mai_n1304_), .Y(mai_mai_n1305_));
  OA220      m1256(.A0(mai_mai_n480_), .A1(mai_mai_n306_), .B0(mai_mai_n373_), .B1(x5), .Y(mai_mai_n1306_));
  OAI220     m1257(.A0(mai_mai_n1306_), .A1(mai_mai_n268_), .B0(mai_mai_n1305_), .B1(mai_mai_n197_), .Y(mai_mai_n1307_));
  AOI210     m1258(.A0(mai_mai_n362_), .A1(mai_mai_n266_), .B0(mai_mai_n1307_), .Y(mai_mai_n1308_));
  AOI210     m1259(.A0(mai_mai_n1308_), .A1(mai_mai_n1303_), .B0(x6), .Y(mai_mai_n1309_));
  NA3        m1260(.A(mai_mai_n484_), .B(mai_mai_n393_), .C(x2), .Y(mai_mai_n1310_));
  NA3        m1261(.A(mai_mai_n939_), .B(mai_mai_n51_), .C(mai_mai_n57_), .Y(mai_mai_n1311_));
  AOI210     m1262(.A0(mai_mai_n1311_), .A1(mai_mai_n1310_), .B0(mai_mai_n726_), .Y(mai_mai_n1312_));
  NA2        m1263(.A(mai_mai_n246_), .B(x6), .Y(mai_mai_n1313_));
  NO2        m1264(.A(x7), .B(mai_mai_n1313_), .Y(mai_mai_n1314_));
  OAI210     m1265(.A0(mai_mai_n1314_), .A1(mai_mai_n1312_), .B0(mai_mai_n53_), .Y(mai_mai_n1315_));
  NO2        m1266(.A(mai_mai_n631_), .B(mai_mai_n239_), .Y(mai_mai_n1316_));
  NO2        m1267(.A(mai_mai_n242_), .B(x3), .Y(mai_mai_n1317_));
  NA2        m1268(.A(mai_mai_n1316_), .B(mai_mai_n1317_), .Y(mai_mai_n1318_));
  AOI210     m1269(.A0(mai_mai_n1013_), .A1(mai_mai_n566_), .B0(x4), .Y(mai_mai_n1319_));
  OAI210     m1270(.A0(mai_mai_n513_), .A1(mai_mai_n552_), .B0(mai_mai_n59_), .Y(mai_mai_n1320_));
  OAI210     m1271(.A0(mai_mai_n572_), .A1(mai_mai_n593_), .B0(mai_mai_n1320_), .Y(mai_mai_n1321_));
  NA2        m1272(.A(mai_mai_n1321_), .B(mai_mai_n150_), .Y(mai_mai_n1322_));
  NA4        m1273(.A(mai_mai_n1322_), .B(mai_mai_n1319_), .C(mai_mai_n1318_), .D(mai_mai_n1315_), .Y(mai_mai_n1323_));
  NO3        m1274(.A(mai_mai_n960_), .B(mai_mai_n124_), .C(mai_mai_n123_), .Y(mai_mai_n1324_));
  OAI210     m1275(.A0(mai_mai_n1324_), .A1(mai_mai_n598_), .B0(mai_mai_n103_), .Y(mai_mai_n1325_));
  NO2        m1276(.A(mai_mai_n1325_), .B(mai_mai_n726_), .Y(mai_mai_n1326_));
  NA3        m1277(.A(mai_mai_n962_), .B(mai_mai_n715_), .C(mai_mai_n317_), .Y(mai_mai_n1327_));
  NA2        m1278(.A(mai_mai_n160_), .B(mai_mai_n713_), .Y(mai_mai_n1328_));
  OAI210     m1279(.A0(mai_mai_n1328_), .A1(mai_mai_n1140_), .B0(mai_mai_n1327_), .Y(mai_mai_n1329_));
  AOI210     m1280(.A0(x2), .A1(mai_mai_n167_), .B0(mai_mai_n1329_), .Y(mai_mai_n1330_));
  OAI210     m1281(.A0(mai_mai_n1330_), .A1(mai_mai_n502_), .B0(x4), .Y(mai_mai_n1331_));
  OAI220     m1282(.A0(mai_mai_n1331_), .A1(mai_mai_n1326_), .B0(mai_mai_n1323_), .B1(mai_mai_n1309_), .Y(mai_mai_n1332_));
  NO2        m1283(.A(mai_mai_n137_), .B(mai_mai_n118_), .Y(mai_mai_n1333_));
  NO2        m1284(.A(mai_mai_n176_), .B(mai_mai_n740_), .Y(mai_mai_n1334_));
  NO2        m1285(.A(mai_mai_n361_), .B(mai_mai_n231_), .Y(mai_mai_n1335_));
  NO2        m1286(.A(mai_mai_n124_), .B(mai_mai_n679_), .Y(mai_mai_n1336_));
  NO2        m1287(.A(mai_mai_n863_), .B(mai_mai_n538_), .Y(mai_mai_n1337_));
  AO220      m1288(.A0(mai_mai_n1337_), .A1(mai_mai_n1336_), .B0(mai_mai_n1335_), .B1(mai_mai_n120_), .Y(mai_mai_n1338_));
  NO3        m1289(.A(mai_mai_n1338_), .B(mai_mai_n1334_), .C(mai_mai_n1333_), .Y(mai_mai_n1339_));
  NA2        m1290(.A(mai_mai_n960_), .B(x3), .Y(mai_mai_n1340_));
  NA2        m1291(.A(mai_mai_n1169_), .B(mai_mai_n125_), .Y(mai_mai_n1341_));
  OAI220     m1292(.A0(mai_mai_n1341_), .A1(mai_mai_n1340_), .B0(mai_mai_n1339_), .B1(x3), .Y(mai_mai_n1342_));
  NO3        m1293(.A(mai_mai_n894_), .B(mai_mai_n631_), .C(mai_mai_n301_), .Y(mai_mai_n1343_));
  AO210      m1294(.A0(mai_mai_n920_), .A1(mai_mai_n272_), .B0(mai_mai_n1343_), .Y(mai_mai_n1344_));
  AOI220     m1295(.A0(mai_mai_n1344_), .A1(x8), .B0(mai_mai_n1169_), .B1(mai_mai_n403_), .Y(mai_mai_n1345_));
  NA2        m1296(.A(mai_mai_n690_), .B(mai_mai_n292_), .Y(mai_mai_n1346_));
  NO4        m1297(.A(mai_mai_n342_), .B(mai_mai_n186_), .C(mai_mai_n312_), .D(x2), .Y(mai_mai_n1347_));
  NA2        m1298(.A(mai_mai_n1216_), .B(mai_mai_n105_), .Y(mai_mai_n1348_));
  NO3        m1299(.A(mai_mai_n1064_), .B(mai_mai_n887_), .C(mai_mai_n1010_), .Y(mai_mai_n1349_));
  AOI210     m1300(.A0(mai_mai_n1349_), .A1(mai_mai_n1348_), .B0(mai_mai_n1347_), .Y(mai_mai_n1350_));
  OA220      m1301(.A0(mai_mai_n1350_), .A1(mai_mai_n863_), .B0(mai_mai_n1346_), .B1(mai_mai_n524_), .Y(mai_mai_n1351_));
  OAI210     m1302(.A0(mai_mai_n1345_), .A1(mai_mai_n383_), .B0(mai_mai_n1351_), .Y(mai_mai_n1352_));
  AOI210     m1303(.A0(mai_mai_n1342_), .A1(mai_mai_n130_), .B0(mai_mai_n1352_), .Y(mai_mai_n1353_));
  NA2        m1304(.A(mai_mai_n1353_), .B(mai_mai_n1332_), .Y(mai19));
  NO2        m1305(.A(mai_mai_n1252_), .B(mai_mai_n235_), .Y(mai_mai_n1355_));
  NA2        m1306(.A(mai_mai_n593_), .B(x3), .Y(mai_mai_n1356_));
  OAI210     m1307(.A0(mai_mai_n143_), .A1(mai_mai_n104_), .B0(mai_mai_n81_), .Y(mai_mai_n1357_));
  NA3        m1308(.A(mai_mai_n1357_), .B(mai_mai_n1356_), .C(mai_mai_n221_), .Y(mai_mai_n1358_));
  NA2        m1309(.A(mai_mai_n1274_), .B(mai_mai_n327_), .Y(mai_mai_n1359_));
  AOI210     m1310(.A0(mai_mai_n1359_), .A1(mai_mai_n1358_), .B0(mai_mai_n56_), .Y(mai_mai_n1360_));
  NO2        m1311(.A(mai_mai_n786_), .B(mai_mai_n1071_), .Y(mai_mai_n1361_));
  OAI210     m1312(.A0(mai_mai_n1360_), .A1(mai_mai_n1355_), .B0(mai_mai_n1361_), .Y(mai_mai_n1362_));
  INV        m1313(.A(mai_mai_n1058_), .Y(mai_mai_n1363_));
  NO2        m1314(.A(mai_mai_n502_), .B(mai_mai_n570_), .Y(mai_mai_n1364_));
  NA2        m1315(.A(mai_mai_n1094_), .B(mai_mai_n50_), .Y(mai_mai_n1365_));
  NO3        m1316(.A(mai_mai_n478_), .B(mai_mai_n280_), .C(mai_mai_n64_), .Y(mai_mai_n1366_));
  NA2        m1317(.A(mai_mai_n1366_), .B(mai_mai_n1365_), .Y(mai_mai_n1367_));
  NA2        m1318(.A(mai_mai_n2219_), .B(mai_mai_n713_), .Y(mai_mai_n1368_));
  AOI210     m1319(.A0(mai_mai_n758_), .A1(mai_mai_n679_), .B0(mai_mai_n703_), .Y(mai_mai_n1369_));
  NO2        m1320(.A(mai_mai_n1369_), .B(x4), .Y(mai_mai_n1370_));
  NA3        m1321(.A(mai_mai_n677_), .B(mai_mai_n234_), .C(x7), .Y(mai_mai_n1371_));
  AOI210     m1322(.A0(mai_mai_n1212_), .A1(mai_mai_n726_), .B0(mai_mai_n645_), .Y(mai_mai_n1372_));
  AOI210     m1323(.A0(mai_mai_n1372_), .A1(mai_mai_n1371_), .B0(mai_mai_n463_), .Y(mai_mai_n1373_));
  OAI210     m1324(.A0(mai_mai_n1373_), .A1(mai_mai_n1370_), .B0(mai_mai_n749_), .Y(mai_mai_n1374_));
  NO2        m1325(.A(mai_mai_n143_), .B(mai_mai_n916_), .Y(mai_mai_n1375_));
  NA2        m1326(.A(mai_mai_n1375_), .B(mai_mai_n1107_), .Y(mai_mai_n1376_));
  AO210      m1327(.A0(mai_mai_n1376_), .A1(mai_mai_n1374_), .B0(x1), .Y(mai_mai_n1377_));
  NA2        m1328(.A(mai_mai_n138_), .B(mai_mai_n106_), .Y(mai_mai_n1378_));
  NOi21      m1329(.An(x1), .B(x6), .Y(mai_mai_n1379_));
  NA2        m1330(.A(mai_mai_n1379_), .B(mai_mai_n84_), .Y(mai_mai_n1380_));
  INV        m1331(.A(mai_mai_n1378_), .Y(mai_mai_n1381_));
  AOI220     m1332(.A0(mai_mai_n1381_), .A1(x3), .B0(mai_mai_n1065_), .B1(mai_mai_n357_), .Y(mai_mai_n1382_));
  NA3        m1333(.A(mai_mai_n1070_), .B(mai_mai_n735_), .C(mai_mai_n554_), .Y(mai_mai_n1383_));
  AOI220     m1334(.A0(mai_mai_n1096_), .A1(mai_mai_n117_), .B0(mai_mai_n837_), .B1(mai_mai_n751_), .Y(mai_mai_n1384_));
  AOI210     m1335(.A0(mai_mai_n1384_), .A1(mai_mai_n1383_), .B0(mai_mai_n296_), .Y(mai_mai_n1385_));
  NA2        m1336(.A(mai_mai_n850_), .B(mai_mai_n50_), .Y(mai_mai_n1386_));
  NA3        m1337(.A(mai_mai_n1058_), .B(mai_mai_n358_), .C(mai_mai_n105_), .Y(mai_mai_n1387_));
  AOI210     m1338(.A0(mai_mai_n1387_), .A1(mai_mai_n1386_), .B0(mai_mai_n872_), .Y(mai_mai_n1388_));
  NO3        m1339(.A(mai_mai_n568_), .B(mai_mai_n477_), .C(mai_mai_n1073_), .Y(mai_mai_n1389_));
  NO3        m1340(.A(mai_mai_n1389_), .B(mai_mai_n1388_), .C(mai_mai_n1385_), .Y(mai_mai_n1390_));
  OAI210     m1341(.A0(mai_mai_n1382_), .A1(mai_mai_n774_), .B0(mai_mai_n1390_), .Y(mai_mai_n1391_));
  NA2        m1342(.A(mai_mai_n1173_), .B(mai_mai_n674_), .Y(mai_mai_n1392_));
  NO2        m1343(.A(mai_mai_n54_), .B(mai_mai_n71_), .Y(mai_mai_n1393_));
  AO220      m1344(.A0(mai_mai_n1393_), .A1(mai_mai_n894_), .B0(mai_mai_n751_), .B1(mai_mai_n862_), .Y(mai_mai_n1394_));
  NA2        m1345(.A(mai_mai_n1044_), .B(mai_mai_n334_), .Y(mai_mai_n1395_));
  NO2        m1346(.A(mai_mai_n887_), .B(mai_mai_n1379_), .Y(mai_mai_n1396_));
  NA2        m1347(.A(mai_mai_n459_), .B(mai_mai_n674_), .Y(mai_mai_n1397_));
  OAI210     m1348(.A0(mai_mai_n1397_), .A1(mai_mai_n1396_), .B0(mai_mai_n1395_), .Y(mai_mai_n1398_));
  AOI210     m1349(.A0(mai_mai_n1394_), .A1(x2), .B0(mai_mai_n1398_), .Y(mai_mai_n1399_));
  OAI220     m1350(.A0(mai_mai_n1399_), .A1(mai_mai_n143_), .B0(mai_mai_n1392_), .B1(mai_mai_n54_), .Y(mai_mai_n1400_));
  OAI210     m1351(.A0(mai_mai_n1400_), .A1(mai_mai_n1391_), .B0(x8), .Y(mai_mai_n1401_));
  NA4        m1352(.A(mai_mai_n1401_), .B(mai_mai_n1377_), .C(mai_mai_n1368_), .D(mai_mai_n1362_), .Y(mai20));
  NA4        m1353(.A(mai_mai_n366_), .B(mai_mai_n255_), .C(mai_mai_n356_), .D(mai_mai_n62_), .Y(mai_mai_n1403_));
  NA2        m1354(.A(mai_mai_n444_), .B(mai_mai_n387_), .Y(mai_mai_n1404_));
  AOI210     m1355(.A0(mai_mai_n1404_), .A1(mai_mai_n1403_), .B0(mai_mai_n87_), .Y(mai_mai_n1405_));
  AOI210     m1356(.A0(mai_mai_n945_), .A1(mai_mai_n62_), .B0(mai_mai_n1364_), .Y(mai_mai_n1406_));
  INV        m1357(.A(mai_mai_n1050_), .Y(mai_mai_n1407_));
  OAI210     m1358(.A0(mai_mai_n1406_), .A1(mai_mai_n627_), .B0(mai_mai_n1407_), .Y(mai_mai_n1408_));
  OAI210     m1359(.A0(mai_mai_n1408_), .A1(mai_mai_n1405_), .B0(mai_mai_n984_), .Y(mai_mai_n1409_));
  NAi21      m1360(.An(mai_mai_n509_), .B(mai_mai_n375_), .Y(mai_mai_n1410_));
  NA3        m1361(.A(mai_mai_n983_), .B(mai_mai_n255_), .C(mai_mai_n537_), .Y(mai_mai_n1411_));
  NO2        m1362(.A(mai_mai_n1411_), .B(mai_mai_n1127_), .Y(mai_mai_n1412_));
  NO2        m1363(.A(mai_mai_n690_), .B(mai_mai_n874_), .Y(mai_mai_n1413_));
  NA2        m1364(.A(mai_mai_n1412_), .B(mai_mai_n301_), .Y(mai_mai_n1414_));
  NO4        m1365(.A(mai_mai_n506_), .B(mai_mai_n216_), .C(x5), .D(x2), .Y(mai_mai_n1415_));
  NA2        m1366(.A(mai_mai_n292_), .B(mai_mai_n93_), .Y(mai_mai_n1416_));
  NA2        m1367(.A(mai_mai_n302_), .B(mai_mai_n103_), .Y(mai_mai_n1417_));
  NA2        m1368(.A(mai_mai_n395_), .B(mai_mai_n52_), .Y(mai_mai_n1418_));
  OAI220     m1369(.A0(mai_mai_n1418_), .A1(mai_mai_n1417_), .B0(mai_mai_n1416_), .B1(mai_mai_n250_), .Y(mai_mai_n1419_));
  OAI210     m1370(.A0(mai_mai_n1419_), .A1(mai_mai_n1415_), .B0(mai_mai_n204_), .Y(mai_mai_n1420_));
  NO2        m1371(.A(mai_mai_n612_), .B(mai_mai_n558_), .Y(mai_mai_n1421_));
  NA2        m1372(.A(mai_mai_n863_), .B(mai_mai_n50_), .Y(mai_mai_n1422_));
  NO3        m1373(.A(mai_mai_n1422_), .B(mai_mai_n340_), .C(mai_mai_n209_), .Y(mai_mai_n1423_));
  NA4        m1374(.A(mai_mai_n313_), .B(mai_mai_n218_), .C(mai_mai_n740_), .D(mai_mai_n64_), .Y(mai_mai_n1424_));
  OAI220     m1375(.A0(mai_mai_n1424_), .A1(mai_mai_n621_), .B0(mai_mai_n1268_), .B1(mai_mai_n928_), .Y(mai_mai_n1425_));
  AOI210     m1376(.A0(mai_mai_n1423_), .A1(mai_mai_n1421_), .B0(mai_mai_n1425_), .Y(mai_mai_n1426_));
  NA4        m1377(.A(mai_mai_n1426_), .B(mai_mai_n1420_), .C(mai_mai_n1414_), .D(mai_mai_n1409_), .Y(mai21));
  NO2        m1378(.A(mai_mai_n946_), .B(mai_mai_n96_), .Y(mai_mai_n1428_));
  NA2        m1379(.A(mai_mai_n1428_), .B(mai_mai_n78_), .Y(mai_mai_n1429_));
  NA2        m1380(.A(mai_mai_n266_), .B(mai_mai_n784_), .Y(mai_mai_n1430_));
  AOI210     m1381(.A0(mai_mai_n1430_), .A1(mai_mai_n282_), .B0(mai_mai_n524_), .Y(mai_mai_n1431_));
  NA2        m1382(.A(mai_mai_n850_), .B(mai_mai_n249_), .Y(mai_mai_n1432_));
  NA2        m1383(.A(mai_mai_n497_), .B(mai_mai_n429_), .Y(mai_mai_n1433_));
  NA3        m1384(.A(mai_mai_n1432_), .B(mai_mai_n1196_), .C(mai_mai_n56_), .Y(mai_mai_n1434_));
  NO3        m1385(.A(x5), .B(mai_mai_n668_), .C(mai_mai_n228_), .Y(mai_mai_n1435_));
  NOi21      m1386(.An(mai_mai_n179_), .B(mai_mai_n974_), .Y(mai_mai_n1436_));
  NO4        m1387(.A(mai_mai_n1436_), .B(mai_mai_n1435_), .C(mai_mai_n1434_), .D(mai_mai_n1431_), .Y(mai_mai_n1437_));
  OAI210     m1388(.A0(mai_mai_n725_), .A1(mai_mai_n542_), .B0(mai_mai_n315_), .Y(mai_mai_n1438_));
  NO2        m1389(.A(mai_mai_n70_), .B(x2), .Y(mai_mai_n1439_));
  INV        m1390(.A(mai_mai_n1438_), .Y(mai_mai_n1440_));
  NA2        m1391(.A(mai_mai_n1440_), .B(x8), .Y(mai_mai_n1441_));
  NO3        m1392(.A(mai_mai_n714_), .B(mai_mai_n571_), .C(mai_mai_n538_), .Y(mai_mai_n1442_));
  NA2        m1393(.A(mai_mai_n55_), .B(mai_mai_n50_), .Y(mai_mai_n1443_));
  MUX2       m1394(.S(mai_mai_n552_), .A(mai_mai_n1443_), .B(mai_mai_n102_), .Y(mai_mai_n1444_));
  NO2        m1395(.A(mai_mai_n1177_), .B(mai_mai_n1444_), .Y(mai_mai_n1445_));
  OAI210     m1396(.A0(mai_mai_n590_), .A1(mai_mai_n537_), .B0(x4), .Y(mai_mai_n1446_));
  NO3        m1397(.A(mai_mai_n1446_), .B(mai_mai_n1445_), .C(mai_mai_n1442_), .Y(mai_mai_n1447_));
  AO220      m1398(.A0(mai_mai_n1447_), .A1(mai_mai_n1441_), .B0(mai_mai_n1437_), .B1(mai_mai_n1429_), .Y(mai_mai_n1448_));
  AN2        m1399(.A(mai_mai_n578_), .B(mai_mai_n296_), .Y(mai_mai_n1449_));
  NO2        m1400(.A(mai_mai_n786_), .B(x0), .Y(mai_mai_n1450_));
  NO3        m1401(.A(mai_mai_n1450_), .B(mai_mai_n507_), .C(mai_mai_n88_), .Y(mai_mai_n1451_));
  NO2        m1402(.A(mai_mai_n149_), .B(x2), .Y(mai_mai_n1452_));
  NA2        m1403(.A(mai_mai_n1452_), .B(mai_mai_n68_), .Y(mai_mai_n1453_));
  OAI210     m1404(.A0(mai_mai_n1451_), .A1(mai_mai_n373_), .B0(mai_mai_n1453_), .Y(mai_mai_n1454_));
  AOI220     m1405(.A0(mai_mai_n1454_), .A1(x5), .B0(mai_mai_n1449_), .B1(mai_mai_n690_), .Y(mai_mai_n1455_));
  AOI210     m1406(.A0(mai_mai_n1455_), .A1(mai_mai_n1448_), .B0(mai_mai_n71_), .Y(mai_mai_n1456_));
  NO2        m1407(.A(mai_mai_n827_), .B(mai_mai_n158_), .Y(mai_mai_n1457_));
  NOi31      m1408(.An(mai_mai_n1236_), .B(mai_mai_n1297_), .C(mai_mai_n1023_), .Y(mai_mai_n1458_));
  NA2        m1409(.A(mai_mai_n1458_), .B(mai_mai_n1457_), .Y(mai_mai_n1459_));
  OAI210     m1410(.A0(mai_mai_n264_), .A1(mai_mai_n147_), .B0(mai_mai_n2218_), .Y(mai_mai_n1460_));
  OAI210     m1411(.A0(mai_mai_n382_), .A1(mai_mai_n396_), .B0(mai_mai_n209_), .Y(mai_mai_n1461_));
  NA2        m1412(.A(x7), .B(mai_mai_n1461_), .Y(mai_mai_n1462_));
  AOI210     m1413(.A0(mai_mai_n1460_), .A1(mai_mai_n1459_), .B0(mai_mai_n1462_), .Y(mai_mai_n1463_));
  NA2        m1414(.A(mai_mai_n700_), .B(mai_mai_n509_), .Y(mai_mai_n1464_));
  AO210      m1415(.A0(mai_mai_n1464_), .A1(mai_mai_n872_), .B0(mai_mai_n50_), .Y(mai_mai_n1465_));
  AOI220     m1416(.A0(x4), .A1(mai_mai_n1033_), .B0(mai_mai_n1152_), .B1(mai_mai_n939_), .Y(mai_mai_n1466_));
  AOI210     m1417(.A0(mai_mai_n1466_), .A1(mai_mai_n1465_), .B0(mai_mai_n105_), .Y(mai_mai_n1467_));
  NO2        m1418(.A(mai_mai_n1467_), .B(mai_mai_n1463_), .Y(mai_mai_n1468_));
  NO2        m1419(.A(mai_mai_n1468_), .B(x6), .Y(mai_mai_n1469_));
  NO2        m1420(.A(mai_mai_n561_), .B(mai_mai_n1297_), .Y(mai_mai_n1470_));
  OAI210     m1421(.A0(mai_mai_n1470_), .A1(mai_mai_n634_), .B0(mai_mai_n56_), .Y(mai_mai_n1471_));
  NO2        m1422(.A(mai_mai_n692_), .B(mai_mai_n54_), .Y(mai_mai_n1472_));
  NO4        m1423(.A(mai_mai_n870_), .B(mai_mai_n253_), .C(mai_mai_n713_), .D(mai_mai_n698_), .Y(mai_mai_n1473_));
  NO2        m1424(.A(mai_mai_n791_), .B(x5), .Y(mai_mai_n1474_));
  NO4        m1425(.A(mai_mai_n1474_), .B(mai_mai_n1473_), .C(mai_mai_n1472_), .D(mai_mai_n857_), .Y(mai_mai_n1475_));
  AOI210     m1426(.A0(mai_mai_n1475_), .A1(mai_mai_n1471_), .B0(mai_mai_n50_), .Y(mai_mai_n1476_));
  NA2        m1427(.A(mai_mai_n149_), .B(mai_mai_n103_), .Y(mai_mai_n1477_));
  OA220      m1428(.A0(mai_mai_n1477_), .A1(mai_mai_n406_), .B0(mai_mai_n434_), .B1(mai_mai_n690_), .Y(mai_mai_n1478_));
  NA3        m1429(.A(mai_mai_n55_), .B(x2), .C(x0), .Y(mai_mai_n1479_));
  AOI220     m1430(.A0(mai_mai_n1479_), .A1(mai_mai_n160_), .B0(mai_mai_n791_), .B1(mai_mai_n145_), .Y(mai_mai_n1480_));
  NO2        m1431(.A(mai_mai_n627_), .B(mai_mai_n234_), .Y(mai_mai_n1481_));
  NO3        m1432(.A(mai_mai_n225_), .B(mai_mai_n207_), .C(mai_mai_n334_), .Y(mai_mai_n1482_));
  NO3        m1433(.A(mai_mai_n1482_), .B(mai_mai_n1481_), .C(mai_mai_n1480_), .Y(mai_mai_n1483_));
  OAI220     m1434(.A0(mai_mai_n1483_), .A1(mai_mai_n56_), .B0(mai_mai_n1478_), .B1(mai_mai_n643_), .Y(mai_mai_n1484_));
  OAI210     m1435(.A0(mai_mai_n1484_), .A1(mai_mai_n1476_), .B0(mai_mai_n111_), .Y(mai_mai_n1485_));
  NO2        m1436(.A(mai_mai_n565_), .B(mai_mai_n277_), .Y(mai_mai_n1486_));
  AOI210     m1437(.A0(mai_mai_n559_), .A1(x5), .B0(mai_mai_n1486_), .Y(mai_mai_n1487_));
  NO2        m1438(.A(mai_mai_n1487_), .B(mai_mai_n105_), .Y(mai_mai_n1488_));
  NA2        m1439(.A(mai_mai_n651_), .B(mai_mai_n81_), .Y(mai_mai_n1489_));
  NA3        m1440(.A(mai_mai_n1489_), .B(mai_mai_n400_), .C(mai_mai_n57_), .Y(mai_mai_n1490_));
  INV        m1441(.A(mai_mai_n1490_), .Y(mai_mai_n1491_));
  OAI210     m1442(.A0(mai_mai_n1491_), .A1(mai_mai_n1488_), .B0(x1), .Y(mai_mai_n1492_));
  NO4        m1443(.A(mai_mai_n391_), .B(mai_mai_n78_), .C(mai_mai_n139_), .D(x3), .Y(mai_mai_n1493_));
  NO2        m1444(.A(mai_mai_n302_), .B(mai_mai_n107_), .Y(mai_mai_n1494_));
  OAI210     m1445(.A0(mai_mai_n1493_), .A1(mai_mai_n1128_), .B0(mai_mai_n1494_), .Y(mai_mai_n1495_));
  NO2        m1446(.A(mai_mai_n60_), .B(mai_mai_n103_), .Y(mai_mai_n1496_));
  NA2        m1447(.A(mai_mai_n1496_), .B(mai_mai_n1334_), .Y(mai_mai_n1497_));
  NA4        m1448(.A(mai_mai_n1497_), .B(mai_mai_n1495_), .C(mai_mai_n1492_), .D(mai_mai_n1485_), .Y(mai_mai_n1498_));
  NO3        m1449(.A(mai_mai_n1498_), .B(mai_mai_n1469_), .C(mai_mai_n1456_), .Y(mai22));
  AOI210     m1450(.A0(mai_mai_n484_), .A1(mai_mai_n71_), .B0(mai_mai_n437_), .Y(mai_mai_n1500_));
  AOI210     m1451(.A0(x5), .A1(x2), .B0(x8), .Y(mai_mai_n1501_));
  NA2        m1452(.A(mai_mai_n1501_), .B(mai_mai_n59_), .Y(mai_mai_n1502_));
  OAI220     m1453(.A0(mai_mai_n1502_), .A1(mai_mai_n293_), .B0(mai_mai_n1500_), .B1(mai_mai_n373_), .Y(mai_mai_n1503_));
  NA2        m1454(.A(mai_mai_n537_), .B(mai_mai_n87_), .Y(mai_mai_n1504_));
  NA2        m1455(.A(mai_mai_n250_), .B(mai_mai_n77_), .Y(mai_mai_n1505_));
  OA220      m1456(.A0(mai_mai_n1505_), .A1(mai_mai_n1504_), .B0(mai_mai_n771_), .B1(mai_mai_n901_), .Y(mai_mai_n1506_));
  NO4        m1457(.A(mai_mai_n361_), .B(mai_mai_n203_), .C(mai_mai_n71_), .D(x3), .Y(mai_mai_n1507_));
  NO3        m1458(.A(mai_mai_n1091_), .B(mai_mai_n87_), .C(x0), .Y(mai_mai_n1508_));
  OAI210     m1459(.A0(mai_mai_n373_), .A1(mai_mai_n188_), .B0(x4), .Y(mai_mai_n1509_));
  NO2        m1460(.A(mai_mai_n1509_), .B(mai_mai_n1507_), .Y(mai_mai_n1510_));
  OAI210     m1461(.A0(mai_mai_n1506_), .A1(mai_mai_n184_), .B0(mai_mai_n1510_), .Y(mai_mai_n1511_));
  AOI210     m1462(.A0(mai_mai_n1503_), .A1(mai_mai_n53_), .B0(mai_mai_n1511_), .Y(mai_mai_n1512_));
  NA2        m1463(.A(mai_mai_n275_), .B(mai_mai_n280_), .Y(mai_mai_n1513_));
  NA3        m1464(.A(mai_mai_n1513_), .B(mai_mai_n204_), .C(mai_mai_n279_), .Y(mai_mai_n1514_));
  NA2        m1465(.A(mai_mai_n532_), .B(mai_mai_n224_), .Y(mai_mai_n1515_));
  NA2        m1466(.A(mai_mai_n1515_), .B(mai_mai_n1514_), .Y(mai_mai_n1516_));
  NO2        m1467(.A(mai_mai_n1091_), .B(x3), .Y(mai_mai_n1517_));
  NA2        m1468(.A(mai_mai_n1517_), .B(mai_mai_n323_), .Y(mai_mai_n1518_));
  OAI210     m1469(.A0(mai_mai_n972_), .A1(mai_mai_n175_), .B0(mai_mai_n56_), .Y(mai_mai_n1519_));
  NO2        m1470(.A(mai_mai_n340_), .B(mai_mai_n196_), .Y(mai_mai_n1520_));
  NO2        m1471(.A(mai_mai_n1520_), .B(mai_mai_n1519_), .Y(mai_mai_n1521_));
  OAI210     m1472(.A0(mai_mai_n1518_), .A1(mai_mai_n234_), .B0(mai_mai_n1521_), .Y(mai_mai_n1522_));
  AOI210     m1473(.A0(mai_mai_n1516_), .A1(mai_mai_n103_), .B0(mai_mai_n1522_), .Y(mai_mai_n1523_));
  OR2        m1474(.A(mai_mai_n1523_), .B(mai_mai_n1512_), .Y(mai_mai_n1524_));
  NA2        m1475(.A(mai_mai_n650_), .B(mai_mai_n638_), .Y(mai_mai_n1525_));
  NO2        m1476(.A(mai_mai_n328_), .B(x0), .Y(mai_mai_n1526_));
  NA3        m1477(.A(mai_mai_n1526_), .B(mai_mai_n323_), .C(mai_mai_n56_), .Y(mai_mai_n1527_));
  AOI210     m1478(.A0(mai_mai_n1527_), .A1(mai_mai_n1525_), .B0(mai_mai_n373_), .Y(mai_mai_n1528_));
  NA2        m1479(.A(mai_mai_n391_), .B(x3), .Y(mai_mai_n1529_));
  NO3        m1480(.A(mai_mai_n786_), .B(mai_mai_n433_), .C(mai_mai_n105_), .Y(mai_mai_n1530_));
  NO2        m1481(.A(mai_mai_n973_), .B(mai_mai_n134_), .Y(mai_mai_n1531_));
  NO3        m1482(.A(mai_mai_n817_), .B(mai_mai_n387_), .C(mai_mai_n276_), .Y(mai_mai_n1532_));
  AOI220     m1483(.A0(mai_mai_n1532_), .A1(mai_mai_n1531_), .B0(mai_mai_n1530_), .B1(mai_mai_n1526_), .Y(mai_mai_n1533_));
  NA3        m1484(.A(mai_mai_n56_), .B(mai_mai_n50_), .C(x0), .Y(mai_mai_n1534_));
  BUFFER     m1485(.A(mai_mai_n83_), .Y(mai_mai_n1535_));
  NA3        m1486(.A(x6), .B(x4), .C(mai_mai_n50_), .Y(mai_mai_n1536_));
  NA2        m1487(.A(mai_mai_n387_), .B(mai_mai_n323_), .Y(mai_mai_n1537_));
  NA2        m1488(.A(mai_mai_n1537_), .B(mai_mai_n1533_), .Y(mai_mai_n1538_));
  AOI210     m1489(.A0(mai_mai_n1538_), .A1(x7), .B0(mai_mai_n1528_), .Y(mai_mai_n1539_));
  OAI210     m1490(.A0(mai_mai_n1524_), .A1(x7), .B0(mai_mai_n1539_), .Y(mai23));
  OR2        m1491(.A(mai_mai_n478_), .B(mai_mai_n204_), .Y(mai_mai_n1541_));
  AOI220     m1492(.A0(mai_mai_n1541_), .A1(mai_mai_n1413_), .B0(mai_mai_n566_), .B1(mai_mai_n269_), .Y(mai_mai_n1542_));
  NO3        m1493(.A(mai_mai_n771_), .B(mai_mai_n546_), .C(mai_mai_n450_), .Y(mai_mai_n1543_));
  NO3        m1494(.A(mai_mai_n864_), .B(mai_mai_n140_), .C(mai_mai_n112_), .Y(mai_mai_n1544_));
  AOI210     m1495(.A0(mai_mai_n1544_), .A1(mai_mai_n923_), .B0(mai_mai_n1543_), .Y(mai_mai_n1545_));
  OAI210     m1496(.A0(mai_mai_n1542_), .A1(mai_mai_n143_), .B0(mai_mai_n1545_), .Y(mai_mai_n1546_));
  NA2        m1497(.A(mai_mai_n1546_), .B(mai_mai_n55_), .Y(mai_mai_n1547_));
  INV        m1498(.A(mai_mai_n476_), .Y(mai_mai_n1548_));
  AN2        m1499(.A(mai_mai_n894_), .B(mai_mai_n690_), .Y(mai_mai_n1549_));
  OAI210     m1500(.A0(mai_mai_n1549_), .A1(mai_mai_n1548_), .B0(mai_mai_n543_), .Y(mai_mai_n1550_));
  INV        m1501(.A(mai_mai_n158_), .Y(mai_mai_n1551_));
  NA2        m1502(.A(mai_mai_n379_), .B(mai_mai_n150_), .Y(mai_mai_n1552_));
  AOI210     m1503(.A0(mai_mai_n1552_), .A1(mai_mai_n1551_), .B0(mai_mai_n216_), .Y(mai_mai_n1553_));
  AOI210     m1504(.A0(mai_mai_n50_), .A1(mai_mai_n461_), .B0(mai_mai_n358_), .Y(mai_mai_n1554_));
  OAI210     m1505(.A0(mai_mai_n1554_), .A1(mai_mai_n1553_), .B0(mai_mai_n272_), .Y(mai_mai_n1555_));
  NA3        m1506(.A(mai_mai_n57_), .B(x4), .C(x3), .Y(mai_mai_n1556_));
  NO3        m1507(.A(mai_mai_n1556_), .B(mai_mai_n688_), .C(mai_mai_n133_), .Y(mai_mai_n1557_));
  INV        m1508(.A(mai_mai_n1557_), .Y(mai_mai_n1558_));
  NA4        m1509(.A(mai_mai_n1558_), .B(mai_mai_n1555_), .C(mai_mai_n1550_), .D(mai_mai_n1547_), .Y(mai24));
  NO2        m1510(.A(mai_mai_n221_), .B(x1), .Y(mai_mai_n1560_));
  NA2        m1511(.A(mai_mai_n313_), .B(mai_mai_n454_), .Y(mai_mai_n1561_));
  NO3        m1512(.A(mai_mai_n960_), .B(mai_mai_n1164_), .C(mai_mai_n941_), .Y(mai_mai_n1562_));
  AOI210     m1513(.A0(mai_mai_n880_), .A1(mai_mai_n56_), .B0(mai_mai_n1258_), .Y(mai_mai_n1563_));
  AN2        m1514(.A(mai_mai_n1563_), .B(mai_mai_n1562_), .Y(mai_mai_n1564_));
  NA2        m1515(.A(mai_mai_n1564_), .B(mai_mai_n923_), .Y(mai_mai_n1565_));
  INV        m1516(.A(mai_mai_n1565_), .Y(mai25));
  NA2        m1517(.A(mai_mai_n302_), .B(mai_mai_n59_), .Y(mai_mai_n1567_));
  NO2        m1518(.A(mai_mai_n687_), .B(mai_mai_n55_), .Y(mai_mai_n1568_));
  NA2        m1519(.A(mai_mai_n1568_), .B(mai_mai_n327_), .Y(mai_mai_n1569_));
  NO2        m1520(.A(mai_mai_n1569_), .B(mai_mai_n625_), .Y(mai_mai_n1570_));
  NO2        m1521(.A(mai_mai_n1206_), .B(mai_mai_n416_), .Y(mai_mai_n1571_));
  NO3        m1522(.A(mai_mai_n1571_), .B(mai_mai_n493_), .C(mai_mai_n98_), .Y(mai_mai_n1572_));
  NA2        m1523(.A(mai_mai_n471_), .B(mai_mai_n55_), .Y(mai_mai_n1573_));
  OAI220     m1524(.A0(mai_mai_n1573_), .A1(mai_mai_n221_), .B0(mai_mai_n540_), .B1(mai_mai_n250_), .Y(mai_mai_n1574_));
  OAI210     m1525(.A0(mai_mai_n1574_), .A1(mai_mai_n1572_), .B0(mai_mai_n582_), .Y(mai_mai_n1575_));
  INV        m1526(.A(mai_mai_n1575_), .Y(mai_mai_n1576_));
  AO210      m1527(.A0(mai_mai_n1576_), .A1(mai_mai_n103_), .B0(mai_mai_n1570_), .Y(mai26));
  NA2        m1528(.A(mai_mai_n573_), .B(mai_mai_n532_), .Y(mai_mai_n1578_));
  OAI210     m1529(.A0(mai_mai_n578_), .A1(mai_mai_n573_), .B0(mai_mai_n690_), .Y(mai_mai_n1579_));
  NO2        m1530(.A(mai_mai_n1064_), .B(mai_mai_n1579_), .Y(mai_mai_n1580_));
  NA2        m1531(.A(mai_mai_n914_), .B(mai_mai_n538_), .Y(mai_mai_n1581_));
  NA2        m1532(.A(mai_mai_n1531_), .B(mai_mai_n1265_), .Y(mai_mai_n1582_));
  NO2        m1533(.A(mai_mai_n973_), .B(mai_mai_n75_), .Y(mai_mai_n1583_));
  NA2        m1534(.A(mai_mai_n749_), .B(mai_mai_n167_), .Y(mai_mai_n1584_));
  NO2        m1535(.A(mai_mai_n1584_), .B(mai_mai_n498_), .Y(mai_mai_n1585_));
  AOI210     m1536(.A0(mai_mai_n1583_), .A1(mai_mai_n539_), .B0(mai_mai_n1585_), .Y(mai_mai_n1586_));
  OAI220     m1537(.A0(mai_mai_n1586_), .A1(mai_mai_n103_), .B0(mai_mai_n1582_), .B1(mai_mai_n53_), .Y(mai_mai_n1587_));
  NA2        m1538(.A(mai_mai_n553_), .B(mai_mai_n471_), .Y(mai_mai_n1588_));
  NO2        m1539(.A(mai_mai_n126_), .B(mai_mai_n124_), .Y(mai_mai_n1589_));
  NA2        m1540(.A(mai_mai_n1589_), .B(mai_mai_n117_), .Y(mai_mai_n1590_));
  NA2        m1541(.A(mai_mai_n690_), .B(x3), .Y(mai_mai_n1591_));
  AOI210     m1542(.A0(mai_mai_n1590_), .A1(mai_mai_n1588_), .B0(mai_mai_n1591_), .Y(mai_mai_n1592_));
  NO2        m1543(.A(mai_mai_n901_), .B(x3), .Y(mai_mai_n1593_));
  NO4        m1544(.A(x0), .B(mai_mai_n1592_), .C(mai_mai_n1587_), .D(mai_mai_n1580_), .Y(mai_mai_n1594_));
  AOI210     m1545(.A0(x8), .A1(x6), .B0(x5), .Y(mai_mai_n1595_));
  AO220      m1546(.A0(mai_mai_n1595_), .A1(mai_mai_n136_), .B0(mai_mai_n546_), .B1(mai_mai_n133_), .Y(mai_mai_n1596_));
  NA2        m1547(.A(mai_mai_n1596_), .B(mai_mai_n415_), .Y(mai_mai_n1597_));
  NA3        m1548(.A(mai_mai_n348_), .B(mai_mai_n784_), .C(mai_mai_n231_), .Y(mai_mai_n1598_));
  NA2        m1549(.A(mai_mai_n1598_), .B(mai_mai_n1597_), .Y(mai_mai_n1599_));
  AOI210     m1550(.A0(mai_mai_n205_), .A1(x2), .B0(mai_mai_n455_), .Y(mai_mai_n1600_));
  NO2        m1551(.A(mai_mai_n1600_), .B(mai_mai_n112_), .Y(mai_mai_n1601_));
  NO2        m1552(.A(mai_mai_n590_), .B(mai_mai_n630_), .Y(mai_mai_n1602_));
  NO2        m1553(.A(mai_mai_n1602_), .B(mai_mai_n1601_), .Y(mai_mai_n1603_));
  OAI210     m1554(.A0(mai_mai_n1603_), .A1(mai_mai_n53_), .B0(x0), .Y(mai_mai_n1604_));
  AOI210     m1555(.A0(mai_mai_n1599_), .A1(x4), .B0(mai_mai_n1604_), .Y(mai_mai_n1605_));
  OR2        m1556(.A(mai_mai_n1605_), .B(mai_mai_n1594_), .Y(mai27));
  NA2        m1557(.A(mai_mai_n1014_), .B(mai_mai_n414_), .Y(mai_mai_n1607_));
  NO2        m1558(.A(mai_mai_n1607_), .B(mai_mai_n273_), .Y(mai_mai_n1608_));
  NA3        m1559(.A(mai_mai_n757_), .B(mai_mai_n337_), .C(mai_mai_n916_), .Y(mai_mai_n1609_));
  NO2        m1560(.A(mai_mai_n1609_), .B(mai_mai_n199_), .Y(mai_mai_n1610_));
  OAI210     m1561(.A0(mai_mai_n1610_), .A1(mai_mai_n1608_), .B0(mai_mai_n646_), .Y(mai_mai_n1611_));
  XO2        m1562(.A(x8), .B(x4), .Y(mai_mai_n1612_));
  NO2        m1563(.A(mai_mai_n368_), .B(mai_mai_n154_), .Y(mai_mai_n1613_));
  NA2        m1564(.A(mai_mai_n1613_), .B(x7), .Y(mai_mai_n1614_));
  AOI210     m1565(.A0(mai_mai_n578_), .A1(mai_mai_n56_), .B0(mai_mai_n1583_), .Y(mai_mai_n1615_));
  OAI220     m1566(.A0(mai_mai_n1615_), .A1(mai_mai_n1094_), .B0(mai_mai_n1063_), .B1(mai_mai_n190_), .Y(mai_mai_n1616_));
  INV        m1567(.A(mai_mai_n643_), .Y(mai_mai_n1617_));
  NO2        m1568(.A(mai_mai_n1049_), .B(mai_mai_n234_), .Y(mai_mai_n1618_));
  AOI220     m1569(.A0(mai_mai_n1618_), .A1(mai_mai_n1617_), .B0(mai_mai_n1616_), .B1(mai_mai_n497_), .Y(mai_mai_n1619_));
  NA3        m1570(.A(mai_mai_n1619_), .B(mai_mai_n1614_), .C(mai_mai_n1611_), .Y(mai28));
  NA2        m1571(.A(mai_mai_n1110_), .B(mai_mai_n538_), .Y(mai_mai_n1621_));
  NA3        m1572(.A(mai_mai_n1045_), .B(mai_mai_n814_), .C(x7), .Y(mai_mai_n1622_));
  NA2        m1573(.A(mai_mai_n1622_), .B(mai_mai_n1621_), .Y(mai_mai_n1623_));
  NA2        m1574(.A(mai_mai_n1091_), .B(mai_mai_n413_), .Y(mai_mai_n1624_));
  NO4        m1575(.A(x6), .B(mai_mai_n56_), .C(x2), .D(x0), .Y(mai_mai_n1625_));
  NO2        m1576(.A(mai_mai_n361_), .B(x7), .Y(mai_mai_n1626_));
  INV        m1577(.A(mai_mai_n81_), .Y(mai_mai_n1627_));
  OAI210     m1578(.A0(mai_mai_n1626_), .A1(mai_mai_n106_), .B0(mai_mai_n1627_), .Y(mai_mai_n1628_));
  NA2        m1579(.A(mai_mai_n1536_), .B(mai_mai_n601_), .Y(mai_mai_n1629_));
  NO2        m1580(.A(mai_mai_n1573_), .B(mai_mai_n77_), .Y(mai_mai_n1630_));
  NA2        m1581(.A(mai_mai_n1630_), .B(mai_mai_n1629_), .Y(mai_mai_n1631_));
  AOI210     m1582(.A0(mai_mai_n1631_), .A1(mai_mai_n1628_), .B0(mai_mai_n59_), .Y(mai_mai_n1632_));
  NA2        m1583(.A(mai_mai_n385_), .B(mai_mai_n423_), .Y(mai_mai_n1633_));
  OAI210     m1584(.A0(mai_mai_n1633_), .A1(mai_mai_n135_), .B0(x1), .Y(mai_mai_n1634_));
  NO2        m1585(.A(mai_mai_n1634_), .B(mai_mai_n1632_), .Y(mai_mai_n1635_));
  NOi21      m1586(.An(mai_mai_n651_), .B(mai_mai_n894_), .Y(mai_mai_n1636_));
  INV        m1587(.A(mai_mai_n971_), .Y(mai_mai_n1637_));
  OAI210     m1588(.A0(mai_mai_n1178_), .A1(mai_mai_n1443_), .B0(mai_mai_n1637_), .Y(mai_mai_n1638_));
  NA2        m1589(.A(mai_mai_n1638_), .B(x7), .Y(mai_mai_n1639_));
  OAI210     m1590(.A0(mai_mai_n413_), .A1(mai_mai_n51_), .B0(mai_mai_n910_), .Y(mai_mai_n1640_));
  AOI220     m1591(.A0(mai_mai_n1640_), .A1(mai_mai_n429_), .B0(mai_mai_n413_), .B1(mai_mai_n362_), .Y(mai_mai_n1641_));
  NO2        m1592(.A(mai_mai_n1641_), .B(mai_mai_n143_), .Y(mai_mai_n1642_));
  NA2        m1593(.A(mai_mai_n152_), .B(mai_mai_n71_), .Y(mai_mai_n1643_));
  OAI210     m1594(.A0(mai_mai_n1581_), .A1(mai_mai_n1643_), .B0(mai_mai_n53_), .Y(mai_mai_n1644_));
  OAI220     m1595(.A0(mai_mai_n631_), .A1(mai_mai_n239_), .B0(mai_mai_n627_), .B1(x6), .Y(mai_mai_n1645_));
  NO2        m1596(.A(mai_mai_n275_), .B(x4), .Y(mai_mai_n1646_));
  AOI220     m1597(.A0(mai_mai_n1646_), .A1(mai_mai_n337_), .B0(mai_mai_n1645_), .B1(x4), .Y(mai_mai_n1647_));
  NO3        m1598(.A(mai_mai_n1647_), .B(mai_mai_n296_), .C(x5), .Y(mai_mai_n1648_));
  NA2        m1599(.A(mai_mai_n1617_), .B(mai_mai_n414_), .Y(mai_mai_n1649_));
  NO2        m1600(.A(mai_mai_n1649_), .B(mai_mai_n234_), .Y(mai_mai_n1650_));
  NO4        m1601(.A(mai_mai_n1650_), .B(mai_mai_n1648_), .C(mai_mai_n1644_), .D(mai_mai_n1642_), .Y(mai_mai_n1651_));
  AOI210     m1602(.A0(mai_mai_n1651_), .A1(mai_mai_n1639_), .B0(mai_mai_n1635_), .Y(mai_mai_n1652_));
  AOI210     m1603(.A0(mai_mai_n1623_), .A1(x3), .B0(mai_mai_n1652_), .Y(mai29));
  OAI210     m1604(.A0(mai_mai_n514_), .A1(mai_mai_n240_), .B0(mai_mai_n674_), .Y(mai_mai_n1654_));
  NA2        m1605(.A(mai_mai_n692_), .B(mai_mai_n939_), .Y(mai_mai_n1655_));
  AO210      m1606(.A0(mai_mai_n1025_), .A1(mai_mai_n1034_), .B0(mai_mai_n1655_), .Y(mai_mai_n1656_));
  AOI210     m1607(.A0(mai_mai_n172_), .A1(mai_mai_n156_), .B0(mai_mai_n651_), .Y(mai_mai_n1657_));
  INV        m1608(.A(mai_mai_n1657_), .Y(mai_mai_n1658_));
  NA3        m1609(.A(mai_mai_n1658_), .B(mai_mai_n1656_), .C(mai_mai_n1654_), .Y(mai_mai_n1659_));
  NO2        m1610(.A(mai_mai_n411_), .B(mai_mai_n58_), .Y(mai_mai_n1660_));
  NA2        m1611(.A(mai_mai_n1660_), .B(mai_mai_n1064_), .Y(mai_mai_n1661_));
  OAI210     m1612(.A0(mai_mai_n133_), .A1(mai_mai_n502_), .B0(mai_mai_n1661_), .Y(mai_mai_n1662_));
  AOI210     m1613(.A0(mai_mai_n1659_), .A1(x6), .B0(mai_mai_n1662_), .Y(mai_mai_n1663_));
  OAI210     m1614(.A0(x8), .A1(x4), .B0(x5), .Y(mai_mai_n1664_));
  NA2        m1615(.A(mai_mai_n1664_), .B(mai_mai_n107_), .Y(mai_mai_n1665_));
  NA4        m1616(.A(x6), .B(mai_mai_n1665_), .C(mai_mai_n610_), .D(mai_mai_n64_), .Y(mai_mai_n1666_));
  AOI210     m1617(.A0(mai_mai_n1145_), .A1(mai_mai_n248_), .B0(mai_mai_n1486_), .Y(mai_mai_n1667_));
  AOI210     m1618(.A0(mai_mai_n1667_), .A1(mai_mai_n1666_), .B0(mai_mai_n811_), .Y(mai_mai_n1668_));
  NA3        m1619(.A(mai_mai_n611_), .B(mai_mai_n280_), .C(mai_mai_n156_), .Y(mai_mai_n1669_));
  NA3        m1620(.A(mai_mai_n577_), .B(mai_mai_n270_), .C(mai_mai_n740_), .Y(mai_mai_n1670_));
  AOI210     m1621(.A0(mai_mai_n1670_), .A1(mai_mai_n1669_), .B0(mai_mai_n1064_), .Y(mai_mai_n1671_));
  NA2        m1622(.A(x8), .B(x7), .Y(mai_mai_n1672_));
  NO2        m1623(.A(mai_mai_n1672_), .B(mai_mai_n122_), .Y(mai_mai_n1673_));
  OAI220     m1624(.A0(mai_mai_n1664_), .A1(mai_mai_n540_), .B0(mai_mai_n1299_), .B1(mai_mai_n368_), .Y(mai_mai_n1674_));
  NO4        m1625(.A(mai_mai_n1674_), .B(mai_mai_n1673_), .C(mai_mai_n1671_), .D(mai_mai_n1668_), .Y(mai_mai_n1675_));
  OAI210     m1626(.A0(mai_mai_n1663_), .A1(x2), .B0(mai_mai_n1675_), .Y(mai_mai_n1676_));
  NA3        m1627(.A(x6), .B(mai_mai_n50_), .C(x2), .Y(mai_mai_n1677_));
  OAI210     m1628(.A0(mai_mai_n1073_), .A1(mai_mai_n327_), .B0(mai_mai_n1677_), .Y(mai_mai_n1678_));
  NA2        m1629(.A(mai_mai_n1678_), .B(mai_mai_n317_), .Y(mai_mai_n1679_));
  NO3        m1630(.A(mai_mai_n644_), .B(mai_mai_n338_), .C(mai_mai_n134_), .Y(mai_mai_n1680_));
  AOI210     m1631(.A0(mai_mai_n673_), .A1(mai_mai_n564_), .B0(mai_mai_n1680_), .Y(mai_mai_n1681_));
  OAI210     m1632(.A0(mai_mai_n1679_), .A1(x7), .B0(mai_mai_n1681_), .Y(mai_mai_n1682_));
  AOI210     m1633(.A0(mai_mai_n975_), .A1(mai_mai_n373_), .B0(mai_mai_n1216_), .Y(mai_mai_n1683_));
  NO2        m1634(.A(mai_mai_n138_), .B(x2), .Y(mai_mai_n1684_));
  OA210      m1635(.A0(mai_mai_n1684_), .A1(mai_mai_n575_), .B0(mai_mai_n611_), .Y(mai_mai_n1685_));
  OAI210     m1636(.A0(mai_mai_n1685_), .A1(mai_mai_n1683_), .B0(mai_mai_n68_), .Y(mai_mai_n1686_));
  NO2        m1637(.A(mai_mai_n184_), .B(mai_mai_n85_), .Y(mai_mai_n1687_));
  OAI210     m1638(.A0(mai_mai_n1687_), .A1(mai_mai_n727_), .B0(mai_mai_n979_), .Y(mai_mai_n1688_));
  NA2        m1639(.A(mai_mai_n1688_), .B(mai_mai_n1686_), .Y(mai_mai_n1689_));
  AOI210     m1640(.A0(mai_mai_n1682_), .A1(x8), .B0(mai_mai_n1689_), .Y(mai_mai_n1690_));
  OAI210     m1641(.A0(mai_mai_n411_), .A1(mai_mai_n226_), .B0(mai_mai_n872_), .Y(mai_mai_n1691_));
  OAI210     m1642(.A0(mai_mai_n1691_), .A1(mai_mai_n994_), .B0(mai_mai_n620_), .Y(mai_mai_n1692_));
  NO2        m1643(.A(mai_mai_n127_), .B(mai_mai_n93_), .Y(mai_mai_n1693_));
  NA2        m1644(.A(mai_mai_n1693_), .B(mai_mai_n541_), .Y(mai_mai_n1694_));
  NA2        m1645(.A(mai_mai_n1694_), .B(mai_mai_n1692_), .Y(mai_mai_n1695_));
  NO3        m1646(.A(mai_mai_n1058_), .B(mai_mai_n463_), .C(mai_mai_n103_), .Y(mai_mai_n1696_));
  NA2        m1647(.A(mai_mai_n1696_), .B(mai_mai_n105_), .Y(mai_mai_n1697_));
  AOI210     m1648(.A0(mai_mai_n279_), .A1(x4), .B0(mai_mai_n178_), .Y(mai_mai_n1698_));
  OAI210     m1649(.A0(mai_mai_n1698_), .A1(mai_mai_n1660_), .B0(mai_mai_n669_), .Y(mai_mai_n1699_));
  OR3        m1650(.A(mai_mai_n1505_), .B(mai_mai_n1234_), .C(mai_mai_n972_), .Y(mai_mai_n1700_));
  NA2        m1651(.A(mai_mai_n1625_), .B(mai_mai_n746_), .Y(mai_mai_n1701_));
  NA3        m1652(.A(mai_mai_n1700_), .B(mai_mai_n1699_), .C(mai_mai_n1697_), .Y(mai_mai_n1702_));
  AOI210     m1653(.A0(mai_mai_n1695_), .A1(mai_mai_n266_), .B0(mai_mai_n1702_), .Y(mai_mai_n1703_));
  OAI210     m1654(.A0(mai_mai_n1690_), .A1(x1), .B0(mai_mai_n1703_), .Y(mai_mai_n1704_));
  AO210      m1655(.A0(mai_mai_n1676_), .A1(x1), .B0(mai_mai_n1704_), .Y(mai30));
  NO3        m1656(.A(mai_mai_n1526_), .B(mai_mai_n530_), .C(mai_mai_n98_), .Y(mai_mai_n1706_));
  NO3        m1657(.A(mai_mai_n1008_), .B(mai_mai_n130_), .C(mai_mai_n358_), .Y(mai_mai_n1707_));
  AOI210     m1658(.A0(mai_mai_n669_), .A1(mai_mai_n231_), .B0(mai_mai_n1707_), .Y(mai_mai_n1708_));
  AOI210     m1659(.A0(mai_mai_n1708_), .A1(mai_mai_n1706_), .B0(mai_mai_n56_), .Y(mai_mai_n1709_));
  NA2        m1660(.A(mai_mai_n751_), .B(mai_mai_n315_), .Y(mai_mai_n1710_));
  INV        m1661(.A(mai_mai_n1710_), .Y(mai_mai_n1711_));
  OAI210     m1662(.A0(mai_mai_n1711_), .A1(mai_mai_n1709_), .B0(mai_mai_n105_), .Y(mai_mai_n1712_));
  OAI210     m1663(.A0(mai_mai_n894_), .A1(mai_mai_n525_), .B0(mai_mai_n620_), .Y(mai_mai_n1713_));
  AOI220     m1664(.A0(mai_mai_n415_), .A1(mai_mai_n850_), .B0(mai_mai_n301_), .B1(mai_mai_n423_), .Y(mai_mai_n1714_));
  AOI210     m1665(.A0(mai_mai_n1714_), .A1(mai_mai_n1713_), .B0(mai_mai_n234_), .Y(mai_mai_n1715_));
  NO2        m1666(.A(mai_mai_n119_), .B(x0), .Y(mai_mai_n1716_));
  AOI210     m1667(.A0(mai_mai_n465_), .A1(x6), .B0(mai_mai_n1716_), .Y(mai_mai_n1717_));
  NO2        m1668(.A(mai_mai_n1717_), .B(mai_mai_n54_), .Y(mai_mai_n1718_));
  NA2        m1669(.A(mai_mai_n153_), .B(mai_mai_n71_), .Y(mai_mai_n1719_));
  AO210      m1670(.A0(mai_mai_n524_), .A1(mai_mai_n479_), .B0(x5), .Y(mai_mai_n1720_));
  AOI210     m1671(.A0(mai_mai_n1719_), .A1(mai_mai_n667_), .B0(mai_mai_n1720_), .Y(mai_mai_n1721_));
  AOI210     m1672(.A0(mai_mai_n1379_), .A1(mai_mai_n50_), .B0(mai_mai_n423_), .Y(mai_mai_n1722_));
  NA2        m1673(.A(mai_mai_n183_), .B(x2), .Y(mai_mai_n1723_));
  OA220      m1674(.A0(mai_mai_n1723_), .A1(mai_mai_n1722_), .B0(mai_mai_n251_), .B1(x6), .Y(mai_mai_n1724_));
  OAI210     m1675(.A0(x7), .A1(x6), .B0(x1), .Y(mai_mai_n1725_));
  NA3        m1676(.A(mai_mai_n57_), .B(x4), .C(mai_mai_n59_), .Y(mai_mai_n1726_));
  AOI220     m1677(.A0(mai_mai_n1726_), .A1(mai_mai_n1184_), .B0(mai_mai_n1725_), .B1(mai_mai_n1556_), .Y(mai_mai_n1727_));
  NO3        m1678(.A(mai_mai_n1181_), .B(mai_mai_n317_), .C(mai_mai_n916_), .Y(mai_mai_n1728_));
  NO3        m1679(.A(mai_mai_n1127_), .B(mai_mai_n212_), .C(mai_mai_n593_), .Y(mai_mai_n1729_));
  NO3        m1680(.A(mai_mai_n1729_), .B(mai_mai_n1728_), .C(mai_mai_n1727_), .Y(mai_mai_n1730_));
  OAI210     m1681(.A0(mai_mai_n1724_), .A1(mai_mai_n698_), .B0(mai_mai_n1730_), .Y(mai_mai_n1731_));
  NO4        m1682(.A(mai_mai_n1731_), .B(mai_mai_n1721_), .C(mai_mai_n1718_), .D(mai_mai_n1715_), .Y(mai_mai_n1732_));
  AOI210     m1683(.A0(mai_mai_n1732_), .A1(mai_mai_n1712_), .B0(x8), .Y(mai_mai_n1733_));
  NO3        m1684(.A(mai_mai_n453_), .B(mai_mai_n724_), .C(mai_mai_n53_), .Y(mai_mai_n1734_));
  OAI220     m1685(.A0(mai_mai_n1534_), .A1(mai_mai_n317_), .B0(mai_mai_n446_), .B1(mai_mai_n537_), .Y(mai_mai_n1735_));
  OAI210     m1686(.A0(mai_mai_n1735_), .A1(mai_mai_n1734_), .B0(x6), .Y(mai_mai_n1736_));
  OAI210     m1687(.A0(mai_mai_n930_), .A1(mai_mai_n497_), .B0(mai_mai_n751_), .Y(mai_mai_n1737_));
  OAI210     m1688(.A0(mai_mai_n1496_), .A1(mai_mai_n304_), .B0(mai_mai_n121_), .Y(mai_mai_n1738_));
  AOI210     m1689(.A0(mai_mai_n353_), .A1(mai_mai_n209_), .B0(mai_mai_n72_), .Y(mai_mai_n1739_));
  AOI210     m1690(.A0(mai_mai_n894_), .A1(mai_mai_n690_), .B0(mai_mai_n1739_), .Y(mai_mai_n1740_));
  NA4        m1691(.A(mai_mai_n1740_), .B(mai_mai_n1738_), .C(mai_mai_n1737_), .D(mai_mai_n1736_), .Y(mai_mai_n1741_));
  NA2        m1692(.A(mai_mai_n1741_), .B(x8), .Y(mai_mai_n1742_));
  NO2        m1693(.A(mai_mai_n1742_), .B(mai_mai_n57_), .Y(mai_mai_n1743_));
  NA2        m1694(.A(mai_mai_n402_), .B(mai_mai_n774_), .Y(mai_mai_n1744_));
  INV        m1695(.A(mai_mai_n607_), .Y(mai_mai_n1745_));
  AOI210     m1696(.A0(mai_mai_n1745_), .A1(mai_mai_n1744_), .B0(mai_mai_n413_), .Y(mai_mai_n1746_));
  NO3        m1697(.A(mai_mai_n582_), .B(mai_mai_n382_), .C(mai_mai_n1008_), .Y(mai_mai_n1747_));
  NO2        m1698(.A(mai_mai_n1747_), .B(mai_mai_n1094_), .Y(mai_mai_n1748_));
  NO2        m1699(.A(mai_mai_n282_), .B(x5), .Y(mai_mai_n1749_));
  INV        m1700(.A(mai_mai_n781_), .Y(mai_mai_n1750_));
  NO2        m1701(.A(mai_mai_n1750_), .B(mai_mai_n950_), .Y(mai_mai_n1751_));
  NO3        m1702(.A(mai_mai_n1751_), .B(mai_mai_n1748_), .C(mai_mai_n1746_), .Y(mai_mai_n1752_));
  NA2        m1703(.A(mai_mai_n870_), .B(mai_mai_n82_), .Y(mai_mai_n1753_));
  AO210      m1704(.A0(mai_mai_n1753_), .A1(mai_mai_n1380_), .B0(x3), .Y(mai_mai_n1754_));
  NO2        m1705(.A(mai_mai_n202_), .B(mai_mai_n56_), .Y(mai_mai_n1755_));
  OAI220     m1706(.A0(mai_mai_n353_), .A1(mai_mai_n1094_), .B0(mai_mai_n328_), .B1(mai_mai_n212_), .Y(mai_mai_n1756_));
  AOI220     m1707(.A0(mai_mai_n1756_), .A1(x2), .B0(mai_mai_n1755_), .B1(mai_mai_n1393_), .Y(mai_mai_n1757_));
  AOI210     m1708(.A0(mai_mai_n1757_), .A1(mai_mai_n1754_), .B0(mai_mai_n239_), .Y(mai_mai_n1758_));
  NO3        m1709(.A(mai_mai_n756_), .B(mai_mai_n645_), .C(mai_mai_n156_), .Y(mai_mai_n1759_));
  NA2        m1710(.A(mai_mai_n1759_), .B(mai_mai_n144_), .Y(mai_mai_n1760_));
  NA3        m1711(.A(x5), .B(x4), .C(mai_mai_n59_), .Y(mai_mai_n1761_));
  AOI210     m1712(.A0(mai_mai_n1761_), .A1(mai_mai_n1135_), .B0(mai_mai_n498_), .Y(mai_mai_n1762_));
  AOI210     m1713(.A0(mai_mai_n1152_), .A1(x2), .B0(mai_mai_n1762_), .Y(mai_mai_n1763_));
  AOI210     m1714(.A0(mai_mai_n1763_), .A1(mai_mai_n1760_), .B0(mai_mai_n50_), .Y(mai_mai_n1764_));
  NA2        m1715(.A(mai_mai_n1275_), .B(mai_mai_n1004_), .Y(mai_mai_n1765_));
  AOI210     m1716(.A0(mai_mai_n1765_), .A1(mai_mai_n1753_), .B0(mai_mai_n561_), .Y(mai_mai_n1766_));
  AOI210     m1717(.A0(mai_mai_n916_), .A1(x1), .B0(mai_mai_n1145_), .Y(mai_mai_n1767_));
  OAI220     m1718(.A0(mai_mai_n280_), .A1(x4), .B0(mai_mai_n51_), .B1(x6), .Y(mai_mai_n1768_));
  NO2        m1719(.A(mai_mai_n117_), .B(mai_mai_n107_), .Y(mai_mai_n1769_));
  AOI220     m1720(.A0(mai_mai_n1769_), .A1(mai_mai_n1768_), .B0(mai_mai_n1027_), .B1(mai_mai_n572_), .Y(mai_mai_n1770_));
  OAI210     m1721(.A0(mai_mai_n1767_), .A1(mai_mai_n448_), .B0(mai_mai_n1770_), .Y(mai_mai_n1771_));
  NO4        m1722(.A(mai_mai_n1771_), .B(mai_mai_n1766_), .C(mai_mai_n1764_), .D(mai_mai_n1758_), .Y(mai_mai_n1772_));
  OAI210     m1723(.A0(mai_mai_n1752_), .A1(mai_mai_n127_), .B0(mai_mai_n1772_), .Y(mai_mai_n1773_));
  NO3        m1724(.A(mai_mai_n1773_), .B(mai_mai_n1743_), .C(mai_mai_n1733_), .Y(mai31));
  NA2        m1725(.A(mai_mai_n880_), .B(mai_mai_n329_), .Y(mai_mai_n1775_));
  NO2        m1726(.A(mai_mai_n416_), .B(mai_mai_n620_), .Y(mai_mai_n1776_));
  AOI210     m1727(.A0(mai_mai_n1776_), .A1(mai_mai_n1775_), .B0(mai_mai_n58_), .Y(mai_mai_n1777_));
  NO2        m1728(.A(mai_mai_n726_), .B(mai_mai_n56_), .Y(mai_mai_n1778_));
  AOI220     m1729(.A0(mai_mai_n1778_), .A1(x2), .B0(mai_mai_n91_), .B1(x0), .Y(mai_mai_n1779_));
  NA3        m1730(.A(mai_mai_n1779_), .B(mai_mai_n1701_), .C(mai_mai_n1578_), .Y(mai_mai_n1780_));
  OAI210     m1731(.A0(mai_mai_n1780_), .A1(mai_mai_n1777_), .B0(mai_mai_n53_), .Y(mai_mai_n1781_));
  NO2        m1732(.A(mai_mai_n400_), .B(mai_mai_n620_), .Y(mai_mai_n1782_));
  NO2        m1733(.A(mai_mai_n1625_), .B(mai_mai_n812_), .Y(mai_mai_n1783_));
  OA220      m1734(.A0(mai_mai_n1783_), .A1(mai_mai_n443_), .B0(mai_mai_n1782_), .B1(mai_mai_n1268_), .Y(mai_mai_n1784_));
  AOI210     m1735(.A0(mai_mai_n1784_), .A1(mai_mai_n1781_), .B0(mai_mai_n103_), .Y(mai_mai_n1785_));
  NO2        m1736(.A(mai_mai_n459_), .B(mai_mai_n75_), .Y(mai_mai_n1786_));
  NA2        m1737(.A(mai_mai_n413_), .B(mai_mai_n57_), .Y(mai_mai_n1787_));
  AOI210     m1738(.A0(mai_mai_n279_), .A1(mai_mai_n86_), .B0(mai_mai_n1787_), .Y(mai_mai_n1788_));
  OAI210     m1739(.A0(mai_mai_n1788_), .A1(mai_mai_n1786_), .B0(mai_mai_n713_), .Y(mai_mai_n1789_));
  NO4        m1740(.A(mai_mai_n1023_), .B(mai_mai_n338_), .C(mai_mai_n1379_), .D(mai_mai_n67_), .Y(mai_mai_n1790_));
  AOI210     m1741(.A0(mai_mai_n1416_), .A1(mai_mai_n1172_), .B0(mai_mai_n411_), .Y(mai_mai_n1791_));
  NO2        m1742(.A(mai_mai_n1791_), .B(mai_mai_n1790_), .Y(mai_mai_n1792_));
  AOI210     m1743(.A0(mai_mai_n1792_), .A1(mai_mai_n1789_), .B0(x5), .Y(mai_mai_n1793_));
  NO2        m1744(.A(mai_mai_n533_), .B(mai_mai_n1073_), .Y(mai_mai_n1794_));
  AOI220     m1745(.A0(mai_mai_n871_), .A1(mai_mai_n679_), .B0(mai_mai_n1008_), .B1(mai_mai_n116_), .Y(mai_mai_n1795_));
  NO2        m1746(.A(mai_mai_n1795_), .B(mai_mai_n361_), .Y(mai_mai_n1796_));
  NO4        m1747(.A(mai_mai_n1796_), .B(mai_mai_n1794_), .C(mai_mai_n1793_), .D(mai_mai_n1785_), .Y(mai_mai_n1797_));
  INV        m1748(.A(mai_mai_n133_), .Y(mai_mai_n1798_));
  NA2        m1749(.A(mai_mai_n1798_), .B(x7), .Y(mai_mai_n1799_));
  NO3        m1750(.A(mai_mai_n353_), .B(mai_mai_n55_), .C(x7), .Y(mai_mai_n1800_));
  OA210      m1751(.A0(mai_mai_n1800_), .A1(mai_mai_n1144_), .B0(mai_mai_n99_), .Y(mai_mai_n1801_));
  NA2        m1752(.A(mai_mai_n973_), .B(mai_mai_n92_), .Y(mai_mai_n1802_));
  AOI210     m1753(.A0(mai_mai_n820_), .A1(mai_mai_n107_), .B0(mai_mai_n1802_), .Y(mai_mai_n1803_));
  NA2        m1754(.A(mai_mai_n1335_), .B(x6), .Y(mai_mai_n1804_));
  AOI210     m1755(.A0(mai_mai_n1804_), .A1(mai_mai_n265_), .B0(mai_mai_n103_), .Y(mai_mai_n1805_));
  NA2        m1756(.A(mai_mai_n1045_), .B(mai_mai_n292_), .Y(mai_mai_n1806_));
  AOI210     m1757(.A0(mai_mai_n1806_), .A1(mai_mai_n590_), .B0(mai_mai_n53_), .Y(mai_mai_n1807_));
  NO4        m1758(.A(mai_mai_n1807_), .B(mai_mai_n1805_), .C(mai_mai_n1803_), .D(mai_mai_n1801_), .Y(mai_mai_n1808_));
  AOI210     m1759(.A0(mai_mai_n1808_), .A1(mai_mai_n1799_), .B0(mai_mai_n630_), .Y(mai_mai_n1809_));
  NO4        m1760(.A(mai_mai_n565_), .B(mai_mai_n541_), .C(mai_mai_n646_), .D(mai_mai_n645_), .Y(mai_mai_n1810_));
  OAI210     m1761(.A0(mai_mai_n1810_), .A1(mai_mai_n968_), .B0(x3), .Y(mai_mai_n1811_));
  NO3        m1762(.A(x6), .B(mai_mai_n56_), .C(x1), .Y(mai_mai_n1812_));
  NA2        m1763(.A(mai_mai_n1812_), .B(mai_mai_n262_), .Y(mai_mai_n1813_));
  NA2        m1764(.A(mai_mai_n1607_), .B(mai_mai_n1813_), .Y(mai_mai_n1814_));
  NA4        m1765(.A(mai_mai_n582_), .B(mai_mai_n168_), .C(x6), .D(mai_mai_n103_), .Y(mai_mai_n1815_));
  NO2        m1766(.A(mai_mai_n782_), .B(mai_mai_n228_), .Y(mai_mai_n1816_));
  NOi31      m1767(.An(mai_mai_n1815_), .B(mai_mai_n1816_), .C(mai_mai_n1814_), .Y(mai_mai_n1817_));
  AOI210     m1768(.A0(mai_mai_n1817_), .A1(mai_mai_n1811_), .B0(mai_mai_n493_), .Y(mai_mai_n1818_));
  OAI210     m1769(.A0(mai_mai_n564_), .A1(mai_mai_n437_), .B0(mai_mai_n850_), .Y(mai_mai_n1819_));
  NO3        m1770(.A(mai_mai_n348_), .B(mai_mai_n77_), .C(mai_mai_n53_), .Y(mai_mai_n1820_));
  NO3        m1771(.A(mai_mai_n429_), .B(mai_mai_n323_), .C(mai_mai_n50_), .Y(mai_mai_n1821_));
  OAI210     m1772(.A0(mai_mai_n1821_), .A1(mai_mai_n1820_), .B0(mai_mai_n1024_), .Y(mai_mai_n1822_));
  AOI210     m1773(.A0(mai_mai_n1822_), .A1(mai_mai_n1819_), .B0(mai_mai_n366_), .Y(mai_mai_n1823_));
  NO2        m1774(.A(mai_mai_n199_), .B(mai_mai_n498_), .Y(mai_mai_n1824_));
  OAI210     m1775(.A0(mai_mai_n130_), .A1(x2), .B0(mai_mai_n1824_), .Y(mai_mai_n1825_));
  NA3        m1776(.A(mai_mai_n382_), .B(mai_mai_n302_), .C(mai_mai_n77_), .Y(mai_mai_n1826_));
  OA210      m1777(.A0(mai_mai_n225_), .A1(mai_mai_n208_), .B0(mai_mai_n1826_), .Y(mai_mai_n1827_));
  AOI210     m1778(.A0(mai_mai_n1827_), .A1(mai_mai_n1825_), .B0(mai_mai_n64_), .Y(mai_mai_n1828_));
  NA2        m1779(.A(mai_mai_n117_), .B(mai_mai_n57_), .Y(mai_mai_n1829_));
  AOI220     m1780(.A0(mai_mai_n1363_), .A1(mai_mai_n827_), .B0(mai_mai_n249_), .B1(x4), .Y(mai_mai_n1830_));
  AOI220     m1781(.A0(mai_mai_n1410_), .A1(mai_mai_n566_), .B0(mai_mai_n668_), .B1(mai_mai_n713_), .Y(mai_mai_n1831_));
  OAI220     m1782(.A0(mai_mai_n1831_), .A1(mai_mai_n1829_), .B0(mai_mai_n1830_), .B1(mai_mai_n176_), .Y(mai_mai_n1832_));
  OR3        m1783(.A(mai_mai_n1832_), .B(mai_mai_n1828_), .C(mai_mai_n1823_), .Y(mai_mai_n1833_));
  NO3        m1784(.A(mai_mai_n1833_), .B(mai_mai_n1818_), .C(mai_mai_n1809_), .Y(mai_mai_n1834_));
  OAI210     m1785(.A0(mai_mai_n1797_), .A1(x3), .B0(mai_mai_n1834_), .Y(mai32));
  NO2        m1786(.A(mai_mai_n1277_), .B(mai_mai_n50_), .Y(mai_mai_n1836_));
  NA3        m1787(.A(mai_mai_n1336_), .B(mai_mai_n741_), .C(mai_mai_n264_), .Y(mai_mai_n1837_));
  INV        m1788(.A(mai_mai_n688_), .Y(mai_mai_n1838_));
  NO2        m1789(.A(mai_mai_n1181_), .B(mai_mai_n537_), .Y(mai_mai_n1839_));
  NO2        m1790(.A(mai_mai_n1839_), .B(mai_mai_n1838_), .Y(mai_mai_n1840_));
  AOI210     m1791(.A0(mai_mai_n1840_), .A1(mai_mai_n1837_), .B0(mai_mai_n134_), .Y(mai_mai_n1841_));
  OAI220     m1792(.A0(mai_mai_n375_), .A1(x7), .B0(mai_mai_n275_), .B1(mai_mai_n270_), .Y(mai_mai_n1842_));
  NA2        m1793(.A(mai_mai_n1842_), .B(mai_mai_n870_), .Y(mai_mai_n1843_));
  NA2        m1794(.A(mai_mai_n490_), .B(mai_mai_n124_), .Y(mai_mai_n1844_));
  AOI210     m1795(.A0(mai_mai_n1844_), .A1(mai_mai_n1843_), .B0(mai_mai_n105_), .Y(mai_mai_n1845_));
  NA3        m1796(.A(mai_mai_n1144_), .B(mai_mai_n1010_), .C(mai_mai_n112_), .Y(mai_mai_n1846_));
  NA2        m1797(.A(mai_mai_n1173_), .B(mai_mai_n646_), .Y(mai_mai_n1847_));
  AOI210     m1798(.A0(mai_mai_n1847_), .A1(mai_mai_n1846_), .B0(mai_mai_n56_), .Y(mai_mai_n1848_));
  NA2        m1799(.A(mai_mai_n870_), .B(mai_mai_n57_), .Y(mai_mai_n1849_));
  NOi21      m1800(.An(mai_mai_n1849_), .B(mai_mai_n124_), .Y(mai_mai_n1850_));
  NO3        m1801(.A(mai_mai_n2217_), .B(mai_mai_n1850_), .C(mai_mai_n59_), .Y(mai_mai_n1851_));
  OR4        m1802(.A(mai_mai_n1851_), .B(mai_mai_n1848_), .C(mai_mai_n1845_), .D(mai_mai_n1841_), .Y(mai_mai_n1852_));
  OAI210     m1803(.A0(mai_mai_n1852_), .A1(mai_mai_n1836_), .B0(mai_mai_n103_), .Y(mai_mai_n1853_));
  NO3        m1804(.A(mai_mai_n1073_), .B(mai_mai_n136_), .C(mai_mai_n120_), .Y(mai_mai_n1854_));
  NO2        m1805(.A(mai_mai_n356_), .B(mai_mai_n55_), .Y(mai_mai_n1855_));
  NA2        m1806(.A(mai_mai_n1855_), .B(mai_mai_n111_), .Y(mai_mai_n1856_));
  INV        m1807(.A(mai_mai_n1856_), .Y(mai_mai_n1857_));
  OAI210     m1808(.A0(mai_mai_n1857_), .A1(mai_mai_n1854_), .B0(x3), .Y(mai_mai_n1858_));
  OAI210     m1809(.A0(mai_mai_n814_), .A1(mai_mai_n248_), .B0(mai_mai_n50_), .Y(mai_mai_n1859_));
  AOI210     m1810(.A0(mai_mai_n62_), .A1(mai_mai_n105_), .B0(mai_mai_n1859_), .Y(mai_mai_n1860_));
  OAI210     m1811(.A0(mai_mai_n1860_), .A1(mai_mai_n1583_), .B0(mai_mai_n645_), .Y(mai_mai_n1861_));
  NO3        m1812(.A(mai_mai_n741_), .B(mai_mai_n336_), .C(mai_mai_n134_), .Y(mai_mai_n1862_));
  NA2        m1813(.A(mai_mai_n1862_), .B(mai_mai_n59_), .Y(mai_mai_n1863_));
  NA2        m1814(.A(mai_mai_n1014_), .B(mai_mai_n71_), .Y(mai_mai_n1864_));
  NO2        m1815(.A(mai_mai_n1626_), .B(mai_mai_n543_), .Y(mai_mai_n1865_));
  NO2        m1816(.A(mai_mai_n1865_), .B(mai_mai_n1864_), .Y(mai_mai_n1866_));
  NO3        m1817(.A(mai_mai_n1137_), .B(mai_mai_n199_), .C(mai_mai_n234_), .Y(mai_mai_n1867_));
  NO3        m1818(.A(mai_mai_n1867_), .B(mai_mai_n1866_), .C(x1), .Y(mai_mai_n1868_));
  NA4        m1819(.A(mai_mai_n1868_), .B(mai_mai_n1863_), .C(mai_mai_n1861_), .D(mai_mai_n1858_), .Y(mai_mai_n1869_));
  OR2        m1820(.A(mai_mai_n370_), .B(mai_mai_n901_), .Y(mai_mai_n1870_));
  NA3        m1821(.A(mai_mai_n1612_), .B(mai_mai_n513_), .C(mai_mai_n250_), .Y(mai_mai_n1871_));
  AOI210     m1822(.A0(mai_mai_n1871_), .A1(mai_mai_n1870_), .B0(mai_mai_n277_), .Y(mai_mai_n1872_));
  NA3        m1823(.A(mai_mai_n1101_), .B(mai_mai_n487_), .C(mai_mai_n361_), .Y(mai_mai_n1873_));
  NO3        m1824(.A(mai_mai_n1234_), .B(mai_mai_n901_), .C(x2), .Y(mai_mai_n1874_));
  NO2        m1825(.A(mai_mai_n1091_), .B(mai_mai_n359_), .Y(mai_mai_n1875_));
  NO2        m1826(.A(mai_mai_n1567_), .B(mai_mai_n64_), .Y(mai_mai_n1876_));
  NO4        m1827(.A(mai_mai_n1876_), .B(mai_mai_n1875_), .C(mai_mai_n1874_), .D(mai_mai_n53_), .Y(mai_mai_n1877_));
  NO2        m1828(.A(mai_mai_n973_), .B(mai_mai_n117_), .Y(mai_mai_n1878_));
  OAI220     m1829(.A0(mai_mai_n630_), .A1(mai_mai_n162_), .B0(mai_mai_n328_), .B1(mai_mai_n134_), .Y(mai_mai_n1879_));
  OAI210     m1830(.A0(mai_mai_n1879_), .A1(mai_mai_n1878_), .B0(mai_mai_n68_), .Y(mai_mai_n1880_));
  NO2        m1831(.A(mai_mai_n1664_), .B(mai_mai_n340_), .Y(mai_mai_n1881_));
  OAI210     m1832(.A0(mai_mai_n1589_), .A1(mai_mai_n559_), .B0(mai_mai_n1881_), .Y(mai_mai_n1882_));
  NA4        m1833(.A(mai_mai_n1882_), .B(mai_mai_n1880_), .C(mai_mai_n1877_), .D(mai_mai_n1873_), .Y(mai_mai_n1883_));
  OAI210     m1834(.A0(mai_mai_n1883_), .A1(mai_mai_n1872_), .B0(mai_mai_n1869_), .Y(mai_mai_n1884_));
  INV        m1835(.A(mai_mai_n344_), .Y(mai_mai_n1885_));
  NA2        m1836(.A(mai_mai_n1218_), .B(mai_mai_n1885_), .Y(mai_mai_n1886_));
  NO3        m1837(.A(x8), .B(mai_mai_n71_), .C(x2), .Y(mai_mai_n1887_));
  NA2        m1838(.A(mai_mai_n906_), .B(mai_mai_n1008_), .Y(mai_mai_n1888_));
  AOI210     m1839(.A0(mai_mai_n617_), .A1(mai_mai_n630_), .B0(mai_mai_n1888_), .Y(mai_mai_n1889_));
  AOI210     m1840(.A0(mai_mai_n541_), .A1(mai_mai_n572_), .B0(mai_mai_n636_), .Y(mai_mai_n1890_));
  NO2        m1841(.A(mai_mai_n1890_), .B(mai_mai_n1556_), .Y(mai_mai_n1891_));
  NO2        m1842(.A(mai_mai_n417_), .B(mai_mai_n400_), .Y(mai_mai_n1892_));
  NOi31      m1843(.An(mai_mai_n1291_), .B(mai_mai_n1892_), .C(mai_mai_n541_), .Y(mai_mai_n1893_));
  NO3        m1844(.A(mai_mai_n1893_), .B(mai_mai_n1891_), .C(mai_mai_n1889_), .Y(mai_mai_n1894_));
  NA4        m1845(.A(mai_mai_n1894_), .B(mai_mai_n1886_), .C(mai_mai_n1884_), .D(mai_mai_n1853_), .Y(mai33));
  OAI210     m1846(.A0(mai_mai_n747_), .A1(x1), .B0(mai_mai_n185_), .Y(mai_mai_n1896_));
  OAI210     m1847(.A0(mai_mai_n1749_), .A1(mai_mai_n167_), .B0(mai_mai_n302_), .Y(mai_mai_n1897_));
  OAI210     m1848(.A0(mai_mai_n1439_), .A1(mai_mai_n327_), .B0(mai_mai_n746_), .Y(mai_mai_n1898_));
  NA3        m1849(.A(mai_mai_n1898_), .B(mai_mai_n1897_), .C(mai_mai_n581_), .Y(mai_mai_n1899_));
  AOI210     m1850(.A0(mai_mai_n1896_), .A1(x5), .B0(mai_mai_n1899_), .Y(mai_mai_n1900_));
  NA2        m1851(.A(mai_mai_n209_), .B(mai_mai_n76_), .Y(mai_mai_n1901_));
  NA4        m1852(.A(mai_mai_n1501_), .B(mai_mai_n520_), .C(mai_mai_n226_), .D(x4), .Y(mai_mai_n1902_));
  AOI210     m1853(.A0(mai_mai_n1902_), .A1(mai_mai_n1901_), .B0(mai_mai_n327_), .Y(mai_mai_n1903_));
  OAI210     m1854(.A0(mai_mai_n402_), .A1(mai_mai_n246_), .B0(mai_mai_n53_), .Y(mai_mai_n1904_));
  AOI210     m1855(.A0(mai_mai_n1904_), .A1(mai_mai_n404_), .B0(mai_mai_n64_), .Y(mai_mai_n1905_));
  NA2        m1856(.A(mai_mai_n1430_), .B(mai_mai_n71_), .Y(mai_mai_n1906_));
  NO3        m1857(.A(mai_mai_n1906_), .B(mai_mai_n1905_), .C(mai_mai_n1903_), .Y(mai_mai_n1907_));
  OAI210     m1858(.A0(mai_mai_n1900_), .A1(x4), .B0(mai_mai_n1907_), .Y(mai_mai_n1908_));
  NO2        m1859(.A(mai_mai_n1849_), .B(mai_mai_n197_), .Y(mai_mai_n1909_));
  OAI210     m1860(.A0(mai_mai_n788_), .A1(mai_mai_n51_), .B0(x6), .Y(mai_mai_n1910_));
  NA3        m1861(.A(mai_mai_n837_), .B(mai_mai_n674_), .C(mai_mai_n55_), .Y(mai_mai_n1911_));
  OAI210     m1862(.A0(mai_mai_n568_), .A1(mai_mai_n465_), .B0(mai_mai_n1911_), .Y(mai_mai_n1912_));
  NO3        m1863(.A(mai_mai_n1912_), .B(mai_mai_n1910_), .C(mai_mai_n1909_), .Y(mai_mai_n1913_));
  INV        m1864(.A(mai_mai_n1913_), .Y(mai_mai_n1914_));
  NA3        m1865(.A(mai_mai_n1914_), .B(mai_mai_n1908_), .C(mai_mai_n59_), .Y(mai_mai_n1915_));
  NA2        m1866(.A(mai_mai_n494_), .B(mai_mai_n104_), .Y(mai_mai_n1916_));
  NO3        m1867(.A(mai_mai_n1348_), .B(mai_mai_n348_), .C(x4), .Y(mai_mai_n1917_));
  AOI210     m1868(.A0(mai_mai_n1917_), .A1(mai_mai_n1916_), .B0(mai_mai_n405_), .Y(mai_mai_n1918_));
  NA2        m1869(.A(mai_mai_n749_), .B(mai_mai_n103_), .Y(mai_mai_n1919_));
  NA2        m1870(.A(mai_mai_n1919_), .B(mai_mai_n428_), .Y(mai_mai_n1920_));
  NO2        m1871(.A(mai_mai_n651_), .B(mai_mai_n349_), .Y(mai_mai_n1921_));
  NA2        m1872(.A(mai_mai_n461_), .B(mai_mai_n53_), .Y(mai_mai_n1922_));
  AOI210     m1873(.A0(mai_mai_n1921_), .A1(mai_mai_n1920_), .B0(mai_mai_n1922_), .Y(mai_mai_n1923_));
  OAI210     m1874(.A0(mai_mai_n1918_), .A1(mai_mai_n59_), .B0(mai_mai_n1923_), .Y(mai_mai_n1924_));
  AOI220     m1875(.A0(mai_mai_n630_), .A1(mai_mai_n216_), .B0(mai_mai_n361_), .B1(mai_mai_n210_), .Y(mai_mai_n1925_));
  NA2        m1876(.A(mai_mai_n675_), .B(mai_mai_n874_), .Y(mai_mai_n1926_));
  OAI210     m1877(.A0(mai_mai_n1926_), .A1(mai_mai_n1925_), .B0(mai_mai_n276_), .Y(mai_mai_n1927_));
  AOI210     m1878(.A0(mai_mai_n1778_), .A1(mai_mai_n198_), .B0(mai_mai_n53_), .Y(mai_mai_n1928_));
  NO2        m1879(.A(mai_mai_n134_), .B(mai_mai_n312_), .Y(mai_mai_n1929_));
  AOI220     m1880(.A0(mai_mai_n1929_), .A1(mai_mai_n887_), .B0(mai_mai_n616_), .B1(mai_mai_n327_), .Y(mai_mai_n1930_));
  NA2        m1881(.A(mai_mai_n413_), .B(mai_mai_n459_), .Y(mai_mai_n1931_));
  NO3        m1882(.A(mai_mai_n1931_), .B(mai_mai_n920_), .C(mai_mai_n172_), .Y(mai_mai_n1932_));
  AOI210     m1883(.A0(mai_mai_n1535_), .A1(mai_mai_n1045_), .B0(mai_mai_n1932_), .Y(mai_mai_n1933_));
  NA4        m1884(.A(mai_mai_n1933_), .B(mai_mai_n1930_), .C(mai_mai_n1928_), .D(mai_mai_n1927_), .Y(mai_mai_n1934_));
  NA3        m1885(.A(mai_mai_n1934_), .B(mai_mai_n1924_), .C(mai_mai_n57_), .Y(mai_mai_n1935_));
  AN2        m1886(.A(mai_mai_n415_), .B(mai_mai_n131_), .Y(mai_mai_n1936_));
  NA3        m1887(.A(mai_mai_n713_), .B(mai_mai_n327_), .C(mai_mai_n60_), .Y(mai_mai_n1937_));
  OAI210     m1888(.A0(mai_mai_n1317_), .A1(mai_mai_n323_), .B0(mai_mai_n106_), .Y(mai_mai_n1938_));
  INV        m1889(.A(mai_mai_n131_), .Y(mai_mai_n1939_));
  OAI210     m1890(.A0(mai_mai_n1939_), .A1(mai_mai_n361_), .B0(mai_mai_n1938_), .Y(mai_mai_n1940_));
  NA2        m1891(.A(mai_mai_n1940_), .B(mai_mai_n100_), .Y(mai_mai_n1941_));
  INV        m1892(.A(mai_mai_n356_), .Y(mai_mai_n1942_));
  NA2        m1893(.A(mai_mai_n1942_), .B(mai_mai_n1560_), .Y(mai_mai_n1943_));
  AOI220     m1894(.A0(mai_mai_n1855_), .A1(mai_mai_n269_), .B0(mai_mai_n1173_), .B1(mai_mai_n1030_), .Y(mai_mai_n1944_));
  NA3        m1895(.A(mai_mai_n1944_), .B(mai_mai_n1943_), .C(mai_mai_n1941_), .Y(mai_mai_n1945_));
  AOI210     m1896(.A0(mai_mai_n1936_), .A1(x7), .B0(mai_mai_n1945_), .Y(mai_mai_n1946_));
  NA3        m1897(.A(mai_mai_n1946_), .B(mai_mai_n1935_), .C(mai_mai_n1915_), .Y(mai34));
  NA2        m1898(.A(mai_mai_n677_), .B(x8), .Y(mai_mai_n1948_));
  AO210      m1899(.A0(mai_mai_n1948_), .A1(mai_mai_n447_), .B0(mai_mai_n606_), .Y(mai_mai_n1949_));
  NA2        m1900(.A(mai_mai_n616_), .B(mai_mai_n575_), .Y(mai_mai_n1950_));
  AOI210     m1901(.A0(mai_mai_n1950_), .A1(mai_mai_n1949_), .B0(mai_mai_n242_), .Y(mai_mai_n1951_));
  NO2        m1902(.A(mai_mai_n1379_), .B(mai_mai_n58_), .Y(mai_mai_n1952_));
  NA3        m1903(.A(mai_mai_n1952_), .B(mai_mai_n313_), .C(x8), .Y(mai_mai_n1953_));
  NO3        m1904(.A(mai_mai_n886_), .B(mai_mai_n651_), .C(mai_mai_n422_), .Y(mai_mai_n1954_));
  INV        m1905(.A(mai_mai_n1954_), .Y(mai_mai_n1955_));
  NA2        m1906(.A(mai_mai_n127_), .B(x0), .Y(mai_mai_n1956_));
  NAi31      m1907(.An(mai_mai_n1956_), .B(mai_mai_n2224_), .C(mai_mai_n735_), .Y(mai_mai_n1957_));
  NA3        m1908(.A(mai_mai_n1375_), .B(mai_mai_n1207_), .C(mai_mai_n50_), .Y(mai_mai_n1958_));
  NA4        m1909(.A(mai_mai_n1958_), .B(mai_mai_n1957_), .C(mai_mai_n1955_), .D(mai_mai_n1953_), .Y(mai_mai_n1959_));
  NA2        m1910(.A(mai_mai_n983_), .B(mai_mai_n690_), .Y(mai_mai_n1960_));
  NA3        m1911(.A(mai_mai_n1010_), .B(mai_mai_n156_), .C(mai_mai_n974_), .Y(mai_mai_n1961_));
  AOI210     m1912(.A0(mai_mai_n1961_), .A1(mai_mai_n1960_), .B0(mai_mai_n699_), .Y(mai_mai_n1962_));
  AOI210     m1913(.A0(mai_mai_n1526_), .A1(mai_mai_n124_), .B0(mai_mai_n1962_), .Y(mai_mai_n1963_));
  NO2        m1914(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n1964_));
  NA3        m1915(.A(mai_mai_n1964_), .B(mai_mai_n677_), .C(mai_mai_n56_), .Y(mai_mai_n1965_));
  OAI210     m1916(.A0(mai_mai_n1963_), .A1(mai_mai_n134_), .B0(mai_mai_n1965_), .Y(mai_mai_n1966_));
  NO3        m1917(.A(mai_mai_n1966_), .B(mai_mai_n1959_), .C(mai_mai_n1951_), .Y(mai_mai_n1967_));
  INV        m1918(.A(mai_mai_n862_), .Y(mai_mai_n1968_));
  NO3        m1919(.A(mai_mai_n1968_), .B(mai_mai_n411_), .C(mai_mai_n301_), .Y(mai_mai_n1969_));
  INV        m1920(.A(mai_mai_n722_), .Y(mai_mai_n1970_));
  INV        m1921(.A(mai_mai_n276_), .Y(mai_mai_n1971_));
  OAI220     m1922(.A0(mai_mai_n1971_), .A1(mai_mai_n1340_), .B0(mai_mai_n1970_), .B1(mai_mai_n1034_), .Y(mai_mai_n1972_));
  OAI210     m1923(.A0(mai_mai_n1972_), .A1(mai_mai_n1969_), .B0(x2), .Y(mai_mai_n1973_));
  INV        m1924(.A(mai_mai_n1973_), .Y(mai_mai_n1974_));
  OAI220     m1925(.A0(mai_mai_n687_), .A1(mai_mai_n55_), .B0(mai_mai_n255_), .B1(mai_mai_n102_), .Y(mai_mai_n1975_));
  NO4        m1926(.A(mai_mai_n414_), .B(mai_mai_n77_), .C(x7), .D(x3), .Y(mai_mai_n1976_));
  NO2        m1927(.A(mai_mai_n983_), .B(mai_mai_n263_), .Y(mai_mai_n1977_));
  NO4        m1928(.A(mai_mai_n1977_), .B(mai_mai_n1976_), .C(mai_mai_n1975_), .D(mai_mai_n2221_), .Y(mai_mai_n1978_));
  NA2        m1929(.A(mai_mai_n1083_), .B(mai_mai_n939_), .Y(mai_mai_n1979_));
  NA4        m1930(.A(mai_mai_n677_), .B(mai_mai_n168_), .C(mai_mai_n57_), .D(mai_mai_n103_), .Y(mai_mai_n1980_));
  NA3        m1931(.A(mai_mai_n1206_), .B(mai_mai_n234_), .C(x7), .Y(mai_mai_n1981_));
  NA3        m1932(.A(mai_mai_n1981_), .B(mai_mai_n1980_), .C(mai_mai_n1979_), .Y(mai_mai_n1982_));
  OAI210     m1933(.A0(mai_mai_n1982_), .A1(mai_mai_n1978_), .B0(mai_mai_n153_), .Y(mai_mai_n1983_));
  NA3        m1934(.A(mai_mai_n1014_), .B(mai_mai_n271_), .C(mai_mai_n539_), .Y(mai_mai_n1984_));
  NA2        m1935(.A(mai_mai_n1018_), .B(mai_mai_n620_), .Y(mai_mai_n1985_));
  OAI210     m1936(.A0(mai_mai_n1985_), .A1(mai_mai_n243_), .B0(mai_mai_n1815_), .Y(mai_mai_n1986_));
  AOI220     m1937(.A0(mai_mai_n1986_), .A1(x7), .B0(mai_mai_n905_), .B1(mai_mai_n607_), .Y(mai_mai_n1987_));
  OAI210     m1938(.A0(mai_mai_n1722_), .A1(mai_mai_n239_), .B0(mai_mai_n680_), .Y(mai_mai_n1988_));
  AOI220     m1939(.A0(mai_mai_n382_), .A1(x8), .B0(mai_mai_n92_), .B1(x2), .Y(mai_mai_n1989_));
  AOI210     m1940(.A0(mai_mai_n247_), .A1(mai_mai_n53_), .B0(mai_mai_n598_), .Y(mai_mai_n1990_));
  OAI220     m1941(.A0(mai_mai_n1990_), .A1(mai_mai_n97_), .B0(mai_mai_n1989_), .B1(mai_mai_n1164_), .Y(mai_mai_n1991_));
  AOI220     m1942(.A0(mai_mai_n1991_), .A1(mai_mai_n1145_), .B0(mai_mai_n1988_), .B1(mai_mai_n1304_), .Y(mai_mai_n1992_));
  NA4        m1943(.A(mai_mai_n1992_), .B(mai_mai_n1987_), .C(mai_mai_n1984_), .D(mai_mai_n1983_), .Y(mai_mai_n1993_));
  AOI210     m1944(.A0(mai_mai_n1974_), .A1(mai_mai_n751_), .B0(mai_mai_n1993_), .Y(mai_mai_n1994_));
  OAI210     m1945(.A0(mai_mai_n1967_), .A1(x2), .B0(mai_mai_n1994_), .Y(mai35));
  NA2        m1946(.A(mai_mai_n465_), .B(mai_mai_n168_), .Y(mai_mai_n1996_));
  AOI220     m1947(.A0(mai_mai_n582_), .A1(mai_mai_n55_), .B0(mai_mai_n713_), .B1(mai_mai_n1071_), .Y(mai_mai_n1997_));
  AOI210     m1948(.A0(mai_mai_n1997_), .A1(mai_mai_n1996_), .B0(mai_mai_n71_), .Y(mai_mai_n1998_));
  NO2        m1949(.A(mai_mai_n473_), .B(mai_mai_n312_), .Y(mai_mai_n1999_));
  OAI210     m1950(.A0(mai_mai_n1999_), .A1(mai_mai_n1998_), .B0(x2), .Y(mai_mai_n2000_));
  AOI210     m1951(.A0(mai_mai_n199_), .A1(x0), .B0(mai_mai_n249_), .Y(mai_mai_n2001_));
  OAI220     m1952(.A0(mai_mai_n2001_), .A1(mai_mai_n612_), .B0(mai_mai_n184_), .B1(x4), .Y(mai_mai_n2002_));
  NA2        m1953(.A(mai_mai_n2002_), .B(mai_mai_n131_), .Y(mai_mai_n2003_));
  NA3        m1954(.A(mai_mai_n382_), .B(x8), .C(mai_mai_n71_), .Y(mai_mai_n2004_));
  AOI210     m1955(.A0(mai_mai_n2004_), .A1(mai_mai_n1479_), .B0(mai_mai_n630_), .Y(mai_mai_n2005_));
  OAI210     m1956(.A0(mai_mai_n1937_), .A1(x6), .B0(mai_mai_n689_), .Y(mai_mai_n2006_));
  NO2        m1957(.A(mai_mai_n2006_), .B(mai_mai_n2005_), .Y(mai_mai_n2007_));
  NA3        m1958(.A(mai_mai_n2007_), .B(mai_mai_n2003_), .C(mai_mai_n2000_), .Y(mai_mai_n2008_));
  NO3        m1959(.A(mai_mai_n625_), .B(mai_mai_n55_), .C(x6), .Y(mai_mai_n2009_));
  OAI210     m1960(.A0(mai_mai_n2009_), .A1(mai_mai_n654_), .B0(mai_mai_n202_), .Y(mai_mai_n2010_));
  NA2        m1961(.A(mai_mai_n1152_), .B(mai_mai_n63_), .Y(mai_mai_n2011_));
  OAI210     m1962(.A0(mai_mai_n962_), .A1(x6), .B0(mai_mai_n438_), .Y(mai_mai_n2012_));
  NA3        m1963(.A(mai_mai_n2012_), .B(mai_mai_n2011_), .C(mai_mai_n2010_), .Y(mai_mai_n2013_));
  NA3        m1964(.A(mai_mai_n1108_), .B(mai_mai_n692_), .C(x3), .Y(mai_mai_n2014_));
  NO3        m1965(.A(mai_mai_n2014_), .B(mai_mai_n627_), .C(mai_mai_n190_), .Y(mai_mai_n2015_));
  AOI210     m1966(.A0(mai_mai_n2013_), .A1(mai_mai_n50_), .B0(mai_mai_n2015_), .Y(mai_mai_n2016_));
  INV        m1967(.A(mai_mai_n2016_), .Y(mai_mai_n2017_));
  AOI210     m1968(.A0(mai_mai_n2008_), .A1(mai_mai_n57_), .B0(mai_mai_n2017_), .Y(mai_mai_n2018_));
  NA2        m1969(.A(mai_mai_n870_), .B(mai_mai_n63_), .Y(mai_mai_n2019_));
  NO2        m1970(.A(mai_mai_n2019_), .B(mai_mai_n50_), .Y(mai_mai_n2020_));
  OAI210     m1971(.A0(mai_mai_n870_), .A1(mai_mai_n232_), .B0(mai_mai_n693_), .Y(mai_mai_n2021_));
  OAI210     m1972(.A0(mai_mai_n232_), .A1(mai_mai_n538_), .B0(mai_mai_n1812_), .Y(mai_mai_n2022_));
  NA2        m1973(.A(mai_mai_n2022_), .B(mai_mai_n2021_), .Y(mai_mai_n2023_));
  OAI210     m1974(.A0(mai_mai_n2023_), .A1(mai_mai_n2020_), .B0(mai_mai_n59_), .Y(mai_mai_n2024_));
  NO4        m1975(.A(mai_mai_n863_), .B(mai_mai_n519_), .C(mai_mai_n336_), .D(mai_mai_n380_), .Y(mai_mai_n2025_));
  XN2        m1976(.A(x4), .B(x3), .Y(mai_mai_n2026_));
  NO3        m1977(.A(mai_mai_n2026_), .B(mai_mai_n611_), .C(mai_mai_n282_), .Y(mai_mai_n2027_));
  NO2        m1978(.A(mai_mai_n2027_), .B(mai_mai_n2025_), .Y(mai_mai_n2028_));
  INV        m1979(.A(mai_mai_n2028_), .Y(mai_mai_n2029_));
  NO3        m1980(.A(mai_mai_n687_), .B(mai_mai_n788_), .C(mai_mai_n250_), .Y(mai_mai_n2030_));
  OAI210     m1981(.A0(mai_mai_n2030_), .A1(mai_mai_n1261_), .B0(mai_mai_n50_), .Y(mai_mai_n2031_));
  INV        m1982(.A(mai_mai_n2031_), .Y(mai_mai_n2032_));
  AOI210     m1983(.A0(mai_mai_n2029_), .A1(mai_mai_n541_), .B0(mai_mai_n2032_), .Y(mai_mai_n2033_));
  NO2        m1984(.A(mai_mai_n589_), .B(mai_mai_n627_), .Y(mai_mai_n2034_));
  NA2        m1985(.A(mai_mai_n558_), .B(mai_mai_n1887_), .Y(mai_mai_n2035_));
  OAI210     m1986(.A0(mai_mai_n1948_), .A1(mai_mai_n57_), .B0(mai_mai_n2035_), .Y(mai_mai_n2036_));
  OAI210     m1987(.A0(mai_mai_n2036_), .A1(mai_mai_n2034_), .B0(mai_mai_n92_), .Y(mai_mai_n2037_));
  NO2        m1988(.A(mai_mai_n263_), .B(x6), .Y(mai_mai_n2038_));
  NA2        m1989(.A(mai_mai_n1530_), .B(mai_mai_n2038_), .Y(mai_mai_n2039_));
  NA4        m1990(.A(mai_mai_n2039_), .B(mai_mai_n2037_), .C(mai_mai_n2033_), .D(mai_mai_n2024_), .Y(mai_mai_n2040_));
  NA3        m1991(.A(mai_mai_n1236_), .B(mai_mai_n1109_), .C(mai_mai_n755_), .Y(mai_mai_n2041_));
  AOI220     m1992(.A0(mai_mai_n1636_), .A1(mai_mai_n131_), .B0(mai_mai_n391_), .B1(mai_mai_n121_), .Y(mai_mai_n2042_));
  AOI210     m1993(.A0(mai_mai_n2042_), .A1(mai_mai_n2041_), .B0(mai_mai_n1299_), .Y(mai_mai_n2043_));
  NO2        m1994(.A(mai_mai_n582_), .B(x3), .Y(mai_mai_n2044_));
  NO3        m1995(.A(mai_mai_n638_), .B(mai_mai_n1379_), .C(x2), .Y(mai_mai_n2045_));
  AOI220     m1996(.A0(mai_mai_n2045_), .A1(mai_mai_n2044_), .B0(mai_mai_n1624_), .B1(mai_mai_n709_), .Y(mai_mai_n2046_));
  NA3        m1997(.A(x6), .B(x4), .C(x0), .Y(mai_mai_n2047_));
  OAI220     m1998(.A0(mai_mai_n2047_), .A1(mai_mai_n183_), .B0(mai_mai_n625_), .B1(mai_mai_n489_), .Y(mai_mai_n2048_));
  NO2        m1999(.A(mai_mai_n348_), .B(mai_mai_n326_), .Y(mai_mai_n2049_));
  AOI220     m2000(.A0(mai_mai_n2049_), .A1(mai_mai_n391_), .B0(mai_mai_n2048_), .B1(mai_mai_n836_), .Y(mai_mai_n2050_));
  OAI210     m2001(.A0(mai_mai_n2046_), .A1(mai_mai_n1025_), .B0(mai_mai_n2050_), .Y(mai_mai_n2051_));
  NO2        m2002(.A(mai_mai_n2051_), .B(mai_mai_n2043_), .Y(mai_mai_n2052_));
  INV        m2003(.A(mai_mai_n2052_), .Y(mai_mai_n2053_));
  AOI210     m2004(.A0(mai_mai_n2040_), .A1(x5), .B0(mai_mai_n2053_), .Y(mai_mai_n2054_));
  OAI210     m2005(.A0(mai_mai_n2018_), .A1(x5), .B0(mai_mai_n2054_), .Y(mai36));
  NA2        m2006(.A(mai_mai_n1855_), .B(mai_mai_n255_), .Y(mai_mai_n2056_));
  NA3        m2007(.A(mai_mai_n413_), .B(mai_mai_n207_), .C(mai_mai_n116_), .Y(mai_mai_n2057_));
  NA2        m2008(.A(mai_mai_n2057_), .B(mai_mai_n2056_), .Y(mai_mai_n2058_));
  NO3        m2009(.A(mai_mai_n105_), .B(mai_mai_n883_), .C(mai_mai_n498_), .Y(mai_mai_n2059_));
  OAI210     m2010(.A0(mai_mai_n394_), .A1(mai_mai_n2059_), .B0(mai_mai_n433_), .Y(mai_mai_n2060_));
  NO2        m2011(.A(mai_mai_n595_), .B(mai_mai_n243_), .Y(mai_mai_n2061_));
  NO3        m2012(.A(mai_mai_n1595_), .B(mai_mai_n1378_), .C(mai_mai_n251_), .Y(mai_mai_n2062_));
  NO2        m2013(.A(mai_mai_n2019_), .B(mai_mai_n209_), .Y(mai_mai_n2063_));
  NO3        m2014(.A(mai_mai_n2063_), .B(mai_mai_n2062_), .C(mai_mai_n2061_), .Y(mai_mai_n2064_));
  INV        m2015(.A(mai_mai_n877_), .Y(mai_mai_n2065_));
  OAI220     m2016(.A0(mai_mai_n1422_), .A1(mai_mai_n1417_), .B0(mai_mai_n877_), .B1(mai_mai_n974_), .Y(mai_mai_n2066_));
  AOI220     m2017(.A0(mai_mai_n2066_), .A1(mai_mai_n115_), .B0(mai_mai_n2065_), .B1(mai_mai_n575_), .Y(mai_mai_n2067_));
  NA3        m2018(.A(mai_mai_n2067_), .B(mai_mai_n2064_), .C(mai_mai_n2060_), .Y(mai_mai_n2068_));
  AOI210     m2019(.A0(mai_mai_n2058_), .A1(mai_mai_n313_), .B0(mai_mai_n2068_), .Y(mai_mai_n2069_));
  OAI210     m2020(.A0(mai_mai_n546_), .A1(mai_mai_n478_), .B0(mai_mai_n157_), .Y(mai_mai_n2070_));
  OAI210     m2021(.A0(mai_mai_n1677_), .A1(mai_mai_n70_), .B0(mai_mai_n2070_), .Y(mai_mai_n2071_));
  OAI210     m2022(.A0(mai_mai_n457_), .A1(mai_mai_n218_), .B0(mai_mai_n232_), .Y(mai_mai_n2072_));
  NO2        m2023(.A(mai_mai_n1684_), .B(mai_mai_n164_), .Y(mai_mai_n2073_));
  NA2        m2024(.A(mai_mai_n1064_), .B(mai_mai_n55_), .Y(mai_mai_n2074_));
  OAI210     m2025(.A0(mai_mai_n2074_), .A1(mai_mai_n2073_), .B0(mai_mai_n2072_), .Y(mai_mai_n2075_));
  OAI210     m2026(.A0(mai_mai_n2075_), .A1(mai_mai_n2071_), .B0(mai_mai_n814_), .Y(mai_mai_n2076_));
  AOI210     m2027(.A0(mai_mai_n102_), .A1(mai_mai_n105_), .B0(mai_mai_n315_), .Y(mai_mai_n2077_));
  NA2        m2028(.A(mai_mai_n616_), .B(mai_mai_n1379_), .Y(mai_mai_n2078_));
  OAI220     m2029(.A0(mai_mai_n2078_), .A1(mai_mai_n2077_), .B0(mai_mai_n689_), .B1(mai_mai_n1094_), .Y(mai_mai_n2079_));
  NO2        m2030(.A(mai_mai_n1207_), .B(mai_mai_n532_), .Y(mai_mai_n2080_));
  NO3        m2031(.A(mai_mai_n2080_), .B(mai_mai_n1534_), .C(mai_mai_n638_), .Y(mai_mai_n2081_));
  NOi31      m2032(.An(mai_mai_n1693_), .B(mai_mai_n1931_), .C(mai_mai_n698_), .Y(mai_mai_n2082_));
  NO3        m2033(.A(mai_mai_n2082_), .B(mai_mai_n2081_), .C(mai_mai_n2079_), .Y(mai_mai_n2083_));
  AOI210     m2034(.A0(mai_mai_n2083_), .A1(mai_mai_n2076_), .B0(x7), .Y(mai_mai_n2084_));
  NA2        m2035(.A(mai_mai_n130_), .B(mai_mai_n63_), .Y(mai_mai_n2085_));
  AOI210     m2036(.A0(mai_mai_n541_), .A1(mai_mai_n572_), .B0(mai_mai_n1045_), .Y(mai_mai_n2086_));
  NA4        m2037(.A(mai_mai_n2086_), .B(mai_mai_n2085_), .C(mai_mai_n886_), .D(mai_mai_n811_), .Y(mai_mai_n2087_));
  NA2        m2038(.A(mai_mai_n2087_), .B(mai_mai_n465_), .Y(mai_mai_n2088_));
  AOI220     m2039(.A0(mai_mai_n1501_), .A1(mai_mai_n235_), .B0(mai_mai_n939_), .B1(mai_mai_n121_), .Y(mai_mai_n2089_));
  NO2        m2040(.A(mai_mai_n2089_), .B(mai_mai_n413_), .Y(mai_mai_n2090_));
  NO2        m2041(.A(mai_mai_n380_), .B(mai_mai_n207_), .Y(mai_mai_n2091_));
  NO3        m2042(.A(mai_mai_n2091_), .B(mai_mai_n1111_), .C(mai_mai_n59_), .Y(mai_mai_n2092_));
  AOI210     m2043(.A0(mai_mai_n1072_), .A1(mai_mai_n381_), .B0(x6), .Y(mai_mai_n2093_));
  NA3        m2044(.A(mai_mai_n1443_), .B(mai_mai_n255_), .C(mai_mai_n247_), .Y(mai_mai_n2094_));
  NA2        m2045(.A(mai_mai_n2094_), .B(mai_mai_n1404_), .Y(mai_mai_n2095_));
  NO4        m2046(.A(mai_mai_n2095_), .B(mai_mai_n2093_), .C(mai_mai_n2092_), .D(mai_mai_n2090_), .Y(mai_mai_n2096_));
  AOI210     m2047(.A0(mai_mai_n2096_), .A1(mai_mai_n2088_), .B0(mai_mai_n422_), .Y(mai_mai_n2097_));
  NO3        m2048(.A(mai_mai_n2026_), .B(mai_mai_n820_), .C(mai_mai_n464_), .Y(mai_mai_n2098_));
  AOI210     m2049(.A0(mai_mai_n1110_), .A1(mai_mai_n246_), .B0(mai_mai_n2098_), .Y(mai_mai_n2099_));
  NO2        m2050(.A(mai_mai_n564_), .B(mai_mai_n105_), .Y(mai_mai_n2100_));
  AN2        m2051(.A(mai_mai_n2100_), .B(x5), .Y(mai_mai_n2101_));
  NO2        m2052(.A(mai_mai_n429_), .B(mai_mai_n392_), .Y(mai_mai_n2102_));
  NA2        m2053(.A(mai_mai_n2102_), .B(mai_mai_n2101_), .Y(mai_mai_n2103_));
  OAI210     m2054(.A0(mai_mai_n2099_), .A1(x1), .B0(mai_mai_n2103_), .Y(mai_mai_n2104_));
  NO3        m2055(.A(mai_mai_n2104_), .B(mai_mai_n2097_), .C(mai_mai_n2084_), .Y(mai_mai_n2105_));
  OAI210     m2056(.A0(mai_mai_n2069_), .A1(mai_mai_n57_), .B0(mai_mai_n2105_), .Y(mai37));
  NA3        m2057(.A(mai_mai_n960_), .B(mai_mai_n133_), .C(x3), .Y(mai_mai_n2107_));
  NO2        m2058(.A(mai_mai_n2107_), .B(mai_mai_n631_), .Y(mai_mai_n2108_));
  NO2        m2059(.A(mai_mai_n960_), .B(mai_mai_n351_), .Y(mai_mai_n2109_));
  OAI210     m2060(.A0(mai_mai_n2109_), .A1(mai_mai_n2108_), .B0(mai_mai_n56_), .Y(mai_mai_n2110_));
  NA2        m2061(.A(mai_mai_n553_), .B(mai_mai_n690_), .Y(mai_mai_n2111_));
  AOI210     m2062(.A0(mai_mai_n2111_), .A1(mai_mai_n940_), .B0(x3), .Y(mai_mai_n2112_));
  AOI220     m2063(.A0(mai_mai_n553_), .A1(mai_mai_n690_), .B0(mai_mai_n433_), .B1(mai_mai_n939_), .Y(mai_mai_n2113_));
  NO2        m2064(.A(mai_mai_n611_), .B(mai_mai_n171_), .Y(mai_mai_n2114_));
  OAI220     m2065(.A0(mai_mai_n2114_), .A1(mai_mai_n766_), .B0(mai_mai_n2113_), .B1(mai_mai_n105_), .Y(mai_mai_n2115_));
  OAI210     m2066(.A0(mai_mai_n2115_), .A1(mai_mai_n2112_), .B0(mai_mai_n71_), .Y(mai_mai_n2116_));
  NA2        m2067(.A(mai_mai_n1047_), .B(mai_mai_n962_), .Y(mai_mai_n2117_));
  OAI210     m2068(.A0(mai_mai_n1066_), .A1(mai_mai_n177_), .B0(mai_mai_n423_), .Y(mai_mai_n2118_));
  NA4        m2069(.A(mai_mai_n2118_), .B(mai_mai_n2117_), .C(mai_mai_n2116_), .D(mai_mai_n2110_), .Y(mai_mai_n2119_));
  NA2        m2070(.A(mai_mai_n2119_), .B(mai_mai_n68_), .Y(mai_mai_n2120_));
  NA2        m2071(.A(mai_mai_n321_), .B(mai_mai_n249_), .Y(mai_mai_n2121_));
  NA2        m2072(.A(mai_mai_n376_), .B(mai_mai_n105_), .Y(mai_mai_n2122_));
  NO2        m2073(.A(mai_mai_n490_), .B(mai_mai_n56_), .Y(mai_mai_n2123_));
  NA3        m2074(.A(mai_mai_n2123_), .B(mai_mai_n2122_), .C(mai_mai_n2121_), .Y(mai_mai_n2124_));
  INV        m2075(.A(mai_mai_n2124_), .Y(mai_mai_n2125_));
  NO2        m2076(.A(mai_mai_n56_), .B(mai_mai_n2125_), .Y(mai_mai_n2126_));
  NA2        m2077(.A(mai_mai_n2126_), .B(mai_mai_n100_), .Y(mai_mai_n2127_));
  NA2        m2078(.A(mai_mai_n638_), .B(mai_mai_n1052_), .Y(mai_mai_n2128_));
  NOi21      m2079(.An(mai_mai_n1178_), .B(mai_mai_n106_), .Y(mai_mai_n2129_));
  NA2        m2080(.A(mai_mai_n2129_), .B(mai_mai_n2128_), .Y(mai_mai_n2130_));
  NO2        m2081(.A(mai_mai_n1864_), .B(mai_mai_n55_), .Y(mai_mai_n2131_));
  OAI210     m2082(.A0(mai_mai_n2131_), .A1(mai_mai_n2130_), .B0(mai_mai_n1560_), .Y(mai_mai_n2132_));
  NA2        m2083(.A(mai_mai_n168_), .B(mai_mai_n103_), .Y(mai_mai_n2133_));
  NA2        m2084(.A(mai_mai_n630_), .B(x6), .Y(mai_mai_n2134_));
  AOI210     m2085(.A0(mai_mai_n2134_), .A1(mai_mai_n447_), .B0(mai_mai_n2133_), .Y(mai_mai_n2135_));
  AOI210     m2086(.A0(mai_mai_n328_), .A1(mai_mai_n133_), .B0(mai_mai_n134_), .Y(mai_mai_n2136_));
  OAI210     m2087(.A0(mai_mai_n2136_), .A1(mai_mai_n2135_), .B0(mai_mai_n321_), .Y(mai_mai_n2137_));
  AOI210     m2088(.A0(mai_mai_n565_), .A1(mai_mai_n402_), .B0(mai_mai_n1119_), .Y(mai_mai_n2138_));
  NO3        m2089(.A(mai_mai_n2138_), .B(mai_mai_n243_), .C(mai_mai_n63_), .Y(mai_mai_n2139_));
  OAI220     m2090(.A0(mai_mai_n1948_), .A1(mai_mai_n446_), .B0(mai_mai_n1761_), .B1(mai_mai_n361_), .Y(mai_mai_n2140_));
  OAI210     m2091(.A0(mai_mai_n2140_), .A1(mai_mai_n2139_), .B0(mai_mai_n53_), .Y(mai_mai_n2141_));
  NO4        m2092(.A(mai_mai_n1956_), .B(mai_mai_n845_), .C(mai_mai_n403_), .D(mai_mai_n204_), .Y(mai_mai_n2142_));
  NO4        m2093(.A(mai_mai_n677_), .B(mai_mai_n554_), .C(mai_mai_n411_), .D(mai_mai_n949_), .Y(mai_mai_n2143_));
  NO3        m2094(.A(mai_mai_n2143_), .B(mai_mai_n2142_), .C(mai_mai_n955_), .Y(mai_mai_n2144_));
  NA4        m2095(.A(mai_mai_n2144_), .B(mai_mai_n2141_), .C(mai_mai_n2137_), .D(mai_mai_n2132_), .Y(mai_mai_n2145_));
  OR2        m2096(.A(mai_mai_n849_), .B(mai_mai_n692_), .Y(mai_mai_n2146_));
  NA2        m2097(.A(mai_mai_n1071_), .B(mai_mai_n55_), .Y(mai_mai_n2147_));
  NOi21      m2098(.An(mai_mai_n2147_), .B(mai_mai_n362_), .Y(mai_mai_n2148_));
  AOI210     m2099(.A0(mai_mai_n2148_), .A1(mai_mai_n2146_), .B0(x1), .Y(mai_mai_n2149_));
  NA2        m2100(.A(mai_mai_n242_), .B(mai_mai_n84_), .Y(mai_mai_n2150_));
  AOI210     m2101(.A0(mai_mai_n1340_), .A1(mai_mai_n375_), .B0(mai_mai_n2150_), .Y(mai_mai_n2151_));
  NA2        m2102(.A(mai_mai_n1018_), .B(mai_mai_n164_), .Y(mai_mai_n2152_));
  INV        m2103(.A(mai_mai_n2152_), .Y(mai_mai_n2153_));
  NO3        m2104(.A(mai_mai_n2153_), .B(mai_mai_n2151_), .C(mai_mai_n2149_), .Y(mai_mai_n2154_));
  NO2        m2105(.A(mai_mai_n2154_), .B(x6), .Y(mai_mai_n2155_));
  AOI220     m2106(.A0(mai_mai_n2155_), .A1(mai_mai_n1265_), .B0(mai_mai_n2145_), .B1(mai_mai_n57_), .Y(mai_mai_n2156_));
  NA3        m2107(.A(mai_mai_n2156_), .B(mai_mai_n2127_), .C(mai_mai_n2120_), .Y(mai38));
  NO2        m2108(.A(mai_mai_n1433_), .B(mai_mai_n874_), .Y(mai_mai_n2158_));
  AOI210     m2109(.A0(mai_mai_n1072_), .A1(mai_mai_n531_), .B0(mai_mai_n973_), .Y(mai_mai_n2159_));
  NO2        m2110(.A(mai_mai_n2147_), .B(mai_mai_n209_), .Y(mai_mai_n2160_));
  NO3        m2111(.A(mai_mai_n2160_), .B(mai_mai_n2159_), .C(mai_mai_n2158_), .Y(mai_mai_n2161_));
  NO2        m2112(.A(mai_mai_n2161_), .B(x6), .Y(mai_mai_n2162_));
  NA4        m2113(.A(mai_mai_n353_), .B(mai_mai_n234_), .C(mai_mai_n176_), .D(x8), .Y(mai_mai_n2163_));
  NA2        m2114(.A(mai_mai_n374_), .B(mai_mai_n103_), .Y(mai_mai_n2164_));
  AOI210     m2115(.A0(mai_mai_n2164_), .A1(mai_mai_n2163_), .B0(mai_mai_n134_), .Y(mai_mai_n2165_));
  NA2        m2116(.A(mai_mai_n2165_), .B(x6), .Y(mai_mai_n2166_));
  NO2        m2117(.A(x3), .B(mai_mai_n234_), .Y(mai_mai_n2167_));
  OAI210     m2118(.A0(mai_mai_n158_), .A1(mai_mai_n2167_), .B0(mai_mai_n751_), .Y(mai_mai_n2168_));
  NO2        m2119(.A(mai_mai_n554_), .B(mai_mai_n251_), .Y(mai_mai_n2169_));
  NA2        m2120(.A(mai_mai_n2169_), .B(mai_mai_n302_), .Y(mai_mai_n2170_));
  OAI210     m2121(.A0(mai_mai_n630_), .A1(x0), .B0(mai_mai_n51_), .Y(mai_mai_n2171_));
  AOI210     m2122(.A0(mai_mai_n537_), .A1(x4), .B0(mai_mai_n208_), .Y(mai_mai_n2172_));
  NA2        m2123(.A(mai_mai_n2172_), .B(mai_mai_n2171_), .Y(mai_mai_n2173_));
  NA4        m2124(.A(mai_mai_n2173_), .B(mai_mai_n2170_), .C(mai_mai_n2168_), .D(mai_mai_n2166_), .Y(mai_mai_n2174_));
  OAI210     m2125(.A0(mai_mai_n2174_), .A1(mai_mai_n2162_), .B0(x7), .Y(mai_mai_n2175_));
  AOI210     m2126(.A0(mai_mai_n349_), .A1(x1), .B0(mai_mai_n1076_), .Y(mai_mai_n2176_));
  NO2        m2127(.A(mai_mai_n2176_), .B(mai_mai_n51_), .Y(mai_mai_n2177_));
  AOI210     m2128(.A0(mai_mai_n92_), .A1(mai_mai_n71_), .B0(mai_mai_n1887_), .Y(mai_mai_n2178_));
  NA2        m2129(.A(mai_mai_n361_), .B(x3), .Y(mai_mai_n2179_));
  NO2        m2130(.A(mai_mai_n1508_), .B(mai_mai_n490_), .Y(mai_mai_n2180_));
  OAI210     m2131(.A0(mai_mai_n2179_), .A1(mai_mai_n2178_), .B0(mai_mai_n2180_), .Y(mai_mai_n2181_));
  OAI210     m2132(.A0(mai_mai_n2181_), .A1(mai_mai_n2177_), .B0(x4), .Y(mai_mai_n2182_));
  NO2        m2133(.A(mai_mai_n1517_), .B(mai_mai_n427_), .Y(mai_mai_n2183_));
  NO3        m2134(.A(mai_mai_n2183_), .B(mai_mai_n375_), .C(mai_mai_n115_), .Y(mai_mai_n2184_));
  AOI210     m2135(.A0(mai_mai_n949_), .A1(mai_mai_n221_), .B0(mai_mai_n368_), .Y(mai_mai_n2185_));
  AO210      m2136(.A0(mai_mai_n1128_), .A1(x6), .B0(mai_mai_n2185_), .Y(mai_mai_n2186_));
  NO2        m2137(.A(mai_mai_n1223_), .B(mai_mai_n131_), .Y(mai_mai_n2187_));
  NA2        m2138(.A(mai_mai_n1646_), .B(mai_mai_n296_), .Y(mai_mai_n2188_));
  OAI220     m2139(.A0(mai_mai_n2188_), .A1(mai_mai_n967_), .B0(mai_mai_n2187_), .B1(mai_mai_n1567_), .Y(mai_mai_n2189_));
  NO3        m2140(.A(mai_mai_n2189_), .B(mai_mai_n2186_), .C(mai_mai_n2184_), .Y(mai_mai_n2190_));
  AOI210     m2141(.A0(mai_mai_n2190_), .A1(mai_mai_n2182_), .B0(mai_mai_n103_), .Y(mai_mai_n2191_));
  NA3        m2142(.A(mai_mai_n1636_), .B(mai_mai_n554_), .C(mai_mai_n153_), .Y(mai_mai_n2192_));
  AOI210     m2143(.A0(mai_mai_n2192_), .A1(mai_mai_n1232_), .B0(mai_mai_n210_), .Y(mai_mai_n2193_));
  AOI210     m2144(.A0(mai_mai_n465_), .A1(mai_mai_n454_), .B0(mai_mai_n626_), .Y(mai_mai_n2194_));
  OAI220     m2145(.A0(mai_mai_n2194_), .A1(mai_mai_n434_), .B0(mai_mai_n184_), .B1(mai_mai_n114_), .Y(mai_mai_n2195_));
  OAI210     m2146(.A0(mai_mai_n2195_), .A1(mai_mai_n2193_), .B0(x0), .Y(mai_mai_n2196_));
  NA3        m2147(.A(mai_mai_n379_), .B(mai_mai_n755_), .C(mai_mai_n251_), .Y(mai_mai_n2197_));
  AOI210     m2148(.A0(mai_mai_n2197_), .A1(mai_mai_n662_), .B0(mai_mai_n2217_), .Y(mai_mai_n2198_));
  NA2        m2149(.A(mai_mai_n995_), .B(mai_mai_n862_), .Y(mai_mai_n2199_));
  NA2        m2150(.A(mai_mai_n168_), .B(x3), .Y(mai_mai_n2200_));
  AOI210     m2151(.A0(mai_mai_n2200_), .A1(mai_mai_n2199_), .B0(mai_mai_n459_), .Y(mai_mai_n2201_));
  NO4        m2152(.A(mai_mai_n1217_), .B(mai_mai_n480_), .C(mai_mai_n1073_), .D(mai_mai_n713_), .Y(mai_mai_n2202_));
  OAI220     m2153(.A0(mai_mai_n1529_), .A1(mai_mai_n1919_), .B0(mai_mai_n208_), .B1(mai_mai_n141_), .Y(mai_mai_n2203_));
  NO4        m2154(.A(mai_mai_n2203_), .B(mai_mai_n2202_), .C(mai_mai_n2201_), .D(mai_mai_n2198_), .Y(mai_mai_n2204_));
  NA2        m2155(.A(mai_mai_n2204_), .B(mai_mai_n2196_), .Y(mai_mai_n2205_));
  OAI210     m2156(.A0(mai_mai_n2205_), .A1(mai_mai_n2191_), .B0(mai_mai_n57_), .Y(mai_mai_n2206_));
  AOI210     m2157(.A0(mai_mai_n1561_), .A1(mai_mai_n251_), .B0(mai_mai_n627_), .Y(mai_mai_n2207_));
  OAI210     m2158(.A0(mai_mai_n1515_), .A1(mai_mai_n197_), .B0(mai_mai_n456_), .Y(mai_mai_n2208_));
  OAI210     m2159(.A0(mai_mai_n2208_), .A1(mai_mai_n2207_), .B0(mai_mai_n577_), .Y(mai_mai_n2209_));
  NA2        m2160(.A(mai_mai_n1593_), .B(mai_mai_n329_), .Y(mai_mai_n2210_));
  OAI220     m2161(.A0(mai_mai_n2210_), .A1(mai_mai_n584_), .B0(mai_mai_n637_), .B1(mai_mai_n141_), .Y(mai_mai_n2211_));
  INV        m2162(.A(mai_mai_n2211_), .Y(mai_mai_n2212_));
  NA4        m2163(.A(mai_mai_n2212_), .B(mai_mai_n2209_), .C(mai_mai_n2206_), .D(mai_mai_n2175_), .Y(mai39));
  INV        m2164(.A(x1), .Y(mai_mai_n2216_));
  INV        m2165(.A(mai_mai_n906_), .Y(mai_mai_n2217_));
  INV        m2166(.A(x4), .Y(mai_mai_n2218_));
  INV        m2167(.A(mai_mai_n1367_), .Y(mai_mai_n2219_));
  INV        m2168(.A(x7), .Y(mai_mai_n2220_));
  INV        m2169(.A(x4), .Y(mai_mai_n2221_));
  INV        m2170(.A(x1), .Y(mai_mai_n2222_));
  INV        m2171(.A(x7), .Y(mai_mai_n2223_));
  INV        m2172(.A(mai_mai_n610_), .Y(mai_mai_n2224_));
  INV        u0000(.A(x3), .Y(men_men_n50_));
  NA2        u0001(.A(men_men_n50_), .B(x2), .Y(men_men_n51_));
  NA2        u0002(.A(x7), .B(x0), .Y(men_men_n52_));
  INV        u0003(.A(x1), .Y(men_men_n53_));
  NA2        u0004(.A(x5), .B(men_men_n53_), .Y(men_men_n54_));
  INV        u0005(.A(x8), .Y(men_men_n55_));
  INV        u0006(.A(x4), .Y(men_men_n56_));
  INV        u0007(.A(x7), .Y(men_men_n57_));
  NA2        u0008(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0009(.A(x0), .Y(men_men_n59_));
  NA2        u0010(.A(x4), .B(men_men_n59_), .Y(men_men_n60_));
  NA2        u0011(.A(men_men_n56_), .B(men_men_n59_), .Y(men_men_n61_));
  NO2        u0012(.A(men_men_n55_), .B(x6), .Y(men_men_n62_));
  NA2        u0013(.A(men_men_n57_), .B(x4), .Y(men_men_n63_));
  NO2        u0014(.A(x8), .B(men_men_n57_), .Y(men_men_n64_));
  NO2        u0015(.A(x7), .B(men_men_n59_), .Y(men_men_n65_));
  NAi21      u0016(.An(x5), .B(x1), .Y(men_men_n66_));
  INV        u0017(.A(x6), .Y(men_men_n67_));
  NA2        u0018(.A(men_men_n67_), .B(x4), .Y(men_men_n68_));
  NA2        u0019(.A(x7), .B(x4), .Y(men_men_n69_));
  NO2        u0020(.A(men_men_n69_), .B(x1), .Y(men_men_n70_));
  NO2        u0021(.A(men_men_n67_), .B(x5), .Y(men_men_n71_));
  NO2        u0022(.A(x8), .B(men_men_n59_), .Y(men_men_n72_));
  NA2        u0023(.A(x5), .B(x3), .Y(men_men_n73_));
  NO2        u0024(.A(x6), .B(x0), .Y(men_men_n74_));
  NO2        u0025(.A(men_men_n74_), .B(x4), .Y(men_men_n75_));
  NO2        u0026(.A(x4), .B(x2), .Y(men_men_n76_));
  NO2        u0027(.A(men_men_n67_), .B(men_men_n59_), .Y(men_men_n77_));
  NO2        u0028(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NA2        u0029(.A(x8), .B(x1), .Y(men_men_n79_));
  NO2        u0030(.A(men_men_n79_), .B(x7), .Y(men_men_n80_));
  OR3        u0031(.A(men_men_n79_), .B(men_men_n78_), .C(men_men_n75_), .Y(men_men_n81_));
  NO3        u0032(.A(x8), .B(men_men_n57_), .C(x6), .Y(men_men_n82_));
  NO2        u0033(.A(x1), .B(men_men_n59_), .Y(men_men_n83_));
  NO2        u0034(.A(men_men_n56_), .B(x2), .Y(men_men_n84_));
  NA2        u0035(.A(men_men_n83_), .B(men_men_n82_), .Y(men_men_n85_));
  AOI210     u0036(.A0(men_men_n85_), .A1(men_men_n81_), .B0(men_men_n73_), .Y(men_men_n86_));
  XO2        u0037(.A(x7), .B(x1), .Y(men_men_n87_));
  NO2        u0038(.A(men_men_n50_), .B(x0), .Y(men_men_n88_));
  NA2        u0039(.A(men_men_n88_), .B(men_men_n55_), .Y(men_men_n89_));
  NO2        u0040(.A(x6), .B(x5), .Y(men_men_n90_));
  NO2        u0041(.A(men_men_n57_), .B(x5), .Y(men_men_n91_));
  NO2        u0042(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n92_));
  NA2        u0043(.A(x6), .B(x1), .Y(men_men_n93_));
  NA2        u0044(.A(men_men_n93_), .B(men_men_n76_), .Y(men_men_n94_));
  NO3        u0045(.A(men_men_n94_), .B(men_men_n92_), .C(men_men_n89_), .Y(men_men_n95_));
  NA2        u0046(.A(x3), .B(x0), .Y(men_men_n96_));
  INV        u0047(.A(x5), .Y(men_men_n97_));
  NA2        u0048(.A(men_men_n67_), .B(men_men_n97_), .Y(men_men_n98_));
  INV        u0049(.A(x2), .Y(men_men_n99_));
  NO2        u0050(.A(men_men_n56_), .B(men_men_n99_), .Y(men_men_n100_));
  NA2        u0051(.A(men_men_n57_), .B(men_men_n97_), .Y(men_men_n101_));
  NA3        u0052(.A(men_men_n101_), .B(men_men_n100_), .C(men_men_n98_), .Y(men_men_n102_));
  NO3        u0053(.A(men_men_n102_), .B(men_men_n96_), .C(men_men_n53_), .Y(men_men_n103_));
  NO3        u0054(.A(men_men_n103_), .B(men_men_n95_), .C(men_men_n86_), .Y(men00));
  NO2        u0055(.A(x7), .B(x6), .Y(men_men_n105_));
  NO2        u0056(.A(men_men_n55_), .B(men_men_n53_), .Y(men_men_n106_));
  NA2        u0057(.A(men_men_n106_), .B(men_men_n56_), .Y(men_men_n107_));
  NO2        u0058(.A(men_men_n107_), .B(x6), .Y(men_men_n108_));
  XN2        u0059(.A(x6), .B(x1), .Y(men_men_n109_));
  INV        u0060(.A(men_men_n109_), .Y(men_men_n110_));
  NO2        u0061(.A(x6), .B(x4), .Y(men_men_n111_));
  NA2        u0062(.A(x6), .B(x4), .Y(men_men_n112_));
  XN2        u0063(.A(x7), .B(x6), .Y(men_men_n113_));
  NO4        u0064(.A(men_men_n113_), .B(men_men_n111_), .C(men_men_n110_), .D(x8), .Y(men_men_n114_));
  NO2        u0065(.A(x3), .B(men_men_n99_), .Y(men_men_n115_));
  NA2        u0066(.A(men_men_n115_), .B(men_men_n97_), .Y(men_men_n116_));
  NO2        u0067(.A(men_men_n116_), .B(men_men_n59_), .Y(men_men_n117_));
  OAI210     u0068(.A0(men_men_n114_), .A1(men_men_n108_), .B0(men_men_n117_), .Y(men_men_n118_));
  NA2        u0069(.A(x3), .B(men_men_n99_), .Y(men_men_n119_));
  NO2        u0070(.A(men_men_n55_), .B(men_men_n57_), .Y(men_men_n120_));
  NA2        u0071(.A(men_men_n120_), .B(men_men_n56_), .Y(men_men_n121_));
  NA2        u0072(.A(men_men_n55_), .B(men_men_n57_), .Y(men_men_n122_));
  NA2        u0073(.A(men_men_n122_), .B(x2), .Y(men_men_n123_));
  NA2        u0074(.A(x8), .B(x3), .Y(men_men_n124_));
  NA2        u0075(.A(men_men_n124_), .B(men_men_n69_), .Y(men_men_n125_));
  OAI220     u0076(.A0(men_men_n125_), .A1(men_men_n123_), .B0(men_men_n121_), .B1(men_men_n119_), .Y(men_men_n126_));
  NO2        u0077(.A(x5), .B(x0), .Y(men_men_n127_));
  NO2        u0078(.A(x6), .B(x1), .Y(men_men_n128_));
  NA3        u0079(.A(men_men_n128_), .B(men_men_n127_), .C(men_men_n126_), .Y(men_men_n129_));
  NA2        u0080(.A(x8), .B(men_men_n97_), .Y(men_men_n130_));
  NA2        u0081(.A(x4), .B(men_men_n50_), .Y(men_men_n131_));
  NO3        u0082(.A(men_men_n131_), .B(men_men_n130_), .C(men_men_n93_), .Y(men_men_n132_));
  NAi21      u0083(.An(x7), .B(x2), .Y(men_men_n133_));
  NO2        u0084(.A(men_men_n133_), .B(x0), .Y(men_men_n134_));
  XO2        u0085(.A(x8), .B(x7), .Y(men_men_n135_));
  NA2        u0086(.A(men_men_n135_), .B(men_men_n99_), .Y(men_men_n136_));
  NA2        u0087(.A(x6), .B(x5), .Y(men_men_n137_));
  NO2        u0088(.A(men_men_n56_), .B(x0), .Y(men_men_n138_));
  NO2        u0089(.A(men_men_n50_), .B(x1), .Y(men_men_n139_));
  NA2        u0090(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NO3        u0091(.A(men_men_n140_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n141_));
  AOI210     u0092(.A0(men_men_n134_), .A1(men_men_n132_), .B0(men_men_n141_), .Y(men_men_n142_));
  NA3        u0093(.A(men_men_n142_), .B(men_men_n129_), .C(men_men_n118_), .Y(men01));
  NA2        u0094(.A(men_men_n57_), .B(men_men_n59_), .Y(men_men_n144_));
  NO2        u0095(.A(x2), .B(x1), .Y(men_men_n145_));
  NA2        u0096(.A(x2), .B(x1), .Y(men_men_n146_));
  NOi21      u0097(.An(men_men_n146_), .B(men_men_n145_), .Y(men_men_n147_));
  NA2        u0098(.A(men_men_n97_), .B(men_men_n53_), .Y(men_men_n148_));
  NO2        u0099(.A(men_men_n148_), .B(x8), .Y(men_men_n149_));
  NAi21      u0100(.An(x8), .B(x1), .Y(men_men_n150_));
  NO2        u0101(.A(men_men_n150_), .B(x3), .Y(men_men_n151_));
  OAI210     u0102(.A0(men_men_n151_), .A1(men_men_n149_), .B0(men_men_n147_), .Y(men_men_n152_));
  NO2        u0103(.A(x5), .B(men_men_n50_), .Y(men_men_n153_));
  NO2        u0104(.A(men_men_n99_), .B(x1), .Y(men_men_n154_));
  NA2        u0105(.A(men_men_n154_), .B(men_men_n153_), .Y(men_men_n155_));
  AOI210     u0106(.A0(men_men_n155_), .A1(men_men_n152_), .B0(men_men_n144_), .Y(men_men_n156_));
  NAi21      u0107(.An(x7), .B(x0), .Y(men_men_n157_));
  NO2        u0108(.A(men_men_n55_), .B(x2), .Y(men_men_n158_));
  NO2        u0109(.A(men_men_n73_), .B(x1), .Y(men_men_n159_));
  NA2        u0110(.A(x5), .B(men_men_n50_), .Y(men_men_n160_));
  NO2        u0111(.A(men_men_n160_), .B(men_men_n150_), .Y(men_men_n161_));
  NA2        u0112(.A(x8), .B(x5), .Y(men_men_n162_));
  NO2        u0113(.A(men_men_n162_), .B(men_men_n51_), .Y(men_men_n163_));
  NO3        u0114(.A(x3), .B(men_men_n99_), .C(men_men_n53_), .Y(men_men_n164_));
  NO3        u0115(.A(men_men_n164_), .B(men_men_n163_), .C(men_men_n161_), .Y(men_men_n165_));
  NO2        u0116(.A(men_men_n165_), .B(men_men_n157_), .Y(men_men_n166_));
  NO2        u0117(.A(men_men_n57_), .B(x3), .Y(men_men_n167_));
  NO2        u0118(.A(men_men_n55_), .B(x0), .Y(men_men_n168_));
  NA3        u0119(.A(men_men_n97_), .B(men_men_n99_), .C(x1), .Y(men_men_n169_));
  NO2        u0120(.A(men_men_n169_), .B(men_men_n168_), .Y(men_men_n170_));
  NO2        u0121(.A(men_men_n79_), .B(men_men_n50_), .Y(men_men_n171_));
  NA2        u0122(.A(men_men_n97_), .B(x0), .Y(men_men_n172_));
  NO2        u0123(.A(men_men_n172_), .B(x2), .Y(men_men_n173_));
  AOI220     u0124(.A0(men_men_n173_), .A1(men_men_n171_), .B0(men_men_n170_), .B1(men_men_n167_), .Y(men_men_n174_));
  NA2        u0125(.A(x7), .B(men_men_n99_), .Y(men_men_n175_));
  NA2        u0126(.A(men_men_n153_), .B(x8), .Y(men_men_n176_));
  NA4        u0127(.A(x5), .B(x3), .C(x1), .D(x0), .Y(men_men_n177_));
  AO210      u0128(.A0(men_men_n177_), .A1(men_men_n176_), .B0(men_men_n175_), .Y(men_men_n178_));
  NAi21      u0129(.An(x1), .B(x2), .Y(men_men_n179_));
  NO2        u0130(.A(men_men_n160_), .B(men_men_n179_), .Y(men_men_n180_));
  NA2        u0131(.A(x8), .B(x7), .Y(men_men_n181_));
  NA2        u0132(.A(men_men_n178_), .B(men_men_n174_), .Y(men_men_n182_));
  NO3        u0133(.A(men_men_n182_), .B(men_men_n166_), .C(men_men_n156_), .Y(men_men_n183_));
  NA2        u0134(.A(x3), .B(x1), .Y(men_men_n184_));
  NA2        u0135(.A(men_men_n50_), .B(men_men_n99_), .Y(men_men_n185_));
  NO2        u0136(.A(men_men_n185_), .B(men_men_n66_), .Y(men_men_n186_));
  OAI210     u0137(.A0(men_men_n186_), .A1(men_men_n180_), .B0(men_men_n64_), .Y(men_men_n187_));
  NA2        u0138(.A(men_men_n120_), .B(men_men_n99_), .Y(men_men_n188_));
  OAI210     u0139(.A0(men_men_n188_), .A1(men_men_n184_), .B0(men_men_n187_), .Y(men_men_n189_));
  XO2        u0140(.A(x5), .B(x3), .Y(men_men_n190_));
  NA2        u0141(.A(men_men_n190_), .B(x8), .Y(men_men_n191_));
  NA2        u0142(.A(x8), .B(men_men_n59_), .Y(men_men_n192_));
  NA2        u0143(.A(x7), .B(men_men_n67_), .Y(men_men_n193_));
  NA2        u0144(.A(men_men_n189_), .B(x0), .Y(men_men_n194_));
  OAI210     u0145(.A0(men_men_n183_), .A1(men_men_n67_), .B0(men_men_n194_), .Y(men_men_n195_));
  NO2        u0146(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n196_));
  NA2        u0147(.A(x8), .B(men_men_n50_), .Y(men_men_n197_));
  NA2        u0148(.A(men_men_n197_), .B(x2), .Y(men_men_n198_));
  NA2        u0149(.A(men_men_n55_), .B(x3), .Y(men_men_n199_));
  NO2        u0150(.A(men_men_n99_), .B(men_men_n59_), .Y(men_men_n200_));
  NA2        u0151(.A(x5), .B(x1), .Y(men_men_n201_));
  NO2        u0152(.A(men_men_n201_), .B(x6), .Y(men_men_n202_));
  NO2        u0153(.A(x3), .B(x1), .Y(men_men_n203_));
  NO2        u0154(.A(men_men_n73_), .B(men_men_n55_), .Y(men_men_n204_));
  NO2        u0155(.A(men_men_n93_), .B(men_men_n50_), .Y(men_men_n205_));
  NO2        u0156(.A(men_men_n205_), .B(men_men_n204_), .Y(men_men_n206_));
  INV        u0157(.A(men_men_n206_), .Y(men_men_n207_));
  NO2        u0158(.A(men_men_n55_), .B(x5), .Y(men_men_n208_));
  NA2        u0159(.A(men_men_n208_), .B(men_men_n67_), .Y(men_men_n209_));
  NAi21      u0160(.An(x2), .B(x5), .Y(men_men_n210_));
  NA2        u0161(.A(x8), .B(x6), .Y(men_men_n211_));
  NA2        u0162(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n212_));
  AN2        u0163(.A(men_men_n207_), .B(men_men_n200_), .Y(men_men_n213_));
  NA2        u0164(.A(men_men_n213_), .B(men_men_n196_), .Y(men_men_n214_));
  NA2        u0165(.A(men_men_n67_), .B(men_men_n56_), .Y(men_men_n215_));
  NO2        u0166(.A(men_men_n215_), .B(x7), .Y(men_men_n216_));
  NO2        u0167(.A(men_men_n97_), .B(men_men_n53_), .Y(men_men_n217_));
  NA2        u0168(.A(men_men_n217_), .B(men_men_n99_), .Y(men_men_n218_));
  NA2        u0169(.A(x3), .B(men_men_n59_), .Y(men_men_n219_));
  NO2        u0170(.A(men_men_n169_), .B(men_men_n219_), .Y(men_men_n220_));
  NO2        u0171(.A(x1), .B(x0), .Y(men_men_n221_));
  NA2        u0172(.A(men_men_n221_), .B(men_men_n99_), .Y(men_men_n222_));
  NA2        u0173(.A(men_men_n97_), .B(men_men_n50_), .Y(men_men_n223_));
  XN2        u0174(.A(x3), .B(x2), .Y(men_men_n224_));
  NA2        u0175(.A(men_men_n224_), .B(men_men_n147_), .Y(men_men_n225_));
  NO2        u0176(.A(men_men_n97_), .B(x0), .Y(men_men_n226_));
  NA2        u0177(.A(x8), .B(men_men_n53_), .Y(men_men_n227_));
  NA2        u0178(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n228_));
  OAI220     u0179(.A0(men_men_n228_), .A1(men_men_n225_), .B0(men_men_n223_), .B1(men_men_n222_), .Y(men_men_n229_));
  NA2        u0180(.A(men_men_n229_), .B(men_men_n216_), .Y(men_men_n230_));
  NO2        u0181(.A(x7), .B(x1), .Y(men_men_n231_));
  NOi21      u0182(.An(x8), .B(x3), .Y(men_men_n232_));
  NA2        u0183(.A(men_men_n232_), .B(men_men_n59_), .Y(men_men_n233_));
  NA2        u0184(.A(x5), .B(x0), .Y(men_men_n234_));
  NAi21      u0185(.An(men_men_n127_), .B(men_men_n234_), .Y(men_men_n235_));
  NA2        u0186(.A(men_men_n67_), .B(men_men_n50_), .Y(men_men_n236_));
  NA2        u0187(.A(x8), .B(men_men_n57_), .Y(men_men_n237_));
  NO2        u0188(.A(men_men_n237_), .B(x5), .Y(men_men_n238_));
  NO2        u0189(.A(men_men_n139_), .B(men_men_n67_), .Y(men_men_n239_));
  NA2        u0190(.A(x1), .B(x0), .Y(men_men_n240_));
  NA2        u0191(.A(men_men_n50_), .B(men_men_n59_), .Y(men_men_n241_));
  NA4        u0192(.A(men_men_n241_), .B(men_men_n240_), .C(men_men_n239_), .D(men_men_n238_), .Y(men_men_n242_));
  NA2        u0193(.A(men_men_n242_), .B(men_men_n177_), .Y(men_men_n243_));
  NO2        u0194(.A(men_men_n97_), .B(x3), .Y(men_men_n244_));
  NO2        u0195(.A(men_men_n99_), .B(x0), .Y(men_men_n245_));
  NA2        u0196(.A(men_men_n245_), .B(men_men_n244_), .Y(men_men_n246_));
  NO2        u0197(.A(men_men_n55_), .B(x7), .Y(men_men_n247_));
  NO3        u0198(.A(x8), .B(men_men_n50_), .C(x0), .Y(men_men_n248_));
  NAi21      u0199(.An(x8), .B(x0), .Y(men_men_n249_));
  NAi21      u0200(.An(x1), .B(x3), .Y(men_men_n250_));
  NO2        u0201(.A(men_men_n250_), .B(men_men_n249_), .Y(men_men_n251_));
  NO2        u0202(.A(x2), .B(men_men_n53_), .Y(men_men_n252_));
  NOi21      u0203(.An(x5), .B(x6), .Y(men_men_n253_));
  NO2        u0204(.A(men_men_n57_), .B(x4), .Y(men_men_n254_));
  NO2        u0205(.A(men_men_n2316_), .B(men_men_n246_), .Y(men_men_n255_));
  AOI210     u0206(.A0(men_men_n243_), .A1(men_men_n100_), .B0(men_men_n255_), .Y(men_men_n256_));
  NA3        u0207(.A(men_men_n256_), .B(men_men_n230_), .C(men_men_n214_), .Y(men_men_n257_));
  AOI210     u0208(.A0(men_men_n195_), .A1(men_men_n56_), .B0(men_men_n257_), .Y(men02));
  NO2        u0209(.A(x8), .B(men_men_n97_), .Y(men_men_n259_));
  XN2        u0210(.A(x7), .B(x3), .Y(men_men_n260_));
  INV        u0211(.A(men_men_n260_), .Y(men_men_n261_));
  NO2        u0212(.A(x2), .B(x0), .Y(men_men_n262_));
  NA2        u0213(.A(men_men_n262_), .B(men_men_n67_), .Y(men_men_n263_));
  NO2        u0214(.A(men_men_n57_), .B(x1), .Y(men_men_n264_));
  NO3        u0215(.A(men_men_n264_), .B(men_men_n263_), .C(men_men_n261_), .Y(men_men_n265_));
  NA2        u0216(.A(men_men_n53_), .B(x0), .Y(men_men_n266_));
  NO2        u0217(.A(men_men_n250_), .B(x6), .Y(men_men_n267_));
  XO2        u0218(.A(x7), .B(x0), .Y(men_men_n268_));
  NO2        u0219(.A(men_men_n268_), .B(men_men_n262_), .Y(men_men_n269_));
  NA2        u0220(.A(men_men_n269_), .B(men_men_n267_), .Y(men_men_n270_));
  AN2        u0221(.A(x7), .B(x2), .Y(men_men_n271_));
  NA2        u0222(.A(men_men_n271_), .B(men_men_n50_), .Y(men_men_n272_));
  NA2        u0223(.A(men_men_n272_), .B(men_men_n270_), .Y(men_men_n273_));
  OAI210     u0224(.A0(men_men_n273_), .A1(men_men_n265_), .B0(men_men_n259_), .Y(men_men_n274_));
  NAi21      u0225(.An(x8), .B(x6), .Y(men_men_n275_));
  NO2        u0226(.A(men_men_n97_), .B(men_men_n59_), .Y(men_men_n276_));
  NA2        u0227(.A(x7), .B(x3), .Y(men_men_n277_));
  NO2        u0228(.A(men_men_n277_), .B(x2), .Y(men_men_n278_));
  NA2        u0229(.A(x2), .B(x0), .Y(men_men_n279_));
  NA2        u0230(.A(men_men_n99_), .B(men_men_n59_), .Y(men_men_n280_));
  NA2        u0231(.A(men_men_n280_), .B(men_men_n279_), .Y(men_men_n281_));
  NAi21      u0232(.An(x7), .B(x1), .Y(men_men_n282_));
  NO2        u0233(.A(men_men_n282_), .B(x3), .Y(men_men_n283_));
  AOI220     u0234(.A0(men_men_n283_), .A1(men_men_n281_), .B0(men_men_n278_), .B1(men_men_n276_), .Y(men_men_n284_));
  NA2        u0235(.A(men_men_n252_), .B(men_men_n50_), .Y(men_men_n285_));
  NA3        u0236(.A(x7), .B(men_men_n97_), .C(x0), .Y(men_men_n286_));
  NA2        u0237(.A(men_men_n245_), .B(men_men_n53_), .Y(men_men_n287_));
  NA2        u0238(.A(men_men_n153_), .B(men_men_n57_), .Y(men_men_n288_));
  OA220      u0239(.A0(men_men_n288_), .A1(men_men_n287_), .B0(men_men_n286_), .B1(men_men_n285_), .Y(men_men_n289_));
  AOI210     u0240(.A0(men_men_n289_), .A1(men_men_n284_), .B0(men_men_n275_), .Y(men_men_n290_));
  INV        u0241(.A(men_men_n268_), .Y(men_men_n291_));
  NO2        u0242(.A(x7), .B(men_men_n67_), .Y(men_men_n292_));
  NA2        u0243(.A(men_men_n97_), .B(x3), .Y(men_men_n293_));
  NO2        u0244(.A(men_men_n293_), .B(men_men_n292_), .Y(men_men_n294_));
  NA2        u0245(.A(men_men_n50_), .B(x0), .Y(men_men_n295_));
  NO2        u0246(.A(men_men_n57_), .B(men_men_n50_), .Y(men_men_n296_));
  NO2        u0247(.A(men_men_n55_), .B(men_men_n99_), .Y(men_men_n297_));
  NA3        u0248(.A(men_men_n297_), .B(men_men_n296_), .C(men_men_n59_), .Y(men_men_n298_));
  NO2        u0249(.A(men_men_n148_), .B(x6), .Y(men_men_n299_));
  NO2        u0250(.A(men_men_n93_), .B(men_men_n97_), .Y(men_men_n300_));
  NA2        u0251(.A(men_men_n57_), .B(men_men_n99_), .Y(men_men_n301_));
  NO2        u0252(.A(men_men_n301_), .B(men_men_n241_), .Y(men_men_n302_));
  OAI210     u0253(.A0(men_men_n300_), .A1(men_men_n299_), .B0(men_men_n302_), .Y(men_men_n303_));
  INV        u0254(.A(men_men_n303_), .Y(men_men_n304_));
  NO2        u0255(.A(men_men_n304_), .B(men_men_n290_), .Y(men_men_n305_));
  AOI210     u0256(.A0(men_men_n305_), .A1(men_men_n274_), .B0(x4), .Y(men_men_n306_));
  NA2        u0257(.A(x8), .B(men_men_n67_), .Y(men_men_n307_));
  NO2        u0258(.A(x3), .B(men_men_n59_), .Y(men_men_n308_));
  NO2        u0259(.A(x3), .B(x0), .Y(men_men_n309_));
  NAi21      u0260(.An(men_men_n309_), .B(men_men_n96_), .Y(men_men_n310_));
  NA2        u0261(.A(x5), .B(x2), .Y(men_men_n311_));
  INV        u0262(.A(men_men_n311_), .Y(men_men_n312_));
  NO2        u0263(.A(men_men_n99_), .B(men_men_n53_), .Y(men_men_n313_));
  NO2        u0264(.A(men_men_n55_), .B(x1), .Y(men_men_n314_));
  NA2        u0265(.A(men_men_n314_), .B(men_men_n99_), .Y(men_men_n315_));
  NO2        u0266(.A(men_men_n50_), .B(x2), .Y(men_men_n316_));
  NAi21      u0267(.An(x6), .B(x5), .Y(men_men_n317_));
  NO2        u0268(.A(x2), .B(men_men_n59_), .Y(men_men_n318_));
  NA2        u0269(.A(men_men_n313_), .B(men_men_n77_), .Y(men_men_n319_));
  NO2        u0270(.A(men_men_n319_), .B(men_men_n69_), .Y(men_men_n320_));
  NO2        u0271(.A(men_men_n97_), .B(men_men_n50_), .Y(men_men_n321_));
  NO2        u0272(.A(men_men_n262_), .B(men_men_n200_), .Y(men_men_n322_));
  XO2        u0273(.A(x7), .B(x2), .Y(men_men_n323_));
  INV        u0274(.A(men_men_n323_), .Y(men_men_n324_));
  XO2        u0275(.A(x6), .B(x2), .Y(men_men_n325_));
  NAi21      u0276(.An(x0), .B(x6), .Y(men_men_n326_));
  NA2        u0277(.A(x7), .B(x5), .Y(men_men_n327_));
  NO2        u0278(.A(x8), .B(x6), .Y(men_men_n328_));
  NAi21      u0279(.An(men_men_n328_), .B(men_men_n211_), .Y(men_men_n329_));
  NO2        u0280(.A(men_men_n83_), .B(x3), .Y(men_men_n330_));
  NA2        u0281(.A(men_men_n97_), .B(x2), .Y(men_men_n331_));
  NO2        u0282(.A(men_men_n331_), .B(men_men_n63_), .Y(men_men_n332_));
  NA2        u0283(.A(x1), .B(men_men_n59_), .Y(men_men_n333_));
  NO2        u0284(.A(men_men_n333_), .B(men_men_n211_), .Y(men_men_n334_));
  OAI210     u0285(.A0(men_men_n334_), .A1(men_men_n50_), .B0(men_men_n332_), .Y(men_men_n335_));
  NA2        u0286(.A(x4), .B(x2), .Y(men_men_n336_));
  NO2        u0287(.A(men_men_n336_), .B(men_men_n97_), .Y(men_men_n337_));
  NAi21      u0288(.An(x1), .B(x6), .Y(men_men_n338_));
  NO2        u0289(.A(men_men_n96_), .B(men_men_n53_), .Y(men_men_n339_));
  NA2        u0290(.A(x8), .B(x2), .Y(men_men_n340_));
  NO2        u0291(.A(men_men_n340_), .B(men_men_n50_), .Y(men_men_n341_));
  INV        u0292(.A(men_men_n202_), .Y(men_men_n342_));
  NO2        u0293(.A(men_men_n342_), .B(men_men_n52_), .Y(men_men_n343_));
  AOI220     u0294(.A0(men_men_n343_), .A1(men_men_n341_), .B0(men_men_n339_), .B1(men_men_n337_), .Y(men_men_n344_));
  OAI210     u0295(.A0(men_men_n335_), .A1(men_men_n330_), .B0(men_men_n344_), .Y(men_men_n345_));
  NO3        u0296(.A(men_men_n345_), .B(men_men_n320_), .C(men_men_n306_), .Y(men03));
  NAi21      u0297(.An(x2), .B(x0), .Y(men_men_n347_));
  NO3        u0298(.A(x8), .B(x6), .C(x4), .Y(men_men_n348_));
  INV        u0299(.A(men_men_n348_), .Y(men_men_n349_));
  NO2        u0300(.A(men_men_n349_), .B(men_men_n347_), .Y(men_men_n350_));
  NA2        u0301(.A(men_men_n100_), .B(men_men_n59_), .Y(men_men_n351_));
  NA2        u0302(.A(men_men_n350_), .B(men_men_n153_), .Y(men_men_n352_));
  NA2        u0303(.A(x3), .B(x2), .Y(men_men_n353_));
  NA2        u0304(.A(x8), .B(x0), .Y(men_men_n354_));
  NO2        u0305(.A(men_men_n354_), .B(x6), .Y(men_men_n355_));
  NO2        u0306(.A(x5), .B(men_men_n59_), .Y(men_men_n356_));
  NO2        u0307(.A(x3), .B(x2), .Y(men_men_n357_));
  NA2        u0308(.A(men_men_n357_), .B(men_men_n356_), .Y(men_men_n358_));
  NO2        u0309(.A(men_men_n53_), .B(x0), .Y(men_men_n359_));
  NA2        u0310(.A(men_men_n359_), .B(x5), .Y(men_men_n360_));
  AOI210     u0311(.A0(men_men_n360_), .A1(men_men_n358_), .B0(men_men_n275_), .Y(men_men_n361_));
  INV        u0312(.A(men_men_n233_), .Y(men_men_n362_));
  NO2        u0313(.A(men_men_n50_), .B(men_men_n59_), .Y(men_men_n363_));
  NO2        u0314(.A(men_men_n67_), .B(x0), .Y(men_men_n364_));
  NO3        u0315(.A(men_men_n364_), .B(x2), .C(men_men_n53_), .Y(men_men_n365_));
  AO210      u0316(.A0(men_men_n365_), .A1(men_men_n362_), .B0(men_men_n361_), .Y(men_men_n366_));
  NA2        u0317(.A(men_men_n366_), .B(x4), .Y(men_men_n367_));
  NO2        u0318(.A(x4), .B(men_men_n53_), .Y(men_men_n368_));
  NA2        u0319(.A(men_men_n368_), .B(men_men_n59_), .Y(men_men_n369_));
  NO3        u0320(.A(men_men_n369_), .B(men_men_n211_), .C(x5), .Y(men_men_n370_));
  NA2        u0321(.A(x7), .B(men_men_n97_), .Y(men_men_n371_));
  NO3        u0322(.A(x5), .B(men_men_n53_), .C(x0), .Y(men_men_n372_));
  INV        u0323(.A(men_men_n372_), .Y(men_men_n373_));
  NO2        u0324(.A(x6), .B(men_men_n56_), .Y(men_men_n374_));
  NO2        u0325(.A(x8), .B(men_men_n50_), .Y(men_men_n375_));
  NA2        u0326(.A(men_men_n375_), .B(men_men_n374_), .Y(men_men_n376_));
  OAI210     u0327(.A0(men_men_n376_), .A1(men_men_n373_), .B0(men_men_n371_), .Y(men_men_n377_));
  AOI210     u0328(.A0(men_men_n370_), .A1(x2), .B0(men_men_n377_), .Y(men_men_n378_));
  AOI220     u0329(.A0(men_men_n378_), .A1(men_men_n367_), .B0(men_men_n352_), .B1(x7), .Y(men_men_n379_));
  NA2        u0330(.A(x7), .B(men_men_n53_), .Y(men_men_n380_));
  NO2        u0331(.A(men_men_n232_), .B(men_men_n99_), .Y(men_men_n381_));
  NO2        u0332(.A(men_men_n55_), .B(men_men_n59_), .Y(men_men_n382_));
  NO3        u0333(.A(men_men_n382_), .B(men_men_n381_), .C(men_men_n137_), .Y(men_men_n383_));
  AOI210     u0334(.A0(x8), .A1(men_men_n90_), .B0(men_men_n383_), .Y(men_men_n384_));
  NO2        u0335(.A(x5), .B(x2), .Y(men_men_n385_));
  NO2        u0336(.A(x8), .B(x3), .Y(men_men_n386_));
  NA2        u0337(.A(men_men_n386_), .B(men_men_n385_), .Y(men_men_n387_));
  NO2        u0338(.A(men_men_n387_), .B(x6), .Y(men_men_n388_));
  AOI210     u0339(.A0(men_men_n2315_), .A1(x8), .B0(men_men_n388_), .Y(men_men_n389_));
  OAI210     u0340(.A0(men_men_n384_), .A1(men_men_n262_), .B0(men_men_n389_), .Y(men_men_n390_));
  NA2        u0341(.A(men_men_n390_), .B(x4), .Y(men_men_n391_));
  NA2        u0342(.A(men_men_n55_), .B(men_men_n59_), .Y(men_men_n392_));
  NO2        u0343(.A(men_men_n392_), .B(x5), .Y(men_men_n393_));
  NAi21      u0344(.An(x4), .B(x6), .Y(men_men_n394_));
  INV        u0345(.A(men_men_n51_), .Y(men_men_n395_));
  NO2        u0346(.A(men_men_n55_), .B(men_men_n67_), .Y(men_men_n396_));
  NO2        u0347(.A(men_men_n50_), .B(men_men_n99_), .Y(men_men_n397_));
  NA2        u0348(.A(men_men_n395_), .B(men_men_n393_), .Y(men_men_n398_));
  AOI210     u0349(.A0(men_men_n398_), .A1(men_men_n391_), .B0(men_men_n380_), .Y(men_men_n399_));
  NA2        u0350(.A(men_men_n57_), .B(men_men_n53_), .Y(men_men_n400_));
  NO2        u0351(.A(men_men_n67_), .B(men_men_n56_), .Y(men_men_n401_));
  NA2        u0352(.A(men_men_n316_), .B(men_men_n59_), .Y(men_men_n402_));
  OAI220     u0353(.A0(men_men_n402_), .A1(men_men_n55_), .B0(men_men_n185_), .B1(men_men_n249_), .Y(men_men_n403_));
  NA2        u0354(.A(men_men_n403_), .B(men_men_n401_), .Y(men_men_n404_));
  NO3        u0355(.A(x6), .B(x4), .C(men_men_n50_), .Y(men_men_n405_));
  NA2        u0356(.A(men_men_n382_), .B(x5), .Y(men_men_n406_));
  NO2        u0357(.A(x8), .B(x5), .Y(men_men_n407_));
  NAi21      u0358(.An(men_men_n407_), .B(men_men_n162_), .Y(men_men_n408_));
  OAI210     u0359(.A0(men_men_n408_), .A1(men_men_n280_), .B0(men_men_n406_), .Y(men_men_n409_));
  NA2        u0360(.A(men_men_n322_), .B(men_men_n71_), .Y(men_men_n410_));
  NOi21      u0361(.An(x3), .B(x4), .Y(men_men_n411_));
  NA2        u0362(.A(men_men_n55_), .B(men_men_n99_), .Y(men_men_n412_));
  NA2        u0363(.A(men_men_n412_), .B(men_men_n411_), .Y(men_men_n413_));
  NO2        u0364(.A(men_men_n51_), .B(x6), .Y(men_men_n414_));
  NO2        u0365(.A(men_men_n137_), .B(men_men_n55_), .Y(men_men_n415_));
  NO3        u0366(.A(men_men_n56_), .B(x2), .C(x0), .Y(men_men_n416_));
  AOI220     u0367(.A0(men_men_n416_), .A1(men_men_n415_), .B0(men_men_n414_), .B1(men_men_n393_), .Y(men_men_n417_));
  OAI210     u0368(.A0(men_men_n413_), .A1(men_men_n410_), .B0(men_men_n417_), .Y(men_men_n418_));
  AOI210     u0369(.A0(men_men_n409_), .A1(men_men_n405_), .B0(men_men_n418_), .Y(men_men_n419_));
  AOI210     u0370(.A0(men_men_n419_), .A1(men_men_n404_), .B0(men_men_n400_), .Y(men_men_n420_));
  NA2        u0371(.A(x7), .B(x1), .Y(men_men_n421_));
  NO3        u0372(.A(x5), .B(x4), .C(x2), .Y(men_men_n422_));
  AN2        u0373(.A(men_men_n422_), .B(men_men_n328_), .Y(men_men_n423_));
  NO3        u0374(.A(men_men_n423_), .B(men_men_n415_), .C(men_men_n337_), .Y(men_men_n424_));
  INV        u0375(.A(men_men_n309_), .Y(men_men_n425_));
  NO2        u0376(.A(men_men_n425_), .B(men_men_n424_), .Y(men_men_n426_));
  NO2        u0377(.A(x4), .B(men_men_n99_), .Y(men_men_n427_));
  NA2        u0378(.A(men_men_n427_), .B(x6), .Y(men_men_n428_));
  NA3        u0379(.A(men_men_n97_), .B(x4), .C(men_men_n99_), .Y(men_men_n429_));
  AOI210     u0380(.A0(men_men_n429_), .A1(men_men_n428_), .B0(men_men_n89_), .Y(men_men_n430_));
  NA2        u0381(.A(men_men_n411_), .B(men_men_n67_), .Y(men_men_n431_));
  NA2        u0382(.A(men_men_n158_), .B(men_men_n59_), .Y(men_men_n432_));
  NA2        u0383(.A(men_men_n397_), .B(x4), .Y(men_men_n433_));
  INV        u0384(.A(men_men_n433_), .Y(men_men_n434_));
  NO3        u0385(.A(men_men_n434_), .B(men_men_n430_), .C(men_men_n426_), .Y(men_men_n435_));
  NA2        u0386(.A(x5), .B(x4), .Y(men_men_n436_));
  NO2        u0387(.A(men_men_n67_), .B(men_men_n53_), .Y(men_men_n437_));
  NO3        u0388(.A(x8), .B(x3), .C(x2), .Y(men_men_n438_));
  NO3        u0389(.A(x6), .B(x5), .C(x2), .Y(men_men_n439_));
  NA3        u0390(.A(men_men_n439_), .B(men_men_n264_), .C(men_men_n72_), .Y(men_men_n440_));
  INV        u0391(.A(men_men_n440_), .Y(men_men_n441_));
  NA2        u0392(.A(men_men_n67_), .B(x2), .Y(men_men_n442_));
  NO3        u0393(.A(x4), .B(x3), .C(men_men_n59_), .Y(men_men_n443_));
  NA2        u0394(.A(men_men_n443_), .B(men_men_n208_), .Y(men_men_n444_));
  XO2        u0395(.A(x4), .B(x0), .Y(men_men_n445_));
  NA2        u0396(.A(men_men_n241_), .B(x5), .Y(men_men_n446_));
  NO2        u0397(.A(men_men_n56_), .B(men_men_n50_), .Y(men_men_n447_));
  NO2        u0398(.A(men_men_n447_), .B(men_men_n62_), .Y(men_men_n448_));
  NO4        u0399(.A(men_men_n448_), .B(men_men_n446_), .C(men_men_n445_), .D(men_men_n146_), .Y(men_men_n449_));
  NO2        u0400(.A(men_men_n449_), .B(men_men_n441_), .Y(men_men_n450_));
  OAI210     u0401(.A0(men_men_n435_), .A1(men_men_n421_), .B0(men_men_n450_), .Y(men_men_n451_));
  NO4        u0402(.A(men_men_n451_), .B(men_men_n420_), .C(men_men_n399_), .D(men_men_n379_), .Y(men04));
  NO2        u0403(.A(x7), .B(x2), .Y(men_men_n453_));
  NO2        u0404(.A(x3), .B(men_men_n53_), .Y(men_men_n454_));
  NO2        u0405(.A(men_men_n454_), .B(men_men_n139_), .Y(men_men_n455_));
  XN2        u0406(.A(x8), .B(x1), .Y(men_men_n456_));
  NO2        u0407(.A(men_men_n456_), .B(men_men_n137_), .Y(men_men_n457_));
  NA2        u0408(.A(men_men_n457_), .B(men_men_n455_), .Y(men_men_n458_));
  NA2        u0409(.A(x6), .B(x3), .Y(men_men_n459_));
  NO2        u0410(.A(men_men_n459_), .B(x5), .Y(men_men_n460_));
  NA2        u0411(.A(men_men_n67_), .B(x1), .Y(men_men_n461_));
  NO2        u0412(.A(men_men_n407_), .B(men_men_n232_), .Y(men_men_n462_));
  NO3        u0413(.A(men_men_n462_), .B(men_men_n386_), .C(men_men_n461_), .Y(men_men_n463_));
  AOI210     u0414(.A0(men_men_n460_), .A1(men_men_n314_), .B0(men_men_n463_), .Y(men_men_n464_));
  AOI210     u0415(.A0(men_men_n464_), .A1(men_men_n458_), .B0(x0), .Y(men_men_n465_));
  NOi21      u0416(.An(men_men_n162_), .B(men_men_n407_), .Y(men_men_n466_));
  NA2        u0417(.A(men_men_n98_), .B(x1), .Y(men_men_n467_));
  NO3        u0418(.A(men_men_n467_), .B(men_men_n466_), .C(men_men_n295_), .Y(men_men_n468_));
  OAI210     u0419(.A0(men_men_n468_), .A1(men_men_n465_), .B0(men_men_n453_), .Y(men_men_n469_));
  NA2        u0420(.A(men_men_n124_), .B(men_men_n219_), .Y(men_men_n470_));
  OR3        u0421(.A(men_men_n470_), .B(men_men_n329_), .C(men_men_n54_), .Y(men_men_n471_));
  OR2        u0422(.A(x6), .B(x0), .Y(men_men_n472_));
  NO3        u0423(.A(men_men_n472_), .B(x3), .C(x1), .Y(men_men_n473_));
  NO2        u0424(.A(men_men_n471_), .B(men_men_n175_), .Y(men_men_n474_));
  NA2        u0425(.A(x7), .B(x2), .Y(men_men_n475_));
  OAI210     u0426(.A0(men_men_n161_), .A1(x3), .B0(men_men_n74_), .Y(men_men_n476_));
  NO3        u0427(.A(x3), .B(x1), .C(x0), .Y(men_men_n477_));
  OR2        u0428(.A(x6), .B(x1), .Y(men_men_n478_));
  NO2        u0429(.A(men_men_n476_), .B(men_men_n475_), .Y(men_men_n479_));
  NA2        u0430(.A(men_men_n67_), .B(x0), .Y(men_men_n480_));
  NOi31      u0431(.An(men_men_n312_), .B(men_men_n480_), .C(men_men_n237_), .Y(men_men_n481_));
  NO4        u0432(.A(men_men_n481_), .B(men_men_n479_), .C(men_men_n474_), .D(men_men_n56_), .Y(men_men_n482_));
  NA2        u0433(.A(men_men_n482_), .B(men_men_n469_), .Y(men_men_n483_));
  NA3        u0434(.A(x8), .B(x7), .C(x0), .Y(men_men_n484_));
  INV        u0435(.A(men_men_n484_), .Y(men_men_n485_));
  AOI210     u0436(.A0(men_men_n247_), .A1(men_men_n88_), .B0(men_men_n485_), .Y(men_men_n486_));
  NO2        u0437(.A(men_men_n486_), .B(men_men_n146_), .Y(men_men_n487_));
  NA2        u0438(.A(men_men_n382_), .B(men_men_n57_), .Y(men_men_n488_));
  NO2        u0439(.A(x8), .B(x0), .Y(men_men_n489_));
  NO2        u0440(.A(men_men_n488_), .B(men_men_n250_), .Y(men_men_n490_));
  OAI210     u0441(.A0(men_men_n490_), .A1(men_men_n487_), .B0(men_men_n253_), .Y(men_men_n491_));
  NO2        u0442(.A(men_men_n67_), .B(men_men_n99_), .Y(men_men_n492_));
  NO2        u0443(.A(men_men_n327_), .B(x8), .Y(men_men_n493_));
  NO2        u0444(.A(men_men_n493_), .B(men_men_n238_), .Y(men_men_n494_));
  NO2        u0445(.A(men_men_n494_), .B(men_men_n333_), .Y(men_men_n495_));
  NO2        u0446(.A(men_men_n261_), .B(x8), .Y(men_men_n496_));
  OAI210     u0447(.A0(men_men_n407_), .A1(men_men_n296_), .B0(men_men_n221_), .Y(men_men_n497_));
  NA2        u0448(.A(men_men_n314_), .B(men_men_n167_), .Y(men_men_n498_));
  OAI220     u0449(.A0(men_men_n498_), .A1(men_men_n59_), .B0(men_men_n497_), .B1(men_men_n496_), .Y(men_men_n499_));
  OAI210     u0450(.A0(men_men_n499_), .A1(men_men_n495_), .B0(men_men_n492_), .Y(men_men_n500_));
  NO2        u0451(.A(x8), .B(x2), .Y(men_men_n501_));
  NO2        u0452(.A(men_men_n203_), .B(men_men_n57_), .Y(men_men_n502_));
  NA3        u0453(.A(men_men_n502_), .B(men_men_n501_), .C(men_men_n310_), .Y(men_men_n503_));
  NO2        u0454(.A(men_men_n222_), .B(men_men_n124_), .Y(men_men_n504_));
  INV        u0455(.A(men_men_n504_), .Y(men_men_n505_));
  AOI210     u0456(.A0(men_men_n505_), .A1(men_men_n503_), .B0(men_men_n98_), .Y(men_men_n506_));
  NA2        u0457(.A(men_men_n308_), .B(x2), .Y(men_men_n507_));
  NO2        u0458(.A(men_men_n57_), .B(men_men_n53_), .Y(men_men_n508_));
  NA2        u0459(.A(men_men_n99_), .B(men_men_n53_), .Y(men_men_n509_));
  NO2        u0460(.A(men_men_n509_), .B(x8), .Y(men_men_n510_));
  NA2        u0461(.A(x7), .B(men_men_n50_), .Y(men_men_n511_));
  NO2        u0462(.A(men_men_n172_), .B(men_men_n511_), .Y(men_men_n512_));
  AN2        u0463(.A(men_men_n512_), .B(men_men_n510_), .Y(men_men_n513_));
  NA2        u0464(.A(men_men_n356_), .B(men_men_n139_), .Y(men_men_n514_));
  NO2        u0465(.A(men_men_n67_), .B(x2), .Y(men_men_n515_));
  NA2        u0466(.A(men_men_n515_), .B(men_men_n247_), .Y(men_men_n516_));
  NO3        u0467(.A(x4), .B(men_men_n513_), .C(men_men_n506_), .Y(men_men_n517_));
  NA3        u0468(.A(men_men_n517_), .B(men_men_n500_), .C(men_men_n491_), .Y(men_men_n518_));
  NA2        u0469(.A(men_men_n53_), .B(men_men_n59_), .Y(men_men_n519_));
  NOi21      u0470(.An(x2), .B(x7), .Y(men_men_n520_));
  NO2        u0471(.A(x6), .B(x3), .Y(men_men_n521_));
  NA2        u0472(.A(men_men_n521_), .B(men_men_n520_), .Y(men_men_n522_));
  NO2        u0473(.A(x6), .B(men_men_n59_), .Y(men_men_n523_));
  NO3        u0474(.A(men_men_n57_), .B(x2), .C(x1), .Y(men_men_n524_));
  NO3        u0475(.A(men_men_n57_), .B(x2), .C(x0), .Y(men_men_n525_));
  AOI220     u0476(.A0(men_men_n525_), .A1(men_men_n205_), .B0(men_men_n524_), .B1(men_men_n523_), .Y(men_men_n526_));
  NA2        u0477(.A(men_men_n522_), .B(men_men_n526_), .Y(men_men_n527_));
  NO2        u0478(.A(men_men_n90_), .B(men_men_n53_), .Y(men_men_n528_));
  NA2        u0479(.A(men_men_n201_), .B(men_men_n57_), .Y(men_men_n529_));
  NA2        u0480(.A(men_men_n528_), .B(men_men_n529_), .Y(men_men_n530_));
  NO3        u0481(.A(men_men_n530_), .B(men_men_n433_), .C(men_men_n59_), .Y(men_men_n531_));
  AO210      u0482(.A0(men_men_n527_), .A1(men_men_n407_), .B0(men_men_n531_), .Y(men_men_n532_));
  AOI210     u0483(.A0(men_men_n518_), .A1(men_men_n483_), .B0(men_men_n532_), .Y(men05));
  AOI210     u0484(.A0(men_men_n153_), .A1(men_men_n55_), .B0(men_men_n447_), .Y(men_men_n534_));
  OR2        u0485(.A(men_men_n534_), .B(men_men_n57_), .Y(men_men_n535_));
  NO2        u0486(.A(x7), .B(men_men_n97_), .Y(men_men_n536_));
  NO2        u0487(.A(x8), .B(men_men_n56_), .Y(men_men_n537_));
  NA2        u0488(.A(x5), .B(men_men_n56_), .Y(men_men_n538_));
  NO2        u0489(.A(men_men_n538_), .B(men_men_n511_), .Y(men_men_n539_));
  NO2        u0490(.A(men_men_n535_), .B(men_men_n99_), .Y(men_men_n540_));
  NO2        u0491(.A(x7), .B(x4), .Y(men_men_n541_));
  NO2        u0492(.A(men_men_n63_), .B(men_men_n55_), .Y(men_men_n542_));
  NO2        u0493(.A(men_men_n185_), .B(x5), .Y(men_men_n543_));
  NA2        u0494(.A(men_men_n97_), .B(men_men_n99_), .Y(men_men_n544_));
  NO2        u0495(.A(men_men_n544_), .B(men_men_n199_), .Y(men_men_n545_));
  AO220      u0496(.A0(men_men_n545_), .A1(men_men_n541_), .B0(men_men_n543_), .B1(men_men_n542_), .Y(men_men_n546_));
  OAI210     u0497(.A0(men_men_n546_), .A1(men_men_n540_), .B0(men_men_n437_), .Y(men_men_n547_));
  NO2        u0498(.A(x6), .B(men_men_n50_), .Y(men_men_n548_));
  NA2        u0499(.A(men_men_n55_), .B(x4), .Y(men_men_n549_));
  NO2        u0500(.A(men_men_n97_), .B(men_men_n99_), .Y(men_men_n550_));
  NA2        u0501(.A(men_men_n385_), .B(men_men_n231_), .Y(men_men_n551_));
  NA2        u0502(.A(men_men_n97_), .B(x4), .Y(men_men_n552_));
  NA3        u0503(.A(x1), .B(men_men_n552_), .C(men_men_n297_), .Y(men_men_n553_));
  NO2        u0504(.A(men_men_n97_), .B(x2), .Y(men_men_n554_));
  NO2        u0505(.A(men_men_n69_), .B(men_men_n55_), .Y(men_men_n555_));
  NA2        u0506(.A(men_men_n555_), .B(men_men_n554_), .Y(men_men_n556_));
  NA2        u0507(.A(men_men_n556_), .B(men_men_n553_), .Y(men_men_n557_));
  NA2        u0508(.A(men_men_n557_), .B(men_men_n548_), .Y(men_men_n558_));
  NO2        u0509(.A(men_men_n67_), .B(men_men_n50_), .Y(men_men_n559_));
  NO2        u0510(.A(men_men_n181_), .B(x4), .Y(men_men_n560_));
  NO2        u0511(.A(x5), .B(men_men_n56_), .Y(men_men_n561_));
  XO2        u0512(.A(x5), .B(x2), .Y(men_men_n562_));
  NO3        u0513(.A(x8), .B(x7), .C(men_men_n99_), .Y(men_men_n563_));
  AN2        u0514(.A(men_men_n562_), .B(men_men_n560_), .Y(men_men_n564_));
  NA3        u0515(.A(men_men_n564_), .B(men_men_n559_), .C(men_men_n53_), .Y(men_men_n565_));
  NA2        u0516(.A(men_men_n244_), .B(men_men_n520_), .Y(men_men_n566_));
  NOi21      u0517(.An(x4), .B(x1), .Y(men_men_n567_));
  NA2        u0518(.A(men_men_n567_), .B(men_men_n62_), .Y(men_men_n568_));
  NA2        u0519(.A(x4), .B(x1), .Y(men_men_n569_));
  NO2        u0520(.A(men_men_n569_), .B(men_men_n50_), .Y(men_men_n570_));
  AOI210     u0521(.A0(men_men_n570_), .A1(men_men_n550_), .B0(men_men_n59_), .Y(men_men_n571_));
  BUFFER     u0522(.A(men_men_n571_), .Y(men_men_n572_));
  NA4        u0523(.A(men_men_n572_), .B(men_men_n565_), .C(men_men_n558_), .D(men_men_n547_), .Y(men_men_n573_));
  NA2        u0524(.A(men_men_n559_), .B(men_men_n56_), .Y(men_men_n574_));
  NA2        u0525(.A(men_men_n501_), .B(men_men_n536_), .Y(men_men_n575_));
  NO2        u0526(.A(men_men_n575_), .B(men_men_n574_), .Y(men_men_n576_));
  NA2        u0527(.A(men_men_n247_), .B(men_men_n111_), .Y(men_men_n577_));
  OAI210     u0528(.A0(men_men_n577_), .A1(men_men_n155_), .B0(men_men_n59_), .Y(men_men_n578_));
  NA2        u0529(.A(men_men_n57_), .B(x6), .Y(men_men_n579_));
  NA2        u0530(.A(men_men_n561_), .B(men_men_n145_), .Y(men_men_n580_));
  NO3        u0531(.A(men_men_n580_), .B(men_men_n57_), .C(men_men_n375_), .Y(men_men_n581_));
  NA2        u0532(.A(men_men_n254_), .B(men_men_n67_), .Y(men_men_n582_));
  NO2        u0533(.A(men_men_n411_), .B(men_men_n97_), .Y(men_men_n583_));
  NO2        u0534(.A(men_men_n509_), .B(x6), .Y(men_men_n584_));
  NO3        u0535(.A(men_men_n581_), .B(men_men_n578_), .C(men_men_n576_), .Y(men_men_n585_));
  NA2        u0536(.A(men_men_n57_), .B(x5), .Y(men_men_n586_));
  NO2        u0537(.A(men_men_n586_), .B(x1), .Y(men_men_n587_));
  NA2        u0538(.A(x8), .B(men_men_n56_), .Y(men_men_n588_));
  NO2        u0539(.A(men_men_n588_), .B(men_men_n119_), .Y(men_men_n589_));
  NA2        u0540(.A(x8), .B(x4), .Y(men_men_n590_));
  NO2        u0541(.A(x8), .B(x4), .Y(men_men_n591_));
  NAi21      u0542(.An(men_men_n591_), .B(men_men_n590_), .Y(men_men_n592_));
  NAi21      u0543(.An(men_men_n501_), .B(men_men_n340_), .Y(men_men_n593_));
  NO4        u0544(.A(men_men_n593_), .B(men_men_n592_), .C(men_men_n375_), .D(men_men_n67_), .Y(men_men_n594_));
  OAI210     u0545(.A0(men_men_n594_), .A1(men_men_n589_), .B0(men_men_n587_), .Y(men_men_n595_));
  NO3        u0546(.A(x8), .B(men_men_n97_), .C(x4), .Y(men_men_n596_));
  INV        u0547(.A(men_men_n596_), .Y(men_men_n597_));
  NO2        u0548(.A(men_men_n597_), .B(men_men_n99_), .Y(men_men_n598_));
  NO2        u0549(.A(x5), .B(x4), .Y(men_men_n599_));
  NA3        u0550(.A(men_men_n599_), .B(men_men_n62_), .C(men_men_n99_), .Y(men_men_n600_));
  NO2        u0551(.A(x6), .B(men_men_n99_), .Y(men_men_n601_));
  INV        u0552(.A(men_men_n600_), .Y(men_men_n602_));
  OAI210     u0553(.A0(men_men_n602_), .A1(men_men_n598_), .B0(men_men_n283_), .Y(men_men_n603_));
  NA3        u0554(.A(men_men_n603_), .B(men_men_n595_), .C(men_men_n585_), .Y(men_men_n604_));
  OR2        u0555(.A(x4), .B(x1), .Y(men_men_n605_));
  NO2        u0556(.A(men_men_n605_), .B(x3), .Y(men_men_n606_));
  NA2        u0557(.A(men_men_n55_), .B(x2), .Y(men_men_n607_));
  NA2        u0558(.A(men_men_n604_), .B(men_men_n573_), .Y(men06));
  NA2        u0559(.A(men_men_n56_), .B(x3), .Y(men_men_n609_));
  NA2        u0560(.A(x6), .B(men_men_n99_), .Y(men_men_n610_));
  NA2        u0561(.A(men_men_n610_), .B(men_men_n55_), .Y(men_men_n611_));
  NA2        u0562(.A(x5), .B(men_men_n59_), .Y(men_men_n612_));
  NO2        u0563(.A(men_men_n612_), .B(men_men_n106_), .Y(men_men_n613_));
  NA3        u0564(.A(men_men_n613_), .B(men_men_n611_), .C(men_men_n442_), .Y(men_men_n614_));
  NO2        u0565(.A(men_men_n340_), .B(x0), .Y(men_men_n615_));
  NA2        u0566(.A(men_men_n307_), .B(x2), .Y(men_men_n616_));
  NOi21      u0567(.An(x6), .B(x8), .Y(men_men_n617_));
  NO2        u0568(.A(men_men_n617_), .B(x2), .Y(men_men_n618_));
  NO3        u0569(.A(men_men_n618_), .B(men_men_n66_), .C(men_men_n59_), .Y(men_men_n619_));
  AOI220     u0570(.A0(men_men_n619_), .A1(men_men_n616_), .B0(men_men_n615_), .B1(men_men_n299_), .Y(men_men_n620_));
  AOI210     u0571(.A0(men_men_n620_), .A1(men_men_n614_), .B0(men_men_n609_), .Y(men_men_n621_));
  NA2        u0572(.A(men_men_n56_), .B(men_men_n50_), .Y(men_men_n622_));
  NA2        u0573(.A(men_men_n326_), .B(men_men_n317_), .Y(men_men_n623_));
  NO2        u0574(.A(men_men_n67_), .B(men_men_n97_), .Y(men_men_n624_));
  NO2        u0575(.A(men_men_n53_), .B(men_men_n59_), .Y(men_men_n625_));
  NO3        u0576(.A(men_men_n607_), .B(men_men_n624_), .C(men_men_n437_), .Y(men_men_n626_));
  AOI220     u0577(.A0(men_men_n626_), .A1(men_men_n623_), .B0(men_men_n372_), .B1(men_men_n62_), .Y(men_men_n627_));
  NO2        u0578(.A(men_men_n627_), .B(men_men_n622_), .Y(men_men_n628_));
  NO2        u0579(.A(men_men_n54_), .B(x0), .Y(men_men_n629_));
  NA2        u0580(.A(x4), .B(x3), .Y(men_men_n630_));
  NA2        u0581(.A(x3), .B(men_men_n629_), .Y(men_men_n631_));
  NO2        u0582(.A(men_men_n93_), .B(men_men_n56_), .Y(men_men_n632_));
  NA2        u0583(.A(men_men_n632_), .B(men_men_n232_), .Y(men_men_n633_));
  AOI210     u0584(.A0(men_men_n633_), .A1(men_men_n631_), .B0(x2), .Y(men_men_n634_));
  INV        u0585(.A(men_men_n337_), .Y(men_men_n635_));
  NO2        u0586(.A(men_men_n359_), .B(x8), .Y(men_men_n636_));
  NO2        u0587(.A(men_men_n233_), .B(men_men_n461_), .Y(men_men_n637_));
  AOI210     u0588(.A0(men_men_n636_), .A1(men_men_n239_), .B0(men_men_n637_), .Y(men_men_n638_));
  NO2        u0589(.A(x5), .B(x3), .Y(men_men_n639_));
  NA3        u0590(.A(men_men_n489_), .B(men_men_n639_), .C(x1), .Y(men_men_n640_));
  NA2        u0591(.A(men_men_n537_), .B(men_men_n492_), .Y(men_men_n641_));
  OA220      u0592(.A0(men_men_n641_), .A1(men_men_n514_), .B0(men_men_n640_), .B1(men_men_n442_), .Y(men_men_n642_));
  OAI210     u0593(.A0(men_men_n638_), .A1(men_men_n635_), .B0(men_men_n642_), .Y(men_men_n643_));
  OR4        u0594(.A(men_men_n643_), .B(men_men_n634_), .C(men_men_n628_), .D(men_men_n621_), .Y(men_men_n644_));
  NA2        u0595(.A(x7), .B(men_men_n56_), .Y(men_men_n645_));
  NO2        u0596(.A(men_men_n550_), .B(men_men_n59_), .Y(men_men_n646_));
  NA2        u0597(.A(men_men_n646_), .B(men_men_n559_), .Y(men_men_n647_));
  NO2        u0598(.A(men_men_n160_), .B(x6), .Y(men_men_n648_));
  NO2        u0599(.A(men_men_n647_), .B(men_men_n645_), .Y(men_men_n649_));
  AN2        u0600(.A(men_men_n416_), .B(men_men_n294_), .Y(men_men_n650_));
  OAI210     u0601(.A0(men_men_n650_), .A1(men_men_n649_), .B0(men_men_n314_), .Y(men_men_n651_));
  NO2        u0602(.A(men_men_n279_), .B(men_men_n97_), .Y(men_men_n652_));
  NO2        u0603(.A(men_men_n56_), .B(x3), .Y(men_men_n653_));
  NA2        u0604(.A(men_men_n653_), .B(men_men_n67_), .Y(men_men_n654_));
  NO2        u0605(.A(men_men_n67_), .B(x3), .Y(men_men_n655_));
  NO2        u0606(.A(men_men_n57_), .B(x6), .Y(men_men_n656_));
  NA2        u0607(.A(men_men_n171_), .B(men_men_n656_), .Y(men_men_n657_));
  INV        u0608(.A(men_men_n657_), .Y(men_men_n658_));
  OR2        u0609(.A(men_men_n658_), .B(men_men_n570_), .Y(men_men_n659_));
  NA2        u0610(.A(men_men_n659_), .B(men_men_n652_), .Y(men_men_n660_));
  NA2        u0611(.A(x7), .B(x6), .Y(men_men_n661_));
  NA3        u0612(.A(x2), .B(x1), .C(x0), .Y(men_men_n662_));
  NO3        u0613(.A(men_men_n662_), .B(men_men_n661_), .C(men_men_n534_), .Y(men_men_n663_));
  NA2        u0614(.A(men_men_n438_), .B(men_men_n138_), .Y(men_men_n664_));
  NO2        u0615(.A(x5), .B(x1), .Y(men_men_n665_));
  NA2        u0616(.A(men_men_n665_), .B(men_men_n656_), .Y(men_men_n666_));
  NA2        u0617(.A(x4), .B(x0), .Y(men_men_n667_));
  NO3        u0618(.A(men_men_n57_), .B(x6), .C(x2), .Y(men_men_n668_));
  NA2        u0619(.A(men_men_n668_), .B(men_men_n204_), .Y(men_men_n669_));
  OAI220     u0620(.A0(men_men_n669_), .A1(men_men_n667_), .B0(men_men_n666_), .B1(men_men_n664_), .Y(men_men_n670_));
  NO2        u0621(.A(men_men_n670_), .B(men_men_n663_), .Y(men_men_n671_));
  NA3        u0622(.A(men_men_n671_), .B(men_men_n660_), .C(men_men_n651_), .Y(men_men_n672_));
  AOI210     u0623(.A0(men_men_n644_), .A1(men_men_n57_), .B0(men_men_n672_), .Y(men07));
  NA2        u0624(.A(men_men_n97_), .B(men_men_n59_), .Y(men_men_n674_));
  NOi21      u0625(.An(men_men_n661_), .B(men_men_n105_), .Y(men_men_n675_));
  NO3        u0626(.A(men_men_n675_), .B(men_men_n227_), .C(men_men_n674_), .Y(men_men_n676_));
  NO3        u0627(.A(men_men_n57_), .B(x5), .C(x1), .Y(men_men_n677_));
  NO2        u0628(.A(men_men_n57_), .B(men_men_n67_), .Y(men_men_n678_));
  NO2        u0629(.A(men_men_n144_), .B(men_men_n98_), .Y(men_men_n679_));
  INV        u0630(.A(men_men_n679_), .Y(men_men_n680_));
  NO2        u0631(.A(men_men_n680_), .B(men_men_n124_), .Y(men_men_n681_));
  OAI210     u0632(.A0(men_men_n681_), .A1(men_men_n676_), .B0(x2), .Y(men_men_n682_));
  NAi21      u0633(.An(men_men_n145_), .B(men_men_n146_), .Y(men_men_n683_));
  NO3        u0634(.A(men_men_n55_), .B(x3), .C(x1), .Y(men_men_n684_));
  NO2        u0635(.A(men_men_n454_), .B(x2), .Y(men_men_n685_));
  AOI210     u0636(.A0(men_men_n685_), .A1(men_men_n456_), .B0(men_men_n684_), .Y(men_men_n686_));
  NO2        u0637(.A(men_men_n686_), .B(men_men_n579_), .Y(men_men_n687_));
  NO2        u0638(.A(x8), .B(men_men_n53_), .Y(men_men_n688_));
  NA2        u0639(.A(men_men_n688_), .B(men_men_n59_), .Y(men_men_n689_));
  NA2        u0640(.A(men_men_n318_), .B(men_men_n314_), .Y(men_men_n690_));
  NO2        u0641(.A(x7), .B(x3), .Y(men_men_n691_));
  NA2        u0642(.A(men_men_n691_), .B(men_men_n90_), .Y(men_men_n692_));
  AOI210     u0643(.A0(men_men_n690_), .A1(men_men_n689_), .B0(men_men_n692_), .Y(men_men_n693_));
  AOI210     u0644(.A0(men_men_n687_), .A1(men_men_n226_), .B0(men_men_n693_), .Y(men_men_n694_));
  AOI210     u0645(.A0(men_men_n694_), .A1(men_men_n682_), .B0(x4), .Y(men_men_n695_));
  NO2        u0646(.A(men_men_n530_), .B(men_men_n99_), .Y(men_men_n696_));
  XO2        u0647(.A(x5), .B(x1), .Y(men_men_n697_));
  NO3        u0648(.A(men_men_n697_), .B(men_men_n193_), .C(men_men_n55_), .Y(men_men_n698_));
  OAI210     u0649(.A0(men_men_n698_), .A1(men_men_n696_), .B0(men_men_n363_), .Y(men_men_n699_));
  NO3        u0650(.A(men_men_n50_), .B(x2), .C(x0), .Y(men_men_n700_));
  NA2        u0651(.A(x6), .B(x0), .Y(men_men_n701_));
  NO2        u0652(.A(men_men_n607_), .B(men_men_n701_), .Y(men_men_n702_));
  NO2        u0653(.A(men_men_n697_), .B(men_men_n617_), .Y(men_men_n703_));
  OAI210     u0654(.A0(men_men_n665_), .A1(men_men_n62_), .B0(men_men_n57_), .Y(men_men_n704_));
  NO2        u0655(.A(men_men_n704_), .B(men_men_n703_), .Y(men_men_n705_));
  NA2        u0656(.A(men_men_n705_), .B(men_men_n700_), .Y(men_men_n706_));
  AOI210     u0657(.A0(men_men_n706_), .A1(men_men_n699_), .B0(men_men_n56_), .Y(men_men_n707_));
  NOi21      u0658(.An(men_men_n211_), .B(men_men_n328_), .Y(men_men_n708_));
  NO3        u0659(.A(men_men_n708_), .B(men_men_n218_), .C(men_men_n64_), .Y(men_men_n709_));
  NO2        u0660(.A(men_men_n179_), .B(men_men_n67_), .Y(men_men_n710_));
  NO2        u0661(.A(men_men_n282_), .B(x6), .Y(men_men_n711_));
  AN2        u0662(.A(men_men_n710_), .B(men_men_n493_), .Y(men_men_n712_));
  OAI210     u0663(.A0(men_men_n712_), .A1(men_men_n709_), .B0(men_men_n59_), .Y(men_men_n713_));
  NAi21      u0664(.An(x8), .B(x7), .Y(men_men_n714_));
  NA2        u0665(.A(men_men_n708_), .B(men_men_n714_), .Y(men_men_n715_));
  NA2        u0666(.A(men_men_n356_), .B(men_men_n99_), .Y(men_men_n716_));
  NO2        u0667(.A(men_men_n617_), .B(x1), .Y(men_men_n717_));
  NO3        u0668(.A(men_men_n717_), .B(men_men_n716_), .C(men_men_n508_), .Y(men_men_n718_));
  NA2        u0669(.A(men_men_n718_), .B(men_men_n715_), .Y(men_men_n719_));
  AOI210     u0670(.A0(men_men_n719_), .A1(men_men_n713_), .B0(men_men_n131_), .Y(men_men_n720_));
  NO2        u0671(.A(x8), .B(x7), .Y(men_men_n721_));
  NO2        u0672(.A(x8), .B(men_men_n99_), .Y(men_men_n722_));
  AOI220     u0673(.A0(men_men_n296_), .A1(men_men_n314_), .B0(men_men_n722_), .B1(men_men_n231_), .Y(men_men_n723_));
  NO2        u0674(.A(men_men_n67_), .B(x4), .Y(men_men_n724_));
  NA2        u0675(.A(men_men_n724_), .B(men_men_n276_), .Y(men_men_n725_));
  NO2        u0676(.A(men_men_n723_), .B(men_men_n725_), .Y(men_men_n726_));
  NO4        u0677(.A(men_men_n726_), .B(men_men_n720_), .C(men_men_n707_), .D(men_men_n695_), .Y(men08));
  NA2        u0678(.A(men_men_n50_), .B(x1), .Y(men_men_n728_));
  XN2        u0679(.A(x5), .B(x4), .Y(men_men_n729_));
  INV        u0680(.A(men_men_n729_), .Y(men_men_n730_));
  AOI220     u0681(.A0(men_men_n730_), .A1(men_men_n318_), .B0(men_men_n127_), .B1(men_men_n56_), .Y(men_men_n731_));
  NO2        u0682(.A(men_men_n219_), .B(men_men_n97_), .Y(men_men_n732_));
  AOI210     u0683(.A0(men_men_n732_), .A1(men_men_n252_), .B0(men_men_n180_), .Y(men_men_n733_));
  OAI220     u0684(.A0(men_men_n733_), .A1(x4), .B0(men_men_n731_), .B1(men_men_n728_), .Y(men_men_n734_));
  NA2        u0685(.A(men_men_n734_), .B(men_men_n247_), .Y(men_men_n735_));
  AOI210     u0686(.A0(men_men_n246_), .A1(men_men_n716_), .B0(men_men_n549_), .Y(men_men_n736_));
  NA2        u0687(.A(men_men_n544_), .B(men_men_n160_), .Y(men_men_n737_));
  OAI220     u0688(.A0(men_men_n737_), .A1(men_men_n588_), .B0(men_men_n429_), .B1(men_men_n50_), .Y(men_men_n738_));
  AO210      u0689(.A0(men_men_n738_), .A1(men_men_n310_), .B0(men_men_n736_), .Y(men_men_n739_));
  NA2        u0690(.A(men_men_n131_), .B(x7), .Y(men_men_n740_));
  OR3        u0691(.A(men_men_n662_), .B(men_men_n411_), .C(men_men_n639_), .Y(men_men_n741_));
  NO2        u0692(.A(men_men_n741_), .B(men_men_n740_), .Y(men_men_n742_));
  AOI210     u0693(.A0(men_men_n739_), .A1(men_men_n264_), .B0(men_men_n742_), .Y(men_men_n743_));
  AOI210     u0694(.A0(men_men_n743_), .A1(men_men_n735_), .B0(men_men_n67_), .Y(men_men_n744_));
  NO2        u0695(.A(men_men_n721_), .B(men_men_n99_), .Y(men_men_n745_));
  NA2        u0696(.A(men_men_n301_), .B(men_men_n53_), .Y(men_men_n746_));
  NO3        u0697(.A(men_men_n359_), .B(men_men_n124_), .C(men_men_n65_), .Y(men_men_n747_));
  NO2        u0698(.A(men_men_n625_), .B(men_men_n221_), .Y(men_men_n748_));
  NO3        u0699(.A(men_men_n502_), .B(men_men_n412_), .C(men_men_n88_), .Y(men_men_n749_));
  AO220      u0700(.A0(men_men_n749_), .A1(men_men_n748_), .B0(men_men_n747_), .B1(men_men_n746_), .Y(men_men_n750_));
  NA2        u0701(.A(x7), .B(men_men_n59_), .Y(men_men_n751_));
  NO2        u0702(.A(men_men_n285_), .B(men_men_n751_), .Y(men_men_n752_));
  AOI210     u0703(.A0(men_men_n750_), .A1(x5), .B0(men_men_n752_), .Y(men_men_n753_));
  NO2        u0704(.A(men_men_n753_), .B(men_men_n68_), .Y(men_men_n754_));
  NO2        u0705(.A(men_men_n66_), .B(x3), .Y(men_men_n755_));
  OAI210     u0706(.A0(men_men_n755_), .A1(men_men_n238_), .B0(men_men_n136_), .Y(men_men_n756_));
  MUX2       u0707(.S(x3), .A(men_men_n154_), .B(men_men_n683_), .Y(men_men_n757_));
  NO3        u0708(.A(x6), .B(x4), .C(x0), .Y(men_men_n758_));
  INV        u0709(.A(men_men_n758_), .Y(men_men_n759_));
  NO2        u0710(.A(men_men_n756_), .B(men_men_n759_), .Y(men_men_n760_));
  NA2        u0711(.A(men_men_n730_), .B(men_men_n281_), .Y(men_men_n761_));
  OR2        u0712(.A(x8), .B(x1), .Y(men_men_n762_));
  NO2        u0713(.A(men_men_n762_), .B(men_men_n761_), .Y(men_men_n763_));
  NAi21      u0714(.An(x4), .B(x1), .Y(men_men_n764_));
  NO2        u0715(.A(men_men_n764_), .B(x0), .Y(men_men_n765_));
  NA3        u0716(.A(men_men_n55_), .B(x1), .C(x0), .Y(men_men_n766_));
  NA2        u0717(.A(men_men_n763_), .B(men_men_n292_), .Y(men_men_n767_));
  AO210      u0718(.A0(men_men_n262_), .A1(men_men_n238_), .B0(men_men_n652_), .Y(men_men_n768_));
  NA2        u0719(.A(men_men_n97_), .B(men_men_n56_), .Y(men_men_n769_));
  NO2        u0720(.A(men_men_n769_), .B(men_men_n236_), .Y(men_men_n770_));
  NO2        u0721(.A(men_men_n57_), .B(x2), .Y(men_men_n771_));
  NO3        u0722(.A(men_men_n297_), .B(men_men_n771_), .C(men_men_n266_), .Y(men_men_n772_));
  AOI220     u0723(.A0(men_men_n772_), .A1(men_men_n770_), .B0(men_men_n768_), .B1(men_men_n570_), .Y(men_men_n773_));
  NA2        u0724(.A(men_men_n773_), .B(men_men_n767_), .Y(men_men_n774_));
  NO4        u0725(.A(men_men_n774_), .B(men_men_n760_), .C(men_men_n754_), .D(men_men_n744_), .Y(men09));
  NO2        u0726(.A(men_men_n519_), .B(men_men_n237_), .Y(men_men_n776_));
  NO2        u0727(.A(men_men_n665_), .B(men_men_n307_), .Y(men_men_n777_));
  NO2        u0728(.A(men_men_n91_), .B(men_men_n99_), .Y(men_men_n778_));
  AO220      u0729(.A0(men_men_n778_), .A1(men_men_n777_), .B0(men_men_n776_), .B1(men_men_n550_), .Y(men_men_n779_));
  NA2        u0730(.A(men_men_n779_), .B(x4), .Y(men_men_n780_));
  OAI220     u0731(.A0(men_men_n326_), .A1(men_men_n133_), .B0(men_men_n347_), .B1(men_men_n253_), .Y(men_men_n781_));
  NO2        u0732(.A(men_men_n179_), .B(men_men_n97_), .Y(men_men_n782_));
  AOI220     u0733(.A0(men_men_n782_), .A1(men_men_n113_), .B0(men_men_n781_), .B1(x1), .Y(men_men_n783_));
  NAi21      u0734(.An(x0), .B(x2), .Y(men_men_n784_));
  NO2        u0735(.A(men_men_n275_), .B(men_men_n784_), .Y(men_men_n785_));
  OAI210     u0736(.A0(men_men_n421_), .A1(men_men_n249_), .B0(men_men_n179_), .Y(men_men_n786_));
  AOI210     u0737(.A0(men_men_n157_), .A1(men_men_n714_), .B0(men_men_n317_), .Y(men_men_n787_));
  NA2        u0738(.A(men_men_n787_), .B(men_men_n786_), .Y(men_men_n788_));
  OAI210     u0739(.A0(men_men_n783_), .A1(men_men_n55_), .B0(men_men_n788_), .Y(men_men_n789_));
  NA2        u0740(.A(men_men_n789_), .B(men_men_n56_), .Y(men_men_n790_));
  NO2        u0741(.A(men_men_n56_), .B(men_men_n59_), .Y(men_men_n791_));
  INV        u0742(.A(men_men_n113_), .Y(men_men_n792_));
  NA2        u0743(.A(men_men_n665_), .B(men_men_n55_), .Y(men_men_n793_));
  NA2        u0744(.A(men_men_n492_), .B(men_men_n55_), .Y(men_men_n794_));
  NO2        u0745(.A(men_men_n210_), .B(men_men_n338_), .Y(men_men_n795_));
  NO2        u0746(.A(men_men_n282_), .B(men_men_n137_), .Y(men_men_n796_));
  OAI220     u0747(.A0(x1), .A1(men_men_n55_), .B0(men_men_n794_), .B1(men_men_n400_), .Y(men_men_n797_));
  NA2        u0748(.A(men_men_n797_), .B(men_men_n791_), .Y(men_men_n798_));
  NO2        u0749(.A(men_men_n354_), .B(men_men_n97_), .Y(men_men_n799_));
  NA2        u0750(.A(men_men_n57_), .B(men_men_n799_), .Y(men_men_n800_));
  NA4        u0751(.A(men_men_n800_), .B(men_men_n798_), .C(men_men_n790_), .D(men_men_n780_), .Y(men_men_n801_));
  NA2        u0752(.A(men_men_n801_), .B(men_men_n50_), .Y(men_men_n802_));
  NO2        u0753(.A(men_men_n331_), .B(men_men_n150_), .Y(men_men_n803_));
  NO3        u0754(.A(men_men_n57_), .B(x5), .C(x2), .Y(men_men_n804_));
  NO2        u0755(.A(men_men_n373_), .B(men_men_n136_), .Y(men_men_n805_));
  NO2        u0756(.A(men_men_n52_), .B(x2), .Y(men_men_n806_));
  NO2        u0757(.A(men_men_n97_), .B(men_men_n56_), .Y(men_men_n807_));
  NA2        u0758(.A(men_men_n807_), .B(x8), .Y(men_men_n808_));
  NA2        u0759(.A(men_men_n808_), .B(men_men_n793_), .Y(men_men_n809_));
  AO210      u0760(.A0(men_men_n809_), .A1(men_men_n806_), .B0(men_men_n805_), .Y(men_men_n810_));
  NA2        u0761(.A(men_men_n810_), .B(men_men_n548_), .Y(men_men_n811_));
  OAI210     u0762(.A0(x4), .A1(x2), .B0(x0), .Y(men_men_n812_));
  NA3        u0763(.A(men_men_n538_), .B(men_men_n549_), .C(men_men_n311_), .Y(men_men_n813_));
  OAI210     u0764(.A0(men_men_n812_), .A1(men_men_n259_), .B0(men_men_n53_), .Y(men_men_n814_));
  AOI210     u0765(.A0(men_men_n813_), .A1(men_men_n812_), .B0(men_men_n814_), .Y(men_men_n815_));
  NA2        u0766(.A(men_men_n815_), .B(men_men_n296_), .Y(men_men_n816_));
  AOI220     u0767(.A0(men_men_n590_), .A1(men_men_n313_), .B0(men_men_n314_), .B1(men_men_n84_), .Y(men_men_n817_));
  NA2        u0768(.A(men_men_n84_), .B(x5), .Y(men_men_n818_));
  OAI220     u0769(.A0(men_men_n818_), .A1(men_men_n762_), .B0(men_men_n817_), .B1(men_men_n293_), .Y(men_men_n819_));
  NA2        u0770(.A(men_men_n819_), .B(men_men_n65_), .Y(men_men_n820_));
  NA2        u0771(.A(men_men_n356_), .B(men_men_n683_), .Y(men_men_n821_));
  NA2        u0772(.A(men_men_n226_), .B(men_men_n154_), .Y(men_men_n822_));
  AO210      u0773(.A0(men_men_n822_), .A1(men_men_n821_), .B0(men_men_n121_), .Y(men_men_n823_));
  NO2        u0774(.A(men_men_n386_), .B(x2), .Y(men_men_n824_));
  NO2        u0775(.A(x7), .B(men_men_n53_), .Y(men_men_n825_));
  NA2        u0776(.A(men_men_n825_), .B(x5), .Y(men_men_n826_));
  NO2        u0777(.A(men_men_n826_), .B(men_men_n60_), .Y(men_men_n827_));
  AOI220     u0778(.A0(men_men_n827_), .A1(men_men_n824_), .B0(men_men_n591_), .B1(men_men_n220_), .Y(men_men_n828_));
  NA4        u0779(.A(men_men_n828_), .B(men_men_n823_), .C(men_men_n820_), .D(men_men_n816_), .Y(men_men_n829_));
  NO4        u0780(.A(men_men_n813_), .B(men_men_n561_), .C(men_men_n400_), .D(men_men_n50_), .Y(men_men_n830_));
  NO2        u0781(.A(men_men_n599_), .B(men_men_n179_), .Y(men_men_n831_));
  NA3        u0782(.A(men_men_n831_), .B(men_men_n592_), .C(x7), .Y(men_men_n832_));
  INV        u0783(.A(men_men_n832_), .Y(men_men_n833_));
  OAI210     u0784(.A0(men_men_n833_), .A1(men_men_n830_), .B0(men_men_n74_), .Y(men_men_n834_));
  NA2        u0785(.A(men_men_n688_), .B(x2), .Y(men_men_n835_));
  NO2        u0786(.A(men_men_n835_), .B(men_men_n58_), .Y(men_men_n836_));
  NO2        u0787(.A(x5), .B(men_men_n53_), .Y(men_men_n837_));
  NAi21      u0788(.An(x1), .B(x4), .Y(men_men_n838_));
  NA2        u0789(.A(men_men_n838_), .B(men_men_n764_), .Y(men_men_n839_));
  NO3        u0790(.A(men_men_n839_), .B(men_men_n188_), .C(men_men_n837_), .Y(men_men_n840_));
  OAI210     u0791(.A0(men_men_n840_), .A1(men_men_n836_), .B0(men_men_n363_), .Y(men_men_n841_));
  NA3        u0792(.A(men_men_n350_), .B(men_men_n665_), .C(men_men_n57_), .Y(men_men_n842_));
  NA3        u0793(.A(men_men_n842_), .B(men_men_n841_), .C(men_men_n834_), .Y(men_men_n843_));
  AOI210     u0794(.A0(men_men_n829_), .A1(x6), .B0(men_men_n843_), .Y(men_men_n844_));
  NA3        u0795(.A(men_men_n844_), .B(men_men_n811_), .C(men_men_n802_), .Y(men10));
  NO2        u0796(.A(x4), .B(x1), .Y(men_men_n846_));
  NO2        u0797(.A(men_men_n846_), .B(men_men_n138_), .Y(men_men_n847_));
  NA3        u0798(.A(x5), .B(x4), .C(x0), .Y(men_men_n848_));
  OAI220     u0799(.A0(men_men_n848_), .A1(men_men_n250_), .B0(men_men_n625_), .B1(men_men_n223_), .Y(men_men_n849_));
  NA2        u0800(.A(men_men_n849_), .B(men_men_n847_), .Y(men_men_n850_));
  NO3        u0801(.A(men_men_n318_), .B(men_men_n293_), .C(men_men_n83_), .Y(men_men_n851_));
  NA3        u0802(.A(men_men_n851_), .B(men_men_n336_), .C(men_men_n61_), .Y(men_men_n852_));
  AOI210     u0803(.A0(men_men_n852_), .A1(men_men_n850_), .B0(men_men_n275_), .Y(men_men_n853_));
  NOi21      u0804(.An(men_men_n234_), .B(men_men_n127_), .Y(men_men_n854_));
  AOI210     u0805(.A0(men_men_n443_), .A1(men_men_n550_), .B0(men_men_n297_), .Y(men_men_n855_));
  NO2        u0806(.A(men_men_n791_), .B(men_men_n309_), .Y(men_men_n856_));
  NOi31      u0807(.An(men_men_n856_), .B(men_men_n855_), .C(men_men_n854_), .Y(men_men_n857_));
  NA2        u0808(.A(x4), .B(men_men_n99_), .Y(men_men_n858_));
  NO2        u0809(.A(men_men_n295_), .B(men_men_n858_), .Y(men_men_n859_));
  NA2        u0810(.A(men_men_n88_), .B(x5), .Y(men_men_n860_));
  NO3        u0811(.A(men_men_n860_), .B(men_men_n100_), .C(men_men_n55_), .Y(men_men_n861_));
  NO3        u0812(.A(men_men_n861_), .B(men_men_n859_), .C(men_men_n857_), .Y(men_men_n862_));
  NA2        u0813(.A(men_men_n537_), .B(men_men_n245_), .Y(men_men_n863_));
  OAI220     u0814(.A0(men_men_n808_), .A1(men_men_n96_), .B0(men_men_n769_), .B1(men_men_n392_), .Y(men_men_n864_));
  NA2        u0815(.A(men_men_n864_), .B(men_men_n252_), .Y(men_men_n865_));
  OAI210     u0816(.A0(men_men_n862_), .A1(men_men_n338_), .B0(men_men_n865_), .Y(men_men_n866_));
  OAI210     u0817(.A0(men_men_n866_), .A1(men_men_n853_), .B0(x7), .Y(men_men_n867_));
  NA2        u0818(.A(men_men_n55_), .B(men_men_n67_), .Y(men_men_n868_));
  AOI210     u0819(.A0(men_men_n392_), .A1(men_men_n317_), .B0(men_men_n858_), .Y(men_men_n869_));
  NO3        u0820(.A(men_men_n394_), .B(men_men_n784_), .C(x5), .Y(men_men_n870_));
  OAI210     u0821(.A0(men_men_n870_), .A1(men_men_n869_), .B0(men_men_n868_), .Y(men_men_n871_));
  NO2        u0822(.A(men_men_n318_), .B(men_men_n130_), .Y(men_men_n872_));
  NA2        u0823(.A(men_men_n872_), .B(men_men_n374_), .Y(men_men_n873_));
  AOI210     u0824(.A0(men_men_n873_), .A1(men_men_n871_), .B0(x3), .Y(men_men_n874_));
  NA2        u0825(.A(men_men_n617_), .B(men_men_n226_), .Y(men_men_n875_));
  NO2        u0826(.A(x5), .B(men_men_n99_), .Y(men_men_n876_));
  NO2        u0827(.A(men_men_n875_), .B(men_men_n630_), .Y(men_men_n877_));
  OAI210     u0828(.A0(men_men_n877_), .A1(men_men_n874_), .B0(men_men_n825_), .Y(men_men_n878_));
  NO2        u0829(.A(x4), .B(x3), .Y(men_men_n879_));
  NA2        u0830(.A(men_men_n251_), .B(men_men_n385_), .Y(men_men_n880_));
  AOI210     u0831(.A0(men_men_n351_), .A1(men_men_n116_), .B0(men_men_n227_), .Y(men_men_n881_));
  NA2        u0832(.A(men_men_n846_), .B(men_men_n55_), .Y(men_men_n882_));
  NO2        u0833(.A(men_men_n466_), .B(men_men_n321_), .Y(men_men_n883_));
  NO3        u0834(.A(x4), .B(men_men_n99_), .C(men_men_n59_), .Y(men_men_n884_));
  NO2        u0835(.A(men_men_n386_), .B(x1), .Y(men_men_n885_));
  NOi31      u0836(.An(men_men_n884_), .B(men_men_n885_), .C(men_men_n883_), .Y(men_men_n886_));
  NA2        u0837(.A(men_men_n55_), .B(x5), .Y(men_men_n887_));
  NO2        u0838(.A(men_men_n886_), .B(men_men_n881_), .Y(men_men_n888_));
  AOI210     u0839(.A0(men_men_n888_), .A1(men_men_n880_), .B0(men_men_n193_), .Y(men_men_n889_));
  NO2        u0840(.A(men_men_n588_), .B(men_men_n442_), .Y(men_men_n890_));
  NO2        u0841(.A(x6), .B(x2), .Y(men_men_n891_));
  NO3        u0842(.A(men_men_n891_), .B(men_men_n617_), .C(men_men_n60_), .Y(men_men_n892_));
  OAI210     u0843(.A0(men_men_n892_), .A1(men_men_n890_), .B0(men_men_n244_), .Y(men_men_n893_));
  NO2        u0844(.A(men_men_n769_), .B(men_men_n392_), .Y(men_men_n894_));
  NA3        u0845(.A(x4), .B(x3), .C(men_men_n99_), .Y(men_men_n895_));
  NO3        u0846(.A(men_men_n895_), .B(men_men_n623_), .C(men_men_n407_), .Y(men_men_n896_));
  AOI210     u0847(.A0(men_men_n894_), .A1(men_men_n414_), .B0(men_men_n896_), .Y(men_men_n897_));
  AOI210     u0848(.A0(men_men_n897_), .A1(men_men_n893_), .B0(men_men_n400_), .Y(men_men_n898_));
  NO2        u0849(.A(men_men_n55_), .B(men_men_n56_), .Y(men_men_n899_));
  OAI220     u0850(.A0(men_men_n730_), .A1(men_men_n402_), .B0(men_men_n667_), .B1(men_men_n116_), .Y(men_men_n900_));
  NOi21      u0851(.An(men_men_n112_), .B(men_men_n111_), .Y(men_men_n901_));
  NO2        u0852(.A(men_men_n311_), .B(men_men_n295_), .Y(men_men_n902_));
  NA2        u0853(.A(men_men_n900_), .B(men_men_n105_), .Y(men_men_n903_));
  INV        u0854(.A(men_men_n903_), .Y(men_men_n904_));
  NA2        u0855(.A(men_men_n459_), .B(men_men_n236_), .Y(men_men_n905_));
  NO2        u0856(.A(men_men_n429_), .B(men_men_n519_), .Y(men_men_n906_));
  NA3        u0857(.A(men_men_n906_), .B(men_men_n905_), .C(men_men_n55_), .Y(men_men_n907_));
  NO2        u0858(.A(men_men_n172_), .B(men_men_n99_), .Y(men_men_n908_));
  NA3        u0859(.A(men_men_n908_), .B(men_men_n171_), .C(men_men_n111_), .Y(men_men_n909_));
  NA2        u0860(.A(men_men_n909_), .B(men_men_n907_), .Y(men_men_n910_));
  NO4        u0861(.A(men_men_n910_), .B(men_men_n904_), .C(men_men_n898_), .D(men_men_n889_), .Y(men_men_n911_));
  NA3        u0862(.A(men_men_n911_), .B(men_men_n878_), .C(men_men_n867_), .Y(men11));
  NA2        u0863(.A(men_men_n329_), .B(men_men_n83_), .Y(men_men_n913_));
  INV        u0864(.A(men_men_n785_), .Y(men_men_n914_));
  OAI220     u0865(.A0(men_men_n914_), .A1(men_men_n53_), .B0(men_men_n913_), .B1(men_men_n325_), .Y(men_men_n915_));
  NO2        u0866(.A(men_men_n683_), .B(x5), .Y(men_men_n916_));
  NO2        u0867(.A(men_men_n158_), .B(men_men_n472_), .Y(men_men_n917_));
  AOI220     u0868(.A0(men_men_n917_), .A1(men_men_n916_), .B0(men_men_n915_), .B1(x5), .Y(men_men_n918_));
  OAI220     u0869(.A0(men_men_n854_), .A1(men_men_n199_), .B0(men_men_n197_), .B1(men_men_n172_), .Y(men_men_n919_));
  NO2        u0870(.A(men_men_n308_), .B(men_men_n375_), .Y(men_men_n920_));
  AOI220     u0871(.A0(men_men_n920_), .A1(men_men_n170_), .B0(men_men_n919_), .B1(men_men_n154_), .Y(men_men_n921_));
  NO2        u0872(.A(men_men_n921_), .B(men_men_n394_), .Y(men_men_n922_));
  NO2        u0873(.A(men_men_n227_), .B(x2), .Y(men_men_n923_));
  OAI210     u0874(.A0(men_men_n803_), .A1(men_men_n923_), .B0(men_men_n364_), .Y(men_men_n924_));
  NO2        u0875(.A(men_men_n55_), .B(men_men_n97_), .Y(men_men_n925_));
  NA2        u0876(.A(men_men_n252_), .B(men_men_n925_), .Y(men_men_n926_));
  NO2        u0877(.A(men_men_n67_), .B(x1), .Y(men_men_n927_));
  NA2        u0878(.A(men_men_n927_), .B(men_men_n72_), .Y(men_men_n928_));
  OA220      u0879(.A0(men_men_n928_), .A1(men_men_n544_), .B0(men_men_n926_), .B1(men_men_n472_), .Y(men_men_n929_));
  AOI210     u0880(.A0(men_men_n929_), .A1(men_men_n924_), .B0(men_men_n630_), .Y(men_men_n930_));
  NO2        u0881(.A(men_men_n276_), .B(men_men_n53_), .Y(men_men_n931_));
  NO2        u0882(.A(men_men_n385_), .B(x3), .Y(men_men_n932_));
  NA3        u0883(.A(men_men_n932_), .B(men_men_n931_), .C(men_men_n784_), .Y(men_men_n933_));
  AOI210     u0884(.A0(men_men_n933_), .A1(men_men_n822_), .B0(men_men_n349_), .Y(men_men_n934_));
  NA2        u0885(.A(men_men_n99_), .B(x1), .Y(men_men_n935_));
  NO2        u0886(.A(men_men_n550_), .B(men_men_n200_), .Y(men_men_n936_));
  NA4        u0887(.A(men_men_n936_), .B(men_men_n777_), .C(men_men_n411_), .D(men_men_n935_), .Y(men_men_n937_));
  NA3        u0888(.A(x6), .B(x5), .C(men_men_n99_), .Y(men_men_n938_));
  NO2        u0889(.A(men_men_n938_), .B(men_men_n250_), .Y(men_men_n939_));
  NO2        u0890(.A(men_men_n394_), .B(x0), .Y(men_men_n940_));
  NOi31      u0891(.An(men_men_n940_), .B(men_men_n162_), .C(men_men_n51_), .Y(men_men_n941_));
  AOI210     u0892(.A0(men_men_n939_), .A1(men_men_n168_), .B0(men_men_n941_), .Y(men_men_n942_));
  NA2        u0893(.A(men_men_n942_), .B(men_men_n937_), .Y(men_men_n943_));
  NO4        u0894(.A(men_men_n943_), .B(men_men_n934_), .C(men_men_n930_), .D(men_men_n922_), .Y(men_men_n944_));
  OAI210     u0895(.A0(men_men_n918_), .A1(men_men_n131_), .B0(men_men_n944_), .Y(men_men_n945_));
  NA2        u0896(.A(men_men_n762_), .B(men_men_n79_), .Y(men_men_n946_));
  NO2        u0897(.A(x8), .B(x1), .Y(men_men_n947_));
  OAI210     u0898(.A0(men_men_n71_), .A1(men_men_n53_), .B0(x1), .Y(men_men_n948_));
  OAI210     u0899(.A0(men_men_n112_), .A1(x3), .B0(men_men_n948_), .Y(men_men_n949_));
  NO2        u0900(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n950_));
  OAI210     u0901(.A0(men_men_n950_), .A1(x2), .B0(men_men_n212_), .Y(men_men_n951_));
  NO2        u0902(.A(men_men_n538_), .B(men_men_n211_), .Y(men_men_n952_));
  INV        u0903(.A(men_men_n952_), .Y(men_men_n953_));
  NO2        u0904(.A(men_men_n459_), .B(x4), .Y(men_men_n954_));
  NO3        u0905(.A(men_men_n55_), .B(x6), .C(x1), .Y(men_men_n955_));
  NA2        u0906(.A(men_men_n954_), .B(men_men_n510_), .Y(men_men_n956_));
  NA2        u0907(.A(men_men_n956_), .B(men_men_n953_), .Y(men_men_n957_));
  AOI210     u0908(.A0(men_men_n949_), .A1(x2), .B0(men_men_n957_), .Y(men_men_n958_));
  NO2        u0909(.A(men_men_n211_), .B(x2), .Y(men_men_n959_));
  NA2        u0910(.A(men_men_n959_), .B(men_men_n879_), .Y(men_men_n960_));
  NOi21      u0911(.An(men_men_n340_), .B(men_men_n501_), .Y(men_men_n961_));
  NO3        u0912(.A(men_men_n961_), .B(men_men_n537_), .C(men_men_n295_), .Y(men_men_n962_));
  NA2        u0913(.A(x8), .B(men_men_n99_), .Y(men_men_n963_));
  OAI220     u0914(.A0(men_men_n630_), .A1(men_men_n963_), .B0(men_men_n295_), .B1(men_men_n336_), .Y(men_men_n964_));
  OAI210     u0915(.A0(men_men_n964_), .A1(men_men_n962_), .B0(men_men_n67_), .Y(men_men_n965_));
  NO2        u0916(.A(men_men_n97_), .B(x1), .Y(men_men_n966_));
  NA2        u0917(.A(men_men_n966_), .B(x7), .Y(men_men_n967_));
  AOI210     u0918(.A0(men_men_n965_), .A1(men_men_n960_), .B0(men_men_n967_), .Y(men_men_n968_));
  INV        u0919(.A(men_men_n224_), .Y(men_men_n969_));
  NA2        u0920(.A(men_men_n969_), .B(men_men_n138_), .Y(men_men_n970_));
  OAI220     u0921(.A0(men_men_n970_), .A1(men_men_n325_), .B0(x6), .B1(men_men_n295_), .Y(men_men_n971_));
  NO2        u0922(.A(men_men_n148_), .B(men_men_n55_), .Y(men_men_n972_));
  AOI210     u0923(.A0(men_men_n972_), .A1(men_men_n971_), .B0(men_men_n968_), .Y(men_men_n973_));
  OAI210     u0924(.A0(men_men_n958_), .A1(men_men_n751_), .B0(men_men_n973_), .Y(men_men_n974_));
  AO210      u0925(.A0(men_men_n945_), .A1(men_men_n57_), .B0(men_men_n974_), .Y(men12));
  NA2        u0926(.A(men_men_n776_), .B(men_men_n223_), .Y(men_men_n976_));
  NA2        u0927(.A(men_men_n622_), .B(men_men_n769_), .Y(men_men_n977_));
  NO2        u0928(.A(men_men_n976_), .B(men_men_n977_), .Y(men_men_n978_));
  NOi21      u0929(.An(men_men_n354_), .B(men_men_n489_), .Y(men_men_n979_));
  NO2        u0930(.A(x7), .B(men_men_n50_), .Y(men_men_n980_));
  NO2        u0931(.A(men_men_n538_), .B(men_men_n980_), .Y(men_men_n981_));
  NO3        u0932(.A(men_men_n764_), .B(men_men_n101_), .C(men_men_n88_), .Y(men_men_n982_));
  AOI210     u0933(.A0(men_men_n981_), .A1(men_men_n885_), .B0(men_men_n982_), .Y(men_men_n983_));
  NA2        u0934(.A(men_men_n925_), .B(men_men_n56_), .Y(men_men_n984_));
  OAI220     u0935(.A0(men_men_n984_), .A1(men_men_n511_), .B0(men_men_n983_), .B1(men_men_n979_), .Y(men_men_n985_));
  OAI210     u0936(.A0(men_men_n985_), .A1(men_men_n978_), .B0(men_men_n515_), .Y(men_men_n986_));
  NA2        u0937(.A(men_men_n79_), .B(x5), .Y(men_men_n987_));
  NA2        u0938(.A(men_men_n295_), .B(men_men_n640_), .Y(men_men_n988_));
  AOI210     u0939(.A0(men_men_n732_), .A1(men_men_n106_), .B0(men_men_n988_), .Y(men_men_n989_));
  NA2        u0940(.A(men_men_n536_), .B(men_men_n53_), .Y(men_men_n990_));
  NA2        u0941(.A(men_men_n259_), .B(men_men_n50_), .Y(men_men_n991_));
  OAI220     u0942(.A0(men_men_n991_), .A1(men_men_n282_), .B0(men_men_n990_), .B1(men_men_n124_), .Y(men_men_n992_));
  INV        u0943(.A(men_men_n454_), .Y(men_men_n993_));
  NO4        u0944(.A(men_men_n217_), .B(men_men_n244_), .C(men_men_n60_), .D(men_men_n57_), .Y(men_men_n994_));
  AOI220     u0945(.A0(men_men_n994_), .A1(men_men_n993_), .B0(men_men_n992_), .B1(men_men_n56_), .Y(men_men_n995_));
  OAI210     u0946(.A0(men_men_n989_), .A1(men_men_n63_), .B0(men_men_n995_), .Y(men_men_n996_));
  NO2        u0947(.A(men_men_n57_), .B(x0), .Y(men_men_n997_));
  NO2        u0948(.A(men_men_n588_), .B(men_men_n293_), .Y(men_men_n998_));
  NO2        u0949(.A(men_men_n667_), .B(x3), .Y(men_men_n999_));
  NO2        u0950(.A(men_men_n586_), .B(x8), .Y(men_men_n1000_));
  AOI220     u0951(.A0(men_men_n1000_), .A1(men_men_n999_), .B0(men_men_n998_), .B1(men_men_n997_), .Y(men_men_n1001_));
  NO2        u0952(.A(men_men_n539_), .B(x8), .Y(men_men_n1002_));
  NA3        u0953(.A(men_men_n584_), .B(men_men_n191_), .C(x0), .Y(men_men_n1003_));
  OAI220     u0954(.A0(men_men_n1003_), .A1(men_men_n1002_), .B0(men_men_n1001_), .B1(men_men_n509_), .Y(men_men_n1004_));
  AOI210     u0955(.A0(men_men_n996_), .A1(men_men_n891_), .B0(men_men_n1004_), .Y(men_men_n1005_));
  NO2        u0956(.A(men_men_n223_), .B(men_men_n55_), .Y(men_men_n1006_));
  NO2        u0957(.A(men_men_n231_), .B(x8), .Y(men_men_n1007_));
  NOi32      u0958(.An(men_men_n1007_), .Bn(men_men_n190_), .C(men_men_n502_), .Y(men_men_n1008_));
  NO2        u0959(.A(men_men_n80_), .B(men_men_n60_), .Y(men_men_n1009_));
  OAI210     u0960(.A0(men_men_n1008_), .A1(men_men_n1006_), .B0(men_men_n1009_), .Y(men_men_n1010_));
  NO2        u0961(.A(men_men_n825_), .B(men_men_n89_), .Y(men_men_n1011_));
  NO2        u0962(.A(men_men_n157_), .B(men_men_n53_), .Y(men_men_n1012_));
  AOI210     u0963(.A0(men_men_n308_), .A1(x8), .B0(men_men_n1012_), .Y(men_men_n1013_));
  AOI210     u0964(.A0(men_men_n199_), .A1(men_men_n87_), .B0(men_men_n1013_), .Y(men_men_n1014_));
  OAI210     u0965(.A0(men_men_n1014_), .A1(men_men_n1011_), .B0(men_men_n599_), .Y(men_men_n1015_));
  NO2        u0966(.A(x7), .B(x0), .Y(men_men_n1016_));
  XN2        u0967(.A(x8), .B(x7), .Y(men_men_n1017_));
  NO2        u0968(.A(men_men_n241_), .B(men_men_n237_), .Y(men_men_n1018_));
  NO2        u0969(.A(men_men_n97_), .B(x4), .Y(men_men_n1019_));
  OAI210     u0970(.A0(men_men_n1018_), .A1(men_men_n251_), .B0(men_men_n1019_), .Y(men_men_n1020_));
  NA3        u0971(.A(men_men_n1020_), .B(men_men_n1015_), .C(men_men_n1010_), .Y(men_men_n1021_));
  NA2        u0972(.A(men_men_n1021_), .B(men_men_n492_), .Y(men_men_n1022_));
  NO2        u0973(.A(men_men_n55_), .B(x4), .Y(men_men_n1023_));
  NA2        u0974(.A(men_men_n1023_), .B(men_men_n153_), .Y(men_men_n1024_));
  NO2        u0975(.A(men_men_n234_), .B(men_men_n380_), .Y(men_men_n1025_));
  OAI220     u0976(.A0(men_men_n261_), .A1(men_men_n249_), .B0(men_men_n237_), .B1(men_men_n219_), .Y(men_men_n1026_));
  NA3        u0977(.A(men_men_n1026_), .B(men_men_n599_), .C(x1), .Y(men_men_n1027_));
  OAI210     u0978(.A0(x8), .A1(x0), .B0(x4), .Y(men_men_n1028_));
  NO2        u0979(.A(x7), .B(men_men_n56_), .Y(men_men_n1029_));
  NO2        u0980(.A(men_men_n65_), .B(men_men_n1029_), .Y(men_men_n1030_));
  NO2        u0981(.A(men_men_n590_), .B(men_men_n295_), .Y(men_men_n1031_));
  NO2        u0982(.A(men_men_n131_), .B(men_men_n130_), .Y(men_men_n1032_));
  NO2        u0983(.A(men_men_n538_), .B(men_men_n392_), .Y(men_men_n1033_));
  OAI210     u0984(.A0(men_men_n1033_), .A1(men_men_n1032_), .B0(men_men_n231_), .Y(men_men_n1034_));
  NA2        u0985(.A(men_men_n296_), .B(men_men_n59_), .Y(men_men_n1035_));
  NA2        u0986(.A(men_men_n1034_), .B(men_men_n1027_), .Y(men_men_n1036_));
  OAI210     u0987(.A0(men_men_n1036_), .A1(men_men_n1025_), .B0(men_men_n601_), .Y(men_men_n1037_));
  NA4        u0988(.A(men_men_n1037_), .B(men_men_n1022_), .C(men_men_n1005_), .D(men_men_n986_), .Y(men13));
  NO2        u0989(.A(men_men_n407_), .B(men_men_n314_), .Y(men_men_n1039_));
  NO2        u0990(.A(men_men_n764_), .B(men_men_n172_), .Y(men_men_n1040_));
  NO2        u0991(.A(men_men_n147_), .B(men_men_n67_), .Y(men_men_n1041_));
  XN2        u0992(.A(x4), .B(x0), .Y(men_men_n1042_));
  NO3        u0993(.A(men_men_n1042_), .B(men_men_n100_), .C(men_men_n371_), .Y(men_men_n1043_));
  AO220      u0994(.A0(men_men_n1043_), .A1(men_men_n1041_), .B0(men_men_n1040_), .B1(men_men_n297_), .Y(men_men_n1044_));
  NA2        u0995(.A(men_men_n1044_), .B(x3), .Y(men_men_n1045_));
  NO2        u0996(.A(men_men_n764_), .B(x6), .Y(men_men_n1046_));
  NO2        u0997(.A(men_men_n991_), .B(men_men_n347_), .Y(men_men_n1047_));
  NO3        u0998(.A(x8), .B(x5), .C(men_men_n99_), .Y(men_men_n1048_));
  NA2        u0999(.A(men_men_n1048_), .B(men_men_n570_), .Y(men_men_n1049_));
  NO2        u1000(.A(men_men_n538_), .B(men_men_n185_), .Y(men_men_n1050_));
  NA2        u1001(.A(men_men_n396_), .B(men_men_n53_), .Y(men_men_n1051_));
  NO2        u1002(.A(men_men_n1051_), .B(men_men_n818_), .Y(men_men_n1052_));
  NA2        u1003(.A(men_men_n56_), .B(men_men_n99_), .Y(men_men_n1053_));
  NA2        u1004(.A(men_men_n1053_), .B(x1), .Y(men_men_n1054_));
  NO2        u1005(.A(men_men_n293_), .B(x6), .Y(men_men_n1055_));
  OAI210     u1006(.A0(men_men_n227_), .A1(men_men_n858_), .B0(men_men_n835_), .Y(men_men_n1056_));
  NA2        u1007(.A(men_men_n1056_), .B(men_men_n1055_), .Y(men_men_n1057_));
  NAi31      u1008(.An(men_men_n1052_), .B(men_men_n1057_), .C(men_men_n1049_), .Y(men_men_n1058_));
  AOI220     u1009(.A0(men_men_n1058_), .A1(men_men_n65_), .B0(men_men_n1047_), .B1(men_men_n1046_), .Y(men_men_n1059_));
  NA2        u1010(.A(men_men_n67_), .B(x3), .Y(men_men_n1060_));
  NA2        u1011(.A(men_men_n1060_), .B(men_men_n793_), .Y(men_men_n1061_));
  OAI220     u1012(.A0(men_men_n275_), .A1(men_men_n728_), .B0(men_men_n79_), .B1(men_men_n71_), .Y(men_men_n1062_));
  AOI210     u1013(.A0(men_men_n987_), .A1(men_men_n548_), .B0(men_men_n858_), .Y(men_men_n1063_));
  OA210      u1014(.A0(men_men_n1062_), .A1(men_men_n1061_), .B0(men_men_n1063_), .Y(men_men_n1064_));
  NA2        u1015(.A(men_men_n550_), .B(men_men_n55_), .Y(men_men_n1065_));
  NA2        u1016(.A(men_men_n447_), .B(men_men_n437_), .Y(men_men_n1066_));
  NA2        u1017(.A(x6), .B(men_men_n50_), .Y(men_men_n1067_));
  NA2        u1018(.A(men_men_n1067_), .B(men_men_n478_), .Y(men_men_n1068_));
  NO2        u1019(.A(men_men_n150_), .B(men_men_n119_), .Y(men_men_n1069_));
  AOI210     u1020(.A0(men_men_n1068_), .A1(men_men_n381_), .B0(men_men_n1069_), .Y(men_men_n1070_));
  OAI220     u1021(.A0(men_men_n1070_), .A1(men_men_n769_), .B0(men_men_n1066_), .B1(men_men_n1065_), .Y(men_men_n1071_));
  OAI210     u1022(.A0(men_men_n1071_), .A1(men_men_n1064_), .B0(men_men_n1016_), .Y(men_men_n1072_));
  NAi21      u1023(.An(men_men_n76_), .B(men_men_n336_), .Y(men_men_n1073_));
  NO2        u1024(.A(men_men_n1073_), .B(men_men_n67_), .Y(men_men_n1074_));
  AOI210     u1025(.A0(men_men_n153_), .A1(x4), .B0(men_men_n164_), .Y(men_men_n1075_));
  NO2        u1026(.A(men_men_n1075_), .B(x0), .Y(men_men_n1076_));
  NO2        u1027(.A(men_men_n160_), .B(men_men_n266_), .Y(men_men_n1077_));
  OAI210     u1028(.A0(men_men_n1077_), .A1(men_men_n1076_), .B0(men_men_n1074_), .Y(men_men_n1078_));
  NO2        u1029(.A(x4), .B(x0), .Y(men_men_n1079_));
  NO3        u1030(.A(men_men_n876_), .B(men_men_n224_), .C(men_men_n478_), .Y(men_men_n1080_));
  OAI210     u1031(.A0(men_men_n1080_), .A1(men_men_n186_), .B0(men_men_n1079_), .Y(men_men_n1081_));
  NA2        u1032(.A(men_men_n1081_), .B(men_men_n1078_), .Y(men_men_n1082_));
  NA2        u1033(.A(men_men_n226_), .B(men_men_n653_), .Y(men_men_n1083_));
  INV        u1034(.A(men_men_n1083_), .Y(men_men_n1084_));
  NA2        u1035(.A(men_men_n56_), .B(x0), .Y(men_men_n1085_));
  NO3        u1036(.A(men_men_n1085_), .B(men_men_n437_), .C(men_men_n73_), .Y(men_men_n1086_));
  OAI210     u1037(.A0(men_men_n1086_), .A1(men_men_n1084_), .B0(x2), .Y(men_men_n1087_));
  NO2        u1038(.A(men_men_n701_), .B(x1), .Y(men_men_n1088_));
  AOI220     u1039(.A0(men_men_n1088_), .A1(men_men_n543_), .B0(men_men_n422_), .B1(men_men_n267_), .Y(men_men_n1089_));
  NA2        u1040(.A(men_men_n1089_), .B(men_men_n1087_), .Y(men_men_n1090_));
  AOI220     u1041(.A0(men_men_n1090_), .A1(men_men_n120_), .B0(men_men_n1082_), .B1(men_men_n64_), .Y(men_men_n1091_));
  NA4        u1042(.A(men_men_n1091_), .B(men_men_n1072_), .C(men_men_n1059_), .D(men_men_n1045_), .Y(men14));
  NO3        u1043(.A(x7), .B(x6), .C(x0), .Y(men_men_n1093_));
  AOI210     u1044(.A0(men_men_n2324_), .A1(men_men_n2313_), .B0(men_men_n146_), .Y(men_men_n1094_));
  AOI220     u1045(.A0(men_men_n328_), .A1(men_men_n751_), .B0(men_men_n396_), .B1(men_men_n371_), .Y(men_men_n1095_));
  NA2        u1046(.A(men_men_n252_), .B(men_men_n854_), .Y(men_men_n1096_));
  OAI220     u1047(.A0(men_men_n1096_), .A1(men_men_n1095_), .B0(men_men_n410_), .B1(men_men_n714_), .Y(men_men_n1097_));
  OA210      u1048(.A0(men_men_n1097_), .A1(men_men_n1094_), .B0(x4), .Y(men_men_n1098_));
  NO2        u1049(.A(men_men_n130_), .B(men_men_n541_), .Y(men_men_n1099_));
  NA2        u1050(.A(x6), .B(x2), .Y(men_men_n1100_));
  INV        u1051(.A(men_men_n1100_), .Y(men_men_n1101_));
  OA210      u1052(.A0(men_men_n1099_), .A1(men_men_n196_), .B0(men_men_n1101_), .Y(men_men_n1102_));
  NO4        u1053(.A(men_men_n538_), .B(men_men_n329_), .C(men_men_n271_), .D(men_men_n105_), .Y(men_men_n1103_));
  OAI210     u1054(.A0(men_men_n1103_), .A1(men_men_n1102_), .B0(men_men_n59_), .Y(men_men_n1104_));
  NA2        u1055(.A(x6), .B(men_men_n97_), .Y(men_men_n1105_));
  NO2        u1056(.A(men_men_n588_), .B(men_men_n1105_), .Y(men_men_n1106_));
  NA2        u1057(.A(men_men_n1106_), .B(men_men_n806_), .Y(men_men_n1107_));
  AOI210     u1058(.A0(men_men_n1000_), .A1(men_men_n884_), .B0(x1), .Y(men_men_n1108_));
  NO2        u1059(.A(men_men_n475_), .B(x5), .Y(men_men_n1109_));
  AN2        u1060(.A(men_men_n1108_), .B(men_men_n1107_), .Y(men_men_n1110_));
  NO2        u1061(.A(men_men_n623_), .B(men_men_n963_), .Y(men_men_n1111_));
  NO2        u1062(.A(men_men_n71_), .B(men_men_n58_), .Y(men_men_n1112_));
  OAI210     u1063(.A0(men_men_n1111_), .A1(men_men_n393_), .B0(men_men_n1112_), .Y(men_men_n1113_));
  AOI220     u1064(.A0(x1), .A1(men_men_n1113_), .B0(men_men_n1110_), .B1(men_men_n1104_), .Y(men_men_n1114_));
  NO2        u1065(.A(men_men_n600_), .B(men_men_n157_), .Y(men_men_n1115_));
  NO3        u1066(.A(men_men_n1115_), .B(men_men_n1114_), .C(men_men_n1098_), .Y(men_men_n1116_));
  NO2        u1067(.A(men_men_n293_), .B(x2), .Y(men_men_n1117_));
  XN2        u1068(.A(x4), .B(x1), .Y(men_men_n1118_));
  NO2        u1069(.A(men_men_n1118_), .B(men_men_n275_), .Y(men_men_n1119_));
  NOi21      u1070(.An(men_men_n1119_), .B(men_men_n359_), .Y(men_men_n1120_));
  NO2        u1071(.A(men_men_n307_), .B(men_men_n60_), .Y(men_men_n1121_));
  OAI210     u1072(.A0(men_men_n1121_), .A1(men_men_n1120_), .B0(men_men_n1117_), .Y(men_men_n1122_));
  NA2        u1073(.A(men_men_n610_), .B(men_men_n56_), .Y(men_men_n1123_));
  AOI220     u1074(.A0(men_men_n127_), .A1(men_men_n56_), .B0(men_men_n84_), .B1(x5), .Y(men_men_n1124_));
  NA2        u1075(.A(men_men_n955_), .B(men_men_n280_), .Y(men_men_n1125_));
  NA2        u1076(.A(men_men_n226_), .B(men_men_n316_), .Y(men_men_n1126_));
  NA2        u1077(.A(men_men_n569_), .B(men_men_n901_), .Y(men_men_n1127_));
  OAI220     u1078(.A0(men_men_n1127_), .A1(men_men_n1126_), .B0(men_men_n1125_), .B1(men_men_n1124_), .Y(men_men_n1128_));
  INV        u1079(.A(men_men_n1128_), .Y(men_men_n1129_));
  AOI210     u1080(.A0(men_men_n1129_), .A1(men_men_n1122_), .B0(x7), .Y(men_men_n1130_));
  NO2        u1081(.A(men_men_n436_), .B(x6), .Y(men_men_n1131_));
  AOI210     u1082(.A0(men_men_n724_), .A1(men_men_n837_), .B0(men_men_n1131_), .Y(men_men_n1132_));
  OAI220     u1083(.A0(men_men_n1132_), .A1(men_men_n55_), .B0(men_men_n436_), .B1(men_men_n93_), .Y(men_men_n1133_));
  NA2        u1084(.A(men_men_n1133_), .B(men_men_n318_), .Y(men_men_n1134_));
  NA3        u1085(.A(men_men_n544_), .B(men_men_n935_), .C(men_men_n66_), .Y(men_men_n1135_));
  NO4        u1086(.A(men_men_n1135_), .B(men_men_n1085_), .C(men_men_n109_), .D(men_men_n55_), .Y(men_men_n1136_));
  NO3        u1087(.A(men_men_n928_), .B(men_men_n730_), .C(men_men_n427_), .Y(men_men_n1137_));
  NO3        u1088(.A(men_men_n1137_), .B(men_men_n1136_), .C(men_men_n906_), .Y(men_men_n1138_));
  AOI210     u1089(.A0(men_men_n1138_), .A1(men_men_n1134_), .B0(men_men_n277_), .Y(men_men_n1139_));
  NA2        u1090(.A(men_men_n791_), .B(men_men_n53_), .Y(men_men_n1140_));
  OAI210     u1091(.A0(men_men_n221_), .A1(men_men_n106_), .B0(x2), .Y(men_men_n1141_));
  NA2        u1092(.A(men_men_n326_), .B(men_men_n56_), .Y(men_men_n1142_));
  OA210      u1093(.A0(men_men_n1142_), .A1(men_men_n1141_), .B0(men_men_n1140_), .Y(men_men_n1143_));
  NA3        u1094(.A(men_men_n906_), .B(men_men_n656_), .C(men_men_n55_), .Y(men_men_n1144_));
  NA2        u1095(.A(men_men_n56_), .B(x2), .Y(men_men_n1145_));
  NO2        u1096(.A(men_men_n1145_), .B(men_men_n184_), .Y(men_men_n1146_));
  NA4        u1097(.A(men_men_n1146_), .B(men_men_n326_), .C(men_men_n234_), .D(men_men_n64_), .Y(men_men_n1147_));
  NA3        u1098(.A(men_men_n1088_), .B(men_men_n550_), .C(men_men_n560_), .Y(men_men_n1148_));
  AN3        u1099(.A(men_men_n1148_), .B(men_men_n1147_), .C(men_men_n1144_), .Y(men_men_n1149_));
  OAI210     u1100(.A0(men_men_n1143_), .A1(men_men_n288_), .B0(men_men_n1149_), .Y(men_men_n1150_));
  NO3        u1101(.A(men_men_n1150_), .B(men_men_n1139_), .C(men_men_n1130_), .Y(men_men_n1151_));
  OAI210     u1102(.A0(men_men_n1116_), .A1(x3), .B0(men_men_n1151_), .Y(men15));
  NA2        u1103(.A(men_men_n520_), .B(men_men_n59_), .Y(men_men_n1153_));
  NAi41      u1104(.An(x2), .B(x7), .C(x6), .D(x0), .Y(men_men_n1154_));
  AOI210     u1105(.A0(men_men_n1154_), .A1(men_men_n1153_), .B0(men_men_n53_), .Y(men_men_n1155_));
  NA3        u1106(.A(men_men_n57_), .B(x6), .C(men_men_n99_), .Y(men_men_n1156_));
  NO2        u1107(.A(men_men_n1156_), .B(men_men_n266_), .Y(men_men_n1157_));
  OAI210     u1108(.A0(men_men_n1157_), .A1(men_men_n1155_), .B0(men_men_n1019_), .Y(men_men_n1158_));
  NA2        u1109(.A(men_men_n101_), .B(men_men_n99_), .Y(men_men_n1159_));
  AOI210     u1110(.A0(men_men_n652_), .A1(men_men_n70_), .B0(x3), .Y(men_men_n1160_));
  NA2        u1111(.A(men_men_n1160_), .B(men_men_n1158_), .Y(men_men_n1161_));
  AOI210     u1112(.A0(men_men_n940_), .A1(men_men_n524_), .B0(men_men_n50_), .Y(men_men_n1162_));
  NO2        u1113(.A(men_men_n215_), .B(x5), .Y(men_men_n1163_));
  NA3        u1114(.A(men_men_n1088_), .B(men_men_n554_), .C(men_men_n1029_), .Y(men_men_n1164_));
  NA2        u1115(.A(men_men_n1164_), .B(men_men_n1162_), .Y(men_men_n1165_));
  NA2        u1116(.A(men_men_n301_), .B(men_men_n309_), .Y(men_men_n1166_));
  AOI210     u1117(.A0(men_men_n1054_), .A1(men_men_n58_), .B0(men_men_n1166_), .Y(men_men_n1167_));
  NA4        u1118(.A(men_men_n1054_), .B(men_men_n622_), .C(men_men_n997_), .D(men_men_n336_), .Y(men_men_n1168_));
  NA2        u1119(.A(men_men_n524_), .B(men_men_n411_), .Y(men_men_n1169_));
  NO2        u1120(.A(men_men_n667_), .B(men_men_n53_), .Y(men_men_n1170_));
  NO2        u1121(.A(men_men_n691_), .B(men_men_n271_), .Y(men_men_n1171_));
  NA2        u1122(.A(men_men_n1171_), .B(men_men_n1170_), .Y(men_men_n1172_));
  NA3        u1123(.A(men_men_n1172_), .B(men_men_n1169_), .C(men_men_n1168_), .Y(men_men_n1173_));
  OAI210     u1124(.A0(men_men_n1173_), .A1(men_men_n1167_), .B0(men_men_n71_), .Y(men_men_n1174_));
  NO2        u1125(.A(men_men_n769_), .B(men_men_n50_), .Y(men_men_n1175_));
  NO2        u1126(.A(men_men_n223_), .B(men_men_n63_), .Y(men_men_n1176_));
  OA210      u1127(.A0(men_men_n1176_), .A1(men_men_n1175_), .B0(men_men_n359_), .Y(men_men_n1177_));
  NA2        u1128(.A(men_men_n57_), .B(x3), .Y(men_men_n1178_));
  NO2        u1129(.A(men_men_n1178_), .B(men_men_n605_), .Y(men_men_n1179_));
  OAI210     u1130(.A0(men_men_n1179_), .A1(men_men_n1177_), .B0(men_men_n891_), .Y(men_men_n1180_));
  NA2        u1131(.A(men_men_n1146_), .B(men_men_n65_), .Y(men_men_n1181_));
  NO2        u1132(.A(men_men_n380_), .B(men_men_n73_), .Y(men_men_n1182_));
  NO2        u1133(.A(men_men_n812_), .B(men_men_n67_), .Y(men_men_n1183_));
  NA2        u1134(.A(men_men_n1183_), .B(men_men_n1182_), .Y(men_men_n1184_));
  NO2        u1135(.A(men_men_n858_), .B(x6), .Y(men_men_n1185_));
  NA4        u1136(.A(men_men_n1185_), .B(men_men_n529_), .C(men_men_n148_), .D(men_men_n363_), .Y(men_men_n1186_));
  AN4        u1137(.A(men_men_n1186_), .B(men_men_n1184_), .C(men_men_n2309_), .D(men_men_n1181_), .Y(men_men_n1187_));
  NA3        u1138(.A(men_men_n1187_), .B(men_men_n1180_), .C(men_men_n1174_), .Y(men_men_n1188_));
  NO2        u1139(.A(men_men_n579_), .B(x2), .Y(men_men_n1189_));
  OAI210     u1140(.A0(men_men_n65_), .A1(men_men_n53_), .B0(men_men_n133_), .Y(men_men_n1190_));
  OAI210     u1141(.A0(men_men_n1189_), .A1(men_men_n77_), .B0(men_men_n1190_), .Y(men_men_n1191_));
  NO2        u1142(.A(men_men_n1191_), .B(men_men_n293_), .Y(men_men_n1192_));
  NO3        u1143(.A(men_men_n1156_), .B(men_men_n240_), .C(men_men_n223_), .Y(men_men_n1193_));
  NA3        u1144(.A(men_men_n57_), .B(x1), .C(x0), .Y(men_men_n1194_));
  NA3        u1145(.A(men_men_n67_), .B(x5), .C(x2), .Y(men_men_n1195_));
  NA4        u1146(.A(x7), .B(x3), .C(men_men_n53_), .D(x0), .Y(men_men_n1196_));
  OAI220     u1147(.A0(men_men_n1196_), .A1(x6), .B0(men_men_n1195_), .B1(men_men_n1194_), .Y(men_men_n1197_));
  NO2        u1148(.A(men_men_n1197_), .B(men_men_n1193_), .Y(men_men_n1198_));
  NAi21      u1149(.An(men_men_n105_), .B(men_men_n661_), .Y(men_men_n1199_));
  NA4        u1150(.A(men_men_n1199_), .B(men_men_n291_), .C(men_men_n261_), .D(men_men_n554_), .Y(men_men_n1200_));
  NA2        u1151(.A(men_men_n74_), .B(men_men_n50_), .Y(men_men_n1201_));
  NA2        u1152(.A(men_men_n1200_), .B(men_men_n1198_), .Y(men_men_n1202_));
  OAI210     u1153(.A0(men_men_n1202_), .A1(men_men_n1192_), .B0(men_men_n56_), .Y(men_men_n1203_));
  OAI220     u1154(.A0(men_men_n53_), .A1(men_men_n272_), .B0(men_men_n895_), .B1(men_men_n826_), .Y(men_men_n1204_));
  NA2        u1155(.A(men_men_n740_), .B(men_men_n356_), .Y(men_men_n1205_));
  OAI210     u1156(.A0(men_men_n1182_), .A1(men_men_n1176_), .B0(men_men_n262_), .Y(men_men_n1206_));
  OAI210     u1157(.A0(men_men_n1205_), .A1(men_men_n746_), .B0(men_men_n1206_), .Y(men_men_n1207_));
  OAI210     u1158(.A0(men_men_n1207_), .A1(men_men_n1204_), .B0(x6), .Y(men_men_n1208_));
  NO2        u1159(.A(men_men_n57_), .B(men_men_n59_), .Y(men_men_n1209_));
  NO2        u1160(.A(x7), .B(x5), .Y(men_men_n1210_));
  AOI220     u1161(.A0(men_men_n755_), .A1(men_men_n1209_), .B0(men_men_n477_), .B1(men_men_n1210_), .Y(men_men_n1211_));
  NA2        u1162(.A(men_men_n677_), .B(men_men_n262_), .Y(men_men_n1212_));
  NA2        u1163(.A(men_men_n1212_), .B(men_men_n1211_), .Y(men_men_n1213_));
  NA2        u1164(.A(men_men_n1213_), .B(men_men_n374_), .Y(men_men_n1214_));
  AOI210     u1165(.A0(men_men_n332_), .A1(men_men_n308_), .B0(men_men_n55_), .Y(men_men_n1215_));
  NA4        u1166(.A(men_men_n1215_), .B(men_men_n1214_), .C(men_men_n1208_), .D(men_men_n1203_), .Y(men_men_n1216_));
  AO220      u1167(.A0(men_men_n1216_), .A1(men_men_n1188_), .B0(men_men_n1165_), .B1(men_men_n1161_), .Y(men16));
  NO2        u1168(.A(x4), .B(men_men_n59_), .Y(men_men_n1218_));
  NA2        u1169(.A(men_men_n587_), .B(x3), .Y(men_men_n1219_));
  NA3        u1170(.A(men_men_n211_), .B(men_men_n381_), .C(men_men_n837_), .Y(men_men_n1220_));
  INV        u1171(.A(men_men_n122_), .Y(men_men_n1221_));
  AOI210     u1172(.A0(men_men_n1220_), .A1(men_men_n1219_), .B0(men_men_n1221_), .Y(men_men_n1222_));
  NO3        u1173(.A(x8), .B(x6), .C(men_men_n50_), .Y(men_men_n1223_));
  NO2        u1174(.A(men_men_n655_), .B(men_men_n175_), .Y(men_men_n1224_));
  OAI210     u1175(.A0(men_men_n1223_), .A1(men_men_n217_), .B0(men_men_n1224_), .Y(men_men_n1225_));
  NO2        u1176(.A(men_men_n150_), .B(x5), .Y(men_men_n1226_));
  NA2        u1177(.A(men_men_n1226_), .B(men_men_n1189_), .Y(men_men_n1227_));
  NA2        u1178(.A(men_men_n1227_), .B(men_men_n1225_), .Y(men_men_n1228_));
  OAI210     u1179(.A0(men_men_n1228_), .A1(men_men_n1222_), .B0(men_men_n1218_), .Y(men_men_n1229_));
  OAI210     u1180(.A0(men_men_n1117_), .A1(men_men_n806_), .B0(men_men_n371_), .Y(men_men_n1230_));
  NO2        u1181(.A(men_men_n293_), .B(x7), .Y(men_men_n1231_));
  NA2        u1182(.A(men_men_n1231_), .B(x0), .Y(men_men_n1232_));
  AOI210     u1183(.A0(men_men_n1232_), .A1(men_men_n1230_), .B0(men_men_n568_), .Y(men_men_n1233_));
  NA2        u1184(.A(men_men_n947_), .B(men_men_n185_), .Y(men_men_n1234_));
  NA2        u1185(.A(men_men_n55_), .B(men_men_n97_), .Y(men_men_n1235_));
  NA2        u1186(.A(men_men_n1235_), .B(men_men_n607_), .Y(men_men_n1236_));
  NA2        u1187(.A(men_men_n331_), .B(men_men_n950_), .Y(men_men_n1237_));
  OA210      u1188(.A0(men_men_n1237_), .A1(men_men_n1236_), .B0(men_men_n1234_), .Y(men_men_n1238_));
  OAI210     u1189(.A0(men_men_n1238_), .A1(men_men_n582_), .B0(men_men_n440_), .Y(men_men_n1239_));
  INV        u1190(.A(men_men_n891_), .Y(men_men_n1240_));
  NO2        u1191(.A(men_men_n1240_), .B(men_men_n61_), .Y(men_men_n1241_));
  AOI220     u1192(.A0(men_men_n1241_), .A1(men_men_n244_), .B0(men_men_n1106_), .B1(men_men_n115_), .Y(men_men_n1242_));
  NO2        u1193(.A(men_men_n1242_), .B(men_men_n282_), .Y(men_men_n1243_));
  NO3        u1194(.A(men_men_n1243_), .B(men_men_n1239_), .C(men_men_n1233_), .Y(men_men_n1244_));
  NO3        u1195(.A(x6), .B(x4), .C(x3), .Y(men_men_n1245_));
  NO2        u1196(.A(men_men_n645_), .B(x3), .Y(men_men_n1246_));
  AOI210     u1197(.A0(men_men_n586_), .A1(men_men_n137_), .B0(men_men_n935_), .Y(men_men_n1247_));
  OA210      u1198(.A0(men_men_n1246_), .A1(men_men_n374_), .B0(men_men_n1247_), .Y(men_men_n1248_));
  NO2        u1199(.A(men_men_n442_), .B(men_men_n69_), .Y(men_men_n1249_));
  INV        u1200(.A(men_men_n453_), .Y(men_men_n1250_));
  NO3        u1201(.A(men_men_n1250_), .B(men_men_n236_), .C(men_men_n145_), .Y(men_men_n1251_));
  NO3        u1202(.A(men_men_n1251_), .B(men_men_n1249_), .C(men_men_n1248_), .Y(men_men_n1252_));
  NA2        u1203(.A(men_men_n357_), .B(men_men_n837_), .Y(men_men_n1253_));
  NA4        u1204(.A(men_men_n427_), .B(men_men_n327_), .C(men_men_n203_), .D(x6), .Y(men_men_n1254_));
  OAI210     u1205(.A0(men_men_n645_), .A1(men_men_n1253_), .B0(men_men_n1254_), .Y(men_men_n1255_));
  NA2        u1206(.A(men_men_n796_), .B(men_men_n1145_), .Y(men_men_n1256_));
  NA2        u1207(.A(men_men_n653_), .B(x7), .Y(men_men_n1257_));
  OAI210     u1208(.A0(men_men_n1257_), .A1(men_men_n342_), .B0(men_men_n1256_), .Y(men_men_n1258_));
  NA2        u1209(.A(men_men_n250_), .B(x2), .Y(men_men_n1259_));
  NO2        u1210(.A(men_men_n1259_), .B(men_men_n68_), .Y(men_men_n1260_));
  OA210      u1211(.A0(men_men_n1105_), .A1(men_men_n58_), .B0(men_men_n692_), .Y(men_men_n1261_));
  NO2        u1212(.A(men_men_n1261_), .B(men_men_n179_), .Y(men_men_n1262_));
  NO4        u1213(.A(men_men_n1262_), .B(men_men_n1260_), .C(men_men_n1258_), .D(men_men_n1255_), .Y(men_men_n1263_));
  OA220      u1214(.A0(men_men_n1263_), .A1(men_men_n392_), .B0(men_men_n1252_), .B1(men_men_n192_), .Y(men_men_n1264_));
  NA2        u1215(.A(men_men_n368_), .B(men_men_n714_), .Y(men_men_n1265_));
  NO2        u1216(.A(men_men_n1265_), .B(x8), .Y(men_men_n1266_));
  NO3        u1217(.A(men_men_n838_), .B(men_men_n301_), .C(x8), .Y(men_men_n1267_));
  OAI210     u1218(.A0(men_men_n1267_), .A1(men_men_n1266_), .B0(x6), .Y(men_men_n1268_));
  OAI210     u1219(.A0(x2), .A1(men_men_n67_), .B0(men_men_n79_), .Y(men_men_n1269_));
  NA2        u1220(.A(men_men_n1269_), .B(men_men_n807_), .Y(men_men_n1270_));
  NA2        u1221(.A(men_men_n771_), .B(men_men_n67_), .Y(men_men_n1271_));
  OAI210     u1222(.A0(men_men_n1271_), .A1(men_men_n148_), .B0(men_men_n882_), .Y(men_men_n1272_));
  AOI210     u1223(.A0(men_men_n442_), .A1(men_men_n57_), .B0(men_men_n562_), .Y(men_men_n1273_));
  NA2        u1224(.A(men_men_n1273_), .B(men_men_n1272_), .Y(men_men_n1274_));
  NA3        u1225(.A(men_men_n1274_), .B(men_men_n1270_), .C(men_men_n1268_), .Y(men_men_n1275_));
  AN2        u1226(.A(x6), .B(men_men_n120_), .Y(men_men_n1276_));
  NO3        u1227(.A(men_men_n394_), .B(men_men_n340_), .C(x7), .Y(men_men_n1277_));
  NO3        u1228(.A(men_men_n150_), .B(men_men_n69_), .C(x2), .Y(men_men_n1278_));
  NO3        u1229(.A(men_men_n1278_), .B(men_men_n1277_), .C(men_men_n1276_), .Y(men_men_n1279_));
  NO2        u1230(.A(men_men_n211_), .B(x1), .Y(men_men_n1280_));
  NA2        u1231(.A(men_men_n1280_), .B(men_men_n453_), .Y(men_men_n1281_));
  NO2        u1232(.A(men_men_n57_), .B(men_men_n97_), .Y(men_men_n1282_));
  NA2        u1233(.A(men_men_n955_), .B(men_men_n1282_), .Y(men_men_n1283_));
  AOI210     u1234(.A0(men_men_n1283_), .A1(men_men_n1281_), .B0(men_men_n56_), .Y(men_men_n1284_));
  AOI220     u1235(.A0(men_men_n678_), .A1(men_men_n688_), .B0(men_men_n456_), .B1(men_men_n253_), .Y(men_men_n1285_));
  NO2        u1236(.A(men_men_n1285_), .B(men_men_n1145_), .Y(men_men_n1286_));
  NA2        u1237(.A(men_men_n825_), .B(x4), .Y(men_men_n1287_));
  OAI220     u1238(.A0(men_men_n1287_), .A1(men_men_n611_), .B0(men_men_n577_), .B1(men_men_n544_), .Y(men_men_n1288_));
  NO3        u1239(.A(men_men_n1288_), .B(men_men_n1286_), .C(men_men_n1284_), .Y(men_men_n1289_));
  OAI210     u1240(.A0(men_men_n1279_), .A1(x5), .B0(men_men_n1289_), .Y(men_men_n1290_));
  AOI220     u1241(.A0(men_men_n1290_), .A1(men_men_n88_), .B0(men_men_n1275_), .B1(men_men_n308_), .Y(men_men_n1291_));
  NA4        u1242(.A(men_men_n1291_), .B(men_men_n1264_), .C(men_men_n1244_), .D(men_men_n1229_), .Y(men17));
  NO4        u1243(.A(men_men_n536_), .B(men_men_n624_), .C(men_men_n91_), .D(men_men_n90_), .Y(men_men_n1293_));
  NO2        u1244(.A(men_men_n113_), .B(men_men_n1029_), .Y(men_men_n1294_));
  AOI220     u1245(.A0(men_men_n1294_), .A1(men_men_n639_), .B0(men_men_n1293_), .B1(men_men_n447_), .Y(men_men_n1295_));
  NA2        u1246(.A(men_men_n154_), .B(men_men_n72_), .Y(men_men_n1296_));
  NOi21      u1247(.An(men_men_n336_), .B(men_men_n76_), .Y(men_men_n1297_));
  OAI210     u1248(.A0(men_men_n554_), .A1(men_men_n55_), .B0(men_men_n1297_), .Y(men_men_n1298_));
  NA2        u1249(.A(men_men_n1073_), .B(men_men_n887_), .Y(men_men_n1299_));
  NA4        u1250(.A(men_men_n1299_), .B(men_men_n1298_), .C(men_men_n655_), .D(men_men_n57_), .Y(men_men_n1300_));
  OA210      u1251(.A0(men_men_n1156_), .A1(men_men_n1024_), .B0(men_men_n669_), .Y(men_men_n1301_));
  NA2        u1252(.A(men_men_n1301_), .B(men_men_n1300_), .Y(men_men_n1302_));
  NA3        u1253(.A(men_men_n153_), .B(men_men_n560_), .C(men_men_n927_), .Y(men_men_n1303_));
  AOI210     u1254(.A0(men_men_n952_), .A1(men_men_n278_), .B0(men_men_n59_), .Y(men_men_n1304_));
  NA2        u1255(.A(men_men_n1304_), .B(men_men_n1303_), .Y(men_men_n1305_));
  AOI210     u1256(.A0(men_men_n1302_), .A1(x1), .B0(men_men_n1305_), .Y(men_men_n1306_));
  NA2        u1257(.A(men_men_n939_), .B(men_men_n541_), .Y(men_men_n1307_));
  NO2        u1258(.A(men_men_n562_), .B(men_men_n467_), .Y(men_men_n1308_));
  OAI210     u1259(.A0(men_men_n1308_), .A1(men_men_n795_), .B0(men_men_n1246_), .Y(men_men_n1309_));
  AOI210     u1260(.A0(men_men_n1309_), .A1(men_men_n1307_), .B0(x8), .Y(men_men_n1310_));
  NA3        u1261(.A(men_men_n562_), .B(men_men_n247_), .C(men_men_n111_), .Y(men_men_n1311_));
  NO2        u1262(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n1312_));
  INV        u1263(.A(x0), .Y(men_men_n1313_));
  OAI210     u1264(.A0(men_men_n1311_), .A1(men_men_n225_), .B0(men_men_n1313_), .Y(men_men_n1314_));
  NO2        u1265(.A(men_men_n1314_), .B(men_men_n1310_), .Y(men_men_n1315_));
  OAI220     u1266(.A0(men_men_n1315_), .A1(men_men_n1306_), .B0(men_men_n1296_), .B1(men_men_n1295_), .Y(men18));
  AOI210     u1267(.A0(x8), .A1(x0), .B0(x5), .Y(men_men_n1317_));
  NA2        u1268(.A(men_men_n536_), .B(men_men_n59_), .Y(men_men_n1318_));
  AOI210     u1269(.A0(men_men_n1234_), .A1(men_men_n315_), .B0(men_men_n1318_), .Y(men_men_n1319_));
  NO4        u1270(.A(men_men_n232_), .B(men_men_n722_), .C(men_men_n144_), .D(men_men_n66_), .Y(men_men_n1320_));
  NO2        u1271(.A(men_men_n1320_), .B(men_men_n1319_), .Y(men_men_n1321_));
  NA3        u1272(.A(men_men_n462_), .B(men_men_n199_), .C(x0), .Y(men_men_n1322_));
  NAi21      u1273(.An(men_men_n341_), .B(men_men_n1322_), .Y(men_men_n1323_));
  NO2        u1274(.A(men_men_n784_), .B(x5), .Y(men_men_n1324_));
  OR2        u1275(.A(men_men_n462_), .B(men_men_n301_), .Y(men_men_n1325_));
  OAI220     u1276(.A0(men_men_n1325_), .A1(men_men_n266_), .B0(men_men_n784_), .B1(men_men_n197_), .Y(men_men_n1326_));
  AOI210     u1277(.A0(men_men_n1323_), .A1(men_men_n264_), .B0(men_men_n1326_), .Y(men_men_n1327_));
  AOI210     u1278(.A0(men_men_n1327_), .A1(men_men_n1321_), .B0(x6), .Y(men_men_n1328_));
  NA3        u1279(.A(men_men_n466_), .B(men_men_n371_), .C(x2), .Y(men_men_n1329_));
  NA3        u1280(.A(men_men_n925_), .B(men_men_n51_), .C(men_men_n57_), .Y(men_men_n1330_));
  AOI210     u1281(.A0(men_men_n1330_), .A1(men_men_n1329_), .B0(men_men_n701_), .Y(men_men_n1331_));
  AOI210     u1282(.A0(men_men_n375_), .A1(men_men_n127_), .B0(men_men_n700_), .Y(men_men_n1332_));
  NA2        u1283(.A(men_men_n244_), .B(x6), .Y(men_men_n1333_));
  OAI210     u1284(.A0(men_men_n168_), .A1(men_men_n99_), .B0(men_men_n1017_), .Y(men_men_n1334_));
  OAI220     u1285(.A0(men_men_n1334_), .A1(men_men_n1333_), .B0(men_men_n1332_), .B1(men_men_n661_), .Y(men_men_n1335_));
  OAI210     u1286(.A0(men_men_n1335_), .A1(men_men_n1331_), .B0(men_men_n53_), .Y(men_men_n1336_));
  NO2        u1287(.A(men_men_n610_), .B(men_men_n237_), .Y(men_men_n1337_));
  NO2        u1288(.A(men_men_n240_), .B(x3), .Y(men_men_n1338_));
  NO3        u1289(.A(men_men_n385_), .B(men_men_n536_), .C(men_men_n745_), .Y(men_men_n1339_));
  OAI210     u1290(.A0(men_men_n1339_), .A1(men_men_n1337_), .B0(men_men_n1338_), .Y(men_men_n1340_));
  AOI210     u1291(.A0(men_men_n1018_), .A1(men_men_n550_), .B0(x4), .Y(men_men_n1341_));
  NA2        u1292(.A(men_men_n536_), .B(men_men_n59_), .Y(men_men_n1342_));
  OAI210     u1293(.A0(men_men_n554_), .A1(men_men_n579_), .B0(men_men_n1342_), .Y(men_men_n1343_));
  AO220      u1294(.A0(men_men_n1109_), .A1(men_men_n655_), .B0(men_men_n493_), .B1(men_men_n318_), .Y(men_men_n1344_));
  AOI220     u1295(.A0(men_men_n1344_), .A1(x1), .B0(men_men_n1343_), .B1(men_men_n151_), .Y(men_men_n1345_));
  NA4        u1296(.A(men_men_n1345_), .B(men_men_n1341_), .C(men_men_n1340_), .D(men_men_n1336_), .Y(men_men_n1346_));
  NO3        u1297(.A(men_men_n946_), .B(men_men_n120_), .C(men_men_n119_), .Y(men_men_n1347_));
  NA2        u1298(.A(men_men_n1347_), .B(men_men_n97_), .Y(men_men_n1348_));
  AOI210     u1299(.A0(men_men_n1348_), .A1(men_men_n498_), .B0(men_men_n701_), .Y(men_men_n1349_));
  NA3        u1300(.A(men_men_n1065_), .B(men_men_n179_), .C(men_men_n130_), .Y(men_men_n1350_));
  NA2        u1301(.A(men_men_n160_), .B(men_men_n688_), .Y(men_men_n1351_));
  NO2        u1302(.A(men_men_n1351_), .B(men_men_n1159_), .Y(men_men_n1352_));
  AOI210     u1303(.A0(men_men_n1350_), .A1(men_men_n167_), .B0(men_men_n1352_), .Y(men_men_n1353_));
  OAI210     u1304(.A0(men_men_n1353_), .A1(men_men_n480_), .B0(x4), .Y(men_men_n1354_));
  OAI220     u1305(.A0(men_men_n1354_), .A1(men_men_n1349_), .B0(men_men_n1346_), .B1(men_men_n1328_), .Y(men_men_n1355_));
  NA2        u1306(.A(men_men_n537_), .B(men_men_n453_), .Y(men_men_n1356_));
  NO2        u1307(.A(men_men_n1356_), .B(x6), .Y(men_men_n1357_));
  NO2        u1308(.A(men_men_n340_), .B(men_men_n231_), .Y(men_men_n1358_));
  NO2        u1309(.A(men_men_n838_), .B(men_men_n520_), .Y(men_men_n1359_));
  AO220      u1310(.A0(men_men_n1359_), .A1(men_men_n57_), .B0(men_men_n1358_), .B1(men_men_n113_), .Y(men_men_n1360_));
  NO2        u1311(.A(men_men_n1360_), .B(men_men_n1357_), .Y(men_men_n1361_));
  NA2        u1312(.A(men_men_n946_), .B(x3), .Y(men_men_n1362_));
  NO2        u1313(.A(men_men_n1361_), .B(x3), .Y(men_men_n1363_));
  NO3        u1314(.A(men_men_n879_), .B(men_men_n610_), .C(men_men_n296_), .Y(men_men_n1364_));
  BUFFER     u1315(.A(men_men_n1364_), .Y(men_men_n1365_));
  AOI220     u1316(.A0(men_men_n1365_), .A1(x8), .B0(men_men_n1185_), .B1(men_men_n386_), .Y(men_men_n1366_));
  NA2        u1317(.A(men_men_n1235_), .B(men_men_n99_), .Y(men_men_n1367_));
  NO2        u1318(.A(men_men_n1366_), .B(men_men_n360_), .Y(men_men_n1368_));
  AOI210     u1319(.A0(men_men_n1363_), .A1(men_men_n127_), .B0(men_men_n1368_), .Y(men_men_n1369_));
  NA2        u1320(.A(men_men_n1369_), .B(men_men_n1355_), .Y(men19));
  NO2        u1321(.A(men_men_n1271_), .B(men_men_n235_), .Y(men_men_n1371_));
  NA2        u1322(.A(men_men_n579_), .B(x3), .Y(men_men_n1372_));
  OAI210     u1323(.A0(men_men_n144_), .A1(men_men_n98_), .B0(men_men_n73_), .Y(men_men_n1373_));
  NA3        u1324(.A(men_men_n1373_), .B(men_men_n1372_), .C(men_men_n219_), .Y(men_men_n1374_));
  NO2        u1325(.A(men_men_n1154_), .B(men_men_n160_), .Y(men_men_n1375_));
  AOI210     u1326(.A0(men_men_n1293_), .A1(men_men_n316_), .B0(men_men_n1375_), .Y(men_men_n1376_));
  AOI210     u1327(.A0(men_men_n1376_), .A1(men_men_n1374_), .B0(men_men_n56_), .Y(men_men_n1377_));
  INV        u1328(.A(men_men_n762_), .Y(men_men_n1378_));
  OAI210     u1329(.A0(men_men_n1377_), .A1(men_men_n1371_), .B0(men_men_n1378_), .Y(men_men_n1379_));
  NOi21      u1330(.An(men_men_n545_), .B(men_men_n582_), .Y(men_men_n1380_));
  AOI210     u1331(.A0(men_men_n316_), .A1(x6), .B0(men_men_n111_), .Y(men_men_n1381_));
  NO2        u1332(.A(men_men_n1381_), .B(men_men_n674_), .Y(men_men_n1382_));
  NA2        u1333(.A(men_men_n1060_), .B(men_men_n112_), .Y(men_men_n1383_));
  NO2        u1334(.A(men_men_n784_), .B(men_men_n71_), .Y(men_men_n1384_));
  NO3        u1335(.A(men_men_n1384_), .B(men_men_n1382_), .C(men_men_n902_), .Y(men_men_n1385_));
  NO2        u1336(.A(men_men_n480_), .B(men_men_n552_), .Y(men_men_n1386_));
  NA2        u1337(.A(men_men_n1105_), .B(men_men_n50_), .Y(men_men_n1387_));
  NO3        u1338(.A(men_men_n460_), .B(men_men_n280_), .C(men_men_n63_), .Y(men_men_n1388_));
  AOI220     u1339(.A0(men_men_n1388_), .A1(men_men_n1387_), .B0(men_men_n1386_), .B1(men_men_n691_), .Y(men_men_n1389_));
  OAI210     u1340(.A0(men_men_n1385_), .A1(men_men_n57_), .B0(men_men_n1389_), .Y(men_men_n1390_));
  AOI210     u1341(.A0(men_men_n1390_), .A1(men_men_n688_), .B0(men_men_n1380_), .Y(men_men_n1391_));
  NO2        u1342(.A(men_men_n98_), .B(x4), .Y(men_men_n1392_));
  INV        u1343(.A(men_men_n1231_), .Y(men_men_n1393_));
  NO2        u1344(.A(men_men_n1393_), .B(men_men_n445_), .Y(men_men_n1394_));
  OAI210     u1345(.A0(men_men_n1394_), .A1(men_men_n1392_), .B0(men_men_n722_), .Y(men_men_n1395_));
  NO2        u1346(.A(men_men_n661_), .B(men_men_n295_), .Y(men_men_n1396_));
  NO2        u1347(.A(men_men_n144_), .B(men_men_n901_), .Y(men_men_n1397_));
  AOI220     u1348(.A0(men_men_n1397_), .A1(men_men_n1117_), .B0(men_men_n1396_), .B1(men_men_n422_), .Y(men_men_n1398_));
  AO210      u1349(.A0(men_men_n1398_), .A1(men_men_n1395_), .B0(x1), .Y(men_men_n1399_));
  NA3        u1350(.A(men_men_n562_), .B(men_men_n927_), .C(men_men_n1053_), .Y(men_men_n1400_));
  NA2        u1351(.A(men_men_n137_), .B(men_men_n100_), .Y(men_men_n1401_));
  NOi21      u1352(.An(x1), .B(x6), .Y(men_men_n1402_));
  NA2        u1353(.A(men_men_n1402_), .B(men_men_n76_), .Y(men_men_n1403_));
  NA3        u1354(.A(men_men_n1403_), .B(men_men_n1401_), .C(men_men_n1400_), .Y(men_men_n1404_));
  NA2        u1355(.A(men_men_n1404_), .B(x3), .Y(men_men_n1405_));
  NA2        u1356(.A(men_men_n825_), .B(men_men_n50_), .Y(men_men_n1406_));
  NA3        u1357(.A(men_men_n1060_), .B(men_men_n338_), .C(men_men_n99_), .Y(men_men_n1407_));
  AOI210     u1358(.A0(men_men_n1407_), .A1(men_men_n1406_), .B0(men_men_n848_), .Y(men_men_n1408_));
  INV        u1359(.A(men_men_n1408_), .Y(men_men_n1409_));
  OAI210     u1360(.A0(men_men_n1405_), .A1(men_men_n751_), .B0(men_men_n1409_), .Y(men_men_n1410_));
  NO2        u1361(.A(men_men_n492_), .B(men_men_n65_), .Y(men_men_n1411_));
  OAI220     u1362(.A0(men_men_n1411_), .A1(men_men_n1372_), .B0(men_men_n279_), .B1(men_men_n792_), .Y(men_men_n1412_));
  AOI220     u1363(.A0(men_men_n1412_), .A1(men_men_n56_), .B0(men_men_n1189_), .B1(men_men_n653_), .Y(men_men_n1413_));
  NO2        u1364(.A(men_men_n54_), .B(men_men_n67_), .Y(men_men_n1414_));
  AO220      u1365(.A0(men_men_n1414_), .A1(men_men_n879_), .B0(men_men_n724_), .B1(men_men_n837_), .Y(men_men_n1415_));
  NA2        u1366(.A(men_men_n1046_), .B(men_men_n321_), .Y(men_men_n1416_));
  NO2        u1367(.A(men_men_n876_), .B(men_men_n1402_), .Y(men_men_n1417_));
  NA2        u1368(.A(men_men_n442_), .B(men_men_n653_), .Y(men_men_n1418_));
  OAI210     u1369(.A0(men_men_n1418_), .A1(men_men_n1417_), .B0(men_men_n1416_), .Y(men_men_n1419_));
  AOI210     u1370(.A0(men_men_n1415_), .A1(x2), .B0(men_men_n1419_), .Y(men_men_n1420_));
  OAI220     u1371(.A0(men_men_n1420_), .A1(men_men_n144_), .B0(men_men_n1413_), .B1(men_men_n54_), .Y(men_men_n1421_));
  OAI210     u1372(.A0(men_men_n1421_), .A1(men_men_n1410_), .B0(x8), .Y(men_men_n1422_));
  NA4        u1373(.A(men_men_n1422_), .B(men_men_n1399_), .C(men_men_n1391_), .D(men_men_n1379_), .Y(men20));
  NA2        u1374(.A(men_men_n422_), .B(men_men_n364_), .Y(men_men_n1424_));
  NO2        u1375(.A(men_men_n1424_), .B(men_men_n79_), .Y(men_men_n1425_));
  AOI210     u1376(.A0(men_men_n931_), .A1(men_men_n61_), .B0(men_men_n1386_), .Y(men_men_n1426_));
  AOI210     u1377(.A0(men_men_n870_), .A1(men_men_n314_), .B0(men_men_n1052_), .Y(men_men_n1427_));
  OAI210     u1378(.A0(men_men_n1426_), .A1(men_men_n607_), .B0(men_men_n1427_), .Y(men_men_n1428_));
  OAI210     u1379(.A0(men_men_n1428_), .A1(men_men_n1425_), .B0(men_men_n980_), .Y(men_men_n1429_));
  NAi21      u1380(.An(men_men_n489_), .B(men_men_n354_), .Y(men_men_n1430_));
  NA3        u1381(.A(men_men_n1430_), .B(men_men_n868_), .C(men_men_n837_), .Y(men_men_n1431_));
  NO2        u1382(.A(men_men_n1431_), .B(men_men_n1145_), .Y(men_men_n1432_));
  NO2        u1383(.A(men_men_n665_), .B(men_men_n858_), .Y(men_men_n1433_));
  NOi31      u1384(.An(men_men_n1433_), .B(men_men_n1039_), .C(men_men_n472_), .Y(men_men_n1434_));
  OAI210     u1385(.A0(men_men_n1434_), .A1(men_men_n1432_), .B0(men_men_n296_), .Y(men_men_n1435_));
  NO3        u1386(.A(men_men_n484_), .B(x5), .C(x2), .Y(men_men_n1436_));
  NA2        u1387(.A(men_men_n292_), .B(men_men_n84_), .Y(men_men_n1437_));
  NA2        u1388(.A(men_men_n297_), .B(men_men_n97_), .Y(men_men_n1438_));
  NA2        u1389(.A(men_men_n374_), .B(men_men_n52_), .Y(men_men_n1439_));
  OAI220     u1390(.A0(men_men_n1439_), .A1(men_men_n1438_), .B0(men_men_n1437_), .B1(men_men_n249_), .Y(men_men_n1440_));
  OAI210     u1391(.A0(men_men_n1440_), .A1(men_men_n1436_), .B0(men_men_n203_), .Y(men_men_n1441_));
  NO2        u1392(.A(men_men_n592_), .B(men_men_n541_), .Y(men_men_n1442_));
  NA2        u1393(.A(men_men_n838_), .B(men_men_n50_), .Y(men_men_n1443_));
  NO3        u1394(.A(men_men_n1443_), .B(men_men_n326_), .C(men_men_n210_), .Y(men_men_n1444_));
  NO2        u1395(.A(men_men_n1287_), .B(men_men_n914_), .Y(men_men_n1445_));
  AOI210     u1396(.A0(men_men_n1444_), .A1(men_men_n1442_), .B0(men_men_n1445_), .Y(men_men_n1446_));
  NA4        u1397(.A(men_men_n1446_), .B(men_men_n1441_), .C(men_men_n1435_), .D(men_men_n1429_), .Y(men21));
  OAI210     u1398(.A0(men_men_n357_), .A1(men_men_n54_), .B0(x7), .Y(men_men_n1448_));
  OAI220     u1399(.A0(men_men_n1448_), .A1(men_men_n1135_), .B0(men_men_n932_), .B1(men_men_n87_), .Y(men_men_n1449_));
  NA2        u1400(.A(men_men_n1449_), .B(men_men_n72_), .Y(men_men_n1450_));
  AOI210     u1401(.A0(men_men_n507_), .A1(men_men_n406_), .B0(men_men_n282_), .Y(men_men_n1451_));
  NA2        u1402(.A(men_men_n825_), .B(men_men_n248_), .Y(men_men_n1452_));
  NA2        u1403(.A(men_men_n477_), .B(men_men_n407_), .Y(men_men_n1453_));
  NA4        u1404(.A(men_men_n1453_), .B(men_men_n1452_), .C(men_men_n1212_), .D(men_men_n56_), .Y(men_men_n1454_));
  NO2        u1405(.A(men_men_n691_), .B(men_men_n385_), .Y(men_men_n1455_));
  NO3        u1406(.A(men_men_n1455_), .B(men_men_n646_), .C(men_men_n227_), .Y(men_men_n1456_));
  NO3        u1407(.A(men_men_n1456_), .B(men_men_n1454_), .C(men_men_n1451_), .Y(men_men_n1457_));
  NO3        u1408(.A(men_men_n385_), .B(men_men_n252_), .C(men_men_n52_), .Y(men_men_n1458_));
  OA210      u1409(.A0(men_men_n1458_), .A1(men_men_n782_), .B0(x3), .Y(men_men_n1459_));
  NO2        u1410(.A(men_men_n66_), .B(x2), .Y(men_men_n1460_));
  OAI210     u1411(.A0(men_men_n167_), .A1(x0), .B0(men_men_n1460_), .Y(men_men_n1461_));
  NA2        u1412(.A(men_men_n134_), .B(men_men_n97_), .Y(men_men_n1462_));
  NA2        u1413(.A(men_men_n1462_), .B(men_men_n1461_), .Y(men_men_n1463_));
  OAI210     u1414(.A0(men_men_n1463_), .A1(men_men_n1459_), .B0(x8), .Y(men_men_n1464_));
  NA2        u1415(.A(men_men_n55_), .B(men_men_n50_), .Y(men_men_n1465_));
  MUX2       u1416(.S(men_men_n536_), .A(men_men_n1465_), .B(men_men_n96_), .Y(men_men_n1466_));
  AOI210     u1417(.A0(men_men_n1194_), .A1(men_men_n218_), .B0(men_men_n1466_), .Y(men_men_n1467_));
  OAI210     u1418(.A0(men_men_n575_), .A1(men_men_n519_), .B0(x4), .Y(men_men_n1468_));
  NO2        u1419(.A(men_men_n1468_), .B(men_men_n1467_), .Y(men_men_n1469_));
  AO220      u1420(.A0(men_men_n1469_), .A1(men_men_n1464_), .B0(men_men_n1457_), .B1(men_men_n1450_), .Y(men_men_n1470_));
  AO220      u1421(.A0(men_men_n563_), .A1(men_men_n295_), .B0(men_men_n525_), .B1(x8), .Y(men_men_n1471_));
  NO2        u1422(.A(men_men_n762_), .B(x0), .Y(men_men_n1472_));
  NO3        u1423(.A(men_men_n1472_), .B(men_men_n485_), .C(men_men_n80_), .Y(men_men_n1473_));
  NO2        u1424(.A(men_men_n150_), .B(x2), .Y(men_men_n1474_));
  NO3        u1425(.A(men_men_n333_), .B(men_men_n232_), .C(men_men_n175_), .Y(men_men_n1475_));
  AOI210     u1426(.A0(men_men_n1474_), .A1(men_men_n65_), .B0(men_men_n1475_), .Y(men_men_n1476_));
  OAI210     u1427(.A0(men_men_n1473_), .A1(men_men_n353_), .B0(men_men_n1476_), .Y(men_men_n1477_));
  AOI220     u1428(.A0(men_men_n1477_), .A1(x5), .B0(men_men_n1471_), .B1(men_men_n665_), .Y(men_men_n1478_));
  AOI210     u1429(.A0(men_men_n1478_), .A1(men_men_n1470_), .B0(men_men_n67_), .Y(men_men_n1479_));
  NO2        u1430(.A(men_men_n799_), .B(men_men_n159_), .Y(men_men_n1480_));
  NOi41      u1431(.An(men_men_n1259_), .B(men_men_n1317_), .C(men_men_n1028_), .D(men_men_n755_), .Y(men_men_n1481_));
  NA2        u1432(.A(men_men_n1481_), .B(men_men_n1480_), .Y(men_men_n1482_));
  NO2        u1433(.A(men_men_n72_), .B(x4), .Y(men_men_n1483_));
  INV        u1434(.A(men_men_n1483_), .Y(men_men_n1484_));
  OAI210     u1435(.A0(men_men_n359_), .A1(men_men_n375_), .B0(men_men_n210_), .Y(men_men_n1485_));
  NO2        u1436(.A(men_men_n234_), .B(men_men_n50_), .Y(men_men_n1486_));
  NO2        u1437(.A(men_men_n1486_), .B(men_men_n57_), .Y(men_men_n1487_));
  NA2        u1438(.A(men_men_n1487_), .B(men_men_n1485_), .Y(men_men_n1488_));
  AOI210     u1439(.A0(men_men_n1484_), .A1(men_men_n1482_), .B0(men_men_n1488_), .Y(men_men_n1489_));
  NA2        u1440(.A(men_men_n271_), .B(men_men_n97_), .Y(men_men_n1490_));
  NA2        u1441(.A(men_men_n791_), .B(men_men_n55_), .Y(men_men_n1491_));
  NO2        u1442(.A(men_men_n1491_), .B(men_men_n1490_), .Y(men_men_n1492_));
  NO2        u1443(.A(men_men_n597_), .B(men_men_n935_), .Y(men_men_n1493_));
  NO3        u1444(.A(men_men_n1493_), .B(men_men_n1492_), .C(men_men_n1489_), .Y(men_men_n1494_));
  NO2        u1445(.A(men_men_n1494_), .B(x6), .Y(men_men_n1495_));
  AOI210     u1446(.A0(men_men_n544_), .A1(men_men_n935_), .B0(men_men_n1317_), .Y(men_men_n1496_));
  OAI210     u1447(.A0(men_men_n1496_), .A1(men_men_n613_), .B0(men_men_n56_), .Y(men_men_n1497_));
  NO2        u1448(.A(men_men_n667_), .B(men_men_n54_), .Y(men_men_n1498_));
  NO4        u1449(.A(men_men_n846_), .B(men_men_n252_), .C(men_men_n688_), .D(men_men_n674_), .Y(men_men_n1499_));
  NO2        u1450(.A(men_men_n766_), .B(x5), .Y(men_men_n1500_));
  NO4        u1451(.A(men_men_n1500_), .B(men_men_n1499_), .C(men_men_n1498_), .D(men_men_n831_), .Y(men_men_n1501_));
  AOI210     u1452(.A0(men_men_n1501_), .A1(men_men_n1497_), .B0(men_men_n50_), .Y(men_men_n1502_));
  NA3        u1453(.A(men_men_n55_), .B(x2), .C(x0), .Y(men_men_n1503_));
  NO2        u1454(.A(men_men_n607_), .B(men_men_n234_), .Y(men_men_n1504_));
  NO3        u1455(.A(men_men_n222_), .B(men_men_n208_), .C(men_men_n321_), .Y(men_men_n1505_));
  NO2        u1456(.A(men_men_n1505_), .B(men_men_n1504_), .Y(men_men_n1506_));
  OAI220     u1457(.A0(men_men_n1506_), .A1(men_men_n56_), .B0(men_men_n412_), .B1(men_men_n622_), .Y(men_men_n1507_));
  OAI210     u1458(.A0(men_men_n1507_), .A1(men_men_n1502_), .B0(men_men_n105_), .Y(men_men_n1508_));
  NO2        u1459(.A(men_men_n549_), .B(men_men_n277_), .Y(men_men_n1509_));
  AOI210     u1460(.A0(men_men_n542_), .A1(x5), .B0(men_men_n1509_), .Y(men_men_n1510_));
  NO2        u1461(.A(men_men_n1510_), .B(men_men_n99_), .Y(men_men_n1511_));
  NA2        u1462(.A(men_men_n630_), .B(men_men_n73_), .Y(men_men_n1512_));
  NA3        u1463(.A(men_men_n1512_), .B(men_men_n382_), .C(men_men_n57_), .Y(men_men_n1513_));
  OAI210     u1464(.A0(men_men_n1491_), .A1(men_men_n1490_), .B0(men_men_n1513_), .Y(men_men_n1514_));
  OAI210     u1465(.A0(men_men_n1514_), .A1(men_men_n1511_), .B0(x1), .Y(men_men_n1515_));
  NO4        u1466(.A(men_men_n368_), .B(men_men_n72_), .C(men_men_n138_), .D(x3), .Y(men_men_n1516_));
  NO2        u1467(.A(men_men_n297_), .B(men_men_n101_), .Y(men_men_n1517_));
  OAI210     u1468(.A0(men_men_n1516_), .A1(men_men_n1146_), .B0(men_men_n1517_), .Y(men_men_n1518_));
  NO4        u1469(.A(men_men_n1490_), .B(men_men_n846_), .C(men_men_n592_), .D(men_men_n50_), .Y(men_men_n1519_));
  INV        u1470(.A(men_men_n1519_), .Y(men_men_n1520_));
  NA4        u1471(.A(men_men_n1520_), .B(men_men_n1518_), .C(men_men_n1515_), .D(men_men_n1508_), .Y(men_men_n1521_));
  NO3        u1472(.A(men_men_n1521_), .B(men_men_n1495_), .C(men_men_n1479_), .Y(men22));
  NO3        u1473(.A(men_men_n1055_), .B(men_men_n492_), .C(men_men_n624_), .Y(men_men_n1523_));
  AOI210     u1474(.A0(x5), .A1(x2), .B0(x8), .Y(men_men_n1524_));
  NA2        u1475(.A(men_men_n1524_), .B(men_men_n59_), .Y(men_men_n1525_));
  OAI220     u1476(.A0(men_men_n1525_), .A1(men_men_n1523_), .B0(men_men_n2317_), .B1(men_men_n353_), .Y(men_men_n1526_));
  NO4        u1477(.A(men_men_n340_), .B(men_men_n201_), .C(men_men_n67_), .D(x3), .Y(men_men_n1527_));
  NO3        u1478(.A(men_men_n1100_), .B(men_men_n79_), .C(x0), .Y(men_men_n1528_));
  OAI210     u1479(.A0(men_men_n353_), .A1(men_men_n192_), .B0(x4), .Y(men_men_n1529_));
  NO3        u1480(.A(men_men_n1529_), .B(men_men_n1528_), .C(men_men_n1527_), .Y(men_men_n1530_));
  INV        u1481(.A(men_men_n1530_), .Y(men_men_n1531_));
  AOI210     u1482(.A0(men_men_n1526_), .A1(men_men_n53_), .B0(men_men_n1531_), .Y(men_men_n1532_));
  NA2        u1483(.A(men_men_n275_), .B(men_men_n280_), .Y(men_men_n1533_));
  NA3        u1484(.A(men_men_n1533_), .B(men_men_n203_), .C(men_men_n279_), .Y(men_men_n1534_));
  NA2        u1485(.A(men_men_n515_), .B(men_men_n221_), .Y(men_men_n1535_));
  NO3        u1486(.A(men_men_n442_), .B(men_men_n240_), .C(men_men_n197_), .Y(men_men_n1536_));
  NAi31      u1487(.An(men_men_n1536_), .B(men_men_n1535_), .C(men_men_n1534_), .Y(men_men_n1537_));
  NO2        u1488(.A(men_men_n412_), .B(men_men_n236_), .Y(men_men_n1538_));
  NO2        u1489(.A(men_men_n1100_), .B(x3), .Y(men_men_n1539_));
  AOI210     u1490(.A0(men_men_n1539_), .A1(men_men_n314_), .B0(men_men_n1538_), .Y(men_men_n1540_));
  OAI210     u1491(.A0(men_men_n961_), .A1(men_men_n177_), .B0(men_men_n56_), .Y(men_men_n1541_));
  NA3        u1492(.A(men_men_n55_), .B(men_men_n67_), .C(x0), .Y(men_men_n1542_));
  NO2        u1493(.A(men_men_n1542_), .B(men_men_n935_), .Y(men_men_n1543_));
  NO2        u1494(.A(men_men_n1543_), .B(men_men_n1541_), .Y(men_men_n1544_));
  OAI210     u1495(.A0(men_men_n1540_), .A1(men_men_n234_), .B0(men_men_n1544_), .Y(men_men_n1545_));
  AOI210     u1496(.A0(men_men_n1537_), .A1(men_men_n97_), .B0(men_men_n1545_), .Y(men_men_n1546_));
  AOI210     u1497(.A0(men_men_n835_), .A1(men_men_n690_), .B0(men_men_n769_), .Y(men_men_n1547_));
  OAI210     u1498(.A0(men_men_n716_), .A1(men_men_n150_), .B0(men_men_n822_), .Y(men_men_n1548_));
  OAI210     u1499(.A0(men_men_n1548_), .A1(men_men_n1547_), .B0(men_men_n548_), .Y(men_men_n1549_));
  OA210      u1500(.A0(men_men_n1546_), .A1(men_men_n1532_), .B0(men_men_n1549_), .Y(men_men_n1550_));
  OAI210     u1501(.A0(men_men_n1040_), .A1(men_men_n629_), .B0(men_men_n617_), .Y(men_men_n1551_));
  NO2        u1502(.A(men_men_n317_), .B(x0), .Y(men_men_n1552_));
  NO2        u1503(.A(men_men_n1551_), .B(men_men_n353_), .Y(men_men_n1553_));
  NO3        u1504(.A(men_men_n160_), .B(men_men_n150_), .C(men_men_n61_), .Y(men_men_n1554_));
  OAI210     u1505(.A0(men_men_n1554_), .A1(men_men_n370_), .B0(men_men_n99_), .Y(men_men_n1555_));
  NA2        u1506(.A(men_men_n130_), .B(men_men_n701_), .Y(men_men_n1556_));
  NA2        u1507(.A(men_men_n368_), .B(x3), .Y(men_men_n1557_));
  NAi31      u1508(.An(men_men_n1557_), .B(men_men_n1556_), .C(men_men_n1367_), .Y(men_men_n1558_));
  NO3        u1509(.A(men_men_n762_), .B(men_men_n411_), .C(men_men_n99_), .Y(men_men_n1559_));
  AOI210     u1510(.A0(men_men_n544_), .A1(men_men_n401_), .B0(men_men_n439_), .Y(men_men_n1560_));
  NA2        u1511(.A(men_men_n1042_), .B(x3), .Y(men_men_n1561_));
  NO2        u1512(.A(men_men_n1561_), .B(men_men_n1560_), .Y(men_men_n1562_));
  NA3        u1513(.A(men_men_n56_), .B(men_men_n50_), .C(x0), .Y(men_men_n1563_));
  NOi21      u1514(.An(men_men_n75_), .B(men_men_n655_), .Y(men_men_n1564_));
  NA2        u1515(.A(men_men_n876_), .B(men_men_n241_), .Y(men_men_n1565_));
  OAI220     u1516(.A0(men_men_n1565_), .A1(men_men_n1564_), .B0(men_men_n938_), .B1(men_men_n1563_), .Y(men_men_n1566_));
  AOI220     u1517(.A0(men_men_n1566_), .A1(men_men_n947_), .B0(men_men_n1562_), .B1(men_men_n314_), .Y(men_men_n1567_));
  NA3        u1518(.A(men_men_n1567_), .B(men_men_n1558_), .C(men_men_n1555_), .Y(men_men_n1568_));
  AOI210     u1519(.A0(men_men_n1568_), .A1(x7), .B0(men_men_n1553_), .Y(men_men_n1569_));
  OAI210     u1520(.A0(men_men_n1550_), .A1(x7), .B0(men_men_n1569_), .Y(men23));
  OR2        u1521(.A(men_men_n460_), .B(men_men_n203_), .Y(men_men_n1571_));
  AOI220     u1522(.A0(men_men_n1571_), .A1(men_men_n1433_), .B0(men_men_n550_), .B1(men_men_n267_), .Y(men_men_n1572_));
  NO3        u1523(.A(men_men_n748_), .B(men_men_n528_), .C(men_men_n433_), .Y(men_men_n1573_));
  INV        u1524(.A(men_men_n1573_), .Y(men_men_n1574_));
  OAI210     u1525(.A0(men_men_n1572_), .A1(men_men_n144_), .B0(men_men_n1574_), .Y(men_men_n1575_));
  NA2        u1526(.A(men_men_n1575_), .B(men_men_n55_), .Y(men_men_n1576_));
  NO2        u1527(.A(men_men_n846_), .B(men_men_n458_), .Y(men_men_n1577_));
  AO220      u1528(.A0(men_men_n1131_), .A1(men_men_n171_), .B0(men_men_n879_), .B1(men_men_n665_), .Y(men_men_n1578_));
  OAI210     u1529(.A0(men_men_n1578_), .A1(men_men_n1577_), .B0(men_men_n525_), .Y(men_men_n1579_));
  NA2        u1530(.A(men_men_n168_), .B(men_men_n159_), .Y(men_men_n1580_));
  NA3        u1531(.A(men_men_n57_), .B(x4), .C(x3), .Y(men_men_n1581_));
  NO3        u1532(.A(men_men_n1581_), .B(men_men_n662_), .C(men_men_n130_), .Y(men_men_n1582_));
  AOI210     u1533(.A0(men_men_n806_), .A1(men_men_n132_), .B0(men_men_n1582_), .Y(men_men_n1583_));
  NA3        u1534(.A(men_men_n1583_), .B(men_men_n1579_), .C(men_men_n1576_), .Y(men24));
  NO2        u1535(.A(men_men_n219_), .B(x1), .Y(men_men_n1585_));
  INV        u1536(.A(men_men_n308_), .Y(men_men_n1586_));
  NAi21      u1537(.An(men_men_n1585_), .B(men_men_n1586_), .Y(men_men_n1587_));
  NO2        u1538(.A(men_men_n480_), .B(men_men_n609_), .Y(men_men_n1588_));
  AOI210     u1539(.A0(men_men_n1587_), .A1(men_men_n84_), .B0(men_men_n1588_), .Y(men_men_n1589_));
  NA2        u1540(.A(men_men_n91_), .B(x8), .Y(men_men_n1590_));
  NO3        u1541(.A(men_men_n946_), .B(men_men_n1178_), .C(men_men_n927_), .Y(men_men_n1591_));
  NA2        u1542(.A(men_men_n868_), .B(men_men_n56_), .Y(men_men_n1592_));
  AO220      u1543(.A0(men_men_n1592_), .A1(men_men_n1591_), .B0(men_men_n1119_), .B1(men_men_n296_), .Y(men_men_n1593_));
  NA2        u1544(.A(men_men_n401_), .B(x8), .Y(men_men_n1594_));
  NA2        u1545(.A(men_men_n593_), .B(men_men_n113_), .Y(men_men_n1595_));
  OAI220     u1546(.A0(men_men_n1595_), .A1(men_men_n1265_), .B0(men_men_n1594_), .B1(men_men_n746_), .Y(men_men_n1596_));
  AOI220     u1547(.A0(men_men_n1596_), .A1(men_men_n1486_), .B0(men_men_n1593_), .B1(men_men_n908_), .Y(men_men_n1597_));
  OAI210     u1548(.A0(men_men_n1590_), .A1(men_men_n1589_), .B0(men_men_n1597_), .Y(men25));
  NA2        u1549(.A(men_men_n297_), .B(men_men_n59_), .Y(men_men_n1599_));
  NO2        u1550(.A(men_men_n1599_), .B(men_men_n293_), .Y(men_men_n1600_));
  OAI210     u1551(.A0(men_men_n1600_), .A1(men_men_n1047_), .B0(men_men_n105_), .Y(men_men_n1601_));
  INV        u1552(.A(men_men_n1126_), .Y(men_men_n1602_));
  NO2        u1553(.A(men_men_n661_), .B(men_men_n55_), .Y(men_men_n1603_));
  AOI220     u1554(.A0(men_men_n1603_), .A1(men_men_n1602_), .B0(men_men_n1396_), .B1(men_men_n1048_), .Y(men_men_n1604_));
  AOI210     u1555(.A0(men_men_n1604_), .A1(men_men_n1601_), .B0(men_men_n605_), .Y(men_men_n1605_));
  NO3        u1556(.A(men_men_n920_), .B(men_men_n133_), .C(men_men_n72_), .Y(men_men_n1606_));
  OAI210     u1557(.A0(men_men_n185_), .A1(men_men_n249_), .B0(men_men_n298_), .Y(men_men_n1607_));
  OAI210     u1558(.A0(men_men_n1607_), .A1(men_men_n1606_), .B0(men_men_n1046_), .Y(men_men_n1608_));
  NA2        u1559(.A(men_men_n453_), .B(men_men_n55_), .Y(men_men_n1609_));
  NO2        u1560(.A(men_men_n1609_), .B(men_men_n219_), .Y(men_men_n1610_));
  NA2        u1561(.A(men_men_n1610_), .B(men_men_n567_), .Y(men_men_n1611_));
  AOI220     u1562(.A0(men_men_n1538_), .A1(men_men_n1012_), .B0(men_men_n1312_), .B1(men_men_n334_), .Y(men_men_n1612_));
  NA3        u1563(.A(men_men_n1612_), .B(men_men_n1611_), .C(men_men_n1608_), .Y(men_men_n1613_));
  AO210      u1564(.A0(men_men_n1613_), .A1(men_men_n97_), .B0(men_men_n1605_), .Y(men26));
  NA2        u1565(.A(men_men_n688_), .B(men_men_n50_), .Y(men_men_n1615_));
  OAI220     u1566(.A0(men_men_n277_), .A1(men_men_n227_), .B0(men_men_n1615_), .B1(x7), .Y(men_men_n1616_));
  AOI220     u1567(.A0(men_men_n1616_), .A1(men_men_n84_), .B0(men_men_n1146_), .B1(men_men_n1017_), .Y(men_men_n1617_));
  NA2        u1568(.A(men_men_n555_), .B(men_men_n515_), .Y(men_men_n1618_));
  INV        u1569(.A(men_men_n665_), .Y(men_men_n1619_));
  NO2        u1570(.A(men_men_n1618_), .B(men_men_n1619_), .Y(men_men_n1620_));
  NA2        u1571(.A(men_men_n899_), .B(men_men_n520_), .Y(men_men_n1621_));
  NO2        u1572(.A(men_men_n1621_), .B(men_men_n1105_), .Y(men_men_n1622_));
  INV        u1573(.A(men_men_n1622_), .Y(men_men_n1623_));
  NA2        u1574(.A(men_men_n722_), .B(men_men_n167_), .Y(men_men_n1624_));
  NO2        u1575(.A(men_men_n1623_), .B(men_men_n53_), .Y(men_men_n1625_));
  NA2        u1576(.A(men_men_n537_), .B(men_men_n453_), .Y(men_men_n1626_));
  NO2        u1577(.A(men_men_n123_), .B(men_men_n120_), .Y(men_men_n1627_));
  NA2        u1578(.A(men_men_n1627_), .B(men_men_n111_), .Y(men_men_n1628_));
  NA2        u1579(.A(men_men_n665_), .B(x3), .Y(men_men_n1629_));
  AOI210     u1580(.A0(men_men_n1628_), .A1(men_men_n1626_), .B0(men_men_n1629_), .Y(men_men_n1630_));
  NO2        u1581(.A(men_men_n887_), .B(x3), .Y(men_men_n1631_));
  AOI210     u1582(.A0(men_men_n396_), .A1(men_men_n97_), .B0(men_men_n1631_), .Y(men_men_n1632_));
  NA3        u1583(.A(men_men_n508_), .B(men_men_n51_), .C(men_men_n56_), .Y(men_men_n1633_));
  AOI210     u1584(.A0(men_men_n1442_), .A1(men_men_n939_), .B0(x0), .Y(men_men_n1634_));
  OAI210     u1585(.A0(men_men_n1633_), .A1(men_men_n1632_), .B0(men_men_n1634_), .Y(men_men_n1635_));
  NO4        u1586(.A(men_men_n1635_), .B(men_men_n1630_), .C(men_men_n1625_), .D(men_men_n1620_), .Y(men_men_n1636_));
  AOI210     u1587(.A0(x8), .A1(x6), .B0(x5), .Y(men_men_n1637_));
  AO220      u1588(.A0(men_men_n1637_), .A1(men_men_n135_), .B0(men_men_n528_), .B1(men_men_n130_), .Y(men_men_n1638_));
  NA2        u1589(.A(men_men_n1638_), .B(men_men_n397_), .Y(men_men_n1639_));
  NO2        u1590(.A(men_men_n675_), .B(men_men_n135_), .Y(men_men_n1640_));
  NA3        u1591(.A(men_men_n1640_), .B(men_men_n1460_), .C(men_men_n124_), .Y(men_men_n1641_));
  NO2        u1592(.A(men_men_n353_), .B(men_men_n1210_), .Y(men_men_n1642_));
  OAI210     u1593(.A0(men_men_n1642_), .A1(men_men_n1182_), .B0(men_men_n396_), .Y(men_men_n1643_));
  NA3        u1594(.A(men_men_n1643_), .B(men_men_n1641_), .C(men_men_n1639_), .Y(men_men_n1644_));
  NA3        u1595(.A(men_men_n724_), .B(men_men_n887_), .C(x7), .Y(men_men_n1645_));
  AOI210     u1596(.A0(men_men_n311_), .A1(men_men_n199_), .B0(men_men_n1645_), .Y(men_men_n1646_));
  OAI220     u1597(.A0(men_men_n794_), .A1(men_men_n277_), .B0(men_men_n575_), .B1(men_men_n609_), .Y(men_men_n1647_));
  NO2        u1598(.A(men_men_n1647_), .B(men_men_n1646_), .Y(men_men_n1648_));
  NA2        u1599(.A(men_men_n593_), .B(men_men_n837_), .Y(men_men_n1649_));
  NA2        u1600(.A(men_men_n1649_), .B(men_men_n575_), .Y(men_men_n1650_));
  NA2        u1601(.A(men_men_n130_), .B(men_men_n122_), .Y(men_men_n1651_));
  OAI210     u1602(.A0(men_men_n1651_), .A1(men_men_n1254_), .B0(x0), .Y(men_men_n1652_));
  AOI210     u1603(.A0(men_men_n1650_), .A1(men_men_n1245_), .B0(men_men_n1652_), .Y(men_men_n1653_));
  OAI210     u1604(.A0(men_men_n1648_), .A1(men_men_n53_), .B0(men_men_n1653_), .Y(men_men_n1654_));
  AOI210     u1605(.A0(men_men_n1644_), .A1(x4), .B0(men_men_n1654_), .Y(men_men_n1655_));
  OA220      u1606(.A0(men_men_n1655_), .A1(men_men_n1636_), .B0(men_men_n1617_), .B1(men_men_n98_), .Y(men27));
  NA2        u1607(.A(men_men_n804_), .B(men_men_n724_), .Y(men_men_n1657_));
  NA3        u1608(.A(men_men_n730_), .B(men_men_n324_), .C(men_men_n901_), .Y(men_men_n1658_));
  AOI210     u1609(.A0(men_men_n1658_), .A1(men_men_n1657_), .B0(men_men_n199_), .Y(men_men_n1659_));
  NA2        u1610(.A(men_men_n1659_), .B(men_men_n625_), .Y(men_men_n1660_));
  XO2        u1611(.A(x8), .B(x4), .Y(men_men_n1661_));
  NO3        u1612(.A(men_men_n1661_), .B(men_men_n396_), .C(men_men_n160_), .Y(men_men_n1662_));
  OA210      u1613(.A0(men_men_n1662_), .A1(men_men_n1106_), .B0(men_men_n252_), .Y(men_men_n1663_));
  NA2        u1614(.A(men_men_n1663_), .B(men_men_n997_), .Y(men_men_n1664_));
  NO2        u1615(.A(men_men_n622_), .B(men_men_n133_), .Y(men_men_n1665_));
  NO2        u1616(.A(men_men_n1051_), .B(men_men_n234_), .Y(men_men_n1666_));
  NA2        u1617(.A(men_men_n1666_), .B(men_men_n1665_), .Y(men_men_n1667_));
  NA3        u1618(.A(men_men_n1667_), .B(men_men_n1664_), .C(men_men_n1660_), .Y(men28));
  NO2        u1619(.A(men_men_n1661_), .B(men_men_n137_), .Y(men_men_n1669_));
  OAI210     u1620(.A0(men_men_n1669_), .A1(men_men_n1121_), .B0(men_men_n520_), .Y(men_men_n1670_));
  NA3        u1621(.A(men_men_n439_), .B(men_men_n72_), .C(men_men_n541_), .Y(men_men_n1671_));
  NA2        u1622(.A(men_men_n1671_), .B(men_men_n1670_), .Y(men_men_n1672_));
  NA2        u1623(.A(men_men_n1100_), .B(men_men_n394_), .Y(men_men_n1673_));
  NA3        u1624(.A(men_men_n1673_), .B(men_men_n1236_), .C(men_men_n363_), .Y(men_men_n1674_));
  NO2        u1625(.A(men_men_n280_), .B(x4), .Y(men_men_n1675_));
  AOI220     u1626(.A0(men_men_n1675_), .A1(men_men_n1631_), .B0(men_men_n998_), .B1(men_men_n601_), .Y(men_men_n1676_));
  NA2        u1627(.A(men_men_n1676_), .B(men_men_n1674_), .Y(men_men_n1677_));
  NO2        u1628(.A(men_men_n1100_), .B(men_men_n1085_), .Y(men_men_n1678_));
  NO4        u1629(.A(x6), .B(men_men_n56_), .C(x2), .D(x0), .Y(men_men_n1679_));
  OAI210     u1630(.A0(men_men_n1679_), .A1(men_men_n1678_), .B0(men_men_n925_), .Y(men_men_n1680_));
  NA2        u1631(.A(men_men_n1042_), .B(men_men_n97_), .Y(men_men_n1681_));
  NA2        u1632(.A(men_men_n959_), .B(men_men_n96_), .Y(men_men_n1682_));
  OAI210     u1633(.A0(men_men_n1682_), .A1(men_men_n1681_), .B0(men_men_n1680_), .Y(men_men_n1683_));
  OAI210     u1634(.A0(men_men_n1683_), .A1(men_men_n1677_), .B0(x7), .Y(men_men_n1684_));
  NO2        u1635(.A(men_men_n340_), .B(x7), .Y(men_men_n1685_));
  NO3        u1636(.A(men_men_n353_), .B(men_men_n247_), .C(men_men_n112_), .Y(men_men_n1686_));
  OAI210     u1637(.A0(men_men_n769_), .A1(men_men_n236_), .B0(men_men_n73_), .Y(men_men_n1687_));
  OAI220     u1638(.A0(men_men_n1687_), .A1(men_men_n1686_), .B0(men_men_n1685_), .B1(men_men_n100_), .Y(men_men_n1688_));
  INV        u1639(.A(men_men_n583_), .Y(men_men_n1689_));
  NO2        u1640(.A(men_men_n1609_), .B(men_men_n71_), .Y(men_men_n1690_));
  AOI220     u1641(.A0(men_men_n1690_), .A1(men_men_n1689_), .B0(men_men_n423_), .B1(men_men_n50_), .Y(men_men_n1691_));
  AOI210     u1642(.A0(men_men_n1691_), .A1(men_men_n1688_), .B0(men_men_n59_), .Y(men_men_n1692_));
  AOI220     u1643(.A0(men_men_n1223_), .A1(men_men_n599_), .B0(men_men_n362_), .B1(men_men_n401_), .Y(men_men_n1693_));
  OAI210     u1644(.A0(men_men_n1693_), .A1(men_men_n133_), .B0(x1), .Y(men_men_n1694_));
  NO2        u1645(.A(men_men_n1694_), .B(men_men_n1692_), .Y(men_men_n1695_));
  AOI210     u1646(.A0(men_men_n1383_), .A1(men_men_n353_), .B0(men_men_n591_), .Y(men_men_n1696_));
  NO2        u1647(.A(men_men_n353_), .B(x5), .Y(men_men_n1697_));
  NO2        u1648(.A(men_men_n1697_), .B(men_men_n208_), .Y(men_men_n1698_));
  NO2        u1649(.A(men_men_n1698_), .B(men_men_n1696_), .Y(men_men_n1699_));
  NOi21      u1650(.An(men_men_n630_), .B(men_men_n879_), .Y(men_men_n1700_));
  NA2        u1651(.A(men_men_n1699_), .B(men_men_n997_), .Y(men_men_n1701_));
  OAI210     u1652(.A0(men_men_n394_), .A1(men_men_n51_), .B0(men_men_n895_), .Y(men_men_n1702_));
  AOI220     u1653(.A0(men_men_n1702_), .A1(men_men_n407_), .B0(men_men_n394_), .B1(men_men_n341_), .Y(men_men_n1703_));
  NO2        u1654(.A(men_men_n1703_), .B(men_men_n144_), .Y(men_men_n1704_));
  NA2        u1655(.A(men_men_n153_), .B(men_men_n67_), .Y(men_men_n1705_));
  OAI210     u1656(.A0(men_men_n1621_), .A1(men_men_n1705_), .B0(men_men_n53_), .Y(men_men_n1706_));
  OAI220     u1657(.A0(men_men_n610_), .A1(men_men_n237_), .B0(men_men_n607_), .B1(x6), .Y(men_men_n1707_));
  NO2        u1658(.A(men_men_n275_), .B(x4), .Y(men_men_n1708_));
  AOI220     u1659(.A0(men_men_n1708_), .A1(men_men_n324_), .B0(men_men_n1707_), .B1(x4), .Y(men_men_n1709_));
  NO3        u1660(.A(men_men_n1709_), .B(men_men_n295_), .C(x5), .Y(men_men_n1710_));
  NO2        u1661(.A(men_men_n630_), .B(men_men_n57_), .Y(men_men_n1711_));
  OAI210     u1662(.A0(men_men_n1711_), .A1(men_men_n1665_), .B0(men_men_n396_), .Y(men_men_n1712_));
  AOI220     u1663(.A0(men_men_n589_), .A1(men_men_n656_), .B0(men_men_n438_), .B1(men_men_n216_), .Y(men_men_n1713_));
  AOI210     u1664(.A0(men_men_n1713_), .A1(men_men_n1712_), .B0(men_men_n234_), .Y(men_men_n1714_));
  NO4        u1665(.A(men_men_n1714_), .B(men_men_n1710_), .C(men_men_n1706_), .D(men_men_n1704_), .Y(men_men_n1715_));
  AOI220     u1666(.A0(men_men_n1715_), .A1(men_men_n1701_), .B0(men_men_n1695_), .B1(men_men_n1684_), .Y(men_men_n1716_));
  AOI210     u1667(.A0(men_men_n1672_), .A1(x3), .B0(men_men_n1716_), .Y(men29));
  OAI210     u1668(.A0(men_men_n493_), .A1(men_men_n238_), .B0(men_men_n653_), .Y(men_men_n1718_));
  NA2        u1669(.A(men_men_n667_), .B(men_men_n925_), .Y(men_men_n1719_));
  AO210      u1670(.A0(men_men_n1030_), .A1(men_men_n1035_), .B0(men_men_n1719_), .Y(men_men_n1720_));
  AOI210     u1671(.A0(men_men_n172_), .A1(men_men_n157_), .B0(men_men_n630_), .Y(men_men_n1721_));
  AOI210     u1672(.A0(men_men_n1246_), .A1(men_men_n72_), .B0(men_men_n1721_), .Y(men_men_n1722_));
  NA3        u1673(.A(men_men_n1722_), .B(men_men_n1720_), .C(men_men_n1718_), .Y(men_men_n1723_));
  NO3        u1674(.A(men_men_n591_), .B(men_men_n1017_), .C(men_men_n50_), .Y(men_men_n1724_));
  NO3        u1675(.A(men_men_n1724_), .B(men_men_n1099_), .C(men_men_n493_), .Y(men_men_n1725_));
  NO2        u1676(.A(men_men_n392_), .B(men_men_n58_), .Y(men_men_n1726_));
  AOI220     u1677(.A0(men_men_n1726_), .A1(men_men_n1067_), .B0(men_men_n596_), .B1(men_men_n1209_), .Y(men_men_n1727_));
  OAI210     u1678(.A0(men_men_n1725_), .A1(men_men_n480_), .B0(men_men_n1727_), .Y(men_men_n1728_));
  AOI210     u1679(.A0(men_men_n1723_), .A1(x6), .B0(men_men_n1728_), .Y(men_men_n1729_));
  OAI210     u1680(.A0(x8), .A1(x4), .B0(x5), .Y(men_men_n1730_));
  NA2        u1681(.A(men_men_n275_), .B(men_men_n137_), .Y(men_men_n1731_));
  NA3        u1682(.A(men_men_n1731_), .B(men_men_n57_), .C(men_men_n63_), .Y(men_men_n1732_));
  NO2        u1683(.A(men_men_n1732_), .B(men_men_n784_), .Y(men_men_n1733_));
  NA2        u1684(.A(men_men_n561_), .B(men_men_n268_), .Y(men_men_n1734_));
  NO2        u1685(.A(men_men_n1734_), .B(men_men_n1067_), .Y(men_men_n1735_));
  OAI210     u1686(.A0(men_men_n791_), .A1(x8), .B0(x7), .Y(men_men_n1736_));
  NO2        u1687(.A(men_men_n1736_), .B(men_men_n116_), .Y(men_men_n1737_));
  OAI210     u1688(.A0(men_men_n1318_), .A1(men_men_n349_), .B0(men_men_n522_), .Y(men_men_n1738_));
  NO4        u1689(.A(men_men_n1738_), .B(men_men_n1737_), .C(men_men_n1735_), .D(men_men_n1733_), .Y(men_men_n1739_));
  OAI210     u1690(.A0(men_men_n1729_), .A1(x2), .B0(men_men_n1739_), .Y(men_men_n1740_));
  NA3        u1691(.A(x6), .B(men_men_n50_), .C(x2), .Y(men_men_n1741_));
  OAI210     u1692(.A0(men_men_n1085_), .A1(men_men_n316_), .B0(men_men_n1741_), .Y(men_men_n1742_));
  NO3        u1693(.A(men_men_n394_), .B(x3), .C(x0), .Y(men_men_n1743_));
  AO220      u1694(.A0(men_men_n1743_), .A1(x5), .B0(men_men_n1679_), .B1(men_men_n73_), .Y(men_men_n1744_));
  AOI210     u1695(.A0(men_men_n1742_), .A1(men_men_n311_), .B0(men_men_n1744_), .Y(men_men_n1745_));
  NO2        u1696(.A(men_men_n1745_), .B(x7), .Y(men_men_n1746_));
  NO2        u1697(.A(men_men_n137_), .B(x2), .Y(men_men_n1747_));
  OA210      u1698(.A0(men_men_n1747_), .A1(men_men_n559_), .B0(men_men_n591_), .Y(men_men_n1748_));
  NA2        u1699(.A(men_men_n1748_), .B(men_men_n65_), .Y(men_men_n1749_));
  NA3        u1700(.A(men_men_n1697_), .B(men_men_n211_), .C(men_men_n75_), .Y(men_men_n1750_));
  NA2        u1701(.A(men_men_n1750_), .B(men_men_n1749_), .Y(men_men_n1751_));
  AOI210     u1702(.A0(men_men_n1746_), .A1(x8), .B0(men_men_n1751_), .Y(men_men_n1752_));
  NA2        u1703(.A(men_men_n2323_), .B(men_men_n50_), .Y(men_men_n1753_));
  NO2        u1704(.A(men_men_n124_), .B(men_men_n84_), .Y(men_men_n1754_));
  AOI220     u1705(.A0(men_men_n1754_), .A1(men_men_n523_), .B0(men_men_n1678_), .B1(men_men_n321_), .Y(men_men_n1755_));
  NOi31      u1706(.An(men_men_n999_), .B(men_men_n1637_), .C(men_men_n554_), .Y(men_men_n1756_));
  NA2        u1707(.A(men_men_n162_), .B(x4), .Y(men_men_n1757_));
  NO3        u1708(.A(men_men_n1297_), .B(men_men_n219_), .C(men_men_n67_), .Y(men_men_n1758_));
  AOI210     u1709(.A0(men_men_n1758_), .A1(men_men_n1757_), .B0(men_men_n1756_), .Y(men_men_n1759_));
  NA3        u1710(.A(men_men_n1759_), .B(men_men_n1755_), .C(men_men_n1753_), .Y(men_men_n1760_));
  NO4        u1711(.A(men_men_n1085_), .B(men_men_n160_), .C(men_men_n55_), .D(men_men_n67_), .Y(men_men_n1761_));
  NO4        u1712(.A(men_men_n1060_), .B(men_men_n445_), .C(men_men_n1209_), .D(men_men_n97_), .Y(men_men_n1762_));
  OAI210     u1713(.A0(men_men_n1762_), .A1(men_men_n1761_), .B0(men_men_n99_), .Y(men_men_n1763_));
  AOI210     u1714(.A0(men_men_n279_), .A1(x4), .B0(men_men_n181_), .Y(men_men_n1764_));
  OAI210     u1715(.A0(men_men_n1764_), .A1(men_men_n1726_), .B0(men_men_n648_), .Y(men_men_n1765_));
  NA2        u1716(.A(men_men_n1679_), .B(men_men_n721_), .Y(men_men_n1766_));
  OA220      u1717(.A0(men_men_n1766_), .A1(men_men_n223_), .B0(men_men_n516_), .B1(men_men_n1563_), .Y(men_men_n1767_));
  NA3        u1718(.A(men_men_n1767_), .B(men_men_n1765_), .C(men_men_n1763_), .Y(men_men_n1768_));
  AOI210     u1719(.A0(men_men_n1760_), .A1(men_men_n264_), .B0(men_men_n1768_), .Y(men_men_n1769_));
  OAI210     u1720(.A0(men_men_n1752_), .A1(x1), .B0(men_men_n1769_), .Y(men_men_n1770_));
  AO210      u1721(.A0(men_men_n1740_), .A1(x1), .B0(men_men_n1770_), .Y(men30));
  NO3        u1722(.A(men_men_n1552_), .B(men_men_n512_), .C(men_men_n88_), .Y(men_men_n1772_));
  AOI210     u1723(.A0(men_men_n338_), .A1(men_men_n1772_), .B0(men_men_n56_), .Y(men_men_n1773_));
  NA2        u1724(.A(men_men_n724_), .B(men_men_n309_), .Y(men_men_n1774_));
  NA2        u1725(.A(men_men_n1774_), .B(men_men_n1196_), .Y(men_men_n1775_));
  OAI210     u1726(.A0(men_men_n1775_), .A1(men_men_n1773_), .B0(men_men_n99_), .Y(men_men_n1776_));
  NO3        u1727(.A(men_men_n254_), .B(men_men_n111_), .C(x0), .Y(men_men_n1777_));
  AOI210     u1728(.A0(men_men_n447_), .A1(x6), .B0(men_men_n1777_), .Y(men_men_n1778_));
  AOI220     u1729(.A0(men_men_n1012_), .A1(men_men_n374_), .B0(men_men_n678_), .B1(men_men_n83_), .Y(men_men_n1779_));
  OAI220     u1730(.A0(men_men_n1779_), .A1(men_men_n223_), .B0(men_men_n1778_), .B1(men_men_n54_), .Y(men_men_n1780_));
  AO210      u1731(.A0(men_men_n507_), .A1(men_men_n461_), .B0(x5), .Y(men_men_n1781_));
  NO2        u1732(.A(men_men_n645_), .B(men_men_n1781_), .Y(men_men_n1782_));
  AOI210     u1733(.A0(men_men_n1402_), .A1(men_men_n50_), .B0(men_men_n401_), .Y(men_men_n1783_));
  OAI210     u1734(.A0(x7), .A1(x6), .B0(x1), .Y(men_men_n1784_));
  NA3        u1735(.A(men_men_n57_), .B(x4), .C(men_men_n59_), .Y(men_men_n1785_));
  AOI220     u1736(.A0(men_men_n1785_), .A1(men_men_n1201_), .B0(men_men_n1784_), .B1(men_men_n1581_), .Y(men_men_n1786_));
  NO2        u1737(.A(men_men_n459_), .B(men_men_n764_), .Y(men_men_n1787_));
  NOi21      u1738(.An(men_men_n1787_), .B(men_men_n751_), .Y(men_men_n1788_));
  NO3        u1739(.A(men_men_n1145_), .B(men_men_n212_), .C(men_men_n579_), .Y(men_men_n1789_));
  NO3        u1740(.A(men_men_n1789_), .B(men_men_n1788_), .C(men_men_n1786_), .Y(men_men_n1790_));
  OAI210     u1741(.A0(men_men_n2314_), .A1(men_men_n674_), .B0(men_men_n1790_), .Y(men_men_n1791_));
  NO3        u1742(.A(men_men_n1791_), .B(men_men_n1782_), .C(men_men_n1780_), .Y(men_men_n1792_));
  AOI210     u1743(.A0(men_men_n1792_), .A1(men_men_n1776_), .B0(x8), .Y(men_men_n1793_));
  NA2        u1744(.A(men_men_n966_), .B(men_men_n59_), .Y(men_men_n1794_));
  AOI210     u1745(.A0(men_men_n807_), .A1(men_men_n437_), .B0(men_men_n606_), .Y(men_men_n1795_));
  OAI220     u1746(.A0(men_men_n1795_), .A1(men_men_n279_), .B0(men_men_n1794_), .B1(men_men_n428_), .Y(men_men_n1796_));
  AOI210     u1747(.A0(men_men_n477_), .A1(x8), .B0(men_men_n1796_), .Y(men_men_n1797_));
  NO2        u1748(.A(men_men_n1797_), .B(men_men_n57_), .Y(men_men_n1798_));
  NO2        u1749(.A(men_men_n806_), .B(men_men_n587_), .Y(men_men_n1799_));
  AOI210     u1750(.A0(men_men_n1799_), .A1(men_men_n2311_), .B0(men_men_n394_), .Y(men_men_n1800_));
  NO3        u1751(.A(men_men_n567_), .B(men_men_n359_), .C(men_men_n1016_), .Y(men_men_n1801_));
  NO3        u1752(.A(men_men_n1801_), .B(men_men_n1105_), .C(men_men_n1209_), .Y(men_men_n1802_));
  AOI210     u1753(.A0(men_men_n276_), .A1(x1), .B0(men_men_n138_), .Y(men_men_n1803_));
  NO2        u1754(.A(men_men_n282_), .B(x5), .Y(men_men_n1804_));
  NO2        u1755(.A(men_men_n1804_), .B(men_men_n758_), .Y(men_men_n1805_));
  OAI220     u1756(.A0(men_men_n1805_), .A1(men_men_n936_), .B0(men_men_n1803_), .B1(men_men_n193_), .Y(men_men_n1806_));
  NO3        u1757(.A(men_men_n1806_), .B(men_men_n1802_), .C(men_men_n1800_), .Y(men_men_n1807_));
  NA2        u1758(.A(men_men_n846_), .B(men_men_n74_), .Y(men_men_n1808_));
  AO210      u1759(.A0(men_men_n1808_), .A1(men_men_n1403_), .B0(x3), .Y(men_men_n1809_));
  NO2        u1760(.A(men_men_n200_), .B(men_men_n56_), .Y(men_men_n1810_));
  OAI220     u1761(.A0(men_men_n333_), .A1(men_men_n1105_), .B0(men_men_n317_), .B1(men_men_n212_), .Y(men_men_n1811_));
  AOI220     u1762(.A0(men_men_n1811_), .A1(x2), .B0(men_men_n1810_), .B1(men_men_n1414_), .Y(men_men_n1812_));
  AOI210     u1763(.A0(men_men_n1812_), .A1(men_men_n1809_), .B0(men_men_n237_), .Y(men_men_n1813_));
  NO2        u1764(.A(men_men_n276_), .B(men_men_n112_), .Y(men_men_n1814_));
  NO3        u1765(.A(men_men_n729_), .B(men_men_n624_), .C(men_men_n157_), .Y(men_men_n1815_));
  OAI210     u1766(.A0(men_men_n1815_), .A1(men_men_n1814_), .B0(men_men_n145_), .Y(men_men_n1816_));
  NA3        u1767(.A(x5), .B(x4), .C(men_men_n59_), .Y(men_men_n1817_));
  NO2        u1768(.A(men_men_n1153_), .B(men_men_n478_), .Y(men_men_n1818_));
  AOI210     u1769(.A0(men_men_n1170_), .A1(x2), .B0(men_men_n1818_), .Y(men_men_n1819_));
  AOI210     u1770(.A0(men_men_n1819_), .A1(men_men_n1816_), .B0(men_men_n50_), .Y(men_men_n1820_));
  NA3        u1771(.A(men_men_n1294_), .B(men_men_n1007_), .C(men_men_n421_), .Y(men_men_n1821_));
  AOI210     u1772(.A0(men_men_n1821_), .A1(men_men_n1808_), .B0(men_men_n544_), .Y(men_men_n1822_));
  AOI210     u1773(.A0(men_men_n901_), .A1(x1), .B0(men_men_n1163_), .Y(men_men_n1823_));
  OAI220     u1774(.A0(men_men_n280_), .A1(x4), .B0(men_men_n51_), .B1(x6), .Y(men_men_n1824_));
  NO2        u1775(.A(men_men_n111_), .B(men_men_n101_), .Y(men_men_n1825_));
  AOI220     u1776(.A0(men_men_n1825_), .A1(men_men_n1824_), .B0(men_men_n1031_), .B1(men_men_n554_), .Y(men_men_n1826_));
  OAI210     u1777(.A0(men_men_n1823_), .A1(men_men_n432_), .B0(men_men_n1826_), .Y(men_men_n1827_));
  NO4        u1778(.A(men_men_n1827_), .B(men_men_n1822_), .C(men_men_n1820_), .D(men_men_n1813_), .Y(men_men_n1828_));
  OAI210     u1779(.A0(men_men_n1807_), .A1(men_men_n124_), .B0(men_men_n1828_), .Y(men_men_n1829_));
  NO3        u1780(.A(men_men_n1829_), .B(men_men_n1798_), .C(men_men_n1793_), .Y(men31));
  NA2        u1781(.A(men_men_n868_), .B(men_men_n318_), .Y(men_men_n1831_));
  AOI210     u1782(.A0(men_men_n2322_), .A1(men_men_n1831_), .B0(men_men_n58_), .Y(men_men_n1832_));
  NO2        u1783(.A(men_men_n701_), .B(men_men_n56_), .Y(men_men_n1833_));
  OAI210     u1784(.A0(men_men_n82_), .A1(men_men_n1832_), .B0(men_men_n53_), .Y(men_men_n1834_));
  OA220      u1785(.A0(men_men_n275_), .A1(men_men_n421_), .B0(men_men_n59_), .B1(men_men_n1287_), .Y(men_men_n1835_));
  AOI210     u1786(.A0(men_men_n1835_), .A1(men_men_n1834_), .B0(men_men_n97_), .Y(men_men_n1836_));
  NA2        u1787(.A(men_men_n394_), .B(men_men_n57_), .Y(men_men_n1837_));
  AOI210     u1788(.A0(men_men_n279_), .A1(men_men_n78_), .B0(men_men_n1837_), .Y(men_men_n1838_));
  NA2        u1789(.A(men_men_n1838_), .B(men_men_n688_), .Y(men_men_n1839_));
  NO4        u1790(.A(men_men_n1028_), .B(men_men_n325_), .C(men_men_n1402_), .D(men_men_n64_), .Y(men_men_n1840_));
  OAI210     u1791(.A0(men_men_n1154_), .A1(men_men_n838_), .B0(men_men_n690_), .Y(men_men_n1841_));
  NO2        u1792(.A(men_men_n1841_), .B(men_men_n1840_), .Y(men_men_n1842_));
  AOI210     u1793(.A0(men_men_n1842_), .A1(men_men_n1839_), .B0(x5), .Y(men_men_n1843_));
  AOI220     u1794(.A0(men_men_n396_), .A1(men_men_n554_), .B0(men_men_n508_), .B1(men_men_n62_), .Y(men_men_n1844_));
  AOI210     u1795(.A0(men_men_n1844_), .A1(men_men_n516_), .B0(men_men_n1085_), .Y(men_men_n1845_));
  AOI220     u1796(.A0(men_men_n847_), .A1(men_men_n656_), .B0(men_men_n1016_), .B1(men_men_n110_), .Y(men_men_n1846_));
  OAI220     u1797(.A0(men_men_n1846_), .A1(men_men_n340_), .B0(men_men_n428_), .B1(men_men_n689_), .Y(men_men_n1847_));
  NO4        u1798(.A(men_men_n1847_), .B(men_men_n1845_), .C(men_men_n1843_), .D(men_men_n1836_), .Y(men_men_n1848_));
  NA2        u1799(.A(men_men_n437_), .B(men_men_n59_), .Y(men_men_n1849_));
  OAI210     u1800(.A0(men_men_n93_), .A1(men_men_n249_), .B0(men_men_n1794_), .Y(men_men_n1850_));
  NA2        u1801(.A(men_men_n1850_), .B(x7), .Y(men_men_n1851_));
  NA2        u1802(.A(men_men_n963_), .B(men_men_n83_), .Y(men_men_n1852_));
  AOI210     u1803(.A0(men_men_n794_), .A1(men_men_n101_), .B0(men_men_n1852_), .Y(men_men_n1853_));
  NA2        u1804(.A(men_men_n1358_), .B(x6), .Y(men_men_n1854_));
  AOI210     u1805(.A0(men_men_n1854_), .A1(men_men_n263_), .B0(men_men_n97_), .Y(men_men_n1855_));
  NA2        u1806(.A(men_men_n1048_), .B(men_men_n292_), .Y(men_men_n1856_));
  AOI210     u1807(.A0(men_men_n1856_), .A1(men_men_n575_), .B0(men_men_n53_), .Y(men_men_n1857_));
  NO3        u1808(.A(men_men_n1857_), .B(men_men_n1855_), .C(men_men_n1853_), .Y(men_men_n1858_));
  AOI210     u1809(.A0(men_men_n1858_), .A1(men_men_n1851_), .B0(men_men_n609_), .Y(men_men_n1859_));
  NOi21      u1810(.An(men_men_n1542_), .B(men_men_n940_), .Y(men_men_n1860_));
  OAI220     u1811(.A0(men_men_n1860_), .A1(men_men_n1681_), .B0(men_men_n808_), .B1(men_men_n1849_), .Y(men_men_n1861_));
  NA2        u1812(.A(men_men_n1861_), .B(x3), .Y(men_men_n1862_));
  AOI210     u1813(.A0(men_men_n1218_), .A1(x8), .B0(x1), .Y(men_men_n1863_));
  NO3        u1814(.A(men_men_n1863_), .B(men_men_n987_), .C(x6), .Y(men_men_n1864_));
  AOI220     u1815(.A0(men_men_n548_), .A1(men_men_n359_), .B0(men_men_n437_), .B1(men_men_n72_), .Y(men_men_n1865_));
  NA2        u1816(.A(men_men_n106_), .B(men_men_n472_), .Y(men_men_n1866_));
  OAI220     u1817(.A0(men_men_n1866_), .A1(men_men_n1681_), .B0(men_men_n1865_), .B1(x4), .Y(men_men_n1867_));
  NO2        u1818(.A(men_men_n1867_), .B(men_men_n1864_), .Y(men_men_n1868_));
  AOI210     u1819(.A0(men_men_n1868_), .A1(men_men_n1862_), .B0(men_men_n175_), .Y(men_men_n1869_));
  NA2        u1820(.A(men_men_n955_), .B(x3), .Y(men_men_n1870_));
  NO4        u1821(.A(men_men_n717_), .B(men_men_n1085_), .C(men_men_n688_), .D(x5), .Y(men_men_n1871_));
  INV        u1822(.A(men_men_n1871_), .Y(men_men_n1872_));
  AOI210     u1823(.A0(men_men_n1872_), .A1(men_men_n1870_), .B0(men_men_n475_), .Y(men_men_n1873_));
  OAI210     u1824(.A0(men_men_n548_), .A1(men_men_n415_), .B0(men_men_n825_), .Y(men_men_n1874_));
  NO3        u1825(.A(men_men_n407_), .B(men_men_n314_), .C(men_men_n50_), .Y(men_men_n1875_));
  NA2        u1826(.A(men_men_n1875_), .B(men_men_n1029_), .Y(men_men_n1876_));
  AOI210     u1827(.A0(men_men_n1876_), .A1(men_men_n1874_), .B0(men_men_n347_), .Y(men_men_n1877_));
  NO2        u1828(.A(men_men_n199_), .B(men_men_n478_), .Y(men_men_n1878_));
  OAI210     u1829(.A0(men_men_n127_), .A1(x2), .B0(men_men_n1878_), .Y(men_men_n1879_));
  NA3        u1830(.A(men_men_n359_), .B(men_men_n297_), .C(men_men_n71_), .Y(men_men_n1880_));
  OA210      u1831(.A0(men_men_n222_), .A1(men_men_n209_), .B0(men_men_n1880_), .Y(men_men_n1881_));
  AOI210     u1832(.A0(men_men_n1881_), .A1(men_men_n1879_), .B0(men_men_n63_), .Y(men_men_n1882_));
  NA2        u1833(.A(men_men_n111_), .B(men_men_n57_), .Y(men_men_n1883_));
  AOI220     u1834(.A0(men_men_n1383_), .A1(men_men_n799_), .B0(men_men_n248_), .B1(x4), .Y(men_men_n1884_));
  AOI220     u1835(.A0(men_men_n1430_), .A1(men_men_n550_), .B0(men_men_n646_), .B1(men_men_n688_), .Y(men_men_n1885_));
  OAI220     u1836(.A0(men_men_n1885_), .A1(men_men_n1883_), .B0(men_men_n1884_), .B1(men_men_n179_), .Y(men_men_n1886_));
  OR3        u1837(.A(men_men_n1886_), .B(men_men_n1882_), .C(men_men_n1877_), .Y(men_men_n1887_));
  NO4        u1838(.A(men_men_n1887_), .B(men_men_n1873_), .C(men_men_n1869_), .D(men_men_n1859_), .Y(men_men_n1888_));
  OAI210     u1839(.A0(men_men_n1848_), .A1(x3), .B0(men_men_n1888_), .Y(men32));
  OAI210     u1840(.A0(men_men_n501_), .A1(men_men_n53_), .B0(men_men_n364_), .Y(men_men_n1890_));
  NA2        u1841(.A(men_men_n456_), .B(x2), .Y(men_men_n1891_));
  AOI210     u1842(.A0(men_men_n1891_), .A1(men_men_n1890_), .B0(men_men_n57_), .Y(men_men_n1892_));
  OAI210     u1843(.A0(men_men_n1892_), .A1(men_men_n702_), .B0(men_men_n56_), .Y(men_men_n1893_));
  NO2        u1844(.A(men_men_n1491_), .B(men_men_n1271_), .Y(men_men_n1894_));
  AOI210     u1845(.A0(men_men_n1833_), .A1(men_men_n252_), .B0(men_men_n1894_), .Y(men_men_n1895_));
  AOI210     u1846(.A0(men_men_n1895_), .A1(men_men_n1893_), .B0(men_men_n50_), .Y(men_men_n1896_));
  NA3        u1847(.A(men_men_n57_), .B(men_men_n715_), .C(men_men_n262_), .Y(men_men_n1897_));
  INV        u1848(.A(men_men_n484_), .Y(men_men_n1898_));
  OAI220     u1849(.A0(men_men_n935_), .A1(men_men_n211_), .B0(men_men_n607_), .B1(men_men_n193_), .Y(men_men_n1899_));
  NO3        u1850(.A(men_men_n329_), .B(men_men_n509_), .C(men_men_n721_), .Y(men_men_n1900_));
  NO3        u1851(.A(men_men_n1900_), .B(men_men_n1899_), .C(men_men_n1898_), .Y(men_men_n1901_));
  AOI210     u1852(.A0(men_men_n1901_), .A1(men_men_n1897_), .B0(men_men_n131_), .Y(men_men_n1902_));
  NA2        u1853(.A(x0), .B(men_men_n846_), .Y(men_men_n1903_));
  NO2        u1854(.A(men_men_n489_), .B(men_men_n764_), .Y(men_men_n1904_));
  NA2        u1855(.A(men_men_n1904_), .B(men_men_n1640_), .Y(men_men_n1905_));
  AOI210     u1856(.A0(men_men_n1905_), .A1(men_men_n1903_), .B0(men_men_n99_), .Y(men_men_n1906_));
  AOI220     u1857(.A0(men_men_n1189_), .A1(men_men_n625_), .B0(men_men_n1093_), .B1(men_men_n923_), .Y(men_men_n1907_));
  NO2        u1858(.A(men_men_n1907_), .B(men_men_n56_), .Y(men_men_n1908_));
  NA2        u1859(.A(men_men_n846_), .B(men_men_n57_), .Y(men_men_n1909_));
  NOi21      u1860(.An(men_men_n1909_), .B(men_men_n120_), .Y(men_men_n1910_));
  NA2        u1861(.A(men_men_n891_), .B(men_men_n227_), .Y(men_men_n1911_));
  NO3        u1862(.A(men_men_n1911_), .B(men_men_n1910_), .C(men_men_n59_), .Y(men_men_n1912_));
  OR4        u1863(.A(men_men_n1912_), .B(men_men_n1908_), .C(men_men_n1906_), .D(men_men_n1902_), .Y(men_men_n1913_));
  OAI210     u1864(.A0(men_men_n1913_), .A1(men_men_n1896_), .B0(men_men_n97_), .Y(men_men_n1914_));
  NO3        u1865(.A(men_men_n1085_), .B(men_men_n135_), .C(men_men_n113_), .Y(men_men_n1915_));
  OAI210     u1866(.A0(men_men_n563_), .A1(men_men_n525_), .B0(men_men_n724_), .Y(men_men_n1916_));
  INV        u1867(.A(men_men_n1916_), .Y(men_men_n1917_));
  OAI210     u1868(.A0(men_men_n1917_), .A1(men_men_n1915_), .B0(x3), .Y(men_men_n1918_));
  NO3        u1869(.A(men_men_n277_), .B(men_men_n162_), .C(men_men_n112_), .Y(men_men_n1919_));
  NO3        u1870(.A(men_men_n715_), .B(men_men_n323_), .C(men_men_n131_), .Y(men_men_n1920_));
  OAI210     u1871(.A0(men_men_n1920_), .A1(men_men_n1919_), .B0(men_men_n59_), .Y(men_men_n1921_));
  NA2        u1872(.A(men_men_n1019_), .B(men_men_n67_), .Y(men_men_n1922_));
  NO2        u1873(.A(men_men_n1685_), .B(men_men_n525_), .Y(men_men_n1923_));
  AOI210     u1874(.A0(men_men_n1923_), .A1(men_men_n1624_), .B0(men_men_n1922_), .Y(men_men_n1924_));
  NO2        u1875(.A(men_men_n249_), .B(men_men_n57_), .Y(men_men_n1925_));
  NO2        u1876(.A(men_men_n1925_), .B(men_men_n884_), .Y(men_men_n1926_));
  NOi31      u1877(.An(men_men_n648_), .B(men_men_n1926_), .C(men_men_n254_), .Y(men_men_n1927_));
  NO3        u1878(.A(men_men_n1156_), .B(men_men_n199_), .C(men_men_n234_), .Y(men_men_n1928_));
  NO4        u1879(.A(men_men_n1928_), .B(men_men_n1927_), .C(men_men_n1924_), .D(x1), .Y(men_men_n1929_));
  NA3        u1880(.A(men_men_n1929_), .B(men_men_n1921_), .C(men_men_n1918_), .Y(men_men_n1930_));
  NA4        u1881(.A(men_men_n1112_), .B(men_men_n470_), .C(men_men_n340_), .D(men_men_n211_), .Y(men_men_n1931_));
  NO2        u1882(.A(men_men_n1599_), .B(men_men_n63_), .Y(men_men_n1932_));
  NO2        u1883(.A(men_men_n1932_), .B(men_men_n53_), .Y(men_men_n1933_));
  NO3        u1884(.A(men_men_n411_), .B(men_men_n963_), .C(men_men_n111_), .Y(men_men_n1934_));
  NO2        u1885(.A(men_men_n609_), .B(men_men_n162_), .Y(men_men_n1935_));
  OAI210     u1886(.A0(men_men_n1935_), .A1(men_men_n1934_), .B0(men_men_n65_), .Y(men_men_n1936_));
  NO2        u1887(.A(men_men_n1730_), .B(men_men_n326_), .Y(men_men_n1937_));
  OAI210     u1888(.A0(men_men_n1627_), .A1(men_men_n542_), .B0(men_men_n1937_), .Y(men_men_n1938_));
  NA4        u1889(.A(men_men_n1938_), .B(men_men_n1936_), .C(men_men_n1933_), .D(men_men_n1931_), .Y(men_men_n1939_));
  NA2        u1890(.A(men_men_n1939_), .B(men_men_n1930_), .Y(men_men_n1940_));
  NO3        u1891(.A(men_men_n1073_), .B(men_men_n96_), .C(men_men_n67_), .Y(men_men_n1941_));
  NO2        u1892(.A(men_men_n501_), .B(men_men_n327_), .Y(men_men_n1942_));
  OAI210     u1893(.A0(men_men_n1941_), .A1(men_men_n1241_), .B0(men_men_n1942_), .Y(men_men_n1943_));
  NO3        u1894(.A(x8), .B(men_men_n67_), .C(x2), .Y(men_men_n1944_));
  OAI220     u1895(.A0(men_men_n1944_), .A1(men_men_n554_), .B0(men_men_n1246_), .B1(men_men_n82_), .Y(men_men_n1945_));
  AOI220     u1896(.A0(men_men_n493_), .A1(men_men_n724_), .B0(men_men_n601_), .B1(men_men_n232_), .Y(men_men_n1946_));
  AOI210     u1897(.A0(men_men_n1946_), .A1(men_men_n1945_), .B0(men_men_n240_), .Y(men_men_n1947_));
  NA2        u1898(.A(men_men_n891_), .B(men_men_n1016_), .Y(men_men_n1948_));
  AOI210     u1899(.A0(men_men_n597_), .A1(men_men_n609_), .B0(men_men_n1948_), .Y(men_men_n1949_));
  AOI210     u1900(.A0(men_men_n523_), .A1(men_men_n554_), .B0(men_men_n615_), .Y(men_men_n1950_));
  NO2        u1901(.A(men_men_n1950_), .B(men_men_n1581_), .Y(men_men_n1951_));
  NO3        u1902(.A(men_men_n1951_), .B(men_men_n1949_), .C(men_men_n1947_), .Y(men_men_n1952_));
  NA4        u1903(.A(men_men_n1952_), .B(men_men_n1943_), .C(men_men_n1940_), .D(men_men_n1914_), .Y(men33));
  OAI210     u1904(.A0(men_men_n2320_), .A1(x1), .B0(men_men_n188_), .Y(men_men_n1954_));
  OAI220     u1905(.A0(men_men_n950_), .A1(men_men_n721_), .B0(men_men_n1460_), .B1(men_men_n316_), .Y(men_men_n1955_));
  NA2        u1906(.A(men_men_n1955_), .B(men_men_n566_), .Y(men_men_n1956_));
  AOI210     u1907(.A0(men_men_n1954_), .A1(x5), .B0(men_men_n1956_), .Y(men_men_n1957_));
  OAI210     u1908(.A0(men_men_n385_), .A1(men_men_n244_), .B0(men_men_n53_), .Y(men_men_n1958_));
  AOI210     u1909(.A0(men_men_n1958_), .A1(men_men_n387_), .B0(men_men_n63_), .Y(men_men_n1959_));
  NO2        u1910(.A(x6), .B(men_men_n1959_), .Y(men_men_n1960_));
  OAI210     u1911(.A0(men_men_n1957_), .A1(x4), .B0(men_men_n1960_), .Y(men_men_n1961_));
  OAI210     u1912(.A0(men_men_n133_), .A1(x5), .B0(men_men_n218_), .Y(men_men_n1962_));
  NA2        u1913(.A(men_men_n175_), .B(x4), .Y(men_men_n1963_));
  NA2        u1914(.A(men_men_n282_), .B(men_men_n259_), .Y(men_men_n1964_));
  NO2        u1915(.A(men_men_n846_), .B(men_men_n208_), .Y(men_men_n1965_));
  OAI220     u1916(.A0(men_men_n2321_), .A1(men_men_n1965_), .B0(men_men_n1964_), .B1(men_men_n1963_), .Y(men_men_n1966_));
  AOI210     u1917(.A0(men_men_n1962_), .A1(men_men_n899_), .B0(men_men_n1966_), .Y(men_men_n1967_));
  NA2        u1918(.A(men_men_n196_), .B(men_men_n837_), .Y(men_men_n1968_));
  AOI210     u1919(.A0(men_men_n1968_), .A1(men_men_n1909_), .B0(men_men_n197_), .Y(men_men_n1969_));
  NO2        u1920(.A(men_men_n1438_), .B(men_men_n838_), .Y(men_men_n1970_));
  OAI210     u1921(.A0(men_men_n764_), .A1(men_men_n51_), .B0(x6), .Y(men_men_n1971_));
  NO2        u1922(.A(men_men_n551_), .B(men_men_n447_), .Y(men_men_n1972_));
  NO4        u1923(.A(men_men_n1972_), .B(men_men_n1971_), .C(men_men_n1970_), .D(men_men_n1969_), .Y(men_men_n1973_));
  OAI210     u1924(.A0(men_men_n1967_), .A1(men_men_n50_), .B0(men_men_n1973_), .Y(men_men_n1974_));
  NA3        u1925(.A(men_men_n1974_), .B(men_men_n1961_), .C(men_men_n59_), .Y(men_men_n1975_));
  NO2        u1926(.A(men_men_n1367_), .B(x4), .Y(men_men_n1976_));
  NO2        u1927(.A(men_men_n1976_), .B(men_men_n388_), .Y(men_men_n1977_));
  NA2        u1928(.A(men_men_n722_), .B(men_men_n97_), .Y(men_men_n1978_));
  NA2        u1929(.A(men_men_n1978_), .B(men_men_n406_), .Y(men_men_n1979_));
  NO2        u1930(.A(men_men_n630_), .B(men_men_n329_), .Y(men_men_n1980_));
  NA2        u1931(.A(men_men_n444_), .B(men_men_n53_), .Y(men_men_n1981_));
  AOI210     u1932(.A0(men_men_n1980_), .A1(men_men_n1979_), .B0(men_men_n1981_), .Y(men_men_n1982_));
  OAI210     u1933(.A0(men_men_n1977_), .A1(men_men_n59_), .B0(men_men_n1982_), .Y(men_men_n1983_));
  AOI220     u1934(.A0(men_men_n609_), .A1(men_men_n215_), .B0(men_men_n340_), .B1(men_men_n211_), .Y(men_men_n1984_));
  NA2        u1935(.A(men_men_n654_), .B(men_men_n858_), .Y(men_men_n1985_));
  OAI210     u1936(.A0(men_men_n1985_), .A1(men_men_n1984_), .B0(men_men_n276_), .Y(men_men_n1986_));
  AOI210     u1937(.A0(men_men_n1833_), .A1(men_men_n198_), .B0(men_men_n53_), .Y(men_men_n1987_));
  NO2        u1938(.A(men_men_n131_), .B(men_men_n307_), .Y(men_men_n1988_));
  AOI220     u1939(.A0(men_men_n1988_), .A1(men_men_n876_), .B0(men_men_n596_), .B1(men_men_n316_), .Y(men_men_n1989_));
  NA2        u1940(.A(men_men_n394_), .B(men_men_n442_), .Y(men_men_n1990_));
  NO3        u1941(.A(men_men_n1990_), .B(men_men_n905_), .C(men_men_n172_), .Y(men_men_n1991_));
  AOI210     u1942(.A0(men_men_n1564_), .A1(men_men_n1048_), .B0(men_men_n1991_), .Y(men_men_n1992_));
  NA4        u1943(.A(men_men_n1992_), .B(men_men_n1989_), .C(men_men_n1987_), .D(men_men_n1986_), .Y(men_men_n1993_));
  NA3        u1944(.A(men_men_n1993_), .B(men_men_n1983_), .C(men_men_n57_), .Y(men_men_n1994_));
  BUFFER     u1945(.A(men_men_n1050_), .Y(men_men_n1995_));
  NA4        u1946(.A(men_men_n569_), .B(men_men_n1145_), .C(men_men_n415_), .D(men_men_n50_), .Y(men_men_n1996_));
  OAI210     u1947(.A0(men_men_n1988_), .A1(men_men_n1787_), .B0(x2), .Y(men_men_n1997_));
  NA4        u1948(.A(men_men_n259_), .B(men_men_n146_), .C(men_men_n250_), .D(men_men_n111_), .Y(men_men_n1998_));
  NA3        u1949(.A(men_men_n1998_), .B(men_men_n1997_), .C(men_men_n1996_), .Y(men_men_n1999_));
  AO220      u1950(.A0(men_men_n1999_), .A1(x0), .B0(men_men_n1995_), .B1(men_men_n128_), .Y(men_men_n2000_));
  NA3        u1951(.A(men_men_n688_), .B(men_men_n316_), .C(men_men_n60_), .Y(men_men_n2001_));
  NO2        u1952(.A(men_men_n1944_), .B(men_men_n363_), .Y(men_men_n2002_));
  NA2        u1953(.A(men_men_n567_), .B(men_men_n459_), .Y(men_men_n2003_));
  OAI220     u1954(.A0(men_men_n2003_), .A1(men_men_n2002_), .B0(men_men_n2001_), .B1(men_men_n67_), .Y(men_men_n2004_));
  AOI210     u1955(.A0(men_men_n523_), .A1(men_men_n411_), .B0(men_men_n128_), .Y(men_men_n2005_));
  NO2        u1956(.A(men_men_n2005_), .B(men_men_n340_), .Y(men_men_n2006_));
  OAI210     u1957(.A0(men_men_n2006_), .A1(men_men_n2004_), .B0(men_men_n91_), .Y(men_men_n2007_));
  NA3        u1958(.A(men_men_n1065_), .B(men_men_n121_), .C(men_men_n336_), .Y(men_men_n2008_));
  NA2        u1959(.A(men_men_n2008_), .B(men_men_n1585_), .Y(men_men_n2009_));
  NA2        u1960(.A(men_men_n1047_), .B(men_men_n632_), .Y(men_men_n2010_));
  NA2        u1961(.A(men_men_n1189_), .B(men_men_n1032_), .Y(men_men_n2011_));
  NA4        u1962(.A(men_men_n2011_), .B(men_men_n2010_), .C(men_men_n2009_), .D(men_men_n2007_), .Y(men_men_n2012_));
  AOI210     u1963(.A0(men_men_n2000_), .A1(x7), .B0(men_men_n2012_), .Y(men_men_n2013_));
  NA3        u1964(.A(men_men_n2013_), .B(men_men_n1994_), .C(men_men_n1975_), .Y(men34));
  NA2        u1965(.A(men_men_n382_), .B(x4), .Y(men_men_n2015_));
  NO2        u1966(.A(men_men_n1708_), .B(men_men_n758_), .Y(men_men_n2016_));
  AOI210     u1967(.A0(men_men_n2016_), .A1(men_men_n2015_), .B0(men_men_n293_), .Y(men_men_n2017_));
  INV        u1968(.A(men_men_n259_), .Y(men_men_n2018_));
  AOI210     u1969(.A0(men_men_n856_), .A1(men_men_n1067_), .B0(men_men_n2018_), .Y(men_men_n2019_));
  AOI210     u1970(.A0(men_men_n1774_), .A1(men_men_n480_), .B0(men_men_n130_), .Y(men_men_n2020_));
  NA2        u1971(.A(men_men_n1708_), .B(x0), .Y(men_men_n2021_));
  OAI210     u1972(.A0(men_men_n1594_), .A1(men_men_n860_), .B0(men_men_n2021_), .Y(men_men_n2022_));
  NO4        u1973(.A(men_men_n2022_), .B(men_men_n2020_), .C(men_men_n2019_), .D(men_men_n2017_), .Y(men_men_n2023_));
  NO2        u1974(.A(men_men_n2023_), .B(men_men_n421_), .Y(men_men_n2024_));
  NA2        u1975(.A(men_men_n655_), .B(x8), .Y(men_men_n2025_));
  AO210      u1976(.A0(men_men_n2025_), .A1(men_men_n431_), .B0(men_men_n586_), .Y(men_men_n2026_));
  NA2        u1977(.A(men_men_n596_), .B(men_men_n559_), .Y(men_men_n2027_));
  AOI210     u1978(.A0(men_men_n2027_), .A1(men_men_n2026_), .B0(men_men_n240_), .Y(men_men_n2028_));
  OAI210     u1979(.A0(men_men_n111_), .A1(men_men_n927_), .B0(men_men_n1282_), .Y(men_men_n2029_));
  OAI210     u1980(.A0(men_men_n1402_), .A1(men_men_n58_), .B0(men_men_n2029_), .Y(men_men_n2030_));
  NA3        u1981(.A(men_men_n2030_), .B(men_men_n308_), .C(x8), .Y(men_men_n2031_));
  NO3        u1982(.A(men_men_n875_), .B(men_men_n630_), .C(men_men_n400_), .Y(men_men_n2032_));
  AOI210     u1983(.A0(men_men_n1386_), .A1(men_men_n296_), .B0(men_men_n2032_), .Y(men_men_n2033_));
  NA2        u1984(.A(men_men_n590_), .B(men_men_n293_), .Y(men_men_n2034_));
  NA2        u1985(.A(men_men_n124_), .B(x0), .Y(men_men_n2035_));
  NAi31      u1986(.An(men_men_n2035_), .B(men_men_n2034_), .C(men_men_n711_), .Y(men_men_n2036_));
  NA3        u1987(.A(men_men_n1397_), .B(men_men_n1226_), .C(men_men_n50_), .Y(men_men_n2037_));
  NA4        u1988(.A(men_men_n2037_), .B(men_men_n2036_), .C(men_men_n2033_), .D(men_men_n2031_), .Y(men_men_n2038_));
  AOI210     u1989(.A0(men_men_n493_), .A1(men_men_n724_), .B0(men_men_n231_), .Y(men_men_n2039_));
  OAI220     u1990(.A0(men_men_n2039_), .A1(men_men_n59_), .B0(men_men_n990_), .B1(men_men_n55_), .Y(men_men_n2040_));
  NA3        u1991(.A(men_men_n2040_), .B(men_men_n655_), .C(men_men_n56_), .Y(men_men_n2041_));
  INV        u1992(.A(men_men_n2041_), .Y(men_men_n2042_));
  NO4        u1993(.A(men_men_n2042_), .B(men_men_n2038_), .C(men_men_n2028_), .D(men_men_n2024_), .Y(men_men_n2043_));
  NO3        u1994(.A(men_men_n53_), .B(men_men_n392_), .C(men_men_n296_), .Y(men_men_n2044_));
  NO3        u1995(.A(men_men_n1925_), .B(men_men_n276_), .C(men_men_n966_), .Y(men_men_n2045_));
  NO2        u1996(.A(men_men_n2045_), .B(men_men_n1362_), .Y(men_men_n2046_));
  OAI210     u1997(.A0(men_men_n2046_), .A1(men_men_n2044_), .B0(x2), .Y(men_men_n2047_));
  OAI210     u1998(.A0(men_men_n766_), .A1(men_men_n327_), .B0(men_men_n2047_), .Y(men_men_n2048_));
  NA2        u1999(.A(men_men_n286_), .B(x4), .Y(men_men_n2049_));
  OAI220     u2000(.A0(men_men_n661_), .A1(men_men_n55_), .B0(men_men_n253_), .B1(men_men_n96_), .Y(men_men_n2050_));
  NO4        u2001(.A(men_men_n396_), .B(men_men_n71_), .C(x7), .D(x3), .Y(men_men_n2051_));
  NO2        u2002(.A(men_men_n979_), .B(men_men_n260_), .Y(men_men_n2052_));
  NO4        u2003(.A(men_men_n2052_), .B(men_men_n2051_), .C(men_men_n2050_), .D(men_men_n2049_), .Y(men_men_n2053_));
  NA4        u2004(.A(men_men_n655_), .B(men_men_n168_), .C(men_men_n57_), .D(men_men_n97_), .Y(men_men_n2054_));
  INV        u2005(.A(men_men_n2054_), .Y(men_men_n2055_));
  OAI210     u2006(.A0(men_men_n2055_), .A1(men_men_n2053_), .B0(men_men_n154_), .Y(men_men_n2056_));
  NA2        u2007(.A(men_men_n79_), .B(x0), .Y(men_men_n2057_));
  NA4        u2008(.A(men_men_n2057_), .B(men_men_n1019_), .C(men_men_n269_), .D(men_men_n521_), .Y(men_men_n2058_));
  NA2        u2009(.A(men_men_n890_), .B(men_men_n587_), .Y(men_men_n2059_));
  NO2        u2010(.A(men_men_n1783_), .B(men_men_n237_), .Y(men_men_n2060_));
  AOI220     u2011(.A0(men_men_n359_), .A1(x8), .B0(men_men_n83_), .B1(x2), .Y(men_men_n2061_));
  NO2        u2012(.A(men_men_n2061_), .B(men_men_n1178_), .Y(men_men_n2062_));
  AOI220     u2013(.A0(men_men_n2062_), .A1(men_men_n1163_), .B0(men_men_n2060_), .B1(men_men_n1324_), .Y(men_men_n2063_));
  NA4        u2014(.A(men_men_n2063_), .B(men_men_n2059_), .C(men_men_n2058_), .D(men_men_n2056_), .Y(men_men_n2064_));
  AOI210     u2015(.A0(men_men_n2048_), .A1(men_men_n724_), .B0(men_men_n2064_), .Y(men_men_n2065_));
  OAI210     u2016(.A0(men_men_n2043_), .A1(x2), .B0(men_men_n2065_), .Y(men35));
  NA2        u2017(.A(men_men_n447_), .B(men_men_n168_), .Y(men_men_n2067_));
  AOI220     u2018(.A0(men_men_n567_), .A1(men_men_n55_), .B0(men_men_n688_), .B1(men_men_n1079_), .Y(men_men_n2068_));
  AOI210     u2019(.A0(men_men_n2068_), .A1(men_men_n2067_), .B0(men_men_n67_), .Y(men_men_n2069_));
  NO3        u2020(.A(men_men_n455_), .B(men_men_n411_), .C(men_men_n307_), .Y(men_men_n2070_));
  OAI210     u2021(.A0(men_men_n2070_), .A1(men_men_n2069_), .B0(x2), .Y(men_men_n2071_));
  AOI210     u2022(.A0(men_men_n199_), .A1(x0), .B0(men_men_n248_), .Y(men_men_n2072_));
  OAI220     u2023(.A0(men_men_n2072_), .A1(men_men_n592_), .B0(men_men_n185_), .B1(x4), .Y(men_men_n2073_));
  NA2        u2024(.A(men_men_n2073_), .B(men_men_n128_), .Y(men_men_n2074_));
  NA3        u2025(.A(men_men_n359_), .B(x8), .C(men_men_n67_), .Y(men_men_n2075_));
  AOI210     u2026(.A0(men_men_n2075_), .A1(men_men_n1503_), .B0(men_men_n609_), .Y(men_men_n2076_));
  OAI210     u2027(.A0(men_men_n2001_), .A1(x6), .B0(men_men_n664_), .Y(men_men_n2077_));
  NO2        u2028(.A(men_men_n2077_), .B(men_men_n2076_), .Y(men_men_n2078_));
  NA3        u2029(.A(men_men_n2078_), .B(men_men_n2074_), .C(men_men_n2071_), .Y(men_men_n2079_));
  NAi21      u2030(.An(men_men_n1474_), .B(men_men_n1141_), .Y(men_men_n2080_));
  NO2        u2031(.A(men_men_n382_), .B(men_men_n375_), .Y(men_men_n2081_));
  AOI210     u2032(.A0(men_men_n2080_), .A1(men_men_n56_), .B0(men_men_n2081_), .Y(men_men_n2082_));
  NA2        u2033(.A(men_men_n678_), .B(men_men_n622_), .Y(men_men_n2083_));
  NA2        u2034(.A(men_men_n1170_), .B(men_men_n62_), .Y(men_men_n2084_));
  OAI210     u2035(.A0(men_men_n947_), .A1(x6), .B0(men_men_n416_), .Y(men_men_n2085_));
  NA2        u2036(.A(men_men_n2085_), .B(men_men_n2084_), .Y(men_men_n2086_));
  NA2        u2037(.A(men_men_n2086_), .B(men_men_n50_), .Y(men_men_n2087_));
  OAI210     u2038(.A0(men_men_n2083_), .A1(men_men_n2082_), .B0(men_men_n2087_), .Y(men_men_n2088_));
  AOI210     u2039(.A0(men_men_n2079_), .A1(men_men_n57_), .B0(men_men_n2088_), .Y(men_men_n2089_));
  NO3        u2040(.A(men_men_n947_), .B(men_men_n501_), .C(men_men_n112_), .Y(men_men_n2090_));
  OAI210     u2041(.A0(men_men_n147_), .A1(men_men_n64_), .B0(men_men_n2090_), .Y(men_men_n2091_));
  NO2        u2042(.A(men_men_n2091_), .B(men_men_n50_), .Y(men_men_n2092_));
  NA4        u2043(.A(men_men_n411_), .B(men_men_n211_), .C(men_men_n771_), .D(men_men_n93_), .Y(men_men_n2093_));
  INV        u2044(.A(men_men_n2093_), .Y(men_men_n2094_));
  OAI210     u2045(.A0(men_men_n2094_), .A1(men_men_n2092_), .B0(men_men_n59_), .Y(men_men_n2095_));
  AOI210     u2046(.A0(men_men_n762_), .A1(men_men_n475_), .B0(men_men_n1661_), .Y(men_men_n2096_));
  AOI210     u2047(.A0(men_men_n501_), .A1(men_men_n541_), .B0(men_men_n2096_), .Y(men_men_n2097_));
  INV        u2048(.A(men_men_n1278_), .Y(men_men_n2098_));
  OAI210     u2049(.A0(men_men_n2097_), .A1(x3), .B0(men_men_n2098_), .Y(men_men_n2099_));
  NA3        u2050(.A(men_men_n954_), .B(men_men_n722_), .C(men_men_n231_), .Y(men_men_n2100_));
  INV        u2051(.A(men_men_n2100_), .Y(men_men_n2101_));
  AOI210     u2052(.A0(men_men_n2099_), .A1(men_men_n523_), .B0(men_men_n2101_), .Y(men_men_n2102_));
  AOI210     u2053(.A0(men_men_n1257_), .A1(men_men_n574_), .B0(men_men_n607_), .Y(men_men_n2103_));
  OAI210     u2054(.A0(men_men_n1711_), .A1(men_men_n541_), .B0(men_men_n1944_), .Y(men_men_n2104_));
  OAI210     u2055(.A0(men_men_n2025_), .A1(x4), .B0(men_men_n2104_), .Y(men_men_n2105_));
  OAI210     u2056(.A0(men_men_n2105_), .A1(men_men_n2103_), .B0(men_men_n83_), .Y(men_men_n2106_));
  NO2        u2057(.A(men_men_n757_), .B(men_men_n588_), .Y(men_men_n2107_));
  NO2        u2058(.A(men_men_n260_), .B(x6), .Y(men_men_n2108_));
  OAI210     u2059(.A0(men_men_n2107_), .A1(men_men_n1559_), .B0(men_men_n2108_), .Y(men_men_n2109_));
  NA4        u2060(.A(men_men_n2109_), .B(men_men_n2106_), .C(men_men_n2102_), .D(men_men_n2095_), .Y(men_men_n2110_));
  AOI210     u2061(.A0(men_men_n99_), .A1(men_men_n376_), .B0(x1), .Y(men_men_n2111_));
  NO2        u2062(.A(men_men_n654_), .B(men_men_n607_), .Y(men_men_n2112_));
  OAI210     u2063(.A0(men_men_n411_), .A1(men_men_n158_), .B0(men_men_n708_), .Y(men_men_n2113_));
  AOI210     u2064(.A0(men_men_n2113_), .A1(men_men_n895_), .B0(men_men_n53_), .Y(men_men_n2114_));
  NO3        u2065(.A(men_men_n2114_), .B(men_men_n2112_), .C(men_men_n2111_), .Y(men_men_n2115_));
  NA3        u2066(.A(men_men_n1259_), .B(men_men_n1119_), .C(men_men_n728_), .Y(men_men_n2116_));
  AOI220     u2067(.A0(men_men_n1700_), .A1(men_men_n128_), .B0(men_men_n368_), .B1(men_men_n115_), .Y(men_men_n2117_));
  AOI210     u2068(.A0(men_men_n2117_), .A1(men_men_n2116_), .B0(men_men_n1318_), .Y(men_men_n2118_));
  NO2        u2069(.A(men_men_n567_), .B(x3), .Y(men_men_n2119_));
  NO3        u2070(.A(men_men_n617_), .B(men_men_n1402_), .C(x2), .Y(men_men_n2120_));
  AOI220     u2071(.A0(men_men_n2120_), .A1(men_men_n2119_), .B0(men_men_n1673_), .B1(men_men_n684_), .Y(men_men_n2121_));
  NO2        u2072(.A(men_men_n1154_), .B(x8), .Y(men_men_n2122_));
  NA2        u2073(.A(men_men_n2122_), .B(men_men_n368_), .Y(men_men_n2123_));
  OAI210     u2074(.A0(men_men_n2121_), .A1(men_men_n1030_), .B0(men_men_n2123_), .Y(men_men_n2124_));
  NO2        u2075(.A(men_men_n2124_), .B(men_men_n2118_), .Y(men_men_n2125_));
  OAI210     u2076(.A0(men_men_n2115_), .A1(men_men_n286_), .B0(men_men_n2125_), .Y(men_men_n2126_));
  AOI210     u2077(.A0(men_men_n2110_), .A1(x5), .B0(men_men_n2126_), .Y(men_men_n2127_));
  OAI210     u2078(.A0(men_men_n2089_), .A1(x5), .B0(men_men_n2127_), .Y(men36));
  NO2        u2079(.A(men_men_n764_), .B(men_men_n275_), .Y(men_men_n2129_));
  NO3        u2080(.A(men_men_n111_), .B(men_men_n927_), .C(men_men_n55_), .Y(men_men_n2130_));
  NO3        u2081(.A(men_men_n2130_), .B(men_men_n1730_), .C(men_men_n947_), .Y(men_men_n2131_));
  OAI210     u2082(.A0(men_men_n2131_), .A1(men_men_n2129_), .B0(men_men_n99_), .Y(men_men_n2132_));
  OR3        u2083(.A(men_men_n717_), .B(men_men_n331_), .C(men_men_n437_), .Y(men_men_n2133_));
  INV        u2084(.A(men_men_n882_), .Y(men_men_n2134_));
  NA2        u2085(.A(men_men_n2134_), .B(men_men_n253_), .Y(men_men_n2135_));
  NA3        u2086(.A(men_men_n2135_), .B(men_men_n2133_), .C(men_men_n2132_), .Y(men_men_n2136_));
  NO3        u2087(.A(men_men_n2310_), .B(men_men_n872_), .C(men_men_n478_), .Y(men_men_n2137_));
  AOI220     u2088(.A0(men_men_n276_), .A1(x1), .B0(men_men_n127_), .B1(x6), .Y(men_men_n2138_));
  AOI210     u2089(.A0(men_men_n966_), .A1(x6), .B0(men_men_n372_), .Y(men_men_n2139_));
  OAI220     u2090(.A0(men_men_n2139_), .A1(men_men_n322_), .B0(men_men_n2138_), .B1(men_men_n412_), .Y(men_men_n2140_));
  OAI210     u2091(.A0(men_men_n2140_), .A1(men_men_n2137_), .B0(men_men_n411_), .Y(men_men_n2141_));
  NA2        u2092(.A(men_men_n596_), .B(men_men_n437_), .Y(men_men_n2142_));
  NO2        u2093(.A(men_men_n2142_), .B(men_men_n241_), .Y(men_men_n2143_));
  NO2        u2094(.A(men_men_n2143_), .B(men_men_n370_), .Y(men_men_n2144_));
  OAI210     u2095(.A0(men_men_n569_), .A1(men_men_n716_), .B0(men_men_n863_), .Y(men_men_n2145_));
  NO2        u2096(.A(men_men_n1443_), .B(men_men_n1438_), .Y(men_men_n2146_));
  AOI220     u2097(.A0(men_men_n2146_), .A1(men_men_n109_), .B0(men_men_n2145_), .B1(men_men_n559_), .Y(men_men_n2147_));
  NA3        u2098(.A(men_men_n2147_), .B(men_men_n2144_), .C(men_men_n2141_), .Y(men_men_n2148_));
  AOI210     u2099(.A0(men_men_n2136_), .A1(men_men_n308_), .B0(men_men_n2148_), .Y(men_men_n2149_));
  OAI210     u2100(.A0(men_men_n528_), .A1(men_men_n460_), .B0(men_men_n158_), .Y(men_men_n2150_));
  OAI210     u2101(.A0(men_men_n1741_), .A1(men_men_n66_), .B0(men_men_n2150_), .Y(men_men_n2151_));
  NA2        u2102(.A(men_men_n217_), .B(men_men_n232_), .Y(men_men_n2152_));
  NO2        u2103(.A(men_men_n1747_), .B(men_men_n164_), .Y(men_men_n2153_));
  NA2        u2104(.A(men_men_n1067_), .B(men_men_n55_), .Y(men_men_n2154_));
  OAI210     u2105(.A0(men_men_n2154_), .A1(men_men_n2153_), .B0(men_men_n2152_), .Y(men_men_n2155_));
  OAI210     u2106(.A0(men_men_n2155_), .A1(men_men_n2151_), .B0(men_men_n791_), .Y(men_men_n2156_));
  AOI210     u2107(.A0(men_men_n96_), .A1(men_men_n99_), .B0(men_men_n309_), .Y(men_men_n2157_));
  NA2        u2108(.A(men_men_n596_), .B(men_men_n1402_), .Y(men_men_n2158_));
  OAI220     u2109(.A0(men_men_n2158_), .A1(men_men_n2157_), .B0(men_men_n664_), .B1(men_men_n1105_), .Y(men_men_n2159_));
  NO2        u2110(.A(men_men_n1226_), .B(men_men_n515_), .Y(men_men_n2160_));
  NO3        u2111(.A(men_men_n2160_), .B(men_men_n1563_), .C(men_men_n617_), .Y(men_men_n2161_));
  NOi31      u2112(.An(men_men_n1754_), .B(men_men_n1990_), .C(men_men_n674_), .Y(men_men_n2162_));
  NO3        u2113(.A(men_men_n2162_), .B(men_men_n2161_), .C(men_men_n2159_), .Y(men_men_n2163_));
  AOI210     u2114(.A0(men_men_n2163_), .A1(men_men_n2156_), .B0(x7), .Y(men_men_n2164_));
  NA2        u2115(.A(men_men_n127_), .B(men_men_n62_), .Y(men_men_n2165_));
  AOI210     u2116(.A0(men_men_n523_), .A1(men_men_n554_), .B0(men_men_n1048_), .Y(men_men_n2166_));
  NA4        u2117(.A(men_men_n2166_), .B(men_men_n2165_), .C(men_men_n875_), .D(men_men_n784_), .Y(men_men_n2167_));
  NA2        u2118(.A(men_men_n2167_), .B(men_men_n447_), .Y(men_men_n2168_));
  AOI220     u2119(.A0(men_men_n1524_), .A1(men_men_n235_), .B0(men_men_n925_), .B1(men_men_n115_), .Y(men_men_n2169_));
  NO2        u2120(.A(men_men_n2169_), .B(men_men_n394_), .Y(men_men_n2170_));
  NO2        u2121(.A(men_men_n357_), .B(men_men_n208_), .Y(men_men_n2171_));
  NO3        u2122(.A(men_men_n2171_), .B(men_men_n1123_), .C(men_men_n59_), .Y(men_men_n2172_));
  AOI210     u2123(.A0(men_men_n1083_), .A1(men_men_n358_), .B0(x6), .Y(men_men_n2173_));
  NA3        u2124(.A(men_men_n1465_), .B(men_men_n253_), .C(men_men_n245_), .Y(men_men_n2174_));
  NA2        u2125(.A(men_men_n2174_), .B(men_men_n1424_), .Y(men_men_n2175_));
  NO4        u2126(.A(men_men_n2175_), .B(men_men_n2173_), .C(men_men_n2172_), .D(men_men_n2170_), .Y(men_men_n2176_));
  AOI210     u2127(.A0(men_men_n2176_), .A1(men_men_n2168_), .B0(men_men_n400_), .Y(men_men_n2177_));
  OAI210     u2128(.A0(men_men_n769_), .A1(men_men_n249_), .B0(men_men_n351_), .Y(men_men_n2178_));
  NA2        u2129(.A(men_men_n1067_), .B(men_men_n162_), .Y(men_men_n2179_));
  NO2        u2130(.A(men_men_n548_), .B(men_men_n99_), .Y(men_men_n2180_));
  AO210      u2131(.A0(men_men_n2180_), .A1(men_men_n2179_), .B0(men_men_n1538_), .Y(men_men_n2181_));
  NO2        u2132(.A(men_men_n407_), .B(men_men_n369_), .Y(men_men_n2182_));
  AOI220     u2133(.A0(men_men_n2182_), .A1(men_men_n2181_), .B0(men_men_n2178_), .B1(men_men_n267_), .Y(men_men_n2183_));
  INV        u2134(.A(men_men_n2183_), .Y(men_men_n2184_));
  NO3        u2135(.A(men_men_n2184_), .B(men_men_n2177_), .C(men_men_n2164_), .Y(men_men_n2185_));
  OAI210     u2136(.A0(men_men_n2149_), .A1(men_men_n57_), .B0(men_men_n2185_), .Y(men37));
  NA3        u2137(.A(men_men_n946_), .B(men_men_n130_), .C(x3), .Y(men_men_n2187_));
  NA3        u2138(.A(men_men_n697_), .B(men_men_n150_), .C(men_men_n50_), .Y(men_men_n2188_));
  AOI210     u2139(.A0(men_men_n2188_), .A1(men_men_n2187_), .B0(men_men_n610_), .Y(men_men_n2189_));
  NO3        u2140(.A(men_men_n946_), .B(men_men_n331_), .C(men_men_n454_), .Y(men_men_n2190_));
  OAI210     u2141(.A0(men_men_n2190_), .A1(men_men_n2189_), .B0(men_men_n56_), .Y(men_men_n2191_));
  NO2        u2142(.A(men_men_n591_), .B(men_men_n171_), .Y(men_men_n2192_));
  NO2        u2143(.A(men_men_n2192_), .B(men_men_n2319_), .Y(men_men_n2193_));
  NA2        u2144(.A(men_men_n2193_), .B(men_men_n67_), .Y(men_men_n2194_));
  NA2        u2145(.A(men_men_n2194_), .B(men_men_n2191_), .Y(men_men_n2195_));
  NA2        u2146(.A(men_men_n375_), .B(men_men_n127_), .Y(men_men_n2196_));
  NO2        u2147(.A(men_men_n1491_), .B(men_men_n98_), .Y(men_men_n2197_));
  AOI210     u2148(.A0(men_men_n1731_), .A1(men_men_n765_), .B0(men_men_n2197_), .Y(men_men_n2198_));
  OAI220     u2149(.A0(men_men_n2198_), .A1(men_men_n51_), .B0(men_men_n1403_), .B1(men_men_n2196_), .Y(men_men_n2199_));
  AOI210     u2150(.A0(men_men_n2195_), .A1(men_men_n65_), .B0(men_men_n2199_), .Y(men_men_n2200_));
  OAI210     u2151(.A0(men_men_n245_), .A1(men_men_n969_), .B0(men_men_n432_), .Y(men_men_n2201_));
  NA2        u2152(.A(men_men_n2201_), .B(men_men_n927_), .Y(men_men_n2202_));
  NA3        u2153(.A(men_men_n355_), .B(men_men_n728_), .C(men_men_n99_), .Y(men_men_n2203_));
  NO2        u2154(.A(men_men_n473_), .B(men_men_n56_), .Y(men_men_n2204_));
  NA2        u2155(.A(men_men_n2204_), .B(men_men_n2203_), .Y(men_men_n2205_));
  AOI210     u2156(.A0(x6), .A1(men_men_n454_), .B0(men_men_n2205_), .Y(men_men_n2206_));
  NO2        u2157(.A(men_men_n1041_), .B(men_men_n249_), .Y(men_men_n2207_));
  OAI210     u2158(.A0(men_men_n267_), .A1(men_men_n239_), .B0(men_men_n2207_), .Y(men_men_n2208_));
  OAI210     u2159(.A0(men_men_n593_), .A1(men_men_n128_), .B0(x3), .Y(men_men_n2209_));
  AOI210     u2160(.A0(men_men_n593_), .A1(men_men_n326_), .B0(men_men_n2209_), .Y(men_men_n2210_));
  OAI210     u2161(.A0(men_men_n53_), .A1(men_men_n354_), .B0(men_men_n56_), .Y(men_men_n2211_));
  NO2        u2162(.A(men_men_n2211_), .B(men_men_n2210_), .Y(men_men_n2212_));
  AOI220     u2163(.A0(men_men_n2212_), .A1(men_men_n2208_), .B0(men_men_n2206_), .B1(men_men_n2202_), .Y(men_men_n2213_));
  OAI210     u2164(.A0(men_men_n2213_), .A1(men_men_n1536_), .B0(men_men_n91_), .Y(men_men_n2214_));
  NA2        u2165(.A(men_men_n617_), .B(men_men_n1053_), .Y(men_men_n2215_));
  NOi21      u2166(.An(men_men_n1195_), .B(men_men_n100_), .Y(men_men_n2216_));
  AOI210     u2167(.A0(men_men_n2216_), .A1(men_men_n2215_), .B0(men_men_n385_), .Y(men_men_n2217_));
  NO2        u2168(.A(men_men_n1922_), .B(men_men_n55_), .Y(men_men_n2218_));
  OAI210     u2169(.A0(men_men_n2218_), .A1(men_men_n2217_), .B0(men_men_n1585_), .Y(men_men_n2219_));
  NA2        u2170(.A(men_men_n168_), .B(men_men_n97_), .Y(men_men_n2220_));
  NA2        u2171(.A(men_men_n609_), .B(x6), .Y(men_men_n2221_));
  AOI210     u2172(.A0(men_men_n2221_), .A1(men_men_n431_), .B0(men_men_n2220_), .Y(men_men_n2222_));
  AOI210     u2173(.A0(men_men_n317_), .A1(men_men_n130_), .B0(men_men_n131_), .Y(men_men_n2223_));
  OAI210     u2174(.A0(men_men_n2223_), .A1(men_men_n2222_), .B0(men_men_n313_), .Y(men_men_n2224_));
  AOI210     u2175(.A0(men_men_n549_), .A1(men_men_n385_), .B0(men_men_n1131_), .Y(men_men_n2225_));
  NO3        u2176(.A(men_men_n2225_), .B(men_men_n241_), .C(men_men_n62_), .Y(men_men_n2226_));
  OAI220     u2177(.A0(men_men_n2025_), .A1(men_men_n429_), .B0(men_men_n1817_), .B1(men_men_n340_), .Y(men_men_n2227_));
  OAI210     u2178(.A0(men_men_n2227_), .A1(men_men_n2226_), .B0(men_men_n53_), .Y(men_men_n2228_));
  NO4        u2179(.A(men_men_n2035_), .B(men_men_n818_), .C(men_men_n386_), .D(men_men_n203_), .Y(men_men_n2229_));
  NO4        u2180(.A(men_men_n655_), .B(men_men_n538_), .C(men_men_n392_), .D(men_men_n935_), .Y(men_men_n2230_));
  NO3        u2181(.A(men_men_n2230_), .B(men_men_n2229_), .C(men_men_n941_), .Y(men_men_n2231_));
  NA4        u2182(.A(men_men_n2231_), .B(men_men_n2228_), .C(men_men_n2224_), .D(men_men_n2219_), .Y(men_men_n2232_));
  NO3        u2183(.A(men_men_n227_), .B(men_men_n316_), .C(men_men_n76_), .Y(men_men_n2233_));
  NO3        u2184(.A(men_men_n53_), .B(men_men_n1067_), .C(men_men_n1085_), .Y(men_men_n2234_));
  OAI220     u2185(.A0(men_men_n2234_), .A1(men_men_n2233_), .B0(men_men_n411_), .B1(men_men_n77_), .Y(men_men_n2235_));
  INV        u2186(.A(men_men_n341_), .Y(men_men_n2236_));
  AOI210     u2187(.A0(men_men_n2236_), .A1(men_men_n2318_), .B0(x1), .Y(men_men_n2237_));
  NA2        u2188(.A(men_men_n240_), .B(men_men_n76_), .Y(men_men_n2238_));
  NO2        u2189(.A(men_men_n354_), .B(men_men_n2238_), .Y(men_men_n2239_));
  NA2        u2190(.A(men_men_n979_), .B(men_men_n61_), .Y(men_men_n2240_));
  NA2        u2191(.A(men_men_n1023_), .B(men_men_n164_), .Y(men_men_n2241_));
  OAI210     u2192(.A0(men_men_n2240_), .A1(men_men_n285_), .B0(men_men_n2241_), .Y(men_men_n2242_));
  NO3        u2193(.A(men_men_n2242_), .B(men_men_n2239_), .C(men_men_n2237_), .Y(men_men_n2243_));
  OAI210     u2194(.A0(men_men_n2243_), .A1(x6), .B0(men_men_n2235_), .Y(men_men_n2244_));
  AOI220     u2195(.A0(men_men_n2244_), .A1(men_men_n1282_), .B0(men_men_n2232_), .B1(men_men_n57_), .Y(men_men_n2245_));
  NA3        u2196(.A(men_men_n2245_), .B(men_men_n2214_), .C(men_men_n2200_), .Y(men38));
  AOI210     u2197(.A0(men_men_n1453_), .A1(men_men_n177_), .B0(men_men_n858_), .Y(men_men_n2247_));
  NO2        u2198(.A(men_men_n514_), .B(men_men_n963_), .Y(men_men_n2248_));
  NO2        u2199(.A(men_men_n1615_), .B(men_men_n210_), .Y(men_men_n2249_));
  NO3        u2200(.A(men_men_n1140_), .B(men_men_n293_), .C(x8), .Y(men_men_n2250_));
  NO4        u2201(.A(men_men_n2250_), .B(men_men_n2249_), .C(men_men_n2248_), .D(men_men_n2247_), .Y(men_men_n2251_));
  NO2        u2202(.A(men_men_n2251_), .B(x6), .Y(men_men_n2252_));
  AOI210     u2203(.A0(men_men_n386_), .A1(men_men_n356_), .B0(men_men_n1512_), .Y(men_men_n2253_));
  NO2        u2204(.A(men_men_n722_), .B(men_men_n83_), .Y(men_men_n2254_));
  OAI210     u2205(.A0(men_men_n899_), .A1(men_men_n138_), .B0(men_men_n321_), .Y(men_men_n2255_));
  OAI220     u2206(.A0(men_men_n2255_), .A1(men_men_n2254_), .B0(men_men_n2253_), .B1(men_men_n179_), .Y(men_men_n2256_));
  NA2        u2207(.A(men_men_n2256_), .B(x6), .Y(men_men_n2257_));
  NO3        u2208(.A(men_men_n2308_), .B(men_men_n1474_), .C(men_men_n234_), .Y(men_men_n2258_));
  NO3        u2209(.A(x3), .B(men_men_n53_), .C(x0), .Y(men_men_n2259_));
  OAI210     u2210(.A0(men_men_n466_), .A1(x2), .B0(men_men_n2259_), .Y(men_men_n2260_));
  NA3        u2211(.A(men_men_n385_), .B(men_men_n375_), .C(men_men_n266_), .Y(men_men_n2261_));
  NA3        u2212(.A(men_men_n2261_), .B(men_men_n2260_), .C(men_men_n1580_), .Y(men_men_n2262_));
  OAI210     u2213(.A0(men_men_n2262_), .A1(men_men_n2258_), .B0(men_men_n724_), .Y(men_men_n2263_));
  AN3        u2214(.A(men_men_n729_), .B(men_men_n697_), .C(x0), .Y(men_men_n2264_));
  NA2        u2215(.A(men_men_n2264_), .B(men_men_n297_), .Y(men_men_n2265_));
  OAI220     u2216(.A0(men_men_n538_), .A1(men_men_n250_), .B0(men_men_n728_), .B1(men_men_n84_), .Y(men_men_n2266_));
  OAI210     u2217(.A0(men_men_n609_), .A1(x0), .B0(men_men_n51_), .Y(men_men_n2267_));
  INV        u2218(.A(men_men_n209_), .Y(men_men_n2268_));
  AOI220     u2219(.A0(men_men_n2268_), .A1(men_men_n2267_), .B0(men_men_n2266_), .B1(men_men_n355_), .Y(men_men_n2269_));
  NA4        u2220(.A(men_men_n2269_), .B(men_men_n2265_), .C(men_men_n2263_), .D(men_men_n2257_), .Y(men_men_n2270_));
  OAI210     u2221(.A0(men_men_n2270_), .A1(men_men_n2252_), .B0(x7), .Y(men_men_n2271_));
  AOI210     u2222(.A0(men_men_n329_), .A1(x1), .B0(men_men_n1088_), .Y(men_men_n2272_));
  NO2        u2223(.A(men_men_n2272_), .B(men_men_n51_), .Y(men_men_n2273_));
  AOI210     u2224(.A0(men_men_n83_), .A1(men_men_n67_), .B0(men_men_n1944_), .Y(men_men_n2274_));
  NO2        u2225(.A(men_men_n1528_), .B(men_men_n473_), .Y(men_men_n2275_));
  OAI210     u2226(.A0(men_men_n2312_), .A1(men_men_n2274_), .B0(men_men_n2275_), .Y(men_men_n2276_));
  OAI210     u2227(.A0(men_men_n2276_), .A1(men_men_n2273_), .B0(x4), .Y(men_men_n2277_));
  NO2        u2228(.A(men_men_n1539_), .B(men_men_n405_), .Y(men_men_n2278_));
  NO3        u2229(.A(men_men_n2278_), .B(men_men_n354_), .C(men_men_n109_), .Y(men_men_n2279_));
  AOI210     u2230(.A0(men_men_n935_), .A1(men_men_n219_), .B0(men_men_n349_), .Y(men_men_n2280_));
  AO210      u2231(.A0(men_men_n1146_), .A1(x6), .B0(men_men_n2280_), .Y(men_men_n2281_));
  NO2        u2232(.A(men_men_n1245_), .B(men_men_n128_), .Y(men_men_n2282_));
  NA2        u2233(.A(men_men_n1708_), .B(men_men_n295_), .Y(men_men_n2283_));
  OAI220     u2234(.A0(men_men_n2283_), .A1(men_men_n951_), .B0(men_men_n2282_), .B1(men_men_n1599_), .Y(men_men_n2284_));
  NO3        u2235(.A(men_men_n2284_), .B(men_men_n2281_), .C(men_men_n2279_), .Y(men_men_n2285_));
  AOI210     u2236(.A0(men_men_n2285_), .A1(men_men_n2277_), .B0(men_men_n97_), .Y(men_men_n2286_));
  NA3        u2237(.A(men_men_n1700_), .B(men_men_n538_), .C(men_men_n154_), .Y(men_men_n2287_));
  AOI210     u2238(.A0(men_men_n2287_), .A1(men_men_n1253_), .B0(men_men_n211_), .Y(men_men_n2288_));
  AOI210     u2239(.A0(men_men_n447_), .A1(men_men_n437_), .B0(men_men_n606_), .Y(men_men_n2289_));
  OAI220     u2240(.A0(men_men_n2289_), .A1(men_men_n412_), .B0(men_men_n185_), .B1(men_men_n107_), .Y(men_men_n2290_));
  OAI210     u2241(.A0(men_men_n2290_), .A1(men_men_n2288_), .B0(x0), .Y(men_men_n2291_));
  NA3        u2242(.A(men_men_n356_), .B(men_men_n728_), .C(men_men_n250_), .Y(men_men_n2292_));
  AOI210     u2243(.A0(men_men_n2292_), .A1(men_men_n640_), .B0(men_men_n1911_), .Y(men_men_n2293_));
  NA2        u2244(.A(men_men_n999_), .B(men_men_n837_), .Y(men_men_n2294_));
  NA4        u2245(.A(men_men_n605_), .B(men_men_n538_), .C(men_men_n168_), .D(x3), .Y(men_men_n2295_));
  AOI210     u2246(.A0(men_men_n2295_), .A1(men_men_n2294_), .B0(men_men_n442_), .Y(men_men_n2296_));
  NO4        u2247(.A(men_men_n1240_), .B(men_men_n462_), .C(men_men_n1085_), .D(men_men_n688_), .Y(men_men_n2297_));
  OAI220     u2248(.A0(men_men_n1557_), .A1(men_men_n1978_), .B0(men_men_n209_), .B1(men_men_n140_), .Y(men_men_n2298_));
  NO4        u2249(.A(men_men_n2298_), .B(men_men_n2297_), .C(men_men_n2296_), .D(men_men_n2293_), .Y(men_men_n2299_));
  NA2        u2250(.A(men_men_n2299_), .B(men_men_n2291_), .Y(men_men_n2300_));
  OAI210     u2251(.A0(men_men_n2300_), .A1(men_men_n2286_), .B0(men_men_n57_), .Y(men_men_n2301_));
  OAI220     u2252(.A0(men_men_n1542_), .A1(men_men_n250_), .B0(men_men_n233_), .B1(men_men_n93_), .Y(men_men_n2302_));
  NO2        u2253(.A(men_men_n616_), .B(men_men_n140_), .Y(men_men_n2303_));
  AOI210     u2254(.A0(men_men_n2302_), .A1(men_men_n876_), .B0(men_men_n2303_), .Y(men_men_n2304_));
  NA3        u2255(.A(men_men_n2304_), .B(men_men_n2301_), .C(men_men_n2271_), .Y(men39));
  INV        u2256(.A(men_men_n224_), .Y(men_men_n2308_));
  INV        u2257(.A(x8), .Y(men_men_n2309_));
  INV        u2258(.A(x8), .Y(men_men_n2310_));
  INV        u2259(.A(men_men_n385_), .Y(men_men_n2311_));
  INV        u2260(.A(x3), .Y(men_men_n2312_));
  INV        u2261(.A(men_men_n1093_), .Y(men_men_n2313_));
  INV        u2262(.A(men_men_n401_), .Y(men_men_n2314_));
  INV        u2263(.A(men_men_n317_), .Y(men_men_n2315_));
  INV        u2264(.A(men_men_n128_), .Y(men_men_n2316_));
  INV        u2265(.A(x5), .Y(men_men_n2317_));
  INV        u2266(.A(men_men_n386_), .Y(men_men_n2318_));
  INV        u2267(.A(men_men_n385_), .Y(men_men_n2319_));
  INV        u2268(.A(x3), .Y(men_men_n2320_));
  INV        u2269(.A(x7), .Y(men_men_n2321_));
  INV        u2270(.A(x8), .Y(men_men_n2322_));
  INV        u2271(.A(men_men_n317_), .Y(men_men_n2323_));
  INV        u2272(.A(men_men_n77_), .Y(men_men_n2324_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
  VOTADOR g14(.A(ori14), .B(mai14), .C(men14), .Y(z14));
  VOTADOR g15(.A(ori15), .B(mai15), .C(men15), .Y(z15));
  VOTADOR g16(.A(ori16), .B(mai16), .C(men16), .Y(z16));
  VOTADOR g17(.A(ori17), .B(mai17), .C(men17), .Y(z17));
  VOTADOR g18(.A(ori18), .B(mai18), .C(men18), .Y(z18));
  VOTADOR g19(.A(ori19), .B(mai19), .C(men19), .Y(z19));
  VOTADOR g20(.A(ori20), .B(mai20), .C(men20), .Y(z20));
  VOTADOR g21(.A(ori21), .B(mai21), .C(men21), .Y(z21));
  VOTADOR g22(.A(ori22), .B(mai22), .C(men22), .Y(z22));
  VOTADOR g23(.A(ori23), .B(mai23), .C(men23), .Y(z23));
  VOTADOR g24(.A(ori24), .B(mai24), .C(men24), .Y(z24));
  VOTADOR g25(.A(ori25), .B(mai25), .C(men25), .Y(z25));
  VOTADOR g26(.A(ori26), .B(mai26), .C(men26), .Y(z26));
  VOTADOR g27(.A(ori27), .B(mai27), .C(men27), .Y(z27));
  VOTADOR g28(.A(ori28), .B(mai28), .C(men28), .Y(z28));
  VOTADOR g29(.A(ori29), .B(mai29), .C(men29), .Y(z29));
  VOTADOR g30(.A(ori30), .B(mai30), .C(men30), .Y(z30));
  VOTADOR g31(.A(ori31), .B(mai31), .C(men31), .Y(z31));
  VOTADOR g32(.A(ori32), .B(mai32), .C(men32), .Y(z32));
  VOTADOR g33(.A(ori33), .B(mai33), .C(men33), .Y(z33));
  VOTADOR g34(.A(ori34), .B(mai34), .C(men34), .Y(z34));
  VOTADOR g35(.A(ori35), .B(mai35), .C(men35), .Y(z35));
  VOTADOR g36(.A(ori36), .B(mai36), .C(men36), .Y(z36));
  VOTADOR g37(.A(ori37), .B(mai37), .C(men37), .Y(z37));
  VOTADOR g38(.A(ori38), .B(mai38), .C(men38), .Y(z38));
  VOTADOR g39(.A(ori39), .B(mai39), .C(men39), .Y(z39));
endmodule