// Benchmark "top" written by ABC on Fri Jun 21 17:49:24 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n140_, new_new_n141_, new_new_n142_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n610_,
    new_new_n611_, new_new_n612_, new_new_n613_, new_new_n614_,
    new_new_n615_, new_new_n616_, new_new_n617_, new_new_n618_,
    new_new_n619_, new_new_n620_, new_new_n621_, new_new_n622_,
    new_new_n623_, new_new_n624_, new_new_n625_, new_new_n626_,
    new_new_n627_, new_new_n628_, new_new_n629_, new_new_n630_,
    new_new_n631_, new_new_n632_, new_new_n633_, new_new_n634_,
    new_new_n635_, new_new_n636_, new_new_n637_, new_new_n638_,
    new_new_n639_, new_new_n640_, new_new_n641_, new_new_n642_,
    new_new_n643_, new_new_n644_, new_new_n645_, new_new_n646_,
    new_new_n647_, new_new_n648_, new_new_n649_, new_new_n650_,
    new_new_n651_, new_new_n652_, new_new_n653_, new_new_n654_,
    new_new_n655_, new_new_n656_, new_new_n657_, new_new_n659_,
    new_new_n660_, new_new_n661_, new_new_n662_, new_new_n663_,
    new_new_n664_, new_new_n665_, new_new_n666_, new_new_n667_,
    new_new_n668_, new_new_n669_, new_new_n670_, new_new_n671_,
    new_new_n672_, new_new_n673_, new_new_n674_, new_new_n675_,
    new_new_n676_, new_new_n677_, new_new_n678_, new_new_n679_,
    new_new_n680_, new_new_n681_, new_new_n682_, new_new_n683_,
    new_new_n684_, new_new_n685_, new_new_n686_, new_new_n687_,
    new_new_n688_, new_new_n689_, new_new_n690_, new_new_n691_,
    new_new_n692_, new_new_n693_, new_new_n694_, new_new_n695_,
    new_new_n696_, new_new_n697_, new_new_n698_, new_new_n699_,
    new_new_n700_, new_new_n701_, new_new_n702_, new_new_n703_,
    new_new_n704_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n870_, new_new_n871_,
    new_new_n872_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n55_));
  NO2        g033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  NO2        g035(.A(new_new_n57_), .B(new_new_n56_), .Y(new_new_n58_));
  NA2        g036(.A(new_new_n58_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g038(.A(i_1_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA3        g040(.A(new_new_n62_), .B(new_new_n60_), .C(new_new_n31_), .Y(new_new_n63_));
  NA2        g041(.A(i_1_), .B(i_10_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NAi31      g043(.An(new_new_n65_), .B(new_new_n63_), .C(new_new_n59_), .Y(new_new_n66_));
  NA2        g044(.A(new_new_n50_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n75_), .Y(new_new_n76_));
  OAI210     g054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g057(.A(new_new_n79_), .B(new_new_n56_), .Y(new_new_n80_));
  NO2        g058(.A(i_3_), .B(i_9_), .Y(new_new_n81_));
  NO2        g059(.A(i_3_), .B(i_7_), .Y(new_new_n82_));
  NO2        g060(.A(new_new_n81_), .B(new_new_n61_), .Y(new_new_n83_));
  INV        g061(.A(i_6_), .Y(new_new_n84_));
  OR4        g062(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n85_));
  INV        g063(.A(new_new_n85_), .Y(new_new_n86_));
  NO2        g064(.A(i_2_), .B(i_7_), .Y(new_new_n87_));
  NO2        g065(.A(new_new_n86_), .B(new_new_n87_), .Y(new_new_n88_));
  OAI210     g066(.A0(new_new_n83_), .A1(new_new_n80_), .B0(new_new_n88_), .Y(new_new_n89_));
  NAi21      g067(.An(i_6_), .B(i_10_), .Y(new_new_n90_));
  NA2        g068(.A(i_6_), .B(i_9_), .Y(new_new_n91_));
  AOI210     g069(.A0(new_new_n91_), .A1(new_new_n90_), .B0(new_new_n61_), .Y(new_new_n92_));
  NA2        g070(.A(i_2_), .B(i_6_), .Y(new_new_n93_));
  NO3        g071(.A(new_new_n93_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n94_));
  NO2        g072(.A(new_new_n94_), .B(new_new_n92_), .Y(new_new_n95_));
  AOI210     g073(.A0(new_new_n95_), .A1(new_new_n89_), .B0(new_new_n78_), .Y(new_new_n96_));
  AN3        g074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n97_));
  NAi21      g075(.An(i_6_), .B(i_11_), .Y(new_new_n98_));
  NO2        g076(.A(i_5_), .B(i_8_), .Y(new_new_n99_));
  NOi21      g077(.An(new_new_n99_), .B(new_new_n98_), .Y(new_new_n100_));
  AOI220     g078(.A0(new_new_n100_), .A1(new_new_n60_), .B0(new_new_n97_), .B1(new_new_n32_), .Y(new_new_n101_));
  INV        g079(.A(i_7_), .Y(new_new_n102_));
  NA2        g080(.A(new_new_n46_), .B(new_new_n102_), .Y(new_new_n103_));
  NO2        g081(.A(i_0_), .B(i_5_), .Y(new_new_n104_));
  NO2        g082(.A(new_new_n104_), .B(new_new_n84_), .Y(new_new_n105_));
  NA2        g083(.A(i_12_), .B(i_3_), .Y(new_new_n106_));
  INV        g084(.A(new_new_n106_), .Y(new_new_n107_));
  NA3        g085(.A(new_new_n107_), .B(new_new_n105_), .C(new_new_n103_), .Y(new_new_n108_));
  NAi21      g086(.An(i_7_), .B(i_11_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n90_), .C(new_new_n53_), .Y(new_new_n110_));
  AN2        g088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g090(.A(new_new_n78_), .B(new_new_n56_), .Y(new_new_n113_));
  NO2        g091(.A(i_8_), .B(new_new_n102_), .Y(new_new_n114_));
  NO3        g092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n61_), .B(new_new_n26_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(i_0_), .Y(new_new_n118_));
  NA2        g096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  OAI210     g097(.A0(new_new_n118_), .A1(new_new_n116_), .B0(new_new_n119_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(new_new_n115_), .Y(new_new_n121_));
  NAi41      g099(.An(new_new_n110_), .B(new_new_n121_), .C(new_new_n108_), .D(new_new_n101_), .Y(new_new_n122_));
  NOi21      g100(.An(i_1_), .B(i_5_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(i_11_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n125_));
  NA2        g103(.A(i_7_), .B(new_new_n25_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(new_new_n125_), .Y(new_new_n127_));
  NO2        g105(.A(new_new_n127_), .B(new_new_n46_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n91_), .B(new_new_n90_), .Y(new_new_n129_));
  NAi21      g107(.An(i_3_), .B(i_8_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n60_), .Y(new_new_n131_));
  NOi31      g109(.An(new_new_n131_), .B(new_new_n129_), .C(new_new_n128_), .Y(new_new_n132_));
  NO2        g110(.A(i_1_), .B(new_new_n84_), .Y(new_new_n133_));
  NO2        g111(.A(i_6_), .B(i_5_), .Y(new_new_n134_));
  NA2        g112(.A(new_new_n134_), .B(i_3_), .Y(new_new_n135_));
  AO210      g113(.A0(new_new_n135_), .A1(new_new_n47_), .B0(new_new_n133_), .Y(new_new_n136_));
  OAI220     g114(.A0(new_new_n136_), .A1(new_new_n109_), .B0(new_new_n132_), .B1(new_new_n124_), .Y(new_new_n137_));
  NO3        g115(.A(new_new_n137_), .B(new_new_n122_), .C(new_new_n96_), .Y(new_new_n138_));
  NA3        g116(.A(new_new_n138_), .B(new_new_n77_), .C(new_new_n55_), .Y(ori2));
  NO2        g117(.A(new_new_n61_), .B(new_new_n37_), .Y(new_new_n140_));
  INV        g118(.A(i_6_), .Y(new_new_n141_));
  NA2        g119(.A(new_new_n141_), .B(new_new_n140_), .Y(new_new_n142_));
  NA4        g120(.A(new_new_n142_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(ori0));
  AN2        g121(.A(i_8_), .B(i_7_), .Y(new_new_n144_));
  NA2        g122(.A(new_new_n144_), .B(i_6_), .Y(new_new_n145_));
  NO2        g123(.A(i_12_), .B(i_13_), .Y(new_new_n146_));
  NAi21      g124(.An(i_5_), .B(i_11_), .Y(new_new_n147_));
  NOi21      g125(.An(new_new_n146_), .B(new_new_n147_), .Y(new_new_n148_));
  NO2        g126(.A(i_0_), .B(i_1_), .Y(new_new_n149_));
  NA2        g127(.A(i_2_), .B(i_3_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n150_), .B(i_4_), .Y(new_new_n151_));
  NA3        g129(.A(new_new_n151_), .B(new_new_n149_), .C(new_new_n148_), .Y(new_new_n152_));
  AN2        g130(.A(new_new_n146_), .B(new_new_n81_), .Y(new_new_n153_));
  NA2        g131(.A(i_1_), .B(i_5_), .Y(new_new_n154_));
  OR2        g132(.A(i_0_), .B(i_1_), .Y(new_new_n155_));
  NO3        g133(.A(new_new_n155_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n156_));
  NAi32      g134(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n157_));
  NAi21      g135(.An(new_new_n157_), .B(new_new_n156_), .Y(new_new_n158_));
  NOi21      g136(.An(i_4_), .B(i_10_), .Y(new_new_n159_));
  NA2        g137(.A(new_new_n159_), .B(new_new_n40_), .Y(new_new_n160_));
  NOi21      g138(.An(i_4_), .B(i_9_), .Y(new_new_n161_));
  NOi21      g139(.An(i_11_), .B(i_13_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  NO2        g141(.A(i_4_), .B(i_5_), .Y(new_new_n164_));
  NAi21      g142(.An(i_12_), .B(i_11_), .Y(new_new_n165_));
  NO2        g143(.A(new_new_n71_), .B(new_new_n61_), .Y(new_new_n166_));
  NA2        g144(.A(new_new_n166_), .B(new_new_n46_), .Y(new_new_n167_));
  NA2        g145(.A(i_3_), .B(i_5_), .Y(new_new_n168_));
  NO2        g146(.A(new_new_n71_), .B(i_5_), .Y(new_new_n169_));
  NO2        g147(.A(i_13_), .B(i_10_), .Y(new_new_n170_));
  NA3        g148(.A(new_new_n170_), .B(new_new_n169_), .C(new_new_n44_), .Y(new_new_n171_));
  NO2        g149(.A(i_2_), .B(i_1_), .Y(new_new_n172_));
  NA2        g150(.A(new_new_n172_), .B(i_3_), .Y(new_new_n173_));
  NAi21      g151(.An(i_4_), .B(i_12_), .Y(new_new_n174_));
  INV        g152(.A(i_8_), .Y(new_new_n175_));
  NO3        g153(.A(i_3_), .B(new_new_n84_), .C(new_new_n48_), .Y(new_new_n176_));
  NA2        g154(.A(new_new_n176_), .B(new_new_n114_), .Y(new_new_n177_));
  NO3        g155(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n178_));
  NO3        g156(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n179_));
  NO2        g157(.A(i_3_), .B(i_8_), .Y(new_new_n180_));
  NO3        g158(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n181_));
  NA3        g159(.A(new_new_n181_), .B(new_new_n180_), .C(new_new_n40_), .Y(new_new_n182_));
  NO2        g160(.A(new_new_n104_), .B(new_new_n56_), .Y(new_new_n183_));
  INV        g161(.A(new_new_n183_), .Y(new_new_n184_));
  NO2        g162(.A(i_13_), .B(i_9_), .Y(new_new_n185_));
  NAi21      g163(.An(i_12_), .B(i_3_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n44_), .B(i_5_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n184_), .B(new_new_n182_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n188_), .B(i_7_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n189_), .B(i_4_), .Y(new_new_n190_));
  NAi21      g168(.An(i_12_), .B(i_7_), .Y(new_new_n191_));
  NA3        g169(.A(i_13_), .B(new_new_n175_), .C(i_10_), .Y(new_new_n192_));
  NO2        g170(.A(new_new_n192_), .B(new_new_n191_), .Y(new_new_n193_));
  NA2        g171(.A(i_0_), .B(i_5_), .Y(new_new_n194_));
  OAI220     g172(.A0(new_new_n84_), .A1(new_new_n173_), .B0(new_new_n167_), .B1(new_new_n135_), .Y(new_new_n195_));
  NAi31      g173(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n36_), .B(i_13_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n198_));
  NO2        g176(.A(new_new_n46_), .B(new_new_n61_), .Y(new_new_n199_));
  NA3        g177(.A(new_new_n199_), .B(new_new_n198_), .C(new_new_n197_), .Y(new_new_n200_));
  INV        g178(.A(i_13_), .Y(new_new_n201_));
  NO2        g179(.A(i_12_), .B(new_new_n201_), .Y(new_new_n202_));
  NA3        g180(.A(new_new_n202_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n203_));
  OAI210     g181(.A0(new_new_n200_), .A1(new_new_n196_), .B0(new_new_n203_), .Y(new_new_n204_));
  AOI220     g182(.A0(new_new_n204_), .A1(new_new_n144_), .B0(new_new_n195_), .B1(new_new_n193_), .Y(new_new_n205_));
  NO2        g183(.A(i_12_), .B(new_new_n37_), .Y(new_new_n206_));
  OR2        g184(.A(i_8_), .B(i_7_), .Y(new_new_n207_));
  INV        g185(.A(i_12_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n44_), .B(new_new_n208_), .Y(new_new_n209_));
  NO3        g187(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n210_));
  NA2        g188(.A(i_2_), .B(i_1_), .Y(new_new_n211_));
  NO3        g189(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n212_));
  NAi21      g190(.An(i_4_), .B(i_3_), .Y(new_new_n213_));
  NO2        g191(.A(i_0_), .B(i_6_), .Y(new_new_n214_));
  NOi41      g192(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n211_), .B(new_new_n168_), .Y(new_new_n216_));
  NO2        g194(.A(i_11_), .B(new_new_n201_), .Y(new_new_n217_));
  NOi21      g195(.An(i_1_), .B(i_6_), .Y(new_new_n218_));
  NAi21      g196(.An(i_3_), .B(i_7_), .Y(new_new_n219_));
  NA2        g197(.A(new_new_n208_), .B(i_9_), .Y(new_new_n220_));
  OR4        g198(.A(new_new_n220_), .B(new_new_n219_), .C(new_new_n218_), .D(new_new_n169_), .Y(new_new_n221_));
  NA2        g199(.A(new_new_n71_), .B(i_5_), .Y(new_new_n222_));
  NA2        g200(.A(i_3_), .B(i_9_), .Y(new_new_n223_));
  NAi21      g201(.An(i_7_), .B(i_10_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n225_));
  NA3        g203(.A(new_new_n225_), .B(new_new_n222_), .C(new_new_n62_), .Y(new_new_n226_));
  NA2        g204(.A(new_new_n226_), .B(new_new_n221_), .Y(new_new_n227_));
  INV        g205(.A(new_new_n145_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n208_), .B(i_13_), .Y(new_new_n229_));
  NO2        g207(.A(new_new_n229_), .B(new_new_n73_), .Y(new_new_n230_));
  AOI220     g208(.A0(new_new_n230_), .A1(new_new_n228_), .B0(new_new_n227_), .B1(new_new_n217_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n207_), .B(new_new_n37_), .Y(new_new_n232_));
  NA2        g210(.A(i_12_), .B(i_6_), .Y(new_new_n233_));
  OR2        g211(.A(i_13_), .B(i_9_), .Y(new_new_n234_));
  NO3        g212(.A(new_new_n234_), .B(new_new_n233_), .C(new_new_n48_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n213_), .B(i_2_), .Y(new_new_n236_));
  NA3        g214(.A(new_new_n236_), .B(new_new_n235_), .C(new_new_n44_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n217_), .B(i_9_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n222_), .B(new_new_n62_), .Y(new_new_n239_));
  OAI210     g217(.A0(new_new_n239_), .A1(new_new_n238_), .B0(new_new_n237_), .Y(new_new_n240_));
  NO3        g218(.A(i_11_), .B(new_new_n201_), .C(new_new_n25_), .Y(new_new_n241_));
  NO2        g219(.A(new_new_n219_), .B(i_8_), .Y(new_new_n242_));
  NO2        g220(.A(i_6_), .B(new_new_n48_), .Y(new_new_n243_));
  NA2        g221(.A(new_new_n240_), .B(new_new_n232_), .Y(new_new_n244_));
  NA3        g222(.A(new_new_n244_), .B(new_new_n231_), .C(new_new_n205_), .Y(new_new_n245_));
  NO3        g223(.A(i_12_), .B(new_new_n201_), .C(new_new_n37_), .Y(new_new_n246_));
  INV        g224(.A(new_new_n246_), .Y(new_new_n247_));
  NO3        g225(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n248_));
  NO2        g226(.A(new_new_n211_), .B(i_0_), .Y(new_new_n249_));
  AOI220     g227(.A0(new_new_n249_), .A1(i_8_), .B0(new_new_n248_), .B1(new_new_n144_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n243_), .B(new_new_n26_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n251_), .B(new_new_n250_), .Y(new_new_n252_));
  INV        g230(.A(new_new_n252_), .Y(new_new_n253_));
  NO2        g231(.A(i_3_), .B(i_10_), .Y(new_new_n254_));
  NO2        g232(.A(i_2_), .B(new_new_n102_), .Y(new_new_n255_));
  NA2        g233(.A(i_1_), .B(new_new_n36_), .Y(new_new_n256_));
  AN2        g234(.A(i_3_), .B(i_10_), .Y(new_new_n257_));
  NO2        g235(.A(i_5_), .B(new_new_n37_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n253_), .B(new_new_n247_), .Y(new_new_n260_));
  NO3        g238(.A(new_new_n260_), .B(new_new_n245_), .C(new_new_n190_), .Y(new_new_n261_));
  NO3        g239(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n262_));
  NO3        g240(.A(i_6_), .B(new_new_n175_), .C(i_7_), .Y(new_new_n263_));
  NO2        g241(.A(i_2_), .B(i_3_), .Y(new_new_n264_));
  OR2        g242(.A(i_0_), .B(i_5_), .Y(new_new_n265_));
  NA2        g243(.A(new_new_n194_), .B(new_new_n265_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n155_), .B(new_new_n46_), .Y(new_new_n267_));
  NO2        g245(.A(i_12_), .B(i_10_), .Y(new_new_n268_));
  NOi21      g246(.An(i_5_), .B(i_0_), .Y(new_new_n269_));
  NO2        g247(.A(i_2_), .B(new_new_n102_), .Y(new_new_n270_));
  NO4        g248(.A(new_new_n270_), .B(new_new_n256_), .C(new_new_n269_), .D(new_new_n130_), .Y(new_new_n271_));
  NA4        g249(.A(new_new_n82_), .B(new_new_n36_), .C(new_new_n84_), .D(i_8_), .Y(new_new_n272_));
  NA2        g250(.A(new_new_n271_), .B(new_new_n268_), .Y(new_new_n273_));
  NO2        g251(.A(i_6_), .B(i_8_), .Y(new_new_n274_));
  NOi21      g252(.An(i_0_), .B(i_2_), .Y(new_new_n275_));
  AN2        g253(.A(new_new_n275_), .B(new_new_n274_), .Y(new_new_n276_));
  NO2        g254(.A(i_1_), .B(i_7_), .Y(new_new_n277_));
  NA3        g255(.A(new_new_n218_), .B(new_new_n255_), .C(new_new_n175_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n278_), .B(new_new_n266_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n279_), .B(i_3_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n175_), .B(i_9_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n281_), .B(new_new_n183_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n282_), .B(new_new_n46_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n283_), .B(new_new_n252_), .Y(new_new_n284_));
  AOI210     g262(.A0(new_new_n284_), .A1(new_new_n280_), .B0(new_new_n160_), .Y(new_new_n285_));
  AOI210     g263(.A0(new_new_n871_), .A1(new_new_n262_), .B0(new_new_n285_), .Y(new_new_n286_));
  NOi32      g264(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n287_));
  INV        g265(.A(new_new_n287_), .Y(new_new_n288_));
  NAi21      g266(.An(i_0_), .B(i_6_), .Y(new_new_n289_));
  NAi21      g267(.An(i_1_), .B(i_5_), .Y(new_new_n290_));
  NAi41      g268(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n291_));
  OAI220     g269(.A0(new_new_n291_), .A1(new_new_n290_), .B0(new_new_n196_), .B1(new_new_n157_), .Y(new_new_n292_));
  AOI210     g270(.A0(new_new_n291_), .A1(new_new_n157_), .B0(new_new_n155_), .Y(new_new_n293_));
  NOi32      g271(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n294_));
  NAi21      g272(.An(i_6_), .B(i_1_), .Y(new_new_n295_));
  NA3        g273(.A(new_new_n295_), .B(new_new_n294_), .C(new_new_n46_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n296_), .B(i_0_), .Y(new_new_n297_));
  OR3        g275(.A(new_new_n297_), .B(new_new_n293_), .C(new_new_n292_), .Y(new_new_n298_));
  NO2        g276(.A(i_1_), .B(new_new_n102_), .Y(new_new_n299_));
  NAi21      g277(.An(i_3_), .B(i_4_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n300_), .B(i_9_), .Y(new_new_n301_));
  AN2        g279(.A(i_6_), .B(i_7_), .Y(new_new_n302_));
  OAI210     g280(.A0(new_new_n302_), .A1(new_new_n299_), .B0(new_new_n301_), .Y(new_new_n303_));
  NA2        g281(.A(i_2_), .B(i_7_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n300_), .B(i_10_), .Y(new_new_n305_));
  NA3        g283(.A(new_new_n305_), .B(new_new_n304_), .C(new_new_n214_), .Y(new_new_n306_));
  AOI210     g284(.A0(new_new_n306_), .A1(new_new_n303_), .B0(new_new_n169_), .Y(new_new_n307_));
  AOI210     g285(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n308_));
  OAI210     g286(.A0(new_new_n308_), .A1(new_new_n172_), .B0(new_new_n305_), .Y(new_new_n309_));
  AOI220     g287(.A0(new_new_n305_), .A1(new_new_n277_), .B0(new_new_n210_), .B1(new_new_n172_), .Y(new_new_n310_));
  AOI210     g288(.A0(new_new_n310_), .A1(new_new_n309_), .B0(i_5_), .Y(new_new_n311_));
  NO3        g289(.A(new_new_n311_), .B(new_new_n307_), .C(new_new_n298_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n312_), .B(new_new_n288_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n314_));
  AN2        g292(.A(i_12_), .B(i_5_), .Y(new_new_n315_));
  NO2        g293(.A(i_4_), .B(new_new_n26_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(new_new_n315_), .Y(new_new_n317_));
  NO2        g295(.A(i_11_), .B(i_6_), .Y(new_new_n318_));
  NA3        g296(.A(new_new_n318_), .B(new_new_n267_), .C(new_new_n201_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n319_), .B(new_new_n317_), .Y(new_new_n320_));
  NO2        g298(.A(i_5_), .B(i_10_), .Y(new_new_n321_));
  NA2        g299(.A(new_new_n321_), .B(new_new_n236_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n146_), .B(new_new_n45_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n323_), .B(new_new_n322_), .Y(new_new_n324_));
  OAI210     g302(.A0(new_new_n324_), .A1(new_new_n320_), .B0(new_new_n314_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n152_), .B(new_new_n84_), .Y(new_new_n327_));
  OAI210     g305(.A0(new_new_n327_), .A1(new_new_n320_), .B0(new_new_n326_), .Y(new_new_n328_));
  NO3        g306(.A(new_new_n84_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n329_));
  NA3        g307(.A(new_new_n254_), .B(new_new_n91_), .C(new_new_n73_), .Y(new_new_n330_));
  NO2        g308(.A(i_11_), .B(i_12_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n331_), .B(new_new_n36_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n330_), .B(new_new_n332_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n321_), .B(new_new_n208_), .Y(new_new_n334_));
  NAi21      g312(.An(i_13_), .B(i_0_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n335_), .B(new_new_n211_), .Y(new_new_n336_));
  NA2        g314(.A(new_new_n333_), .B(new_new_n336_), .Y(new_new_n337_));
  NA3        g315(.A(new_new_n337_), .B(new_new_n328_), .C(new_new_n325_), .Y(new_new_n338_));
  NA2        g316(.A(new_new_n44_), .B(new_new_n201_), .Y(new_new_n339_));
  NO3        g317(.A(i_1_), .B(i_12_), .C(new_new_n84_), .Y(new_new_n340_));
  NO2        g318(.A(i_0_), .B(i_11_), .Y(new_new_n341_));
  NOi21      g319(.An(i_2_), .B(i_12_), .Y(new_new_n342_));
  NAi21      g320(.An(i_9_), .B(i_4_), .Y(new_new_n343_));
  OR2        g321(.A(i_13_), .B(i_10_), .Y(new_new_n344_));
  NO3        g322(.A(new_new_n344_), .B(new_new_n119_), .C(new_new_n343_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n163_), .B(new_new_n125_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n102_), .B(new_new_n25_), .Y(new_new_n347_));
  NO2        g325(.A(new_new_n168_), .B(new_new_n84_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n175_), .B(i_10_), .Y(new_new_n349_));
  NA3        g327(.A(new_new_n222_), .B(new_new_n62_), .C(i_2_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n350_), .B(new_new_n349_), .Y(new_new_n351_));
  NO2        g329(.A(i_3_), .B(new_new_n48_), .Y(new_new_n352_));
  NA3        g330(.A(new_new_n277_), .B(new_new_n276_), .C(new_new_n352_), .Y(new_new_n353_));
  NA2        g331(.A(new_new_n263_), .B(new_new_n266_), .Y(new_new_n354_));
  OAI210     g332(.A0(new_new_n354_), .A1(new_new_n173_), .B0(new_new_n353_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n355_), .B(new_new_n351_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n356_), .B(new_new_n238_), .Y(new_new_n357_));
  NO3        g335(.A(new_new_n357_), .B(new_new_n338_), .C(new_new_n313_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n71_), .B(i_13_), .Y(new_new_n359_));
  NO2        g337(.A(i_10_), .B(i_9_), .Y(new_new_n360_));
  NAi21      g338(.An(i_12_), .B(i_8_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n361_), .B(i_3_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n46_), .B(i_4_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n363_), .B(new_new_n105_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n364_), .B(new_new_n182_), .Y(new_new_n365_));
  NA2        g343(.A(new_new_n259_), .B(i_0_), .Y(new_new_n366_));
  NO3        g344(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n367_));
  NA2        g345(.A(new_new_n233_), .B(new_new_n98_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n368_), .B(new_new_n367_), .Y(new_new_n369_));
  NA2        g347(.A(i_8_), .B(i_9_), .Y(new_new_n370_));
  AOI210     g348(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n371_));
  OR2        g349(.A(new_new_n371_), .B(new_new_n370_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n246_), .B(new_new_n183_), .Y(new_new_n373_));
  OAI220     g351(.A0(new_new_n373_), .A1(new_new_n372_), .B0(new_new_n369_), .B1(new_new_n366_), .Y(new_new_n374_));
  NA2        g352(.A(new_new_n217_), .B(new_new_n258_), .Y(new_new_n375_));
  NO3        g353(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n376_));
  INV        g354(.A(new_new_n376_), .Y(new_new_n377_));
  NA3        g355(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n378_));
  NA4        g356(.A(new_new_n147_), .B(new_new_n117_), .C(new_new_n78_), .D(new_new_n23_), .Y(new_new_n379_));
  OAI220     g357(.A0(new_new_n379_), .A1(new_new_n378_), .B0(new_new_n377_), .B1(new_new_n375_), .Y(new_new_n380_));
  NO3        g358(.A(new_new_n380_), .B(new_new_n374_), .C(new_new_n365_), .Y(new_new_n381_));
  OR2        g359(.A(new_new_n282_), .B(new_new_n102_), .Y(new_new_n382_));
  OR2        g360(.A(new_new_n382_), .B(new_new_n160_), .Y(new_new_n383_));
  NA2        g361(.A(new_new_n97_), .B(i_13_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n348_), .B(new_new_n314_), .Y(new_new_n385_));
  NO2        g363(.A(i_2_), .B(i_13_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n385_), .B(new_new_n384_), .Y(new_new_n387_));
  NO3        g365(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n388_));
  NO2        g366(.A(i_6_), .B(i_7_), .Y(new_new_n389_));
  NO2        g367(.A(i_11_), .B(i_1_), .Y(new_new_n390_));
  OR2        g368(.A(i_11_), .B(i_8_), .Y(new_new_n391_));
  NOi21      g369(.An(i_2_), .B(i_7_), .Y(new_new_n392_));
  NO2        g370(.A(i_6_), .B(i_10_), .Y(new_new_n393_));
  NA3        g371(.A(new_new_n215_), .B(new_new_n162_), .C(new_new_n134_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n155_), .B(i_3_), .Y(new_new_n396_));
  NAi31      g374(.An(new_new_n395_), .B(new_new_n396_), .C(new_new_n202_), .Y(new_new_n397_));
  NA3        g375(.A(new_new_n326_), .B(new_new_n166_), .C(new_new_n151_), .Y(new_new_n398_));
  NA3        g376(.A(new_new_n398_), .B(new_new_n397_), .C(new_new_n394_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(new_new_n387_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n367_), .B(new_new_n315_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n376_), .B(new_new_n321_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n402_), .B(new_new_n200_), .Y(new_new_n403_));
  NAi21      g381(.An(new_new_n192_), .B(new_new_n331_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n277_), .B(new_new_n194_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n405_), .B(new_new_n404_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n27_), .B(i_10_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n262_), .B(new_new_n210_), .Y(new_new_n408_));
  OAI220     g386(.A0(new_new_n408_), .A1(new_new_n350_), .B0(new_new_n407_), .B1(new_new_n384_), .Y(new_new_n409_));
  NO3        g387(.A(new_new_n409_), .B(new_new_n406_), .C(new_new_n403_), .Y(new_new_n410_));
  NA4        g388(.A(new_new_n410_), .B(new_new_n400_), .C(new_new_n383_), .D(new_new_n381_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n124_), .B(new_new_n113_), .Y(new_new_n412_));
  AN2        g390(.A(new_new_n412_), .B(new_new_n367_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n413_), .B(new_new_n259_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n287_), .B(new_new_n71_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n302_), .B(new_new_n294_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n36_), .B(i_8_), .Y(new_new_n417_));
  AOI210     g395(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n345_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n222_), .B(new_new_n62_), .Y(new_new_n419_));
  OAI210     g397(.A0(i_8_), .A1(new_new_n419_), .B0(new_new_n136_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n420_), .B(new_new_n346_), .Y(new_new_n421_));
  NA3        g399(.A(new_new_n421_), .B(new_new_n418_), .C(new_new_n414_), .Y(new_new_n422_));
  NO2        g400(.A(i_12_), .B(new_new_n175_), .Y(new_new_n423_));
  NO2        g401(.A(i_8_), .B(i_7_), .Y(new_new_n424_));
  AOI220     g402(.A0(new_new_n348_), .A1(new_new_n267_), .B0(new_new_n216_), .B1(new_new_n214_), .Y(new_new_n425_));
  OAI220     g403(.A0(new_new_n425_), .A1(new_new_n229_), .B0(new_new_n384_), .B1(new_new_n135_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n426_), .B(new_new_n232_), .Y(new_new_n427_));
  NA3        g405(.A(new_new_n257_), .B(new_new_n164_), .C(new_new_n97_), .Y(new_new_n428_));
  NO2        g406(.A(new_new_n197_), .B(new_new_n44_), .Y(new_new_n429_));
  NO2        g407(.A(new_new_n155_), .B(i_5_), .Y(new_new_n430_));
  NA3        g408(.A(new_new_n430_), .B(new_new_n339_), .C(new_new_n264_), .Y(new_new_n431_));
  OAI210     g409(.A0(new_new_n431_), .A1(new_new_n429_), .B0(new_new_n428_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n432_), .B(new_new_n376_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n433_), .B(new_new_n427_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n199_), .B(new_new_n198_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n360_), .B(new_new_n197_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n435_), .B(new_new_n436_), .Y(new_new_n437_));
  AOI210     g415(.A0(new_new_n295_), .A1(new_new_n46_), .B0(new_new_n299_), .Y(new_new_n438_));
  NA2        g416(.A(i_0_), .B(new_new_n48_), .Y(new_new_n439_));
  NA3        g417(.A(new_new_n423_), .B(new_new_n241_), .C(new_new_n439_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n438_), .B(new_new_n440_), .Y(new_new_n441_));
  NO2        g419(.A(new_new_n441_), .B(new_new_n437_), .Y(new_new_n442_));
  NO4        g420(.A(new_new_n218_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n443_));
  NO3        g421(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n207_), .B(new_new_n36_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n344_), .B(i_1_), .Y(new_new_n446_));
  NOi31      g424(.An(new_new_n446_), .B(new_new_n368_), .C(new_new_n71_), .Y(new_new_n447_));
  NOi21      g425(.An(i_10_), .B(i_6_), .Y(new_new_n448_));
  NO2        g426(.A(new_new_n84_), .B(new_new_n25_), .Y(new_new_n449_));
  AOI220     g427(.A0(new_new_n246_), .A1(new_new_n449_), .B0(new_new_n241_), .B1(new_new_n448_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n450_), .B(new_new_n366_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n178_), .B(new_new_n37_), .Y(new_new_n453_));
  NOi31      g431(.An(new_new_n148_), .B(new_new_n453_), .C(new_new_n272_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n454_), .B(new_new_n451_), .Y(new_new_n455_));
  NO2        g433(.A(new_new_n415_), .B(new_new_n310_), .Y(new_new_n456_));
  INV        g434(.A(new_new_n264_), .Y(new_new_n457_));
  NO2        g435(.A(i_12_), .B(new_new_n84_), .Y(new_new_n458_));
  NA3        g436(.A(new_new_n458_), .B(new_new_n241_), .C(new_new_n439_), .Y(new_new_n459_));
  NA3        g437(.A(new_new_n318_), .B(new_new_n246_), .C(new_new_n194_), .Y(new_new_n460_));
  AOI210     g438(.A0(new_new_n460_), .A1(new_new_n459_), .B0(new_new_n457_), .Y(new_new_n461_));
  OR2        g439(.A(i_2_), .B(i_5_), .Y(new_new_n462_));
  OR2        g440(.A(new_new_n462_), .B(i_6_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n304_), .B(new_new_n214_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n464_), .B(new_new_n404_), .Y(new_new_n465_));
  NO3        g443(.A(new_new_n465_), .B(new_new_n461_), .C(new_new_n456_), .Y(new_new_n466_));
  NA3        g444(.A(new_new_n466_), .B(new_new_n455_), .C(new_new_n442_), .Y(new_new_n467_));
  NO4        g445(.A(new_new_n467_), .B(new_new_n434_), .C(new_new_n422_), .D(new_new_n411_), .Y(new_new_n468_));
  NA4        g446(.A(new_new_n468_), .B(new_new_n358_), .C(new_new_n286_), .D(new_new_n261_), .Y(ori7));
  NO2        g447(.A(new_new_n93_), .B(new_new_n54_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n109_), .B(new_new_n90_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n316_), .B(new_new_n471_), .Y(new_new_n472_));
  NA2        g450(.A(new_new_n393_), .B(new_new_n82_), .Y(new_new_n473_));
  NA2        g451(.A(i_11_), .B(new_new_n175_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n146_), .B(new_new_n474_), .Y(new_new_n475_));
  OAI210     g453(.A0(new_new_n475_), .A1(new_new_n473_), .B0(new_new_n472_), .Y(new_new_n476_));
  NO2        g454(.A(new_new_n208_), .B(i_4_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n477_), .B(i_8_), .Y(new_new_n478_));
  NA2        g456(.A(i_2_), .B(new_new_n84_), .Y(new_new_n479_));
  OAI210     g457(.A0(new_new_n87_), .A1(new_new_n180_), .B0(new_new_n181_), .Y(new_new_n480_));
  NO2        g458(.A(i_7_), .B(new_new_n37_), .Y(new_new_n481_));
  NA2        g459(.A(i_4_), .B(i_8_), .Y(new_new_n482_));
  AOI210     g460(.A0(new_new_n482_), .A1(new_new_n257_), .B0(new_new_n481_), .Y(new_new_n483_));
  OAI220     g461(.A0(new_new_n483_), .A1(new_new_n479_), .B0(new_new_n480_), .B1(i_13_), .Y(new_new_n484_));
  NO3        g462(.A(new_new_n484_), .B(new_new_n476_), .C(new_new_n470_), .Y(new_new_n485_));
  AOI210     g463(.A0(new_new_n130_), .A1(new_new_n60_), .B0(i_10_), .Y(new_new_n486_));
  AOI210     g464(.A0(new_new_n486_), .A1(new_new_n208_), .B0(new_new_n159_), .Y(new_new_n487_));
  OR2        g465(.A(i_6_), .B(i_10_), .Y(new_new_n488_));
  OR3        g466(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n489_));
  INV        g467(.A(new_new_n179_), .Y(new_new_n490_));
  OR2        g468(.A(new_new_n487_), .B(new_new_n234_), .Y(new_new_n491_));
  AOI210     g469(.A0(new_new_n491_), .A1(new_new_n485_), .B0(new_new_n61_), .Y(new_new_n492_));
  NOi21      g470(.An(i_11_), .B(i_7_), .Y(new_new_n493_));
  AO210      g471(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n494_), .B(new_new_n493_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n495_), .B(new_new_n185_), .Y(new_new_n496_));
  NA3        g474(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n497_));
  NAi31      g475(.An(new_new_n497_), .B(new_new_n191_), .C(i_11_), .Y(new_new_n498_));
  AOI210     g476(.A0(new_new_n498_), .A1(new_new_n496_), .B0(new_new_n61_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n86_), .B(new_new_n61_), .Y(new_new_n500_));
  AO210      g478(.A0(new_new_n500_), .A1(new_new_n310_), .B0(new_new_n41_), .Y(new_new_n501_));
  NO3        g479(.A(new_new_n224_), .B(new_new_n186_), .C(new_new_n474_), .Y(new_new_n502_));
  OAI210     g480(.A0(new_new_n502_), .A1(new_new_n202_), .B0(new_new_n61_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n342_), .B(new_new_n31_), .Y(new_new_n504_));
  OR2        g482(.A(new_new_n186_), .B(new_new_n109_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n505_), .B(new_new_n504_), .Y(new_new_n506_));
  NO2        g484(.A(new_new_n61_), .B(i_9_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(i_4_), .Y(new_new_n508_));
  NA2        g486(.A(new_new_n508_), .B(new_new_n506_), .Y(new_new_n509_));
  NO2        g487(.A(i_1_), .B(i_12_), .Y(new_new_n510_));
  NA3        g488(.A(new_new_n510_), .B(new_new_n111_), .C(new_new_n24_), .Y(new_new_n511_));
  BUFFER     g489(.A(new_new_n511_), .Y(new_new_n512_));
  NA4        g490(.A(new_new_n512_), .B(new_new_n509_), .C(new_new_n503_), .D(new_new_n501_), .Y(new_new_n513_));
  OAI210     g491(.A0(new_new_n513_), .A1(new_new_n499_), .B0(i_6_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n208_), .B(new_new_n84_), .Y(new_new_n515_));
  NO2        g493(.A(new_new_n515_), .B(i_11_), .Y(new_new_n516_));
  INV        g494(.A(new_new_n369_), .Y(new_new_n517_));
  NO3        g495(.A(new_new_n488_), .B(new_new_n207_), .C(new_new_n23_), .Y(new_new_n518_));
  AOI210     g496(.A0(i_1_), .A1(new_new_n225_), .B0(new_new_n518_), .Y(new_new_n519_));
  NO2        g497(.A(new_new_n519_), .B(new_new_n44_), .Y(new_new_n520_));
  NA3        g498(.A(new_new_n424_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n521_));
  INV        g499(.A(i_2_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n140_), .B(i_9_), .Y(new_new_n523_));
  NA3        g501(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n46_), .B(i_1_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n523_), .B(new_new_n522_), .Y(new_new_n526_));
  NA3        g504(.A(new_new_n507_), .B(new_new_n264_), .C(i_6_), .Y(new_new_n527_));
  NO2        g505(.A(new_new_n527_), .B(new_new_n23_), .Y(new_new_n528_));
  AOI210     g506(.A0(new_new_n390_), .A1(new_new_n347_), .B0(new_new_n212_), .Y(new_new_n529_));
  NO2        g507(.A(new_new_n529_), .B(new_new_n479_), .Y(new_new_n530_));
  NAi21      g508(.An(new_new_n521_), .B(new_new_n92_), .Y(new_new_n531_));
  NA2        g509(.A(new_new_n525_), .B(new_new_n233_), .Y(new_new_n532_));
  NO2        g510(.A(i_11_), .B(new_new_n37_), .Y(new_new_n533_));
  NA2        g511(.A(new_new_n533_), .B(new_new_n24_), .Y(new_new_n534_));
  OAI210     g512(.A0(new_new_n534_), .A1(new_new_n532_), .B0(new_new_n531_), .Y(new_new_n535_));
  OR4        g513(.A(new_new_n535_), .B(new_new_n530_), .C(new_new_n528_), .D(new_new_n526_), .Y(new_new_n536_));
  NO3        g514(.A(new_new_n536_), .B(new_new_n520_), .C(new_new_n517_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n208_), .B(new_new_n102_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n538_), .B(new_new_n493_), .Y(new_new_n539_));
  NA2        g517(.A(new_new_n539_), .B(i_1_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n540_), .B(new_new_n489_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n343_), .B(new_new_n84_), .Y(new_new_n542_));
  NA2        g520(.A(new_new_n541_), .B(new_new_n46_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n207_), .B(new_new_n44_), .Y(new_new_n544_));
  NO3        g522(.A(new_new_n544_), .B(new_new_n259_), .C(new_new_n209_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n119_), .B(new_new_n37_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n546_), .B(i_6_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n84_), .B(i_9_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n548_), .B(new_new_n61_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n549_), .B(new_new_n510_), .Y(new_new_n550_));
  NO4        g528(.A(new_new_n550_), .B(new_new_n547_), .C(new_new_n545_), .D(i_4_), .Y(new_new_n551_));
  NA2        g529(.A(i_1_), .B(i_3_), .Y(new_new_n552_));
  INV        g530(.A(new_new_n551_), .Y(new_new_n553_));
  NA4        g531(.A(new_new_n553_), .B(new_new_n543_), .C(new_new_n537_), .D(new_new_n514_), .Y(new_new_n554_));
  NO3        g532(.A(new_new_n391_), .B(i_3_), .C(i_7_), .Y(new_new_n555_));
  NOi21      g533(.An(new_new_n555_), .B(i_10_), .Y(new_new_n556_));
  OA210      g534(.A0(new_new_n556_), .A1(new_new_n215_), .B0(new_new_n84_), .Y(new_new_n557_));
  NA3        g535(.A(new_new_n393_), .B(new_new_n417_), .C(new_new_n46_), .Y(new_new_n558_));
  NO3        g536(.A(new_new_n392_), .B(new_new_n482_), .C(new_new_n84_), .Y(new_new_n559_));
  NA2        g537(.A(new_new_n559_), .B(new_new_n25_), .Y(new_new_n560_));
  NA3        g538(.A(new_new_n159_), .B(new_new_n82_), .C(new_new_n84_), .Y(new_new_n561_));
  NA3        g539(.A(new_new_n561_), .B(new_new_n560_), .C(new_new_n558_), .Y(new_new_n562_));
  OAI210     g540(.A0(new_new_n562_), .A1(new_new_n557_), .B0(i_1_), .Y(new_new_n563_));
  AOI210     g541(.A0(new_new_n233_), .A1(new_new_n98_), .B0(i_1_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n300_), .B(i_2_), .Y(new_new_n565_));
  NA2        g543(.A(new_new_n565_), .B(new_new_n564_), .Y(new_new_n566_));
  OAI210     g544(.A0(new_new_n527_), .A1(new_new_n361_), .B0(new_new_n566_), .Y(new_new_n567_));
  INV        g545(.A(new_new_n567_), .Y(new_new_n568_));
  AOI210     g546(.A0(new_new_n568_), .A1(new_new_n563_), .B0(i_13_), .Y(new_new_n569_));
  OR2        g547(.A(i_11_), .B(i_7_), .Y(new_new_n570_));
  NA3        g548(.A(new_new_n570_), .B(new_new_n107_), .C(new_new_n140_), .Y(new_new_n571_));
  AOI220     g549(.A0(new_new_n386_), .A1(new_new_n159_), .B0(new_new_n363_), .B1(new_new_n140_), .Y(new_new_n572_));
  OAI210     g550(.A0(new_new_n572_), .A1(new_new_n44_), .B0(new_new_n571_), .Y(new_new_n573_));
  NO2        g551(.A(new_new_n54_), .B(i_12_), .Y(new_new_n574_));
  NO2        g552(.A(new_new_n392_), .B(new_new_n24_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n575_), .B(new_new_n542_), .Y(new_new_n576_));
  OAI220     g554(.A0(new_new_n576_), .A1(new_new_n41_), .B0(new_new_n870_), .B1(new_new_n93_), .Y(new_new_n577_));
  AOI210     g555(.A0(new_new_n573_), .A1(new_new_n274_), .B0(new_new_n577_), .Y(new_new_n578_));
  INV        g556(.A(new_new_n116_), .Y(new_new_n579_));
  AOI220     g557(.A0(new_new_n579_), .A1(new_new_n70_), .B0(new_new_n318_), .B1(new_new_n525_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n580_), .B(new_new_n213_), .Y(new_new_n581_));
  NA2        g559(.A(new_new_n129_), .B(i_13_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n524_), .B(new_new_n116_), .Y(new_new_n583_));
  INV        g561(.A(new_new_n583_), .Y(new_new_n584_));
  OAI220     g562(.A0(new_new_n584_), .A1(new_new_n69_), .B0(new_new_n582_), .B1(new_new_n564_), .Y(new_new_n585_));
  NO3        g563(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n102_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n26_), .B(new_new_n175_), .Y(new_new_n587_));
  INV        g565(.A(i_7_), .Y(new_new_n588_));
  AOI220     g566(.A0(new_new_n318_), .A1(new_new_n525_), .B0(new_new_n92_), .B1(new_new_n103_), .Y(new_new_n589_));
  OAI220     g567(.A0(new_new_n589_), .A1(new_new_n478_), .B0(new_new_n872_), .B1(new_new_n490_), .Y(new_new_n590_));
  NO3        g568(.A(new_new_n590_), .B(new_new_n585_), .C(new_new_n581_), .Y(new_new_n591_));
  OR2        g569(.A(i_11_), .B(i_6_), .Y(new_new_n592_));
  NA3        g570(.A(new_new_n477_), .B(new_new_n587_), .C(i_7_), .Y(new_new_n593_));
  AOI210     g571(.A0(new_new_n593_), .A1(new_new_n584_), .B0(new_new_n592_), .Y(new_new_n594_));
  NA3        g572(.A(new_new_n342_), .B(new_new_n481_), .C(new_new_n98_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n516_), .B(i_13_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n103_), .B(new_new_n587_), .Y(new_new_n597_));
  NAi21      g575(.An(i_11_), .B(i_12_), .Y(new_new_n598_));
  NOi41      g576(.An(new_new_n112_), .B(new_new_n598_), .C(i_13_), .D(new_new_n84_), .Y(new_new_n599_));
  NO3        g577(.A(new_new_n392_), .B(new_new_n458_), .C(new_new_n482_), .Y(new_new_n600_));
  AOI220     g578(.A0(new_new_n600_), .A1(new_new_n262_), .B0(new_new_n599_), .B1(new_new_n597_), .Y(new_new_n601_));
  NA3        g579(.A(new_new_n601_), .B(new_new_n596_), .C(new_new_n595_), .Y(new_new_n602_));
  OAI210     g580(.A0(new_new_n602_), .A1(new_new_n594_), .B0(new_new_n61_), .Y(new_new_n603_));
  NO2        g581(.A(i_2_), .B(i_12_), .Y(new_new_n604_));
  NA2        g582(.A(new_new_n299_), .B(new_new_n604_), .Y(new_new_n605_));
  INV        g583(.A(new_new_n605_), .Y(new_new_n606_));
  NA3        g584(.A(new_new_n606_), .B(new_new_n45_), .C(new_new_n201_), .Y(new_new_n607_));
  NA4        g585(.A(new_new_n607_), .B(new_new_n603_), .C(new_new_n591_), .D(new_new_n578_), .Y(new_new_n608_));
  OR4        g586(.A(new_new_n608_), .B(new_new_n569_), .C(new_new_n554_), .D(new_new_n492_), .Y(ori5));
  NA2        g587(.A(new_new_n539_), .B(new_new_n236_), .Y(new_new_n610_));
  AN2        g588(.A(new_new_n24_), .B(i_10_), .Y(new_new_n611_));
  NA3        g589(.A(new_new_n611_), .B(new_new_n604_), .C(new_new_n109_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n478_), .B(i_11_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n87_), .B(new_new_n613_), .Y(new_new_n614_));
  NA3        g592(.A(new_new_n614_), .B(new_new_n612_), .C(new_new_n610_), .Y(new_new_n615_));
  NO3        g593(.A(i_11_), .B(new_new_n208_), .C(i_13_), .Y(new_new_n616_));
  NO2        g594(.A(new_new_n126_), .B(new_new_n23_), .Y(new_new_n617_));
  NA2        g595(.A(i_12_), .B(i_8_), .Y(new_new_n618_));
  OAI210     g596(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n618_), .Y(new_new_n619_));
  INV        g597(.A(new_new_n360_), .Y(new_new_n620_));
  AOI220     g598(.A0(new_new_n264_), .A1(new_new_n452_), .B0(new_new_n619_), .B1(new_new_n617_), .Y(new_new_n621_));
  INV        g599(.A(new_new_n621_), .Y(new_new_n622_));
  NO2        g600(.A(new_new_n622_), .B(new_new_n615_), .Y(new_new_n623_));
  INV        g601(.A(new_new_n162_), .Y(new_new_n624_));
  INV        g602(.A(new_new_n215_), .Y(new_new_n625_));
  OAI210     g603(.A0(new_new_n565_), .A1(new_new_n362_), .B0(new_new_n112_), .Y(new_new_n626_));
  AOI210     g604(.A0(new_new_n626_), .A1(new_new_n625_), .B0(new_new_n624_), .Y(new_new_n627_));
  NO2        g605(.A(new_new_n370_), .B(new_new_n26_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n628_), .B(new_new_n347_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n629_), .B(i_2_), .Y(new_new_n630_));
  INV        g608(.A(new_new_n630_), .Y(new_new_n631_));
  AOI210     g609(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n344_), .Y(new_new_n632_));
  AOI210     g610(.A0(new_new_n632_), .A1(new_new_n631_), .B0(new_new_n627_), .Y(new_new_n633_));
  NO2        g611(.A(new_new_n174_), .B(new_new_n127_), .Y(new_new_n634_));
  OAI210     g612(.A0(new_new_n634_), .A1(new_new_n617_), .B0(i_2_), .Y(new_new_n635_));
  INV        g613(.A(new_new_n163_), .Y(new_new_n636_));
  NO3        g614(.A(new_new_n494_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n637_));
  AOI210     g615(.A0(new_new_n636_), .A1(new_new_n87_), .B0(new_new_n637_), .Y(new_new_n638_));
  AOI210     g616(.A0(new_new_n638_), .A1(new_new_n635_), .B0(new_new_n175_), .Y(new_new_n639_));
  OA210      g617(.A0(new_new_n495_), .A1(new_new_n128_), .B0(i_13_), .Y(new_new_n640_));
  NA2        g618(.A(new_new_n179_), .B(new_new_n180_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n153_), .B(new_new_n474_), .Y(new_new_n642_));
  AOI210     g620(.A0(new_new_n642_), .A1(new_new_n641_), .B0(new_new_n304_), .Y(new_new_n643_));
  AOI210     g621(.A0(new_new_n186_), .A1(new_new_n150_), .B0(new_new_n417_), .Y(new_new_n644_));
  NA2        g622(.A(new_new_n644_), .B(new_new_n347_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n103_), .B(new_new_n44_), .Y(new_new_n646_));
  INV        g624(.A(new_new_n255_), .Y(new_new_n647_));
  NA4        g625(.A(new_new_n647_), .B(new_new_n257_), .C(new_new_n126_), .D(new_new_n42_), .Y(new_new_n648_));
  OAI210     g626(.A0(new_new_n648_), .A1(new_new_n646_), .B0(new_new_n645_), .Y(new_new_n649_));
  NO4        g627(.A(new_new_n649_), .B(new_new_n643_), .C(new_new_n640_), .D(new_new_n639_), .Y(new_new_n650_));
  NA2        g628(.A(new_new_n452_), .B(new_new_n28_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n616_), .B(new_new_n242_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n652_), .B(new_new_n651_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n60_), .B(i_12_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n654_), .B(new_new_n128_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n655_), .B(new_new_n474_), .Y(new_new_n656_));
  AOI220     g634(.A0(new_new_n656_), .A1(new_new_n36_), .B0(new_new_n653_), .B1(new_new_n46_), .Y(new_new_n657_));
  NA4        g635(.A(new_new_n657_), .B(new_new_n650_), .C(new_new_n633_), .D(new_new_n623_), .Y(ori6));
  NO2        g636(.A(new_new_n196_), .B(new_new_n395_), .Y(new_new_n659_));
  NO2        g637(.A(i_11_), .B(i_9_), .Y(new_new_n660_));
  INV        g638(.A(new_new_n269_), .Y(new_new_n661_));
  OR2        g639(.A(new_new_n661_), .B(i_12_), .Y(new_new_n662_));
  NA2        g640(.A(new_new_n305_), .B(new_new_n277_), .Y(new_new_n663_));
  NA2        g641(.A(new_new_n458_), .B(new_new_n61_), .Y(new_new_n664_));
  NA2        g642(.A(new_new_n556_), .B(new_new_n69_), .Y(new_new_n665_));
  BUFFER     g643(.A(new_new_n500_), .Y(new_new_n666_));
  NA4        g644(.A(new_new_n666_), .B(new_new_n665_), .C(new_new_n664_), .D(new_new_n663_), .Y(new_new_n667_));
  INV        g645(.A(new_new_n177_), .Y(new_new_n668_));
  AOI220     g646(.A0(new_new_n668_), .A1(new_new_n660_), .B0(new_new_n667_), .B1(new_new_n71_), .Y(new_new_n669_));
  INV        g647(.A(new_new_n268_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n73_), .B(new_new_n133_), .Y(new_new_n671_));
  INV        g649(.A(new_new_n126_), .Y(new_new_n672_));
  NA2        g650(.A(new_new_n672_), .B(new_new_n46_), .Y(new_new_n673_));
  AOI210     g651(.A0(new_new_n673_), .A1(new_new_n671_), .B0(new_new_n670_), .Y(new_new_n674_));
  NO2        g652(.A(new_new_n218_), .B(i_9_), .Y(new_new_n675_));
  NA2        g653(.A(new_new_n675_), .B(new_new_n654_), .Y(new_new_n676_));
  AOI210     g654(.A0(new_new_n676_), .A1(new_new_n416_), .B0(new_new_n169_), .Y(new_new_n677_));
  NO2        g655(.A(new_new_n32_), .B(i_11_), .Y(new_new_n678_));
  NA3        g656(.A(new_new_n678_), .B(new_new_n389_), .C(new_new_n321_), .Y(new_new_n679_));
  NAi32      g657(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n592_), .B(new_new_n680_), .Y(new_new_n681_));
  OAI210     g659(.A0(new_new_n555_), .A1(new_new_n445_), .B0(new_new_n444_), .Y(new_new_n682_));
  NAi31      g660(.An(new_new_n681_), .B(new_new_n682_), .C(new_new_n679_), .Y(new_new_n683_));
  OR3        g661(.A(new_new_n683_), .B(new_new_n677_), .C(new_new_n674_), .Y(new_new_n684_));
  NO2        g662(.A(new_new_n570_), .B(i_2_), .Y(new_new_n685_));
  OR2        g663(.A(new_new_n495_), .B(new_new_n362_), .Y(new_new_n686_));
  NA3        g664(.A(new_new_n686_), .B(new_new_n149_), .C(new_new_n67_), .Y(new_new_n687_));
  AO210      g665(.A0(new_new_n402_), .A1(new_new_n620_), .B0(new_new_n36_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n688_), .B(new_new_n687_), .Y(new_new_n689_));
  OAI210     g667(.A0(new_new_n515_), .A1(i_11_), .B0(new_new_n85_), .Y(new_new_n690_));
  AOI220     g668(.A0(new_new_n690_), .A1(new_new_n444_), .B0(new_new_n659_), .B1(new_new_n588_), .Y(new_new_n691_));
  NA3        g669(.A(new_new_n304_), .B(new_new_n210_), .C(new_new_n149_), .Y(new_new_n692_));
  NA2        g670(.A(new_new_n329_), .B(new_new_n68_), .Y(new_new_n693_));
  NA4        g671(.A(new_new_n693_), .B(new_new_n692_), .C(new_new_n691_), .D(new_new_n480_), .Y(new_new_n694_));
  AO210      g672(.A0(new_new_n417_), .A1(new_new_n46_), .B0(new_new_n86_), .Y(new_new_n695_));
  NA3        g673(.A(new_new_n695_), .B(new_new_n393_), .C(new_new_n194_), .Y(new_new_n696_));
  AOI210     g674(.A0(new_new_n362_), .A1(new_new_n360_), .B0(new_new_n443_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n488_), .B(new_new_n103_), .Y(new_new_n698_));
  OAI210     g676(.A0(new_new_n698_), .A1(new_new_n113_), .B0(new_new_n341_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n214_), .B(new_new_n46_), .Y(new_new_n700_));
  INV        g678(.A(new_new_n463_), .Y(new_new_n701_));
  NA3        g679(.A(new_new_n701_), .B(new_new_n268_), .C(i_7_), .Y(new_new_n702_));
  NA4        g680(.A(new_new_n702_), .B(new_new_n699_), .C(new_new_n697_), .D(new_new_n696_), .Y(new_new_n703_));
  NO4        g681(.A(new_new_n703_), .B(new_new_n694_), .C(new_new_n689_), .D(new_new_n684_), .Y(new_new_n704_));
  NA4        g682(.A(new_new_n704_), .B(new_new_n669_), .C(new_new_n662_), .D(new_new_n312_), .Y(ori3));
  NA2        g683(.A(i_12_), .B(i_10_), .Y(new_new_n706_));
  NO2        g684(.A(i_11_), .B(new_new_n208_), .Y(new_new_n707_));
  NA3        g685(.A(new_new_n692_), .B(new_new_n480_), .C(new_new_n303_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n708_), .B(new_new_n40_), .Y(new_new_n709_));
  NOi21      g687(.An(new_new_n97_), .B(new_new_n629_), .Y(new_new_n710_));
  NO3        g688(.A(new_new_n505_), .B(new_new_n370_), .C(new_new_n133_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n342_), .B(new_new_n45_), .Y(new_new_n712_));
  NO2        g690(.A(new_new_n711_), .B(new_new_n710_), .Y(new_new_n713_));
  AOI210     g691(.A0(new_new_n713_), .A1(new_new_n709_), .B0(new_new_n48_), .Y(new_new_n714_));
  NO4        g692(.A(new_new_n308_), .B(new_new_n315_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n715_));
  NA2        g693(.A(new_new_n169_), .B(new_new_n448_), .Y(new_new_n716_));
  NOi21      g694(.An(new_new_n716_), .B(new_new_n715_), .Y(new_new_n717_));
  NO2        g695(.A(new_new_n717_), .B(new_new_n61_), .Y(new_new_n718_));
  NOi21      g696(.An(i_5_), .B(i_9_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n719_), .B(new_new_n359_), .Y(new_new_n720_));
  BUFFER     g698(.A(new_new_n233_), .Y(new_new_n721_));
  AOI210     g699(.A0(new_new_n721_), .A1(new_new_n390_), .B0(new_new_n559_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n722_), .B(new_new_n720_), .Y(new_new_n723_));
  NO3        g701(.A(new_new_n723_), .B(new_new_n718_), .C(new_new_n714_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n169_), .B(new_new_n24_), .Y(new_new_n725_));
  NO2        g703(.A(new_new_n546_), .B(new_new_n471_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n726_), .B(new_new_n725_), .Y(new_new_n727_));
  NA2        g705(.A(new_new_n262_), .B(new_new_n131_), .Y(new_new_n728_));
  NAi21      g706(.An(new_new_n160_), .B(new_new_n352_), .Y(new_new_n729_));
  OAI220     g707(.A0(new_new_n729_), .A1(new_new_n700_), .B0(new_new_n728_), .B1(new_new_n334_), .Y(new_new_n730_));
  NO2        g708(.A(new_new_n730_), .B(new_new_n727_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n449_), .B(i_0_), .Y(new_new_n732_));
  NO3        g710(.A(new_new_n732_), .B(new_new_n317_), .C(new_new_n87_), .Y(new_new_n733_));
  NO4        g711(.A(new_new_n462_), .B(new_new_n191_), .C(new_new_n344_), .D(i_6_), .Y(new_new_n734_));
  AOI210     g712(.A0(new_new_n734_), .A1(i_11_), .B0(new_new_n733_), .Y(new_new_n735_));
  INV        g713(.A(new_new_n389_), .Y(new_new_n736_));
  NA2        g714(.A(new_new_n616_), .B(new_new_n269_), .Y(new_new_n737_));
  AOI210     g715(.A0(new_new_n393_), .A1(new_new_n87_), .B0(new_new_n56_), .Y(new_new_n738_));
  NO2        g716(.A(new_new_n738_), .B(new_new_n737_), .Y(new_new_n739_));
  NO2        g717(.A(new_new_n220_), .B(new_new_n154_), .Y(new_new_n740_));
  NA2        g718(.A(i_0_), .B(i_10_), .Y(new_new_n741_));
  AN2        g719(.A(new_new_n740_), .B(i_6_), .Y(new_new_n742_));
  NO2        g720(.A(new_new_n742_), .B(new_new_n739_), .Y(new_new_n743_));
  NA3        g721(.A(new_new_n743_), .B(new_new_n735_), .C(new_new_n731_), .Y(new_new_n744_));
  NO2        g722(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n745_));
  NA2        g723(.A(i_11_), .B(i_9_), .Y(new_new_n746_));
  NO3        g724(.A(i_12_), .B(new_new_n746_), .C(new_new_n479_), .Y(new_new_n747_));
  AN2        g725(.A(new_new_n747_), .B(new_new_n745_), .Y(new_new_n748_));
  NO2        g726(.A(new_new_n48_), .B(i_7_), .Y(new_new_n749_));
  NA2        g727(.A(new_new_n326_), .B(new_new_n166_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n750_), .B(new_new_n158_), .Y(new_new_n751_));
  NO2        g729(.A(new_new_n746_), .B(new_new_n71_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n165_), .B(i_0_), .Y(new_new_n753_));
  INV        g731(.A(new_new_n340_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n754_), .B(new_new_n720_), .Y(new_new_n755_));
  NO3        g733(.A(new_new_n755_), .B(new_new_n751_), .C(new_new_n748_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n533_), .B(new_new_n123_), .Y(new_new_n757_));
  NO2        g735(.A(i_6_), .B(new_new_n757_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n162_), .B(new_new_n104_), .Y(new_new_n759_));
  NA2        g737(.A(new_new_n481_), .B(new_new_n269_), .Y(new_new_n760_));
  NO2        g738(.A(new_new_n760_), .B(new_new_n712_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n761_), .B(new_new_n758_), .Y(new_new_n762_));
  NOi21      g740(.An(i_7_), .B(i_5_), .Y(new_new_n763_));
  NOi31      g741(.An(new_new_n763_), .B(i_0_), .C(new_new_n598_), .Y(new_new_n764_));
  NA3        g742(.A(new_new_n764_), .B(new_new_n316_), .C(i_6_), .Y(new_new_n765_));
  BUFFER     g743(.A(new_new_n765_), .Y(new_new_n766_));
  INV        g744(.A(new_new_n265_), .Y(new_new_n767_));
  NA3        g745(.A(new_new_n766_), .B(new_new_n762_), .C(new_new_n756_), .Y(new_new_n768_));
  NO2        g746(.A(new_new_n706_), .B(new_new_n264_), .Y(new_new_n769_));
  OA210      g747(.A0(new_new_n389_), .A1(new_new_n199_), .B0(new_new_n388_), .Y(new_new_n770_));
  NA2        g748(.A(new_new_n769_), .B(new_new_n752_), .Y(new_new_n771_));
  NA3        g749(.A(new_new_n388_), .B(new_new_n342_), .C(new_new_n45_), .Y(new_new_n772_));
  OAI210     g750(.A0(new_new_n729_), .A1(new_new_n736_), .B0(new_new_n772_), .Y(new_new_n773_));
  NA2        g751(.A(new_new_n752_), .B(new_new_n257_), .Y(new_new_n774_));
  OAI210     g752(.A0(i_3_), .A1(new_new_n171_), .B0(new_new_n774_), .Y(new_new_n775_));
  AOI220     g753(.A0(new_new_n775_), .A1(new_new_n389_), .B0(new_new_n773_), .B1(new_new_n71_), .Y(new_new_n776_));
  NA3        g754(.A(i_5_), .B(new_new_n314_), .C(new_new_n515_), .Y(new_new_n777_));
  NA2        g755(.A(new_new_n93_), .B(new_new_n44_), .Y(new_new_n778_));
  NO2        g756(.A(new_new_n73_), .B(new_new_n618_), .Y(new_new_n779_));
  AOI220     g757(.A0(new_new_n779_), .A1(new_new_n778_), .B0(new_new_n164_), .B1(new_new_n471_), .Y(new_new_n780_));
  AOI210     g758(.A0(new_new_n780_), .A1(new_new_n777_), .B0(new_new_n47_), .Y(new_new_n781_));
  NO3        g759(.A(new_new_n462_), .B(new_new_n289_), .C(new_new_n24_), .Y(new_new_n782_));
  AOI210     g760(.A0(new_new_n575_), .A1(new_new_n430_), .B0(new_new_n782_), .Y(new_new_n783_));
  NAi21      g761(.An(i_9_), .B(i_5_), .Y(new_new_n784_));
  NO2        g762(.A(new_new_n784_), .B(new_new_n335_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n785_), .B(new_new_n495_), .Y(new_new_n786_));
  OAI220     g764(.A0(new_new_n786_), .A1(new_new_n84_), .B0(new_new_n783_), .B1(new_new_n163_), .Y(new_new_n787_));
  NO2        g765(.A(new_new_n787_), .B(new_new_n781_), .Y(new_new_n788_));
  NA3        g766(.A(new_new_n788_), .B(new_new_n776_), .C(new_new_n771_), .Y(new_new_n789_));
  NO3        g767(.A(new_new_n789_), .B(new_new_n768_), .C(new_new_n744_), .Y(new_new_n790_));
  NO2        g768(.A(i_0_), .B(new_new_n598_), .Y(new_new_n791_));
  NO2        g769(.A(new_new_n664_), .B(new_new_n759_), .Y(new_new_n792_));
  INV        g770(.A(new_new_n792_), .Y(new_new_n793_));
  NO2        g771(.A(new_new_n682_), .B(new_new_n335_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n214_), .B(new_new_n206_), .Y(new_new_n795_));
  AOI210     g773(.A0(new_new_n795_), .A1(new_new_n732_), .B0(new_new_n154_), .Y(new_new_n796_));
  NO2        g774(.A(new_new_n796_), .B(new_new_n794_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n797_), .B(new_new_n793_), .Y(new_new_n798_));
  NO3        g776(.A(new_new_n741_), .B(new_new_n719_), .C(new_new_n174_), .Y(new_new_n799_));
  AOI220     g777(.A0(new_new_n799_), .A1(i_11_), .B0(new_new_n447_), .B1(new_new_n73_), .Y(new_new_n800_));
  NO3        g778(.A(new_new_n187_), .B(new_new_n315_), .C(i_0_), .Y(new_new_n801_));
  OAI210     g779(.A0(new_new_n801_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n802_), .B(new_new_n800_), .Y(new_new_n803_));
  NO2        g781(.A(new_new_n213_), .B(new_new_n93_), .Y(new_new_n804_));
  AOI210     g782(.A0(new_new_n804_), .A1(new_new_n791_), .B0(new_new_n110_), .Y(new_new_n805_));
  OR2        g783(.A(new_new_n805_), .B(i_5_), .Y(new_new_n806_));
  AOI210     g784(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n165_), .Y(new_new_n807_));
  NA2        g785(.A(new_new_n807_), .B(new_new_n770_), .Y(new_new_n808_));
  INV        g786(.A(new_new_n428_), .Y(new_new_n809_));
  NO3        g787(.A(new_new_n712_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n401_), .B(new_new_n394_), .Y(new_new_n811_));
  NO3        g789(.A(new_new_n811_), .B(new_new_n810_), .C(new_new_n809_), .Y(new_new_n812_));
  NA3        g790(.A(new_new_n321_), .B(new_new_n162_), .C(new_new_n161_), .Y(new_new_n813_));
  NA3        g791(.A(new_new_n749_), .B(new_new_n249_), .C(new_new_n206_), .Y(new_new_n814_));
  NA2        g792(.A(new_new_n814_), .B(new_new_n813_), .Y(new_new_n815_));
  NA3        g793(.A(new_new_n321_), .B(new_new_n276_), .C(new_new_n197_), .Y(new_new_n816_));
  INV        g794(.A(new_new_n816_), .Y(new_new_n817_));
  NO3        g795(.A(new_new_n746_), .B(new_new_n194_), .C(new_new_n174_), .Y(new_new_n818_));
  NO3        g796(.A(new_new_n818_), .B(new_new_n817_), .C(new_new_n815_), .Y(new_new_n819_));
  NA4        g797(.A(new_new_n819_), .B(new_new_n812_), .C(new_new_n808_), .D(new_new_n806_), .Y(new_new_n820_));
  NO2        g798(.A(new_new_n84_), .B(i_5_), .Y(new_new_n821_));
  NA3        g799(.A(new_new_n707_), .B(new_new_n111_), .C(new_new_n126_), .Y(new_new_n822_));
  INV        g800(.A(new_new_n822_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n823_), .B(new_new_n821_), .Y(new_new_n824_));
  NA3        g802(.A(new_new_n257_), .B(i_5_), .C(new_new_n175_), .Y(new_new_n825_));
  NAi31      g803(.An(new_new_n212_), .B(new_new_n825_), .C(new_new_n213_), .Y(new_new_n826_));
  NO4        g804(.A(new_new_n211_), .B(new_new_n187_), .C(i_0_), .D(i_12_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n827_), .B(new_new_n826_), .Y(new_new_n828_));
  AN2        g806(.A(new_new_n741_), .B(new_new_n154_), .Y(new_new_n829_));
  NO4        g807(.A(new_new_n829_), .B(i_12_), .C(new_new_n521_), .D(new_new_n133_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n830_), .B(new_new_n194_), .Y(new_new_n831_));
  NA2        g809(.A(new_new_n763_), .B(new_new_n386_), .Y(new_new_n832_));
  NA2        g810(.A(new_new_n62_), .B(new_new_n102_), .Y(new_new_n833_));
  OAI220     g811(.A0(new_new_n833_), .A1(new_new_n825_), .B0(new_new_n832_), .B1(new_new_n549_), .Y(new_new_n834_));
  NA2        g812(.A(new_new_n834_), .B(new_new_n753_), .Y(new_new_n835_));
  NA4        g813(.A(new_new_n835_), .B(new_new_n831_), .C(new_new_n828_), .D(new_new_n824_), .Y(new_new_n836_));
  NO4        g814(.A(new_new_n836_), .B(new_new_n820_), .C(new_new_n803_), .D(new_new_n798_), .Y(new_new_n837_));
  OAI210     g815(.A0(new_new_n685_), .A1(new_new_n678_), .B0(new_new_n37_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n838_), .B(new_new_n487_), .Y(new_new_n839_));
  NA2        g817(.A(new_new_n839_), .B(new_new_n185_), .Y(new_new_n840_));
  NAi31      g818(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n841_));
  AOI210     g819(.A0(new_new_n119_), .A1(new_new_n68_), .B0(new_new_n841_), .Y(new_new_n842_));
  NO2        g820(.A(new_new_n842_), .B(new_new_n518_), .Y(new_new_n843_));
  INV        g821(.A(new_new_n843_), .Y(new_new_n844_));
  AOI210     g822(.A0(new_new_n844_), .A1(new_new_n48_), .B0(new_new_n734_), .Y(new_new_n845_));
  AOI210     g823(.A0(new_new_n845_), .A1(new_new_n840_), .B0(new_new_n71_), .Y(new_new_n846_));
  INV        g824(.A(new_new_n311_), .Y(new_new_n847_));
  NO2        g825(.A(new_new_n847_), .B(new_new_n624_), .Y(new_new_n848_));
  OAI210     g826(.A0(new_new_n78_), .A1(new_new_n54_), .B0(new_new_n109_), .Y(new_new_n849_));
  NA2        g827(.A(new_new_n849_), .B(new_new_n74_), .Y(new_new_n850_));
  AOI210     g828(.A0(new_new_n807_), .A1(new_new_n749_), .B0(new_new_n764_), .Y(new_new_n851_));
  AOI210     g829(.A0(new_new_n851_), .A1(new_new_n850_), .B0(new_new_n552_), .Y(new_new_n852_));
  INV        g830(.A(new_new_n852_), .Y(new_new_n853_));
  OAI210     g831(.A0(new_new_n235_), .A1(new_new_n156_), .B0(new_new_n87_), .Y(new_new_n854_));
  NA3        g832(.A(new_new_n628_), .B(new_new_n249_), .C(new_new_n78_), .Y(new_new_n855_));
  AOI210     g833(.A0(new_new_n855_), .A1(new_new_n854_), .B0(i_11_), .Y(new_new_n856_));
  NO3        g834(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n857_));
  OAI210     g835(.A0(new_new_n767_), .A1(new_new_n258_), .B0(new_new_n857_), .Y(new_new_n858_));
  NO2        g836(.A(new_new_n858_), .B(new_new_n598_), .Y(new_new_n859_));
  NO4        g837(.A(new_new_n784_), .B(new_new_n391_), .C(new_new_n219_), .D(new_new_n218_), .Y(new_new_n860_));
  NO2        g838(.A(new_new_n860_), .B(new_new_n443_), .Y(new_new_n861_));
  INV        g839(.A(new_new_n292_), .Y(new_new_n862_));
  AOI210     g840(.A0(new_new_n862_), .A1(new_new_n861_), .B0(new_new_n41_), .Y(new_new_n863_));
  NO3        g841(.A(new_new_n863_), .B(new_new_n859_), .C(new_new_n856_), .Y(new_new_n864_));
  OAI210     g842(.A0(new_new_n853_), .A1(i_4_), .B0(new_new_n864_), .Y(new_new_n865_));
  NO3        g843(.A(new_new_n865_), .B(new_new_n848_), .C(new_new_n846_), .Y(new_new_n866_));
  NA4        g844(.A(new_new_n866_), .B(new_new_n837_), .C(new_new_n790_), .D(new_new_n724_), .Y(ori4));
  INV        g845(.A(new_new_n574_), .Y(new_new_n870_));
  INV        g846(.A(new_new_n273_), .Y(new_new_n871_));
  INV        g847(.A(new_new_n586_), .Y(new_new_n872_));
endmodule


