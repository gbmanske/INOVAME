//Benchmark atmr_9sym_175_0.0313

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n167_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n166_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n171_, men_men_n172_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  NA2        o002(.A(i_4_), .B(ori_ori_n12_), .Y(ori_ori_n13_));
  INV        o003(.A(i_5_), .Y(ori_ori_n14_));
  NOi21      o004(.An(i_3_), .B(i_7_), .Y(ori_ori_n15_));
  NA3        o005(.A(ori_ori_n15_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n16_));
  INV        o006(.A(i_0_), .Y(ori_ori_n17_));
  NOi21      o007(.An(i_1_), .B(i_3_), .Y(ori_ori_n18_));
  NO2        o008(.A(ori_ori_n16_), .B(ori_ori_n13_), .Y(ori_ori_n19_));
  INV        o009(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o010(.A(i_0_), .B(ori_ori_n20_), .Y(ori_ori_n21_));
  INV        o011(.A(i_7_), .Y(ori_ori_n22_));
  NA3        o012(.A(i_6_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n23_));
  NOi21      o013(.An(i_8_), .B(i_6_), .Y(ori_ori_n24_));
  NOi21      o014(.An(i_1_), .B(i_8_), .Y(ori_ori_n25_));
  AOI220     o015(.A0(ori_ori_n25_), .A1(i_2_), .B0(ori_ori_n24_), .B1(i_5_), .Y(ori_ori_n26_));
  AOI210     o016(.A0(ori_ori_n26_), .A1(ori_ori_n23_), .B0(ori_ori_n21_), .Y(ori_ori_n27_));
  AOI210     o017(.A0(ori_ori_n27_), .A1(ori_ori_n11_), .B0(ori_ori_n19_), .Y(ori_ori_n28_));
  NA2        o018(.A(i_0_), .B(ori_ori_n14_), .Y(ori_ori_n29_));
  NA2        o019(.A(ori_ori_n17_), .B(i_5_), .Y(ori_ori_n30_));
  NO2        o020(.A(i_2_), .B(i_4_), .Y(ori_ori_n31_));
  NA3        o021(.A(ori_ori_n31_), .B(i_6_), .C(i_8_), .Y(ori_ori_n32_));
  AOI210     o022(.A0(ori_ori_n30_), .A1(ori_ori_n29_), .B0(ori_ori_n32_), .Y(ori_ori_n33_));
  INV        o023(.A(i_2_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_5_), .B(i_0_), .Y(ori_ori_n35_));
  NOi21      o025(.An(i_6_), .B(i_8_), .Y(ori_ori_n36_));
  NOi21      o026(.An(i_7_), .B(i_1_), .Y(ori_ori_n37_));
  NOi21      o027(.An(i_5_), .B(i_6_), .Y(ori_ori_n38_));
  AOI220     o028(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n36_), .B1(ori_ori_n35_), .Y(ori_ori_n39_));
  NO3        o029(.A(ori_ori_n39_), .B(ori_ori_n34_), .C(i_4_), .Y(ori_ori_n40_));
  NOi21      o030(.An(i_0_), .B(i_4_), .Y(ori_ori_n41_));
  XO2        o031(.A(i_1_), .B(i_3_), .Y(ori_ori_n42_));
  NOi21      o032(.An(i_7_), .B(i_5_), .Y(ori_ori_n43_));
  AN3        o033(.A(ori_ori_n43_), .B(ori_ori_n42_), .C(ori_ori_n41_), .Y(ori_ori_n44_));
  INV        o034(.A(i_1_), .Y(ori_ori_n45_));
  NOi21      o035(.An(i_3_), .B(i_0_), .Y(ori_ori_n46_));
  NA2        o036(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o037(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n48_));
  NO4        o038(.A(ori_ori_n48_), .B(ori_ori_n44_), .C(ori_ori_n40_), .D(ori_ori_n33_), .Y(ori_ori_n49_));
  NOi21      o039(.An(i_4_), .B(i_0_), .Y(ori_ori_n50_));
  NO2        o040(.A(ori_ori_n24_), .B(ori_ori_n15_), .Y(ori_ori_n51_));
  NA2        o041(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n52_));
  NOi21      o042(.An(i_2_), .B(i_8_), .Y(ori_ori_n53_));
  NO2        o043(.A(ori_ori_n53_), .B(ori_ori_n41_), .Y(ori_ori_n54_));
  NO3        o044(.A(ori_ori_n54_), .B(ori_ori_n52_), .C(ori_ori_n51_), .Y(ori_ori_n55_));
  INV        o045(.A(ori_ori_n55_), .Y(ori_ori_n56_));
  NOi31      o046(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n57_));
  NA2        o047(.A(ori_ori_n57_), .B(i_0_), .Y(ori_ori_n58_));
  NOi21      o048(.An(i_4_), .B(i_3_), .Y(ori_ori_n59_));
  NOi21      o049(.An(i_1_), .B(i_4_), .Y(ori_ori_n60_));
  OAI210     o050(.A0(ori_ori_n60_), .A1(ori_ori_n59_), .B0(ori_ori_n53_), .Y(ori_ori_n61_));
  NA2        o051(.A(ori_ori_n61_), .B(ori_ori_n58_), .Y(ori_ori_n62_));
  AN2        o052(.A(i_8_), .B(i_7_), .Y(ori_ori_n63_));
  INV        o053(.A(ori_ori_n63_), .Y(ori_ori_n64_));
  NOi21      o054(.An(i_8_), .B(i_7_), .Y(ori_ori_n65_));
  NA3        o055(.A(ori_ori_n65_), .B(ori_ori_n59_), .C(i_6_), .Y(ori_ori_n66_));
  OAI210     o056(.A0(ori_ori_n64_), .A1(ori_ori_n52_), .B0(ori_ori_n66_), .Y(ori_ori_n67_));
  AOI220     o057(.A0(ori_ori_n67_), .A1(ori_ori_n34_), .B0(ori_ori_n62_), .B1(ori_ori_n38_), .Y(ori_ori_n68_));
  NA4        o058(.A(ori_ori_n68_), .B(ori_ori_n56_), .C(ori_ori_n49_), .D(ori_ori_n28_), .Y(ori_ori_n69_));
  INV        o059(.A(i_8_), .Y(ori_ori_n70_));
  NO3        o060(.A(ori_ori_n70_), .B(ori_ori_n13_), .C(i_1_), .Y(ori_ori_n71_));
  NA2        o061(.A(i_8_), .B(ori_ori_n22_), .Y(ori_ori_n72_));
  AOI220     o062(.A0(ori_ori_n46_), .A1(i_1_), .B0(ori_ori_n42_), .B1(i_2_), .Y(ori_ori_n73_));
  NOi21      o063(.An(i_1_), .B(i_2_), .Y(ori_ori_n74_));
  NO2        o064(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n75_));
  OAI210     o065(.A0(ori_ori_n75_), .A1(ori_ori_n71_), .B0(ori_ori_n14_), .Y(ori_ori_n76_));
  NA2        o066(.A(ori_ori_n65_), .B(ori_ori_n12_), .Y(ori_ori_n77_));
  NA2        o067(.A(ori_ori_n25_), .B(ori_ori_n14_), .Y(ori_ori_n78_));
  NA2        o068(.A(ori_ori_n78_), .B(ori_ori_n77_), .Y(ori_ori_n79_));
  NOi32      o069(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(ori_ori_n80_));
  NA2        o070(.A(ori_ori_n18_), .B(i_6_), .Y(ori_ori_n81_));
  INV        o071(.A(ori_ori_n81_), .Y(ori_ori_n82_));
  INV        o072(.A(i_0_), .Y(ori_ori_n83_));
  AOI220     o073(.A0(ori_ori_n83_), .A1(ori_ori_n82_), .B0(ori_ori_n79_), .B1(ori_ori_n59_), .Y(ori_ori_n84_));
  NA2        o074(.A(ori_ori_n84_), .B(ori_ori_n76_), .Y(ori_ori_n85_));
  NAi21      o075(.An(i_3_), .B(i_6_), .Y(ori_ori_n86_));
  NA2        o076(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n87_));
  NOi21      o077(.An(i_7_), .B(i_8_), .Y(ori_ori_n88_));
  NOi21      o078(.An(i_6_), .B(i_5_), .Y(ori_ori_n89_));
  AOI210     o079(.A0(ori_ori_n88_), .A1(ori_ori_n12_), .B0(ori_ori_n89_), .Y(ori_ori_n90_));
  OAI210     o080(.A0(ori_ori_n90_), .A1(ori_ori_n11_), .B0(ori_ori_n87_), .Y(ori_ori_n91_));
  NA2        o081(.A(ori_ori_n91_), .B(ori_ori_n74_), .Y(ori_ori_n92_));
  AOI220     o082(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n18_), .B1(ori_ori_n34_), .Y(ori_ori_n93_));
  NA3        o083(.A(ori_ori_n20_), .B(i_5_), .C(i_7_), .Y(ori_ori_n94_));
  NO2        o084(.A(ori_ori_n94_), .B(ori_ori_n93_), .Y(ori_ori_n95_));
  INV        o085(.A(ori_ori_n95_), .Y(ori_ori_n96_));
  NA3        o086(.A(ori_ori_n65_), .B(ori_ori_n34_), .C(i_3_), .Y(ori_ori_n97_));
  NA2        o087(.A(ori_ori_n45_), .B(i_6_), .Y(ori_ori_n98_));
  AOI210     o088(.A0(ori_ori_n98_), .A1(ori_ori_n21_), .B0(ori_ori_n97_), .Y(ori_ori_n99_));
  NOi21      o089(.An(i_2_), .B(i_1_), .Y(ori_ori_n100_));
  AN3        o090(.A(ori_ori_n88_), .B(ori_ori_n100_), .C(ori_ori_n50_), .Y(ori_ori_n101_));
  NAi21      o091(.An(i_6_), .B(i_0_), .Y(ori_ori_n102_));
  NA3        o092(.A(ori_ori_n60_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n103_));
  NOi21      o093(.An(i_4_), .B(i_6_), .Y(ori_ori_n104_));
  INV        o094(.A(i_3_), .Y(ori_ori_n105_));
  NA2        o095(.A(ori_ori_n74_), .B(ori_ori_n104_), .Y(ori_ori_n106_));
  OAI210     o096(.A0(ori_ori_n103_), .A1(ori_ori_n102_), .B0(ori_ori_n106_), .Y(ori_ori_n107_));
  NA2        o097(.A(ori_ori_n74_), .B(ori_ori_n36_), .Y(ori_ori_n108_));
  NO3        o098(.A(ori_ori_n107_), .B(ori_ori_n101_), .C(ori_ori_n99_), .Y(ori_ori_n109_));
  NOi31      o099(.An(ori_ori_n50_), .B(ori_ori_n167_), .C(i_2_), .Y(ori_ori_n110_));
  NA2        o100(.A(ori_ori_n65_), .B(ori_ori_n12_), .Y(ori_ori_n111_));
  NA2        o101(.A(ori_ori_n36_), .B(ori_ori_n14_), .Y(ori_ori_n112_));
  NOi21      o102(.An(i_3_), .B(i_1_), .Y(ori_ori_n113_));
  NA2        o103(.A(ori_ori_n113_), .B(i_4_), .Y(ori_ori_n114_));
  AOI210     o104(.A0(ori_ori_n112_), .A1(ori_ori_n111_), .B0(ori_ori_n114_), .Y(ori_ori_n115_));
  NOi31      o105(.An(ori_ori_n46_), .B(i_5_), .C(ori_ori_n34_), .Y(ori_ori_n116_));
  NO3        o106(.A(ori_ori_n116_), .B(ori_ori_n115_), .C(ori_ori_n110_), .Y(ori_ori_n117_));
  NA4        o107(.A(ori_ori_n117_), .B(ori_ori_n109_), .C(ori_ori_n96_), .D(ori_ori_n92_), .Y(ori_ori_n118_));
  NA2        o108(.A(ori_ori_n53_), .B(ori_ori_n15_), .Y(ori_ori_n119_));
  NOi31      o109(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n120_));
  NOi31      o110(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n121_));
  OAI210     o111(.A0(ori_ori_n121_), .A1(ori_ori_n120_), .B0(i_7_), .Y(ori_ori_n122_));
  NA2        o112(.A(ori_ori_n36_), .B(ori_ori_n14_), .Y(ori_ori_n123_));
  NA4        o113(.A(ori_ori_n123_), .B(ori_ori_n122_), .C(ori_ori_n119_), .D(ori_ori_n108_), .Y(ori_ori_n124_));
  NA2        o114(.A(ori_ori_n124_), .B(ori_ori_n41_), .Y(ori_ori_n125_));
  NA2        o115(.A(ori_ori_n59_), .B(ori_ori_n37_), .Y(ori_ori_n126_));
  AOI210     o116(.A0(ori_ori_n126_), .A1(ori_ori_n77_), .B0(ori_ori_n30_), .Y(ori_ori_n127_));
  NA3        o117(.A(ori_ori_n63_), .B(ori_ori_n17_), .C(ori_ori_n12_), .Y(ori_ori_n128_));
  NAi31      o118(.An(ori_ori_n102_), .B(ori_ori_n88_), .C(ori_ori_n100_), .Y(ori_ori_n129_));
  NA3        o119(.A(ori_ori_n65_), .B(ori_ori_n57_), .C(i_6_), .Y(ori_ori_n130_));
  NA3        o120(.A(ori_ori_n130_), .B(ori_ori_n129_), .C(ori_ori_n128_), .Y(ori_ori_n131_));
  NOi21      o121(.An(i_0_), .B(i_2_), .Y(ori_ori_n132_));
  NA3        o122(.A(ori_ori_n132_), .B(ori_ori_n37_), .C(ori_ori_n104_), .Y(ori_ori_n133_));
  NOi32      o123(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n134_));
  NA2        o124(.A(ori_ori_n134_), .B(ori_ori_n120_), .Y(ori_ori_n135_));
  NA3        o125(.A(ori_ori_n132_), .B(ori_ori_n59_), .C(ori_ori_n36_), .Y(ori_ori_n136_));
  NA3        o126(.A(ori_ori_n136_), .B(ori_ori_n135_), .C(ori_ori_n133_), .Y(ori_ori_n137_));
  NA4        o127(.A(ori_ori_n57_), .B(i_6_), .C(ori_ori_n14_), .D(i_7_), .Y(ori_ori_n138_));
  NA4        o128(.A(ori_ori_n60_), .B(ori_ori_n46_), .C(i_5_), .D(ori_ori_n22_), .Y(ori_ori_n139_));
  NA2        o129(.A(ori_ori_n139_), .B(ori_ori_n138_), .Y(ori_ori_n140_));
  NO4        o130(.A(ori_ori_n140_), .B(ori_ori_n137_), .C(ori_ori_n131_), .D(ori_ori_n127_), .Y(ori_ori_n141_));
  INV        o131(.A(i_2_), .Y(ori_ori_n142_));
  AOI220     o132(.A0(ori_ori_n142_), .A1(ori_ori_n88_), .B0(ori_ori_n63_), .B1(ori_ori_n31_), .Y(ori_ori_n143_));
  AOI210     o133(.A0(ori_ori_n143_), .A1(ori_ori_n119_), .B0(ori_ori_n98_), .Y(ori_ori_n144_));
  NO4        o134(.A(i_2_), .B(ori_ori_n20_), .C(ori_ori_n11_), .D(ori_ori_n14_), .Y(ori_ori_n145_));
  NA2        o135(.A(i_2_), .B(i_4_), .Y(ori_ori_n146_));
  AOI210     o136(.A0(ori_ori_n102_), .A1(ori_ori_n86_), .B0(ori_ori_n146_), .Y(ori_ori_n147_));
  NO2        o137(.A(i_8_), .B(i_7_), .Y(ori_ori_n148_));
  OA210      o138(.A0(ori_ori_n147_), .A1(ori_ori_n145_), .B0(ori_ori_n148_), .Y(ori_ori_n149_));
  NA4        o139(.A(ori_ori_n113_), .B(i_0_), .C(i_5_), .D(ori_ori_n22_), .Y(ori_ori_n150_));
  NO2        o140(.A(ori_ori_n150_), .B(i_4_), .Y(ori_ori_n151_));
  NO3        o141(.A(ori_ori_n151_), .B(ori_ori_n149_), .C(ori_ori_n144_), .Y(ori_ori_n152_));
  NA2        o142(.A(ori_ori_n88_), .B(ori_ori_n12_), .Y(ori_ori_n153_));
  NA3        o143(.A(i_2_), .B(i_1_), .C(ori_ori_n14_), .Y(ori_ori_n154_));
  NA2        o144(.A(ori_ori_n50_), .B(i_3_), .Y(ori_ori_n155_));
  AOI210     o145(.A0(ori_ori_n155_), .A1(ori_ori_n154_), .B0(ori_ori_n153_), .Y(ori_ori_n156_));
  NA4        o146(.A(ori_ori_n105_), .B(ori_ori_n63_), .C(ori_ori_n45_), .D(ori_ori_n20_), .Y(ori_ori_n157_));
  NA3        o147(.A(ori_ori_n53_), .B(ori_ori_n35_), .C(ori_ori_n15_), .Y(ori_ori_n158_));
  NOi31      o148(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n159_));
  OAI210     o149(.A0(ori_ori_n134_), .A1(ori_ori_n80_), .B0(ori_ori_n159_), .Y(ori_ori_n160_));
  NA3        o150(.A(ori_ori_n160_), .B(ori_ori_n158_), .C(ori_ori_n157_), .Y(ori_ori_n161_));
  NO2        o151(.A(ori_ori_n161_), .B(ori_ori_n156_), .Y(ori_ori_n162_));
  NA4        o152(.A(ori_ori_n162_), .B(ori_ori_n152_), .C(ori_ori_n141_), .D(ori_ori_n125_), .Y(ori_ori_n163_));
  OR4        o153(.A(ori_ori_n163_), .B(ori_ori_n118_), .C(ori_ori_n85_), .D(ori_ori_n69_), .Y(ori00));
  INV        o154(.A(i_8_), .Y(ori_ori_n167_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  INV        m002(.A(i_5_), .Y(mai_mai_n13_));
  NOi21      m003(.An(i_3_), .B(i_7_), .Y(mai_mai_n14_));
  INV        m004(.A(i_0_), .Y(mai_mai_n15_));
  NOi21      m005(.An(i_1_), .B(i_3_), .Y(mai_mai_n16_));
  INV        m006(.A(i_4_), .Y(mai_mai_n17_));
  NA2        m007(.A(i_0_), .B(mai_mai_n17_), .Y(mai_mai_n18_));
  INV        m008(.A(i_7_), .Y(mai_mai_n19_));
  NA3        m009(.A(i_6_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n20_));
  NOi21      m010(.An(i_8_), .B(i_6_), .Y(mai_mai_n21_));
  NOi21      m011(.An(i_1_), .B(i_8_), .Y(mai_mai_n22_));
  AOI220     m012(.A0(mai_mai_n22_), .A1(i_2_), .B0(mai_mai_n21_), .B1(i_5_), .Y(mai_mai_n23_));
  AOI210     m013(.A0(mai_mai_n23_), .A1(mai_mai_n20_), .B0(mai_mai_n18_), .Y(mai_mai_n24_));
  NA2        m014(.A(mai_mai_n24_), .B(mai_mai_n11_), .Y(mai_mai_n25_));
  NA2        m015(.A(i_0_), .B(mai_mai_n13_), .Y(mai_mai_n26_));
  NA2        m016(.A(mai_mai_n15_), .B(i_5_), .Y(mai_mai_n27_));
  NO2        m017(.A(i_2_), .B(i_4_), .Y(mai_mai_n28_));
  NA3        m018(.A(mai_mai_n28_), .B(i_6_), .C(i_8_), .Y(mai_mai_n29_));
  AOI210     m019(.A0(mai_mai_n27_), .A1(mai_mai_n26_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  INV        m020(.A(i_2_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_5_), .B(i_0_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_6_), .B(i_8_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_7_), .B(i_1_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_5_), .B(i_6_), .Y(mai_mai_n35_));
  AOI220     m025(.A0(mai_mai_n35_), .A1(mai_mai_n34_), .B0(mai_mai_n33_), .B1(mai_mai_n32_), .Y(mai_mai_n36_));
  NO3        m026(.A(mai_mai_n36_), .B(mai_mai_n31_), .C(i_4_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_0_), .B(i_4_), .Y(mai_mai_n38_));
  NOi21      m028(.An(i_7_), .B(i_5_), .Y(mai_mai_n39_));
  AN2        m029(.A(mai_mai_n39_), .B(mai_mai_n38_), .Y(mai_mai_n40_));
  INV        m030(.A(i_1_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_3_), .B(i_0_), .Y(mai_mai_n42_));
  NA2        m032(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA3        m033(.A(i_6_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n44_));
  AOI210     m034(.A0(mai_mai_n44_), .A1(mai_mai_n20_), .B0(mai_mai_n43_), .Y(mai_mai_n45_));
  NO4        m035(.A(mai_mai_n45_), .B(mai_mai_n40_), .C(mai_mai_n37_), .D(mai_mai_n30_), .Y(mai_mai_n46_));
  INV        m036(.A(i_8_), .Y(mai_mai_n47_));
  NA2        m037(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n48_));
  NO4        m038(.A(mai_mai_n48_), .B(mai_mai_n26_), .C(i_2_), .D(mai_mai_n47_), .Y(mai_mai_n49_));
  NOi21      m039(.An(i_4_), .B(i_0_), .Y(mai_mai_n50_));
  AOI210     m040(.A0(mai_mai_n50_), .A1(mai_mai_n21_), .B0(mai_mai_n14_), .Y(mai_mai_n51_));
  NA2        m041(.A(i_1_), .B(mai_mai_n13_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_2_), .B(i_8_), .Y(mai_mai_n53_));
  NO2        m043(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n54_));
  NO2        m044(.A(mai_mai_n54_), .B(mai_mai_n49_), .Y(mai_mai_n55_));
  NOi31      m045(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n56_));
  NA2        m046(.A(mai_mai_n56_), .B(i_0_), .Y(mai_mai_n57_));
  NOi21      m047(.An(i_4_), .B(i_3_), .Y(mai_mai_n58_));
  NOi21      m048(.An(i_1_), .B(i_4_), .Y(mai_mai_n59_));
  OAI210     m049(.A0(mai_mai_n59_), .A1(mai_mai_n58_), .B0(mai_mai_n53_), .Y(mai_mai_n60_));
  NA2        m050(.A(mai_mai_n60_), .B(mai_mai_n57_), .Y(mai_mai_n61_));
  AN2        m051(.A(i_8_), .B(i_7_), .Y(mai_mai_n62_));
  NA2        m052(.A(mai_mai_n62_), .B(mai_mai_n12_), .Y(mai_mai_n63_));
  NOi21      m053(.An(i_8_), .B(i_7_), .Y(mai_mai_n64_));
  NA3        m054(.A(mai_mai_n64_), .B(mai_mai_n58_), .C(i_6_), .Y(mai_mai_n65_));
  OAI210     m055(.A0(mai_mai_n63_), .A1(mai_mai_n52_), .B0(mai_mai_n65_), .Y(mai_mai_n66_));
  AOI220     m056(.A0(mai_mai_n66_), .A1(mai_mai_n31_), .B0(mai_mai_n61_), .B1(mai_mai_n35_), .Y(mai_mai_n67_));
  NA4        m057(.A(mai_mai_n67_), .B(mai_mai_n55_), .C(mai_mai_n46_), .D(mai_mai_n25_), .Y(mai_mai_n68_));
  NA2        m058(.A(i_8_), .B(mai_mai_n19_), .Y(mai_mai_n69_));
  NOi21      m059(.An(i_1_), .B(i_2_), .Y(mai_mai_n70_));
  NA3        m060(.A(mai_mai_n70_), .B(mai_mai_n50_), .C(i_6_), .Y(mai_mai_n71_));
  OAI210     m061(.A0(mai_mai_n166_), .A1(mai_mai_n69_), .B0(mai_mai_n71_), .Y(mai_mai_n72_));
  NA2        m062(.A(mai_mai_n72_), .B(mai_mai_n13_), .Y(mai_mai_n73_));
  NA3        m063(.A(mai_mai_n64_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n74_));
  NA3        m064(.A(mai_mai_n22_), .B(i_0_), .C(mai_mai_n13_), .Y(mai_mai_n75_));
  NA2        m065(.A(mai_mai_n75_), .B(mai_mai_n74_), .Y(mai_mai_n76_));
  NOi32      m066(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n77_));
  NA2        m067(.A(mai_mai_n77_), .B(i_3_), .Y(mai_mai_n78_));
  NA3        m068(.A(mai_mai_n16_), .B(i_2_), .C(i_6_), .Y(mai_mai_n79_));
  NA2        m069(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  NO2        m070(.A(i_0_), .B(i_4_), .Y(mai_mai_n81_));
  AOI220     m071(.A0(mai_mai_n81_), .A1(mai_mai_n80_), .B0(mai_mai_n76_), .B1(mai_mai_n58_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n82_), .B(mai_mai_n73_), .Y(mai_mai_n83_));
  NAi21      m073(.An(i_3_), .B(i_6_), .Y(mai_mai_n84_));
  NO3        m074(.A(mai_mai_n84_), .B(i_0_), .C(mai_mai_n47_), .Y(mai_mai_n85_));
  NA2        m075(.A(mai_mai_n33_), .B(mai_mai_n32_), .Y(mai_mai_n86_));
  NOi21      m076(.An(i_7_), .B(i_8_), .Y(mai_mai_n87_));
  NA2        m077(.A(mai_mai_n87_), .B(mai_mai_n12_), .Y(mai_mai_n88_));
  OAI210     m078(.A0(mai_mai_n88_), .A1(mai_mai_n11_), .B0(mai_mai_n86_), .Y(mai_mai_n89_));
  OAI210     m079(.A0(mai_mai_n89_), .A1(mai_mai_n85_), .B0(mai_mai_n70_), .Y(mai_mai_n90_));
  NA3        m080(.A(mai_mai_n21_), .B(i_2_), .C(mai_mai_n13_), .Y(mai_mai_n91_));
  NO2        m081(.A(mai_mai_n48_), .B(mai_mai_n91_), .Y(mai_mai_n92_));
  AOI220     m082(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n16_), .B1(mai_mai_n31_), .Y(mai_mai_n93_));
  NA3        m083(.A(mai_mai_n17_), .B(i_5_), .C(i_7_), .Y(mai_mai_n94_));
  NO2        m084(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n95_));
  NO2        m085(.A(mai_mai_n95_), .B(mai_mai_n92_), .Y(mai_mai_n96_));
  NA3        m086(.A(mai_mai_n64_), .B(mai_mai_n31_), .C(i_3_), .Y(mai_mai_n97_));
  NA2        m087(.A(mai_mai_n41_), .B(i_6_), .Y(mai_mai_n98_));
  AOI210     m088(.A0(mai_mai_n98_), .A1(mai_mai_n18_), .B0(mai_mai_n97_), .Y(mai_mai_n99_));
  NAi21      m089(.An(i_6_), .B(i_0_), .Y(mai_mai_n100_));
  NA3        m090(.A(mai_mai_n59_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n101_));
  NOi21      m091(.An(i_4_), .B(i_6_), .Y(mai_mai_n102_));
  NOi21      m092(.An(i_5_), .B(i_3_), .Y(mai_mai_n103_));
  NA3        m093(.A(mai_mai_n103_), .B(mai_mai_n70_), .C(mai_mai_n102_), .Y(mai_mai_n104_));
  OAI210     m094(.A0(mai_mai_n101_), .A1(mai_mai_n100_), .B0(mai_mai_n104_), .Y(mai_mai_n105_));
  NA2        m095(.A(mai_mai_n70_), .B(mai_mai_n33_), .Y(mai_mai_n106_));
  NOi21      m096(.An(mai_mai_n39_), .B(mai_mai_n106_), .Y(mai_mai_n107_));
  NO3        m097(.A(mai_mai_n107_), .B(mai_mai_n105_), .C(mai_mai_n99_), .Y(mai_mai_n108_));
  NOi21      m098(.An(i_6_), .B(i_1_), .Y(mai_mai_n109_));
  AOI220     m099(.A0(mai_mai_n109_), .A1(i_7_), .B0(mai_mai_n21_), .B1(i_5_), .Y(mai_mai_n110_));
  NOi31      m100(.An(mai_mai_n50_), .B(mai_mai_n110_), .C(i_2_), .Y(mai_mai_n111_));
  NOi21      m101(.An(i_3_), .B(i_1_), .Y(mai_mai_n112_));
  NA2        m102(.A(mai_mai_n112_), .B(i_4_), .Y(mai_mai_n113_));
  AOI210     m103(.A0(i_8_), .A1(i_6_), .B0(mai_mai_n113_), .Y(mai_mai_n114_));
  NA2        m104(.A(mai_mai_n87_), .B(mai_mai_n13_), .Y(mai_mai_n115_));
  NOi31      m105(.An(mai_mai_n42_), .B(mai_mai_n115_), .C(mai_mai_n31_), .Y(mai_mai_n116_));
  NO3        m106(.A(mai_mai_n116_), .B(mai_mai_n114_), .C(mai_mai_n111_), .Y(mai_mai_n117_));
  NA4        m107(.A(mai_mai_n117_), .B(mai_mai_n108_), .C(mai_mai_n96_), .D(mai_mai_n90_), .Y(mai_mai_n118_));
  NA2        m108(.A(mai_mai_n53_), .B(mai_mai_n14_), .Y(mai_mai_n119_));
  NOi31      m109(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n120_));
  NA2        m110(.A(mai_mai_n120_), .B(i_7_), .Y(mai_mai_n121_));
  NA3        m111(.A(mai_mai_n33_), .B(i_2_), .C(mai_mai_n13_), .Y(mai_mai_n122_));
  NA4        m112(.A(mai_mai_n122_), .B(mai_mai_n121_), .C(mai_mai_n119_), .D(mai_mai_n106_), .Y(mai_mai_n123_));
  NA2        m113(.A(mai_mai_n123_), .B(mai_mai_n38_), .Y(mai_mai_n124_));
  NA2        m114(.A(mai_mai_n58_), .B(mai_mai_n34_), .Y(mai_mai_n125_));
  AOI210     m115(.A0(mai_mai_n125_), .A1(mai_mai_n74_), .B0(mai_mai_n27_), .Y(mai_mai_n126_));
  NA3        m116(.A(mai_mai_n64_), .B(mai_mai_n56_), .C(i_6_), .Y(mai_mai_n127_));
  INV        m117(.A(mai_mai_n127_), .Y(mai_mai_n128_));
  NOi21      m118(.An(i_0_), .B(i_2_), .Y(mai_mai_n129_));
  NA3        m119(.A(mai_mai_n129_), .B(mai_mai_n34_), .C(mai_mai_n102_), .Y(mai_mai_n130_));
  NA3        m120(.A(mai_mai_n50_), .B(mai_mai_n39_), .C(mai_mai_n16_), .Y(mai_mai_n131_));
  NOi32      m121(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(mai_mai_n132_));
  NA3        m122(.A(mai_mai_n129_), .B(mai_mai_n58_), .C(mai_mai_n33_), .Y(mai_mai_n133_));
  NA3        m123(.A(mai_mai_n133_), .B(mai_mai_n131_), .C(mai_mai_n130_), .Y(mai_mai_n134_));
  NA3        m124(.A(mai_mai_n56_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n135_));
  NA4        m125(.A(mai_mai_n59_), .B(mai_mai_n35_), .C(mai_mai_n15_), .D(i_8_), .Y(mai_mai_n136_));
  NA4        m126(.A(mai_mai_n59_), .B(mai_mai_n42_), .C(i_5_), .D(mai_mai_n19_), .Y(mai_mai_n137_));
  NA3        m127(.A(mai_mai_n137_), .B(mai_mai_n136_), .C(mai_mai_n135_), .Y(mai_mai_n138_));
  NO4        m128(.A(mai_mai_n138_), .B(mai_mai_n134_), .C(mai_mai_n128_), .D(mai_mai_n126_), .Y(mai_mai_n139_));
  AOI220     m129(.A0(i_5_), .A1(mai_mai_n87_), .B0(mai_mai_n62_), .B1(mai_mai_n28_), .Y(mai_mai_n140_));
  AOI210     m130(.A0(mai_mai_n140_), .A1(mai_mai_n119_), .B0(mai_mai_n98_), .Y(mai_mai_n141_));
  NO3        m131(.A(i_2_), .B(mai_mai_n17_), .C(mai_mai_n11_), .Y(mai_mai_n142_));
  NA2        m132(.A(i_2_), .B(i_4_), .Y(mai_mai_n143_));
  AOI210     m133(.A0(mai_mai_n100_), .A1(mai_mai_n84_), .B0(mai_mai_n143_), .Y(mai_mai_n144_));
  NO2        m134(.A(i_8_), .B(i_7_), .Y(mai_mai_n145_));
  OA210      m135(.A0(mai_mai_n144_), .A1(mai_mai_n142_), .B0(mai_mai_n145_), .Y(mai_mai_n146_));
  NA3        m136(.A(mai_mai_n112_), .B(i_0_), .C(mai_mai_n19_), .Y(mai_mai_n147_));
  NO2        m137(.A(mai_mai_n147_), .B(i_4_), .Y(mai_mai_n148_));
  NO3        m138(.A(mai_mai_n148_), .B(mai_mai_n146_), .C(mai_mai_n141_), .Y(mai_mai_n149_));
  NA2        m139(.A(mai_mai_n87_), .B(mai_mai_n12_), .Y(mai_mai_n150_));
  NA2        m140(.A(i_2_), .B(mai_mai_n13_), .Y(mai_mai_n151_));
  NA2        m141(.A(mai_mai_n50_), .B(i_3_), .Y(mai_mai_n152_));
  AOI210     m142(.A0(mai_mai_n152_), .A1(mai_mai_n151_), .B0(mai_mai_n150_), .Y(mai_mai_n153_));
  NA3        m143(.A(mai_mai_n129_), .B(mai_mai_n64_), .C(mai_mai_n102_), .Y(mai_mai_n154_));
  OAI210     m144(.A0(mai_mai_n97_), .A1(mai_mai_n27_), .B0(mai_mai_n154_), .Y(mai_mai_n155_));
  NA4        m145(.A(mai_mai_n103_), .B(mai_mai_n62_), .C(mai_mai_n41_), .D(mai_mai_n17_), .Y(mai_mai_n156_));
  NA3        m146(.A(mai_mai_n53_), .B(mai_mai_n32_), .C(mai_mai_n14_), .Y(mai_mai_n157_));
  NOi31      m147(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n158_));
  OAI210     m148(.A0(mai_mai_n132_), .A1(mai_mai_n77_), .B0(mai_mai_n158_), .Y(mai_mai_n159_));
  NA3        m149(.A(mai_mai_n159_), .B(mai_mai_n157_), .C(mai_mai_n156_), .Y(mai_mai_n160_));
  NO3        m150(.A(mai_mai_n160_), .B(mai_mai_n155_), .C(mai_mai_n153_), .Y(mai_mai_n161_));
  NA4        m151(.A(mai_mai_n161_), .B(mai_mai_n149_), .C(mai_mai_n139_), .D(mai_mai_n124_), .Y(mai_mai_n162_));
  OR4        m152(.A(mai_mai_n162_), .B(mai_mai_n118_), .C(mai_mai_n83_), .D(mai_mai_n68_), .Y(mai00));
  INV        m153(.A(i_2_), .Y(mai_mai_n166_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  AOI210     u014(.A0(men_men_n171_), .A1(men_men_n172_), .B0(men_men_n22_), .Y(men_men_n25_));
  AOI210     u015(.A0(men_men_n25_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n26_));
  NA2        u016(.A(i_0_), .B(men_men_n14_), .Y(men_men_n27_));
  NA2        u017(.A(men_men_n17_), .B(i_5_), .Y(men_men_n28_));
  NO2        u018(.A(i_2_), .B(i_4_), .Y(men_men_n29_));
  NA3        u019(.A(men_men_n29_), .B(i_6_), .C(i_8_), .Y(men_men_n30_));
  AOI210     u020(.A0(men_men_n28_), .A1(men_men_n27_), .B0(men_men_n30_), .Y(men_men_n31_));
  INV        u021(.A(i_2_), .Y(men_men_n32_));
  NOi21      u022(.An(i_5_), .B(i_0_), .Y(men_men_n33_));
  NOi21      u023(.An(i_6_), .B(i_8_), .Y(men_men_n34_));
  NOi21      u024(.An(i_7_), .B(i_1_), .Y(men_men_n35_));
  NOi21      u025(.An(i_5_), .B(i_6_), .Y(men_men_n36_));
  AOI220     u026(.A0(men_men_n36_), .A1(men_men_n35_), .B0(men_men_n34_), .B1(men_men_n33_), .Y(men_men_n37_));
  NO3        u027(.A(men_men_n37_), .B(men_men_n32_), .C(i_4_), .Y(men_men_n38_));
  NOi21      u028(.An(i_0_), .B(i_4_), .Y(men_men_n39_));
  XO2        u029(.A(i_1_), .B(i_3_), .Y(men_men_n40_));
  NOi21      u030(.An(i_7_), .B(i_5_), .Y(men_men_n41_));
  AN3        u031(.A(men_men_n41_), .B(men_men_n40_), .C(men_men_n39_), .Y(men_men_n42_));
  INV        u032(.A(i_1_), .Y(men_men_n43_));
  NOi21      u033(.An(i_3_), .B(i_0_), .Y(men_men_n44_));
  NA2        u034(.A(men_men_n44_), .B(men_men_n43_), .Y(men_men_n45_));
  NO2        u035(.A(men_men_n172_), .B(men_men_n45_), .Y(men_men_n46_));
  NO4        u036(.A(men_men_n46_), .B(men_men_n42_), .C(men_men_n38_), .D(men_men_n31_), .Y(men_men_n47_));
  NOi21      u037(.An(i_4_), .B(i_0_), .Y(men_men_n48_));
  AOI210     u038(.A0(men_men_n48_), .A1(men_men_n24_), .B0(men_men_n15_), .Y(men_men_n49_));
  NA2        u039(.A(i_1_), .B(men_men_n14_), .Y(men_men_n50_));
  NOi21      u040(.An(i_2_), .B(i_8_), .Y(men_men_n51_));
  NO3        u041(.A(men_men_n51_), .B(men_men_n48_), .C(men_men_n39_), .Y(men_men_n52_));
  NO3        u042(.A(men_men_n52_), .B(men_men_n50_), .C(men_men_n49_), .Y(men_men_n53_));
  INV        u043(.A(men_men_n53_), .Y(men_men_n54_));
  NOi31      u044(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n55_));
  NA2        u045(.A(men_men_n55_), .B(i_0_), .Y(men_men_n56_));
  NOi21      u046(.An(i_4_), .B(i_3_), .Y(men_men_n57_));
  NOi21      u047(.An(i_1_), .B(i_4_), .Y(men_men_n58_));
  OAI210     u048(.A0(men_men_n58_), .A1(men_men_n57_), .B0(men_men_n51_), .Y(men_men_n59_));
  NA2        u049(.A(men_men_n59_), .B(men_men_n56_), .Y(men_men_n60_));
  AN2        u050(.A(i_8_), .B(i_7_), .Y(men_men_n61_));
  NA2        u051(.A(men_men_n61_), .B(men_men_n12_), .Y(men_men_n62_));
  NOi21      u052(.An(i_8_), .B(i_7_), .Y(men_men_n63_));
  NA3        u053(.A(men_men_n63_), .B(men_men_n57_), .C(i_6_), .Y(men_men_n64_));
  OAI210     u054(.A0(men_men_n62_), .A1(men_men_n50_), .B0(men_men_n64_), .Y(men_men_n65_));
  AOI220     u055(.A0(men_men_n65_), .A1(men_men_n32_), .B0(men_men_n60_), .B1(men_men_n36_), .Y(men_men_n66_));
  NA4        u056(.A(men_men_n66_), .B(men_men_n54_), .C(men_men_n47_), .D(men_men_n26_), .Y(men_men_n67_));
  NA2        u057(.A(i_8_), .B(i_7_), .Y(men_men_n68_));
  NO3        u058(.A(men_men_n68_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n69_));
  NA2        u059(.A(i_8_), .B(men_men_n23_), .Y(men_men_n70_));
  NA2        u060(.A(men_men_n40_), .B(i_2_), .Y(men_men_n71_));
  NOi21      u061(.An(i_1_), .B(i_2_), .Y(men_men_n72_));
  NA3        u062(.A(men_men_n72_), .B(men_men_n48_), .C(i_6_), .Y(men_men_n73_));
  OAI210     u063(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n73_), .Y(men_men_n74_));
  OAI210     u064(.A0(men_men_n74_), .A1(men_men_n69_), .B0(men_men_n14_), .Y(men_men_n75_));
  NA3        u065(.A(men_men_n63_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n76_));
  NA3        u066(.A(i_1_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n77_));
  NA2        u067(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NOi32      u068(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n79_));
  NA2        u069(.A(men_men_n79_), .B(i_3_), .Y(men_men_n80_));
  NA3        u070(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n81_));
  NA2        u071(.A(men_men_n81_), .B(men_men_n80_), .Y(men_men_n82_));
  NO2        u072(.A(i_0_), .B(i_4_), .Y(men_men_n83_));
  AOI220     u073(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n78_), .B1(men_men_n57_), .Y(men_men_n84_));
  NA2        u074(.A(men_men_n84_), .B(men_men_n75_), .Y(men_men_n85_));
  INV        u075(.A(i_6_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n87_));
  NOi21      u077(.An(i_7_), .B(i_8_), .Y(men_men_n88_));
  NOi31      u078(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n89_));
  AOI210     u079(.A0(men_men_n88_), .A1(men_men_n12_), .B0(men_men_n89_), .Y(men_men_n90_));
  OAI210     u080(.A0(men_men_n90_), .A1(men_men_n11_), .B0(men_men_n87_), .Y(men_men_n91_));
  NA2        u081(.A(men_men_n91_), .B(men_men_n72_), .Y(men_men_n92_));
  NA3        u082(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n93_));
  NO2        u083(.A(men_men_n22_), .B(men_men_n93_), .Y(men_men_n94_));
  NA2        u084(.A(i_4_), .B(i_5_), .Y(men_men_n95_));
  NA3        u085(.A(men_men_n68_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n96_));
  NO2        u086(.A(men_men_n96_), .B(men_men_n95_), .Y(men_men_n97_));
  NO2        u087(.A(men_men_n97_), .B(men_men_n94_), .Y(men_men_n98_));
  NA3        u088(.A(men_men_n63_), .B(men_men_n32_), .C(i_3_), .Y(men_men_n99_));
  NA2        u089(.A(men_men_n43_), .B(i_6_), .Y(men_men_n100_));
  AOI210     u090(.A0(men_men_n100_), .A1(men_men_n22_), .B0(men_men_n99_), .Y(men_men_n101_));
  NOi21      u091(.An(i_2_), .B(i_1_), .Y(men_men_n102_));
  NAi21      u092(.An(i_6_), .B(i_0_), .Y(men_men_n103_));
  NOi21      u093(.An(i_4_), .B(i_6_), .Y(men_men_n104_));
  NOi21      u094(.An(i_5_), .B(i_3_), .Y(men_men_n105_));
  NA3        u095(.A(men_men_n105_), .B(men_men_n72_), .C(men_men_n104_), .Y(men_men_n106_));
  INV        u096(.A(men_men_n106_), .Y(men_men_n107_));
  NA2        u097(.A(men_men_n72_), .B(men_men_n34_), .Y(men_men_n108_));
  NOi21      u098(.An(men_men_n41_), .B(men_men_n108_), .Y(men_men_n109_));
  NO3        u099(.A(men_men_n109_), .B(men_men_n107_), .C(men_men_n101_), .Y(men_men_n110_));
  NOi21      u100(.An(i_6_), .B(i_1_), .Y(men_men_n111_));
  AOI220     u101(.A0(men_men_n111_), .A1(i_7_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n112_));
  NOi31      u102(.An(men_men_n48_), .B(men_men_n112_), .C(i_2_), .Y(men_men_n113_));
  NA2        u103(.A(men_men_n63_), .B(men_men_n12_), .Y(men_men_n114_));
  NA2        u104(.A(men_men_n34_), .B(men_men_n14_), .Y(men_men_n115_));
  NOi21      u105(.An(i_3_), .B(i_1_), .Y(men_men_n116_));
  NA2        u106(.A(men_men_n116_), .B(i_4_), .Y(men_men_n117_));
  AOI210     u107(.A0(men_men_n115_), .A1(men_men_n114_), .B0(men_men_n117_), .Y(men_men_n118_));
  AOI220     u108(.A0(men_men_n88_), .A1(men_men_n14_), .B0(men_men_n104_), .B1(men_men_n23_), .Y(men_men_n119_));
  NOi31      u109(.An(men_men_n44_), .B(men_men_n119_), .C(men_men_n32_), .Y(men_men_n120_));
  NO3        u110(.A(men_men_n120_), .B(men_men_n118_), .C(men_men_n113_), .Y(men_men_n121_));
  NA4        u111(.A(men_men_n121_), .B(men_men_n110_), .C(men_men_n98_), .D(men_men_n92_), .Y(men_men_n122_));
  NA2        u112(.A(men_men_n51_), .B(men_men_n15_), .Y(men_men_n123_));
  NOi31      u113(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n124_));
  NOi31      u114(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n125_));
  OAI210     u115(.A0(men_men_n125_), .A1(men_men_n124_), .B0(i_7_), .Y(men_men_n126_));
  NA3        u116(.A(men_men_n34_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n127_));
  NA4        u117(.A(men_men_n127_), .B(men_men_n126_), .C(men_men_n123_), .D(men_men_n108_), .Y(men_men_n128_));
  NA2        u118(.A(men_men_n128_), .B(men_men_n39_), .Y(men_men_n129_));
  NO2        u119(.A(men_men_n76_), .B(men_men_n28_), .Y(men_men_n130_));
  NA3        u120(.A(men_men_n61_), .B(men_men_n102_), .C(men_men_n17_), .Y(men_men_n131_));
  NAi31      u121(.An(men_men_n103_), .B(men_men_n88_), .C(men_men_n102_), .Y(men_men_n132_));
  NA3        u122(.A(men_men_n63_), .B(men_men_n55_), .C(i_6_), .Y(men_men_n133_));
  NA3        u123(.A(men_men_n133_), .B(men_men_n132_), .C(men_men_n131_), .Y(men_men_n134_));
  NOi21      u124(.An(i_0_), .B(i_2_), .Y(men_men_n135_));
  NA3        u125(.A(men_men_n135_), .B(men_men_n35_), .C(men_men_n104_), .Y(men_men_n136_));
  NA3        u126(.A(men_men_n48_), .B(men_men_n41_), .C(men_men_n18_), .Y(men_men_n137_));
  NOi32      u127(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n138_));
  NA2        u128(.A(men_men_n138_), .B(men_men_n124_), .Y(men_men_n139_));
  NA3        u129(.A(men_men_n135_), .B(men_men_n57_), .C(men_men_n34_), .Y(men_men_n140_));
  NA4        u130(.A(men_men_n140_), .B(men_men_n139_), .C(men_men_n137_), .D(men_men_n136_), .Y(men_men_n141_));
  NA4        u131(.A(men_men_n55_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n142_));
  NA3        u132(.A(men_men_n58_), .B(men_men_n17_), .C(i_8_), .Y(men_men_n143_));
  NA2        u133(.A(men_men_n143_), .B(men_men_n142_), .Y(men_men_n144_));
  NO4        u134(.A(men_men_n144_), .B(men_men_n141_), .C(men_men_n134_), .D(men_men_n130_), .Y(men_men_n145_));
  NOi21      u135(.An(i_5_), .B(i_2_), .Y(men_men_n146_));
  AOI220     u136(.A0(men_men_n146_), .A1(men_men_n88_), .B0(men_men_n61_), .B1(men_men_n29_), .Y(men_men_n147_));
  AOI210     u137(.A0(men_men_n147_), .A1(men_men_n123_), .B0(men_men_n100_), .Y(men_men_n148_));
  NO3        u138(.A(i_2_), .B(men_men_n11_), .C(men_men_n14_), .Y(men_men_n149_));
  NA2        u139(.A(i_2_), .B(i_4_), .Y(men_men_n150_));
  AOI210     u140(.A0(men_men_n103_), .A1(men_men_n86_), .B0(men_men_n150_), .Y(men_men_n151_));
  NO2        u141(.A(i_8_), .B(i_7_), .Y(men_men_n152_));
  OA210      u142(.A0(men_men_n151_), .A1(men_men_n149_), .B0(men_men_n152_), .Y(men_men_n153_));
  NA3        u143(.A(men_men_n116_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n154_));
  NO2        u144(.A(men_men_n154_), .B(i_4_), .Y(men_men_n155_));
  NO3        u145(.A(men_men_n155_), .B(men_men_n153_), .C(men_men_n148_), .Y(men_men_n156_));
  NA2        u146(.A(men_men_n88_), .B(men_men_n12_), .Y(men_men_n157_));
  NA3        u147(.A(i_2_), .B(i_1_), .C(men_men_n14_), .Y(men_men_n158_));
  INV        u148(.A(men_men_n48_), .Y(men_men_n159_));
  AOI210     u149(.A0(men_men_n159_), .A1(men_men_n158_), .B0(men_men_n157_), .Y(men_men_n160_));
  NA3        u150(.A(men_men_n135_), .B(men_men_n63_), .C(men_men_n104_), .Y(men_men_n161_));
  OAI210     u151(.A0(men_men_n99_), .A1(men_men_n28_), .B0(men_men_n161_), .Y(men_men_n162_));
  NOi31      u152(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n163_));
  OAI210     u153(.A0(men_men_n138_), .A1(men_men_n79_), .B0(men_men_n163_), .Y(men_men_n164_));
  INV        u154(.A(men_men_n164_), .Y(men_men_n165_));
  NO3        u155(.A(men_men_n165_), .B(men_men_n162_), .C(men_men_n160_), .Y(men_men_n166_));
  NA4        u156(.A(men_men_n166_), .B(men_men_n156_), .C(men_men_n145_), .D(men_men_n129_), .Y(men_men_n167_));
  OR4        u157(.A(men_men_n167_), .B(men_men_n122_), .C(men_men_n85_), .D(men_men_n67_), .Y(men00));
  INV        u158(.A(i_1_), .Y(men_men_n171_));
  INV        u159(.A(i_5_), .Y(men_men_n172_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule