// Benchmark "top" written by ABC on Fri Jun 21 17:49:29 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n132_, new_new_n133_, new_new_n134_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n962_, new_new_n963_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g021(.A(new_new_n35_), .Y(mai1));
  INV        g022(.A(i_11_), .Y(new_new_n45_));
  NO2        g023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g024(.A(i_2_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NA3        g030(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n53_));
  NO2        g031(.A(i_1_), .B(i_6_), .Y(new_new_n54_));
  NA2        g032(.A(i_8_), .B(i_7_), .Y(new_new_n55_));
  OAI210     g033(.A0(new_new_n55_), .A1(new_new_n54_), .B0(new_new_n53_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n56_), .B(i_12_), .Y(new_new_n57_));
  NAi21      g035(.An(i_2_), .B(i_7_), .Y(new_new_n58_));
  INV        g036(.A(i_1_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_6_), .Y(new_new_n60_));
  NA3        g038(.A(new_new_n60_), .B(new_new_n58_), .C(new_new_n31_), .Y(new_new_n61_));
  NA2        g039(.A(i_1_), .B(i_10_), .Y(new_new_n62_));
  NO2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NAi31      g041(.An(new_new_n63_), .B(new_new_n61_), .C(new_new_n57_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n50_), .B(i_2_), .Y(new_new_n65_));
  AOI210     g043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_6_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(new_new_n25_), .Y(new_new_n68_));
  INV        g046(.A(i_0_), .Y(new_new_n69_));
  NAi21      g047(.An(i_5_), .B(i_10_), .Y(new_new_n70_));
  NA2        g048(.A(i_5_), .B(i_9_), .Y(new_new_n71_));
  AOI210     g049(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n69_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n72_), .B(new_new_n68_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n66_), .A1(new_new_n65_), .B0(new_new_n73_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n74_), .A1(new_new_n64_), .B0(i_0_), .Y(new_new_n75_));
  NA2        g053(.A(i_12_), .B(i_5_), .Y(new_new_n76_));
  NA2        g054(.A(i_2_), .B(i_8_), .Y(new_new_n77_));
  NO2        g055(.A(new_new_n77_), .B(new_new_n54_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_9_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_7_), .Y(new_new_n80_));
  NO3        g058(.A(new_new_n80_), .B(new_new_n79_), .C(new_new_n59_), .Y(new_new_n81_));
  INV        g059(.A(i_6_), .Y(new_new_n82_));
  OR4        g060(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n83_));
  INV        g061(.A(new_new_n83_), .Y(new_new_n84_));
  NO2        g062(.A(i_2_), .B(i_7_), .Y(new_new_n85_));
  OAI210     g063(.A0(new_new_n81_), .A1(new_new_n78_), .B0(i_2_), .Y(new_new_n86_));
  NAi21      g064(.An(i_6_), .B(i_10_), .Y(new_new_n87_));
  NA2        g065(.A(i_6_), .B(i_9_), .Y(new_new_n88_));
  AOI210     g066(.A0(new_new_n88_), .A1(new_new_n87_), .B0(new_new_n59_), .Y(new_new_n89_));
  NA2        g067(.A(i_2_), .B(i_6_), .Y(new_new_n90_));
  INV        g068(.A(new_new_n89_), .Y(new_new_n91_));
  AOI210     g069(.A0(new_new_n91_), .A1(new_new_n86_), .B0(new_new_n76_), .Y(new_new_n92_));
  AN3        g070(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n93_));
  NAi21      g071(.An(i_6_), .B(i_11_), .Y(new_new_n94_));
  NO2        g072(.A(i_5_), .B(i_8_), .Y(new_new_n95_));
  NOi21      g073(.An(new_new_n95_), .B(new_new_n94_), .Y(new_new_n96_));
  AOI220     g074(.A0(new_new_n96_), .A1(new_new_n58_), .B0(new_new_n93_), .B1(new_new_n32_), .Y(new_new_n97_));
  INV        g075(.A(i_7_), .Y(new_new_n98_));
  NA2        g076(.A(new_new_n47_), .B(new_new_n98_), .Y(new_new_n99_));
  NO2        g077(.A(i_0_), .B(i_5_), .Y(new_new_n100_));
  NO2        g078(.A(new_new_n100_), .B(new_new_n82_), .Y(new_new_n101_));
  NA2        g079(.A(i_12_), .B(i_3_), .Y(new_new_n102_));
  INV        g080(.A(new_new_n102_), .Y(new_new_n103_));
  NA3        g081(.A(new_new_n103_), .B(new_new_n101_), .C(new_new_n99_), .Y(new_new_n104_));
  NAi21      g082(.An(i_7_), .B(i_11_), .Y(new_new_n105_));
  AN2        g083(.A(i_2_), .B(i_10_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(i_7_), .Y(new_new_n107_));
  OR2        g085(.A(new_new_n76_), .B(new_new_n54_), .Y(new_new_n108_));
  NO2        g086(.A(i_8_), .B(new_new_n98_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n108_), .C(new_new_n107_), .Y(new_new_n110_));
  NA2        g088(.A(i_12_), .B(i_7_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n59_), .B(new_new_n26_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n112_), .B(i_0_), .Y(new_new_n113_));
  NA2        g091(.A(i_11_), .B(i_12_), .Y(new_new_n114_));
  OAI210     g092(.A0(new_new_n113_), .A1(new_new_n111_), .B0(new_new_n114_), .Y(new_new_n115_));
  NO2        g093(.A(new_new_n115_), .B(new_new_n110_), .Y(new_new_n116_));
  NA3        g094(.A(new_new_n116_), .B(new_new_n104_), .C(new_new_n97_), .Y(new_new_n117_));
  NOi21      g095(.An(i_1_), .B(i_5_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n118_), .B(i_11_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n98_), .B(new_new_n37_), .Y(new_new_n120_));
  NA2        g098(.A(i_7_), .B(new_new_n25_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n121_), .B(new_new_n120_), .Y(new_new_n122_));
  NO2        g100(.A(new_new_n122_), .B(new_new_n47_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n88_), .B(new_new_n87_), .Y(new_new_n124_));
  INV        g102(.A(new_new_n124_), .Y(new_new_n125_));
  NO2        g103(.A(i_1_), .B(new_new_n82_), .Y(new_new_n126_));
  NO2        g104(.A(i_6_), .B(i_5_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(i_3_), .Y(new_new_n128_));
  OAI220     g106(.A0(new_new_n128_), .A1(new_new_n105_), .B0(new_new_n125_), .B1(new_new_n119_), .Y(new_new_n129_));
  NO3        g107(.A(new_new_n129_), .B(new_new_n117_), .C(new_new_n92_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n75_), .Y(mai2));
  NO2        g109(.A(new_new_n59_), .B(new_new_n37_), .Y(new_new_n132_));
  NA2        g110(.A(i_6_), .B(new_new_n25_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(new_new_n132_), .Y(new_new_n134_));
  NA4        g112(.A(new_new_n134_), .B(new_new_n73_), .C(new_new_n65_), .D(new_new_n30_), .Y(mai0));
  AN2        g113(.A(i_8_), .B(i_7_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(i_6_), .Y(new_new_n137_));
  NO2        g115(.A(i_12_), .B(i_13_), .Y(new_new_n138_));
  NAi21      g116(.An(i_5_), .B(i_11_), .Y(new_new_n139_));
  NOi21      g117(.An(new_new_n138_), .B(new_new_n139_), .Y(new_new_n140_));
  NO2        g118(.A(i_0_), .B(i_1_), .Y(new_new_n141_));
  NA2        g119(.A(i_2_), .B(i_3_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n142_), .B(i_4_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(new_new_n140_), .Y(new_new_n144_));
  AN2        g122(.A(new_new_n138_), .B(new_new_n79_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(new_new_n27_), .Y(new_new_n146_));
  NA2        g124(.A(i_1_), .B(i_5_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n69_), .B(new_new_n47_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n36_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  OR2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NO3        g129(.A(new_new_n151_), .B(new_new_n76_), .C(i_13_), .Y(new_new_n152_));
  NAi32      g130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n153_));
  NAi21      g131(.An(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  NOi21      g132(.An(i_4_), .B(i_10_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n40_), .Y(new_new_n156_));
  NO2        g134(.A(i_3_), .B(i_5_), .Y(new_new_n157_));
  NO3        g135(.A(new_new_n69_), .B(i_2_), .C(i_1_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n157_), .Y(new_new_n159_));
  OAI210     g137(.A0(new_new_n159_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n160_), .B(new_new_n150_), .Y(new_new_n161_));
  AOI210     g139(.A0(new_new_n161_), .A1(new_new_n144_), .B0(new_new_n137_), .Y(new_new_n162_));
  NA3        g140(.A(new_new_n69_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n163_));
  NOi21      g141(.An(i_4_), .B(i_9_), .Y(new_new_n164_));
  NOi21      g142(.An(i_11_), .B(i_13_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  NO2        g144(.A(i_4_), .B(i_5_), .Y(new_new_n167_));
  NAi21      g145(.An(i_12_), .B(i_11_), .Y(new_new_n168_));
  NO2        g146(.A(new_new_n168_), .B(i_13_), .Y(new_new_n169_));
  NA3        g147(.A(new_new_n169_), .B(new_new_n167_), .C(new_new_n79_), .Y(new_new_n170_));
  AOI210     g148(.A0(new_new_n170_), .A1(new_new_n166_), .B0(new_new_n163_), .Y(new_new_n171_));
  NO2        g149(.A(new_new_n69_), .B(new_new_n59_), .Y(new_new_n172_));
  INV        g150(.A(new_new_n172_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n36_), .B(i_5_), .Y(new_new_n174_));
  NAi31      g152(.An(new_new_n174_), .B(new_new_n145_), .C(i_11_), .Y(new_new_n175_));
  NA2        g153(.A(i_3_), .B(i_5_), .Y(new_new_n176_));
  OR2        g154(.A(new_new_n176_), .B(new_new_n166_), .Y(new_new_n177_));
  AOI210     g155(.A0(new_new_n177_), .A1(new_new_n175_), .B0(new_new_n173_), .Y(new_new_n178_));
  NO2        g156(.A(new_new_n69_), .B(i_5_), .Y(new_new_n179_));
  NO2        g157(.A(i_13_), .B(i_10_), .Y(new_new_n180_));
  NA3        g158(.A(new_new_n180_), .B(new_new_n179_), .C(new_new_n45_), .Y(new_new_n181_));
  NO2        g159(.A(i_2_), .B(i_1_), .Y(new_new_n182_));
  NAi21      g160(.An(i_4_), .B(i_12_), .Y(new_new_n183_));
  NO3        g161(.A(new_new_n183_), .B(i_2_), .C(new_new_n181_), .Y(new_new_n184_));
  NO3        g162(.A(new_new_n184_), .B(new_new_n178_), .C(new_new_n171_), .Y(new_new_n185_));
  INV        g163(.A(i_8_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n186_), .B(i_7_), .Y(new_new_n187_));
  NA2        g165(.A(new_new_n187_), .B(i_6_), .Y(new_new_n188_));
  NO3        g166(.A(i_3_), .B(new_new_n82_), .C(new_new_n48_), .Y(new_new_n189_));
  NA2        g167(.A(new_new_n189_), .B(new_new_n109_), .Y(new_new_n190_));
  NO3        g168(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n191_));
  NA3        g169(.A(new_new_n191_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n192_));
  NO3        g170(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n193_));
  OAI210     g171(.A0(new_new_n93_), .A1(i_12_), .B0(new_new_n193_), .Y(new_new_n194_));
  AOI210     g172(.A0(new_new_n194_), .A1(new_new_n192_), .B0(new_new_n190_), .Y(new_new_n195_));
  NO2        g173(.A(i_3_), .B(i_8_), .Y(new_new_n196_));
  NO3        g174(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n197_));
  NA3        g175(.A(new_new_n197_), .B(new_new_n196_), .C(new_new_n40_), .Y(new_new_n198_));
  NO2        g176(.A(new_new_n100_), .B(new_new_n54_), .Y(new_new_n199_));
  NO2        g177(.A(i_13_), .B(i_9_), .Y(new_new_n200_));
  NA3        g178(.A(new_new_n200_), .B(i_6_), .C(new_new_n186_), .Y(new_new_n201_));
  NAi21      g179(.An(i_12_), .B(i_3_), .Y(new_new_n202_));
  BUFFER     g180(.A(new_new_n201_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n45_), .B(i_5_), .Y(new_new_n204_));
  NO3        g182(.A(i_0_), .B(i_2_), .C(new_new_n59_), .Y(new_new_n205_));
  NA3        g183(.A(new_new_n205_), .B(new_new_n204_), .C(i_10_), .Y(new_new_n206_));
  OAI220     g184(.A0(new_new_n206_), .A1(new_new_n203_), .B0(new_new_n100_), .B1(new_new_n198_), .Y(new_new_n207_));
  AOI210     g185(.A0(new_new_n207_), .A1(i_7_), .B0(new_new_n195_), .Y(new_new_n208_));
  OAI220     g186(.A0(new_new_n208_), .A1(i_4_), .B0(new_new_n188_), .B1(new_new_n185_), .Y(new_new_n209_));
  NAi21      g187(.An(i_12_), .B(i_7_), .Y(new_new_n210_));
  NA3        g188(.A(i_13_), .B(new_new_n186_), .C(i_10_), .Y(new_new_n211_));
  NA2        g189(.A(i_0_), .B(i_5_), .Y(new_new_n212_));
  NAi31      g190(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n36_), .B(i_13_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n69_), .B(new_new_n26_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n47_), .B(new_new_n59_), .Y(new_new_n216_));
  INV        g194(.A(i_13_), .Y(new_new_n217_));
  NO2        g195(.A(i_12_), .B(new_new_n217_), .Y(new_new_n218_));
  NO2        g196(.A(i_12_), .B(new_new_n37_), .Y(new_new_n219_));
  NO2        g197(.A(new_new_n176_), .B(i_4_), .Y(new_new_n220_));
  NA2        g198(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n221_));
  OR2        g199(.A(i_8_), .B(i_7_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n222_), .B(new_new_n82_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n51_), .B(i_1_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n224_), .B(new_new_n223_), .Y(new_new_n225_));
  INV        g203(.A(i_12_), .Y(new_new_n226_));
  NO3        g204(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n227_));
  NA2        g205(.A(i_2_), .B(i_1_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n225_), .B(new_new_n221_), .Y(new_new_n229_));
  NAi21      g207(.An(i_4_), .B(i_3_), .Y(new_new_n230_));
  INV        g208(.A(new_new_n71_), .Y(new_new_n231_));
  NO2        g209(.A(i_0_), .B(i_6_), .Y(new_new_n232_));
  NOi41      g210(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n233_));
  NA2        g211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  NAi21      g212(.An(new_new_n234_), .B(i_5_), .Y(new_new_n235_));
  INV        g213(.A(new_new_n235_), .Y(new_new_n236_));
  AOI210     g214(.A0(new_new_n236_), .A1(new_new_n40_), .B0(new_new_n229_), .Y(new_new_n237_));
  NO2        g215(.A(i_11_), .B(new_new_n217_), .Y(new_new_n238_));
  NOi21      g216(.An(i_1_), .B(i_6_), .Y(new_new_n239_));
  NAi21      g217(.An(i_3_), .B(i_7_), .Y(new_new_n240_));
  NA2        g218(.A(new_new_n226_), .B(i_9_), .Y(new_new_n241_));
  OR4        g219(.A(new_new_n241_), .B(new_new_n240_), .C(new_new_n239_), .D(new_new_n179_), .Y(new_new_n242_));
  NO2        g220(.A(i_12_), .B(i_3_), .Y(new_new_n243_));
  NA2        g221(.A(new_new_n69_), .B(i_5_), .Y(new_new_n244_));
  NA2        g222(.A(i_3_), .B(i_9_), .Y(new_new_n245_));
  NAi21      g223(.An(i_7_), .B(i_10_), .Y(new_new_n246_));
  NO2        g224(.A(new_new_n246_), .B(new_new_n245_), .Y(new_new_n247_));
  NA3        g225(.A(new_new_n247_), .B(new_new_n244_), .C(new_new_n60_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n248_), .B(new_new_n242_), .Y(new_new_n249_));
  NA3        g227(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n250_));
  INV        g228(.A(new_new_n137_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n226_), .B(i_13_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n252_), .B(new_new_n71_), .Y(new_new_n253_));
  AOI220     g231(.A0(new_new_n253_), .A1(new_new_n251_), .B0(new_new_n249_), .B1(new_new_n238_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n222_), .B(new_new_n37_), .Y(new_new_n255_));
  NA2        g233(.A(i_12_), .B(i_6_), .Y(new_new_n256_));
  OR2        g234(.A(i_13_), .B(i_9_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n230_), .B(i_2_), .Y(new_new_n258_));
  NA2        g236(.A(new_new_n238_), .B(i_9_), .Y(new_new_n259_));
  NA2        g237(.A(new_new_n148_), .B(new_new_n59_), .Y(new_new_n260_));
  NO3        g238(.A(i_11_), .B(new_new_n217_), .C(new_new_n25_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n240_), .B(i_8_), .Y(new_new_n262_));
  NA3        g240(.A(i_5_), .B(new_new_n262_), .C(new_new_n261_), .Y(new_new_n263_));
  NA3        g241(.A(i_6_), .B(new_new_n255_), .C(new_new_n218_), .Y(new_new_n264_));
  AOI210     g242(.A0(new_new_n264_), .A1(new_new_n263_), .B0(new_new_n260_), .Y(new_new_n265_));
  INV        g243(.A(new_new_n265_), .Y(new_new_n266_));
  NA3        g244(.A(new_new_n266_), .B(new_new_n254_), .C(new_new_n237_), .Y(new_new_n267_));
  NO3        g245(.A(i_12_), .B(new_new_n217_), .C(new_new_n37_), .Y(new_new_n268_));
  INV        g246(.A(new_new_n268_), .Y(new_new_n269_));
  NA2        g247(.A(i_8_), .B(new_new_n98_), .Y(new_new_n270_));
  NOi21      g248(.An(new_new_n157_), .B(new_new_n82_), .Y(new_new_n271_));
  NO3        g249(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n272_));
  AOI220     g250(.A0(new_new_n272_), .A1(new_new_n189_), .B0(new_new_n271_), .B1(new_new_n224_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n273_), .B(new_new_n270_), .Y(new_new_n274_));
  NO3        g252(.A(i_0_), .B(i_2_), .C(new_new_n59_), .Y(new_new_n275_));
  NO2        g253(.A(new_new_n228_), .B(i_0_), .Y(new_new_n276_));
  AOI220     g254(.A0(new_new_n276_), .A1(new_new_n187_), .B0(new_new_n275_), .B1(new_new_n136_), .Y(new_new_n277_));
  NA2        g255(.A(i_5_), .B(new_new_n26_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n278_), .B(new_new_n277_), .Y(new_new_n279_));
  NA2        g257(.A(i_0_), .B(i_1_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(i_2_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n55_), .B(i_6_), .Y(new_new_n282_));
  NA3        g260(.A(new_new_n282_), .B(new_new_n281_), .C(new_new_n157_), .Y(new_new_n283_));
  OAI210     g261(.A0(new_new_n159_), .A1(new_new_n137_), .B0(new_new_n283_), .Y(new_new_n284_));
  NO3        g262(.A(new_new_n284_), .B(new_new_n279_), .C(new_new_n274_), .Y(new_new_n285_));
  NO2        g263(.A(i_3_), .B(i_10_), .Y(new_new_n286_));
  NA3        g264(.A(new_new_n286_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n287_));
  NO2        g265(.A(i_2_), .B(new_new_n98_), .Y(new_new_n288_));
  NO2        g266(.A(i_4_), .B(i_8_), .Y(new_new_n289_));
  NOi21      g267(.An(new_new_n212_), .B(new_new_n100_), .Y(new_new_n290_));
  NA3        g268(.A(new_new_n290_), .B(new_new_n289_), .C(new_new_n288_), .Y(new_new_n291_));
  AN2        g269(.A(i_3_), .B(i_10_), .Y(new_new_n292_));
  NA4        g270(.A(new_new_n292_), .B(new_new_n191_), .C(new_new_n169_), .D(new_new_n167_), .Y(new_new_n293_));
  NO2        g271(.A(i_5_), .B(new_new_n37_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n295_));
  OR2        g273(.A(new_new_n291_), .B(new_new_n287_), .Y(new_new_n296_));
  OAI220     g274(.A0(new_new_n296_), .A1(i_6_), .B0(new_new_n285_), .B1(new_new_n269_), .Y(new_new_n297_));
  NO4        g275(.A(new_new_n297_), .B(new_new_n267_), .C(new_new_n209_), .D(new_new_n162_), .Y(new_new_n298_));
  NO3        g276(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n55_), .B(new_new_n82_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n276_), .B(new_new_n300_), .Y(new_new_n301_));
  NO3        g279(.A(i_6_), .B(new_new_n186_), .C(i_7_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n302_), .B(new_new_n191_), .Y(new_new_n303_));
  AOI210     g281(.A0(new_new_n303_), .A1(new_new_n301_), .B0(i_5_), .Y(new_new_n304_));
  NO2        g282(.A(i_2_), .B(i_3_), .Y(new_new_n305_));
  NA3        g283(.A(new_new_n223_), .B(new_new_n305_), .C(i_1_), .Y(new_new_n306_));
  NA3        g284(.A(new_new_n276_), .B(new_new_n271_), .C(new_new_n109_), .Y(new_new_n307_));
  NO2        g285(.A(i_8_), .B(i_6_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n151_), .B(new_new_n47_), .Y(new_new_n309_));
  NA3        g287(.A(new_new_n309_), .B(new_new_n308_), .C(new_new_n157_), .Y(new_new_n310_));
  NA3        g288(.A(new_new_n310_), .B(new_new_n307_), .C(new_new_n306_), .Y(new_new_n311_));
  OAI210     g289(.A0(new_new_n311_), .A1(new_new_n304_), .B0(i_4_), .Y(new_new_n312_));
  NO2        g290(.A(i_12_), .B(i_10_), .Y(new_new_n313_));
  NOi21      g291(.An(i_5_), .B(i_0_), .Y(new_new_n314_));
  NA4        g292(.A(new_new_n80_), .B(new_new_n36_), .C(new_new_n82_), .D(i_8_), .Y(new_new_n315_));
  NO2        g293(.A(i_6_), .B(i_8_), .Y(new_new_n316_));
  AN2        g294(.A(i_0_), .B(new_new_n316_), .Y(new_new_n317_));
  NO2        g295(.A(i_1_), .B(i_7_), .Y(new_new_n318_));
  NA3        g296(.A(new_new_n316_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n319_));
  NA2        g297(.A(new_new_n319_), .B(new_new_n312_), .Y(new_new_n320_));
  NO3        g298(.A(new_new_n222_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n321_));
  NO3        g299(.A(i_8_), .B(i_2_), .C(i_1_), .Y(new_new_n322_));
  OAI210     g300(.A0(new_new_n322_), .A1(new_new_n321_), .B0(i_6_), .Y(new_new_n323_));
  INV        g301(.A(new_new_n323_), .Y(new_new_n324_));
  NOi21      g302(.An(new_new_n147_), .B(new_new_n101_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n325_), .B(new_new_n121_), .Y(new_new_n326_));
  OAI210     g304(.A0(new_new_n326_), .A1(new_new_n324_), .B0(i_3_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n280_), .B(new_new_n77_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n328_), .B(new_new_n127_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n90_), .B(new_new_n186_), .Y(new_new_n330_));
  NA3        g308(.A(new_new_n290_), .B(new_new_n330_), .C(new_new_n59_), .Y(new_new_n331_));
  AOI210     g309(.A0(new_new_n331_), .A1(new_new_n329_), .B0(i_7_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n186_), .B(i_9_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n333_), .B(new_new_n199_), .Y(new_new_n334_));
  NO2        g312(.A(new_new_n334_), .B(new_new_n47_), .Y(new_new_n335_));
  NO3        g313(.A(new_new_n335_), .B(new_new_n332_), .C(new_new_n279_), .Y(new_new_n336_));
  AOI210     g314(.A0(new_new_n336_), .A1(new_new_n327_), .B0(new_new_n156_), .Y(new_new_n337_));
  AOI210     g315(.A0(new_new_n320_), .A1(new_new_n299_), .B0(new_new_n337_), .Y(new_new_n338_));
  NOi32      g316(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n339_));
  INV        g317(.A(new_new_n339_), .Y(new_new_n340_));
  NAi21      g318(.An(i_1_), .B(i_5_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n341_), .B(i_0_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n342_), .B(new_new_n25_), .Y(new_new_n343_));
  OAI210     g321(.A0(new_new_n343_), .A1(new_new_n153_), .B0(new_new_n234_), .Y(new_new_n344_));
  NAi41      g322(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n345_));
  OAI220     g323(.A0(new_new_n345_), .A1(new_new_n341_), .B0(new_new_n213_), .B1(new_new_n153_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n153_), .B(new_new_n151_), .Y(new_new_n347_));
  NOi32      g325(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n348_));
  NAi21      g326(.An(i_6_), .B(i_1_), .Y(new_new_n349_));
  NA3        g327(.A(new_new_n349_), .B(new_new_n348_), .C(new_new_n47_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n350_), .B(i_0_), .Y(new_new_n351_));
  OR3        g329(.A(new_new_n351_), .B(new_new_n347_), .C(new_new_n346_), .Y(new_new_n352_));
  NO2        g330(.A(i_1_), .B(new_new_n98_), .Y(new_new_n353_));
  NAi21      g331(.An(i_3_), .B(i_4_), .Y(new_new_n354_));
  NO2        g332(.A(new_new_n354_), .B(i_9_), .Y(new_new_n355_));
  AN2        g333(.A(i_6_), .B(i_7_), .Y(new_new_n356_));
  NA2        g334(.A(i_2_), .B(i_7_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n354_), .B(i_10_), .Y(new_new_n358_));
  NA3        g336(.A(new_new_n358_), .B(new_new_n357_), .C(new_new_n232_), .Y(new_new_n359_));
  INV        g337(.A(new_new_n359_), .Y(new_new_n360_));
  AOI220     g338(.A0(new_new_n358_), .A1(new_new_n318_), .B0(new_new_n227_), .B1(new_new_n182_), .Y(new_new_n361_));
  NO3        g339(.A(new_new_n360_), .B(new_new_n352_), .C(new_new_n344_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n362_), .B(new_new_n340_), .Y(new_new_n363_));
  AN2        g341(.A(i_12_), .B(i_5_), .Y(new_new_n364_));
  NO2        g342(.A(i_11_), .B(i_6_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n230_), .B(i_5_), .Y(new_new_n366_));
  NO2        g344(.A(i_5_), .B(i_10_), .Y(new_new_n367_));
  AOI220     g345(.A0(new_new_n367_), .A1(new_new_n258_), .B0(new_new_n366_), .B1(new_new_n191_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n138_), .B(new_new_n46_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n369_), .B(new_new_n368_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n370_), .B(i_7_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n372_));
  NO3        g350(.A(new_new_n82_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n373_));
  INV        g351(.A(i_3_), .Y(new_new_n374_));
  NA3        g352(.A(new_new_n286_), .B(new_new_n88_), .C(new_new_n52_), .Y(new_new_n375_));
  NO2        g353(.A(i_11_), .B(i_12_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n376_), .B(new_new_n36_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n375_), .B(new_new_n377_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n42_), .B(i_11_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n213_), .Y(new_new_n380_));
  NAi21      g358(.An(i_13_), .B(i_0_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n381_), .B(new_new_n228_), .Y(new_new_n382_));
  OAI210     g360(.A0(new_new_n380_), .A1(new_new_n378_), .B0(new_new_n382_), .Y(new_new_n383_));
  NA2        g361(.A(new_new_n383_), .B(new_new_n371_), .Y(new_new_n384_));
  NO3        g362(.A(i_1_), .B(i_12_), .C(new_new_n82_), .Y(new_new_n385_));
  NO2        g363(.A(i_0_), .B(i_11_), .Y(new_new_n386_));
  AN2        g364(.A(i_1_), .B(i_6_), .Y(new_new_n387_));
  NOi21      g365(.An(i_2_), .B(i_12_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n388_), .B(new_new_n387_), .Y(new_new_n389_));
  INV        g367(.A(new_new_n389_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n136_), .B(i_9_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n391_), .B(i_4_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n390_), .B(new_new_n392_), .Y(new_new_n393_));
  NAi21      g371(.An(i_9_), .B(i_4_), .Y(new_new_n394_));
  OR2        g372(.A(i_13_), .B(i_10_), .Y(new_new_n395_));
  NO3        g373(.A(new_new_n395_), .B(new_new_n114_), .C(new_new_n394_), .Y(new_new_n396_));
  OR2        g374(.A(new_new_n211_), .B(new_new_n210_), .Y(new_new_n397_));
  NO2        g375(.A(new_new_n98_), .B(new_new_n25_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n268_), .B(new_new_n398_), .Y(new_new_n399_));
  NA2        g377(.A(i_5_), .B(new_new_n205_), .Y(new_new_n400_));
  OAI220     g378(.A0(new_new_n400_), .A1(new_new_n397_), .B0(new_new_n399_), .B1(new_new_n325_), .Y(new_new_n401_));
  INV        g379(.A(new_new_n401_), .Y(new_new_n402_));
  AOI210     g380(.A0(new_new_n402_), .A1(new_new_n393_), .B0(new_new_n26_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n307_), .B(new_new_n306_), .Y(new_new_n404_));
  AOI220     g382(.A0(new_new_n282_), .A1(new_new_n272_), .B0(new_new_n276_), .B1(new_new_n300_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n405_), .B(i_5_), .Y(new_new_n406_));
  AOI220     g384(.A0(i_3_), .A1(new_new_n281_), .B0(i_6_), .B1(new_new_n205_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n407_), .B(new_new_n270_), .Y(new_new_n408_));
  NO3        g386(.A(new_new_n408_), .B(new_new_n406_), .C(new_new_n404_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n189_), .B(new_new_n93_), .Y(new_new_n410_));
  NA3        g388(.A(new_new_n309_), .B(new_new_n157_), .C(new_new_n82_), .Y(new_new_n411_));
  AOI210     g389(.A0(new_new_n411_), .A1(new_new_n410_), .B0(i_8_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n186_), .B(i_10_), .Y(new_new_n413_));
  NA3        g391(.A(new_new_n244_), .B(new_new_n60_), .C(i_2_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n282_), .B(new_new_n224_), .Y(new_new_n415_));
  OAI220     g393(.A0(new_new_n415_), .A1(new_new_n176_), .B0(new_new_n414_), .B1(new_new_n413_), .Y(new_new_n416_));
  NO2        g394(.A(i_3_), .B(new_new_n48_), .Y(new_new_n417_));
  NA3        g395(.A(new_new_n318_), .B(new_new_n317_), .C(new_new_n417_), .Y(new_new_n418_));
  INV        g396(.A(new_new_n418_), .Y(new_new_n419_));
  NO3        g397(.A(new_new_n419_), .B(new_new_n416_), .C(new_new_n412_), .Y(new_new_n420_));
  AOI210     g398(.A0(new_new_n420_), .A1(new_new_n409_), .B0(new_new_n259_), .Y(new_new_n421_));
  NO4        g399(.A(new_new_n421_), .B(new_new_n403_), .C(new_new_n384_), .D(new_new_n363_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n69_), .B(i_13_), .Y(new_new_n423_));
  NO2        g401(.A(i_10_), .B(i_9_), .Y(new_new_n424_));
  NAi21      g402(.An(i_12_), .B(i_8_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n425_), .B(i_3_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n295_), .B(i_0_), .Y(new_new_n427_));
  NO3        g405(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n428_));
  NA2        g406(.A(new_new_n256_), .B(new_new_n94_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n429_), .B(new_new_n428_), .Y(new_new_n430_));
  NA2        g408(.A(i_8_), .B(i_9_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n268_), .B(new_new_n199_), .Y(new_new_n432_));
  OAI220     g410(.A0(new_new_n432_), .A1(new_new_n431_), .B0(new_new_n430_), .B1(new_new_n427_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n238_), .B(new_new_n294_), .Y(new_new_n434_));
  NO3        g412(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n435_));
  INV        g413(.A(new_new_n435_), .Y(new_new_n436_));
  NA3        g414(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n437_));
  NA4        g415(.A(new_new_n139_), .B(new_new_n112_), .C(new_new_n76_), .D(new_new_n23_), .Y(new_new_n438_));
  OAI220     g416(.A0(new_new_n438_), .A1(new_new_n437_), .B0(new_new_n436_), .B1(new_new_n434_), .Y(new_new_n439_));
  NO2        g417(.A(new_new_n439_), .B(new_new_n433_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n281_), .B(new_new_n105_), .Y(new_new_n441_));
  OR2        g419(.A(new_new_n441_), .B(new_new_n201_), .Y(new_new_n442_));
  BUFFER     g420(.A(new_new_n283_), .Y(new_new_n443_));
  OA220      g421(.A0(new_new_n443_), .A1(new_new_n156_), .B0(new_new_n442_), .B1(new_new_n221_), .Y(new_new_n444_));
  NA2        g422(.A(new_new_n93_), .B(i_13_), .Y(new_new_n445_));
  NO3        g423(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n446_));
  NO2        g424(.A(i_6_), .B(i_7_), .Y(new_new_n447_));
  NA2        g425(.A(new_new_n447_), .B(new_new_n446_), .Y(new_new_n448_));
  NO2        g426(.A(i_11_), .B(i_1_), .Y(new_new_n449_));
  OR2        g427(.A(i_11_), .B(i_8_), .Y(new_new_n450_));
  NOi21      g428(.An(i_2_), .B(i_7_), .Y(new_new_n451_));
  NAi31      g429(.An(new_new_n450_), .B(new_new_n451_), .C(i_0_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n395_), .B(i_6_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n453_), .B(i_1_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n454_), .B(new_new_n452_), .Y(new_new_n455_));
  NO2        g433(.A(i_3_), .B(new_new_n186_), .Y(new_new_n456_));
  NO2        g434(.A(i_6_), .B(i_10_), .Y(new_new_n457_));
  NA4        g435(.A(new_new_n457_), .B(new_new_n299_), .C(new_new_n456_), .D(new_new_n226_), .Y(new_new_n458_));
  NO2        g436(.A(new_new_n458_), .B(new_new_n149_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n151_), .B(i_3_), .Y(new_new_n461_));
  NAi31      g439(.An(new_new_n460_), .B(new_new_n461_), .C(new_new_n218_), .Y(new_new_n462_));
  INV        g440(.A(new_new_n462_), .Y(new_new_n463_));
  NO3        g441(.A(new_new_n463_), .B(new_new_n459_), .C(new_new_n455_), .Y(new_new_n464_));
  NA2        g442(.A(new_new_n428_), .B(new_new_n364_), .Y(new_new_n465_));
  NAi21      g443(.An(new_new_n211_), .B(new_new_n376_), .Y(new_new_n466_));
  NO2        g444(.A(new_new_n26_), .B(i_5_), .Y(new_new_n467_));
  NA3        g445(.A(i_6_), .B(new_new_n467_), .C(new_new_n136_), .Y(new_new_n468_));
  OR3        g446(.A(i_4_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n469_));
  NO2        g447(.A(new_new_n469_), .B(new_new_n468_), .Y(new_new_n470_));
  NA2        g448(.A(new_new_n27_), .B(i_10_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n299_), .B(new_new_n227_), .Y(new_new_n472_));
  OAI220     g450(.A0(new_new_n472_), .A1(new_new_n414_), .B0(new_new_n471_), .B1(new_new_n445_), .Y(new_new_n473_));
  NA4        g451(.A(new_new_n292_), .B(new_new_n216_), .C(new_new_n69_), .D(new_new_n226_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n474_), .B(new_new_n448_), .Y(new_new_n475_));
  NO3        g453(.A(new_new_n475_), .B(new_new_n473_), .C(new_new_n470_), .Y(new_new_n476_));
  NA4        g454(.A(new_new_n476_), .B(new_new_n464_), .C(new_new_n444_), .D(new_new_n440_), .Y(new_new_n477_));
  NA3        g455(.A(new_new_n292_), .B(new_new_n169_), .C(new_new_n167_), .Y(new_new_n478_));
  OAI210     g456(.A0(new_new_n287_), .A1(new_new_n174_), .B0(new_new_n478_), .Y(new_new_n479_));
  AN2        g457(.A(new_new_n272_), .B(new_new_n223_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n480_), .B(new_new_n479_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n299_), .B(new_new_n158_), .Y(new_new_n482_));
  OAI210     g460(.A0(new_new_n482_), .A1(new_new_n221_), .B0(new_new_n293_), .Y(new_new_n483_));
  NA2        g461(.A(new_new_n483_), .B(new_new_n308_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n364_), .B(new_new_n217_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n339_), .B(new_new_n69_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n356_), .B(new_new_n348_), .Y(new_new_n487_));
  OR2        g465(.A(new_new_n485_), .B(new_new_n487_), .Y(new_new_n488_));
  NO2        g466(.A(new_new_n36_), .B(i_8_), .Y(new_new_n489_));
  NAi41      g467(.An(new_new_n486_), .B(new_new_n457_), .C(new_new_n489_), .D(new_new_n47_), .Y(new_new_n490_));
  AOI210     g468(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n396_), .Y(new_new_n491_));
  NA3        g469(.A(new_new_n491_), .B(new_new_n490_), .C(new_new_n488_), .Y(new_new_n492_));
  INV        g470(.A(new_new_n492_), .Y(new_new_n493_));
  AOI210     g471(.A0(new_new_n187_), .A1(i_9_), .B0(new_new_n255_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n494_), .B(new_new_n192_), .Y(new_new_n495_));
  NO2        g473(.A(new_new_n176_), .B(new_new_n82_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n496_), .B(new_new_n495_), .Y(new_new_n497_));
  NA4        g475(.A(new_new_n497_), .B(new_new_n493_), .C(new_new_n484_), .D(new_new_n481_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n366_), .B(new_new_n281_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n163_), .B(new_new_n499_), .Y(new_new_n500_));
  NO2        g478(.A(i_12_), .B(new_new_n186_), .Y(new_new_n501_));
  NO3        g479(.A(i_10_), .B(new_new_n186_), .C(new_new_n441_), .Y(new_new_n502_));
  NOi31      g480(.An(new_new_n302_), .B(new_new_n395_), .C(new_new_n38_), .Y(new_new_n503_));
  OAI210     g481(.A0(new_new_n503_), .A1(new_new_n502_), .B0(new_new_n500_), .Y(new_new_n504_));
  NO2        g482(.A(i_8_), .B(i_7_), .Y(new_new_n505_));
  OAI210     g483(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n506_), .B(new_new_n216_), .Y(new_new_n507_));
  AOI220     g485(.A0(new_new_n309_), .A1(new_new_n40_), .B0(new_new_n224_), .B1(new_new_n200_), .Y(new_new_n508_));
  OAI220     g486(.A0(new_new_n508_), .A1(new_new_n176_), .B0(new_new_n507_), .B1(new_new_n230_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n45_), .B(i_10_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n510_), .B(i_6_), .Y(new_new_n511_));
  NA3        g489(.A(new_new_n511_), .B(new_new_n509_), .C(new_new_n505_), .Y(new_new_n512_));
  NO2        g490(.A(new_new_n445_), .B(new_new_n128_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n513_), .B(new_new_n255_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n287_), .B(new_new_n174_), .Y(new_new_n515_));
  NA2        g493(.A(new_new_n515_), .B(new_new_n435_), .Y(new_new_n516_));
  NA4        g494(.A(new_new_n516_), .B(new_new_n514_), .C(new_new_n512_), .D(new_new_n504_), .Y(new_new_n517_));
  NA3        g495(.A(new_new_n212_), .B(new_new_n67_), .C(new_new_n45_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n268_), .B(new_new_n80_), .Y(new_new_n519_));
  AOI210     g497(.A0(new_new_n518_), .A1(new_new_n329_), .B0(new_new_n519_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n282_), .B(new_new_n272_), .Y(new_new_n521_));
  NO2        g499(.A(new_new_n521_), .B(new_new_n166_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n424_), .B(new_new_n214_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n523_), .B(new_new_n524_), .Y(new_new_n525_));
  NA2        g503(.A(i_0_), .B(new_new_n48_), .Y(new_new_n526_));
  NA3        g504(.A(new_new_n501_), .B(new_new_n261_), .C(new_new_n526_), .Y(new_new_n527_));
  NO2        g505(.A(i_2_), .B(new_new_n527_), .Y(new_new_n528_));
  NO4        g506(.A(new_new_n528_), .B(new_new_n525_), .C(new_new_n522_), .D(new_new_n520_), .Y(new_new_n529_));
  NO4        g507(.A(new_new_n239_), .B(new_new_n43_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n530_));
  NO3        g508(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n222_), .B(new_new_n36_), .Y(new_new_n532_));
  AN2        g510(.A(new_new_n532_), .B(new_new_n531_), .Y(new_new_n533_));
  AN2        g511(.A(new_new_n530_), .B(new_new_n339_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n395_), .B(i_1_), .Y(new_new_n535_));
  NOi31      g513(.An(new_new_n535_), .B(new_new_n429_), .C(new_new_n69_), .Y(new_new_n536_));
  AN4        g514(.A(new_new_n536_), .B(new_new_n392_), .C(new_new_n467_), .D(i_2_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n405_), .B(new_new_n170_), .Y(new_new_n538_));
  NO3        g516(.A(new_new_n538_), .B(new_new_n537_), .C(new_new_n534_), .Y(new_new_n539_));
  NOi21      g517(.An(i_10_), .B(i_6_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n111_), .B(new_new_n23_), .Y(new_new_n541_));
  NA2        g519(.A(new_new_n302_), .B(new_new_n158_), .Y(new_new_n542_));
  AOI220     g520(.A0(new_new_n542_), .A1(new_new_n415_), .B0(new_new_n177_), .B1(new_new_n175_), .Y(new_new_n543_));
  NOi21      g521(.An(new_new_n140_), .B(new_new_n315_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n544_), .B(new_new_n543_), .Y(new_new_n545_));
  INV        g523(.A(new_new_n305_), .Y(new_new_n546_));
  NO2        g524(.A(i_12_), .B(new_new_n82_), .Y(new_new_n547_));
  NA2        g525(.A(new_new_n167_), .B(i_0_), .Y(new_new_n548_));
  NO3        g526(.A(new_new_n548_), .B(new_new_n323_), .C(new_new_n287_), .Y(new_new_n549_));
  OR2        g527(.A(i_2_), .B(i_5_), .Y(new_new_n550_));
  OR2        g528(.A(new_new_n550_), .B(new_new_n387_), .Y(new_new_n551_));
  AOI210     g529(.A0(new_new_n357_), .A1(new_new_n232_), .B0(new_new_n191_), .Y(new_new_n552_));
  AOI210     g530(.A0(new_new_n552_), .A1(new_new_n551_), .B0(new_new_n466_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n553_), .B(new_new_n549_), .Y(new_new_n554_));
  NA4        g532(.A(new_new_n554_), .B(new_new_n545_), .C(new_new_n539_), .D(new_new_n529_), .Y(new_new_n555_));
  NO4        g533(.A(new_new_n555_), .B(new_new_n517_), .C(new_new_n498_), .D(new_new_n477_), .Y(new_new_n556_));
  NA4        g534(.A(new_new_n556_), .B(new_new_n422_), .C(new_new_n338_), .D(new_new_n298_), .Y(mai7));
  NO2        g535(.A(new_new_n90_), .B(new_new_n52_), .Y(new_new_n558_));
  NA2        g536(.A(new_new_n457_), .B(new_new_n80_), .Y(new_new_n559_));
  NA2        g537(.A(i_11_), .B(new_new_n186_), .Y(new_new_n560_));
  NA3        g538(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n226_), .B(i_4_), .Y(new_new_n562_));
  NO2        g540(.A(new_new_n102_), .B(new_new_n561_), .Y(new_new_n563_));
  NA2        g541(.A(i_2_), .B(new_new_n82_), .Y(new_new_n564_));
  OAI210     g542(.A0(new_new_n85_), .A1(new_new_n196_), .B0(new_new_n197_), .Y(new_new_n565_));
  NO2        g543(.A(i_7_), .B(new_new_n37_), .Y(new_new_n566_));
  NA2        g544(.A(i_4_), .B(i_8_), .Y(new_new_n567_));
  AOI210     g545(.A0(new_new_n567_), .A1(new_new_n292_), .B0(new_new_n566_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n568_), .B(new_new_n564_), .Y(new_new_n569_));
  NO3        g547(.A(new_new_n569_), .B(new_new_n563_), .C(new_new_n558_), .Y(new_new_n570_));
  AOI210     g548(.A0(i_3_), .A1(new_new_n58_), .B0(i_10_), .Y(new_new_n571_));
  AOI210     g549(.A0(new_new_n571_), .A1(new_new_n226_), .B0(new_new_n155_), .Y(new_new_n572_));
  OR2        g550(.A(i_6_), .B(i_10_), .Y(new_new_n573_));
  NO2        g551(.A(new_new_n573_), .B(new_new_n23_), .Y(new_new_n574_));
  OR3        g552(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n575_));
  NO3        g553(.A(new_new_n575_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n576_));
  INV        g554(.A(new_new_n193_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n576_), .B(new_new_n574_), .Y(new_new_n578_));
  OA220      g556(.A0(new_new_n578_), .A1(new_new_n546_), .B0(new_new_n572_), .B1(new_new_n257_), .Y(new_new_n579_));
  AOI210     g557(.A0(new_new_n579_), .A1(new_new_n570_), .B0(new_new_n59_), .Y(new_new_n580_));
  NOi21      g558(.An(i_11_), .B(i_7_), .Y(new_new_n581_));
  AO210      g559(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n582_), .B(new_new_n581_), .Y(new_new_n583_));
  NA2        g561(.A(new_new_n84_), .B(new_new_n59_), .Y(new_new_n584_));
  AO210      g562(.A0(new_new_n584_), .A1(new_new_n361_), .B0(new_new_n41_), .Y(new_new_n585_));
  NA2        g563(.A(new_new_n218_), .B(new_new_n59_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n388_), .B(new_new_n31_), .Y(new_new_n587_));
  OR2        g565(.A(new_new_n202_), .B(new_new_n105_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n588_), .B(new_new_n587_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n59_), .B(i_9_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n590_), .B(i_4_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(new_new_n589_), .Y(new_new_n592_));
  NO2        g570(.A(i_1_), .B(i_12_), .Y(new_new_n593_));
  NA3        g571(.A(new_new_n593_), .B(new_new_n106_), .C(new_new_n24_), .Y(new_new_n594_));
  BUFFER     g572(.A(new_new_n594_), .Y(new_new_n595_));
  NA4        g573(.A(new_new_n595_), .B(new_new_n592_), .C(new_new_n586_), .D(new_new_n585_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n596_), .B(i_6_), .Y(new_new_n597_));
  NO2        g575(.A(i_6_), .B(i_11_), .Y(new_new_n598_));
  INV        g576(.A(new_new_n430_), .Y(new_new_n599_));
  NO4        g577(.A(new_new_n210_), .B(i_3_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n600_), .B(new_new_n590_), .Y(new_new_n601_));
  NA2        g579(.A(i_1_), .B(new_new_n247_), .Y(new_new_n602_));
  OAI210     g580(.A0(new_new_n602_), .A1(new_new_n45_), .B0(new_new_n601_), .Y(new_new_n603_));
  INV        g581(.A(i_2_), .Y(new_new_n604_));
  NA2        g582(.A(new_new_n132_), .B(i_9_), .Y(new_new_n605_));
  NA3        g583(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n606_));
  NO2        g584(.A(new_new_n47_), .B(i_1_), .Y(new_new_n607_));
  NA3        g585(.A(new_new_n607_), .B(new_new_n256_), .C(new_new_n45_), .Y(new_new_n608_));
  OAI220     g586(.A0(new_new_n608_), .A1(new_new_n606_), .B0(new_new_n605_), .B1(new_new_n604_), .Y(new_new_n609_));
  NO2        g587(.A(i_11_), .B(new_new_n37_), .Y(new_new_n610_));
  NA2        g588(.A(new_new_n610_), .B(new_new_n24_), .Y(new_new_n611_));
  NO3        g589(.A(new_new_n609_), .B(new_new_n603_), .C(new_new_n599_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n226_), .B(new_new_n98_), .Y(new_new_n613_));
  NO2        g591(.A(new_new_n613_), .B(new_new_n581_), .Y(new_new_n614_));
  NA2        g592(.A(new_new_n614_), .B(i_1_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n615_), .B(new_new_n575_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n616_), .B(new_new_n47_), .Y(new_new_n617_));
  NA2        g595(.A(i_3_), .B(new_new_n186_), .Y(new_new_n618_));
  NO2        g596(.A(new_new_n618_), .B(new_new_n111_), .Y(new_new_n619_));
  AN2        g597(.A(new_new_n619_), .B(new_new_n511_), .Y(new_new_n620_));
  NO2        g598(.A(new_new_n222_), .B(new_new_n45_), .Y(new_new_n621_));
  NO3        g599(.A(new_new_n621_), .B(new_new_n295_), .C(i_12_), .Y(new_new_n622_));
  NO2        g600(.A(new_new_n114_), .B(new_new_n37_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n623_), .B(i_6_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n82_), .B(i_9_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n59_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n626_), .B(new_new_n593_), .Y(new_new_n627_));
  NO4        g605(.A(new_new_n627_), .B(new_new_n624_), .C(new_new_n622_), .D(i_4_), .Y(new_new_n628_));
  NA2        g606(.A(i_1_), .B(i_3_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n431_), .B(new_new_n90_), .Y(new_new_n630_));
  AOI210     g608(.A0(new_new_n621_), .A1(new_new_n540_), .B0(new_new_n630_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n631_), .B(new_new_n629_), .Y(new_new_n632_));
  NO3        g610(.A(new_new_n632_), .B(new_new_n628_), .C(new_new_n620_), .Y(new_new_n633_));
  NA4        g611(.A(new_new_n633_), .B(new_new_n617_), .C(new_new_n612_), .D(new_new_n597_), .Y(new_new_n634_));
  NO3        g612(.A(new_new_n450_), .B(i_3_), .C(i_7_), .Y(new_new_n635_));
  NOi21      g613(.An(new_new_n635_), .B(i_10_), .Y(new_new_n636_));
  OA210      g614(.A0(new_new_n636_), .A1(new_new_n233_), .B0(new_new_n82_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n356_), .B(new_new_n355_), .Y(new_new_n638_));
  NA3        g616(.A(new_new_n457_), .B(new_new_n489_), .C(new_new_n47_), .Y(new_new_n639_));
  NO3        g617(.A(new_new_n451_), .B(new_new_n567_), .C(new_new_n82_), .Y(new_new_n640_));
  NA2        g618(.A(new_new_n640_), .B(new_new_n25_), .Y(new_new_n641_));
  NA3        g619(.A(new_new_n155_), .B(new_new_n80_), .C(new_new_n82_), .Y(new_new_n642_));
  NA3        g620(.A(new_new_n642_), .B(new_new_n641_), .C(new_new_n639_), .Y(new_new_n643_));
  OAI210     g621(.A0(new_new_n643_), .A1(new_new_n637_), .B0(i_1_), .Y(new_new_n644_));
  AOI210     g622(.A0(new_new_n256_), .A1(new_new_n94_), .B0(i_1_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n354_), .B(i_2_), .Y(new_new_n646_));
  NA2        g624(.A(new_new_n646_), .B(new_new_n645_), .Y(new_new_n647_));
  AOI210     g625(.A0(new_new_n647_), .A1(new_new_n644_), .B0(i_13_), .Y(new_new_n648_));
  OR2        g626(.A(i_11_), .B(i_7_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n52_), .B(i_12_), .Y(new_new_n650_));
  INV        g628(.A(new_new_n650_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n233_), .B(new_new_n126_), .Y(new_new_n652_));
  OAI220     g630(.A0(new_new_n652_), .A1(new_new_n41_), .B0(new_new_n651_), .B1(new_new_n90_), .Y(new_new_n653_));
  INV        g631(.A(new_new_n653_), .Y(new_new_n654_));
  NA2        g632(.A(new_new_n365_), .B(new_new_n607_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n655_), .B(new_new_n230_), .Y(new_new_n656_));
  AOI210     g634(.A0(new_new_n425_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n657_));
  NOi31      g635(.An(new_new_n657_), .B(new_new_n559_), .C(new_new_n45_), .Y(new_new_n658_));
  NA2        g636(.A(new_new_n124_), .B(i_13_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n606_), .B(new_new_n111_), .Y(new_new_n660_));
  INV        g638(.A(new_new_n660_), .Y(new_new_n661_));
  OAI220     g639(.A0(new_new_n661_), .A1(new_new_n67_), .B0(new_new_n659_), .B1(new_new_n645_), .Y(new_new_n662_));
  NA2        g640(.A(new_new_n26_), .B(new_new_n186_), .Y(new_new_n663_));
  NA2        g641(.A(new_new_n663_), .B(i_7_), .Y(new_new_n664_));
  NO3        g642(.A(new_new_n451_), .B(new_new_n226_), .C(new_new_n82_), .Y(new_new_n665_));
  NA2        g643(.A(new_new_n665_), .B(new_new_n664_), .Y(new_new_n666_));
  NO2        g644(.A(new_new_n666_), .B(new_new_n577_), .Y(new_new_n667_));
  NO4        g645(.A(new_new_n667_), .B(new_new_n662_), .C(new_new_n658_), .D(new_new_n656_), .Y(new_new_n668_));
  OR2        g646(.A(i_11_), .B(i_6_), .Y(new_new_n669_));
  NA2        g647(.A(new_new_n562_), .B(i_7_), .Y(new_new_n670_));
  AOI210     g648(.A0(new_new_n670_), .A1(new_new_n661_), .B0(new_new_n669_), .Y(new_new_n671_));
  NA3        g649(.A(new_new_n388_), .B(new_new_n566_), .C(new_new_n94_), .Y(new_new_n672_));
  NA2        g650(.A(new_new_n598_), .B(i_13_), .Y(new_new_n673_));
  NA2        g651(.A(new_new_n99_), .B(new_new_n663_), .Y(new_new_n674_));
  NAi21      g652(.An(i_11_), .B(i_12_), .Y(new_new_n675_));
  NOi41      g653(.An(new_new_n107_), .B(new_new_n675_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n676_));
  NO3        g654(.A(new_new_n451_), .B(new_new_n547_), .C(new_new_n567_), .Y(new_new_n677_));
  AOI220     g655(.A0(new_new_n677_), .A1(new_new_n299_), .B0(new_new_n676_), .B1(new_new_n674_), .Y(new_new_n678_));
  NA3        g656(.A(new_new_n678_), .B(new_new_n673_), .C(new_new_n672_), .Y(new_new_n679_));
  OAI210     g657(.A0(new_new_n679_), .A1(new_new_n671_), .B0(new_new_n59_), .Y(new_new_n680_));
  NO3        g658(.A(i_9_), .B(i_3_), .C(new_new_n562_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n681_), .B(new_new_n353_), .Y(new_new_n682_));
  NO2        g660(.A(i_3_), .B(i_2_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n683_), .B(new_new_n593_), .Y(new_new_n684_));
  NA2        g662(.A(new_new_n684_), .B(new_new_n682_), .Y(new_new_n685_));
  NA3        g663(.A(new_new_n685_), .B(new_new_n46_), .C(new_new_n217_), .Y(new_new_n686_));
  NA4        g664(.A(new_new_n686_), .B(new_new_n680_), .C(new_new_n668_), .D(new_new_n654_), .Y(new_new_n687_));
  OR4        g665(.A(new_new_n687_), .B(new_new_n648_), .C(new_new_n634_), .D(new_new_n580_), .Y(mai5));
  NA2        g666(.A(new_new_n614_), .B(new_new_n258_), .Y(new_new_n689_));
  INV        g667(.A(new_new_n689_), .Y(new_new_n690_));
  NO3        g668(.A(i_11_), .B(new_new_n226_), .C(i_13_), .Y(new_new_n691_));
  NO2        g669(.A(new_new_n121_), .B(new_new_n23_), .Y(new_new_n692_));
  INV        g670(.A(new_new_n424_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n305_), .B(new_new_n541_), .Y(new_new_n694_));
  INV        g672(.A(new_new_n694_), .Y(new_new_n695_));
  NO2        g673(.A(new_new_n695_), .B(new_new_n690_), .Y(new_new_n696_));
  INV        g674(.A(new_new_n165_), .Y(new_new_n697_));
  INV        g675(.A(new_new_n233_), .Y(new_new_n698_));
  OAI210     g676(.A0(new_new_n646_), .A1(new_new_n426_), .B0(new_new_n107_), .Y(new_new_n699_));
  AOI210     g677(.A0(new_new_n699_), .A1(new_new_n698_), .B0(new_new_n697_), .Y(new_new_n700_));
  NO2        g678(.A(new_new_n431_), .B(new_new_n26_), .Y(new_new_n701_));
  NO2        g679(.A(new_new_n701_), .B(new_new_n398_), .Y(new_new_n702_));
  NA2        g680(.A(new_new_n702_), .B(i_2_), .Y(new_new_n703_));
  INV        g681(.A(new_new_n703_), .Y(new_new_n704_));
  AOI210     g682(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n395_), .Y(new_new_n705_));
  AOI210     g683(.A0(new_new_n705_), .A1(new_new_n704_), .B0(new_new_n700_), .Y(new_new_n706_));
  NO2        g684(.A(new_new_n183_), .B(new_new_n122_), .Y(new_new_n707_));
  OAI210     g685(.A0(new_new_n707_), .A1(new_new_n692_), .B0(i_2_), .Y(new_new_n708_));
  INV        g686(.A(new_new_n166_), .Y(new_new_n709_));
  NO3        g687(.A(new_new_n582_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n710_));
  AOI210     g688(.A0(new_new_n709_), .A1(new_new_n85_), .B0(new_new_n710_), .Y(new_new_n711_));
  AOI210     g689(.A0(new_new_n711_), .A1(new_new_n708_), .B0(new_new_n186_), .Y(new_new_n712_));
  OA210      g690(.A0(new_new_n583_), .A1(new_new_n123_), .B0(i_13_), .Y(new_new_n713_));
  NA2        g691(.A(new_new_n193_), .B(new_new_n196_), .Y(new_new_n714_));
  INV        g692(.A(new_new_n145_), .Y(new_new_n715_));
  AOI210     g693(.A0(new_new_n715_), .A1(new_new_n714_), .B0(new_new_n357_), .Y(new_new_n716_));
  AOI210     g694(.A0(new_new_n202_), .A1(new_new_n142_), .B0(new_new_n489_), .Y(new_new_n717_));
  NA2        g695(.A(new_new_n717_), .B(new_new_n398_), .Y(new_new_n718_));
  NO2        g696(.A(new_new_n99_), .B(new_new_n45_), .Y(new_new_n719_));
  INV        g697(.A(new_new_n288_), .Y(new_new_n720_));
  NA4        g698(.A(new_new_n720_), .B(new_new_n292_), .C(new_new_n121_), .D(new_new_n43_), .Y(new_new_n721_));
  OAI210     g699(.A0(new_new_n721_), .A1(new_new_n719_), .B0(new_new_n718_), .Y(new_new_n722_));
  NO4        g700(.A(new_new_n722_), .B(new_new_n716_), .C(new_new_n713_), .D(new_new_n712_), .Y(new_new_n723_));
  NA2        g701(.A(new_new_n541_), .B(new_new_n28_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n691_), .B(new_new_n262_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n725_), .B(new_new_n724_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n58_), .B(i_12_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n727_), .B(new_new_n123_), .Y(new_new_n728_));
  NO2        g706(.A(new_new_n728_), .B(new_new_n560_), .Y(new_new_n729_));
  AOI220     g707(.A0(new_new_n729_), .A1(new_new_n36_), .B0(new_new_n726_), .B1(new_new_n47_), .Y(new_new_n730_));
  NA4        g708(.A(new_new_n730_), .B(new_new_n723_), .C(new_new_n706_), .D(new_new_n696_), .Y(mai6));
  NO3        g709(.A(i_9_), .B(new_new_n294_), .C(i_1_), .Y(new_new_n732_));
  NO2        g710(.A(new_new_n179_), .B(new_new_n133_), .Y(new_new_n733_));
  OAI210     g711(.A0(new_new_n733_), .A1(new_new_n732_), .B0(new_new_n683_), .Y(new_new_n734_));
  NA4        g712(.A(new_new_n367_), .B(new_new_n456_), .C(new_new_n67_), .D(new_new_n98_), .Y(new_new_n735_));
  INV        g713(.A(new_new_n735_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n213_), .B(new_new_n460_), .Y(new_new_n737_));
  NO2        g715(.A(i_11_), .B(i_9_), .Y(new_new_n738_));
  NO2        g716(.A(new_new_n736_), .B(new_new_n314_), .Y(new_new_n739_));
  AO210      g717(.A0(new_new_n739_), .A1(new_new_n734_), .B0(i_12_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n358_), .B(new_new_n318_), .Y(new_new_n741_));
  NA2        g719(.A(new_new_n547_), .B(new_new_n59_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n636_), .B(new_new_n67_), .Y(new_new_n743_));
  BUFFER     g721(.A(new_new_n584_), .Y(new_new_n744_));
  NA4        g722(.A(new_new_n744_), .B(new_new_n743_), .C(new_new_n742_), .D(new_new_n741_), .Y(new_new_n745_));
  INV        g723(.A(new_new_n190_), .Y(new_new_n746_));
  AOI220     g724(.A0(new_new_n746_), .A1(new_new_n738_), .B0(new_new_n745_), .B1(new_new_n69_), .Y(new_new_n747_));
  INV        g725(.A(new_new_n313_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n71_), .B(new_new_n126_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n749_), .B(new_new_n748_), .Y(new_new_n750_));
  NO2        g728(.A(new_new_n239_), .B(i_9_), .Y(new_new_n751_));
  NA2        g729(.A(new_new_n751_), .B(new_new_n727_), .Y(new_new_n752_));
  AOI210     g730(.A0(new_new_n752_), .A1(new_new_n487_), .B0(new_new_n179_), .Y(new_new_n753_));
  NAi32      g731(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n669_), .B(new_new_n754_), .Y(new_new_n755_));
  OAI210     g733(.A0(new_new_n635_), .A1(new_new_n532_), .B0(new_new_n531_), .Y(new_new_n756_));
  NAi21      g734(.An(new_new_n755_), .B(new_new_n756_), .Y(new_new_n757_));
  OR3        g735(.A(new_new_n757_), .B(new_new_n753_), .C(new_new_n750_), .Y(new_new_n758_));
  NO2        g736(.A(new_new_n649_), .B(i_2_), .Y(new_new_n759_));
  NA2        g737(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n760_));
  NO2        g738(.A(new_new_n760_), .B(new_new_n387_), .Y(new_new_n761_));
  NA2        g739(.A(new_new_n761_), .B(new_new_n759_), .Y(new_new_n762_));
  AO220      g740(.A0(new_new_n342_), .A1(new_new_n333_), .B0(new_new_n373_), .B1(new_new_n560_), .Y(new_new_n763_));
  NA3        g741(.A(new_new_n763_), .B(new_new_n243_), .C(i_7_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n426_), .B(new_new_n141_), .Y(new_new_n765_));
  OR2        g743(.A(new_new_n693_), .B(new_new_n36_), .Y(new_new_n766_));
  NA4        g744(.A(new_new_n766_), .B(new_new_n765_), .C(new_new_n764_), .D(new_new_n762_), .Y(new_new_n767_));
  OAI210     g745(.A0(i_6_), .A1(i_11_), .B0(new_new_n83_), .Y(new_new_n768_));
  AOI220     g746(.A0(new_new_n768_), .A1(new_new_n531_), .B0(new_new_n737_), .B1(new_new_n664_), .Y(new_new_n769_));
  NA2        g747(.A(new_new_n373_), .B(new_new_n66_), .Y(new_new_n770_));
  NA3        g748(.A(new_new_n770_), .B(new_new_n769_), .C(new_new_n565_), .Y(new_new_n771_));
  AO210      g749(.A0(new_new_n489_), .A1(new_new_n47_), .B0(new_new_n84_), .Y(new_new_n772_));
  NA3        g750(.A(new_new_n772_), .B(new_new_n457_), .C(new_new_n212_), .Y(new_new_n773_));
  AOI210     g751(.A0(new_new_n426_), .A1(new_new_n424_), .B0(new_new_n530_), .Y(new_new_n774_));
  NA2        g752(.A(new_new_n108_), .B(new_new_n386_), .Y(new_new_n775_));
  INV        g753(.A(new_new_n551_), .Y(new_new_n776_));
  NA3        g754(.A(new_new_n776_), .B(new_new_n313_), .C(i_7_), .Y(new_new_n777_));
  NA4        g755(.A(new_new_n777_), .B(new_new_n775_), .C(new_new_n774_), .D(new_new_n773_), .Y(new_new_n778_));
  NO4        g756(.A(new_new_n778_), .B(new_new_n771_), .C(new_new_n767_), .D(new_new_n758_), .Y(new_new_n779_));
  NA4        g757(.A(new_new_n779_), .B(new_new_n747_), .C(new_new_n740_), .D(new_new_n362_), .Y(mai3));
  NA2        g758(.A(i_12_), .B(i_10_), .Y(new_new_n781_));
  NA2        g759(.A(i_6_), .B(i_7_), .Y(new_new_n782_));
  NO2        g760(.A(new_new_n782_), .B(i_0_), .Y(new_new_n783_));
  NO2        g761(.A(i_11_), .B(new_new_n226_), .Y(new_new_n784_));
  NA2        g762(.A(new_new_n276_), .B(new_new_n784_), .Y(new_new_n785_));
  NO2        g763(.A(new_new_n785_), .B(new_new_n186_), .Y(new_new_n786_));
  NO3        g764(.A(new_new_n427_), .B(new_new_n87_), .C(new_new_n45_), .Y(new_new_n787_));
  OA210      g765(.A0(new_new_n787_), .A1(new_new_n786_), .B0(new_new_n167_), .Y(new_new_n788_));
  NO2        g766(.A(new_new_n588_), .B(new_new_n431_), .Y(new_new_n789_));
  NA2        g767(.A(new_new_n388_), .B(new_new_n46_), .Y(new_new_n790_));
  NO2        g768(.A(new_new_n962_), .B(new_new_n48_), .Y(new_new_n791_));
  NA2        g769(.A(new_new_n657_), .B(new_new_n625_), .Y(new_new_n792_));
  NA2        g770(.A(i_0_), .B(new_new_n417_), .Y(new_new_n793_));
  NO2        g771(.A(new_new_n793_), .B(new_new_n792_), .Y(new_new_n794_));
  NOi21      g772(.An(i_5_), .B(i_9_), .Y(new_new_n795_));
  NA2        g773(.A(new_new_n795_), .B(new_new_n423_), .Y(new_new_n796_));
  BUFFER     g774(.A(new_new_n256_), .Y(new_new_n797_));
  AOI210     g775(.A0(new_new_n797_), .A1(new_new_n449_), .B0(new_new_n640_), .Y(new_new_n798_));
  NO3        g776(.A(new_new_n391_), .B(new_new_n256_), .C(new_new_n69_), .Y(new_new_n799_));
  NO2        g777(.A(new_new_n168_), .B(new_new_n142_), .Y(new_new_n800_));
  AOI210     g778(.A0(new_new_n800_), .A1(new_new_n232_), .B0(new_new_n799_), .Y(new_new_n801_));
  OAI220     g779(.A0(new_new_n801_), .A1(new_new_n174_), .B0(new_new_n798_), .B1(new_new_n796_), .Y(new_new_n802_));
  NO4        g780(.A(new_new_n802_), .B(new_new_n794_), .C(new_new_n791_), .D(new_new_n788_), .Y(new_new_n803_));
  NA2        g781(.A(new_new_n179_), .B(new_new_n24_), .Y(new_new_n804_));
  NAi21      g782(.An(new_new_n156_), .B(new_new_n417_), .Y(new_new_n805_));
  NO2        g783(.A(new_new_n805_), .B(i_2_), .Y(new_new_n806_));
  INV        g784(.A(new_new_n806_), .Y(new_new_n807_));
  INV        g785(.A(new_new_n280_), .Y(new_new_n808_));
  NA2        g786(.A(new_new_n808_), .B(new_new_n660_), .Y(new_new_n809_));
  NO4        g787(.A(new_new_n550_), .B(new_new_n210_), .C(new_new_n395_), .D(new_new_n387_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n810_), .B(i_11_), .Y(new_new_n811_));
  AN2        g789(.A(new_new_n93_), .B(new_new_n231_), .Y(new_new_n812_));
  NA2        g790(.A(new_new_n691_), .B(new_new_n314_), .Y(new_new_n813_));
  INV        g791(.A(new_new_n54_), .Y(new_new_n814_));
  OAI220     g792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n611_), .B1(new_new_n507_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n241_), .B(new_new_n147_), .Y(new_new_n816_));
  INV        g794(.A(new_new_n510_), .Y(new_new_n817_));
  NO4        g795(.A(new_new_n111_), .B(new_new_n54_), .C(new_new_n618_), .D(i_5_), .Y(new_new_n818_));
  AO220      g796(.A0(new_new_n818_), .A1(new_new_n817_), .B0(new_new_n816_), .B1(i_6_), .Y(new_new_n819_));
  NA2        g797(.A(new_new_n179_), .B(new_new_n80_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n535_), .B(i_4_), .Y(new_new_n821_));
  NA2        g799(.A(new_new_n182_), .B(new_new_n196_), .Y(new_new_n822_));
  OAI220     g800(.A0(new_new_n822_), .A1(new_new_n813_), .B0(new_new_n821_), .B1(new_new_n820_), .Y(new_new_n823_));
  NO4        g801(.A(new_new_n823_), .B(new_new_n819_), .C(new_new_n815_), .D(new_new_n812_), .Y(new_new_n824_));
  NA4        g802(.A(new_new_n824_), .B(new_new_n811_), .C(new_new_n809_), .D(new_new_n807_), .Y(new_new_n825_));
  NA2        g803(.A(i_11_), .B(i_9_), .Y(new_new_n826_));
  NO2        g804(.A(new_new_n48_), .B(i_7_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n372_), .B(new_new_n172_), .Y(new_new_n828_));
  NA2        g806(.A(new_new_n828_), .B(new_new_n154_), .Y(new_new_n829_));
  NO2        g807(.A(new_new_n826_), .B(new_new_n69_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n447_), .B(new_new_n220_), .Y(new_new_n831_));
  AOI210     g809(.A0(new_new_n356_), .A1(new_new_n42_), .B0(new_new_n385_), .Y(new_new_n832_));
  OAI220     g810(.A0(new_new_n832_), .A1(new_new_n796_), .B0(new_new_n831_), .B1(new_new_n168_), .Y(new_new_n833_));
  NO2        g811(.A(new_new_n833_), .B(new_new_n829_), .Y(new_new_n834_));
  NA2        g812(.A(new_new_n610_), .B(new_new_n118_), .Y(new_new_n835_));
  NO2        g813(.A(i_6_), .B(new_new_n835_), .Y(new_new_n836_));
  AOI210     g814(.A0(new_new_n425_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n837_));
  NA2        g815(.A(new_new_n165_), .B(new_new_n100_), .Y(new_new_n838_));
  NOi32      g816(.An(new_new_n837_), .Bn(new_new_n182_), .C(new_new_n838_), .Y(new_new_n839_));
  NA2        g817(.A(new_new_n566_), .B(new_new_n314_), .Y(new_new_n840_));
  NO2        g818(.A(new_new_n840_), .B(new_new_n790_), .Y(new_new_n841_));
  NO3        g819(.A(new_new_n841_), .B(new_new_n839_), .C(new_new_n836_), .Y(new_new_n842_));
  INV        g820(.A(i_5_), .Y(new_new_n843_));
  OR2        g821(.A(new_new_n838_), .B(new_new_n487_), .Y(new_new_n844_));
  NO3        g822(.A(new_new_n381_), .B(new_new_n345_), .C(new_new_n341_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n250_), .B(i_5_), .Y(new_new_n846_));
  NO2        g824(.A(new_new_n675_), .B(new_new_n245_), .Y(new_new_n847_));
  AOI210     g825(.A0(new_new_n847_), .A1(new_new_n846_), .B0(new_new_n845_), .Y(new_new_n848_));
  NA4        g826(.A(new_new_n848_), .B(new_new_n844_), .C(new_new_n842_), .D(new_new_n834_), .Y(new_new_n849_));
  NO2        g827(.A(new_new_n804_), .B(new_new_n228_), .Y(new_new_n850_));
  AN2        g828(.A(new_new_n316_), .B(new_new_n314_), .Y(new_new_n851_));
  AN2        g829(.A(new_new_n851_), .B(new_new_n800_), .Y(new_new_n852_));
  OAI210     g830(.A0(new_new_n852_), .A1(new_new_n850_), .B0(i_10_), .Y(new_new_n853_));
  INV        g831(.A(new_new_n781_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n854_), .B(new_new_n830_), .Y(new_new_n855_));
  NA3        g833(.A(new_new_n446_), .B(new_new_n388_), .C(new_new_n46_), .Y(new_new_n856_));
  OAI210     g834(.A0(new_new_n805_), .A1(i_7_), .B0(new_new_n856_), .Y(new_new_n857_));
  NA2        g835(.A(new_new_n830_), .B(new_new_n292_), .Y(new_new_n858_));
  OAI210     g836(.A0(i_2_), .A1(new_new_n181_), .B0(new_new_n858_), .Y(new_new_n859_));
  AOI220     g837(.A0(new_new_n859_), .A1(new_new_n447_), .B0(new_new_n857_), .B1(new_new_n69_), .Y(new_new_n860_));
  NAi21      g838(.An(i_9_), .B(i_5_), .Y(new_new_n861_));
  NO2        g839(.A(new_new_n861_), .B(new_new_n381_), .Y(new_new_n862_));
  NO2        g840(.A(new_new_n561_), .B(new_new_n102_), .Y(new_new_n863_));
  AOI220     g841(.A0(new_new_n863_), .A1(i_0_), .B0(new_new_n862_), .B1(new_new_n583_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n864_), .B(new_new_n82_), .Y(new_new_n865_));
  NO2        g843(.A(new_new_n865_), .B(new_new_n492_), .Y(new_new_n866_));
  NA4        g844(.A(new_new_n866_), .B(new_new_n860_), .C(new_new_n855_), .D(new_new_n853_), .Y(new_new_n867_));
  NO3        g845(.A(new_new_n867_), .B(new_new_n849_), .C(new_new_n825_), .Y(new_new_n868_));
  NO2        g846(.A(i_0_), .B(new_new_n675_), .Y(new_new_n869_));
  NA2        g847(.A(new_new_n69_), .B(new_new_n45_), .Y(new_new_n870_));
  NO3        g848(.A(new_new_n102_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n871_));
  AO220      g849(.A0(new_new_n871_), .A1(new_new_n45_), .B0(new_new_n869_), .B1(new_new_n167_), .Y(new_new_n872_));
  AOI210     g850(.A0(new_new_n742_), .A1(new_new_n638_), .B0(new_new_n838_), .Y(new_new_n873_));
  AOI210     g851(.A0(new_new_n872_), .A1(new_new_n330_), .B0(new_new_n873_), .Y(new_new_n874_));
  NA3        g852(.A(new_new_n140_), .B(new_new_n625_), .C(new_new_n69_), .Y(new_new_n875_));
  NO2        g853(.A(new_new_n756_), .B(new_new_n381_), .Y(new_new_n876_));
  NA3        g854(.A(new_new_n783_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n877_));
  NA2        g855(.A(new_new_n784_), .B(i_9_), .Y(new_new_n878_));
  AOI210     g856(.A0(new_new_n877_), .A1(new_new_n468_), .B0(new_new_n878_), .Y(new_new_n879_));
  NA2        g857(.A(new_new_n232_), .B(new_new_n219_), .Y(new_new_n880_));
  NO2        g858(.A(new_new_n880_), .B(new_new_n147_), .Y(new_new_n881_));
  NO3        g859(.A(new_new_n881_), .B(new_new_n879_), .C(new_new_n876_), .Y(new_new_n882_));
  NA3        g860(.A(new_new_n882_), .B(new_new_n875_), .C(new_new_n874_), .Y(new_new_n883_));
  NA2        g861(.A(new_new_n851_), .B(new_new_n357_), .Y(new_new_n884_));
  AOI210     g862(.A0(new_new_n287_), .A1(new_new_n156_), .B0(new_new_n884_), .Y(new_new_n885_));
  NA3        g863(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n886_));
  NA2        g864(.A(new_new_n827_), .B(new_new_n461_), .Y(new_new_n887_));
  AOI210     g865(.A0(new_new_n886_), .A1(new_new_n156_), .B0(new_new_n887_), .Y(new_new_n888_));
  NO2        g866(.A(new_new_n888_), .B(new_new_n885_), .Y(new_new_n889_));
  NA2        g867(.A(new_new_n536_), .B(new_new_n71_), .Y(new_new_n890_));
  NO3        g868(.A(new_new_n204_), .B(new_new_n364_), .C(i_0_), .Y(new_new_n891_));
  OAI210     g869(.A0(new_new_n891_), .A1(new_new_n72_), .B0(i_13_), .Y(new_new_n892_));
  INV        g870(.A(new_new_n212_), .Y(new_new_n893_));
  NO2        g871(.A(i_12_), .B(new_new_n577_), .Y(new_new_n894_));
  NA3        g872(.A(new_new_n894_), .B(new_new_n374_), .C(new_new_n893_), .Y(new_new_n895_));
  NA4        g873(.A(new_new_n895_), .B(new_new_n892_), .C(new_new_n890_), .D(new_new_n889_), .Y(new_new_n896_));
  NA2        g874(.A(new_new_n843_), .B(new_new_n461_), .Y(new_new_n897_));
  NA2        g875(.A(new_new_n333_), .B(new_new_n169_), .Y(new_new_n898_));
  OR2        g876(.A(new_new_n898_), .B(new_new_n897_), .Y(new_new_n899_));
  NA3        g877(.A(new_new_n574_), .B(new_new_n179_), .C(new_new_n80_), .Y(new_new_n900_));
  INV        g878(.A(new_new_n900_), .Y(new_new_n901_));
  NO3        g879(.A(new_new_n790_), .B(new_new_n52_), .C(new_new_n48_), .Y(new_new_n902_));
  INV        g880(.A(new_new_n465_), .Y(new_new_n903_));
  NO3        g881(.A(new_new_n903_), .B(new_new_n902_), .C(new_new_n901_), .Y(new_new_n904_));
  NA3        g882(.A(new_new_n367_), .B(new_new_n165_), .C(new_new_n164_), .Y(new_new_n905_));
  NA3        g883(.A(new_new_n827_), .B(new_new_n276_), .C(new_new_n219_), .Y(new_new_n906_));
  NA2        g884(.A(new_new_n906_), .B(new_new_n905_), .Y(new_new_n907_));
  NA3        g885(.A(new_new_n367_), .B(new_new_n317_), .C(new_new_n214_), .Y(new_new_n908_));
  INV        g886(.A(new_new_n908_), .Y(new_new_n909_));
  NOi31      g887(.An(new_new_n366_), .B(new_new_n870_), .C(new_new_n228_), .Y(new_new_n910_));
  NO3        g888(.A(new_new_n826_), .B(new_new_n212_), .C(new_new_n183_), .Y(new_new_n911_));
  NO4        g889(.A(new_new_n911_), .B(new_new_n910_), .C(new_new_n909_), .D(new_new_n907_), .Y(new_new_n912_));
  NA3        g890(.A(new_new_n912_), .B(new_new_n904_), .C(new_new_n899_), .Y(new_new_n913_));
  INV        g891(.A(new_new_n576_), .Y(new_new_n914_));
  NO3        g892(.A(new_new_n914_), .B(new_new_n526_), .C(i_7_), .Y(new_new_n915_));
  INV        g893(.A(new_new_n915_), .Y(new_new_n916_));
  NA2        g894(.A(new_new_n736_), .B(new_new_n169_), .Y(new_new_n917_));
  NA3        g895(.A(new_new_n95_), .B(new_new_n540_), .C(i_11_), .Y(new_new_n918_));
  NO2        g896(.A(new_new_n918_), .B(new_new_n149_), .Y(new_new_n919_));
  INV        g897(.A(new_new_n919_), .Y(new_new_n920_));
  NA3        g898(.A(new_new_n920_), .B(new_new_n917_), .C(new_new_n916_), .Y(new_new_n921_));
  NO4        g899(.A(new_new_n921_), .B(new_new_n913_), .C(new_new_n896_), .D(new_new_n883_), .Y(new_new_n922_));
  NA2        g900(.A(new_new_n759_), .B(new_new_n37_), .Y(new_new_n923_));
  NA3        g901(.A(new_new_n837_), .B(new_new_n353_), .C(i_5_), .Y(new_new_n924_));
  NA3        g902(.A(new_new_n924_), .B(new_new_n923_), .C(new_new_n572_), .Y(new_new_n925_));
  NA2        g903(.A(new_new_n925_), .B(new_new_n200_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n180_), .B(new_new_n182_), .Y(new_new_n927_));
  OAI210     g905(.A0(new_new_n576_), .A1(new_new_n574_), .B0(new_new_n305_), .Y(new_new_n928_));
  NAi31      g906(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n929_));
  NO2        g907(.A(new_new_n66_), .B(new_new_n929_), .Y(new_new_n930_));
  INV        g908(.A(new_new_n930_), .Y(new_new_n931_));
  NA3        g909(.A(new_new_n931_), .B(new_new_n928_), .C(new_new_n927_), .Y(new_new_n932_));
  NO2        g910(.A(new_new_n437_), .B(new_new_n256_), .Y(new_new_n933_));
  NO4        g911(.A(new_new_n222_), .B(new_new_n139_), .C(new_new_n629_), .D(new_new_n37_), .Y(new_new_n934_));
  NO3        g912(.A(new_new_n934_), .B(new_new_n933_), .C(new_new_n810_), .Y(new_new_n935_));
  NA2        g913(.A(new_new_n918_), .B(new_new_n935_), .Y(new_new_n936_));
  AOI210     g914(.A0(new_new_n932_), .A1(new_new_n48_), .B0(new_new_n936_), .Y(new_new_n937_));
  AOI210     g915(.A0(new_new_n937_), .A1(new_new_n926_), .B0(new_new_n69_), .Y(new_new_n938_));
  INV        g916(.A(new_new_n533_), .Y(new_new_n939_));
  NO2        g917(.A(new_new_n939_), .B(new_new_n697_), .Y(new_new_n940_));
  NA2        g918(.A(new_new_n250_), .B(new_new_n53_), .Y(new_new_n941_));
  NA2        g919(.A(new_new_n941_), .B(new_new_n72_), .Y(new_new_n942_));
  NO2        g920(.A(new_new_n942_), .B(new_new_n226_), .Y(new_new_n943_));
  NA3        g921(.A(new_new_n93_), .B(new_new_n294_), .C(new_new_n31_), .Y(new_new_n944_));
  INV        g922(.A(new_new_n944_), .Y(new_new_n945_));
  NO2        g923(.A(new_new_n945_), .B(new_new_n943_), .Y(new_new_n946_));
  NA2        g924(.A(new_new_n152_), .B(new_new_n85_), .Y(new_new_n947_));
  NO2        g925(.A(new_new_n947_), .B(i_11_), .Y(new_new_n948_));
  OAI210     g926(.A0(new_new_n963_), .A1(new_new_n837_), .B0(new_new_n200_), .Y(new_new_n949_));
  NA2        g927(.A(new_new_n158_), .B(i_5_), .Y(new_new_n950_));
  NO2        g928(.A(new_new_n949_), .B(new_new_n950_), .Y(new_new_n951_));
  NO4        g929(.A(new_new_n861_), .B(new_new_n450_), .C(new_new_n240_), .D(new_new_n239_), .Y(new_new_n952_));
  NO2        g930(.A(new_new_n952_), .B(new_new_n530_), .Y(new_new_n953_));
  INV        g931(.A(new_new_n346_), .Y(new_new_n954_));
  AOI210     g932(.A0(new_new_n954_), .A1(new_new_n953_), .B0(new_new_n41_), .Y(new_new_n955_));
  NO3        g933(.A(new_new_n955_), .B(new_new_n951_), .C(new_new_n948_), .Y(new_new_n956_));
  OAI210     g934(.A0(new_new_n946_), .A1(i_4_), .B0(new_new_n956_), .Y(new_new_n957_));
  NO3        g935(.A(new_new_n957_), .B(new_new_n940_), .C(new_new_n938_), .Y(new_new_n958_));
  NA4        g936(.A(new_new_n958_), .B(new_new_n922_), .C(new_new_n868_), .D(new_new_n803_), .Y(mai4));
  INV        g937(.A(new_new_n789_), .Y(new_new_n962_));
  INV        g938(.A(i_12_), .Y(new_new_n963_));
endmodule


