//Benchmark atmr_5xp1_76_0.5

module atmr_5xp1(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
 wire ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n49_, ori_ori_n53_, ori_ori_n55_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n48_, mai_mai_n52_, mai_mai_n53_, mai_mai_n55_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n76_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n57_, men_men_n61_, men_men_n62_, men_men_n64_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09;
  INV        o00(.A(i_5_), .Y(ori_ori_n18_));
  INV        o01(.A(i_4_), .Y(ori_ori_n19_));
  NA2        o02(.A(ori_ori_n19_), .B(i_5_), .Y(ori_ori_n20_));
  INV        o03(.A(i_1_), .Y(ori_ori_n21_));
  AOI210     o04(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(ori_ori_n22_));
  INV        o05(.A(ori_ori_n20_), .Y(ori_ori_n23_));
  INV        o06(.A(i_6_), .Y(ori_ori_n24_));
  NO2        o07(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n25_));
  INV        o08(.A(i_0_), .Y(ori_ori_n26_));
  NO2        o09(.A(ori_ori_n19_), .B(i_5_), .Y(ori_ori_n27_));
  NO2        o10(.A(i_2_), .B(i_3_), .Y(ori_ori_n28_));
  NO3        o11(.A(ori_ori_n28_), .B(ori_ori_n26_), .C(ori_ori_n21_), .Y(ori_ori_n29_));
  AO210      o12(.A0(ori_ori_n29_), .A1(ori_ori_n27_), .B0(ori_ori_n25_), .Y(ori_ori_n30_));
  NA2        o13(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n31_));
  NA2        o14(.A(i_2_), .B(i_3_), .Y(ori_ori_n32_));
  NO2        o15(.A(ori_ori_n31_), .B(i_0_), .Y(ori_ori_n33_));
  OR3        o16(.A(ori_ori_n33_), .B(ori_ori_n30_), .C(ori_ori_n23_), .Y(ori01));
  NA2        o17(.A(i_0_), .B(i_1_), .Y(ori_ori_n35_));
  AOI210     o18(.A0(ori_ori_n22_), .A1(ori_ori_n21_), .B0(ori_ori_n24_), .Y(ori_ori_n36_));
  AOI220     o19(.A0(ori_ori_n36_), .A1(i_0_), .B0(ori_ori_n35_), .B1(ori_ori_n24_), .Y(ori_ori_n37_));
  NO2        o20(.A(ori_ori_n37_), .B(i_4_), .Y(ori_ori_n38_));
  NA2        o21(.A(i_0_), .B(i_6_), .Y(ori_ori_n39_));
  NO2        o22(.A(ori_ori_n70_), .B(ori_ori_n19_), .Y(ori_ori_n40_));
  NA2        o23(.A(ori_ori_n26_), .B(ori_ori_n24_), .Y(ori_ori_n41_));
  NO2        o24(.A(ori_ori_n41_), .B(ori_ori_n19_), .Y(ori_ori_n42_));
  INV        o25(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  OAI210     o26(.A0(ori_ori_n40_), .A1(ori_ori_n38_), .B0(ori_ori_n43_), .Y(ori02));
  NAi21      o27(.An(ori_ori_n20_), .B(ori_ori_n36_), .Y(ori_ori_n45_));
  NA3        o28(.A(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n46_));
  NO2        o29(.A(ori_ori_n42_), .B(ori_ori_n27_), .Y(ori_ori_n47_));
  NA2        o30(.A(ori_ori_n47_), .B(ori_ori_n45_), .Y(ori00));
  NA2        o31(.A(ori_ori_n41_), .B(i_5_), .Y(ori_ori_n49_));
  NO2        o32(.A(ori_ori_n49_), .B(ori_ori_n19_), .Y(ori09));
  NOi21      o33(.An(ori_ori_n32_), .B(ori_ori_n28_), .Y(ori07));
  INV        o34(.A(i_3_), .Y(ori08));
  INV        o35(.A(ori07), .Y(ori_ori_n53_));
  XO2        o36(.A(ori_ori_n53_), .B(ori_ori_n26_), .Y(ori05));
  NO2        o37(.A(i_2_), .B(ori08), .Y(ori_ori_n55_));
  XO2        o38(.A(ori_ori_n55_), .B(i_1_), .Y(ori06));
  NO2        o39(.A(i_1_), .B(i_6_), .Y(ori_ori_n57_));
  NO3        o40(.A(ori_ori_n57_), .B(i_0_), .C(ori_ori_n32_), .Y(ori_ori_n58_));
  NO2        o41(.A(ori_ori_n72_), .B(i_0_), .Y(ori_ori_n59_));
  INV        o42(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  NA3        o43(.A(ori_ori_n60_), .B(ori_ori_n18_), .C(ori_ori_n71_), .Y(ori03));
  NA2        o44(.A(ori_ori_n26_), .B(ori08), .Y(ori_ori_n62_));
  OAI210     o45(.A0(ori_ori_n62_), .A1(i_1_), .B0(ori_ori_n46_), .Y(ori_ori_n63_));
  OAI210     o46(.A0(ori_ori_n63_), .A1(ori_ori_n29_), .B0(i_6_), .Y(ori_ori_n64_));
  NA2        o47(.A(ori_ori_n62_), .B(ori_ori_n57_), .Y(ori_ori_n65_));
  NA3        o48(.A(ori_ori_n22_), .B(i_1_), .C(ori_ori_n24_), .Y(ori_ori_n66_));
  NA3        o49(.A(ori_ori_n66_), .B(ori_ori_n65_), .C(ori_ori_n64_), .Y(ori04));
  INV        o50(.A(ori_ori_n39_), .Y(ori_ori_n70_));
  INV        o51(.A(ori_ori_n58_), .Y(ori_ori_n71_));
  INV        o52(.A(i_6_), .Y(ori_ori_n72_));
  INV        m00(.A(i_5_), .Y(mai_mai_n18_));
  NO3        m01(.A(i_4_), .B(i_6_), .C(mai_mai_n18_), .Y(mai_mai_n19_));
  INV        m02(.A(i_4_), .Y(mai_mai_n20_));
  INV        m03(.A(i_1_), .Y(mai_mai_n21_));
  INV        m04(.A(i_6_), .Y(mai_mai_n22_));
  INV        m05(.A(i_0_), .Y(mai_mai_n23_));
  NO2        m06(.A(i_2_), .B(i_1_), .Y(mai_mai_n24_));
  NO2        m07(.A(mai_mai_n20_), .B(i_5_), .Y(mai00));
  NO2        m08(.A(i_2_), .B(i_3_), .Y(mai_mai_n26_));
  NO3        m09(.A(mai_mai_n26_), .B(mai_mai_n23_), .C(mai_mai_n21_), .Y(mai_mai_n27_));
  NA2        m10(.A(i_2_), .B(i_3_), .Y(mai_mai_n28_));
  OR2        m11(.A(mai00), .B(mai_mai_n19_), .Y(mai01));
  OR2        m12(.A(i_2_), .B(i_3_), .Y(mai_mai_n30_));
  NA3        m13(.A(mai_mai_n30_), .B(i_0_), .C(i_1_), .Y(mai_mai_n31_));
  NA2        m14(.A(mai_mai_n23_), .B(mai_mai_n18_), .Y(mai_mai_n32_));
  AOI220     m15(.A0(i_6_), .A1(mai_mai_n32_), .B0(mai_mai_n31_), .B1(mai_mai_n22_), .Y(mai_mai_n33_));
  NA2        m16(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n34_));
  OAI220     m17(.A0(mai_mai_n34_), .A1(mai_mai_n22_), .B0(mai_mai_n76_), .B1(mai_mai_n23_), .Y(mai_mai_n35_));
  NO3        m18(.A(mai_mai_n35_), .B(mai_mai_n33_), .C(i_4_), .Y(mai_mai_n36_));
  NA2        m19(.A(i_0_), .B(i_6_), .Y(mai_mai_n37_));
  OAI210     m20(.A0(i_0_), .A1(i_1_), .B0(mai_mai_n37_), .Y(mai_mai_n38_));
  NOi21      m21(.An(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n39_));
  NA3        m22(.A(i_1_), .B(i_6_), .C(i_5_), .Y(mai_mai_n40_));
  AOI210     m23(.A0(mai_mai_n40_), .A1(mai_mai_n37_), .B0(mai_mai_n24_), .Y(mai_mai_n41_));
  NO3        m24(.A(mai_mai_n30_), .B(i_6_), .C(i_5_), .Y(mai_mai_n42_));
  NO4        m25(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n39_), .D(mai_mai_n20_), .Y(mai_mai_n43_));
  AOI210     m26(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(mai_mai_n44_));
  AO220      m27(.A0(mai_mai_n44_), .A1(mai00), .B0(i_1_), .B1(mai_mai_n19_), .Y(mai_mai_n45_));
  INV        m28(.A(mai_mai_n45_), .Y(mai_mai_n46_));
  OAI210     m29(.A0(mai_mai_n43_), .A1(mai_mai_n36_), .B0(mai_mai_n46_), .Y(mai02));
  INV        m30(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m31(.A(mai_mai_n48_), .B(mai_mai_n20_), .Y(mai09));
  NOi21      m32(.An(mai_mai_n28_), .B(mai_mai_n26_), .Y(mai07));
  INV        m33(.A(i_3_), .Y(mai08));
  INV        m34(.A(mai_mai_n24_), .Y(mai_mai_n52_));
  NA2        m35(.A(mai07), .B(mai_mai_n52_), .Y(mai_mai_n53_));
  XO2        m36(.A(mai_mai_n53_), .B(mai_mai_n23_), .Y(mai05));
  NO2        m37(.A(i_2_), .B(mai08), .Y(mai_mai_n55_));
  XO2        m38(.A(mai_mai_n55_), .B(i_1_), .Y(mai06));
  NAi21      m39(.An(mai_mai_n42_), .B(mai_mai_n34_), .Y(mai_mai_n57_));
  NA2        m40(.A(mai_mai_n57_), .B(i_0_), .Y(mai_mai_n58_));
  NO2        m41(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NO3        m42(.A(mai_mai_n59_), .B(mai_mai_n32_), .C(mai_mai_n28_), .Y(mai_mai_n60_));
  INV        m43(.A(mai_mai_n60_), .Y(mai_mai_n61_));
  OR2        m44(.A(mai_mai_n31_), .B(mai_mai_n18_), .Y(mai_mai_n62_));
  NO2        m45(.A(mai_mai_n24_), .B(mai_mai_n23_), .Y(mai_mai_n63_));
  NO2        m46(.A(mai_mai_n22_), .B(mai_mai_n18_), .Y(mai_mai_n64_));
  OAI210     m47(.A0(mai_mai_n21_), .A1(i_6_), .B0(mai_mai_n18_), .Y(mai_mai_n65_));
  NO2        m48(.A(mai_mai_n65_), .B(mai_mai_n38_), .Y(mai_mai_n66_));
  AOI210     m49(.A0(mai_mai_n64_), .A1(mai_mai_n63_), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  NA4        m50(.A(mai_mai_n67_), .B(mai_mai_n62_), .C(mai_mai_n61_), .D(mai_mai_n58_), .Y(mai03));
  NA2        m51(.A(mai_mai_n27_), .B(i_6_), .Y(mai_mai_n69_));
  AOI210     m52(.A0(mai_mai_n26_), .A1(mai_mai_n22_), .B0(mai_mai_n24_), .Y(mai_mai_n70_));
  OR2        m53(.A(mai_mai_n70_), .B(mai_mai_n59_), .Y(mai_mai_n71_));
  NA2        m54(.A(mai_mai_n59_), .B(i_2_), .Y(mai_mai_n72_));
  NA3        m55(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(mai_mai_n69_), .Y(mai04));
  INV        m56(.A(i_5_), .Y(mai_mai_n76_));
  INV        u00(.A(i_5_), .Y(men_men_n18_));
  NO3        u01(.A(i_4_), .B(i_6_), .C(men_men_n18_), .Y(men_men_n19_));
  INV        u02(.A(i_4_), .Y(men_men_n20_));
  NA2        u03(.A(men_men_n20_), .B(i_5_), .Y(men_men_n21_));
  INV        u04(.A(i_1_), .Y(men_men_n22_));
  AOI210     u05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(men_men_n23_));
  NA2        u06(.A(men_men_n23_), .B(men_men_n22_), .Y(men_men_n24_));
  NO2        u07(.A(men_men_n24_), .B(men_men_n21_), .Y(men_men_n25_));
  INV        u08(.A(i_6_), .Y(men_men_n26_));
  NO2        u09(.A(men_men_n26_), .B(i_5_), .Y(men_men_n27_));
  INV        u10(.A(i_0_), .Y(men_men_n28_));
  NO2        u11(.A(i_2_), .B(i_1_), .Y(men_men_n29_));
  OAI210     u12(.A0(men_men_n29_), .A1(men_men_n28_), .B0(men_men_n20_), .Y(men_men_n30_));
  NO2        u13(.A(men_men_n20_), .B(i_5_), .Y(men_men_n31_));
  NO2        u14(.A(i_2_), .B(i_3_), .Y(men_men_n32_));
  AN2        u15(.A(men_men_n30_), .B(men_men_n27_), .Y(men_men_n33_));
  NA2        u16(.A(men_men_n26_), .B(i_5_), .Y(men_men_n34_));
  NA2        u17(.A(i_2_), .B(i_3_), .Y(men_men_n35_));
  NO2        u18(.A(men_men_n35_), .B(men_men_n22_), .Y(men_men_n36_));
  NO3        u19(.A(men_men_n36_), .B(men_men_n34_), .C(i_0_), .Y(men_men_n37_));
  OR4        u20(.A(men_men_n37_), .B(men_men_n33_), .C(men_men_n25_), .D(men_men_n19_), .Y(men01));
  AOI210     u21(.A0(men_men_n23_), .A1(men_men_n22_), .B0(men_men_n26_), .Y(men_men_n39_));
  NO2        u22(.A(men_men_n39_), .B(men_men_n26_), .Y(men_men_n40_));
  NA2        u23(.A(men_men_n29_), .B(men_men_n18_), .Y(men_men_n41_));
  OAI220     u24(.A0(men_men_n41_), .A1(men_men_n26_), .B0(men_men_n34_), .B1(men_men_n28_), .Y(men_men_n42_));
  NO3        u25(.A(men_men_n42_), .B(men_men_n40_), .C(i_4_), .Y(men_men_n43_));
  NOi31      u26(.An(i_6_), .B(men_men_n23_), .C(men_men_n18_), .Y(men_men_n44_));
  NA2        u27(.A(i_1_), .B(i_6_), .Y(men_men_n45_));
  NO2        u28(.A(men_men_n45_), .B(men_men_n29_), .Y(men_men_n46_));
  NO2        u29(.A(i_6_), .B(i_5_), .Y(men_men_n47_));
  NO4        u30(.A(men_men_n47_), .B(men_men_n46_), .C(men_men_n44_), .D(men_men_n20_), .Y(men_men_n48_));
  NO2        u31(.A(i_6_), .B(men_men_n20_), .Y(men_men_n49_));
  AN2        u32(.A(men_men_n36_), .B(men_men_n19_), .Y(men_men_n50_));
  AOI210     u33(.A0(men_men_n49_), .A1(men_men_n35_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u34(.A0(men_men_n48_), .A1(men_men_n43_), .B0(men_men_n51_), .Y(men02));
  NAi21      u35(.An(men_men_n21_), .B(men_men_n39_), .Y(men_men_n53_));
  NA3        u36(.A(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n54_));
  AOI210     u37(.A0(men_men_n49_), .A1(men_men_n54_), .B0(men_men_n31_), .Y(men_men_n55_));
  NA2        u38(.A(men_men_n55_), .B(men_men_n53_), .Y(men00));
  OAI210     u39(.A0(i_6_), .A1(men_men_n36_), .B0(i_5_), .Y(men_men_n57_));
  NO2        u40(.A(men_men_n57_), .B(men_men_n20_), .Y(men09));
  NOi21      u41(.An(men_men_n35_), .B(men_men_n32_), .Y(men07));
  INV        u42(.A(i_3_), .Y(men08));
  INV        u43(.A(men_men_n29_), .Y(men_men_n61_));
  NA2        u44(.A(men07), .B(men_men_n61_), .Y(men_men_n62_));
  XO2        u45(.A(men_men_n62_), .B(men_men_n28_), .Y(men05));
  NO2        u46(.A(i_2_), .B(men08), .Y(men_men_n64_));
  XO2        u47(.A(men_men_n64_), .B(i_1_), .Y(men06));
  NAi21      u48(.An(men_men_n47_), .B(men_men_n41_), .Y(men_men_n66_));
  NA2        u49(.A(men_men_n66_), .B(i_0_), .Y(men_men_n67_));
  NO2        u50(.A(i_1_), .B(i_6_), .Y(men_men_n68_));
  INV        u51(.A(men_men_n37_), .Y(men_men_n69_));
  OR2        u52(.A(men_men_n24_), .B(men_men_n18_), .Y(men_men_n70_));
  NO2        u53(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n71_));
  NO2        u54(.A(men_men_n26_), .B(men_men_n18_), .Y(men_men_n72_));
  NA2        u55(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n73_));
  NA4        u56(.A(men_men_n73_), .B(men_men_n70_), .C(men_men_n69_), .D(men_men_n67_), .Y(men03));
  INV        u57(.A(men_men_n68_), .Y(men04));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
endmodule