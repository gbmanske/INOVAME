//Benchmark atmr_misex3_1774_0.5

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n68_, ori_ori_n69_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  INV        o00(.A(n), .Y(ori_ori_n29_));
  NOi21      o01(.An(k), .B(m), .Y(ori_ori_n30_));
  INV        o02(.A(f), .Y(ori_ori_n31_));
  OR3        o03(.A(n), .B(m), .C(k), .Y(ori_ori_n32_));
  NO2        o04(.A(n), .B(m), .Y(ori_ori_n33_));
  BUFFER     o05(.A(f), .Y(ori_ori_n34_));
  NOi32      o06(.An(f), .Bn(c), .C(e), .Y(ori_ori_n35_));
  NOi31      o07(.An(k), .B(n), .C(m), .Y(ori12));
  NOi21      o08(.An(ori12), .B(ori_ori_n34_), .Y(ori_ori_n37_));
  INV        o09(.A(ori_ori_n37_), .Y(ori_ori_n38_));
  NAi31      o10(.An(f), .B(e), .C(c), .Y(ori_ori_n39_));
  NO2        o11(.A(ori_ori_n39_), .B(ori_ori_n32_), .Y(ori_ori_n40_));
  INV        o12(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  AN2        o13(.A(ori_ori_n41_), .B(ori_ori_n38_), .Y(ori_ori_n42_));
  NA2        o14(.A(ori_ori_n30_), .B(i), .Y(ori_ori_n43_));
  NA2        o15(.A(ori_ori_n33_), .B(ori_ori_n35_), .Y(ori_ori_n44_));
  NO2        o16(.A(n), .B(m), .Y(ori_ori_n45_));
  NA2        o17(.A(ori_ori_n44_), .B(ori_ori_n42_), .Y(ori10));
  NOi32      o18(.An(f), .Bn(d), .C(c), .Y(ori_ori_n47_));
  NA2        o19(.A(ori_ori_n33_), .B(ori_ori_n82_), .Y(ori_ori_n48_));
  INV        o20(.A(f), .Y(ori_ori_n49_));
  NA2        o21(.A(ori12), .B(i), .Y(ori_ori_n50_));
  NA2        o22(.A(ori_ori_n42_), .B(ori_ori_n48_), .Y(ori11));
  NOi32      o23(.An(e), .Bn(c), .C(f), .Y(ori_ori_n52_));
  NO2        o24(.A(ori_ori_n47_), .B(ori_ori_n35_), .Y(ori_ori_n53_));
  NA2        o25(.A(ori_ori_n53_), .B(ori_ori_n39_), .Y(ori_ori_n54_));
  NA2        o26(.A(ori_ori_n54_), .B(ori_ori_n33_), .Y(ori_ori_n55_));
  INV        o27(.A(ori_ori_n55_), .Y(ori08));
  NO2        o28(.A(ori_ori_n81_), .B(m), .Y(ori_ori_n57_));
  NA2        o29(.A(ori_ori_n52_), .B(ori_ori_n29_), .Y(ori_ori_n58_));
  INV        o30(.A(ori_ori_n58_), .Y(ori_ori_n59_));
  NA2        o31(.A(ori_ori_n59_), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o32(.A(ori_ori_n60_), .Y(ori_ori_n61_));
  NA3        o33(.A(ori_ori_n54_), .B(ori_ori_n45_), .C(k), .Y(ori_ori_n62_));
  INV        o34(.A(ori_ori_n62_), .Y(ori_ori_n63_));
  NO2        o35(.A(ori_ori_n63_), .B(ori_ori_n61_), .Y(ori_ori_n64_));
  NO2        o36(.A(ori_ori_n53_), .B(n), .Y(ori_ori_n65_));
  NA2        o37(.A(ori_ori_n65_), .B(ori_ori_n57_), .Y(ori_ori_n66_));
  NA2        o38(.A(ori_ori_n66_), .B(ori_ori_n64_), .Y(ori09));
  INV        o39(.A(ori_ori_n39_), .Y(ori_ori_n68_));
  NA2        o40(.A(ori_ori_n68_), .B(ori12), .Y(ori_ori_n69_));
  INV        o41(.A(ori_ori_n69_), .Y(ori06));
  NO2        o42(.A(ori_ori_n50_), .B(ori_ori_n31_), .Y(ori_ori_n71_));
  INV        o43(.A(ori_ori_n71_), .Y(ori_ori_n72_));
  OAI220     o44(.A0(ori_ori_n58_), .A1(ori_ori_n43_), .B0(ori_ori_n49_), .B1(ori_ori_n50_), .Y(ori_ori_n73_));
  NA2        o45(.A(ori_ori_n78_), .B(ori_ori_n72_), .Y(ori07));
  OR2        o46(.A(ori_ori_n80_), .B(ori_ori_n79_), .Y(ori04));
  INV        o47(.A(ori_ori_n73_), .Y(ori_ori_n78_));
  INV        o48(.A(n), .Y(ori_ori_n79_));
  INV        o49(.A(m), .Y(ori_ori_n80_));
  INV        o50(.A(j), .Y(ori_ori_n81_));
  INV        o51(.A(e), .Y(ori_ori_n82_));
  ZERO       o52(.Y(ori13));
  ZERO       o53(.Y(ori02));
  ZERO       o54(.Y(ori03));
  ZERO       o55(.Y(ori00));
  ZERO       o56(.Y(ori01));
  ZERO       o57(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  AN2        m0001(.A(f), .B(e), .Y(mai_mai_n30_));
  NA2        m0002(.A(mai_mai_n30_), .B(mai_mai_n29_), .Y(mai_mai_n31_));
  NOi32      m0003(.An(m), .Bn(l), .C(n), .Y(mai_mai_n32_));
  NOi32      m0004(.An(i), .Bn(m), .C(h), .Y(mai_mai_n33_));
  NOi32      m0005(.An(j), .Bn(m), .C(k), .Y(mai_mai_n34_));
  INV        m0006(.A(h), .Y(mai_mai_n35_));
  NAi21      m0007(.An(n), .B(m), .Y(mai_mai_n36_));
  INV        m0008(.A(i), .Y(mai_mai_n37_));
  AN2        m0009(.A(h), .B(m), .Y(mai_mai_n38_));
  NAi21      m0010(.An(n), .B(m), .Y(mai_mai_n39_));
  NOi32      m0011(.An(k), .Bn(h), .C(l), .Y(mai_mai_n40_));
  NOi32      m0012(.An(k), .Bn(h), .C(m), .Y(mai_mai_n41_));
  INV        m0013(.A(mai_mai_n39_), .Y(mai_mai_n42_));
  NO2        m0014(.A(mai_mai_n39_), .B(mai_mai_n31_), .Y(mai_mai_n43_));
  INV        m0015(.A(c), .Y(mai_mai_n44_));
  NA2        m0016(.A(e), .B(b), .Y(mai_mai_n45_));
  INV        m0017(.A(d), .Y(mai_mai_n46_));
  NAi21      m0018(.An(i), .B(h), .Y(mai_mai_n47_));
  NAi32      m0019(.An(n), .Bn(k), .C(m), .Y(mai_mai_n48_));
  NAi31      m0020(.An(l), .B(m), .C(k), .Y(mai_mai_n49_));
  NAi41      m0021(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n50_));
  INV        m0022(.A(m), .Y(mai_mai_n51_));
  NOi21      m0023(.An(k), .B(l), .Y(mai_mai_n52_));
  NA2        m0024(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  AN4        m0025(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n54_));
  NOi31      m0026(.An(h), .B(m), .C(f), .Y(mai_mai_n55_));
  NA2        m0027(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NAi32      m0028(.An(m), .Bn(k), .C(j), .Y(mai_mai_n57_));
  NOi32      m0029(.An(h), .Bn(m), .C(f), .Y(mai_mai_n58_));
  NA2        m0030(.A(mai_mai_n58_), .B(mai_mai_n54_), .Y(mai_mai_n59_));
  OA220      m0031(.A0(mai_mai_n59_), .A1(mai_mai_n57_), .B0(mai_mai_n56_), .B1(mai_mai_n53_), .Y(mai_mai_n60_));
  INV        m0032(.A(mai_mai_n60_), .Y(mai_mai_n61_));
  INV        m0033(.A(n), .Y(mai_mai_n62_));
  NOi32      m0034(.An(e), .Bn(b), .C(d), .Y(mai_mai_n63_));
  INV        m0035(.A(j), .Y(mai_mai_n64_));
  AN3        m0036(.A(m), .B(k), .C(i), .Y(mai_mai_n65_));
  NA3        m0037(.A(mai_mai_n65_), .B(mai_mai_n64_), .C(m), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(f), .Y(mai_mai_n67_));
  NAi32      m0039(.An(m), .Bn(f), .C(h), .Y(mai_mai_n68_));
  NAi31      m0040(.An(j), .B(m), .C(l), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NA2        m0042(.A(m), .B(l), .Y(mai_mai_n71_));
  NAi31      m0043(.An(k), .B(j), .C(m), .Y(mai_mai_n72_));
  NO3        m0044(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(f), .Y(mai_mai_n73_));
  NOi21      m0045(.An(m), .B(i), .Y(mai_mai_n74_));
  NOi32      m0046(.An(m), .Bn(j), .C(k), .Y(mai_mai_n75_));
  NA2        m0047(.A(m), .B(m), .Y(mai_mai_n76_));
  NO2        m0048(.A(mai_mai_n76_), .B(f), .Y(mai_mai_n77_));
  NAi41      m0049(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n78_));
  AN2        m0050(.A(e), .B(b), .Y(mai_mai_n79_));
  NOi31      m0051(.An(c), .B(h), .C(f), .Y(mai_mai_n80_));
  NA2        m0052(.A(mai_mai_n80_), .B(mai_mai_n79_), .Y(mai_mai_n81_));
  NOi21      m0053(.An(m), .B(f), .Y(mai_mai_n82_));
  NOi21      m0054(.An(i), .B(h), .Y(mai_mai_n83_));
  INV        m0055(.A(a), .Y(mai_mai_n84_));
  NA2        m0056(.A(mai_mai_n79_), .B(mai_mai_n84_), .Y(mai_mai_n85_));
  INV        m0057(.A(l), .Y(mai_mai_n86_));
  NOi21      m0058(.An(m), .B(n), .Y(mai_mai_n87_));
  AN2        m0059(.A(k), .B(h), .Y(mai_mai_n88_));
  INV        m0060(.A(b), .Y(mai_mai_n89_));
  NA2        m0061(.A(l), .B(j), .Y(mai_mai_n90_));
  NOi32      m0062(.An(c), .Bn(a), .C(d), .Y(mai_mai_n91_));
  NA2        m0063(.A(mai_mai_n91_), .B(mai_mai_n87_), .Y(mai_mai_n92_));
  NOi31      m0064(.An(k), .B(m), .C(j), .Y(mai_mai_n93_));
  NA3        m0065(.A(mai_mai_n93_), .B(mai_mai_n55_), .C(mai_mai_n54_), .Y(mai_mai_n94_));
  NOi31      m0066(.An(k), .B(m), .C(i), .Y(mai_mai_n95_));
  NA3        m0067(.A(mai_mai_n95_), .B(mai_mai_n58_), .C(mai_mai_n54_), .Y(mai_mai_n96_));
  NA2        m0068(.A(mai_mai_n96_), .B(mai_mai_n94_), .Y(mai_mai_n97_));
  NOi32      m0069(.An(f), .Bn(b), .C(e), .Y(mai_mai_n98_));
  NAi21      m0070(.An(m), .B(n), .Y(mai_mai_n99_));
  NAi21      m0071(.An(j), .B(k), .Y(mai_mai_n100_));
  NO3        m0072(.A(mai_mai_n100_), .B(mai_mai_n99_), .C(m), .Y(mai_mai_n101_));
  NAi41      m0073(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n102_));
  NAi31      m0074(.An(j), .B(k), .C(h), .Y(mai_mai_n103_));
  NO3        m0075(.A(mai_mai_n103_), .B(mai_mai_n102_), .C(mai_mai_n99_), .Y(mai_mai_n104_));
  AOI210     m0076(.A0(mai_mai_n101_), .A1(mai_mai_n98_), .B0(mai_mai_n104_), .Y(mai_mai_n105_));
  NO2        m0077(.A(k), .B(j), .Y(mai_mai_n106_));
  NO2        m0078(.A(mai_mai_n106_), .B(mai_mai_n99_), .Y(mai_mai_n107_));
  AN2        m0079(.A(k), .B(j), .Y(mai_mai_n108_));
  NAi21      m0080(.An(c), .B(b), .Y(mai_mai_n109_));
  NA2        m0081(.A(f), .B(d), .Y(mai_mai_n110_));
  NO4        m0082(.A(mai_mai_n110_), .B(mai_mai_n109_), .C(mai_mai_n108_), .D(m), .Y(mai_mai_n111_));
  NAi31      m0083(.An(f), .B(e), .C(b), .Y(mai_mai_n112_));
  NA2        m0084(.A(mai_mai_n111_), .B(mai_mai_n107_), .Y(mai_mai_n113_));
  NA2        m0085(.A(d), .B(b), .Y(mai_mai_n114_));
  NAi21      m0086(.An(e), .B(f), .Y(mai_mai_n115_));
  NA2        m0087(.A(b), .B(a), .Y(mai_mai_n116_));
  NAi21      m0088(.An(e), .B(m), .Y(mai_mai_n117_));
  NAi21      m0089(.An(c), .B(d), .Y(mai_mai_n118_));
  NAi31      m0090(.An(l), .B(k), .C(h), .Y(mai_mai_n119_));
  NO2        m0091(.A(mai_mai_n99_), .B(mai_mai_n119_), .Y(mai_mai_n120_));
  NAi31      m0092(.An(mai_mai_n97_), .B(mai_mai_n113_), .C(mai_mai_n105_), .Y(mai_mai_n121_));
  NAi31      m0093(.An(e), .B(f), .C(b), .Y(mai_mai_n122_));
  NOi21      m0094(.An(m), .B(d), .Y(mai_mai_n123_));
  NO2        m0095(.A(mai_mai_n123_), .B(mai_mai_n122_), .Y(mai_mai_n124_));
  NOi21      m0096(.An(h), .B(i), .Y(mai_mai_n125_));
  NOi21      m0097(.An(k), .B(m), .Y(mai_mai_n126_));
  NA3        m0098(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(n), .Y(mai_mai_n127_));
  NOi21      m0099(.An(mai_mai_n124_), .B(mai_mai_n127_), .Y(mai_mai_n128_));
  NOi21      m0100(.An(h), .B(m), .Y(mai_mai_n129_));
  INV        m0101(.A(mai_mai_n109_), .Y(mai_mai_n130_));
  NA2        m0102(.A(mai_mai_n130_), .B(mai_mai_n129_), .Y(mai_mai_n131_));
  NOi32      m0103(.An(n), .Bn(k), .C(m), .Y(mai_mai_n132_));
  NA2        m0104(.A(l), .B(i), .Y(mai_mai_n133_));
  NA2        m0105(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n134_));
  NO2        m0106(.A(mai_mai_n134_), .B(mai_mai_n131_), .Y(mai_mai_n135_));
  NAi31      m0107(.An(d), .B(f), .C(c), .Y(mai_mai_n136_));
  NAi31      m0108(.An(e), .B(f), .C(c), .Y(mai_mai_n137_));
  NA2        m0109(.A(j), .B(h), .Y(mai_mai_n138_));
  OR3        m0110(.A(n), .B(m), .C(k), .Y(mai_mai_n139_));
  NO2        m0111(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n140_));
  NAi32      m0112(.An(m), .Bn(k), .C(n), .Y(mai_mai_n141_));
  NO2        m0113(.A(mai_mai_n141_), .B(mai_mai_n138_), .Y(mai_mai_n142_));
  AOI220     m0114(.A0(mai_mai_n142_), .A1(mai_mai_n124_), .B0(mai_mai_n140_), .B1(f), .Y(mai_mai_n143_));
  NO2        m0115(.A(n), .B(m), .Y(mai_mai_n144_));
  NA2        m0116(.A(mai_mai_n144_), .B(mai_mai_n40_), .Y(mai_mai_n145_));
  NAi21      m0117(.An(f), .B(e), .Y(mai_mai_n146_));
  NA2        m0118(.A(d), .B(c), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n147_), .B(mai_mai_n146_), .Y(mai_mai_n148_));
  NOi21      m0120(.An(mai_mai_n148_), .B(mai_mai_n145_), .Y(mai_mai_n149_));
  NAi31      m0121(.An(m), .B(n), .C(b), .Y(mai_mai_n150_));
  NA2        m0122(.A(k), .B(i), .Y(mai_mai_n151_));
  NAi21      m0123(.An(h), .B(f), .Y(mai_mai_n152_));
  INV        m0124(.A(mai_mai_n152_), .Y(mai_mai_n153_));
  NO2        m0125(.A(mai_mai_n150_), .B(mai_mai_n118_), .Y(mai_mai_n154_));
  NA2        m0126(.A(mai_mai_n154_), .B(mai_mai_n153_), .Y(mai_mai_n155_));
  NOi32      m0127(.An(f), .Bn(c), .C(d), .Y(mai_mai_n156_));
  NOi32      m0128(.An(f), .Bn(c), .C(e), .Y(mai_mai_n157_));
  NO2        m0129(.A(mai_mai_n157_), .B(mai_mai_n156_), .Y(mai_mai_n158_));
  NO3        m0130(.A(n), .B(m), .C(j), .Y(mai_mai_n159_));
  NA2        m0131(.A(mai_mai_n159_), .B(mai_mai_n88_), .Y(mai_mai_n160_));
  AO210      m0132(.A0(mai_mai_n160_), .A1(mai_mai_n145_), .B0(mai_mai_n158_), .Y(mai_mai_n161_));
  NAi41      m0133(.An(mai_mai_n149_), .B(mai_mai_n161_), .C(mai_mai_n155_), .D(mai_mai_n143_), .Y(mai_mai_n162_));
  OR3        m0134(.A(mai_mai_n162_), .B(mai_mai_n135_), .C(mai_mai_n121_), .Y(mai_mai_n163_));
  NO3        m0135(.A(mai_mai_n163_), .B(mai_mai_n61_), .C(mai_mai_n43_), .Y(mai_mai_n164_));
  NAi31      m0136(.An(n), .B(h), .C(m), .Y(mai_mai_n165_));
  NOi32      m0137(.An(m), .Bn(k), .C(l), .Y(mai_mai_n166_));
  NA3        m0138(.A(mai_mai_n166_), .B(mai_mai_n64_), .C(m), .Y(mai_mai_n167_));
  NOi21      m0139(.An(k), .B(j), .Y(mai_mai_n168_));
  AN2        m0140(.A(i), .B(m), .Y(mai_mai_n169_));
  NAi41      m0141(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n170_));
  INV        m0142(.A(mai_mai_n170_), .Y(mai_mai_n171_));
  INV        m0143(.A(f), .Y(mai_mai_n172_));
  INV        m0144(.A(m), .Y(mai_mai_n173_));
  NOi31      m0145(.An(i), .B(j), .C(h), .Y(mai_mai_n174_));
  NOi21      m0146(.An(l), .B(m), .Y(mai_mai_n175_));
  NA2        m0147(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n176_), .B(mai_mai_n173_), .Y(mai_mai_n177_));
  NA2        m0149(.A(mai_mai_n177_), .B(mai_mai_n171_), .Y(mai_mai_n178_));
  INV        m0150(.A(mai_mai_n178_), .Y(mai_mai_n179_));
  NOi21      m0151(.An(n), .B(m), .Y(mai_mai_n180_));
  NA2        m0152(.A(i), .B(mai_mai_n180_), .Y(mai_mai_n181_));
  OA220      m0153(.A0(mai_mai_n181_), .A1(mai_mai_n81_), .B0(mai_mai_n57_), .B1(mai_mai_n56_), .Y(mai_mai_n182_));
  NAi21      m0154(.An(j), .B(h), .Y(mai_mai_n183_));
  XN2        m0155(.A(i), .B(h), .Y(mai_mai_n184_));
  NA2        m0156(.A(mai_mai_n184_), .B(mai_mai_n183_), .Y(mai_mai_n185_));
  NOi31      m0157(.An(k), .B(n), .C(m), .Y(mai_mai_n186_));
  NOi31      m0158(.An(mai_mai_n186_), .B(mai_mai_n147_), .C(mai_mai_n146_), .Y(mai_mai_n187_));
  NA2        m0159(.A(mai_mai_n187_), .B(mai_mai_n185_), .Y(mai_mai_n188_));
  NAi31      m0160(.An(f), .B(e), .C(c), .Y(mai_mai_n189_));
  NO4        m0161(.A(mai_mai_n189_), .B(mai_mai_n139_), .C(mai_mai_n138_), .D(mai_mai_n46_), .Y(mai_mai_n190_));
  NA4        m0162(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n191_));
  NAi32      m0163(.An(m), .Bn(i), .C(k), .Y(mai_mai_n192_));
  NO3        m0164(.A(mai_mai_n192_), .B(mai_mai_n68_), .C(mai_mai_n191_), .Y(mai_mai_n193_));
  NA2        m0165(.A(k), .B(h), .Y(mai_mai_n194_));
  NO2        m0166(.A(mai_mai_n193_), .B(mai_mai_n190_), .Y(mai_mai_n195_));
  NAi21      m0167(.An(n), .B(a), .Y(mai_mai_n196_));
  NAi41      m0168(.An(m), .B(m), .C(k), .D(h), .Y(mai_mai_n197_));
  AN3        m0169(.A(mai_mai_n195_), .B(mai_mai_n188_), .C(mai_mai_n182_), .Y(mai_mai_n198_));
  OR2        m0170(.A(h), .B(m), .Y(mai_mai_n199_));
  NO2        m0171(.A(mai_mai_n199_), .B(mai_mai_n78_), .Y(mai_mai_n200_));
  NA2        m0172(.A(mai_mai_n200_), .B(mai_mai_n98_), .Y(mai_mai_n201_));
  NAi41      m0173(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n202_));
  NO2        m0174(.A(mai_mai_n202_), .B(mai_mai_n172_), .Y(mai_mai_n203_));
  NA2        m0175(.A(mai_mai_n126_), .B(mai_mai_n83_), .Y(mai_mai_n204_));
  NAi21      m0176(.An(mai_mai_n204_), .B(mai_mai_n203_), .Y(mai_mai_n205_));
  NO2        m0177(.A(n), .B(a), .Y(mai_mai_n206_));
  NAi31      m0178(.An(mai_mai_n197_), .B(mai_mai_n206_), .C(mai_mai_n79_), .Y(mai_mai_n207_));
  AN2        m0179(.A(mai_mai_n207_), .B(mai_mai_n205_), .Y(mai_mai_n208_));
  NAi21      m0180(.An(h), .B(i), .Y(mai_mai_n209_));
  NA2        m0181(.A(mai_mai_n144_), .B(k), .Y(mai_mai_n210_));
  NO2        m0182(.A(mai_mai_n210_), .B(mai_mai_n209_), .Y(mai_mai_n211_));
  NA2        m0183(.A(mai_mai_n211_), .B(mai_mai_n156_), .Y(mai_mai_n212_));
  NA3        m0184(.A(mai_mai_n212_), .B(mai_mai_n208_), .C(mai_mai_n201_), .Y(mai_mai_n213_));
  NOi21      m0185(.An(m), .B(e), .Y(mai_mai_n214_));
  NO2        m0186(.A(mai_mai_n50_), .B(mai_mai_n51_), .Y(mai_mai_n215_));
  NO2        m0187(.A(mai_mai_n100_), .B(mai_mai_n39_), .Y(mai_mai_n216_));
  NOi31      m0188(.An(mai_mai_n198_), .B(mai_mai_n213_), .C(mai_mai_n179_), .Y(mai_mai_n217_));
  NO2        m0189(.A(mai_mai_n36_), .B(mai_mai_n85_), .Y(mai_mai_n218_));
  NA3        m0190(.A(mai_mai_n46_), .B(c), .C(b), .Y(mai_mai_n219_));
  OR4        m0191(.A(h), .B(mai_mai_n219_), .C(mai_mai_n181_), .D(e), .Y(mai_mai_n220_));
  NO2        m0192(.A(mai_mai_n204_), .B(f), .Y(mai_mai_n221_));
  NAi31      m0193(.An(m), .B(k), .C(h), .Y(mai_mai_n222_));
  NO3        m0194(.A(mai_mai_n99_), .B(mai_mai_n222_), .C(l), .Y(mai_mai_n223_));
  NAi31      m0195(.An(e), .B(d), .C(a), .Y(mai_mai_n224_));
  NA2        m0196(.A(mai_mai_n223_), .B(mai_mai_n98_), .Y(mai_mai_n225_));
  NA2        m0197(.A(mai_mai_n225_), .B(mai_mai_n220_), .Y(mai_mai_n226_));
  NA4        m0198(.A(mai_mai_n126_), .B(mai_mai_n58_), .C(mai_mai_n54_), .D(mai_mai_n90_), .Y(mai_mai_n227_));
  NA3        m0199(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(mai_mai_n62_), .Y(mai_mai_n228_));
  NO2        m0200(.A(mai_mai_n228_), .B(mai_mai_n158_), .Y(mai_mai_n229_));
  NOi21      m0201(.An(mai_mai_n227_), .B(mai_mai_n229_), .Y(mai_mai_n230_));
  NA3        m0202(.A(e), .B(c), .C(b), .Y(mai_mai_n231_));
  NAi32      m0203(.An(k), .Bn(i), .C(j), .Y(mai_mai_n232_));
  NOi21      m0204(.An(l), .B(j), .Y(mai_mai_n233_));
  OR3        m0205(.A(mai_mai_n50_), .B(mai_mai_n51_), .C(e), .Y(mai_mai_n234_));
  NAi32      m0206(.An(j), .Bn(h), .C(i), .Y(mai_mai_n235_));
  NAi21      m0207(.An(m), .B(l), .Y(mai_mai_n236_));
  NO3        m0208(.A(mai_mai_n236_), .B(mai_mai_n235_), .C(mai_mai_n62_), .Y(mai_mai_n237_));
  NA2        m0209(.A(h), .B(m), .Y(mai_mai_n238_));
  NA2        m0210(.A(mai_mai_n132_), .B(mai_mai_n37_), .Y(mai_mai_n239_));
  NA3        m0211(.A(mai_mai_n239_), .B(mai_mai_n234_), .C(mai_mai_n230_), .Y(mai_mai_n240_));
  NO2        m0212(.A(mai_mai_n112_), .B(d), .Y(mai_mai_n241_));
  NA2        m0213(.A(mai_mai_n241_), .B(mai_mai_n42_), .Y(mai_mai_n242_));
  NAi32      m0214(.An(n), .Bn(m), .C(l), .Y(mai_mai_n243_));
  NO2        m0215(.A(mai_mai_n243_), .B(mai_mai_n235_), .Y(mai_mai_n244_));
  NA2        m0216(.A(mai_mai_n244_), .B(mai_mai_n148_), .Y(mai_mai_n245_));
  NA2        m0217(.A(mai_mai_n245_), .B(mai_mai_n242_), .Y(mai_mai_n246_));
  NO4        m0218(.A(mai_mai_n246_), .B(mai_mai_n240_), .C(mai_mai_n226_), .D(mai_mai_n218_), .Y(mai_mai_n247_));
  NA2        m0219(.A(mai_mai_n211_), .B(mai_mai_n157_), .Y(mai_mai_n248_));
  NAi21      m0220(.An(m), .B(k), .Y(mai_mai_n249_));
  NO2        m0221(.A(mai_mai_n184_), .B(mai_mai_n249_), .Y(mai_mai_n250_));
  NAi41      m0222(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n251_));
  NO2        m0223(.A(mai_mai_n251_), .B(mai_mai_n117_), .Y(mai_mai_n252_));
  NA2        m0224(.A(mai_mai_n252_), .B(mai_mai_n250_), .Y(mai_mai_n253_));
  NA2        m0225(.A(e), .B(c), .Y(mai_mai_n254_));
  NO3        m0226(.A(mai_mai_n254_), .B(n), .C(d), .Y(mai_mai_n255_));
  NOi21      m0227(.An(f), .B(h), .Y(mai_mai_n256_));
  NA2        m0228(.A(mai_mai_n256_), .B(k), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n257_), .B(mai_mai_n173_), .Y(mai_mai_n258_));
  NAi31      m0230(.An(d), .B(e), .C(b), .Y(mai_mai_n259_));
  NO2        m0231(.A(mai_mai_n99_), .B(mai_mai_n259_), .Y(mai_mai_n260_));
  NA2        m0232(.A(mai_mai_n260_), .B(mai_mai_n258_), .Y(mai_mai_n261_));
  NA3        m0233(.A(mai_mai_n261_), .B(mai_mai_n253_), .C(mai_mai_n248_), .Y(mai_mai_n262_));
  NO4        m0234(.A(mai_mai_n251_), .B(mai_mai_n57_), .C(e), .D(mai_mai_n173_), .Y(mai_mai_n263_));
  NA2        m0235(.A(mai_mai_n206_), .B(mai_mai_n79_), .Y(mai_mai_n264_));
  NOi31      m0236(.An(l), .B(n), .C(m), .Y(mai_mai_n265_));
  NA2        m0237(.A(mai_mai_n265_), .B(mai_mai_n174_), .Y(mai_mai_n266_));
  NO2        m0238(.A(mai_mai_n266_), .B(mai_mai_n158_), .Y(mai_mai_n267_));
  OR2        m0239(.A(mai_mai_n267_), .B(mai_mai_n263_), .Y(mai_mai_n268_));
  NAi32      m0240(.An(m), .Bn(j), .C(k), .Y(mai_mai_n269_));
  NAi41      m0241(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n270_));
  NA2        m0242(.A(mai_mai_n170_), .B(mai_mai_n270_), .Y(mai_mai_n271_));
  NOi31      m0243(.An(j), .B(m), .C(k), .Y(mai_mai_n272_));
  NO2        m0244(.A(mai_mai_n93_), .B(mai_mai_n272_), .Y(mai_mai_n273_));
  AN3        m0245(.A(h), .B(m), .C(f), .Y(mai_mai_n274_));
  NAi31      m0246(.An(mai_mai_n273_), .B(mai_mai_n274_), .C(mai_mai_n271_), .Y(mai_mai_n275_));
  NO2        m0247(.A(mai_mai_n236_), .B(mai_mai_n235_), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n176_), .B(m), .Y(mai_mai_n277_));
  NO2        m0249(.A(mai_mai_n122_), .B(mai_mai_n62_), .Y(mai_mai_n278_));
  AOI220     m0250(.A0(mai_mai_n278_), .A1(mai_mai_n277_), .B0(mai_mai_n203_), .B1(mai_mai_n276_), .Y(mai_mai_n279_));
  INV        m0251(.A(mai_mai_n192_), .Y(mai_mai_n280_));
  NA2        m0252(.A(mai_mai_n280_), .B(mai_mai_n171_), .Y(mai_mai_n281_));
  NA3        m0253(.A(mai_mai_n281_), .B(mai_mai_n279_), .C(mai_mai_n275_), .Y(mai_mai_n282_));
  NA3        m0254(.A(h), .B(m), .C(f), .Y(mai_mai_n283_));
  NO2        m0255(.A(mai_mai_n283_), .B(mai_mai_n53_), .Y(mai_mai_n284_));
  NA2        m0256(.A(n), .B(mai_mai_n284_), .Y(mai_mai_n285_));
  NA2        m0257(.A(m), .B(mai_mai_n87_), .Y(mai_mai_n286_));
  NOi32      m0258(.An(e), .Bn(b), .C(a), .Y(mai_mai_n287_));
  AN2        m0259(.A(l), .B(j), .Y(mai_mai_n288_));
  NO2        m0260(.A(mai_mai_n249_), .B(mai_mai_n288_), .Y(mai_mai_n289_));
  NO3        m0261(.A(mai_mai_n251_), .B(e), .C(mai_mai_n173_), .Y(mai_mai_n290_));
  NA2        m0262(.A(mai_mai_n290_), .B(mai_mai_n289_), .Y(mai_mai_n291_));
  NO2        m0263(.A(mai_mai_n259_), .B(n), .Y(mai_mai_n292_));
  NA2        m0264(.A(mai_mai_n169_), .B(k), .Y(mai_mai_n293_));
  NA3        m0265(.A(m), .B(mai_mai_n86_), .C(mai_mai_n172_), .Y(mai_mai_n294_));
  NA4        m0266(.A(mai_mai_n166_), .B(mai_mai_n64_), .C(m), .D(mai_mai_n172_), .Y(mai_mai_n295_));
  NAi41      m0267(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n41_), .B(mai_mai_n87_), .Y(mai_mai_n297_));
  NO2        m0269(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n298_));
  NA2        m0270(.A(mai_mai_n166_), .B(mai_mai_n292_), .Y(mai_mai_n299_));
  NA3        m0271(.A(mai_mai_n299_), .B(mai_mai_n291_), .C(mai_mai_n285_), .Y(mai_mai_n300_));
  NO4        m0272(.A(mai_mai_n300_), .B(mai_mai_n282_), .C(mai_mai_n268_), .D(mai_mai_n262_), .Y(mai_mai_n301_));
  NA4        m0273(.A(mai_mai_n301_), .B(mai_mai_n247_), .C(mai_mai_n217_), .D(mai_mai_n164_), .Y(mai10));
  NA3        m0274(.A(m), .B(k), .C(i), .Y(mai_mai_n303_));
  NO3        m0275(.A(mai_mai_n303_), .B(j), .C(mai_mai_n173_), .Y(mai_mai_n304_));
  NOi21      m0276(.An(e), .B(f), .Y(mai_mai_n305_));
  NO4        m0277(.A(mai_mai_n118_), .B(mai_mai_n305_), .C(n), .D(mai_mai_n84_), .Y(mai_mai_n306_));
  NAi31      m0278(.An(b), .B(f), .C(c), .Y(mai_mai_n307_));
  INV        m0279(.A(mai_mai_n307_), .Y(mai_mai_n308_));
  NOi32      m0280(.An(k), .Bn(h), .C(j), .Y(mai_mai_n309_));
  NA2        m0281(.A(mai_mai_n309_), .B(mai_mai_n180_), .Y(mai_mai_n310_));
  NA2        m0282(.A(mai_mai_n127_), .B(mai_mai_n310_), .Y(mai_mai_n311_));
  AOI220     m0283(.A0(mai_mai_n311_), .A1(mai_mai_n308_), .B0(mai_mai_n306_), .B1(mai_mai_n304_), .Y(mai_mai_n312_));
  AN2        m0284(.A(j), .B(h), .Y(mai_mai_n313_));
  NO3        m0285(.A(n), .B(m), .C(k), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n314_), .B(mai_mai_n313_), .Y(mai_mai_n315_));
  NO3        m0287(.A(mai_mai_n315_), .B(mai_mai_n118_), .C(mai_mai_n172_), .Y(mai_mai_n316_));
  OR2        m0288(.A(m), .B(k), .Y(mai_mai_n317_));
  NO2        m0289(.A(mai_mai_n138_), .B(mai_mai_n317_), .Y(mai_mai_n318_));
  NA4        m0290(.A(n), .B(f), .C(c), .D(mai_mai_n89_), .Y(mai_mai_n319_));
  NOi21      m0291(.An(mai_mai_n318_), .B(mai_mai_n319_), .Y(mai_mai_n320_));
  NOi32      m0292(.An(d), .Bn(a), .C(c), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n321_), .B(mai_mai_n146_), .Y(mai_mai_n322_));
  NO2        m0294(.A(mai_mai_n320_), .B(mai_mai_n316_), .Y(mai_mai_n323_));
  NO2        m0295(.A(mai_mai_n319_), .B(mai_mai_n236_), .Y(mai_mai_n324_));
  NOi32      m0296(.An(f), .Bn(d), .C(c), .Y(mai_mai_n325_));
  AOI220     m0297(.A0(mai_mai_n325_), .A1(mai_mai_n244_), .B0(mai_mai_n324_), .B1(mai_mai_n174_), .Y(mai_mai_n326_));
  NA3        m0298(.A(mai_mai_n326_), .B(mai_mai_n323_), .C(mai_mai_n312_), .Y(mai_mai_n327_));
  INV        m0299(.A(e), .Y(mai_mai_n328_));
  NO2        m0300(.A(mai_mai_n1204_), .B(mai_mai_n1200_), .Y(mai_mai_n329_));
  AN2        m0301(.A(m), .B(e), .Y(mai_mai_n330_));
  INV        m0302(.A(mai_mai_n329_), .Y(mai_mai_n331_));
  NOi32      m0303(.An(h), .Bn(e), .C(m), .Y(mai_mai_n332_));
  NA3        m0304(.A(mai_mai_n332_), .B(mai_mai_n233_), .C(m), .Y(mai_mai_n333_));
  NOi21      m0305(.An(m), .B(h), .Y(mai_mai_n334_));
  NA3        m0306(.A(m), .B(mai_mai_n334_), .C(e), .Y(mai_mai_n335_));
  NA3        m0307(.A(mai_mai_n34_), .B(m), .C(e), .Y(mai_mai_n336_));
  NA3        m0308(.A(mai_mai_n321_), .B(mai_mai_n146_), .C(mai_mai_n62_), .Y(mai_mai_n337_));
  NAi31      m0309(.An(b), .B(c), .C(a), .Y(mai_mai_n338_));
  NO2        m0310(.A(mai_mai_n338_), .B(n), .Y(mai_mai_n339_));
  INV        m0311(.A(mai_mai_n327_), .Y(mai_mai_n340_));
  NO2        m0312(.A(mai_mai_n224_), .B(c), .Y(mai_mai_n341_));
  NOi21      m0313(.An(a), .B(n), .Y(mai_mai_n342_));
  NOi21      m0314(.An(d), .B(c), .Y(mai_mai_n343_));
  NA2        m0315(.A(mai_mai_n343_), .B(mai_mai_n342_), .Y(mai_mai_n344_));
  NA3        m0316(.A(m), .B(mai_mai_n334_), .C(mai_mai_n146_), .Y(mai_mai_n345_));
  NO2        m0317(.A(mai_mai_n345_), .B(mai_mai_n344_), .Y(mai_mai_n346_));
  INV        m0318(.A(mai_mai_n346_), .Y(mai_mai_n347_));
  OR2        m0319(.A(n), .B(m), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n348_), .B(mai_mai_n119_), .Y(mai_mai_n349_));
  NO2        m0321(.A(mai_mai_n147_), .B(mai_mai_n115_), .Y(mai_mai_n350_));
  OAI210     m0322(.A0(mai_mai_n349_), .A1(mai_mai_n140_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  NA3        m0323(.A(mai_mai_n87_), .B(mai_mai_n287_), .C(d), .Y(mai_mai_n352_));
  NO2        m0324(.A(mai_mai_n338_), .B(mai_mai_n39_), .Y(mai_mai_n353_));
  NAi21      m0325(.An(k), .B(j), .Y(mai_mai_n354_));
  NAi21      m0326(.An(e), .B(d), .Y(mai_mai_n355_));
  INV        m0327(.A(mai_mai_n355_), .Y(mai_mai_n356_));
  NO2        m0328(.A(mai_mai_n210_), .B(mai_mai_n172_), .Y(mai_mai_n357_));
  NA3        m0329(.A(mai_mai_n357_), .B(mai_mai_n356_), .C(mai_mai_n185_), .Y(mai_mai_n358_));
  NA3        m0330(.A(mai_mai_n358_), .B(mai_mai_n352_), .C(mai_mai_n351_), .Y(mai_mai_n359_));
  NO2        m0331(.A(mai_mai_n266_), .B(mai_mai_n172_), .Y(mai_mai_n360_));
  NA2        m0332(.A(mai_mai_n360_), .B(mai_mai_n356_), .Y(mai_mai_n361_));
  NOi31      m0333(.An(n), .B(m), .C(k), .Y(mai_mai_n362_));
  AOI220     m0334(.A0(mai_mai_n362_), .A1(mai_mai_n313_), .B0(mai_mai_n180_), .B1(mai_mai_n40_), .Y(mai_mai_n363_));
  NAi31      m0335(.An(m), .B(f), .C(c), .Y(mai_mai_n364_));
  NA2        m0336(.A(mai_mai_n361_), .B(mai_mai_n245_), .Y(mai_mai_n365_));
  NO2        m0337(.A(mai_mai_n365_), .B(mai_mai_n359_), .Y(mai_mai_n366_));
  NOi32      m0338(.An(c), .Bn(a), .C(b), .Y(mai_mai_n367_));
  NA2        m0339(.A(mai_mai_n367_), .B(mai_mai_n87_), .Y(mai_mai_n368_));
  AN2        m0340(.A(e), .B(d), .Y(mai_mai_n369_));
  NO2        m0341(.A(mai_mai_n115_), .B(mai_mai_n368_), .Y(mai_mai_n370_));
  NOi21      m0342(.An(a), .B(b), .Y(mai_mai_n371_));
  NA3        m0343(.A(e), .B(d), .C(c), .Y(mai_mai_n372_));
  BUFFER     m0344(.A(mai_mai_n372_), .Y(mai_mai_n373_));
  NO2        m0345(.A(mai_mai_n36_), .B(mai_mai_n373_), .Y(mai_mai_n374_));
  NO4        m0346(.A(mai_mai_n152_), .B(mai_mai_n78_), .C(mai_mai_n44_), .D(b), .Y(mai_mai_n375_));
  NA2        m0347(.A(mai_mai_n308_), .B(mai_mai_n120_), .Y(mai_mai_n376_));
  OR2        m0348(.A(k), .B(j), .Y(mai_mai_n377_));
  NA2        m0349(.A(l), .B(k), .Y(mai_mai_n378_));
  NA3        m0350(.A(mai_mai_n378_), .B(mai_mai_n377_), .C(mai_mai_n180_), .Y(mai_mai_n379_));
  NA3        m0351(.A(mai_mai_n227_), .B(mai_mai_n96_), .C(mai_mai_n94_), .Y(mai_mai_n380_));
  NA2        m0352(.A(mai_mai_n321_), .B(mai_mai_n87_), .Y(mai_mai_n381_));
  NO3        m0353(.A(mai_mai_n337_), .B(mai_mai_n69_), .C(m), .Y(mai_mai_n382_));
  NO2        m0354(.A(mai_mai_n382_), .B(mai_mai_n380_), .Y(mai_mai_n383_));
  NA2        m0355(.A(mai_mai_n383_), .B(mai_mai_n376_), .Y(mai_mai_n384_));
  NO4        m0356(.A(mai_mai_n384_), .B(mai_mai_n375_), .C(mai_mai_n374_), .D(mai_mai_n370_), .Y(mai_mai_n385_));
  NOi21      m0357(.An(d), .B(e), .Y(mai_mai_n386_));
  OAI210     m0358(.A0(j), .A1(mai_mai_n99_), .B0(mai_mai_n78_), .Y(mai_mai_n387_));
  NO2        m0359(.A(mai_mai_n322_), .B(mai_mai_n297_), .Y(mai_mai_n388_));
  NO2        m0360(.A(mai_mai_n388_), .B(mai_mai_n149_), .Y(mai_mai_n389_));
  NA2        m0361(.A(mai_mai_n389_), .B(mai_mai_n198_), .Y(mai_mai_n390_));
  OAI210     m0362(.A0(mai_mai_n95_), .A1(mai_mai_n93_), .B0(n), .Y(mai_mai_n391_));
  XO2        m0363(.A(i), .B(h), .Y(mai_mai_n392_));
  NA3        m0364(.A(mai_mai_n392_), .B(mai_mai_n126_), .C(n), .Y(mai_mai_n393_));
  NAi41      m0365(.An(mai_mai_n237_), .B(mai_mai_n393_), .C(mai_mai_n363_), .D(mai_mai_n310_), .Y(mai_mai_n394_));
  AN2        m0366(.A(mai_mai_n394_), .B(mai_mai_n1206_), .Y(mai_mai_n395_));
  NAi31      m0367(.An(c), .B(f), .C(d), .Y(mai_mai_n396_));
  AOI210     m0368(.A0(mai_mai_n228_), .A1(mai_mai_n160_), .B0(mai_mai_n396_), .Y(mai_mai_n397_));
  NOi21      m0369(.An(mai_mai_n60_), .B(mai_mai_n397_), .Y(mai_mai_n398_));
  NA3        m0370(.A(mai_mai_n306_), .B(m), .C(m), .Y(mai_mai_n399_));
  NA2        m0371(.A(mai_mai_n186_), .B(mai_mai_n83_), .Y(mai_mai_n400_));
  AOI210     m0372(.A0(mai_mai_n400_), .A1(mai_mai_n145_), .B0(mai_mai_n396_), .Y(mai_mai_n401_));
  NOi21      m0373(.An(mai_mai_n399_), .B(mai_mai_n401_), .Y(mai_mai_n402_));
  NA3        m0374(.A(mai_mai_n34_), .B(m), .C(f), .Y(mai_mai_n403_));
  NA3        m0375(.A(mai_mai_n234_), .B(mai_mai_n402_), .C(mai_mai_n398_), .Y(mai_mai_n404_));
  NO3        m0376(.A(mai_mai_n404_), .B(mai_mai_n395_), .C(mai_mai_n390_), .Y(mai_mai_n405_));
  NA4        m0377(.A(mai_mai_n405_), .B(mai_mai_n385_), .C(mai_mai_n366_), .D(mai_mai_n340_), .Y(mai11));
  NO2        m0378(.A(mai_mai_n50_), .B(f), .Y(mai_mai_n407_));
  NA3        m0379(.A(m), .B(k), .C(j), .Y(mai_mai_n408_));
  NA2        m0380(.A(m), .B(mai_mai_n407_), .Y(mai_mai_n409_));
  NOi32      m0381(.An(e), .Bn(b), .C(f), .Y(mai_mai_n410_));
  NA2        m0382(.A(mai_mai_n38_), .B(j), .Y(mai_mai_n411_));
  NO2        m0383(.A(mai_mai_n411_), .B(mai_mai_n239_), .Y(mai_mai_n412_));
  NAi31      m0384(.An(d), .B(e), .C(a), .Y(mai_mai_n413_));
  NO2        m0385(.A(mai_mai_n413_), .B(n), .Y(mai_mai_n414_));
  AOI210     m0386(.A0(mai_mai_n414_), .A1(mai_mai_n77_), .B0(mai_mai_n412_), .Y(mai_mai_n415_));
  NAi41      m0387(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n416_));
  AN2        m0388(.A(mai_mai_n416_), .B(mai_mai_n296_), .Y(mai_mai_n417_));
  NA2        m0389(.A(j), .B(i), .Y(mai_mai_n418_));
  NAi31      m0390(.An(n), .B(m), .C(k), .Y(mai_mai_n419_));
  NO4        m0391(.A(n), .B(d), .C(mai_mai_n89_), .D(a), .Y(mai_mai_n420_));
  OR2        m0392(.A(n), .B(c), .Y(mai_mai_n421_));
  NO2        m0393(.A(mai_mai_n421_), .B(mai_mai_n116_), .Y(mai_mai_n422_));
  INV        m0394(.A(mai_mai_n422_), .Y(mai_mai_n423_));
  NOi32      m0395(.An(m), .Bn(f), .C(i), .Y(mai_mai_n424_));
  NO2        m0396(.A(mai_mai_n408_), .B(mai_mai_n423_), .Y(mai_mai_n425_));
  INV        m0397(.A(mai_mai_n425_), .Y(mai_mai_n426_));
  NA2        m0398(.A(mai_mai_n108_), .B(mai_mai_n33_), .Y(mai_mai_n427_));
  OAI220     m0399(.A0(mai_mai_n427_), .A1(m), .B0(mai_mai_n411_), .B1(mai_mai_n192_), .Y(mai_mai_n428_));
  NOi41      m0400(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n429_));
  NAi32      m0401(.An(e), .Bn(b), .C(c), .Y(mai_mai_n430_));
  OR2        m0402(.A(mai_mai_n430_), .B(mai_mai_n62_), .Y(mai_mai_n431_));
  AN2        m0403(.A(mai_mai_n270_), .B(mai_mai_n251_), .Y(mai_mai_n432_));
  NA2        m0404(.A(mai_mai_n432_), .B(mai_mai_n431_), .Y(mai_mai_n433_));
  AN2        m0405(.A(mai_mai_n429_), .B(mai_mai_n428_), .Y(mai_mai_n434_));
  NAi31      m0406(.An(d), .B(c), .C(a), .Y(mai_mai_n435_));
  NO2        m0407(.A(mai_mai_n435_), .B(n), .Y(mai_mai_n436_));
  NA3        m0408(.A(mai_mai_n436_), .B(m), .C(e), .Y(mai_mai_n437_));
  NO3        m0409(.A(i), .B(mai_mai_n39_), .C(mai_mai_n173_), .Y(mai_mai_n438_));
  NO2        m0410(.A(mai_mai_n189_), .B(mai_mai_n84_), .Y(mai_mai_n439_));
  NA2        m0411(.A(mai_mai_n438_), .B(mai_mai_n439_), .Y(mai_mai_n440_));
  NA2        m0412(.A(mai_mai_n440_), .B(mai_mai_n437_), .Y(mai_mai_n441_));
  NO2        m0413(.A(mai_mai_n224_), .B(n), .Y(mai_mai_n442_));
  NO2        m0414(.A(mai_mai_n339_), .B(mai_mai_n442_), .Y(mai_mai_n443_));
  NA2        m0415(.A(m), .B(f), .Y(mai_mai_n444_));
  NAi32      m0416(.An(d), .Bn(a), .C(b), .Y(mai_mai_n445_));
  NO2        m0417(.A(mai_mai_n445_), .B(mai_mai_n39_), .Y(mai_mai_n446_));
  NA2        m0418(.A(h), .B(f), .Y(mai_mai_n447_));
  NO2        m0419(.A(mai_mai_n447_), .B(mai_mai_n72_), .Y(mai_mai_n448_));
  NO3        m0420(.A(mai_mai_n141_), .B(mai_mai_n138_), .C(m), .Y(mai_mai_n449_));
  AOI210     m0421(.A0(mai_mai_n449_), .A1(c), .B0(mai_mai_n446_), .Y(mai_mai_n450_));
  OAI210     m0422(.A0(mai_mai_n444_), .A1(mai_mai_n443_), .B0(mai_mai_n450_), .Y(mai_mai_n451_));
  NO2        m0423(.A(mai_mai_n114_), .B(c), .Y(mai_mai_n452_));
  NA3        m0424(.A(mai_mai_n452_), .B(j), .C(mai_mai_n362_), .Y(mai_mai_n453_));
  NA3        m0425(.A(f), .B(d), .C(b), .Y(mai_mai_n454_));
  INV        m0426(.A(mai_mai_n453_), .Y(mai_mai_n455_));
  NO4        m0427(.A(mai_mai_n455_), .B(mai_mai_n451_), .C(mai_mai_n441_), .D(mai_mai_n434_), .Y(mai_mai_n456_));
  AN4        m0428(.A(mai_mai_n456_), .B(mai_mai_n426_), .C(mai_mai_n415_), .D(mai_mai_n409_), .Y(mai_mai_n457_));
  INV        m0429(.A(k), .Y(mai_mai_n458_));
  NA4        m0430(.A(mai_mai_n321_), .B(mai_mai_n334_), .C(mai_mai_n146_), .D(mai_mai_n87_), .Y(mai_mai_n459_));
  NAi32      m0431(.An(h), .Bn(f), .C(m), .Y(mai_mai_n460_));
  NAi41      m0432(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n461_));
  OAI210     m0433(.A0(mai_mai_n413_), .A1(n), .B0(mai_mai_n461_), .Y(mai_mai_n462_));
  NA2        m0434(.A(mai_mai_n462_), .B(m), .Y(mai_mai_n463_));
  NAi31      m0435(.An(h), .B(m), .C(f), .Y(mai_mai_n464_));
  OR3        m0436(.A(mai_mai_n464_), .B(mai_mai_n224_), .C(mai_mai_n39_), .Y(mai_mai_n465_));
  NA4        m0437(.A(mai_mai_n334_), .B(mai_mai_n91_), .C(mai_mai_n87_), .D(e), .Y(mai_mai_n466_));
  AN2        m0438(.A(mai_mai_n466_), .B(mai_mai_n465_), .Y(mai_mai_n467_));
  OA210      m0439(.A0(mai_mai_n463_), .A1(mai_mai_n460_), .B0(mai_mai_n467_), .Y(mai_mai_n468_));
  NO3        m0440(.A(mai_mai_n460_), .B(mai_mai_n50_), .C(mai_mai_n51_), .Y(mai_mai_n469_));
  NO4        m0441(.A(mai_mai_n464_), .B(mai_mai_n421_), .C(mai_mai_n116_), .D(mai_mai_n51_), .Y(mai_mai_n470_));
  OR2        m0442(.A(mai_mai_n470_), .B(mai_mai_n469_), .Y(mai_mai_n471_));
  NAi21      m0443(.An(mai_mai_n471_), .B(mai_mai_n468_), .Y(mai_mai_n472_));
  NAi31      m0444(.An(f), .B(h), .C(m), .Y(mai_mai_n473_));
  NOi32      m0445(.An(b), .Bn(a), .C(c), .Y(mai_mai_n474_));
  NOi32      m0446(.An(d), .Bn(a), .C(e), .Y(mai_mai_n475_));
  NA2        m0447(.A(mai_mai_n475_), .B(mai_mai_n87_), .Y(mai_mai_n476_));
  NO2        m0448(.A(n), .B(c), .Y(mai_mai_n477_));
  NA3        m0449(.A(mai_mai_n477_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n478_));
  NAi32      m0450(.An(n), .Bn(f), .C(m), .Y(mai_mai_n479_));
  NOi32      m0451(.An(e), .Bn(a), .C(d), .Y(mai_mai_n480_));
  INV        m0452(.A(mai_mai_n472_), .Y(mai_mai_n481_));
  NO3        m0453(.A(mai_mai_n249_), .B(mai_mai_n47_), .C(n), .Y(mai_mai_n482_));
  NA3        m0454(.A(mai_mai_n396_), .B(mai_mai_n137_), .C(mai_mai_n136_), .Y(mai_mai_n483_));
  NA2        m0455(.A(mai_mai_n364_), .B(mai_mai_n189_), .Y(mai_mai_n484_));
  OR2        m0456(.A(mai_mai_n484_), .B(mai_mai_n483_), .Y(mai_mai_n485_));
  NA2        m0457(.A(mai_mai_n52_), .B(mai_mai_n87_), .Y(mai_mai_n486_));
  NA2        m0458(.A(mai_mai_n485_), .B(mai_mai_n482_), .Y(mai_mai_n487_));
  NO2        m0459(.A(mai_mai_n487_), .B(mai_mai_n64_), .Y(mai_mai_n488_));
  NA3        m0460(.A(mai_mai_n429_), .B(mai_mai_n272_), .C(mai_mai_n38_), .Y(mai_mai_n489_));
  NOi32      m0461(.An(e), .Bn(c), .C(f), .Y(mai_mai_n490_));
  NOi21      m0462(.An(f), .B(m), .Y(mai_mai_n491_));
  NO2        m0463(.A(mai_mai_n491_), .B(mai_mai_n170_), .Y(mai_mai_n492_));
  AOI220     m0464(.A0(mai_mai_n492_), .A1(mai_mai_n318_), .B0(mai_mai_n490_), .B1(mai_mai_n140_), .Y(mai_mai_n493_));
  NA3        m0465(.A(mai_mai_n493_), .B(mai_mai_n489_), .C(mai_mai_n143_), .Y(mai_mai_n494_));
  AOI210     m0466(.A0(mai_mai_n417_), .A1(mai_mai_n322_), .B0(mai_mai_n238_), .Y(mai_mai_n495_));
  NAi21      m0467(.An(k), .B(h), .Y(mai_mai_n496_));
  NO2        m0468(.A(mai_mai_n496_), .B(f), .Y(mai_mai_n497_));
  NA2        m0469(.A(mai_mai_n497_), .B(j), .Y(mai_mai_n498_));
  OR2        m0470(.A(mai_mai_n498_), .B(mai_mai_n463_), .Y(mai_mai_n499_));
  NOi31      m0471(.An(m), .B(n), .C(k), .Y(mai_mai_n500_));
  NA2        m0472(.A(j), .B(mai_mai_n500_), .Y(mai_mai_n501_));
  AOI210     m0473(.A0(mai_mai_n322_), .A1(mai_mai_n296_), .B0(mai_mai_n238_), .Y(mai_mai_n502_));
  NAi21      m0474(.An(mai_mai_n501_), .B(mai_mai_n502_), .Y(mai_mai_n503_));
  NO2        m0475(.A(mai_mai_n224_), .B(mai_mai_n39_), .Y(mai_mai_n504_));
  INV        m0476(.A(mai_mai_n39_), .Y(mai_mai_n505_));
  NA2        m0477(.A(mai_mai_n504_), .B(mai_mai_n448_), .Y(mai_mai_n506_));
  NA3        m0478(.A(mai_mai_n506_), .B(mai_mai_n503_), .C(mai_mai_n499_), .Y(mai_mai_n507_));
  NA2        m0479(.A(mai_mai_n83_), .B(m), .Y(mai_mai_n508_));
  NO2        m0480(.A(mai_mai_n410_), .B(mai_mai_n287_), .Y(mai_mai_n509_));
  NO2        m0481(.A(mai_mai_n509_), .B(n), .Y(mai_mai_n510_));
  NAi31      m0482(.An(mai_mai_n508_), .B(mai_mai_n510_), .C(m), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n411_), .B(mai_mai_n141_), .Y(mai_mai_n512_));
  NA3        m0484(.A(mai_mai_n430_), .B(mai_mai_n219_), .C(mai_mai_n112_), .Y(mai_mai_n513_));
  NO3        m0485(.A(mai_mai_n319_), .B(m), .C(mai_mai_n64_), .Y(mai_mai_n514_));
  AOI210     m0486(.A0(mai_mai_n513_), .A1(mai_mai_n512_), .B0(mai_mai_n514_), .Y(mai_mai_n515_));
  OAI210     m0487(.A0(d), .A1(mai_mai_n98_), .B0(n), .Y(mai_mai_n516_));
  NA3        m0488(.A(mai_mai_n392_), .B(mai_mai_n126_), .C(mai_mai_n173_), .Y(mai_mai_n517_));
  AOI210     m0489(.A0(mai_mai_n516_), .A1(mai_mai_n191_), .B0(mai_mai_n517_), .Y(mai_mai_n518_));
  NAi31      m0490(.An(m), .B(n), .C(k), .Y(mai_mai_n519_));
  OR2        m0491(.A(mai_mai_n102_), .B(mai_mai_n47_), .Y(mai_mai_n520_));
  INV        m0492(.A(mai_mai_n207_), .Y(mai_mai_n521_));
  OAI210     m0493(.A0(mai_mai_n521_), .A1(mai_mai_n518_), .B0(j), .Y(mai_mai_n522_));
  NA3        m0494(.A(mai_mai_n522_), .B(mai_mai_n515_), .C(mai_mai_n511_), .Y(mai_mai_n523_));
  NO4        m0495(.A(mai_mai_n523_), .B(mai_mai_n507_), .C(mai_mai_n494_), .D(mai_mai_n488_), .Y(mai_mai_n524_));
  INV        m0496(.A(mai_mai_n306_), .Y(mai_mai_n525_));
  OR3        m0497(.A(m), .B(mai_mai_n224_), .C(n), .Y(mai_mai_n526_));
  NA3        m0498(.A(mai_mai_n332_), .B(mai_mai_n91_), .C(mai_mai_n62_), .Y(mai_mai_n527_));
  OAI210     m0499(.A0(n), .A1(mai_mai_n68_), .B0(mai_mai_n527_), .Y(mai_mai_n528_));
  NOi21      m0500(.An(mai_mai_n526_), .B(mai_mai_n528_), .Y(mai_mai_n529_));
  AOI210     m0501(.A0(mai_mai_n529_), .A1(mai_mai_n525_), .B0(mai_mai_n408_), .Y(mai_mai_n530_));
  NO3        m0502(.A(m), .B(mai_mai_n172_), .C(mai_mai_n44_), .Y(mai_mai_n531_));
  NO2        m0503(.A(mai_mai_n400_), .B(mai_mai_n64_), .Y(mai_mai_n532_));
  OAI210     m0504(.A0(mai_mai_n532_), .A1(mai_mai_n318_), .B0(mai_mai_n531_), .Y(mai_mai_n533_));
  OR2        m0505(.A(mai_mai_n50_), .B(mai_mai_n51_), .Y(mai_mai_n534_));
  NA2        m0506(.A(mai_mai_n474_), .B(mai_mai_n274_), .Y(mai_mai_n535_));
  OA220      m0507(.A0(mai_mai_n501_), .A1(mai_mai_n535_), .B0(mai_mai_n498_), .B1(mai_mai_n534_), .Y(mai_mai_n536_));
  AN2        m0508(.A(h), .B(f), .Y(mai_mai_n537_));
  NA2        m0509(.A(mai_mai_n537_), .B(mai_mai_n34_), .Y(mai_mai_n538_));
  NA2        m0510(.A(mai_mai_n75_), .B(mai_mai_n38_), .Y(mai_mai_n539_));
  NO2        m0511(.A(mai_mai_n538_), .B(mai_mai_n368_), .Y(mai_mai_n540_));
  AOI210     m0512(.A0(mai_mai_n445_), .A1(mai_mai_n338_), .B0(mai_mai_n39_), .Y(mai_mai_n541_));
  NA2        m0513(.A(mai_mai_n536_), .B(mai_mai_n533_), .Y(mai_mai_n542_));
  NO2        m0514(.A(mai_mai_n209_), .B(f), .Y(mai_mai_n543_));
  NO2        m0515(.A(mai_mai_n491_), .B(mai_mai_n47_), .Y(mai_mai_n544_));
  NO2        m0516(.A(mai_mai_n544_), .B(mai_mai_n543_), .Y(mai_mai_n545_));
  INV        m0517(.A(mai_mai_n260_), .Y(mai_mai_n546_));
  OA220      m0518(.A0(mai_mai_n99_), .A1(mai_mai_n427_), .B0(mai_mai_n286_), .B1(mai_mai_n85_), .Y(mai_mai_n547_));
  OAI210     m0519(.A0(mai_mai_n546_), .A1(mai_mai_n545_), .B0(mai_mai_n547_), .Y(mai_mai_n548_));
  NO3        m0520(.A(mai_mai_n325_), .B(mai_mai_n157_), .C(mai_mai_n156_), .Y(mai_mai_n549_));
  NA2        m0521(.A(mai_mai_n549_), .B(mai_mai_n189_), .Y(mai_mai_n550_));
  NA3        m0522(.A(mai_mai_n550_), .B(mai_mai_n211_), .C(j), .Y(mai_mai_n551_));
  NO3        m0523(.A(mai_mai_n364_), .B(mai_mai_n138_), .C(i), .Y(mai_mai_n552_));
  NA2        m0524(.A(mai_mai_n367_), .B(mai_mai_n62_), .Y(mai_mai_n553_));
  NA3        m0525(.A(mai_mai_n551_), .B(mai_mai_n399_), .C(mai_mai_n323_), .Y(mai_mai_n554_));
  NO4        m0526(.A(mai_mai_n554_), .B(mai_mai_n548_), .C(mai_mai_n542_), .D(mai_mai_n530_), .Y(mai_mai_n555_));
  NA4        m0527(.A(mai_mai_n555_), .B(mai_mai_n524_), .C(mai_mai_n481_), .D(mai_mai_n457_), .Y(mai08));
  NO2        m0528(.A(k), .B(h), .Y(mai_mai_n557_));
  AO210      m0529(.A0(mai_mai_n209_), .A1(mai_mai_n354_), .B0(mai_mai_n557_), .Y(mai_mai_n558_));
  NO2        m0530(.A(mai_mai_n558_), .B(mai_mai_n236_), .Y(mai_mai_n559_));
  NA2        m0531(.A(mai_mai_n490_), .B(mai_mai_n62_), .Y(mai_mai_n560_));
  NA2        m0532(.A(mai_mai_n560_), .B(mai_mai_n364_), .Y(mai_mai_n561_));
  AOI210     m0533(.A0(mai_mai_n561_), .A1(mai_mai_n559_), .B0(mai_mai_n382_), .Y(mai_mai_n562_));
  NA2        m0534(.A(mai_mai_n62_), .B(mai_mai_n84_), .Y(mai_mai_n563_));
  NO2        m0535(.A(mai_mai_n563_), .B(mai_mai_n45_), .Y(mai_mai_n564_));
  NA2        m0536(.A(mai_mai_n454_), .B(mai_mai_n191_), .Y(mai_mai_n565_));
  AOI220     m0537(.A0(mai_mai_n565_), .A1(mai_mai_n277_), .B0(m), .B1(mai_mai_n564_), .Y(mai_mai_n566_));
  AOI210     m0538(.A0(mai_mai_n454_), .A1(mai_mai_n122_), .B0(mai_mai_n62_), .Y(mai_mai_n567_));
  NA4        m0539(.A(mai_mai_n175_), .B(mai_mai_n108_), .C(mai_mai_n37_), .D(h), .Y(mai_mai_n568_));
  AN2        m0540(.A(l), .B(k), .Y(mai_mai_n569_));
  NA4        m0541(.A(mai_mai_n569_), .B(mai_mai_n83_), .C(mai_mai_n51_), .D(mai_mai_n173_), .Y(mai_mai_n570_));
  OAI210     m0542(.A0(mai_mai_n568_), .A1(m), .B0(mai_mai_n570_), .Y(mai_mai_n571_));
  NA2        m0543(.A(mai_mai_n571_), .B(mai_mai_n567_), .Y(mai_mai_n572_));
  NA4        m0544(.A(mai_mai_n572_), .B(mai_mai_n566_), .C(mai_mai_n562_), .D(mai_mai_n279_), .Y(mai_mai_n573_));
  NO4        m0545(.A(mai_mai_n138_), .B(mai_mai_n317_), .C(mai_mai_n86_), .D(m), .Y(mai_mai_n574_));
  NA2        m0546(.A(mai_mai_n574_), .B(mai_mai_n565_), .Y(mai_mai_n575_));
  NA2        m0547(.A(mai_mai_n492_), .B(mai_mai_n276_), .Y(mai_mai_n576_));
  NAi31      m0548(.An(mai_mai_n73_), .B(mai_mai_n576_), .C(mai_mai_n575_), .Y(mai_mai_n577_));
  NA2        m0549(.A(mai_mai_n430_), .B(mai_mai_n520_), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n378_), .B(mai_mai_n99_), .Y(mai_mai_n579_));
  NA2        m0551(.A(mai_mai_n579_), .B(mai_mai_n578_), .Y(mai_mai_n580_));
  NO3        m0552(.A(mai_mai_n249_), .B(m), .C(j), .Y(mai_mai_n581_));
  NAi21      m0553(.An(mai_mai_n581_), .B(mai_mai_n570_), .Y(mai_mai_n582_));
  NA2        m0554(.A(mai_mai_n558_), .B(mai_mai_n103_), .Y(mai_mai_n583_));
  AOI220     m0555(.A0(mai_mai_n583_), .A1(mai_mai_n324_), .B0(mai_mai_n582_), .B1(mai_mai_n54_), .Y(mai_mai_n584_));
  OAI210     m0556(.A0(mai_mai_n580_), .A1(mai_mai_n64_), .B0(mai_mai_n584_), .Y(mai_mai_n585_));
  NA3        m0557(.A(mai_mai_n550_), .B(mai_mai_n265_), .C(mai_mai_n309_), .Y(mai_mai_n586_));
  NA2        m0558(.A(mai_mai_n569_), .B(mai_mai_n180_), .Y(mai_mai_n587_));
  NO2        m0559(.A(mai_mai_n587_), .B(mai_mai_n259_), .Y(mai_mai_n588_));
  NA2        m0560(.A(mai_mai_n588_), .B(mai_mai_n543_), .Y(mai_mai_n589_));
  NA3        m0561(.A(m), .B(l), .C(k), .Y(mai_mai_n590_));
  AOI210     m0562(.A0(mai_mai_n527_), .A1(mai_mai_n526_), .B0(mai_mai_n590_), .Y(mai_mai_n591_));
  NA4        m0563(.A(mai_mai_n87_), .B(l), .C(k), .D(mai_mai_n64_), .Y(mai_mai_n592_));
  NA3        m0564(.A(mai_mai_n91_), .B(mai_mai_n330_), .C(i), .Y(mai_mai_n593_));
  NO2        m0565(.A(mai_mai_n593_), .B(mai_mai_n592_), .Y(mai_mai_n594_));
  NO2        m0566(.A(mai_mai_n594_), .B(mai_mai_n591_), .Y(mai_mai_n595_));
  NA3        m0567(.A(mai_mai_n595_), .B(mai_mai_n589_), .C(mai_mai_n586_), .Y(mai_mai_n596_));
  NO4        m0568(.A(mai_mai_n596_), .B(mai_mai_n585_), .C(mai_mai_n577_), .D(mai_mai_n573_), .Y(mai_mai_n597_));
  NA2        m0569(.A(mai_mai_n492_), .B(mai_mai_n318_), .Y(mai_mai_n598_));
  NOi31      m0570(.An(m), .B(h), .C(f), .Y(mai_mai_n599_));
  NA2        m0571(.A(mai_mai_n505_), .B(mai_mai_n599_), .Y(mai_mai_n600_));
  AOI210     m0572(.A0(mai_mai_n321_), .A1(mai_mai_n87_), .B0(mai_mai_n388_), .Y(mai_mai_n601_));
  NA4        m0573(.A(mai_mai_n601_), .B(mai_mai_n600_), .C(mai_mai_n598_), .D(mai_mai_n208_), .Y(mai_mai_n602_));
  NA2        m0574(.A(mai_mai_n569_), .B(mai_mai_n51_), .Y(mai_mai_n603_));
  NO4        m0575(.A(mai_mai_n549_), .B(mai_mai_n138_), .C(n), .D(i), .Y(mai_mai_n604_));
  NOi21      m0576(.An(h), .B(j), .Y(mai_mai_n605_));
  NA2        m0577(.A(mai_mai_n605_), .B(f), .Y(mai_mai_n606_));
  NO2        m0578(.A(mai_mai_n606_), .B(mai_mai_n202_), .Y(mai_mai_n607_));
  NO3        m0579(.A(mai_mai_n607_), .B(mai_mai_n604_), .C(mai_mai_n552_), .Y(mai_mai_n608_));
  OAI210     m0580(.A0(mai_mai_n608_), .A1(mai_mai_n603_), .B0(mai_mai_n467_), .Y(mai_mai_n609_));
  NO2        m0581(.A(mai_mai_n602_), .B(mai_mai_n609_), .Y(mai_mai_n610_));
  NO2        m0582(.A(j), .B(i), .Y(mai_mai_n611_));
  NA3        m0583(.A(mai_mai_n611_), .B(mai_mai_n58_), .C(l), .Y(mai_mai_n612_));
  NA2        m0584(.A(mai_mai_n611_), .B(mai_mai_n32_), .Y(mai_mai_n613_));
  NA2        m0585(.A(e), .B(mai_mai_n91_), .Y(mai_mai_n614_));
  OA220      m0586(.A0(mai_mai_n614_), .A1(mai_mai_n613_), .B0(mai_mai_n612_), .B1(mai_mai_n463_), .Y(mai_mai_n615_));
  NO3        m0587(.A(mai_mai_n118_), .B(mai_mai_n39_), .C(mai_mai_n84_), .Y(mai_mai_n616_));
  NO3        m0588(.A(mai_mai_n421_), .B(mai_mai_n116_), .C(mai_mai_n51_), .Y(mai_mai_n617_));
  NA2        m0589(.A(k), .B(j), .Y(mai_mai_n618_));
  NO3        m0590(.A(mai_mai_n236_), .B(mai_mai_n618_), .C(mai_mai_n35_), .Y(mai_mai_n619_));
  AOI210     m0591(.A0(mai_mai_n410_), .A1(n), .B0(mai_mai_n429_), .Y(mai_mai_n620_));
  NA2        m0592(.A(mai_mai_n620_), .B(mai_mai_n432_), .Y(mai_mai_n621_));
  AN3        m0593(.A(mai_mai_n621_), .B(mai_mai_n619_), .C(mai_mai_n74_), .Y(mai_mai_n622_));
  NO3        m0594(.A(mai_mai_n138_), .B(mai_mai_n317_), .C(mai_mai_n86_), .Y(mai_mai_n623_));
  AOI220     m0595(.A0(mai_mai_n623_), .A1(mai_mai_n203_), .B0(mai_mai_n484_), .B1(mai_mai_n244_), .Y(mai_mai_n624_));
  NA2        m0596(.A(mai_mai_n70_), .B(mai_mai_n62_), .Y(mai_mai_n625_));
  NA2        m0597(.A(mai_mai_n625_), .B(mai_mai_n624_), .Y(mai_mai_n626_));
  NO2        m0598(.A(mai_mai_n236_), .B(mai_mai_n103_), .Y(mai_mai_n627_));
  AOI220     m0599(.A0(mai_mai_n627_), .A1(mai_mai_n492_), .B0(mai_mai_n581_), .B1(mai_mai_n567_), .Y(mai_mai_n628_));
  NO2        m0600(.A(mai_mai_n590_), .B(mai_mai_n68_), .Y(mai_mai_n629_));
  NA2        m0601(.A(mai_mai_n629_), .B(mai_mai_n462_), .Y(mai_mai_n630_));
  NA2        m0602(.A(mai_mai_n1205_), .B(mai_mai_n541_), .Y(mai_mai_n631_));
  NA3        m0603(.A(mai_mai_n631_), .B(mai_mai_n630_), .C(mai_mai_n628_), .Y(mai_mai_n632_));
  OR3        m0604(.A(mai_mai_n632_), .B(mai_mai_n626_), .C(mai_mai_n622_), .Y(mai_mai_n633_));
  NA3        m0605(.A(mai_mai_n620_), .B(mai_mai_n432_), .C(mai_mai_n431_), .Y(mai_mai_n634_));
  NA4        m0606(.A(mai_mai_n634_), .B(mai_mai_n175_), .C(mai_mai_n354_), .D(mai_mai_n33_), .Y(mai_mai_n635_));
  NO3        m0607(.A(mai_mai_n378_), .B(j), .C(f), .Y(mai_mai_n636_));
  NO2        m0608(.A(mai_mai_n568_), .B(mai_mai_n560_), .Y(mai_mai_n637_));
  INV        m0609(.A(mai_mai_n637_), .Y(mai_mai_n638_));
  NA3        m0610(.A(mai_mai_n424_), .B(mai_mai_n233_), .C(h), .Y(mai_mai_n639_));
  NOi21      m0611(.An(mai_mai_n541_), .B(mai_mai_n639_), .Y(mai_mai_n640_));
  INV        m0612(.A(mai_mai_n69_), .Y(mai_mai_n641_));
  NO2        m0613(.A(mai_mai_n639_), .B(mai_mai_n478_), .Y(mai_mai_n642_));
  AOI210     m0614(.A0(mai_mai_n641_), .A1(mai_mai_n510_), .B0(mai_mai_n642_), .Y(mai_mai_n643_));
  NA2        m0615(.A(mai_mai_n638_), .B(mai_mai_n635_), .Y(mai_mai_n644_));
  NO2        m0616(.A(n), .B(mai_mai_n51_), .Y(mai_mai_n645_));
  AOI210     m0617(.A0(mai_mai_n636_), .A1(mai_mai_n645_), .B0(mai_mai_n267_), .Y(mai_mai_n646_));
  OAI210     m0618(.A0(mai_mai_n590_), .A1(m), .B0(mai_mai_n403_), .Y(mai_mai_n647_));
  NA3        m0619(.A(mai_mai_n206_), .B(mai_mai_n46_), .C(b), .Y(mai_mai_n648_));
  AOI220     m0620(.A0(mai_mai_n477_), .A1(mai_mai_n29_), .B0(mai_mai_n367_), .B1(mai_mai_n62_), .Y(mai_mai_n649_));
  NA2        m0621(.A(mai_mai_n649_), .B(mai_mai_n648_), .Y(mai_mai_n650_));
  NO2        m0622(.A(mai_mai_n639_), .B(mai_mai_n381_), .Y(mai_mai_n651_));
  AOI210     m0623(.A0(mai_mai_n650_), .A1(mai_mai_n647_), .B0(mai_mai_n651_), .Y(mai_mai_n652_));
  NA3        m0624(.A(mai_mai_n652_), .B(mai_mai_n646_), .C(mai_mai_n1201_), .Y(mai_mai_n653_));
  NOi41      m0625(.An(mai_mai_n615_), .B(mai_mai_n653_), .C(mai_mai_n644_), .D(mai_mai_n633_), .Y(mai_mai_n654_));
  OR2        m0626(.A(mai_mai_n568_), .B(mai_mai_n191_), .Y(mai_mai_n655_));
  NO3        m0627(.A(mai_mai_n273_), .B(mai_mai_n238_), .C(mai_mai_n86_), .Y(mai_mai_n656_));
  NA2        m0628(.A(mai_mai_n656_), .B(mai_mai_n621_), .Y(mai_mai_n657_));
  NO2        m0629(.A(mai_mai_n613_), .B(mai_mai_n224_), .Y(mai_mai_n658_));
  NA3        m0630(.A(mai_mai_n657_), .B(mai_mai_n655_), .C(mai_mai_n326_), .Y(mai_mai_n659_));
  NOi31      m0631(.An(b), .B(d), .C(a), .Y(mai_mai_n660_));
  NO2        m0632(.A(mai_mai_n660_), .B(mai_mai_n475_), .Y(mai_mai_n661_));
  NO2        m0633(.A(mai_mai_n661_), .B(n), .Y(mai_mai_n662_));
  NOi21      m0634(.An(mai_mai_n649_), .B(mai_mai_n662_), .Y(mai_mai_n663_));
  NO2        m0635(.A(mai_mai_n663_), .B(mai_mai_n69_), .Y(mai_mai_n664_));
  NO2        m0636(.A(mai_mai_n430_), .B(mai_mai_n62_), .Y(mai_mai_n665_));
  NO3        m0637(.A(mai_mai_n491_), .B(mai_mai_n259_), .C(mai_mai_n90_), .Y(mai_mai_n666_));
  NOi21      m0638(.An(mai_mai_n666_), .B(mai_mai_n127_), .Y(mai_mai_n667_));
  AOI210     m0639(.A0(mai_mai_n656_), .A1(mai_mai_n665_), .B0(mai_mai_n667_), .Y(mai_mai_n668_));
  OAI210     m0640(.A0(mai_mai_n568_), .A1(mai_mai_n319_), .B0(mai_mai_n668_), .Y(mai_mai_n669_));
  NO2        m0641(.A(mai_mai_n549_), .B(n), .Y(mai_mai_n670_));
  AOI220     m0642(.A0(mai_mai_n627_), .A1(mai_mai_n531_), .B0(mai_mai_n670_), .B1(mai_mai_n559_), .Y(mai_mai_n671_));
  NA2        m0643(.A(mai_mai_n91_), .B(mai_mai_n62_), .Y(mai_mai_n672_));
  AOI210     m0644(.A0(mai_mai_n336_), .A1(mai_mai_n333_), .B0(mai_mai_n672_), .Y(mai_mai_n673_));
  NA2        m0645(.A(mai_mai_n588_), .B(mai_mai_n33_), .Y(mai_mai_n674_));
  NAi21      m0646(.An(mai_mai_n592_), .B(mai_mai_n341_), .Y(mai_mai_n675_));
  NA2        m0647(.A(mai_mai_n574_), .B(mai_mai_n278_), .Y(mai_mai_n676_));
  NO2        m0648(.A(mai_mai_n470_), .B(mai_mai_n469_), .Y(mai_mai_n677_));
  AN3        m0649(.A(mai_mai_n677_), .B(mai_mai_n676_), .C(mai_mai_n675_), .Y(mai_mai_n678_));
  NAi41      m0650(.An(mai_mai_n673_), .B(mai_mai_n678_), .C(mai_mai_n674_), .D(mai_mai_n671_), .Y(mai_mai_n679_));
  NO4        m0651(.A(mai_mai_n679_), .B(mai_mai_n669_), .C(mai_mai_n664_), .D(mai_mai_n659_), .Y(mai_mai_n680_));
  NA4        m0652(.A(mai_mai_n680_), .B(mai_mai_n654_), .C(mai_mai_n610_), .D(mai_mai_n597_), .Y(mai09));
  INV        m0653(.A(mai_mai_n92_), .Y(mai_mai_n682_));
  NA2        m0654(.A(mai_mai_n349_), .B(e), .Y(mai_mai_n683_));
  NO2        m0655(.A(mai_mai_n683_), .B(mai_mai_n396_), .Y(mai_mai_n684_));
  AOI210     m0656(.A0(e), .A1(mai_mai_n682_), .B0(mai_mai_n684_), .Y(mai_mai_n685_));
  OA210      m0657(.A0(m), .A1(m), .B0(mai_mai_n662_), .Y(mai_mai_n686_));
  INV        m0658(.A(mai_mai_n270_), .Y(mai_mai_n687_));
  NO2        m0659(.A(mai_mai_n95_), .B(mai_mai_n93_), .Y(mai_mai_n688_));
  NOi31      m0660(.An(k), .B(m), .C(l), .Y(mai_mai_n689_));
  NO2        m0661(.A(mai_mai_n272_), .B(mai_mai_n689_), .Y(mai_mai_n690_));
  AOI210     m0662(.A0(mai_mai_n690_), .A1(mai_mai_n688_), .B0(mai_mai_n473_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n691_), .B(mai_mai_n687_), .Y(mai_mai_n692_));
  NA2        m0664(.A(mai_mai_n133_), .B(mai_mai_n88_), .Y(mai_mai_n693_));
  NA3        m0665(.A(mai_mai_n693_), .B(mai_mai_n558_), .C(mai_mai_n103_), .Y(mai_mai_n694_));
  NA3        m0666(.A(mai_mai_n694_), .B(mai_mai_n154_), .C(mai_mai_n30_), .Y(mai_mai_n695_));
  NA4        m0667(.A(mai_mai_n695_), .B(mai_mai_n692_), .C(mai_mai_n493_), .D(mai_mai_n60_), .Y(mai_mai_n696_));
  NO2        m0668(.A(mai_mai_n460_), .B(j), .Y(mai_mai_n697_));
  NA2        m0669(.A(mai_mai_n697_), .B(mai_mai_n154_), .Y(mai_mai_n698_));
  NOi21      m0670(.An(f), .B(d), .Y(mai_mai_n699_));
  NA2        m0671(.A(mai_mai_n699_), .B(m), .Y(mai_mai_n700_));
  INV        m0672(.A(mai_mai_n700_), .Y(mai_mai_n701_));
  NA2        m0673(.A(mai_mai_n701_), .B(mai_mai_n422_), .Y(mai_mai_n702_));
  NA3        m0674(.A(mai_mai_n371_), .B(d), .C(mai_mai_n62_), .Y(mai_mai_n703_));
  NO2        m0675(.A(mai_mai_n232_), .B(mai_mai_n44_), .Y(mai_mai_n704_));
  NAi31      m0676(.An(mai_mai_n380_), .B(mai_mai_n702_), .C(mai_mai_n698_), .Y(mai_mai_n705_));
  NO4        m0677(.A(mai_mai_n491_), .B(mai_mai_n99_), .C(mai_mai_n259_), .D(mai_mai_n119_), .Y(mai_mai_n706_));
  NO2        m0678(.A(mai_mai_n519_), .B(mai_mai_n259_), .Y(mai_mai_n707_));
  AN2        m0679(.A(mai_mai_n707_), .B(mai_mai_n543_), .Y(mai_mai_n708_));
  NO3        m0680(.A(mai_mai_n708_), .B(mai_mai_n706_), .C(mai_mai_n193_), .Y(mai_mai_n709_));
  NA2        m0681(.A(mai_mai_n475_), .B(mai_mai_n62_), .Y(mai_mai_n710_));
  NA3        m0682(.A(mai_mai_n126_), .B(mai_mai_n83_), .C(mai_mai_n82_), .Y(mai_mai_n711_));
  NO2        m0683(.A(mai_mai_n270_), .B(mai_mai_n711_), .Y(mai_mai_n712_));
  NOi21      m0684(.An(mai_mai_n182_), .B(mai_mai_n712_), .Y(mai_mai_n713_));
  NA2        m0685(.A(c), .B(mai_mai_n89_), .Y(mai_mai_n714_));
  INV        m0686(.A(mai_mai_n714_), .Y(mai_mai_n715_));
  NA3        m0687(.A(mai_mai_n715_), .B(mai_mai_n394_), .C(f), .Y(mai_mai_n716_));
  OR2        m0688(.A(m), .B(mai_mai_n419_), .Y(mai_mai_n717_));
  INV        m0689(.A(mai_mai_n717_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n661_), .B(mai_mai_n85_), .Y(mai_mai_n719_));
  NA2        m0691(.A(mai_mai_n719_), .B(mai_mai_n718_), .Y(mai_mai_n720_));
  NA4        m0692(.A(mai_mai_n720_), .B(mai_mai_n716_), .C(mai_mai_n713_), .D(mai_mai_n709_), .Y(mai_mai_n721_));
  NO4        m0693(.A(mai_mai_n721_), .B(mai_mai_n705_), .C(mai_mai_n696_), .D(mai_mai_n686_), .Y(mai_mai_n722_));
  OR2        m0694(.A(mai_mai_n703_), .B(mai_mai_n51_), .Y(mai_mai_n723_));
  INV        m0695(.A(mai_mai_n723_), .Y(mai_mai_n724_));
  NO2        m0696(.A(mai_mai_n103_), .B(mai_mai_n99_), .Y(mai_mai_n725_));
  NO2        m0697(.A(mai_mai_n189_), .B(mai_mai_n183_), .Y(mai_mai_n726_));
  AOI220     m0698(.A0(mai_mai_n726_), .A1(mai_mai_n186_), .B0(mai_mai_n241_), .B1(mai_mai_n725_), .Y(mai_mai_n727_));
  INV        m0699(.A(mai_mai_n727_), .Y(mai_mai_n728_));
  NA2        m0700(.A(e), .B(d), .Y(mai_mai_n729_));
  OAI220     m0701(.A0(mai_mai_n729_), .A1(c), .B0(mai_mai_n254_), .B1(d), .Y(mai_mai_n730_));
  NA3        m0702(.A(mai_mai_n730_), .B(mai_mai_n357_), .C(mai_mai_n392_), .Y(mai_mai_n731_));
  AOI210     m0703(.A0(mai_mai_n400_), .A1(mai_mai_n145_), .B0(mai_mai_n189_), .Y(mai_mai_n732_));
  AOI210     m0704(.A0(mai_mai_n492_), .A1(mai_mai_n276_), .B0(mai_mai_n732_), .Y(mai_mai_n733_));
  NA3        m0705(.A(mai_mai_n132_), .B(mai_mai_n63_), .C(mai_mai_n33_), .Y(mai_mai_n734_));
  NA3        m0706(.A(mai_mai_n734_), .B(mai_mai_n733_), .C(mai_mai_n731_), .Y(mai_mai_n735_));
  NO3        m0707(.A(mai_mai_n735_), .B(mai_mai_n728_), .C(mai_mai_n724_), .Y(mai_mai_n736_));
  NA2        m0708(.A(mai_mai_n687_), .B(mai_mai_n30_), .Y(mai_mai_n737_));
  AO210      m0709(.A0(mai_mai_n737_), .A1(mai_mai_n560_), .B0(mai_mai_n176_), .Y(mai_mai_n738_));
  OAI220     m0710(.A0(mai_mai_n491_), .A1(mai_mai_n47_), .B0(mai_mai_n238_), .B1(j), .Y(mai_mai_n739_));
  AOI220     m0711(.A0(mai_mai_n739_), .A1(mai_mai_n707_), .B0(mai_mai_n482_), .B1(mai_mai_n490_), .Y(mai_mai_n740_));
  OAI210     m0712(.A0(mai_mai_n683_), .A1(mai_mai_n136_), .B0(mai_mai_n740_), .Y(mai_mai_n741_));
  INV        m0713(.A(mai_mai_n741_), .Y(mai_mai_n742_));
  AO220      m0714(.A0(mai_mai_n357_), .A1(mai_mai_n605_), .B0(mai_mai_n140_), .B1(f), .Y(mai_mai_n743_));
  OAI210     m0715(.A0(mai_mai_n743_), .A1(mai_mai_n360_), .B0(mai_mai_n730_), .Y(mai_mai_n744_));
  INV        m0716(.A(mai_mai_n49_), .Y(mai_mai_n745_));
  OAI210     m0717(.A0(m), .A1(mai_mai_n745_), .B0(mai_mai_n564_), .Y(mai_mai_n746_));
  AN4        m0718(.A(mai_mai_n746_), .B(mai_mai_n744_), .C(mai_mai_n742_), .D(mai_mai_n738_), .Y(mai_mai_n747_));
  NA4        m0719(.A(mai_mai_n747_), .B(mai_mai_n736_), .C(mai_mai_n722_), .D(mai_mai_n685_), .Y(mai12));
  NO2        m0720(.A(mai_mai_n355_), .B(c), .Y(mai_mai_n749_));
  NO3        m0721(.A(mai_mai_n348_), .B(mai_mai_n209_), .C(mai_mai_n173_), .Y(mai_mai_n750_));
  NA2        m0722(.A(mai_mai_n750_), .B(mai_mai_n749_), .Y(mai_mai_n751_));
  NA2        m0723(.A(mai_mai_n422_), .B(mai_mai_n745_), .Y(mai_mai_n752_));
  NO2        m0724(.A(mai_mai_n355_), .B(mai_mai_n89_), .Y(mai_mai_n753_));
  NO2        m0725(.A(m), .B(mai_mai_n303_), .Y(mai_mai_n754_));
  NA3        m0726(.A(mai_mai_n752_), .B(mai_mai_n751_), .C(mai_mai_n347_), .Y(mai_mai_n755_));
  AOI210     m0727(.A0(mai_mai_n192_), .A1(mai_mai_n269_), .B0(mai_mai_n165_), .Y(mai_mai_n756_));
  OAI210     m0728(.A0(mai_mai_n314_), .A1(mai_mai_n1213_), .B0(mai_mai_n325_), .Y(mai_mai_n757_));
  NO2        m0729(.A(mai_mai_n508_), .B(f), .Y(mai_mai_n758_));
  INV        m0730(.A(mai_mai_n464_), .Y(mai_mai_n759_));
  NA2        m0731(.A(mai_mai_n759_), .B(mai_mai_n442_), .Y(mai_mai_n760_));
  NO2        m0732(.A(mai_mai_n118_), .B(mai_mai_n196_), .Y(mai_mai_n761_));
  NA2        m0733(.A(mai_mai_n760_), .B(mai_mai_n757_), .Y(mai_mai_n762_));
  NO3        m0734(.A(mai_mai_n99_), .B(mai_mai_n119_), .C(mai_mai_n173_), .Y(mai_mai_n763_));
  INV        m0735(.A(mai_mai_n763_), .Y(mai_mai_n764_));
  NA4        m0736(.A(mai_mai_n349_), .B(mai_mai_n343_), .C(mai_mai_n146_), .D(m), .Y(mai_mai_n765_));
  NA2        m0737(.A(mai_mai_n765_), .B(mai_mai_n764_), .Y(mai_mai_n766_));
  NO2        m0738(.A(mai_mai_n529_), .B(mai_mai_n69_), .Y(mai_mai_n767_));
  NO4        m0739(.A(mai_mai_n767_), .B(mai_mai_n766_), .C(mai_mai_n762_), .D(mai_mai_n755_), .Y(mai_mai_n768_));
  NA2        m0740(.A(mai_mai_n430_), .B(mai_mai_n112_), .Y(mai_mai_n769_));
  NOi21      m0741(.An(mai_mai_n33_), .B(mai_mai_n519_), .Y(mai_mai_n770_));
  NA2        m0742(.A(mai_mai_n770_), .B(mai_mai_n769_), .Y(mai_mai_n771_));
  INV        m0743(.A(mai_mai_n771_), .Y(mai_mai_n772_));
  NO3        m0744(.A(mai_mai_n672_), .B(mai_mai_n66_), .C(mai_mai_n328_), .Y(mai_mai_n773_));
  NO2        m0745(.A(mai_mai_n391_), .B(mai_mai_n238_), .Y(mai_mai_n774_));
  INV        m0746(.A(mai_mai_n291_), .Y(mai_mai_n775_));
  NO4        m0747(.A(mai_mai_n775_), .B(mai_mai_n774_), .C(mai_mai_n773_), .D(mai_mai_n772_), .Y(mai_mai_n776_));
  NA2        m0748(.A(mai_mai_n276_), .B(m), .Y(mai_mai_n777_));
  NA2        m0749(.A(mai_mai_n38_), .B(i), .Y(mai_mai_n778_));
  NO2        m0750(.A(mai_mai_n112_), .B(mai_mai_n62_), .Y(mai_mai_n779_));
  OR2        m0751(.A(mai_mai_n779_), .B(mai_mai_n429_), .Y(mai_mai_n780_));
  NA2        m0752(.A(mai_mai_n430_), .B(mai_mai_n307_), .Y(mai_mai_n781_));
  AOI210     m0753(.A0(mai_mai_n781_), .A1(n), .B0(mai_mai_n780_), .Y(mai_mai_n782_));
  OAI220     m0754(.A0(mai_mai_n782_), .A1(mai_mai_n777_), .B0(mai_mai_n1200_), .B1(mai_mai_n264_), .Y(mai_mai_n783_));
  NO2        m0755(.A(m), .B(j), .Y(mai_mai_n784_));
  INV        m0756(.A(mai_mai_n1208_), .Y(mai_mai_n785_));
  OAI220     m0757(.A0(mai_mai_n785_), .A1(mai_mai_n784_), .B0(mai_mai_n541_), .B1(mai_mai_n617_), .Y(mai_mai_n786_));
  NA2        m0758(.A(mai_mai_n480_), .B(mai_mai_n87_), .Y(mai_mai_n787_));
  NA3        m0759(.A(j), .B(mai_mai_n58_), .C(i), .Y(mai_mai_n788_));
  OR2        m0760(.A(mai_mai_n788_), .B(mai_mai_n787_), .Y(mai_mai_n789_));
  NO2        m0761(.A(mai_mai_n1214_), .B(m), .Y(mai_mai_n790_));
  NA2        m0762(.A(mai_mai_n790_), .B(mai_mai_n255_), .Y(mai_mai_n791_));
  NA2        m0763(.A(mai_mai_n553_), .B(mai_mai_n710_), .Y(mai_mai_n792_));
  NA2        m0764(.A(i), .B(mai_mai_n55_), .Y(mai_mai_n793_));
  NA2        m0765(.A(mai_mai_n793_), .B(mai_mai_n788_), .Y(mai_mai_n794_));
  AOI220     m0766(.A0(mai_mai_n794_), .A1(mai_mai_n215_), .B0(mai_mai_n65_), .B1(mai_mai_n792_), .Y(mai_mai_n795_));
  NA4        m0767(.A(mai_mai_n795_), .B(mai_mai_n791_), .C(mai_mai_n789_), .D(mai_mai_n786_), .Y(mai_mai_n796_));
  NA2        m0768(.A(mai_mai_n758_), .B(mai_mai_n1215_), .Y(mai_mai_n797_));
  NA2        m0769(.A(mai_mai_n528_), .B(mai_mai_n65_), .Y(mai_mai_n798_));
  NO2        m0770(.A(mai_mai_n363_), .B(mai_mai_n173_), .Y(mai_mai_n799_));
  NA2        m0771(.A(mai_mai_n799_), .B(mai_mai_n308_), .Y(mai_mai_n800_));
  AOI220     m0772(.A0(mai_mai_n754_), .A1(mai_mai_n761_), .B0(mai_mai_n462_), .B1(mai_mai_n67_), .Y(mai_mai_n801_));
  NA4        m0773(.A(mai_mai_n801_), .B(mai_mai_n800_), .C(mai_mai_n798_), .D(mai_mai_n797_), .Y(mai_mai_n802_));
  OAI210     m0774(.A0(mai_mai_n65_), .A1(mai_mai_n759_), .B0(mai_mai_n420_), .Y(mai_mai_n803_));
  NO2        m0775(.A(mai_mai_n335_), .B(mai_mai_n672_), .Y(mai_mai_n804_));
  INV        m0776(.A(mai_mai_n804_), .Y(mai_mai_n805_));
  NA2        m0777(.A(mai_mai_n790_), .B(mai_mai_n753_), .Y(mai_mai_n806_));
  NO2        m0778(.A(mai_mai_n1198_), .B(mai_mai_n39_), .Y(mai_mai_n807_));
  AOI220     m0779(.A0(mai_mai_n807_), .A1(mai_mai_n495_), .B0(mai_mai_n512_), .B1(mai_mai_n410_), .Y(mai_mai_n808_));
  NA4        m0780(.A(mai_mai_n808_), .B(mai_mai_n806_), .C(mai_mai_n805_), .D(mai_mai_n803_), .Y(mai_mai_n809_));
  NO4        m0781(.A(mai_mai_n809_), .B(mai_mai_n802_), .C(mai_mai_n796_), .D(mai_mai_n783_), .Y(mai_mai_n810_));
  NAi31      m0782(.An(mai_mai_n109_), .B(e), .C(n), .Y(mai_mai_n811_));
  NO3        m0783(.A(mai_mai_n93_), .B(mai_mai_n272_), .C(mai_mai_n689_), .Y(mai_mai_n812_));
  NO2        m0784(.A(mai_mai_n812_), .B(mai_mai_n811_), .Y(mai_mai_n813_));
  NO3        m0785(.A(h), .B(mai_mai_n109_), .C(mai_mai_n328_), .Y(mai_mai_n814_));
  AOI210     m0786(.A0(mai_mai_n814_), .A1(mai_mai_n387_), .B0(mai_mai_n813_), .Y(mai_mai_n815_));
  NA2        m0787(.A(mai_mai_n382_), .B(i), .Y(mai_mai_n816_));
  NA2        m0788(.A(mai_mai_n816_), .B(mai_mai_n815_), .Y(mai_mai_n817_));
  NA2        m0789(.A(mai_mai_n189_), .B(mai_mai_n137_), .Y(mai_mai_n818_));
  NOi31      m0790(.An(mai_mai_n818_), .B(mai_mai_n348_), .C(mai_mai_n173_), .Y(mai_mai_n819_));
  NAi21      m0791(.An(mai_mai_n430_), .B(mai_mai_n799_), .Y(mai_mai_n820_));
  NA2        m0792(.A(mai_mai_n375_), .B(m), .Y(mai_mai_n821_));
  NA2        m0793(.A(mai_mai_n821_), .B(mai_mai_n820_), .Y(mai_mai_n822_));
  NO2        m0794(.A(mai_mai_n1208_), .B(mai_mai_n476_), .Y(mai_mai_n823_));
  NA2        m0795(.A(mai_mai_n756_), .B(mai_mai_n749_), .Y(mai_mai_n824_));
  NO3        m0796(.A(mai_mai_n421_), .B(mai_mai_n116_), .C(mai_mai_n172_), .Y(mai_mai_n825_));
  OAI210     m0797(.A0(mai_mai_n825_), .A1(mai_mai_n407_), .B0(mai_mai_n304_), .Y(mai_mai_n826_));
  OAI220     m0798(.A0(mai_mai_n754_), .A1(mai_mai_n759_), .B0(mai_mai_n422_), .B1(mai_mai_n339_), .Y(mai_mai_n827_));
  NA4        m0799(.A(mai_mai_n827_), .B(mai_mai_n826_), .C(mai_mai_n824_), .D(mai_mai_n489_), .Y(mai_mai_n828_));
  AOI210     m0800(.A0(mai_mai_n306_), .A1(mai_mai_n304_), .B0(mai_mai_n263_), .Y(mai_mai_n829_));
  NA2        m0801(.A(mai_mai_n829_), .B(mai_mai_n220_), .Y(mai_mai_n830_));
  OR3        m0802(.A(mai_mai_n830_), .B(mai_mai_n828_), .C(mai_mai_n823_), .Y(mai_mai_n831_));
  NO4        m0803(.A(mai_mai_n831_), .B(mai_mai_n822_), .C(mai_mai_n819_), .D(mai_mai_n817_), .Y(mai_mai_n832_));
  NA4        m0804(.A(mai_mai_n832_), .B(mai_mai_n810_), .C(mai_mai_n776_), .D(mai_mai_n768_), .Y(mai13));
  NA3        m0805(.A(mai_mai_n206_), .B(b), .C(m), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n386_), .B(f), .Y(mai_mai_n835_));
  NO4        m0807(.A(mai_mai_n835_), .B(mai_mai_n834_), .C(j), .D(k), .Y(mai_mai_n836_));
  NO4        m0808(.A(mai_mai_n48_), .B(mai_mai_n835_), .C(m), .D(a), .Y(mai_mai_n837_));
  NAi32      m0809(.An(d), .Bn(c), .C(e), .Y(mai_mai_n838_));
  NO4        m0810(.A(i), .B(mai_mai_n838_), .C(mai_mai_n464_), .D(mai_mai_n243_), .Y(mai_mai_n839_));
  NA2        m0811(.A(mai_mai_n330_), .B(mai_mai_n172_), .Y(mai_mai_n840_));
  NA2        m0812(.A(c), .B(mai_mai_n89_), .Y(mai_mai_n841_));
  NO3        m0813(.A(mai_mai_n841_), .B(mai_mai_n840_), .C(mai_mai_n141_), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n386_), .B(c), .Y(mai_mai_n843_));
  NO4        m0815(.A(i), .B(mai_mai_n460_), .C(mai_mai_n843_), .D(mai_mai_n243_), .Y(mai_mai_n844_));
  OR2        m0816(.A(mai_mai_n842_), .B(mai_mai_n844_), .Y(mai_mai_n845_));
  OR4        m0817(.A(mai_mai_n845_), .B(mai_mai_n839_), .C(mai_mai_n837_), .D(mai_mai_n836_), .Y(mai_mai_n846_));
  NAi32      m0818(.An(f), .Bn(e), .C(c), .Y(mai_mai_n847_));
  NO2        m0819(.A(mai_mai_n847_), .B(mai_mai_n114_), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n848_), .B(m), .Y(mai_mai_n849_));
  NO2        m0821(.A(mai_mai_n141_), .B(mai_mai_n849_), .Y(mai_mai_n850_));
  NO2        m0822(.A(mai_mai_n843_), .B(mai_mai_n243_), .Y(mai_mai_n851_));
  NO2        m0823(.A(j), .B(mai_mai_n37_), .Y(mai_mai_n852_));
  NA2        m0824(.A(mai_mai_n497_), .B(mai_mai_n852_), .Y(mai_mai_n853_));
  NOi21      m0825(.An(mai_mai_n851_), .B(mai_mai_n853_), .Y(mai_mai_n854_));
  NO2        m0826(.A(mai_mai_n618_), .B(mai_mai_n86_), .Y(mai_mai_n855_));
  NOi41      m0827(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n856_));
  NO2        m0828(.A(h), .B(mai_mai_n849_), .Y(mai_mai_n857_));
  OR3        m0829(.A(e), .B(d), .C(c), .Y(mai_mai_n858_));
  NA3        m0830(.A(k), .B(j), .C(i), .Y(mai_mai_n859_));
  NO3        m0831(.A(mai_mai_n859_), .B(mai_mai_n243_), .C(mai_mai_n68_), .Y(mai_mai_n860_));
  NOi21      m0832(.An(mai_mai_n860_), .B(mai_mai_n858_), .Y(mai_mai_n861_));
  OR4        m0833(.A(mai_mai_n861_), .B(mai_mai_n857_), .C(mai_mai_n854_), .D(mai_mai_n850_), .Y(mai_mai_n862_));
  NA3        m0834(.A(mai_mai_n369_), .B(mai_mai_n265_), .C(mai_mai_n44_), .Y(mai_mai_n863_));
  NO2        m0835(.A(mai_mai_n863_), .B(mai_mai_n853_), .Y(mai_mai_n864_));
  NO3        m0836(.A(mai_mai_n863_), .B(mai_mai_n460_), .C(mai_mai_n354_), .Y(mai_mai_n865_));
  NO2        m0837(.A(f), .B(c), .Y(mai_mai_n866_));
  NOi21      m0838(.An(mai_mai_n866_), .B(mai_mai_n348_), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n867_), .B(mai_mai_n46_), .Y(mai_mai_n868_));
  NO3        m0840(.A(i), .B(mai_mai_n199_), .C(l), .Y(mai_mai_n869_));
  NOi31      m0841(.An(mai_mai_n869_), .B(mai_mai_n868_), .C(j), .Y(mai_mai_n870_));
  OR3        m0842(.A(mai_mai_n870_), .B(mai_mai_n865_), .C(mai_mai_n864_), .Y(mai_mai_n871_));
  OR3        m0843(.A(mai_mai_n871_), .B(mai_mai_n862_), .C(mai_mai_n846_), .Y(mai02));
  OR3        m0844(.A(n), .B(m), .C(i), .Y(mai_mai_n873_));
  NO4        m0845(.A(mai_mai_n873_), .B(h), .C(l), .D(mai_mai_n858_), .Y(mai_mai_n874_));
  NOi31      m0846(.An(e), .B(d), .C(c), .Y(mai_mai_n875_));
  AOI210     m0847(.A0(mai_mai_n860_), .A1(mai_mai_n875_), .B0(mai_mai_n839_), .Y(mai_mai_n876_));
  AN3        m0848(.A(m), .B(f), .C(c), .Y(mai_mai_n877_));
  OR2        m0849(.A(mai_mai_n859_), .B(mai_mai_n243_), .Y(mai_mai_n878_));
  OR2        m0850(.A(mai_mai_n878_), .B(mai_mai_n1212_), .Y(mai_mai_n879_));
  NO3        m0851(.A(mai_mai_n863_), .B(i), .C(mai_mai_n460_), .Y(mai_mai_n880_));
  NO2        m0852(.A(mai_mai_n880_), .B(mai_mai_n850_), .Y(mai_mai_n881_));
  NA3        m0853(.A(l), .B(k), .C(j), .Y(mai_mai_n882_));
  NA2        m0854(.A(i), .B(h), .Y(mai_mai_n883_));
  NO3        m0855(.A(mai_mai_n883_), .B(mai_mai_n882_), .C(mai_mai_n99_), .Y(mai_mai_n884_));
  NO3        m0856(.A(mai_mai_n110_), .B(mai_mai_n231_), .C(mai_mai_n173_), .Y(mai_mai_n885_));
  AOI210     m0857(.A0(mai_mai_n885_), .A1(mai_mai_n884_), .B0(mai_mai_n854_), .Y(mai_mai_n886_));
  NA3        m0858(.A(c), .B(b), .C(a), .Y(mai_mai_n887_));
  NO3        m0859(.A(mai_mai_n859_), .B(mai_mai_n238_), .C(mai_mai_n39_), .Y(mai_mai_n888_));
  AOI210     m0860(.A0(mai_mai_n888_), .A1(a), .B0(mai_mai_n864_), .Y(mai_mai_n889_));
  AN4        m0861(.A(mai_mai_n889_), .B(mai_mai_n886_), .C(mai_mai_n881_), .D(mai_mai_n879_), .Y(mai_mai_n890_));
  NO2        m0862(.A(mai_mai_n841_), .B(mai_mai_n840_), .Y(mai_mai_n891_));
  NA2        m0863(.A(h), .B(mai_mai_n141_), .Y(mai_mai_n892_));
  AOI210     m0864(.A0(mai_mai_n892_), .A1(mai_mai_n891_), .B0(mai_mai_n836_), .Y(mai_mai_n893_));
  NAi41      m0865(.An(mai_mai_n874_), .B(mai_mai_n893_), .C(mai_mai_n890_), .D(mai_mai_n876_), .Y(mai03));
  NO2        m0866(.A(mai_mai_n1202_), .B(mai_mai_n553_), .Y(mai_mai_n895_));
  NA4        m0867(.A(i), .B(mai_mai_n875_), .C(mai_mai_n274_), .D(mai_mai_n265_), .Y(mai_mai_n896_));
  NOi31      m0868(.An(m), .B(n), .C(f), .Y(mai_mai_n897_));
  NA2        m0869(.A(mai_mai_n897_), .B(mai_mai_n41_), .Y(mai_mai_n898_));
  NO2        m0870(.A(mai_mai_n717_), .B(mai_mai_n338_), .Y(mai_mai_n899_));
  INV        m0871(.A(mai_mai_n839_), .Y(mai_mai_n900_));
  NO2        m0872(.A(mai_mai_n883_), .B(mai_mai_n378_), .Y(mai_mai_n901_));
  NO2        m0873(.A(mai_mai_n64_), .B(m), .Y(mai_mai_n902_));
  NO2        m0874(.A(mai_mai_n901_), .B(mai_mai_n869_), .Y(mai_mai_n903_));
  OR2        m0875(.A(mai_mai_n903_), .B(mai_mai_n868_), .Y(mai_mai_n904_));
  NA3        m0876(.A(mai_mai_n904_), .B(mai_mai_n900_), .C(mai_mai_n896_), .Y(mai_mai_n905_));
  NO3        m0877(.A(mai_mai_n905_), .B(mai_mai_n895_), .C(mai_mai_n441_), .Y(mai_mai_n906_));
  NA2        m0878(.A(c), .B(b), .Y(mai_mai_n907_));
  NO2        m0879(.A(mai_mai_n563_), .B(mai_mai_n907_), .Y(mai_mai_n908_));
  NA2        m0880(.A(mai_mai_n700_), .B(mai_mai_n331_), .Y(mai_mai_n909_));
  NA2        m0881(.A(mai_mai_n909_), .B(mai_mai_n908_), .Y(mai_mai_n910_));
  NAi21      m0882(.An(f), .B(d), .Y(mai_mai_n911_));
  NO2        m0883(.A(mai_mai_n911_), .B(mai_mai_n887_), .Y(mai_mai_n912_));
  NA2        m0884(.A(mai_mai_n912_), .B(mai_mai_n87_), .Y(mai_mai_n913_));
  NO2        m0885(.A(mai_mai_n147_), .B(mai_mai_n196_), .Y(mai_mai_n914_));
  NA2        m0886(.A(mai_mai_n914_), .B(m), .Y(mai_mai_n915_));
  NO2        m0887(.A(mai_mai_n115_), .B(mai_mai_n915_), .Y(mai_mai_n916_));
  INV        m0888(.A(mai_mai_n916_), .Y(mai_mai_n917_));
  NA4        m0889(.A(mai_mai_n917_), .B(mai_mai_n913_), .C(mai_mai_n910_), .D(mai_mai_n906_), .Y(mai00));
  NO3        m0890(.A(mai_mai_n880_), .B(mai_mai_n773_), .C(mai_mai_n73_), .Y(mai_mai_n919_));
  NA3        m0891(.A(mai_mai_n919_), .B(mai_mai_n896_), .C(mai_mai_n805_), .Y(mai_mai_n920_));
  NA2        m0892(.A(mai_mai_n394_), .B(f), .Y(mai_mai_n921_));
  INV        m0893(.A(mai_mai_n812_), .Y(mai_mai_n922_));
  NA2        m0894(.A(mai_mai_n922_), .B(n), .Y(mai_mai_n923_));
  AOI210     m0895(.A0(mai_mai_n923_), .A1(mai_mai_n921_), .B0(mai_mai_n841_), .Y(mai_mai_n924_));
  NO4        m0896(.A(mai_mai_n924_), .B(mai_mai_n920_), .C(mai_mai_n223_), .D(mai_mai_n862_), .Y(mai_mai_n925_));
  NA3        m0897(.A(mai_mai_n132_), .B(mai_mai_n38_), .C(mai_mai_n37_), .Y(mai_mai_n926_));
  NOi31      m0898(.An(n), .B(m), .C(i), .Y(mai_mai_n927_));
  NA3        m0899(.A(mai_mai_n927_), .B(d), .C(mai_mai_n41_), .Y(mai_mai_n928_));
  NA2        m0900(.A(mai_mai_n926_), .B(mai_mai_n928_), .Y(mai_mai_n929_));
  INV        m0901(.A(mai_mai_n453_), .Y(mai_mai_n930_));
  NO2        m0902(.A(mai_mai_n930_), .B(mai_mai_n929_), .Y(mai_mai_n931_));
  NO3        m0903(.A(mai_mai_n379_), .B(mai_mai_n1207_), .C(mai_mai_n907_), .Y(mai_mai_n932_));
  NA3        m0904(.A(mai_mai_n309_), .B(mai_mai_n180_), .C(m), .Y(mai_mai_n933_));
  NO2        m0905(.A(h), .B(m), .Y(mai_mai_n934_));
  NA3        m0906(.A(mai_mai_n387_), .B(mai_mai_n934_), .C(b), .Y(mai_mai_n935_));
  AOI220     m0907(.A0(m), .A1(mai_mai_n414_), .B0(mai_mai_n763_), .B1(mai_mai_n452_), .Y(mai_mai_n936_));
  NA2        m0908(.A(mai_mai_n250_), .B(mai_mai_n203_), .Y(mai_mai_n937_));
  NA4        m0909(.A(mai_mai_n937_), .B(mai_mai_n936_), .C(mai_mai_n935_), .D(mai_mai_n933_), .Y(mai_mai_n938_));
  NO2        m0910(.A(mai_mai_n938_), .B(mai_mai_n932_), .Y(mai_mai_n939_));
  NA2        m0911(.A(mai_mai_n203_), .B(mai_mai_n276_), .Y(mai_mai_n940_));
  INV        m0912(.A(mai_mai_n940_), .Y(mai_mai_n941_));
  NOi31      m0913(.An(mai_mai_n704_), .B(h), .C(mai_mai_n1211_), .Y(mai_mai_n942_));
  NAi31      m0914(.An(mai_mai_n150_), .B(mai_mai_n697_), .C(mai_mai_n369_), .Y(mai_mai_n943_));
  NAi21      m0915(.An(mai_mai_n942_), .B(mai_mai_n943_), .Y(mai_mai_n944_));
  INV        m0916(.A(mai_mai_n874_), .Y(mai_mai_n945_));
  NAi21      m0917(.An(mai_mai_n844_), .B(mai_mai_n945_), .Y(mai_mai_n946_));
  NO3        m0918(.A(mai_mai_n946_), .B(mai_mai_n944_), .C(mai_mai_n941_), .Y(mai_mai_n947_));
  AN3        m0919(.A(mai_mai_n947_), .B(mai_mai_n939_), .C(mai_mai_n931_), .Y(mai_mai_n948_));
  NA4        m0920(.A(d), .B(mai_mai_n168_), .C(mai_mai_n180_), .D(mai_mai_n129_), .Y(mai_mai_n949_));
  NA2        m0921(.A(mai_mai_n949_), .B(mai_mai_n234_), .Y(mai_mai_n950_));
  OR4        m0922(.A(mai_mai_n841_), .B(h), .C(mai_mai_n181_), .D(e), .Y(mai_mai_n951_));
  INV        m0923(.A(mai_mai_n114_), .Y(mai_mai_n952_));
  AOI220     m0924(.A0(mai_mai_n952_), .A1(mai_mai_n221_), .B0(mai_mai_n687_), .B1(mai_mai_n174_), .Y(mai_mai_n953_));
  NA2        m0925(.A(e), .B(mai_mai_n353_), .Y(mai_mai_n954_));
  NA3        m0926(.A(mai_mai_n954_), .B(mai_mai_n953_), .C(mai_mai_n951_), .Y(mai_mai_n955_));
  AOI220     m0927(.A0(mai_mai_n770_), .A1(mai_mai_n452_), .B0(d), .B1(mai_mai_n200_), .Y(mai_mai_n956_));
  NO3        m0928(.A(mai_mai_n841_), .B(mai_mai_n840_), .C(mai_mai_n587_), .Y(mai_mai_n957_));
  INV        m0929(.A(mai_mai_n957_), .Y(mai_mai_n958_));
  NA3        m0930(.A(mai_mai_n958_), .B(mai_mai_n956_), .C(mai_mai_n702_), .Y(mai_mai_n959_));
  NO3        m0931(.A(mai_mai_n959_), .B(mai_mai_n955_), .C(mai_mai_n950_), .Y(mai_mai_n960_));
  NA2        m0932(.A(e), .B(mai_mai_n616_), .Y(mai_mai_n961_));
  NA4        m0933(.A(mai_mai_n961_), .B(mai_mai_n960_), .C(mai_mai_n948_), .D(mai_mai_n925_), .Y(mai01));
  AN2        m0934(.A(mai_mai_n826_), .B(mai_mai_n824_), .Y(mai_mai_n963_));
  NO3        m0935(.A(mai_mai_n658_), .B(mai_mai_n651_), .C(mai_mai_n229_), .Y(mai_mai_n964_));
  NA2        m0936(.A(mai_mai_n320_), .B(i), .Y(mai_mai_n965_));
  NA3        m0937(.A(mai_mai_n965_), .B(mai_mai_n964_), .C(mai_mai_n963_), .Y(mai_mai_n966_));
  NA2        m0938(.A(mai_mai_n462_), .B(mai_mai_n67_), .Y(mai_mai_n967_));
  NA2        m0939(.A(mai_mai_n967_), .B(mai_mai_n740_), .Y(mai_mai_n968_));
  NA2        m0940(.A(mai_mai_n569_), .B(m), .Y(mai_mai_n969_));
  NO2        m0941(.A(mai_mai_n969_), .B(mai_mai_n1197_), .Y(mai_mai_n970_));
  INV        m0942(.A(mai_mai_n949_), .Y(mai_mai_n971_));
  AOI210     m0943(.A0(mai_mai_n970_), .A1(mai_mai_n504_), .B0(mai_mai_n971_), .Y(mai_mai_n972_));
  OA220      m0944(.A0(mai_mai_n1199_), .A1(mai_mai_n459_), .B0(n), .B1(mai_mai_n295_), .Y(mai_mai_n973_));
  NAi41      m0945(.An(mai_mai_n128_), .B(mai_mai_n973_), .C(mai_mai_n972_), .D(mai_mai_n727_), .Y(mai_mai_n974_));
  NO3        m0946(.A(mai_mai_n640_), .B(mai_mai_n540_), .C(mai_mai_n397_), .Y(mai_mai_n975_));
  NA3        m0947(.A(mai_mai_n569_), .B(mai_mai_n37_), .C(mai_mai_n172_), .Y(mai_mai_n976_));
  OA220      m0948(.A0(mai_mai_n976_), .A1(mai_mai_n534_), .B0(mai_mai_n160_), .B1(mai_mai_n158_), .Y(mai_mai_n977_));
  NA3        m0949(.A(mai_mai_n977_), .B(mai_mai_n975_), .C(mai_mai_n105_), .Y(mai_mai_n978_));
  NO4        m0950(.A(mai_mai_n978_), .B(mai_mai_n974_), .C(mai_mai_n968_), .D(mai_mai_n966_), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n417_), .B(mai_mai_n322_), .Y(mai_mai_n980_));
  NOi21      m0952(.An(mai_mai_n438_), .B(mai_mai_n458_), .Y(mai_mai_n981_));
  NA2        m0953(.A(mai_mai_n981_), .B(mai_mai_n980_), .Y(mai_mai_n982_));
  AOI210     m0954(.A0(mai_mai_n167_), .A1(mai_mai_n66_), .B0(mai_mai_n172_), .Y(mai_mai_n983_));
  OAI210     m0955(.A0(mai_mai_n662_), .A1(mai_mai_n339_), .B0(mai_mai_n983_), .Y(mai_mai_n984_));
  OR2        m0956(.A(mai_mai_n1203_), .B(mai_mai_n264_), .Y(mai_mai_n985_));
  NA3        m0957(.A(mai_mai_n985_), .B(mai_mai_n984_), .C(mai_mai_n982_), .Y(mai_mai_n986_));
  NA2        m0958(.A(mai_mai_n471_), .B(k), .Y(mai_mai_n987_));
  OAI210     m0959(.A0(mai_mai_n1199_), .A1(mai_mai_n468_), .B0(mai_mai_n987_), .Y(mai_mai_n988_));
  NA2        m0960(.A(mai_mai_n228_), .B(mai_mai_n160_), .Y(mai_mai_n989_));
  OAI210     m0961(.A0(mai_mai_n989_), .A1(mai_mai_n311_), .B0(mai_mai_n531_), .Y(mai_mai_n990_));
  INV        m0962(.A(mai_mai_n773_), .Y(mai_mai_n991_));
  OAI210     m0963(.A0(mai_mai_n970_), .A1(mai_mai_n258_), .B0(mai_mai_n541_), .Y(mai_mai_n992_));
  NA4        m0964(.A(mai_mai_n992_), .B(mai_mai_n991_), .C(mai_mai_n990_), .D(mai_mai_n643_), .Y(mai_mai_n993_));
  NO3        m0965(.A(mai_mai_n993_), .B(mai_mai_n988_), .C(mai_mai_n986_), .Y(mai_mai_n994_));
  NA3        m0966(.A(mai_mai_n477_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n995_));
  NO2        m0967(.A(mai_mai_n995_), .B(mai_mai_n167_), .Y(mai_mai_n996_));
  INV        m0968(.A(mai_mai_n996_), .Y(mai_mai_n997_));
  OR3        m0969(.A(mai_mai_n969_), .B(mai_mai_n478_), .C(mai_mai_n1197_), .Y(mai_mai_n998_));
  NO2        m0970(.A(mai_mai_n976_), .B(mai_mai_n787_), .Y(mai_mai_n999_));
  NO2        m0971(.A(mai_mai_n999_), .B(mai_mai_n929_), .Y(mai_mai_n1000_));
  NA4        m0972(.A(mai_mai_n1000_), .B(mai_mai_n998_), .C(mai_mai_n997_), .D(mai_mai_n615_), .Y(mai_mai_n1001_));
  NO2        m0973(.A(m), .B(mai_mai_n191_), .Y(mai_mai_n1002_));
  NO2        m0974(.A(mai_mai_n778_), .B(mai_mai_n432_), .Y(mai_mai_n1003_));
  OAI210     m0975(.A0(mai_mai_n1003_), .A1(mai_mai_n1002_), .B0(mai_mai_n272_), .Y(mai_mai_n1004_));
  NA2        m0976(.A(mai_mai_n448_), .B(mai_mai_n446_), .Y(mai_mai_n1005_));
  NO3        m0977(.A(mai_mai_n57_), .B(mai_mai_n238_), .C(mai_mai_n37_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n1006_), .B(mai_mai_n429_), .Y(mai_mai_n1007_));
  NA3        m0979(.A(mai_mai_n1007_), .B(mai_mai_n1005_), .C(mai_mai_n536_), .Y(mai_mai_n1008_));
  BUFFER     m0980(.A(mai_mai_n933_), .Y(mai_mai_n1009_));
  NO2        m0981(.A(mai_mai_n295_), .B(mai_mai_n50_), .Y(mai_mai_n1010_));
  INV        m0982(.A(mai_mai_n1010_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(mai_mai_n1006_), .B(mai_mai_n665_), .Y(mai_mai_n1012_));
  NA4        m0984(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .C(mai_mai_n1009_), .D(mai_mai_n312_), .Y(mai_mai_n1013_));
  NOi41      m0985(.An(mai_mai_n1004_), .B(mai_mai_n1013_), .C(mai_mai_n1008_), .D(mai_mai_n1001_), .Y(mai_mai_n1014_));
  AO220      m0986(.A0(i), .A1(mai_mai_n492_), .B0(mai_mai_n1209_), .B1(mai_mai_n567_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(mai_mai_n1015_), .B(mai_mai_n272_), .Y(mai_mai_n1016_));
  NA2        m0988(.A(mai_mai_n364_), .B(mai_mai_n102_), .Y(mai_mai_n1017_));
  NO3        m0989(.A(mai_mai_n883_), .B(mai_mai_n141_), .C(mai_mai_n64_), .Y(mai_mai_n1018_));
  AOI220     m0990(.A0(mai_mai_n1018_), .A1(mai_mai_n1017_), .B0(mai_mai_n1006_), .B1(mai_mai_n779_), .Y(mai_mai_n1019_));
  NA2        m0991(.A(mai_mai_n1019_), .B(mai_mai_n1016_), .Y(mai_mai_n1020_));
  NO2        m0992(.A(mai_mai_n484_), .B(mai_mai_n483_), .Y(mai_mai_n1021_));
  NO4        m0993(.A(mai_mai_n883_), .B(mai_mai_n1021_), .C(mai_mai_n139_), .D(mai_mai_n64_), .Y(mai_mai_n1022_));
  NO3        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1020_), .C(mai_mai_n507_), .Y(mai_mai_n1023_));
  NA4        m0995(.A(mai_mai_n1023_), .B(mai_mai_n1014_), .C(mai_mai_n994_), .D(mai_mai_n979_), .Y(mai06));
  NO2        m0996(.A(mai_mai_n1204_), .B(mai_mai_n435_), .Y(mai_mai_n1025_));
  NA2        m0997(.A(mai_mai_n216_), .B(mai_mai_n1025_), .Y(mai_mai_n1026_));
  NO2        m0998(.A(mai_mai_n183_), .B(mai_mai_n78_), .Y(mai_mai_n1027_));
  OAI210     m0999(.A0(mai_mai_n1027_), .A1(mai_mai_n1018_), .B0(mai_mai_n308_), .Y(mai_mai_n1028_));
  NO3        m1000(.A(mai_mai_n474_), .B(mai_mai_n660_), .C(mai_mai_n475_), .Y(mai_mai_n1029_));
  OR2        m1001(.A(mai_mai_n1029_), .B(mai_mai_n717_), .Y(mai_mai_n1030_));
  NA4        m1002(.A(mai_mai_n1030_), .B(mai_mai_n1028_), .C(mai_mai_n1026_), .D(mai_mai_n1004_), .Y(mai_mai_n1031_));
  NO3        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1008_), .C(mai_mai_n213_), .Y(mai_mai_n1032_));
  NA2        m1004(.A(i), .B(mai_mai_n780_), .Y(mai_mai_n1033_));
  AOI210     m1005(.A0(i), .A1(mai_mai_n433_), .B0(mai_mai_n1015_), .Y(mai_mai_n1034_));
  AOI210     m1006(.A0(mai_mai_n1034_), .A1(mai_mai_n1033_), .B0(mai_mai_n269_), .Y(mai_mai_n1035_));
  INV        m1007(.A(mai_mai_n539_), .Y(mai_mai_n1036_));
  NA2        m1008(.A(mai_mai_n1036_), .B(mai_mai_n510_), .Y(mai_mai_n1037_));
  NO2        m1009(.A(mai_mai_n400_), .B(mai_mai_n137_), .Y(mai_mai_n1038_));
  INV        m1010(.A(mai_mai_n898_), .Y(mai_mai_n1039_));
  OAI210     m1011(.A0(mai_mai_n364_), .A1(mai_mai_n204_), .B0(mai_mai_n734_), .Y(mai_mai_n1040_));
  NO4        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1039_), .C(mai_mai_n104_), .D(mai_mai_n1038_), .Y(mai_mai_n1041_));
  NO2        m1013(.A(mai_mai_n294_), .B(mai_mai_n103_), .Y(mai_mai_n1042_));
  NA2        m1014(.A(mai_mai_n1042_), .B(mai_mai_n462_), .Y(mai_mai_n1043_));
  NA3        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1041_), .C(mai_mai_n1037_), .Y(mai_mai_n1044_));
  NO2        m1016(.A(mai_mai_n606_), .B(mai_mai_n293_), .Y(mai_mai_n1045_));
  NO2        m1017(.A(mai_mai_n541_), .B(mai_mai_n617_), .Y(mai_mai_n1046_));
  NOi21      m1018(.An(mai_mai_n1045_), .B(mai_mai_n1046_), .Y(mai_mai_n1047_));
  AN2        m1019(.A(mai_mai_n770_), .B(mai_mai_n513_), .Y(mai_mai_n1048_));
  NO4        m1020(.A(mai_mai_n1048_), .B(mai_mai_n1047_), .C(mai_mai_n1044_), .D(mai_mai_n1035_), .Y(mai_mai_n1049_));
  INV        m1021(.A(mai_mai_n224_), .Y(mai_mai_n1050_));
  OAI210     m1022(.A0(mai_mai_n183_), .A1(mai_mai_n486_), .B0(mai_mai_n592_), .Y(mai_mai_n1051_));
  OAI210     m1023(.A0(mai_mai_n224_), .A1(c), .B0(mai_mai_n509_), .Y(mai_mai_n1052_));
  AOI220     m1024(.A0(mai_mai_n1052_), .A1(mai_mai_n1051_), .B0(mai_mai_n1050_), .B1(mai_mai_n216_), .Y(mai_mai_n1053_));
  OAI220     m1025(.A0(mai_mai_n560_), .A1(mai_mai_n204_), .B0(mai_mai_n396_), .B1(mai_mai_n400_), .Y(mai_mai_n1054_));
  OAI210     m1026(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1055_));
  NO3        m1027(.A(mai_mai_n1055_), .B(mai_mai_n473_), .C(j), .Y(mai_mai_n1056_));
  NOi21      m1028(.An(mai_mai_n1056_), .B(mai_mai_n534_), .Y(mai_mai_n1057_));
  NO3        m1029(.A(mai_mai_n1057_), .B(mai_mai_n1054_), .C(mai_mai_n899_), .Y(mai_mai_n1058_));
  NA3        m1030(.A(mai_mai_n649_), .B(mai_mai_n648_), .C(mai_mai_n344_), .Y(mai_mai_n1059_));
  NAi31      m1031(.An(mai_mai_n606_), .B(mai_mai_n1059_), .C(mai_mai_n166_), .Y(mai_mai_n1060_));
  NA4        m1032(.A(mai_mai_n1060_), .B(mai_mai_n1058_), .C(mai_mai_n1053_), .D(mai_mai_n956_), .Y(mai_mai_n1061_));
  OR2        m1033(.A(mai_mai_n639_), .B(mai_mai_n419_), .Y(mai_mai_n1062_));
  OR3        m1034(.A(mai_mai_n296_), .B(mai_mai_n183_), .C(mai_mai_n486_), .Y(mai_mai_n1063_));
  AOI210     m1035(.A0(mai_mai_n448_), .A1(mai_mai_n353_), .B0(mai_mai_n298_), .Y(mai_mai_n1064_));
  NA2        m1036(.A(mai_mai_n1056_), .B(mai_mai_n645_), .Y(mai_mai_n1065_));
  NA4        m1037(.A(mai_mai_n1065_), .B(mai_mai_n1064_), .C(mai_mai_n1063_), .D(mai_mai_n1062_), .Y(mai_mai_n1066_));
  NA2        m1038(.A(mai_mai_n1045_), .B(mai_mai_n616_), .Y(mai_mai_n1067_));
  AO220      m1039(.A0(mai_mai_n1027_), .A1(mai_mai_n531_), .B0(mai_mai_n750_), .B1(mai_mai_n749_), .Y(mai_mai_n1068_));
  NO4        m1040(.A(mai_mai_n1068_), .B(mai_mai_n708_), .C(mai_mai_n388_), .D(mai_mai_n375_), .Y(mai_mai_n1069_));
  NA3        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1067_), .C(mai_mai_n1012_), .Y(mai_mai_n1070_));
  NAi21      m1042(.An(j), .B(i), .Y(mai_mai_n1071_));
  NO4        m1043(.A(mai_mai_n1021_), .B(mai_mai_n1071_), .C(mai_mai_n348_), .D(mai_mai_n194_), .Y(mai_mai_n1072_));
  NO4        m1044(.A(mai_mai_n1072_), .B(mai_mai_n1070_), .C(mai_mai_n1066_), .D(mai_mai_n1061_), .Y(mai_mai_n1073_));
  NA4        m1045(.A(mai_mai_n1073_), .B(mai_mai_n1049_), .C(mai_mai_n1032_), .D(mai_mai_n1023_), .Y(mai07));
  NOi21      m1046(.An(j), .B(k), .Y(mai_mai_n1075_));
  NA4        m1047(.A(mai_mai_n144_), .B(mai_mai_n83_), .C(mai_mai_n1075_), .D(f), .Y(mai_mai_n1076_));
  NAi32      m1048(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1077_));
  NO3        m1049(.A(mai_mai_n1077_), .B(m), .C(f), .Y(mai_mai_n1078_));
  OAI210     m1050(.A0(i), .A1(mai_mai_n377_), .B0(mai_mai_n1078_), .Y(mai_mai_n1079_));
  NAi21      m1051(.An(f), .B(c), .Y(mai_mai_n1080_));
  OR2        m1052(.A(e), .B(d), .Y(mai_mai_n1081_));
  NO2        m1053(.A(mai_mai_n496_), .B(mai_mai_n254_), .Y(mai_mai_n1082_));
  NA3        m1054(.A(mai_mai_n1082_), .B(mai_mai_n852_), .C(mai_mai_n144_), .Y(mai_mai_n1083_));
  NOi31      m1055(.An(n), .B(m), .C(b), .Y(mai_mai_n1084_));
  NO3        m1056(.A(mai_mai_n99_), .B(mai_mai_n354_), .C(h), .Y(mai_mai_n1085_));
  NA3        m1057(.A(mai_mai_n1083_), .B(mai_mai_n1079_), .C(mai_mai_n1076_), .Y(mai_mai_n1086_));
  NO2        m1058(.A(k), .B(i), .Y(mai_mai_n1087_));
  NA3        m1059(.A(mai_mai_n1087_), .B(mai_mai_n726_), .C(mai_mai_n144_), .Y(mai_mai_n1088_));
  NO2        m1060(.A(mai_mai_n859_), .B(mai_mai_n243_), .Y(mai_mai_n1089_));
  INV        m1061(.A(mai_mai_n1088_), .Y(mai_mai_n1090_));
  NO2        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1086_), .Y(mai_mai_n1091_));
  NO3        m1063(.A(e), .B(d), .C(c), .Y(mai_mai_n1092_));
  OAI210     m1064(.A0(mai_mai_n99_), .A1(mai_mai_n173_), .B0(mai_mai_n479_), .Y(mai_mai_n1093_));
  NA2        m1065(.A(mai_mai_n1093_), .B(mai_mai_n1092_), .Y(mai_mai_n1094_));
  INV        m1066(.A(mai_mai_n1094_), .Y(mai_mai_n1095_));
  NO2        m1067(.A(l), .B(k), .Y(mai_mai_n1096_));
  NOi41      m1068(.An(mai_mai_n424_), .B(mai_mai_n1096_), .C(mai_mai_n372_), .D(mai_mai_n348_), .Y(mai_mai_n1097_));
  NO3        m1069(.A(mai_mai_n348_), .B(d), .C(c), .Y(mai_mai_n1098_));
  NO2        m1070(.A(mai_mai_n1097_), .B(mai_mai_n1095_), .Y(mai_mai_n1099_));
  NO2        m1071(.A(m), .B(c), .Y(mai_mai_n1100_));
  NA3        m1072(.A(mai_mai_n1100_), .B(mai_mai_n110_), .C(mai_mai_n151_), .Y(mai_mai_n1101_));
  NO2        m1073(.A(mai_mai_n1101_), .B(mai_mai_n1196_), .Y(mai_mai_n1102_));
  NA2        m1074(.A(mai_mai_n1102_), .B(mai_mai_n144_), .Y(mai_mai_n1103_));
  NO2        m1075(.A(mai_mai_n355_), .B(a), .Y(mai_mai_n1104_));
  NA3        m1076(.A(mai_mai_n1104_), .B(k), .C(mai_mai_n87_), .Y(mai_mai_n1105_));
  NO2        m1077(.A(i), .B(h), .Y(mai_mai_n1106_));
  NA2        m1078(.A(mai_mai_n911_), .B(h), .Y(mai_mai_n1107_));
  NA2        m1079(.A(mai_mai_n106_), .B(mai_mai_n180_), .Y(mai_mai_n1108_));
  NO2        m1080(.A(mai_mai_n1108_), .B(mai_mai_n1107_), .Y(mai_mai_n1109_));
  NOi31      m1081(.An(m), .B(n), .C(b), .Y(mai_mai_n1110_));
  NOi31      m1082(.An(f), .B(d), .C(c), .Y(mai_mai_n1111_));
  NA2        m1083(.A(mai_mai_n1111_), .B(mai_mai_n1110_), .Y(mai_mai_n1112_));
  INV        m1084(.A(mai_mai_n1112_), .Y(mai_mai_n1113_));
  NO2        m1085(.A(mai_mai_n1113_), .B(mai_mai_n1109_), .Y(mai_mai_n1114_));
  NA2        m1086(.A(mai_mai_n877_), .B(mai_mai_n369_), .Y(mai_mai_n1115_));
  NO4        m1087(.A(mai_mai_n1115_), .B(mai_mai_n855_), .C(mai_mai_n348_), .D(mai_mai_n37_), .Y(mai_mai_n1116_));
  NA2        m1088(.A(mai_mai_n147_), .B(mai_mai_n856_), .Y(mai_mai_n1117_));
  INV        m1089(.A(mai_mai_n1117_), .Y(mai_mai_n1118_));
  NO2        m1090(.A(mai_mai_n1118_), .B(mai_mai_n1116_), .Y(mai_mai_n1119_));
  AN4        m1091(.A(mai_mai_n1119_), .B(mai_mai_n1114_), .C(mai_mai_n1105_), .D(mai_mai_n1103_), .Y(mai_mai_n1120_));
  NA2        m1092(.A(mai_mai_n1084_), .B(mai_mai_n305_), .Y(mai_mai_n1121_));
  NA2        m1093(.A(mai_mai_n1098_), .B(mai_mai_n174_), .Y(mai_mai_n1122_));
  NA2        m1094(.A(mai_mai_n884_), .B(mai_mai_n1115_), .Y(mai_mai_n1123_));
  NA2        m1095(.A(mai_mai_n1123_), .B(mai_mai_n1122_), .Y(mai_mai_n1124_));
  NO4        m1096(.A(mai_mai_n99_), .B(m), .C(f), .D(e), .Y(mai_mai_n1125_));
  NA3        m1097(.A(mai_mai_n1087_), .B(mai_mai_n233_), .C(h), .Y(mai_mai_n1126_));
  OR2        m1098(.A(e), .B(a), .Y(mai_mai_n1127_));
  NO2        m1099(.A(mai_mai_n1081_), .B(mai_mai_n1080_), .Y(mai_mai_n1128_));
  INV        m1100(.A(mai_mai_n1128_), .Y(mai_mai_n1129_));
  NO2        m1101(.A(mai_mai_n1129_), .B(mai_mai_n873_), .Y(mai_mai_n1130_));
  NO2        m1102(.A(mai_mai_n1130_), .B(mai_mai_n1124_), .Y(mai_mai_n1131_));
  NA4        m1103(.A(mai_mai_n1131_), .B(mai_mai_n1120_), .C(mai_mai_n1099_), .D(mai_mai_n1091_), .Y(mai_mai_n1132_));
  NO2        m1104(.A(mai_mai_n317_), .B(j), .Y(mai_mai_n1133_));
  NAi41      m1105(.An(mai_mai_n1106_), .B(mai_mai_n867_), .C(mai_mai_n133_), .D(mai_mai_n117_), .Y(mai_mai_n1134_));
  INV        m1106(.A(mai_mai_n1134_), .Y(mai_mai_n1135_));
  NA3        m1107(.A(m), .B(mai_mai_n1133_), .C(mai_mai_n125_), .Y(mai_mai_n1136_));
  INV        m1108(.A(mai_mai_n1136_), .Y(mai_mai_n1137_));
  NO3        m1109(.A(mai_mai_n606_), .B(mai_mai_n139_), .C(mai_mai_n330_), .Y(mai_mai_n1138_));
  NO3        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1137_), .C(mai_mai_n1135_), .Y(mai_mai_n1139_));
  OR2        m1111(.A(n), .B(i), .Y(mai_mai_n1140_));
  NO2        m1112(.A(mai_mai_n1140_), .B(mai_mai_n866_), .Y(mai_mai_n1141_));
  NA2        m1113(.A(mai_mai_n1141_), .B(mai_mai_n934_), .Y(mai_mai_n1142_));
  NO3        m1114(.A(mai_mai_n887_), .B(mai_mai_n1081_), .C(mai_mai_n39_), .Y(mai_mai_n1143_));
  NO2        m1115(.A(mai_mai_n873_), .B(h), .Y(mai_mai_n1144_));
  NA3        m1116(.A(mai_mai_n1144_), .B(d), .C(mai_mai_n840_), .Y(mai_mai_n1145_));
  NO2        m1117(.A(mai_mai_n1145_), .B(c), .Y(mai_mai_n1146_));
  NA2        m1118(.A(mai_mai_n144_), .B(mai_mai_n86_), .Y(mai_mai_n1147_));
  INV        m1119(.A(mai_mai_n1146_), .Y(mai_mai_n1148_));
  NA3        m1120(.A(mai_mai_n1148_), .B(mai_mai_n1142_), .C(mai_mai_n1139_), .Y(mai_mai_n1149_));
  NO3        m1121(.A(mai_mai_n877_), .B(mai_mai_n866_), .C(mai_mai_n35_), .Y(mai_mai_n1150_));
  NA2        m1122(.A(mai_mai_n1150_), .B(mai_mai_n1089_), .Y(mai_mai_n1151_));
  OAI210     m1123(.A0(mai_mai_n1125_), .A1(mai_mai_n1084_), .B0(mai_mai_n714_), .Y(mai_mai_n1152_));
  NO2        m1124(.A(mai_mai_n838_), .B(mai_mai_n99_), .Y(mai_mai_n1153_));
  NA2        m1125(.A(mai_mai_n1153_), .B(mai_mai_n491_), .Y(mai_mai_n1154_));
  NA3        m1126(.A(mai_mai_n1154_), .B(mai_mai_n1152_), .C(mai_mai_n1151_), .Y(mai_mai_n1155_));
  OAI220     m1127(.A0(mai_mai_n118_), .A1(mai_mai_n146_), .B0(mai_mai_n354_), .B1(m), .Y(mai_mai_n1156_));
  OAI210     m1128(.A0(mai_mai_n1156_), .A1(mai_mai_n84_), .B0(mai_mai_n1110_), .Y(mai_mai_n1157_));
  INV        m1129(.A(mai_mai_n1157_), .Y(mai_mai_n1158_));
  NO2        m1130(.A(mai_mai_n1158_), .B(mai_mai_n1155_), .Y(mai_mai_n1159_));
  NO2        m1131(.A(mai_mai_n1080_), .B(e), .Y(mai_mai_n1160_));
  NO2        m1132(.A(mai_mai_n146_), .B(c), .Y(mai_mai_n1161_));
  OAI210     m1133(.A0(mai_mai_n1161_), .A1(mai_mai_n1160_), .B0(mai_mai_n144_), .Y(mai_mai_n1162_));
  AOI220     m1134(.A0(mai_mai_n1162_), .A1(mai_mai_n868_), .B0(mai_mai_n411_), .B1(mai_mai_n293_), .Y(mai_mai_n1163_));
  INV        m1135(.A(mai_mai_n1143_), .Y(mai_mai_n1164_));
  NO2        m1136(.A(mai_mai_n1127_), .B(f), .Y(mai_mai_n1165_));
  AOI210     m1137(.A0(mai_mai_n902_), .A1(a), .B0(mai_mai_n1165_), .Y(mai_mai_n1166_));
  OAI210     m1138(.A0(mai_mai_n1166_), .A1(mai_mai_n48_), .B0(mai_mai_n1164_), .Y(mai_mai_n1167_));
  AOI210     m1139(.A0(mai_mai_n729_), .A1(mai_mai_n334_), .B0(mai_mai_n80_), .Y(mai_mai_n1168_));
  OR2        m1140(.A(mai_mai_n1168_), .B(mai_mai_n418_), .Y(mai_mai_n1169_));
  NO2        m1141(.A(mai_mai_n1169_), .B(mai_mai_n139_), .Y(mai_mai_n1170_));
  NA4        m1142(.A(mai_mai_n885_), .B(mai_mai_n882_), .C(mai_mai_n180_), .D(i), .Y(mai_mai_n1171_));
  NA2        m1143(.A(mai_mai_n1085_), .B(mai_mai_n147_), .Y(mai_mai_n1172_));
  NO2        m1144(.A(mai_mai_n39_), .B(l), .Y(mai_mai_n1173_));
  OAI210     m1145(.A0(mai_mai_n1127_), .A1(mai_mai_n699_), .B0(mai_mai_n377_), .Y(mai_mai_n1174_));
  NA2        m1146(.A(mai_mai_n1174_), .B(mai_mai_n1173_), .Y(mai_mai_n1175_));
  NA3        m1147(.A(mai_mai_n1175_), .B(mai_mai_n1172_), .C(mai_mai_n1171_), .Y(mai_mai_n1176_));
  NO4        m1148(.A(mai_mai_n1176_), .B(mai_mai_n1170_), .C(mai_mai_n1167_), .D(mai_mai_n1163_), .Y(mai_mai_n1177_));
  NA2        m1149(.A(mai_mai_n1177_), .B(mai_mai_n1159_), .Y(mai_mai_n1178_));
  AO210      m1150(.A0(mai_mai_n100_), .A1(l), .B0(mai_mai_n1121_), .Y(mai_mai_n1179_));
  NO4        m1151(.A(mai_mai_n183_), .B(mai_mai_n150_), .C(mai_mai_n214_), .D(k), .Y(mai_mai_n1180_));
  AOI210     m1152(.A0(mai_mai_n123_), .A1(mai_mai_n44_), .B0(mai_mai_n1160_), .Y(mai_mai_n1181_));
  NO2        m1153(.A(mai_mai_n1181_), .B(mai_mai_n1147_), .Y(mai_mai_n1182_));
  NOi21      m1154(.An(mai_mai_n1085_), .B(e), .Y(mai_mai_n1183_));
  NO3        m1155(.A(mai_mai_n1183_), .B(mai_mai_n1182_), .C(mai_mai_n1180_), .Y(mai_mai_n1184_));
  NA2        m1156(.A(mai_mai_n1184_), .B(mai_mai_n1179_), .Y(mai_mai_n1185_));
  OR4        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1178_), .C(mai_mai_n1149_), .D(mai_mai_n1132_), .Y(mai04));
  NOi31      m1158(.An(mai_mai_n1125_), .B(mai_mai_n1126_), .C(mai_mai_n841_), .Y(mai_mai_n1187_));
  NO3        m1159(.A(h), .B(mai_mai_n834_), .C(j), .Y(mai_mai_n1188_));
  OR3        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1187_), .C(mai_mai_n857_), .Y(mai_mai_n1189_));
  AOI210     m1161(.A0(mai_mai_n1210_), .A1(mai_mai_n851_), .B0(mai_mai_n942_), .Y(mai_mai_n1190_));
  NA2        m1162(.A(mai_mai_n1190_), .B(mai_mai_n958_), .Y(mai_mai_n1191_));
  NO4        m1163(.A(mai_mai_n1191_), .B(mai_mai_n1189_), .C(mai_mai_n865_), .D(mai_mai_n846_), .Y(mai_mai_n1192_));
  NA4        m1164(.A(mai_mai_n1192_), .B(mai_mai_n904_), .C(mai_mai_n896_), .D(mai_mai_n890_), .Y(mai05));
  INV        m1165(.A(l), .Y(mai_mai_n1196_));
  INV        m1166(.A(f), .Y(mai_mai_n1197_));
  INV        m1167(.A(j), .Y(mai_mai_n1198_));
  INV        m1168(.A(k), .Y(mai_mai_n1199_));
  INV        m1169(.A(m), .Y(mai_mai_n1200_));
  INV        m1170(.A(mai_mai_n504_), .Y(mai_mai_n1201_));
  INV        m1171(.A(m), .Y(mai_mai_n1202_));
  INV        m1172(.A(m), .Y(mai_mai_n1203_));
  INV        m1173(.A(e), .Y(mai_mai_n1204_));
  INV        m1174(.A(h), .Y(mai_mai_n1205_));
  INV        m1175(.A(e), .Y(mai_mai_n1206_));
  INV        m1176(.A(h), .Y(mai_mai_n1207_));
  INV        m1177(.A(j), .Y(mai_mai_n1208_));
  INV        m1178(.A(m), .Y(mai_mai_n1209_));
  INV        m1179(.A(m), .Y(mai_mai_n1210_));
  INV        m1180(.A(m), .Y(mai_mai_n1211_));
  INV        m1181(.A(f), .Y(mai_mai_n1212_));
  INV        m1182(.A(mai_mai_n348_), .Y(mai_mai_n1213_));
  INV        m1183(.A(f), .Y(mai_mai_n1214_));
  INV        m1184(.A(n), .Y(mai_mai_n1215_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  NA3        u0002(.A(e), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n31_));
  NOi32      u0003(.An(m), .Bn(l), .C(n), .Y(men_men_n32_));
  NOi32      u0004(.An(i), .Bn(u), .C(h), .Y(men_men_n33_));
  NA2        u0005(.A(men_men_n33_), .B(men_men_n32_), .Y(men_men_n34_));
  AN2        u0006(.A(m), .B(l), .Y(men_men_n35_));
  NOi32      u0007(.An(j), .Bn(u), .C(k), .Y(men_men_n36_));
  NA2        u0008(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n37_));
  NO2        u0009(.A(men_men_n37_), .B(n), .Y(men_men_n38_));
  INV        u0010(.A(h), .Y(men_men_n39_));
  NAi21      u0011(.An(j), .B(l), .Y(men_men_n40_));
  NAi32      u0012(.An(n), .Bn(u), .C(m), .Y(men_men_n41_));
  NO3        u0013(.A(men_men_n41_), .B(men_men_n40_), .C(men_men_n39_), .Y(men_men_n42_));
  NAi31      u0014(.An(n), .B(m), .C(l), .Y(men_men_n43_));
  INV        u0015(.A(i), .Y(men_men_n44_));
  AN2        u0016(.A(h), .B(u), .Y(men_men_n45_));
  NA2        u0017(.A(men_men_n45_), .B(men_men_n44_), .Y(men_men_n46_));
  NO2        u0018(.A(men_men_n46_), .B(men_men_n43_), .Y(men_men_n47_));
  NAi21      u0019(.An(n), .B(m), .Y(men_men_n48_));
  NOi32      u0020(.An(k), .Bn(h), .C(l), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(u), .Y(men_men_n50_));
  NO2        u0022(.A(men_men_n50_), .B(men_men_n49_), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n48_), .Y(men_men_n52_));
  NO4        u0024(.A(men_men_n52_), .B(men_men_n47_), .C(men_men_n42_), .D(men_men_n38_), .Y(men_men_n53_));
  AOI210     u0025(.A0(men_men_n53_), .A1(men_men_n34_), .B0(men_men_n31_), .Y(men_men_n54_));
  INV        u0026(.A(c), .Y(men_men_n55_));
  NA2        u0027(.A(e), .B(b), .Y(men_men_n56_));
  NO2        u0028(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  INV        u0029(.A(d), .Y(men_men_n58_));
  NA2        u0030(.A(u), .B(men_men_n58_), .Y(men_men_n59_));
  NAi21      u0031(.An(i), .B(h), .Y(men_men_n60_));
  NAi31      u0032(.An(i), .B(l), .C(j), .Y(men_men_n61_));
  OAI220     u0033(.A0(men_men_n61_), .A1(men_men_n48_), .B0(men_men_n60_), .B1(men_men_n43_), .Y(men_men_n62_));
  NAi31      u0034(.An(men_men_n59_), .B(men_men_n62_), .C(men_men_n57_), .Y(men_men_n63_));
  NAi41      u0035(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n64_));
  NA2        u0036(.A(u), .B(f), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi21      u0038(.An(i), .B(j), .Y(men_men_n67_));
  NAi32      u0039(.An(n), .Bn(k), .C(m), .Y(men_men_n68_));
  NO2        u0040(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi31      u0041(.An(l), .B(m), .C(k), .Y(men_men_n70_));
  NAi21      u0042(.An(e), .B(h), .Y(men_men_n71_));
  NAi41      u0043(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n73_));
  INV        u0045(.A(m), .Y(men_men_n74_));
  NOi21      u0046(.An(k), .B(l), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  AN4        u0048(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n77_));
  NA2        u0049(.A(h), .B(men_men_n77_), .Y(men_men_n78_));
  NOi32      u0050(.An(h), .Bn(u), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n80_));
  INV        u0052(.A(n), .Y(men_men_n81_));
  INV        u0053(.A(j), .Y(men_men_n82_));
  AN3        u0054(.A(m), .B(k), .C(i), .Y(men_men_n83_));
  NA3        u0055(.A(men_men_n83_), .B(men_men_n82_), .C(u), .Y(men_men_n84_));
  NO2        u0056(.A(men_men_n84_), .B(f), .Y(men_men_n85_));
  NAi32      u0057(.An(u), .Bn(f), .C(h), .Y(men_men_n86_));
  NAi31      u0058(.An(j), .B(m), .C(l), .Y(men_men_n87_));
  NO2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  NA2        u0060(.A(m), .B(l), .Y(men_men_n89_));
  NAi31      u0061(.An(k), .B(j), .C(u), .Y(men_men_n90_));
  NO3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(f), .Y(men_men_n91_));
  AN2        u0063(.A(j), .B(u), .Y(men_men_n92_));
  NOi32      u0064(.An(m), .Bn(l), .C(i), .Y(men_men_n93_));
  NOi21      u0065(.An(u), .B(i), .Y(men_men_n94_));
  NOi32      u0066(.An(m), .Bn(j), .C(k), .Y(men_men_n95_));
  AOI220     u0067(.A0(men_men_n95_), .A1(men_men_n94_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n96_));
  NO2        u0068(.A(men_men_n96_), .B(f), .Y(men_men_n97_));
  NAi41      u0069(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n98_));
  AN2        u0070(.A(e), .B(b), .Y(men_men_n99_));
  NA2        u0071(.A(c), .B(men_men_n99_), .Y(men_men_n100_));
  NO3        u0072(.A(men_men_n100_), .B(men_men_n98_), .C(u), .Y(men_men_n101_));
  NOi21      u0073(.An(u), .B(f), .Y(men_men_n102_));
  NOi21      u0074(.An(i), .B(h), .Y(men_men_n103_));
  NA3        u0075(.A(men_men_n103_), .B(men_men_n102_), .C(men_men_n35_), .Y(men_men_n104_));
  INV        u0076(.A(a), .Y(men_men_n105_));
  NA2        u0077(.A(men_men_n99_), .B(men_men_n105_), .Y(men_men_n106_));
  INV        u0078(.A(l), .Y(men_men_n107_));
  NOi21      u0079(.An(m), .B(n), .Y(men_men_n108_));
  AN2        u0080(.A(k), .B(h), .Y(men_men_n109_));
  INV        u0081(.A(b), .Y(men_men_n110_));
  NA2        u0082(.A(l), .B(j), .Y(men_men_n111_));
  AN2        u0083(.A(k), .B(i), .Y(men_men_n112_));
  NA2        u0084(.A(men_men_n112_), .B(men_men_n111_), .Y(men_men_n113_));
  NA2        u0085(.A(u), .B(e), .Y(men_men_n114_));
  NOi32      u0086(.An(c), .Bn(a), .C(d), .Y(men_men_n115_));
  NA2        u0087(.A(men_men_n115_), .B(men_men_n108_), .Y(men_men_n116_));
  NO4        u0088(.A(men_men_n116_), .B(men_men_n114_), .C(men_men_n113_), .D(men_men_n110_), .Y(men_men_n117_));
  NO2        u0089(.A(men_men_n117_), .B(men_men_n101_), .Y(men_men_n118_));
  INV        u0090(.A(men_men_n118_), .Y(men_men_n119_));
  NOi31      u0091(.An(k), .B(m), .C(j), .Y(men_men_n120_));
  NOi31      u0092(.An(k), .B(m), .C(i), .Y(men_men_n121_));
  NA3        u0093(.A(men_men_n121_), .B(men_men_n79_), .C(men_men_n77_), .Y(men_men_n122_));
  INV        u0094(.A(men_men_n122_), .Y(men_men_n123_));
  NOi32      u0095(.An(f), .Bn(b), .C(e), .Y(men_men_n124_));
  NAi21      u0096(.An(u), .B(h), .Y(men_men_n125_));
  NAi21      u0097(.An(m), .B(n), .Y(men_men_n126_));
  NO3        u0098(.A(j), .B(men_men_n126_), .C(men_men_n125_), .Y(men_men_n127_));
  NAi41      u0099(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n128_));
  NAi31      u0100(.An(j), .B(k), .C(h), .Y(men_men_n129_));
  NO3        u0101(.A(men_men_n129_), .B(men_men_n128_), .C(men_men_n126_), .Y(men_men_n130_));
  AOI210     u0102(.A0(men_men_n127_), .A1(men_men_n124_), .B0(men_men_n130_), .Y(men_men_n131_));
  NO2        u0103(.A(k), .B(j), .Y(men_men_n132_));
  AN2        u0104(.A(k), .B(j), .Y(men_men_n133_));
  NAi21      u0105(.An(c), .B(b), .Y(men_men_n134_));
  NA2        u0106(.A(f), .B(d), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n125_), .Y(men_men_n136_));
  NA2        u0108(.A(h), .B(c), .Y(men_men_n137_));
  NAi31      u0109(.An(f), .B(e), .C(b), .Y(men_men_n138_));
  NA2        u0110(.A(men_men_n136_), .B(n), .Y(men_men_n139_));
  NA2        u0111(.A(d), .B(b), .Y(men_men_n140_));
  NAi21      u0112(.An(e), .B(f), .Y(men_men_n141_));
  NO2        u0113(.A(men_men_n141_), .B(men_men_n140_), .Y(men_men_n142_));
  NA2        u0114(.A(b), .B(a), .Y(men_men_n143_));
  NAi21      u0115(.An(e), .B(u), .Y(men_men_n144_));
  NAi21      u0116(.An(c), .B(d), .Y(men_men_n145_));
  NAi31      u0117(.An(l), .B(k), .C(h), .Y(men_men_n146_));
  NO2        u0118(.A(men_men_n126_), .B(men_men_n146_), .Y(men_men_n147_));
  NA2        u0119(.A(men_men_n147_), .B(men_men_n142_), .Y(men_men_n148_));
  NAi41      u0120(.An(men_men_n123_), .B(men_men_n148_), .C(men_men_n139_), .D(men_men_n131_), .Y(men_men_n149_));
  NAi31      u0121(.An(e), .B(f), .C(b), .Y(men_men_n150_));
  NOi21      u0122(.An(u), .B(d), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n151_), .B(men_men_n150_), .Y(men_men_n152_));
  NOi21      u0124(.An(h), .B(i), .Y(men_men_n153_));
  NOi21      u0125(.An(k), .B(m), .Y(men_men_n154_));
  NA3        u0126(.A(men_men_n154_), .B(men_men_n153_), .C(n), .Y(men_men_n155_));
  NOi21      u0127(.An(men_men_n152_), .B(men_men_n155_), .Y(men_men_n156_));
  NOi21      u0128(.An(h), .B(u), .Y(men_men_n157_));
  NO2        u0129(.A(men_men_n135_), .B(men_men_n134_), .Y(men_men_n158_));
  NAi31      u0130(.An(l), .B(j), .C(h), .Y(men_men_n159_));
  NO2        u0131(.A(men_men_n159_), .B(men_men_n48_), .Y(men_men_n160_));
  NA2        u0132(.A(men_men_n160_), .B(men_men_n66_), .Y(men_men_n161_));
  NA2        u0133(.A(l), .B(i), .Y(men_men_n162_));
  INV        u0134(.A(men_men_n161_), .Y(men_men_n163_));
  NAi31      u0135(.An(d), .B(f), .C(c), .Y(men_men_n164_));
  NAi31      u0136(.An(e), .B(f), .C(c), .Y(men_men_n165_));
  NA2        u0137(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  NA2        u0138(.A(j), .B(h), .Y(men_men_n167_));
  OR3        u0139(.A(n), .B(m), .C(k), .Y(men_men_n168_));
  NO2        u0140(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  NAi32      u0141(.An(m), .Bn(k), .C(n), .Y(men_men_n170_));
  NO2        u0142(.A(men_men_n170_), .B(men_men_n167_), .Y(men_men_n171_));
  AOI220     u0143(.A0(men_men_n171_), .A1(men_men_n152_), .B0(men_men_n169_), .B1(men_men_n166_), .Y(men_men_n172_));
  NO2        u0144(.A(n), .B(m), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n49_), .Y(men_men_n174_));
  NAi21      u0146(.An(f), .B(e), .Y(men_men_n175_));
  NA2        u0147(.A(d), .B(c), .Y(men_men_n176_));
  NO2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  NOi21      u0149(.An(men_men_n177_), .B(men_men_n174_), .Y(men_men_n178_));
  NAi21      u0150(.An(d), .B(c), .Y(men_men_n179_));
  NAi31      u0151(.An(m), .B(n), .C(b), .Y(men_men_n180_));
  NA2        u0152(.A(k), .B(i), .Y(men_men_n181_));
  NAi21      u0153(.An(h), .B(f), .Y(men_men_n182_));
  NO2        u0154(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  NA2        u0155(.A(n), .B(men_men_n183_), .Y(men_men_n184_));
  NOi32      u0156(.An(f), .Bn(c), .C(d), .Y(men_men_n185_));
  NOi32      u0157(.An(f), .Bn(c), .C(e), .Y(men_men_n186_));
  NO3        u0158(.A(n), .B(m), .C(j), .Y(men_men_n187_));
  NA2        u0159(.A(men_men_n187_), .B(men_men_n109_), .Y(men_men_n188_));
  AO210      u0160(.A0(men_men_n188_), .A1(men_men_n174_), .B0(men_men_n1359_), .Y(men_men_n189_));
  NAi41      u0161(.An(men_men_n178_), .B(men_men_n189_), .C(men_men_n184_), .D(men_men_n172_), .Y(men_men_n190_));
  OR4        u0162(.A(men_men_n190_), .B(men_men_n163_), .C(men_men_n156_), .D(men_men_n149_), .Y(men_men_n191_));
  NO4        u0163(.A(men_men_n191_), .B(men_men_n119_), .C(men_men_n80_), .D(men_men_n54_), .Y(men_men_n192_));
  NA3        u0164(.A(m), .B(men_men_n107_), .C(j), .Y(men_men_n193_));
  NAi31      u0165(.An(n), .B(h), .C(u), .Y(men_men_n194_));
  NO2        u0166(.A(men_men_n194_), .B(men_men_n193_), .Y(men_men_n195_));
  NOi32      u0167(.An(m), .Bn(k), .C(l), .Y(men_men_n196_));
  NA3        u0168(.A(men_men_n196_), .B(men_men_n82_), .C(u), .Y(men_men_n197_));
  NO2        u0169(.A(men_men_n197_), .B(n), .Y(men_men_n198_));
  NOi21      u0170(.An(k), .B(j), .Y(men_men_n199_));
  NA4        u0171(.A(men_men_n199_), .B(men_men_n108_), .C(i), .D(u), .Y(men_men_n200_));
  AN2        u0172(.A(i), .B(u), .Y(men_men_n201_));
  NA3        u0173(.A(men_men_n75_), .B(men_men_n201_), .C(men_men_n108_), .Y(men_men_n202_));
  NA2        u0174(.A(men_men_n202_), .B(men_men_n200_), .Y(men_men_n203_));
  NO3        u0175(.A(men_men_n203_), .B(men_men_n198_), .C(men_men_n195_), .Y(men_men_n204_));
  NAi41      u0176(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n205_));
  INV        u0177(.A(men_men_n205_), .Y(men_men_n206_));
  INV        u0178(.A(f), .Y(men_men_n207_));
  INV        u0179(.A(u), .Y(men_men_n208_));
  NOi31      u0180(.An(i), .B(j), .C(h), .Y(men_men_n209_));
  NOi21      u0181(.An(l), .B(m), .Y(men_men_n210_));
  NA2        u0182(.A(men_men_n210_), .B(men_men_n209_), .Y(men_men_n211_));
  NO3        u0183(.A(men_men_n211_), .B(men_men_n208_), .C(men_men_n207_), .Y(men_men_n212_));
  NA2        u0184(.A(men_men_n212_), .B(men_men_n206_), .Y(men_men_n213_));
  OAI210     u0185(.A0(men_men_n204_), .A1(men_men_n31_), .B0(men_men_n213_), .Y(men_men_n214_));
  NOi21      u0186(.An(n), .B(m), .Y(men_men_n215_));
  NOi32      u0187(.An(l), .Bn(i), .C(j), .Y(men_men_n216_));
  NA2        u0188(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  OA220      u0189(.A0(men_men_n217_), .A1(men_men_n100_), .B0(k), .B1(men_men_n78_), .Y(men_men_n218_));
  NAi21      u0190(.An(j), .B(h), .Y(men_men_n219_));
  XN2        u0191(.A(i), .B(h), .Y(men_men_n220_));
  NOi31      u0192(.An(k), .B(n), .C(m), .Y(men_men_n221_));
  NAi31      u0193(.An(f), .B(e), .C(c), .Y(men_men_n222_));
  NA4        u0194(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n223_));
  NAi32      u0195(.An(m), .Bn(i), .C(k), .Y(men_men_n224_));
  NO3        u0196(.A(men_men_n224_), .B(men_men_n86_), .C(men_men_n223_), .Y(men_men_n225_));
  INV        u0197(.A(k), .Y(men_men_n226_));
  INV        u0198(.A(men_men_n225_), .Y(men_men_n227_));
  NAi21      u0199(.An(n), .B(a), .Y(men_men_n228_));
  NO2        u0200(.A(men_men_n228_), .B(men_men_n140_), .Y(men_men_n229_));
  NAi41      u0201(.An(u), .B(m), .C(k), .D(h), .Y(men_men_n230_));
  NO2        u0202(.A(men_men_n230_), .B(e), .Y(men_men_n231_));
  NO3        u0203(.A(men_men_n141_), .B(men_men_n90_), .C(men_men_n89_), .Y(men_men_n232_));
  OAI210     u0204(.A0(men_men_n232_), .A1(men_men_n231_), .B0(men_men_n229_), .Y(men_men_n233_));
  AN3        u0205(.A(men_men_n233_), .B(men_men_n227_), .C(men_men_n218_), .Y(men_men_n234_));
  NO2        u0206(.A(h), .B(men_men_n98_), .Y(men_men_n235_));
  NA2        u0207(.A(men_men_n235_), .B(men_men_n124_), .Y(men_men_n236_));
  NAi41      u0208(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n237_));
  NO2        u0209(.A(men_men_n237_), .B(men_men_n207_), .Y(men_men_n238_));
  NA2        u0210(.A(men_men_n154_), .B(men_men_n103_), .Y(men_men_n239_));
  NO2        u0211(.A(n), .B(a), .Y(men_men_n240_));
  NAi31      u0212(.An(men_men_n230_), .B(men_men_n240_), .C(men_men_n99_), .Y(men_men_n241_));
  NAi21      u0213(.An(h), .B(i), .Y(men_men_n242_));
  NA2        u0214(.A(men_men_n173_), .B(k), .Y(men_men_n243_));
  NO2        u0215(.A(men_men_n243_), .B(men_men_n242_), .Y(men_men_n244_));
  NA2        u0216(.A(men_men_n244_), .B(men_men_n185_), .Y(men_men_n245_));
  NA3        u0217(.A(men_men_n245_), .B(men_men_n241_), .C(men_men_n236_), .Y(men_men_n246_));
  NOi21      u0218(.An(u), .B(e), .Y(men_men_n247_));
  NO2        u0219(.A(men_men_n72_), .B(men_men_n74_), .Y(men_men_n248_));
  NA2        u0220(.A(men_men_n248_), .B(men_men_n247_), .Y(men_men_n249_));
  NOi32      u0221(.An(l), .Bn(j), .C(i), .Y(men_men_n250_));
  AOI210     u0222(.A0(men_men_n75_), .A1(men_men_n82_), .B0(men_men_n250_), .Y(men_men_n251_));
  NO2        u0223(.A(men_men_n242_), .B(men_men_n43_), .Y(men_men_n252_));
  NAi21      u0224(.An(f), .B(u), .Y(men_men_n253_));
  NO2        u0225(.A(men_men_n253_), .B(men_men_n64_), .Y(men_men_n254_));
  NO2        u0226(.A(men_men_n68_), .B(men_men_n111_), .Y(men_men_n255_));
  AOI220     u0227(.A0(men_men_n255_), .A1(men_men_n254_), .B0(men_men_n252_), .B1(men_men_n66_), .Y(men_men_n256_));
  OAI210     u0228(.A0(men_men_n251_), .A1(men_men_n249_), .B0(men_men_n256_), .Y(men_men_n257_));
  NOi41      u0229(.An(men_men_n234_), .B(men_men_n257_), .C(men_men_n246_), .D(men_men_n214_), .Y(men_men_n258_));
  NO4        u0230(.A(men_men_n195_), .B(men_men_n47_), .C(men_men_n42_), .D(men_men_n38_), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n259_), .B(men_men_n106_), .Y(men_men_n260_));
  NA3        u0232(.A(men_men_n58_), .B(c), .C(b), .Y(men_men_n261_));
  NAi21      u0233(.An(h), .B(u), .Y(men_men_n262_));
  OR4        u0234(.A(men_men_n262_), .B(men_men_n261_), .C(men_men_n217_), .D(e), .Y(men_men_n263_));
  NO2        u0235(.A(men_men_n239_), .B(men_men_n253_), .Y(men_men_n264_));
  NA2        u0236(.A(men_men_n264_), .B(men_men_n77_), .Y(men_men_n265_));
  NAi31      u0237(.An(u), .B(k), .C(h), .Y(men_men_n266_));
  NO3        u0238(.A(men_men_n126_), .B(men_men_n266_), .C(l), .Y(men_men_n267_));
  NAi31      u0239(.An(e), .B(d), .C(a), .Y(men_men_n268_));
  NA2        u0240(.A(men_men_n267_), .B(men_men_n124_), .Y(men_men_n269_));
  NA3        u0241(.A(men_men_n269_), .B(men_men_n265_), .C(men_men_n263_), .Y(men_men_n270_));
  NA4        u0242(.A(men_men_n154_), .B(men_men_n79_), .C(men_men_n77_), .D(men_men_n111_), .Y(men_men_n271_));
  NA3        u0243(.A(men_men_n154_), .B(men_men_n153_), .C(men_men_n81_), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n272_), .B(men_men_n1359_), .Y(men_men_n273_));
  NOi21      u0245(.An(men_men_n271_), .B(men_men_n273_), .Y(men_men_n274_));
  NA3        u0246(.A(e), .B(c), .C(b), .Y(men_men_n275_));
  NO2        u0247(.A(men_men_n59_), .B(men_men_n275_), .Y(men_men_n276_));
  NAi32      u0248(.An(k), .Bn(i), .C(j), .Y(men_men_n277_));
  NAi31      u0249(.An(h), .B(l), .C(i), .Y(men_men_n278_));
  NA3        u0250(.A(men_men_n278_), .B(men_men_n277_), .C(men_men_n159_), .Y(men_men_n279_));
  NOi21      u0251(.An(men_men_n279_), .B(men_men_n48_), .Y(men_men_n280_));
  OAI210     u0252(.A0(men_men_n254_), .A1(men_men_n276_), .B0(men_men_n280_), .Y(men_men_n281_));
  NAi21      u0253(.An(l), .B(k), .Y(men_men_n282_));
  NO2        u0254(.A(men_men_n282_), .B(men_men_n48_), .Y(men_men_n283_));
  NOi21      u0255(.An(l), .B(j), .Y(men_men_n284_));
  NA2        u0256(.A(men_men_n157_), .B(men_men_n284_), .Y(men_men_n285_));
  NA3        u0257(.A(men_men_n112_), .B(men_men_n111_), .C(u), .Y(men_men_n286_));
  OR3        u0258(.A(men_men_n72_), .B(men_men_n74_), .C(e), .Y(men_men_n287_));
  AOI210     u0259(.A0(men_men_n286_), .A1(men_men_n285_), .B0(men_men_n287_), .Y(men_men_n288_));
  INV        u0260(.A(men_men_n288_), .Y(men_men_n289_));
  NAi32      u0261(.An(j), .Bn(h), .C(i), .Y(men_men_n290_));
  NAi21      u0262(.An(m), .B(l), .Y(men_men_n291_));
  NO3        u0263(.A(men_men_n291_), .B(men_men_n290_), .C(men_men_n81_), .Y(men_men_n292_));
  NA2        u0264(.A(h), .B(u), .Y(men_men_n293_));
  NO2        u0265(.A(men_men_n1356_), .B(men_men_n293_), .Y(men_men_n294_));
  OAI210     u0266(.A0(men_men_n294_), .A1(men_men_n292_), .B0(men_men_n158_), .Y(men_men_n295_));
  NA4        u0267(.A(men_men_n295_), .B(men_men_n289_), .C(men_men_n281_), .D(men_men_n274_), .Y(men_men_n296_));
  NO2        u0268(.A(men_men_n100_), .B(men_men_n98_), .Y(men_men_n297_));
  NAi32      u0269(.An(n), .Bn(m), .C(l), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n298_), .B(men_men_n290_), .Y(men_men_n299_));
  NA2        u0271(.A(men_men_n299_), .B(men_men_n177_), .Y(men_men_n300_));
  NO2        u0272(.A(men_men_n116_), .B(men_men_n110_), .Y(men_men_n301_));
  NAi31      u0273(.An(k), .B(l), .C(j), .Y(men_men_n302_));
  OAI210     u0274(.A0(men_men_n282_), .A1(j), .B0(men_men_n302_), .Y(men_men_n303_));
  NOi21      u0275(.An(men_men_n303_), .B(men_men_n114_), .Y(men_men_n304_));
  NA2        u0276(.A(men_men_n304_), .B(men_men_n301_), .Y(men_men_n305_));
  NA2        u0277(.A(men_men_n305_), .B(men_men_n300_), .Y(men_men_n306_));
  NO4        u0278(.A(men_men_n306_), .B(men_men_n296_), .C(men_men_n270_), .D(men_men_n260_), .Y(men_men_n307_));
  NAi21      u0279(.An(m), .B(k), .Y(men_men_n308_));
  NO2        u0280(.A(men_men_n220_), .B(men_men_n308_), .Y(men_men_n309_));
  NAi41      u0281(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n310_));
  NO2        u0282(.A(men_men_n310_), .B(men_men_n144_), .Y(men_men_n311_));
  NA2        u0283(.A(men_men_n311_), .B(men_men_n309_), .Y(men_men_n312_));
  NAi31      u0284(.An(i), .B(l), .C(h), .Y(men_men_n313_));
  NO4        u0285(.A(men_men_n313_), .B(men_men_n144_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n314_));
  NA2        u0286(.A(e), .B(c), .Y(men_men_n315_));
  NO3        u0287(.A(men_men_n315_), .B(n), .C(d), .Y(men_men_n316_));
  NOi21      u0288(.An(f), .B(h), .Y(men_men_n317_));
  NA2        u0289(.A(men_men_n317_), .B(men_men_n112_), .Y(men_men_n318_));
  NO2        u0290(.A(men_men_n318_), .B(men_men_n208_), .Y(men_men_n319_));
  NAi31      u0291(.An(d), .B(e), .C(b), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n126_), .B(men_men_n320_), .Y(men_men_n321_));
  NA2        u0293(.A(men_men_n321_), .B(men_men_n319_), .Y(men_men_n322_));
  NAi31      u0294(.An(men_men_n314_), .B(men_men_n322_), .C(men_men_n312_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n240_), .B(men_men_n99_), .Y(men_men_n324_));
  OR2        u0296(.A(men_men_n324_), .B(men_men_n197_), .Y(men_men_n325_));
  NOi31      u0297(.An(l), .B(n), .C(m), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n326_), .B(men_men_n209_), .Y(men_men_n327_));
  NO2        u0299(.A(men_men_n327_), .B(men_men_n1359_), .Y(men_men_n328_));
  NAi21      u0300(.An(men_men_n328_), .B(men_men_n325_), .Y(men_men_n329_));
  NAi32      u0301(.An(m), .Bn(j), .C(k), .Y(men_men_n330_));
  NAi41      u0302(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n331_));
  NOi31      u0303(.An(j), .B(m), .C(k), .Y(men_men_n332_));
  INV        u0304(.A(men_men_n120_), .Y(men_men_n333_));
  AN3        u0305(.A(h), .B(u), .C(f), .Y(men_men_n334_));
  NOi32      u0306(.An(m), .Bn(j), .C(l), .Y(men_men_n335_));
  NO2        u0307(.A(men_men_n335_), .B(men_men_n93_), .Y(men_men_n336_));
  NO2        u0308(.A(men_men_n291_), .B(men_men_n290_), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n211_), .B(u), .Y(men_men_n338_));
  AOI220     u0310(.A0(f), .A1(men_men_n338_), .B0(men_men_n238_), .B1(men_men_n337_), .Y(men_men_n339_));
  NA2        u0311(.A(men_men_n334_), .B(men_men_n206_), .Y(men_men_n340_));
  NA2        u0312(.A(men_men_n340_), .B(men_men_n339_), .Y(men_men_n341_));
  NA3        u0313(.A(h), .B(u), .C(f), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n342_), .B(men_men_n76_), .Y(men_men_n343_));
  NA2        u0315(.A(men_men_n157_), .B(e), .Y(men_men_n344_));
  NO2        u0316(.A(men_men_n344_), .B(men_men_n40_), .Y(men_men_n345_));
  NA2        u0317(.A(men_men_n345_), .B(men_men_n301_), .Y(men_men_n346_));
  NOi32      u0318(.An(j), .Bn(u), .C(i), .Y(men_men_n347_));
  NA3        u0319(.A(men_men_n347_), .B(men_men_n282_), .C(men_men_n108_), .Y(men_men_n348_));
  AO210      u0320(.A0(men_men_n106_), .A1(men_men_n31_), .B0(men_men_n348_), .Y(men_men_n349_));
  NOi32      u0321(.An(e), .Bn(b), .C(a), .Y(men_men_n350_));
  AN2        u0322(.A(l), .B(j), .Y(men_men_n351_));
  NO3        u0323(.A(men_men_n310_), .B(men_men_n71_), .C(men_men_n208_), .Y(men_men_n352_));
  NA3        u0324(.A(men_men_n202_), .B(men_men_n200_), .C(men_men_n34_), .Y(men_men_n353_));
  AOI210     u0325(.A0(men_men_n353_), .A1(men_men_n350_), .B0(men_men_n352_), .Y(men_men_n354_));
  NA2        u0326(.A(men_men_n201_), .B(k), .Y(men_men_n355_));
  NA3        u0327(.A(m), .B(men_men_n107_), .C(men_men_n207_), .Y(men_men_n356_));
  NA4        u0328(.A(men_men_n196_), .B(men_men_n82_), .C(u), .D(men_men_n207_), .Y(men_men_n357_));
  NAi41      u0329(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n358_));
  NA2        u0330(.A(men_men_n50_), .B(men_men_n108_), .Y(men_men_n359_));
  NO2        u0331(.A(men_men_n359_), .B(men_men_n358_), .Y(men_men_n360_));
  INV        u0332(.A(men_men_n360_), .Y(men_men_n361_));
  NA4        u0333(.A(men_men_n361_), .B(men_men_n354_), .C(men_men_n349_), .D(men_men_n346_), .Y(men_men_n362_));
  NO4        u0334(.A(men_men_n362_), .B(men_men_n341_), .C(men_men_n329_), .D(men_men_n323_), .Y(men_men_n363_));
  NA4        u0335(.A(men_men_n363_), .B(men_men_n307_), .C(men_men_n258_), .D(men_men_n192_), .Y(men10));
  NA3        u0336(.A(m), .B(k), .C(i), .Y(men_men_n365_));
  NO3        u0337(.A(men_men_n365_), .B(j), .C(men_men_n208_), .Y(men_men_n366_));
  NOi21      u0338(.An(e), .B(f), .Y(men_men_n367_));
  NO4        u0339(.A(men_men_n145_), .B(men_men_n367_), .C(n), .D(men_men_n105_), .Y(men_men_n368_));
  NAi31      u0340(.An(b), .B(f), .C(c), .Y(men_men_n369_));
  INV        u0341(.A(men_men_n369_), .Y(men_men_n370_));
  NA2        u0342(.A(h), .B(men_men_n215_), .Y(men_men_n371_));
  INV        u0343(.A(men_men_n371_), .Y(men_men_n372_));
  AOI220     u0344(.A0(men_men_n372_), .A1(men_men_n370_), .B0(men_men_n368_), .B1(men_men_n366_), .Y(men_men_n373_));
  AN2        u0345(.A(j), .B(h), .Y(men_men_n374_));
  NO3        u0346(.A(n), .B(m), .C(k), .Y(men_men_n375_));
  NA2        u0347(.A(men_men_n375_), .B(men_men_n374_), .Y(men_men_n376_));
  NO3        u0348(.A(men_men_n376_), .B(men_men_n145_), .C(men_men_n207_), .Y(men_men_n377_));
  OR2        u0349(.A(m), .B(k), .Y(men_men_n378_));
  NO2        u0350(.A(men_men_n167_), .B(men_men_n378_), .Y(men_men_n379_));
  NA4        u0351(.A(n), .B(f), .C(c), .D(men_men_n110_), .Y(men_men_n380_));
  NOi32      u0352(.An(d), .Bn(a), .C(c), .Y(men_men_n381_));
  NA2        u0353(.A(men_men_n381_), .B(men_men_n175_), .Y(men_men_n382_));
  NAi21      u0354(.An(i), .B(u), .Y(men_men_n383_));
  NAi31      u0355(.An(k), .B(m), .C(j), .Y(men_men_n384_));
  NO3        u0356(.A(men_men_n384_), .B(men_men_n383_), .C(n), .Y(men_men_n385_));
  NOi21      u0357(.An(men_men_n385_), .B(men_men_n382_), .Y(men_men_n386_));
  NO2        u0358(.A(men_men_n386_), .B(men_men_n377_), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n380_), .B(men_men_n291_), .Y(men_men_n388_));
  NOi32      u0360(.An(f), .Bn(d), .C(c), .Y(men_men_n389_));
  NA2        u0361(.A(men_men_n388_), .B(men_men_n209_), .Y(men_men_n390_));
  NA3        u0362(.A(men_men_n390_), .B(men_men_n387_), .C(men_men_n373_), .Y(men_men_n391_));
  NO2        u0363(.A(men_men_n58_), .B(men_men_n110_), .Y(men_men_n392_));
  NA2        u0364(.A(men_men_n240_), .B(men_men_n392_), .Y(men_men_n393_));
  INV        u0365(.A(e), .Y(men_men_n394_));
  NA2        u0366(.A(men_men_n45_), .B(e), .Y(men_men_n395_));
  OAI220     u0367(.A0(men_men_n395_), .A1(men_men_n193_), .B0(men_men_n197_), .B1(men_men_n394_), .Y(men_men_n396_));
  AN2        u0368(.A(u), .B(e), .Y(men_men_n397_));
  NA3        u0369(.A(men_men_n397_), .B(men_men_n196_), .C(i), .Y(men_men_n398_));
  OAI210     u0370(.A0(men_men_n84_), .A1(men_men_n394_), .B0(men_men_n398_), .Y(men_men_n399_));
  NO2        u0371(.A(men_men_n96_), .B(men_men_n394_), .Y(men_men_n400_));
  NO3        u0372(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n396_), .Y(men_men_n401_));
  NOi32      u0373(.An(h), .Bn(e), .C(u), .Y(men_men_n402_));
  NA3        u0374(.A(men_men_n402_), .B(men_men_n284_), .C(m), .Y(men_men_n403_));
  NOi21      u0375(.An(u), .B(h), .Y(men_men_n404_));
  AN3        u0376(.A(m), .B(l), .C(i), .Y(men_men_n405_));
  NA3        u0377(.A(men_men_n405_), .B(men_men_n404_), .C(e), .Y(men_men_n406_));
  AN3        u0378(.A(h), .B(u), .C(e), .Y(men_men_n407_));
  NA2        u0379(.A(men_men_n407_), .B(men_men_n93_), .Y(men_men_n408_));
  AN3        u0380(.A(men_men_n408_), .B(men_men_n406_), .C(men_men_n403_), .Y(men_men_n409_));
  AOI210     u0381(.A0(men_men_n409_), .A1(men_men_n401_), .B0(men_men_n393_), .Y(men_men_n410_));
  NA3        u0382(.A(men_men_n36_), .B(men_men_n35_), .C(e), .Y(men_men_n411_));
  NO2        u0383(.A(men_men_n411_), .B(men_men_n393_), .Y(men_men_n412_));
  NA2        u0384(.A(men_men_n381_), .B(men_men_n175_), .Y(men_men_n413_));
  NAi31      u0385(.An(b), .B(c), .C(a), .Y(men_men_n414_));
  NO2        u0386(.A(men_men_n414_), .B(n), .Y(men_men_n415_));
  OAI210     u0387(.A0(men_men_n50_), .A1(men_men_n49_), .B0(m), .Y(men_men_n416_));
  NO2        u0388(.A(men_men_n416_), .B(men_men_n141_), .Y(men_men_n417_));
  NA2        u0389(.A(men_men_n417_), .B(men_men_n415_), .Y(men_men_n418_));
  INV        u0390(.A(men_men_n418_), .Y(men_men_n419_));
  NO4        u0391(.A(men_men_n419_), .B(men_men_n412_), .C(men_men_n410_), .D(men_men_n391_), .Y(men_men_n420_));
  NA2        u0392(.A(i), .B(u), .Y(men_men_n421_));
  NO3        u0393(.A(men_men_n268_), .B(men_men_n421_), .C(c), .Y(men_men_n422_));
  NOi21      u0394(.An(d), .B(c), .Y(men_men_n423_));
  NA2        u0395(.A(men_men_n423_), .B(a), .Y(men_men_n424_));
  NA3        u0396(.A(i), .B(u), .C(f), .Y(men_men_n425_));
  OR2        u0397(.A(men_men_n425_), .B(men_men_n70_), .Y(men_men_n426_));
  NA3        u0398(.A(men_men_n405_), .B(men_men_n404_), .C(men_men_n175_), .Y(men_men_n427_));
  AOI210     u0399(.A0(men_men_n427_), .A1(men_men_n426_), .B0(men_men_n424_), .Y(men_men_n428_));
  AOI210     u0400(.A0(men_men_n422_), .A1(men_men_n283_), .B0(men_men_n428_), .Y(men_men_n429_));
  OR2        u0401(.A(n), .B(m), .Y(men_men_n430_));
  NO2        u0402(.A(men_men_n430_), .B(men_men_n146_), .Y(men_men_n431_));
  NO2        u0403(.A(men_men_n176_), .B(men_men_n141_), .Y(men_men_n432_));
  OAI210     u0404(.A0(men_men_n431_), .A1(men_men_n169_), .B0(men_men_n432_), .Y(men_men_n433_));
  INV        u0405(.A(men_men_n359_), .Y(men_men_n434_));
  NA3        u0406(.A(men_men_n434_), .B(men_men_n350_), .C(d), .Y(men_men_n435_));
  NO2        u0407(.A(men_men_n414_), .B(men_men_n48_), .Y(men_men_n436_));
  NO3        u0408(.A(men_men_n65_), .B(men_men_n107_), .C(e), .Y(men_men_n437_));
  NAi21      u0409(.An(k), .B(j), .Y(men_men_n438_));
  NA2        u0410(.A(men_men_n242_), .B(men_men_n438_), .Y(men_men_n439_));
  NA3        u0411(.A(men_men_n439_), .B(men_men_n437_), .C(men_men_n436_), .Y(men_men_n440_));
  NAi21      u0412(.An(e), .B(d), .Y(men_men_n441_));
  NO2        u0413(.A(men_men_n243_), .B(men_men_n207_), .Y(men_men_n442_));
  NA3        u0414(.A(men_men_n440_), .B(men_men_n435_), .C(men_men_n433_), .Y(men_men_n443_));
  NO2        u0415(.A(men_men_n327_), .B(men_men_n207_), .Y(men_men_n444_));
  NA2        u0416(.A(men_men_n444_), .B(d), .Y(men_men_n445_));
  NA2        u0417(.A(n), .B(men_men_n374_), .Y(men_men_n446_));
  NAi31      u0418(.An(u), .B(f), .C(c), .Y(men_men_n447_));
  OR3        u0419(.A(men_men_n447_), .B(men_men_n446_), .C(e), .Y(men_men_n448_));
  NA3        u0420(.A(men_men_n448_), .B(men_men_n445_), .C(men_men_n300_), .Y(men_men_n449_));
  NOi41      u0421(.An(men_men_n429_), .B(men_men_n449_), .C(men_men_n443_), .D(men_men_n257_), .Y(men_men_n450_));
  NOi32      u0422(.An(c), .Bn(a), .C(b), .Y(men_men_n451_));
  NA2        u0423(.A(men_men_n451_), .B(men_men_n108_), .Y(men_men_n452_));
  INV        u0424(.A(men_men_n266_), .Y(men_men_n453_));
  AN2        u0425(.A(e), .B(d), .Y(men_men_n454_));
  NA2        u0426(.A(men_men_n454_), .B(men_men_n453_), .Y(men_men_n455_));
  INV        u0427(.A(men_men_n141_), .Y(men_men_n456_));
  NO2        u0428(.A(men_men_n125_), .B(men_men_n40_), .Y(men_men_n457_));
  NO2        u0429(.A(men_men_n65_), .B(e), .Y(men_men_n458_));
  NOi31      u0430(.An(j), .B(k), .C(i), .Y(men_men_n459_));
  NOi21      u0431(.An(men_men_n159_), .B(men_men_n459_), .Y(men_men_n460_));
  NA4        u0432(.A(men_men_n313_), .B(men_men_n460_), .C(men_men_n251_), .D(men_men_n113_), .Y(men_men_n461_));
  AOI220     u0433(.A0(men_men_n461_), .A1(men_men_n458_), .B0(men_men_n457_), .B1(men_men_n456_), .Y(men_men_n462_));
  AOI210     u0434(.A0(men_men_n462_), .A1(men_men_n455_), .B0(men_men_n452_), .Y(men_men_n463_));
  NO2        u0435(.A(men_men_n203_), .B(men_men_n198_), .Y(men_men_n464_));
  NOi21      u0436(.An(a), .B(b), .Y(men_men_n465_));
  NA3        u0437(.A(e), .B(d), .C(c), .Y(men_men_n466_));
  NAi21      u0438(.An(men_men_n466_), .B(men_men_n465_), .Y(men_men_n467_));
  NO2        u0439(.A(men_men_n413_), .B(men_men_n197_), .Y(men_men_n468_));
  NOi21      u0440(.An(men_men_n467_), .B(men_men_n468_), .Y(men_men_n469_));
  AOI210     u0441(.A0(men_men_n259_), .A1(men_men_n464_), .B0(men_men_n469_), .Y(men_men_n470_));
  NO3        u0442(.A(men_men_n182_), .B(men_men_n98_), .C(men_men_n55_), .Y(men_men_n471_));
  OR2        u0443(.A(k), .B(j), .Y(men_men_n472_));
  NA2        u0444(.A(l), .B(k), .Y(men_men_n473_));
  NA2        u0445(.A(men_men_n224_), .B(men_men_n330_), .Y(men_men_n474_));
  OR3        u0446(.A(men_men_n1353_), .B(men_men_n137_), .C(men_men_n128_), .Y(men_men_n475_));
  NA2        u0447(.A(men_men_n271_), .B(men_men_n122_), .Y(men_men_n476_));
  NA2        u0448(.A(men_men_n381_), .B(men_men_n108_), .Y(men_men_n477_));
  NO4        u0449(.A(men_men_n477_), .B(men_men_n90_), .C(men_men_n107_), .D(e), .Y(men_men_n478_));
  NO3        u0450(.A(men_men_n413_), .B(men_men_n87_), .C(men_men_n125_), .Y(men_men_n479_));
  NO4        u0451(.A(men_men_n479_), .B(men_men_n478_), .C(men_men_n476_), .D(men_men_n314_), .Y(men_men_n480_));
  NA2        u0452(.A(men_men_n480_), .B(men_men_n475_), .Y(men_men_n481_));
  NO4        u0453(.A(men_men_n481_), .B(men_men_n471_), .C(men_men_n470_), .D(men_men_n463_), .Y(men_men_n482_));
  NA2        u0454(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n483_));
  NAi31      u0455(.An(j), .B(l), .C(i), .Y(men_men_n484_));
  OAI210     u0456(.A0(men_men_n484_), .A1(men_men_n126_), .B0(men_men_n98_), .Y(men_men_n485_));
  NO3        u0457(.A(men_men_n382_), .B(men_men_n336_), .C(men_men_n194_), .Y(men_men_n486_));
  NO2        u0458(.A(men_men_n382_), .B(men_men_n359_), .Y(men_men_n487_));
  NO4        u0459(.A(men_men_n487_), .B(men_men_n486_), .C(men_men_n178_), .D(men_men_n297_), .Y(men_men_n488_));
  NA3        u0460(.A(men_men_n488_), .B(men_men_n483_), .C(men_men_n234_), .Y(men_men_n489_));
  OAI210     u0461(.A0(men_men_n121_), .A1(men_men_n120_), .B0(n), .Y(men_men_n490_));
  NO2        u0462(.A(men_men_n490_), .B(men_men_n125_), .Y(men_men_n491_));
  BUFFER     u0463(.A(men_men_n292_), .Y(men_men_n492_));
  OA210      u0464(.A0(men_men_n492_), .A1(men_men_n491_), .B0(men_men_n186_), .Y(men_men_n493_));
  XO2        u0465(.A(i), .B(h), .Y(men_men_n494_));
  NA3        u0466(.A(men_men_n494_), .B(men_men_n154_), .C(n), .Y(men_men_n495_));
  NAi31      u0467(.An(men_men_n292_), .B(men_men_n495_), .C(men_men_n371_), .Y(men_men_n496_));
  NOi32      u0468(.An(men_men_n496_), .Bn(men_men_n458_), .C(men_men_n261_), .Y(men_men_n497_));
  NAi31      u0469(.An(c), .B(f), .C(d), .Y(men_men_n498_));
  AOI210     u0470(.A0(men_men_n272_), .A1(men_men_n188_), .B0(men_men_n498_), .Y(men_men_n499_));
  INV        u0471(.A(men_men_n499_), .Y(men_men_n500_));
  NA3        u0472(.A(men_men_n368_), .B(men_men_n93_), .C(men_men_n92_), .Y(men_men_n501_));
  NA2        u0473(.A(men_men_n221_), .B(men_men_n103_), .Y(men_men_n502_));
  AOI210     u0474(.A0(men_men_n502_), .A1(men_men_n174_), .B0(men_men_n498_), .Y(men_men_n503_));
  AOI210     u0475(.A0(men_men_n348_), .A1(men_men_n34_), .B0(men_men_n467_), .Y(men_men_n504_));
  NOi31      u0476(.An(men_men_n501_), .B(men_men_n504_), .C(men_men_n503_), .Y(men_men_n505_));
  AO220      u0477(.A0(men_men_n280_), .A1(men_men_n254_), .B0(men_men_n160_), .B1(men_men_n66_), .Y(men_men_n506_));
  NA3        u0478(.A(men_men_n36_), .B(men_men_n35_), .C(f), .Y(men_men_n507_));
  NO2        u0479(.A(men_men_n507_), .B(men_men_n424_), .Y(men_men_n508_));
  NO2        u0480(.A(men_men_n508_), .B(men_men_n288_), .Y(men_men_n509_));
  NAi41      u0481(.An(men_men_n506_), .B(men_men_n509_), .C(men_men_n505_), .D(men_men_n500_), .Y(men_men_n510_));
  NO4        u0482(.A(men_men_n510_), .B(men_men_n497_), .C(men_men_n493_), .D(men_men_n489_), .Y(men_men_n511_));
  NA4        u0483(.A(men_men_n511_), .B(men_men_n482_), .C(men_men_n450_), .D(men_men_n420_), .Y(men11));
  NO2        u0484(.A(men_men_n72_), .B(f), .Y(men_men_n513_));
  NA2        u0485(.A(j), .B(u), .Y(men_men_n514_));
  NAi31      u0486(.An(i), .B(m), .C(l), .Y(men_men_n515_));
  NA3        u0487(.A(m), .B(k), .C(j), .Y(men_men_n516_));
  OAI220     u0488(.A0(men_men_n516_), .A1(men_men_n125_), .B0(men_men_n515_), .B1(men_men_n514_), .Y(men_men_n517_));
  NA2        u0489(.A(men_men_n517_), .B(men_men_n513_), .Y(men_men_n518_));
  NOi32      u0490(.An(e), .Bn(b), .C(f), .Y(men_men_n519_));
  NA2        u0491(.A(men_men_n250_), .B(men_men_n108_), .Y(men_men_n520_));
  NA2        u0492(.A(men_men_n45_), .B(j), .Y(men_men_n521_));
  NO2        u0493(.A(men_men_n521_), .B(men_men_n1356_), .Y(men_men_n522_));
  NAi31      u0494(.An(d), .B(e), .C(a), .Y(men_men_n523_));
  NO2        u0495(.A(men_men_n523_), .B(n), .Y(men_men_n524_));
  NA2        u0496(.A(men_men_n522_), .B(men_men_n519_), .Y(men_men_n525_));
  NAi41      u0497(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n526_));
  BUFFER     u0498(.A(men_men_n526_), .Y(men_men_n527_));
  AOI210     u0499(.A0(men_men_n527_), .A1(men_men_n382_), .B0(men_men_n262_), .Y(men_men_n528_));
  NA2        u0500(.A(j), .B(i), .Y(men_men_n529_));
  NAi31      u0501(.An(n), .B(m), .C(k), .Y(men_men_n530_));
  NO3        u0502(.A(men_men_n530_), .B(men_men_n529_), .C(men_men_n107_), .Y(men_men_n531_));
  NO2        u0503(.A(c), .B(men_men_n143_), .Y(men_men_n532_));
  NOi32      u0504(.An(u), .Bn(f), .C(i), .Y(men_men_n533_));
  NA2        u0505(.A(men_men_n517_), .B(f), .Y(men_men_n534_));
  NO2        u0506(.A(men_men_n266_), .B(men_men_n48_), .Y(men_men_n535_));
  NO2        u0507(.A(men_men_n534_), .B(n), .Y(men_men_n536_));
  AOI210     u0508(.A0(men_men_n531_), .A1(men_men_n528_), .B0(men_men_n536_), .Y(men_men_n537_));
  NA2        u0509(.A(men_men_n133_), .B(men_men_n33_), .Y(men_men_n538_));
  OAI220     u0510(.A0(men_men_n538_), .A1(m), .B0(men_men_n521_), .B1(men_men_n224_), .Y(men_men_n539_));
  NOi41      u0511(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n540_));
  NAi32      u0512(.An(e), .Bn(b), .C(c), .Y(men_men_n541_));
  AN2        u0513(.A(men_men_n331_), .B(men_men_n310_), .Y(men_men_n542_));
  NA2        u0514(.A(men_men_n542_), .B(men_men_n541_), .Y(men_men_n543_));
  AN2        u0515(.A(men_men_n543_), .B(men_men_n539_), .Y(men_men_n544_));
  OAI220     u0516(.A0(men_men_n384_), .A1(men_men_n383_), .B0(men_men_n515_), .B1(men_men_n514_), .Y(men_men_n545_));
  NAi31      u0517(.An(d), .B(c), .C(a), .Y(men_men_n546_));
  NO2        u0518(.A(men_men_n546_), .B(n), .Y(men_men_n547_));
  NA3        u0519(.A(men_men_n547_), .B(men_men_n545_), .C(e), .Y(men_men_n548_));
  NO3        u0520(.A(men_men_n61_), .B(men_men_n48_), .C(men_men_n208_), .Y(men_men_n549_));
  OAI210     u0521(.A0(men_men_n549_), .A1(men_men_n385_), .B0(e), .Y(men_men_n550_));
  NA2        u0522(.A(men_men_n550_), .B(men_men_n548_), .Y(men_men_n551_));
  NA2        u0523(.A(men_men_n545_), .B(f), .Y(men_men_n552_));
  NA2        u0524(.A(h), .B(f), .Y(men_men_n553_));
  NO2        u0525(.A(men_men_n553_), .B(men_men_n90_), .Y(men_men_n554_));
  NO3        u0526(.A(men_men_n170_), .B(men_men_n167_), .C(u), .Y(men_men_n555_));
  AOI220     u0527(.A0(men_men_n555_), .A1(men_men_n57_), .B0(men_men_n554_), .B1(m), .Y(men_men_n556_));
  OAI210     u0528(.A0(men_men_n552_), .A1(n), .B0(men_men_n556_), .Y(men_men_n557_));
  AN3        u0529(.A(j), .B(h), .C(u), .Y(men_men_n558_));
  NA3        u0530(.A(f), .B(d), .C(b), .Y(men_men_n559_));
  NO4        u0531(.A(men_men_n559_), .B(men_men_n170_), .C(men_men_n167_), .D(u), .Y(men_men_n560_));
  NO4        u0532(.A(men_men_n560_), .B(men_men_n557_), .C(men_men_n551_), .D(men_men_n544_), .Y(men_men_n561_));
  AN4        u0533(.A(men_men_n561_), .B(men_men_n537_), .C(men_men_n525_), .D(men_men_n518_), .Y(men_men_n562_));
  INV        u0534(.A(k), .Y(men_men_n563_));
  NA3        u0535(.A(l), .B(men_men_n563_), .C(i), .Y(men_men_n564_));
  INV        u0536(.A(men_men_n564_), .Y(men_men_n565_));
  NA4        u0537(.A(men_men_n381_), .B(men_men_n404_), .C(men_men_n175_), .D(men_men_n108_), .Y(men_men_n566_));
  NAi32      u0538(.An(h), .Bn(f), .C(u), .Y(men_men_n567_));
  NAi41      u0539(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n568_));
  OAI210     u0540(.A0(men_men_n523_), .A1(n), .B0(men_men_n568_), .Y(men_men_n569_));
  NA2        u0541(.A(men_men_n569_), .B(m), .Y(men_men_n570_));
  NAi31      u0542(.An(h), .B(u), .C(f), .Y(men_men_n571_));
  OR2        u0543(.A(men_men_n570_), .B(men_men_n567_), .Y(men_men_n572_));
  NO3        u0544(.A(men_men_n567_), .B(men_men_n72_), .C(men_men_n74_), .Y(men_men_n573_));
  NAi31      u0545(.An(men_men_n573_), .B(men_men_n572_), .C(men_men_n566_), .Y(men_men_n574_));
  NAi31      u0546(.An(f), .B(h), .C(u), .Y(men_men_n575_));
  NO4        u0547(.A(men_men_n302_), .B(men_men_n575_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n576_));
  NOi32      u0548(.An(b), .Bn(a), .C(c), .Y(men_men_n577_));
  NOi32      u0549(.An(d), .Bn(a), .C(e), .Y(men_men_n578_));
  NO2        u0550(.A(n), .B(c), .Y(men_men_n579_));
  NOi32      u0551(.An(e), .Bn(a), .C(d), .Y(men_men_n580_));
  AOI210     u0552(.A0(men_men_n29_), .A1(d), .B0(men_men_n580_), .Y(men_men_n581_));
  AOI210     u0553(.A0(men_men_n581_), .A1(men_men_n207_), .B0(men_men_n538_), .Y(men_men_n582_));
  AOI210     u0554(.A0(men_men_n582_), .A1(men_men_n108_), .B0(men_men_n576_), .Y(men_men_n583_));
  INV        u0555(.A(men_men_n583_), .Y(men_men_n584_));
  AOI210     u0556(.A0(men_men_n574_), .A1(men_men_n565_), .B0(men_men_n584_), .Y(men_men_n585_));
  NO3        u0557(.A(men_men_n308_), .B(men_men_n60_), .C(n), .Y(men_men_n586_));
  NA3        u0558(.A(men_men_n498_), .B(men_men_n165_), .C(men_men_n164_), .Y(men_men_n587_));
  NA2        u0559(.A(men_men_n447_), .B(men_men_n222_), .Y(men_men_n588_));
  NA2        u0560(.A(men_men_n75_), .B(men_men_n108_), .Y(men_men_n589_));
  NO2        u0561(.A(men_men_n589_), .B(men_men_n44_), .Y(men_men_n590_));
  AOI210     u0562(.A0(men_men_n590_), .A1(men_men_n528_), .B0(men_men_n586_), .Y(men_men_n591_));
  NO2        u0563(.A(men_men_n591_), .B(men_men_n82_), .Y(men_men_n592_));
  NA3        u0564(.A(men_men_n540_), .B(men_men_n332_), .C(men_men_n45_), .Y(men_men_n593_));
  NOi32      u0565(.An(e), .Bn(c), .C(f), .Y(men_men_n594_));
  INV        u0566(.A(men_men_n205_), .Y(men_men_n595_));
  AOI220     u0567(.A0(men_men_n595_), .A1(men_men_n379_), .B0(men_men_n594_), .B1(men_men_n169_), .Y(men_men_n596_));
  NA3        u0568(.A(men_men_n596_), .B(men_men_n593_), .C(men_men_n172_), .Y(men_men_n597_));
  AOI210     u0569(.A0(men_men_n527_), .A1(men_men_n382_), .B0(men_men_n293_), .Y(men_men_n598_));
  NA2        u0570(.A(men_men_n598_), .B(men_men_n255_), .Y(men_men_n599_));
  NOi21      u0571(.An(j), .B(l), .Y(men_men_n600_));
  NAi21      u0572(.An(k), .B(h), .Y(men_men_n601_));
  NO2        u0573(.A(men_men_n601_), .B(men_men_n253_), .Y(men_men_n602_));
  NA2        u0574(.A(men_men_n602_), .B(men_men_n600_), .Y(men_men_n603_));
  OR2        u0575(.A(men_men_n603_), .B(men_men_n570_), .Y(men_men_n604_));
  NOi31      u0576(.An(m), .B(n), .C(k), .Y(men_men_n605_));
  NA2        u0577(.A(men_men_n600_), .B(men_men_n605_), .Y(men_men_n606_));
  NO2        u0578(.A(men_men_n382_), .B(men_men_n293_), .Y(men_men_n607_));
  NAi21      u0579(.An(men_men_n606_), .B(men_men_n607_), .Y(men_men_n608_));
  NO2        u0580(.A(men_men_n302_), .B(men_men_n575_), .Y(men_men_n609_));
  NO2        u0581(.A(men_men_n523_), .B(men_men_n48_), .Y(men_men_n610_));
  NA2        u0582(.A(men_men_n610_), .B(men_men_n609_), .Y(men_men_n611_));
  NA4        u0583(.A(men_men_n611_), .B(men_men_n608_), .C(men_men_n604_), .D(men_men_n599_), .Y(men_men_n612_));
  NA2        u0584(.A(men_men_n103_), .B(men_men_n35_), .Y(men_men_n613_));
  NO2        u0585(.A(k), .B(men_men_n208_), .Y(men_men_n614_));
  NAi31      u0586(.An(men_men_n613_), .B(men_men_n350_), .C(men_men_n614_), .Y(men_men_n615_));
  NO2        u0587(.A(men_men_n521_), .B(men_men_n170_), .Y(men_men_n616_));
  NA2        u0588(.A(men_men_n494_), .B(men_men_n154_), .Y(men_men_n617_));
  NO3        u0589(.A(men_men_n380_), .B(men_men_n617_), .C(men_men_n82_), .Y(men_men_n618_));
  NO2        u0590(.A(men_men_n616_), .B(men_men_n618_), .Y(men_men_n619_));
  AN3        u0591(.A(f), .B(d), .C(b), .Y(men_men_n620_));
  OAI210     u0592(.A0(men_men_n620_), .A1(men_men_n124_), .B0(n), .Y(men_men_n621_));
  NA3        u0593(.A(men_men_n494_), .B(men_men_n154_), .C(men_men_n208_), .Y(men_men_n622_));
  AOI210     u0594(.A0(men_men_n621_), .A1(men_men_n223_), .B0(men_men_n622_), .Y(men_men_n623_));
  NAi31      u0595(.An(m), .B(n), .C(k), .Y(men_men_n624_));
  OAI210     u0596(.A0(men_men_n128_), .A1(men_men_n624_), .B0(men_men_n241_), .Y(men_men_n625_));
  OAI210     u0597(.A0(men_men_n625_), .A1(men_men_n623_), .B0(j), .Y(men_men_n626_));
  NA3        u0598(.A(men_men_n626_), .B(men_men_n619_), .C(men_men_n615_), .Y(men_men_n627_));
  NO4        u0599(.A(men_men_n627_), .B(men_men_n612_), .C(men_men_n597_), .D(men_men_n592_), .Y(men_men_n628_));
  NA2        u0600(.A(men_men_n368_), .B(men_men_n157_), .Y(men_men_n629_));
  NAi31      u0601(.An(u), .B(h), .C(f), .Y(men_men_n630_));
  OA210      u0602(.A0(men_men_n523_), .A1(n), .B0(men_men_n568_), .Y(men_men_n631_));
  NO2        u0603(.A(men_men_n631_), .B(men_men_n86_), .Y(men_men_n632_));
  INV        u0604(.A(men_men_n632_), .Y(men_men_n633_));
  AOI210     u0605(.A0(men_men_n633_), .A1(men_men_n629_), .B0(men_men_n516_), .Y(men_men_n634_));
  NO3        u0606(.A(u), .B(men_men_n207_), .C(men_men_n55_), .Y(men_men_n635_));
  NAi21      u0607(.An(h), .B(j), .Y(men_men_n636_));
  NA2        u0608(.A(men_men_n379_), .B(men_men_n635_), .Y(men_men_n637_));
  OR2        u0609(.A(men_men_n603_), .B(men_men_n72_), .Y(men_men_n638_));
  NA3        u0610(.A(men_men_n513_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n639_));
  NA2        u0611(.A(h), .B(men_men_n36_), .Y(men_men_n640_));
  NA2        u0612(.A(men_men_n95_), .B(men_men_n45_), .Y(men_men_n641_));
  NO2        u0613(.A(men_men_n641_), .B(men_men_n324_), .Y(men_men_n642_));
  OAI220     u0614(.A0(men_men_n571_), .A1(men_men_n564_), .B0(men_men_n318_), .B1(men_men_n514_), .Y(men_men_n643_));
  AOI210     u0615(.A0(men_men_n643_), .A1(m), .B0(men_men_n642_), .Y(men_men_n644_));
  NA4        u0616(.A(men_men_n644_), .B(men_men_n639_), .C(men_men_n638_), .D(men_men_n637_), .Y(men_men_n645_));
  NA2        u0617(.A(men_men_n321_), .B(men_men_n133_), .Y(men_men_n646_));
  OR2        u0618(.A(men_men_n1352_), .B(men_men_n538_), .Y(men_men_n647_));
  NA2        u0619(.A(men_men_n646_), .B(men_men_n647_), .Y(men_men_n648_));
  NA2        u0620(.A(men_men_n244_), .B(j), .Y(men_men_n649_));
  NA3        u0621(.A(men_men_n649_), .B(men_men_n501_), .C(men_men_n387_), .Y(men_men_n650_));
  NO4        u0622(.A(men_men_n650_), .B(men_men_n648_), .C(men_men_n645_), .D(men_men_n634_), .Y(men_men_n651_));
  NA4        u0623(.A(men_men_n651_), .B(men_men_n628_), .C(men_men_n585_), .D(men_men_n562_), .Y(men08));
  NO2        u0624(.A(k), .B(h), .Y(men_men_n653_));
  AO210      u0625(.A0(men_men_n242_), .A1(men_men_n438_), .B0(men_men_n653_), .Y(men_men_n654_));
  NO2        u0626(.A(men_men_n654_), .B(men_men_n291_), .Y(men_men_n655_));
  INV        u0627(.A(men_men_n594_), .Y(men_men_n656_));
  AOI210     u0628(.A0(f), .A1(men_men_n655_), .B0(men_men_n479_), .Y(men_men_n657_));
  NO2        u0629(.A(n), .B(men_men_n56_), .Y(men_men_n658_));
  NO4        u0630(.A(men_men_n365_), .B(men_men_n107_), .C(j), .D(men_men_n208_), .Y(men_men_n659_));
  AOI220     u0631(.A0(e), .A1(men_men_n338_), .B0(men_men_n659_), .B1(men_men_n658_), .Y(men_men_n660_));
  AOI210     u0632(.A0(men_men_n559_), .A1(men_men_n150_), .B0(men_men_n81_), .Y(men_men_n661_));
  NA3        u0633(.A(men_men_n210_), .B(men_men_n44_), .C(h), .Y(men_men_n662_));
  AN2        u0634(.A(l), .B(k), .Y(men_men_n663_));
  NA4        u0635(.A(men_men_n663_), .B(men_men_n103_), .C(men_men_n74_), .D(men_men_n208_), .Y(men_men_n664_));
  OAI210     u0636(.A0(men_men_n662_), .A1(u), .B0(men_men_n664_), .Y(men_men_n665_));
  NA2        u0637(.A(men_men_n665_), .B(men_men_n661_), .Y(men_men_n666_));
  NA4        u0638(.A(men_men_n666_), .B(men_men_n660_), .C(men_men_n657_), .D(men_men_n339_), .Y(men_men_n667_));
  AN2        u0639(.A(men_men_n524_), .B(men_men_n91_), .Y(men_men_n668_));
  NO3        u0640(.A(men_men_n167_), .B(men_men_n378_), .C(men_men_n107_), .Y(men_men_n669_));
  NO2        u0641(.A(men_men_n527_), .B(men_men_n34_), .Y(men_men_n670_));
  INV        u0642(.A(men_men_n128_), .Y(men_men_n671_));
  NO2        u0643(.A(men_men_n473_), .B(men_men_n126_), .Y(men_men_n672_));
  AOI210     u0644(.A0(men_men_n672_), .A1(men_men_n671_), .B0(men_men_n670_), .Y(men_men_n673_));
  NO3        u0645(.A(men_men_n308_), .B(men_men_n125_), .C(men_men_n40_), .Y(men_men_n674_));
  NAi21      u0646(.An(men_men_n674_), .B(men_men_n664_), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n675_), .B(men_men_n77_), .Y(men_men_n676_));
  OAI210     u0648(.A0(men_men_n673_), .A1(men_men_n82_), .B0(men_men_n676_), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n350_), .B(men_men_n42_), .Y(men_men_n678_));
  NA2        u0650(.A(men_men_n663_), .B(men_men_n215_), .Y(men_men_n679_));
  NO2        u0651(.A(men_men_n679_), .B(men_men_n320_), .Y(men_men_n680_));
  AOI210     u0652(.A0(men_men_n680_), .A1(i), .B0(men_men_n478_), .Y(men_men_n681_));
  NA3        u0653(.A(m), .B(l), .C(k), .Y(men_men_n682_));
  NO2        u0654(.A(men_men_n526_), .B(men_men_n262_), .Y(men_men_n683_));
  NOi21      u0655(.An(men_men_n683_), .B(men_men_n520_), .Y(men_men_n684_));
  NA4        u0656(.A(men_men_n108_), .B(l), .C(k), .D(men_men_n82_), .Y(men_men_n685_));
  INV        u0657(.A(men_men_n684_), .Y(men_men_n686_));
  NA3        u0658(.A(men_men_n686_), .B(men_men_n681_), .C(men_men_n678_), .Y(men_men_n687_));
  NO4        u0659(.A(men_men_n687_), .B(men_men_n677_), .C(men_men_n669_), .D(men_men_n667_), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n610_), .B(u), .Y(men_men_n689_));
  OR2        u0661(.A(men_men_n689_), .B(men_men_n529_), .Y(men_men_n690_));
  NO3        u0662(.A(men_men_n382_), .B(men_men_n514_), .C(h), .Y(men_men_n691_));
  AOI210     u0663(.A0(men_men_n691_), .A1(men_men_n108_), .B0(men_men_n487_), .Y(men_men_n692_));
  NA3        u0664(.A(men_men_n692_), .B(men_men_n690_), .C(men_men_n241_), .Y(men_men_n693_));
  NA2        u0665(.A(men_men_n663_), .B(men_men_n74_), .Y(men_men_n694_));
  NO3        u0666(.A(men_men_n167_), .B(n), .C(i), .Y(men_men_n695_));
  NOi21      u0667(.An(h), .B(j), .Y(men_men_n696_));
  NA2        u0668(.A(men_men_n696_), .B(f), .Y(men_men_n697_));
  INV        u0669(.A(men_men_n695_), .Y(men_men_n698_));
  NO2        u0670(.A(men_men_n698_), .B(men_men_n694_), .Y(men_men_n699_));
  AOI210     u0671(.A0(men_men_n693_), .A1(l), .B0(men_men_n699_), .Y(men_men_n700_));
  NO2        u0672(.A(j), .B(i), .Y(men_men_n701_));
  NA3        u0673(.A(men_men_n701_), .B(men_men_n79_), .C(l), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n701_), .B(men_men_n32_), .Y(men_men_n703_));
  OR2        u0675(.A(men_men_n702_), .B(men_men_n570_), .Y(men_men_n704_));
  NO3        u0676(.A(men_men_n145_), .B(men_men_n48_), .C(men_men_n105_), .Y(men_men_n705_));
  NO3        u0677(.A(men_men_n473_), .B(men_men_n425_), .C(j), .Y(men_men_n706_));
  NO2        u0678(.A(men_men_n689_), .B(men_men_n61_), .Y(men_men_n707_));
  NA2        u0679(.A(k), .B(j), .Y(men_men_n708_));
  NO2        u0680(.A(men_men_n291_), .B(men_men_n39_), .Y(men_men_n709_));
  NA2        u0681(.A(f), .B(men_men_n542_), .Y(men_men_n710_));
  AN3        u0682(.A(men_men_n710_), .B(men_men_n709_), .C(men_men_n94_), .Y(men_men_n711_));
  NAi21      u0683(.An(men_men_n581_), .B(men_men_n88_), .Y(men_men_n712_));
  INV        u0684(.A(men_men_n712_), .Y(men_men_n713_));
  NO2        u0685(.A(men_men_n291_), .B(men_men_n129_), .Y(men_men_n714_));
  AOI220     u0686(.A0(men_men_n714_), .A1(men_men_n595_), .B0(men_men_n674_), .B1(men_men_n661_), .Y(men_men_n715_));
  NO2        u0687(.A(men_men_n682_), .B(men_men_n86_), .Y(men_men_n716_));
  NA2        u0688(.A(men_men_n716_), .B(men_men_n569_), .Y(men_men_n717_));
  NO2        u0689(.A(men_men_n571_), .B(men_men_n111_), .Y(men_men_n718_));
  OAI210     u0690(.A0(men_men_n718_), .A1(men_men_n706_), .B0(m), .Y(men_men_n719_));
  NA3        u0691(.A(men_men_n719_), .B(men_men_n717_), .C(men_men_n715_), .Y(men_men_n720_));
  OR4        u0692(.A(men_men_n720_), .B(men_men_n713_), .C(men_men_n711_), .D(men_men_n707_), .Y(men_men_n721_));
  NA3        u0693(.A(men_men_n210_), .B(men_men_n438_), .C(men_men_n33_), .Y(men_men_n722_));
  NO4        u0694(.A(men_men_n473_), .B(men_men_n421_), .C(j), .D(f), .Y(men_men_n723_));
  OAI220     u0695(.A0(men_men_n662_), .A1(men_men_n656_), .B0(men_men_n324_), .B1(men_men_n37_), .Y(men_men_n724_));
  AOI210     u0696(.A0(men_men_n723_), .A1(men_men_n248_), .B0(men_men_n724_), .Y(men_men_n725_));
  NA3        u0697(.A(men_men_n533_), .B(men_men_n284_), .C(h), .Y(men_men_n726_));
  NO2        u0698(.A(men_men_n87_), .B(men_men_n46_), .Y(men_men_n727_));
  NO2        u0699(.A(men_men_n702_), .B(men_men_n72_), .Y(men_men_n728_));
  AOI210     u0700(.A0(men_men_n727_), .A1(men_men_n350_), .B0(men_men_n728_), .Y(men_men_n729_));
  NA3        u0701(.A(men_men_n729_), .B(men_men_n725_), .C(men_men_n722_), .Y(men_men_n730_));
  OR2        u0702(.A(men_men_n716_), .B(men_men_n91_), .Y(men_men_n731_));
  NA2        u0703(.A(men_men_n731_), .B(men_men_n229_), .Y(men_men_n732_));
  NO2        u0704(.A(men_men_n631_), .B(men_men_n74_), .Y(men_men_n733_));
  AOI210     u0705(.A0(men_men_n723_), .A1(men_men_n733_), .B0(men_men_n328_), .Y(men_men_n734_));
  OAI210     u0706(.A0(men_men_n682_), .A1(men_men_n630_), .B0(men_men_n507_), .Y(men_men_n735_));
  INV        u0707(.A(men_men_n735_), .Y(men_men_n736_));
  NA3        u0708(.A(men_men_n736_), .B(men_men_n734_), .C(men_men_n732_), .Y(men_men_n737_));
  NOi41      u0709(.An(men_men_n704_), .B(men_men_n737_), .C(men_men_n730_), .D(men_men_n721_), .Y(men_men_n738_));
  NO3        u0710(.A(men_men_n333_), .B(men_men_n293_), .C(men_men_n107_), .Y(men_men_n739_));
  INV        u0711(.A(men_men_n739_), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n45_), .B(men_men_n55_), .Y(men_men_n741_));
  NO3        u0713(.A(men_men_n741_), .B(men_men_n703_), .C(men_men_n268_), .Y(men_men_n742_));
  NO3        u0714(.A(men_men_n514_), .B(men_men_n89_), .C(h), .Y(men_men_n743_));
  AOI210     u0715(.A0(men_men_n743_), .A1(men_men_n658_), .B0(men_men_n742_), .Y(men_men_n744_));
  NA3        u0716(.A(men_men_n744_), .B(men_men_n740_), .C(men_men_n390_), .Y(men_men_n745_));
  OR2        u0717(.A(men_men_n630_), .B(men_men_n87_), .Y(men_men_n746_));
  NOi31      u0718(.An(b), .B(d), .C(a), .Y(men_men_n747_));
  OAI220     u0719(.A0(n), .A1(men_men_n746_), .B0(men_men_n726_), .B1(n), .Y(men_men_n748_));
  NO2        u0720(.A(men_men_n320_), .B(men_men_n111_), .Y(men_men_n749_));
  NOi21      u0721(.An(men_men_n749_), .B(men_men_n155_), .Y(men_men_n750_));
  INV        u0722(.A(men_men_n750_), .Y(men_men_n751_));
  OAI210     u0723(.A0(men_men_n662_), .A1(men_men_n380_), .B0(men_men_n751_), .Y(men_men_n752_));
  NA2        u0724(.A(men_men_n714_), .B(men_men_n635_), .Y(men_men_n753_));
  NO2        u0725(.A(men_men_n315_), .B(men_men_n228_), .Y(men_men_n754_));
  OAI210     u0726(.A0(men_men_n91_), .A1(men_men_n88_), .B0(men_men_n754_), .Y(men_men_n755_));
  NA2        u0727(.A(men_men_n115_), .B(men_men_n81_), .Y(men_men_n756_));
  AOI210     u0728(.A0(men_men_n411_), .A1(men_men_n403_), .B0(men_men_n756_), .Y(men_men_n757_));
  INV        u0729(.A(men_men_n755_), .Y(men_men_n758_));
  NAi21      u0730(.An(men_men_n685_), .B(men_men_n422_), .Y(men_men_n759_));
  NO2        u0731(.A(men_men_n262_), .B(i), .Y(men_men_n760_));
  NA2        u0732(.A(men_men_n573_), .B(men_men_n351_), .Y(men_men_n761_));
  AN2        u0733(.A(men_men_n761_), .B(men_men_n759_), .Y(men_men_n762_));
  NAi31      u0734(.An(men_men_n758_), .B(men_men_n762_), .C(men_men_n753_), .Y(men_men_n763_));
  NO4        u0735(.A(men_men_n763_), .B(men_men_n752_), .C(men_men_n748_), .D(men_men_n745_), .Y(men_men_n764_));
  NA4        u0736(.A(men_men_n764_), .B(men_men_n738_), .C(men_men_n700_), .D(men_men_n688_), .Y(men09));
  NA2        u0737(.A(f), .B(e), .Y(men_men_n766_));
  NO2        u0738(.A(men_men_n220_), .B(men_men_n107_), .Y(men_men_n767_));
  NA2        u0739(.A(men_men_n767_), .B(u), .Y(men_men_n768_));
  NA4        u0740(.A(men_men_n302_), .B(men_men_n460_), .C(men_men_n251_), .D(men_men_n113_), .Y(men_men_n769_));
  AOI210     u0741(.A0(men_men_n769_), .A1(u), .B0(men_men_n457_), .Y(men_men_n770_));
  AOI210     u0742(.A0(men_men_n770_), .A1(men_men_n768_), .B0(men_men_n766_), .Y(men_men_n771_));
  NA2        u0743(.A(men_men_n431_), .B(e), .Y(men_men_n772_));
  NO2        u0744(.A(men_men_n772_), .B(men_men_n498_), .Y(men_men_n773_));
  INV        u0745(.A(men_men_n773_), .Y(men_men_n774_));
  NO2        u0746(.A(men_men_n197_), .B(men_men_n207_), .Y(men_men_n775_));
  NA3        u0747(.A(m), .B(l), .C(i), .Y(men_men_n776_));
  OAI220     u0748(.A0(men_men_n571_), .A1(men_men_n776_), .B0(men_men_n342_), .B1(men_men_n515_), .Y(men_men_n777_));
  NA4        u0749(.A(men_men_n83_), .B(men_men_n82_), .C(u), .D(f), .Y(men_men_n778_));
  NA3        u0750(.A(men_men_n746_), .B(men_men_n552_), .C(men_men_n507_), .Y(men_men_n779_));
  OR2        u0751(.A(men_men_n779_), .B(men_men_n775_), .Y(men_men_n780_));
  INV        u0752(.A(men_men_n331_), .Y(men_men_n781_));
  NO2        u0753(.A(men_men_n121_), .B(men_men_n120_), .Y(men_men_n782_));
  NO2        u0754(.A(m), .B(men_men_n575_), .Y(men_men_n783_));
  NA2        u0755(.A(men_men_n334_), .B(men_men_n335_), .Y(men_men_n784_));
  NA2        u0756(.A(men_men_n783_), .B(men_men_n781_), .Y(men_men_n785_));
  NA2        u0757(.A(men_men_n785_), .B(men_men_n596_), .Y(men_men_n786_));
  NO2        u0758(.A(men_men_n567_), .B(men_men_n484_), .Y(men_men_n787_));
  NA2        u0759(.A(f), .B(m), .Y(men_men_n788_));
  NO2        u0760(.A(men_men_n788_), .B(men_men_n51_), .Y(men_men_n789_));
  NOi32      u0761(.An(u), .Bn(f), .C(d), .Y(men_men_n790_));
  NA4        u0762(.A(men_men_n790_), .B(men_men_n579_), .C(men_men_n29_), .D(m), .Y(men_men_n791_));
  NOi21      u0763(.An(men_men_n303_), .B(men_men_n791_), .Y(men_men_n792_));
  AOI210     u0764(.A0(men_men_n789_), .A1(men_men_n532_), .B0(men_men_n792_), .Y(men_men_n793_));
  AN2        u0765(.A(f), .B(d), .Y(men_men_n794_));
  BUFFER     u0766(.A(men_men_n476_), .Y(men_men_n795_));
  NO2        u0767(.A(men_men_n624_), .B(men_men_n320_), .Y(men_men_n796_));
  NO2        u0768(.A(men_men_n796_), .B(men_men_n225_), .Y(men_men_n797_));
  OAI220     u0769(.A0(men_men_n784_), .A1(n), .B0(n), .B1(men_men_n426_), .Y(men_men_n798_));
  NA3        u0770(.A(men_men_n154_), .B(men_men_n103_), .C(men_men_n102_), .Y(men_men_n799_));
  NO2        u0771(.A(men_men_n331_), .B(men_men_n799_), .Y(men_men_n800_));
  NOi41      u0772(.An(men_men_n218_), .B(men_men_n800_), .C(men_men_n798_), .D(men_men_n297_), .Y(men_men_n801_));
  NA3        u0773(.A(e), .B(men_men_n496_), .C(f), .Y(men_men_n802_));
  OR2        u0774(.A(men_men_n630_), .B(men_men_n530_), .Y(men_men_n803_));
  NA4        u0775(.A(men_men_n803_), .B(men_men_n802_), .C(men_men_n801_), .D(men_men_n797_), .Y(men_men_n804_));
  NO4        u0776(.A(men_men_n804_), .B(men_men_n795_), .C(men_men_n786_), .D(men_men_n780_), .Y(men_men_n805_));
  NO2        u0777(.A(n), .B(men_men_n778_), .Y(men_men_n806_));
  NO2        u0778(.A(men_men_n416_), .B(men_men_n766_), .Y(men_men_n807_));
  NA2        u0779(.A(e), .B(d), .Y(men_men_n808_));
  OAI220     u0780(.A0(men_men_n808_), .A1(c), .B0(men_men_n315_), .B1(d), .Y(men_men_n809_));
  NA3        u0781(.A(men_men_n809_), .B(men_men_n442_), .C(men_men_n494_), .Y(men_men_n810_));
  AOI210     u0782(.A0(men_men_n502_), .A1(men_men_n174_), .B0(men_men_n222_), .Y(men_men_n811_));
  AOI210     u0783(.A0(men_men_n595_), .A1(men_men_n337_), .B0(men_men_n811_), .Y(men_men_n812_));
  NA2        u0784(.A(men_men_n812_), .B(men_men_n810_), .Y(men_men_n813_));
  NO2        u0785(.A(men_men_n813_), .B(men_men_n806_), .Y(men_men_n814_));
  AO210      u0786(.A0(men_men_n331_), .A1(men_men_n656_), .B0(men_men_n211_), .Y(men_men_n815_));
  AOI220     u0787(.A0(h), .A1(men_men_n796_), .B0(men_men_n586_), .B1(men_men_n594_), .Y(men_men_n816_));
  OAI210     u0788(.A0(men_men_n772_), .A1(men_men_n164_), .B0(men_men_n816_), .Y(men_men_n817_));
  AOI210     u0789(.A0(men_men_n112_), .A1(men_men_n111_), .B0(men_men_n250_), .Y(men_men_n818_));
  NOi31      u0790(.An(men_men_n532_), .B(men_men_n788_), .C(men_men_n285_), .Y(men_men_n819_));
  NO2        u0791(.A(men_men_n777_), .B(men_men_n817_), .Y(men_men_n820_));
  AO210      u0792(.A0(men_men_n442_), .A1(men_men_n696_), .B0(men_men_n169_), .Y(men_men_n821_));
  OAI210     u0793(.A0(men_men_n821_), .A1(men_men_n444_), .B0(men_men_n809_), .Y(men_men_n822_));
  AN3        u0794(.A(men_men_n822_), .B(men_men_n820_), .C(men_men_n815_), .Y(men_men_n823_));
  NA4        u0795(.A(men_men_n823_), .B(men_men_n814_), .C(men_men_n805_), .D(men_men_n774_), .Y(men12));
  NO2        u0796(.A(men_men_n441_), .B(c), .Y(men_men_n825_));
  NO4        u0797(.A(men_men_n430_), .B(men_men_n242_), .C(men_men_n563_), .D(men_men_n208_), .Y(men_men_n826_));
  NA2        u0798(.A(men_men_n826_), .B(men_men_n825_), .Y(men_men_n827_));
  NO2        u0799(.A(men_men_n441_), .B(men_men_n110_), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n782_), .B(men_men_n342_), .Y(men_men_n829_));
  NO2        u0801(.A(men_men_n630_), .B(men_men_n365_), .Y(men_men_n830_));
  AOI210     u0802(.A0(men_men_n829_), .A1(men_men_n828_), .B0(men_men_n830_), .Y(men_men_n831_));
  NA3        u0803(.A(men_men_n831_), .B(men_men_n827_), .C(men_men_n429_), .Y(men_men_n832_));
  AOI210     u0804(.A0(men_men_n224_), .A1(men_men_n330_), .B0(men_men_n194_), .Y(men_men_n833_));
  OR2        u0805(.A(men_men_n833_), .B(men_men_n826_), .Y(men_men_n834_));
  AOI210     u0806(.A0(men_men_n327_), .A1(men_men_n376_), .B0(men_men_n208_), .Y(men_men_n835_));
  OAI210     u0807(.A0(men_men_n835_), .A1(men_men_n834_), .B0(men_men_n389_), .Y(men_men_n836_));
  NO2        u0808(.A(men_men_n613_), .B(men_men_n253_), .Y(men_men_n837_));
  NO2        u0809(.A(men_men_n571_), .B(men_men_n776_), .Y(men_men_n838_));
  NA2        u0810(.A(men_men_n754_), .B(men_men_n837_), .Y(men_men_n839_));
  NO2        u0811(.A(men_men_n145_), .B(men_men_n228_), .Y(men_men_n840_));
  NA3        u0812(.A(men_men_n840_), .B(men_men_n231_), .C(i), .Y(men_men_n841_));
  NA3        u0813(.A(men_men_n841_), .B(men_men_n839_), .C(men_men_n836_), .Y(men_men_n842_));
  OR2        u0814(.A(men_men_n316_), .B(men_men_n828_), .Y(men_men_n843_));
  NA2        u0815(.A(men_men_n843_), .B(men_men_n343_), .Y(men_men_n844_));
  NO3        u0816(.A(men_men_n126_), .B(men_men_n146_), .C(men_men_n208_), .Y(men_men_n845_));
  NA2        u0817(.A(men_men_n845_), .B(men_men_n519_), .Y(men_men_n846_));
  NA2        u0818(.A(men_men_n431_), .B(u), .Y(men_men_n847_));
  NA3        u0819(.A(men_men_n847_), .B(men_men_n846_), .C(men_men_n844_), .Y(men_men_n848_));
  NO3        u0820(.A(men_men_n633_), .B(men_men_n87_), .C(men_men_n44_), .Y(men_men_n849_));
  NO4        u0821(.A(men_men_n849_), .B(men_men_n848_), .C(men_men_n842_), .D(men_men_n832_), .Y(men_men_n850_));
  NO2        u0822(.A(men_men_n356_), .B(men_men_n355_), .Y(men_men_n851_));
  NA2        u0823(.A(men_men_n568_), .B(men_men_n72_), .Y(men_men_n852_));
  NOi21      u0824(.An(men_men_n33_), .B(men_men_n624_), .Y(men_men_n853_));
  AOI220     u0825(.A0(men_men_n853_), .A1(c), .B0(men_men_n852_), .B1(men_men_n851_), .Y(men_men_n854_));
  OAI210     u0826(.A0(men_men_n241_), .A1(men_men_n44_), .B0(men_men_n854_), .Y(men_men_n855_));
  NA2        u0827(.A(men_men_n422_), .B(men_men_n255_), .Y(men_men_n856_));
  NO3        u0828(.A(men_men_n756_), .B(men_men_n84_), .C(men_men_n394_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n856_), .B(men_men_n312_), .Y(men_men_n858_));
  NO2        u0830(.A(men_men_n48_), .B(men_men_n44_), .Y(men_men_n859_));
  NO2        u0831(.A(men_men_n490_), .B(men_men_n293_), .Y(men_men_n860_));
  NO2        u0832(.A(men_men_n860_), .B(men_men_n353_), .Y(men_men_n861_));
  NO2        u0833(.A(men_men_n861_), .B(men_men_n138_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n605_), .B(men_men_n351_), .Y(men_men_n863_));
  NO4        u0835(.A(men_men_n352_), .B(men_men_n862_), .C(men_men_n858_), .D(men_men_n855_), .Y(men_men_n864_));
  NA2        u0836(.A(men_men_n337_), .B(u), .Y(men_men_n865_));
  NA2        u0837(.A(men_men_n157_), .B(i), .Y(men_men_n866_));
  NA2        u0838(.A(men_men_n45_), .B(i), .Y(men_men_n867_));
  OAI220     u0839(.A0(men_men_n867_), .A1(men_men_n193_), .B0(men_men_n866_), .B1(men_men_n87_), .Y(men_men_n868_));
  AOI210     u0840(.A0(men_men_n405_), .A1(men_men_n36_), .B0(men_men_n868_), .Y(men_men_n869_));
  NA2        u0841(.A(men_men_n541_), .B(men_men_n369_), .Y(men_men_n870_));
  NO2        u0842(.A(n), .B(men_men_n1354_), .Y(men_men_n871_));
  OAI220     u0843(.A0(men_men_n871_), .A1(men_men_n865_), .B0(men_men_n869_), .B1(men_men_n324_), .Y(men_men_n872_));
  NO2        u0844(.A(men_men_n630_), .B(men_men_n484_), .Y(men_men_n873_));
  NA3        u0845(.A(men_men_n334_), .B(men_men_n600_), .C(i), .Y(men_men_n874_));
  NA2        u0846(.A(men_men_n873_), .B(m), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n580_), .B(men_men_n108_), .Y(men_men_n876_));
  OR3        u0848(.A(men_men_n302_), .B(men_men_n421_), .C(f), .Y(men_men_n877_));
  NA3        u0849(.A(men_men_n600_), .B(men_men_n79_), .C(i), .Y(men_men_n878_));
  OA220      u0850(.A0(men_men_n878_), .A1(men_men_n876_), .B0(men_men_n877_), .B1(men_men_n570_), .Y(men_men_n879_));
  NA3        u0851(.A(men_men_n317_), .B(men_men_n112_), .C(u), .Y(men_men_n880_));
  AOI210     u0852(.A0(men_men_n640_), .A1(men_men_n880_), .B0(m), .Y(men_men_n881_));
  OAI210     u0853(.A0(men_men_n881_), .A1(men_men_n829_), .B0(men_men_n316_), .Y(men_men_n882_));
  NA2        u0854(.A(men_men_n778_), .B(men_men_n426_), .Y(men_men_n883_));
  NA2        u0855(.A(men_men_n216_), .B(h), .Y(men_men_n884_));
  NA3        u0856(.A(men_men_n884_), .B(men_men_n878_), .C(men_men_n877_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n885_), .B(men_men_n248_), .Y(men_men_n886_));
  NA4        u0858(.A(men_men_n886_), .B(men_men_n882_), .C(men_men_n879_), .D(men_men_n875_), .Y(men_men_n887_));
  NO2        u0859(.A(men_men_n365_), .B(men_men_n86_), .Y(men_men_n888_));
  OAI210     u0860(.A0(men_men_n888_), .A1(men_men_n837_), .B0(men_men_n229_), .Y(men_men_n889_));
  NA2        u0861(.A(men_men_n632_), .B(men_men_n83_), .Y(men_men_n890_));
  NO2        u0862(.A(men_men_n446_), .B(men_men_n208_), .Y(men_men_n891_));
  AOI220     u0863(.A0(men_men_n891_), .A1(men_men_n370_), .B0(men_men_n843_), .B1(men_men_n212_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n569_), .B(men_men_n85_), .Y(men_men_n893_));
  NA4        u0865(.A(men_men_n893_), .B(men_men_n892_), .C(men_men_n890_), .D(men_men_n889_), .Y(men_men_n894_));
  NO2        u0866(.A(men_men_n883_), .B(men_men_n838_), .Y(men_men_n895_));
  AOI210     u0867(.A0(men_men_n406_), .A1(men_men_n398_), .B0(men_men_n756_), .Y(men_men_n896_));
  OAI210     u0868(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n104_), .Y(men_men_n897_));
  AOI210     u0869(.A0(men_men_n897_), .A1(men_men_n524_), .B0(men_men_n896_), .Y(men_men_n898_));
  NA2        u0870(.A(men_men_n881_), .B(men_men_n828_), .Y(men_men_n899_));
  NO3        u0871(.A(l), .B(men_men_n48_), .C(men_men_n44_), .Y(men_men_n900_));
  AOI220     u0872(.A0(men_men_n900_), .A1(men_men_n598_), .B0(men_men_n616_), .B1(men_men_n519_), .Y(men_men_n901_));
  NA4        u0873(.A(men_men_n901_), .B(men_men_n899_), .C(men_men_n898_), .D(men_men_n895_), .Y(men_men_n902_));
  NO4        u0874(.A(men_men_n902_), .B(men_men_n894_), .C(men_men_n887_), .D(men_men_n872_), .Y(men_men_n903_));
  NAi31      u0875(.An(men_men_n134_), .B(men_men_n407_), .C(n), .Y(men_men_n904_));
  NO2        u0876(.A(m), .B(men_men_n904_), .Y(men_men_n905_));
  NO2        u0877(.A(men_men_n262_), .B(men_men_n134_), .Y(men_men_n906_));
  AOI210     u0878(.A0(men_men_n906_), .A1(men_men_n485_), .B0(men_men_n905_), .Y(men_men_n907_));
  NA2        u0879(.A(men_men_n479_), .B(i), .Y(men_men_n908_));
  NA2        u0880(.A(men_men_n908_), .B(men_men_n907_), .Y(men_men_n909_));
  NA2        u0881(.A(men_men_n222_), .B(men_men_n165_), .Y(men_men_n910_));
  NO3        u0882(.A(men_men_n299_), .B(men_men_n431_), .C(men_men_n169_), .Y(men_men_n911_));
  NOi31      u0883(.An(men_men_n910_), .B(men_men_n911_), .C(men_men_n208_), .Y(men_men_n912_));
  NAi21      u0884(.An(men_men_n541_), .B(men_men_n891_), .Y(men_men_n913_));
  NO3        u0885(.A(men_men_n425_), .B(men_men_n302_), .C(men_men_n74_), .Y(men_men_n914_));
  INV        u0886(.A(men_men_n914_), .Y(men_men_n915_));
  NA2        u0887(.A(men_men_n915_), .B(men_men_n913_), .Y(men_men_n916_));
  NO2        u0888(.A(men_men_n874_), .B(n), .Y(men_men_n917_));
  NA2        u0889(.A(men_men_n833_), .B(men_men_n825_), .Y(men_men_n918_));
  NA2        u0890(.A(men_men_n513_), .B(men_men_n366_), .Y(men_men_n919_));
  NA2        u0891(.A(men_men_n918_), .B(men_men_n593_), .Y(men_men_n920_));
  OAI210     u0892(.A0(men_men_n833_), .A1(men_men_n826_), .B0(men_men_n910_), .Y(men_men_n921_));
  NA3        u0893(.A(men_men_n870_), .B(men_men_n474_), .C(men_men_n45_), .Y(men_men_n922_));
  NA2        u0894(.A(men_men_n368_), .B(men_men_n366_), .Y(men_men_n923_));
  NA4        u0895(.A(men_men_n923_), .B(men_men_n922_), .C(men_men_n921_), .D(men_men_n263_), .Y(men_men_n924_));
  OR3        u0896(.A(men_men_n924_), .B(men_men_n920_), .C(men_men_n917_), .Y(men_men_n925_));
  NO4        u0897(.A(men_men_n925_), .B(men_men_n916_), .C(men_men_n912_), .D(men_men_n909_), .Y(men_men_n926_));
  NA4        u0898(.A(men_men_n926_), .B(men_men_n903_), .C(men_men_n864_), .D(men_men_n850_), .Y(men13));
  NA2        u0899(.A(men_men_n45_), .B(men_men_n82_), .Y(men_men_n928_));
  AN2        u0900(.A(c), .B(b), .Y(men_men_n929_));
  NO4        u0901(.A(e), .B(men_men_n1358_), .C(men_men_n928_), .D(men_men_n564_), .Y(men_men_n930_));
  NA2        u0902(.A(men_men_n255_), .B(men_men_n929_), .Y(men_men_n931_));
  NO4        u0903(.A(men_men_n931_), .B(e), .C(men_men_n866_), .D(a), .Y(men_men_n932_));
  NA2        u0904(.A(men_men_n133_), .B(men_men_n44_), .Y(men_men_n933_));
  NO4        u0905(.A(men_men_n933_), .B(d), .C(men_men_n571_), .D(men_men_n298_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n636_), .B(men_men_n219_), .Y(men_men_n935_));
  AN2        u0907(.A(d), .B(c), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n936_), .B(men_men_n110_), .Y(men_men_n937_));
  NO3        u0909(.A(men_men_n937_), .B(men_men_n170_), .C(men_men_n162_), .Y(men_men_n938_));
  NO3        u0910(.A(men_men_n933_), .B(men_men_n567_), .C(men_men_n298_), .Y(men_men_n939_));
  AO210      u0911(.A0(men_men_n938_), .A1(men_men_n935_), .B0(men_men_n939_), .Y(men_men_n940_));
  OR4        u0912(.A(men_men_n940_), .B(men_men_n934_), .C(men_men_n932_), .D(men_men_n930_), .Y(men_men_n941_));
  NAi32      u0913(.An(f), .Bn(e), .C(c), .Y(men_men_n942_));
  OR3        u0914(.A(men_men_n219_), .B(men_men_n170_), .C(men_men_n162_), .Y(men_men_n943_));
  NO2        u0915(.A(men_men_n943_), .B(men_men_n942_), .Y(men_men_n944_));
  INV        u0916(.A(men_men_n298_), .Y(men_men_n945_));
  NA2        u0917(.A(men_men_n602_), .B(men_men_n1351_), .Y(men_men_n946_));
  NOi21      u0918(.An(men_men_n945_), .B(men_men_n946_), .Y(men_men_n947_));
  NO2        u0919(.A(men_men_n708_), .B(men_men_n107_), .Y(men_men_n948_));
  NOi41      u0920(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n949_));
  NA2        u0921(.A(men_men_n949_), .B(men_men_n948_), .Y(men_men_n950_));
  NO2        u0922(.A(men_men_n950_), .B(men_men_n942_), .Y(men_men_n951_));
  NA3        u0923(.A(k), .B(j), .C(i), .Y(men_men_n952_));
  NO3        u0924(.A(men_men_n952_), .B(men_men_n298_), .C(men_men_n86_), .Y(men_men_n953_));
  OR4        u0925(.A(men_men_n953_), .B(men_men_n951_), .C(men_men_n947_), .D(men_men_n944_), .Y(men_men_n954_));
  NA3        u0926(.A(men_men_n454_), .B(men_men_n326_), .C(men_men_n55_), .Y(men_men_n955_));
  NO3        u0927(.A(men_men_n955_), .B(men_men_n567_), .C(men_men_n44_), .Y(men_men_n956_));
  NO2        u0928(.A(f), .B(c), .Y(men_men_n957_));
  NOi21      u0929(.An(men_men_n957_), .B(men_men_n430_), .Y(men_men_n958_));
  NA2        u0930(.A(men_men_n958_), .B(men_men_n58_), .Y(men_men_n959_));
  NO3        u0931(.A(k), .B(h), .C(l), .Y(men_men_n960_));
  NOi21      u0932(.An(men_men_n960_), .B(men_men_n959_), .Y(men_men_n961_));
  OR2        u0933(.A(men_men_n961_), .B(men_men_n956_), .Y(men_men_n962_));
  OR3        u0934(.A(men_men_n962_), .B(men_men_n954_), .C(men_men_n941_), .Y(men02));
  OR2        u0935(.A(l), .B(k), .Y(men_men_n964_));
  OR3        u0936(.A(h), .B(u), .C(f), .Y(men_men_n965_));
  OR3        u0937(.A(n), .B(m), .C(i), .Y(men_men_n966_));
  NO4        u0938(.A(men_men_n966_), .B(men_men_n965_), .C(men_men_n964_), .D(e), .Y(men_men_n967_));
  NO2        u0939(.A(men_men_n953_), .B(men_men_n934_), .Y(men_men_n968_));
  AN3        u0940(.A(u), .B(f), .C(c), .Y(men_men_n969_));
  NA3        u0941(.A(men_men_n969_), .B(men_men_n454_), .C(h), .Y(men_men_n970_));
  OR2        u0942(.A(men_men_n298_), .B(men_men_n970_), .Y(men_men_n971_));
  NO3        u0943(.A(men_men_n955_), .B(men_men_n933_), .C(men_men_n567_), .Y(men_men_n972_));
  NO2        u0944(.A(men_men_n972_), .B(men_men_n944_), .Y(men_men_n973_));
  NA2        u0945(.A(i), .B(h), .Y(men_men_n974_));
  NO2        u0946(.A(men_men_n974_), .B(men_men_n126_), .Y(men_men_n975_));
  NO3        u0947(.A(men_men_n135_), .B(men_men_n275_), .C(men_men_n208_), .Y(men_men_n976_));
  AOI210     u0948(.A0(men_men_n976_), .A1(men_men_n975_), .B0(men_men_n947_), .Y(men_men_n977_));
  NA3        u0949(.A(c), .B(b), .C(a), .Y(men_men_n978_));
  NO3        u0950(.A(men_men_n978_), .B(men_men_n808_), .C(men_men_n207_), .Y(men_men_n979_));
  NO3        u0951(.A(men_men_n952_), .B(men_men_n48_), .C(men_men_n107_), .Y(men_men_n980_));
  NA2        u0952(.A(men_men_n980_), .B(men_men_n979_), .Y(men_men_n981_));
  AN4        u0953(.A(men_men_n981_), .B(men_men_n977_), .C(men_men_n973_), .D(men_men_n971_), .Y(men_men_n982_));
  NA2        u0954(.A(men_men_n950_), .B(men_men_n943_), .Y(men_men_n983_));
  AOI210     u0955(.A0(men_men_n983_), .A1(men_men_n936_), .B0(men_men_n930_), .Y(men_men_n984_));
  NAi41      u0956(.An(men_men_n967_), .B(men_men_n984_), .C(men_men_n982_), .D(men_men_n968_), .Y(men03));
  NA4        u0957(.A(men_men_n83_), .B(men_men_n82_), .C(u), .D(men_men_n207_), .Y(men_men_n986_));
  NA4        u0958(.A(men_men_n558_), .B(m), .C(men_men_n107_), .D(men_men_n207_), .Y(men_men_n987_));
  NA3        u0959(.A(men_men_n987_), .B(men_men_n357_), .C(men_men_n986_), .Y(men_men_n988_));
  NOi31      u0960(.An(i), .B(k), .C(j), .Y(men_men_n989_));
  NA4        u0961(.A(men_men_n989_), .B(e), .C(men_men_n334_), .D(men_men_n326_), .Y(men_men_n990_));
  OAI210     u0962(.A0(men_men_n756_), .A1(men_men_n408_), .B0(men_men_n990_), .Y(men_men_n991_));
  NOi31      u0963(.An(m), .B(n), .C(f), .Y(men_men_n992_));
  NA2        u0964(.A(men_men_n992_), .B(men_men_n50_), .Y(men_men_n993_));
  AN2        u0965(.A(e), .B(c), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n994_), .B(a), .Y(men_men_n995_));
  NO2        u0967(.A(men_men_n995_), .B(men_men_n993_), .Y(men_men_n996_));
  NA2        u0968(.A(men_men_n494_), .B(l), .Y(men_men_n997_));
  INV        u0969(.A(men_men_n934_), .Y(men_men_n998_));
  NO2        u0970(.A(men_men_n82_), .B(u), .Y(men_men_n999_));
  AOI210     u0971(.A0(men_men_n999_), .A1(i), .B0(men_men_n960_), .Y(men_men_n1000_));
  OR2        u0972(.A(men_men_n1000_), .B(men_men_n959_), .Y(men_men_n1001_));
  NA3        u0973(.A(men_men_n1001_), .B(men_men_n998_), .C(men_men_n990_), .Y(men_men_n1002_));
  NO2        u0974(.A(men_men_n1002_), .B(men_men_n777_), .Y(men_men_n1003_));
  NA2        u0975(.A(c), .B(b), .Y(men_men_n1004_));
  OAI210     u0976(.A0(men_men_n788_), .A1(men_men_n770_), .B0(men_men_n401_), .Y(men_men_n1005_));
  OAI210     u0977(.A0(men_men_n1005_), .A1(men_men_n789_), .B0(c), .Y(men_men_n1006_));
  BUFFER     u0978(.A(men_men_n409_), .Y(men_men_n1007_));
  NA3        u0979(.A(men_men_n415_), .B(men_men_n545_), .C(f), .Y(men_men_n1008_));
  OAI210     u0980(.A0(men_men_n535_), .A1(men_men_n38_), .B0(e), .Y(men_men_n1009_));
  NA3        u0981(.A(men_men_n1009_), .B(men_men_n1008_), .C(men_men_n1007_), .Y(men_men_n1010_));
  NA2        u0982(.A(men_men_n251_), .B(men_men_n113_), .Y(men_men_n1011_));
  OAI210     u0983(.A0(men_men_n1011_), .A1(men_men_n279_), .B0(u), .Y(men_men_n1012_));
  AOI210     u0984(.A0(men_men_n1012_), .A1(men_men_n285_), .B0(men_men_n978_), .Y(men_men_n1013_));
  AOI210     u0985(.A0(men_men_n1013_), .A1(men_men_n108_), .B0(men_men_n1010_), .Y(men_men_n1014_));
  NO2        u0986(.A(men_men_n176_), .B(men_men_n228_), .Y(men_men_n1015_));
  NA3        u0987(.A(men_men_n818_), .B(men_men_n997_), .C(men_men_n460_), .Y(men_men_n1016_));
  NA2        u0988(.A(men_men_n153_), .B(men_men_n32_), .Y(men_men_n1017_));
  AOI210     u0989(.A0(men_men_n863_), .A1(men_men_n1017_), .B0(men_men_n208_), .Y(men_men_n1018_));
  OAI210     u0990(.A0(men_men_n1018_), .A1(men_men_n434_), .B0(b), .Y(men_men_n1019_));
  NO2        u0991(.A(men_men_n359_), .B(men_men_n358_), .Y(men_men_n1020_));
  NA4        u0992(.A(men_men_n1019_), .B(men_men_n1014_), .C(men_men_n1006_), .D(men_men_n1003_), .Y(men00));
  NO2        u0993(.A(men_men_n292_), .B(men_men_n267_), .Y(men_men_n1022_));
  NO2        u0994(.A(men_men_n1022_), .B(men_men_n559_), .Y(men_men_n1023_));
  AOI210     u0995(.A0(men_men_n807_), .A1(men_men_n840_), .B0(men_men_n991_), .Y(men_men_n1024_));
  NO2        u0996(.A(men_men_n857_), .B(men_men_n668_), .Y(men_men_n1025_));
  NA3        u0997(.A(men_men_n1025_), .B(men_men_n1024_), .C(men_men_n898_), .Y(men_men_n1026_));
  NA2        u0998(.A(men_men_n496_), .B(f), .Y(men_men_n1027_));
  OAI210     u0999(.A0(m), .A1(men_men_n39_), .B0(men_men_n617_), .Y(men_men_n1028_));
  NA3        u1000(.A(men_men_n1028_), .B(men_men_n247_), .C(n), .Y(men_men_n1029_));
  AOI210     u1001(.A0(men_men_n1029_), .A1(men_men_n1027_), .B0(men_men_n937_), .Y(men_men_n1030_));
  NO4        u1002(.A(men_men_n1030_), .B(men_men_n1026_), .C(men_men_n1023_), .D(men_men_n954_), .Y(men_men_n1031_));
  NA3        u1003(.A(d), .B(men_men_n55_), .C(b), .Y(men_men_n1032_));
  NOi31      u1004(.An(n), .B(m), .C(i), .Y(men_men_n1033_));
  NA3        u1005(.A(men_men_n1033_), .B(men_men_n620_), .C(men_men_n50_), .Y(men_men_n1034_));
  INV        u1006(.A(men_men_n1034_), .Y(men_men_n1035_));
  NO3        u1007(.A(men_men_n1035_), .B(men_men_n1020_), .C(men_men_n819_), .Y(men_men_n1036_));
  NO4        u1008(.A(men_men_n1353_), .B(men_men_n344_), .C(men_men_n1004_), .D(men_men_n58_), .Y(men_men_n1037_));
  NA3        u1009(.A(h), .B(men_men_n215_), .C(u), .Y(men_men_n1038_));
  OA220      u1010(.A0(men_men_n1038_), .A1(men_men_n1032_), .B0(men_men_n371_), .B1(men_men_n128_), .Y(men_men_n1039_));
  NO2        u1011(.A(h), .B(u), .Y(men_men_n1040_));
  NA4        u1012(.A(men_men_n485_), .B(men_men_n454_), .C(men_men_n1040_), .D(men_men_n929_), .Y(men_men_n1041_));
  OAI220     u1013(.A0(men_men_n515_), .A1(men_men_n575_), .B0(men_men_n87_), .B1(men_men_n86_), .Y(men_men_n1042_));
  NA2        u1014(.A(men_men_n1042_), .B(men_men_n524_), .Y(men_men_n1043_));
  NA3        u1015(.A(men_men_n1043_), .B(men_men_n1041_), .C(men_men_n1039_), .Y(men_men_n1044_));
  NO3        u1016(.A(men_men_n1044_), .B(men_men_n1037_), .C(men_men_n257_), .Y(men_men_n1045_));
  INV        u1017(.A(men_men_n314_), .Y(men_men_n1046_));
  AOI210     u1018(.A0(men_men_n238_), .A1(men_men_n337_), .B0(men_men_n560_), .Y(men_men_n1047_));
  NA3        u1019(.A(men_men_n1047_), .B(men_men_n1046_), .C(men_men_n148_), .Y(men_men_n1048_));
  NO2        u1020(.A(men_men_n230_), .B(men_men_n175_), .Y(men_men_n1049_));
  NA2        u1021(.A(men_men_n1049_), .B(men_men_n415_), .Y(men_men_n1050_));
  NA3        u1022(.A(men_men_n173_), .B(men_men_n107_), .C(u), .Y(men_men_n1051_));
  NA3        u1023(.A(men_men_n454_), .B(men_men_n39_), .C(f), .Y(men_men_n1052_));
  NOi31      u1024(.An(j), .B(men_men_n1052_), .C(men_men_n1051_), .Y(men_men_n1053_));
  NAi31      u1025(.An(men_men_n180_), .B(men_men_n787_), .C(men_men_n454_), .Y(men_men_n1054_));
  NAi31      u1026(.An(men_men_n1053_), .B(men_men_n1054_), .C(men_men_n1050_), .Y(men_men_n1055_));
  NO2        u1027(.A(men_men_n266_), .B(men_men_n74_), .Y(men_men_n1056_));
  NO3        u1028(.A(men_men_n414_), .B(men_men_n766_), .C(n), .Y(men_men_n1057_));
  AOI210     u1029(.A0(men_men_n1057_), .A1(men_men_n1056_), .B0(men_men_n967_), .Y(men_men_n1058_));
  NAi31      u1030(.An(men_men_n939_), .B(men_men_n1058_), .C(men_men_n73_), .Y(men_men_n1059_));
  NO4        u1031(.A(men_men_n1059_), .B(men_men_n1055_), .C(men_men_n1048_), .D(men_men_n506_), .Y(men_men_n1060_));
  AN3        u1032(.A(men_men_n1060_), .B(men_men_n1045_), .C(men_men_n1036_), .Y(men_men_n1061_));
  NA2        u1033(.A(men_men_n524_), .B(men_men_n97_), .Y(men_men_n1062_));
  NA3        u1034(.A(men_men_n992_), .B(men_men_n580_), .C(men_men_n453_), .Y(men_men_n1063_));
  NA4        u1035(.A(men_men_n1063_), .B(men_men_n548_), .C(men_men_n1062_), .D(men_men_n233_), .Y(men_men_n1064_));
  NA2        u1036(.A(men_men_n988_), .B(men_men_n524_), .Y(men_men_n1065_));
  NA4        u1037(.A(men_men_n620_), .B(men_men_n199_), .C(men_men_n215_), .D(men_men_n157_), .Y(men_men_n1066_));
  NA3        u1038(.A(men_men_n1066_), .B(men_men_n1065_), .C(men_men_n289_), .Y(men_men_n1067_));
  OAI210     u1039(.A0(men_men_n452_), .A1(men_men_n114_), .B0(men_men_n791_), .Y(men_men_n1068_));
  AOI220     u1040(.A0(men_men_n1068_), .A1(men_men_n1016_), .B0(men_men_n547_), .B1(men_men_n396_), .Y(men_men_n1069_));
  OR4        u1041(.A(men_men_n937_), .B(men_men_n262_), .C(men_men_n217_), .D(e), .Y(men_men_n1070_));
  NO2        u1042(.A(men_men_n211_), .B(men_men_n208_), .Y(men_men_n1071_));
  NA2        u1043(.A(n), .B(e), .Y(men_men_n1072_));
  NO2        u1044(.A(men_men_n1072_), .B(men_men_n140_), .Y(men_men_n1073_));
  AOI220     u1045(.A0(men_men_n1073_), .A1(men_men_n264_), .B0(men_men_n781_), .B1(men_men_n1071_), .Y(men_men_n1074_));
  OAI210     u1046(.A0(men_men_n345_), .A1(men_men_n304_), .B0(men_men_n436_), .Y(men_men_n1075_));
  NA4        u1047(.A(men_men_n1075_), .B(men_men_n1074_), .C(men_men_n1070_), .D(men_men_n1069_), .Y(men_men_n1076_));
  AOI210     u1048(.A0(men_men_n1073_), .A1(men_men_n783_), .B0(men_men_n757_), .Y(men_men_n1077_));
  AOI220     u1049(.A0(men_men_n853_), .A1(men_men_n1357_), .B0(men_men_n620_), .B1(men_men_n235_), .Y(men_men_n1078_));
  NO2        u1050(.A(men_men_n67_), .B(h), .Y(men_men_n1079_));
  NO2        u1051(.A(men_men_n937_), .B(men_men_n679_), .Y(men_men_n1080_));
  NO2        u1052(.A(men_men_n964_), .B(men_men_n126_), .Y(men_men_n1081_));
  AN2        u1053(.A(men_men_n1081_), .B(men_men_n976_), .Y(men_men_n1082_));
  OAI210     u1054(.A0(men_men_n1082_), .A1(men_men_n1080_), .B0(men_men_n1079_), .Y(men_men_n1083_));
  NA4        u1055(.A(men_men_n1083_), .B(men_men_n1078_), .C(men_men_n1077_), .D(men_men_n793_), .Y(men_men_n1084_));
  NO4        u1056(.A(men_men_n1084_), .B(men_men_n1076_), .C(men_men_n1067_), .D(men_men_n1064_), .Y(men_men_n1085_));
  NA2        u1057(.A(men_men_n771_), .B(men_men_n705_), .Y(men_men_n1086_));
  NA4        u1058(.A(men_men_n1086_), .B(men_men_n1085_), .C(men_men_n1061_), .D(men_men_n1031_), .Y(men01));
  NO3        u1059(.A(men_men_n742_), .B(men_men_n468_), .C(men_men_n273_), .Y(men_men_n1088_));
  NA2        u1060(.A(men_men_n1088_), .B(men_men_n919_), .Y(men_men_n1089_));
  NA2        u1061(.A(men_men_n569_), .B(men_men_n85_), .Y(men_men_n1090_));
  NA2        u1062(.A(men_men_n541_), .B(men_men_n261_), .Y(men_men_n1091_));
  NA2        u1063(.A(men_men_n860_), .B(men_men_n1091_), .Y(men_men_n1092_));
  NA4        u1064(.A(men_men_n1092_), .B(men_men_n1090_), .C(men_men_n816_), .D(men_men_n325_), .Y(men_men_n1093_));
  NA2        u1065(.A(men_men_n663_), .B(men_men_n92_), .Y(men_men_n1094_));
  NO2        u1066(.A(men_men_n1094_), .B(i), .Y(men_men_n1095_));
  OAI210     u1067(.A0(men_men_n726_), .A1(n), .B0(men_men_n1066_), .Y(men_men_n1096_));
  INV        u1068(.A(men_men_n1096_), .Y(men_men_n1097_));
  NA2        u1069(.A(men_men_n112_), .B(l), .Y(men_men_n1098_));
  OR2        u1070(.A(men_men_n631_), .B(men_men_n357_), .Y(men_men_n1099_));
  NAi31      u1071(.An(men_men_n156_), .B(men_men_n1099_), .C(men_men_n1097_), .Y(men_men_n1100_));
  NA3        u1072(.A(men_men_n188_), .B(men_men_n641_), .C(men_men_n131_), .Y(men_men_n1101_));
  NO4        u1073(.A(men_men_n1101_), .B(men_men_n1100_), .C(men_men_n1093_), .D(men_men_n1089_), .Y(men_men_n1102_));
  NA2        u1074(.A(men_men_n1038_), .B(men_men_n200_), .Y(men_men_n1103_));
  OAI210     u1075(.A0(men_men_n1103_), .A1(men_men_n294_), .B0(men_men_n519_), .Y(men_men_n1104_));
  NO2        u1076(.A(men_men_n566_), .B(men_men_n1355_), .Y(men_men_n1105_));
  INV        u1077(.A(men_men_n1105_), .Y(men_men_n1106_));
  AOI210     u1078(.A0(men_men_n197_), .A1(men_men_n84_), .B0(men_men_n207_), .Y(men_men_n1107_));
  INV        u1079(.A(men_men_n1107_), .Y(men_men_n1108_));
  AN3        u1080(.A(m), .B(l), .C(k), .Y(men_men_n1109_));
  OAI210     u1081(.A0(men_men_n347_), .A1(men_men_n33_), .B0(men_men_n1109_), .Y(men_men_n1110_));
  NA2        u1082(.A(men_men_n196_), .B(men_men_n33_), .Y(men_men_n1111_));
  AO210      u1083(.A0(men_men_n1111_), .A1(men_men_n1110_), .B0(men_men_n324_), .Y(men_men_n1112_));
  NA4        u1084(.A(men_men_n1112_), .B(men_men_n1108_), .C(men_men_n1106_), .D(men_men_n1104_), .Y(men_men_n1113_));
  AOI210     u1085(.A0(men_men_n573_), .A1(men_men_n112_), .B0(men_men_n576_), .Y(men_men_n1114_));
  OAI210     u1086(.A0(men_men_n1098_), .A1(men_men_n572_), .B0(men_men_n1114_), .Y(men_men_n1115_));
  OAI210     u1087(.A0(men_men_n1095_), .A1(men_men_n319_), .B0(m), .Y(men_men_n1116_));
  NA3        u1088(.A(men_men_n1116_), .B(men_men_n272_), .C(men_men_n729_), .Y(men_men_n1117_));
  NO3        u1089(.A(men_men_n1117_), .B(men_men_n1115_), .C(men_men_n1113_), .Y(men_men_n1118_));
  NA2        u1090(.A(men_men_n491_), .B(men_men_n57_), .Y(men_men_n1119_));
  NA3        u1091(.A(u), .B(men_men_n75_), .C(i), .Y(men_men_n1120_));
  NO2        u1092(.A(men_men_n1120_), .B(men_men_n876_), .Y(men_men_n1121_));
  NO2        u1093(.A(men_men_n1121_), .B(men_men_n1035_), .Y(men_men_n1122_));
  NA3        u1094(.A(men_men_n1122_), .B(men_men_n1119_), .C(men_men_n704_), .Y(men_men_n1123_));
  NO2        u1095(.A(men_men_n866_), .B(men_men_n223_), .Y(men_men_n1124_));
  NA2        u1096(.A(men_men_n554_), .B(m), .Y(men_men_n1125_));
  NO3        u1097(.A(k), .B(men_men_n293_), .C(men_men_n44_), .Y(men_men_n1126_));
  NA2        u1098(.A(men_men_n1126_), .B(men_men_n540_), .Y(men_men_n1127_));
  NA3        u1099(.A(men_men_n1127_), .B(men_men_n1125_), .C(men_men_n638_), .Y(men_men_n1128_));
  OR2        u1100(.A(men_men_n1038_), .B(men_men_n1032_), .Y(men_men_n1129_));
  NO2        u1101(.A(men_men_n357_), .B(men_men_n72_), .Y(men_men_n1130_));
  AOI210     u1102(.A0(men_men_n683_), .A1(men_men_n590_), .B0(men_men_n1130_), .Y(men_men_n1131_));
  NA3        u1103(.A(men_men_n1131_), .B(men_men_n1129_), .C(men_men_n373_), .Y(men_men_n1132_));
  NO3        u1104(.A(men_men_n1132_), .B(men_men_n1128_), .C(men_men_n1123_), .Y(men_men_n1133_));
  AN2        u1105(.A(i), .B(men_men_n661_), .Y(men_men_n1134_));
  NO3        u1106(.A(men_men_n974_), .B(men_men_n170_), .C(men_men_n82_), .Y(men_men_n1135_));
  NO2        u1107(.A(men_men_n588_), .B(men_men_n587_), .Y(men_men_n1136_));
  NO4        u1108(.A(men_men_n974_), .B(men_men_n1136_), .C(men_men_n168_), .D(men_men_n82_), .Y(men_men_n1137_));
  NO3        u1109(.A(men_men_n1137_), .B(men_men_n1135_), .C(men_men_n612_), .Y(men_men_n1138_));
  NA4        u1110(.A(men_men_n1138_), .B(men_men_n1133_), .C(men_men_n1118_), .D(men_men_n1102_), .Y(men06));
  NO2        u1111(.A(men_men_n395_), .B(men_men_n546_), .Y(men_men_n1140_));
  OAI210     u1112(.A0(men_men_n108_), .A1(m), .B0(men_men_n1140_), .Y(men_men_n1141_));
  OAI210     u1113(.A0(n), .A1(men_men_n1135_), .B0(men_men_n370_), .Y(men_men_n1142_));
  NO3        u1114(.A(men_men_n577_), .B(men_men_n747_), .C(men_men_n578_), .Y(men_men_n1143_));
  BUFFER     u1115(.A(men_men_n803_), .Y(men_men_n1144_));
  NA3        u1116(.A(men_men_n1144_), .B(men_men_n1142_), .C(men_men_n1141_), .Y(men_men_n1145_));
  NO3        u1117(.A(men_men_n1145_), .B(men_men_n1128_), .C(men_men_n246_), .Y(men_men_n1146_));
  AOI210     u1118(.A0(u), .A1(men_men_n1354_), .B0(men_men_n1124_), .Y(men_men_n1147_));
  INV        u1119(.A(men_men_n1134_), .Y(men_men_n1148_));
  AOI210     u1120(.A0(men_men_n1148_), .A1(men_men_n1147_), .B0(men_men_n330_), .Y(men_men_n1149_));
  OAI210     u1121(.A0(men_men_n84_), .A1(men_men_n39_), .B0(men_men_n641_), .Y(men_men_n1150_));
  NA2        u1122(.A(men_men_n1150_), .B(men_men_n350_), .Y(men_men_n1151_));
  NO2        u1123(.A(men_men_n581_), .B(men_men_n993_), .Y(men_men_n1152_));
  NO2        u1124(.A(men_men_n447_), .B(men_men_n239_), .Y(men_men_n1153_));
  NO2        u1125(.A(men_men_n1153_), .B(men_men_n1152_), .Y(men_men_n1154_));
  INV        u1126(.A(men_men_n576_), .Y(men_men_n1155_));
  NA3        u1127(.A(men_men_n1155_), .B(men_men_n1154_), .C(men_men_n1151_), .Y(men_men_n1156_));
  NO2        u1128(.A(men_men_n697_), .B(men_men_n355_), .Y(men_men_n1157_));
  NOi21      u1129(.An(men_men_n1157_), .B(men_men_n48_), .Y(men_men_n1158_));
  BUFFER     u1130(.A(men_men_n853_), .Y(men_men_n1159_));
  NO4        u1131(.A(men_men_n1159_), .B(men_men_n1158_), .C(men_men_n1156_), .D(men_men_n1149_), .Y(men_men_n1160_));
  NO2        u1132(.A(men_men_n741_), .B(men_men_n268_), .Y(men_men_n1161_));
  OAI220     u1133(.A0(men_men_n685_), .A1(men_men_n46_), .B0(men_men_n219_), .B1(men_men_n589_), .Y(men_men_n1162_));
  AOI220     u1134(.A0(men_men_n350_), .A1(men_men_n1162_), .B0(men_men_n1161_), .B1(m), .Y(men_men_n1163_));
  NO3        u1135(.A(h), .B(men_men_n98_), .C(men_men_n275_), .Y(men_men_n1164_));
  NO2        u1136(.A(men_men_n575_), .B(j), .Y(men_men_n1165_));
  NOi21      u1137(.An(men_men_n1165_), .B(men_men_n72_), .Y(men_men_n1166_));
  NO3        u1138(.A(men_men_n1166_), .B(men_men_n1164_), .C(men_men_n996_), .Y(men_men_n1167_));
  NAi21      u1139(.An(men_men_n697_), .B(men_men_n196_), .Y(men_men_n1168_));
  NA4        u1140(.A(men_men_n1168_), .B(men_men_n1167_), .C(men_men_n1163_), .D(men_men_n1078_), .Y(men_men_n1169_));
  NOi31      u1141(.An(men_men_n1143_), .B(men_men_n451_), .C(men_men_n381_), .Y(men_men_n1170_));
  OR3        u1142(.A(men_men_n1170_), .B(men_men_n726_), .C(men_men_n530_), .Y(men_men_n1171_));
  NA2        u1143(.A(men_men_n1165_), .B(men_men_n733_), .Y(men_men_n1172_));
  NA2        u1144(.A(men_men_n1172_), .B(men_men_n1171_), .Y(men_men_n1173_));
  AN2        u1145(.A(men_men_n826_), .B(men_men_n825_), .Y(men_men_n1174_));
  NO3        u1146(.A(men_men_n1174_), .B(men_men_n796_), .C(men_men_n487_), .Y(men_men_n1175_));
  INV        u1147(.A(men_men_n1175_), .Y(men_men_n1176_));
  NO4        u1148(.A(men_men_n1136_), .B(j), .C(men_men_n430_), .D(men_men_n226_), .Y(men_men_n1177_));
  NO4        u1149(.A(men_men_n1177_), .B(men_men_n1176_), .C(men_men_n1173_), .D(men_men_n1169_), .Y(men_men_n1178_));
  NA4        u1150(.A(men_men_n1178_), .B(men_men_n1160_), .C(men_men_n1146_), .D(men_men_n1138_), .Y(men07));
  NOi21      u1151(.An(j), .B(k), .Y(men_men_n1180_));
  NAi32      u1152(.An(m), .Bn(b), .C(n), .Y(men_men_n1181_));
  NAi21      u1153(.An(f), .B(c), .Y(men_men_n1182_));
  OR2        u1154(.A(e), .B(d), .Y(men_men_n1183_));
  NOi31      u1155(.An(n), .B(m), .C(b), .Y(men_men_n1184_));
  NOi41      u1156(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1185_));
  NA3        u1157(.A(men_men_n1185_), .B(men_men_n794_), .C(men_men_n397_), .Y(men_men_n1186_));
  NO2        u1158(.A(men_men_n1186_), .B(men_men_n55_), .Y(men_men_n1187_));
  NA2        u1159(.A(men_men_n976_), .B(men_men_n215_), .Y(men_men_n1188_));
  NO2        u1160(.A(men_men_n1188_), .B(men_men_n60_), .Y(men_men_n1189_));
  NO2        u1161(.A(k), .B(i), .Y(men_men_n1190_));
  NA2        u1162(.A(men_men_n82_), .B(men_men_n44_), .Y(men_men_n1191_));
  NO2        u1163(.A(men_men_n942_), .B(men_men_n430_), .Y(men_men_n1192_));
  NA3        u1164(.A(men_men_n1192_), .B(men_men_n1191_), .C(men_men_n208_), .Y(men_men_n1193_));
  NO2        u1165(.A(men_men_n952_), .B(men_men_n298_), .Y(men_men_n1194_));
  NA2        u1166(.A(men_men_n531_), .B(men_men_n79_), .Y(men_men_n1195_));
  NA2        u1167(.A(men_men_n1079_), .B(men_men_n283_), .Y(men_men_n1196_));
  NA3        u1168(.A(men_men_n1196_), .B(men_men_n1195_), .C(men_men_n1193_), .Y(men_men_n1197_));
  NO3        u1169(.A(men_men_n1197_), .B(men_men_n1189_), .C(men_men_n1187_), .Y(men_men_n1198_));
  OR2        u1170(.A(h), .B(f), .Y(men_men_n1199_));
  NO3        u1171(.A(n), .B(m), .C(i), .Y(men_men_n1200_));
  OAI210     u1172(.A0(men_men_n994_), .A1(men_men_n151_), .B0(men_men_n1200_), .Y(men_men_n1201_));
  NO2        u1173(.A(i), .B(u), .Y(men_men_n1202_));
  OR3        u1174(.A(men_men_n1202_), .B(men_men_n1181_), .C(men_men_n71_), .Y(men_men_n1203_));
  OAI220     u1175(.A0(men_men_n1203_), .A1(men_men_n472_), .B0(men_men_n1201_), .B1(men_men_n1199_), .Y(men_men_n1204_));
  NA2        u1176(.A(men_men_n653_), .B(men_men_n107_), .Y(men_men_n1205_));
  NA3        u1177(.A(men_men_n1184_), .B(men_men_n948_), .C(h), .Y(men_men_n1206_));
  AOI210     u1178(.A0(men_men_n1206_), .A1(men_men_n1205_), .B0(men_men_n44_), .Y(men_men_n1207_));
  NA2        u1179(.A(men_men_n1200_), .B(men_men_n614_), .Y(men_men_n1208_));
  NO3        u1180(.A(men_men_n430_), .B(d), .C(c), .Y(men_men_n1209_));
  NO2        u1181(.A(men_men_n1207_), .B(men_men_n1204_), .Y(men_men_n1210_));
  NO2        u1182(.A(men_men_n141_), .B(h), .Y(men_men_n1211_));
  NO2        u1183(.A(u), .B(c), .Y(men_men_n1212_));
  NO2        u1184(.A(men_men_n441_), .B(a), .Y(men_men_n1213_));
  NA3        u1185(.A(men_men_n1213_), .B(men_men_n1350_), .C(men_men_n108_), .Y(men_men_n1214_));
  NO2        u1186(.A(i), .B(h), .Y(men_men_n1215_));
  NA2        u1187(.A(men_men_n1215_), .B(men_men_n215_), .Y(men_men_n1216_));
  AOI210     u1188(.A0(men_men_n247_), .A1(men_men_n110_), .B0(men_men_n519_), .Y(men_men_n1217_));
  NO2        u1189(.A(men_men_n1217_), .B(men_men_n1216_), .Y(men_men_n1218_));
  NO2        u1190(.A(men_men_n703_), .B(men_men_n182_), .Y(men_men_n1219_));
  NOi31      u1191(.An(f), .B(d), .C(c), .Y(men_men_n1220_));
  NO2        u1192(.A(men_men_n1219_), .B(men_men_n1218_), .Y(men_men_n1221_));
  NA2        u1193(.A(men_men_n514_), .B(men_men_n949_), .Y(men_men_n1222_));
  NO3        u1194(.A(men_men_n40_), .B(i), .C(h), .Y(men_men_n1223_));
  AN3        u1195(.A(men_men_n1222_), .B(men_men_n1221_), .C(men_men_n1214_), .Y(men_men_n1224_));
  NA2        u1196(.A(men_men_n1184_), .B(men_men_n367_), .Y(men_men_n1225_));
  NO2        u1197(.A(men_men_n1225_), .B(men_men_n935_), .Y(men_men_n1226_));
  NO2        u1198(.A(men_men_n182_), .B(b), .Y(men_men_n1227_));
  NA2        u1199(.A(men_men_n1033_), .B(men_men_n1227_), .Y(men_men_n1228_));
  NO2        u1200(.A(i), .B(men_men_n207_), .Y(men_men_n1229_));
  NA4        u1201(.A(men_men_n1015_), .B(men_men_n1229_), .C(men_men_n99_), .D(m), .Y(men_men_n1230_));
  NAi31      u1202(.An(men_men_n1226_), .B(men_men_n1230_), .C(men_men_n1228_), .Y(men_men_n1231_));
  NO4        u1203(.A(men_men_n126_), .B(u), .C(f), .D(e), .Y(men_men_n1232_));
  NA2        u1204(.A(men_men_n187_), .B(men_men_n94_), .Y(men_men_n1233_));
  OR2        u1205(.A(e), .B(a), .Y(men_men_n1234_));
  NA2        u1206(.A(men_men_n30_), .B(h), .Y(men_men_n1235_));
  NO2        u1207(.A(men_men_n1235_), .B(men_men_n966_), .Y(men_men_n1236_));
  NOi41      u1208(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1237_));
  NA2        u1209(.A(men_men_n1237_), .B(men_men_n108_), .Y(men_men_n1238_));
  INV        u1210(.A(men_men_n1238_), .Y(men_men_n1239_));
  OR3        u1211(.A(men_men_n530_), .B(men_men_n529_), .C(men_men_n107_), .Y(men_men_n1240_));
  NA2        u1212(.A(men_men_n992_), .B(men_men_n394_), .Y(men_men_n1241_));
  OAI220     u1213(.A0(men_men_n1241_), .A1(men_men_n423_), .B0(men_men_n1240_), .B1(men_men_n293_), .Y(men_men_n1242_));
  AO210      u1214(.A0(men_men_n1242_), .A1(men_men_n110_), .B0(men_men_n1239_), .Y(men_men_n1243_));
  NO3        u1215(.A(men_men_n1243_), .B(men_men_n1236_), .C(men_men_n1231_), .Y(men_men_n1244_));
  NA4        u1216(.A(men_men_n1244_), .B(men_men_n1224_), .C(men_men_n1210_), .D(men_men_n1198_), .Y(men_men_n1245_));
  NO2        u1217(.A(men_men_n1004_), .B(men_men_n105_), .Y(men_men_n1246_));
  NA2        u1218(.A(men_men_n367_), .B(men_men_n55_), .Y(men_men_n1247_));
  AOI210     u1219(.A0(men_men_n1247_), .A1(men_men_n942_), .B0(men_men_n1208_), .Y(men_men_n1248_));
  NA2        u1220(.A(men_men_n209_), .B(men_men_n173_), .Y(men_men_n1249_));
  AOI210     u1221(.A0(men_men_n1249_), .A1(men_men_n1051_), .B0(men_men_n1247_), .Y(men_men_n1250_));
  NO2        u1222(.A(men_men_n970_), .B(men_men_n966_), .Y(men_men_n1251_));
  NO3        u1223(.A(men_men_n1251_), .B(men_men_n1250_), .C(men_men_n1248_), .Y(men_men_n1252_));
  NA2        u1224(.A(men_men_n1223_), .B(men_men_n1183_), .Y(men_men_n1253_));
  NO3        u1225(.A(men_men_n966_), .B(men_men_n563_), .C(u), .Y(men_men_n1254_));
  NOi21      u1226(.An(men_men_n1249_), .B(men_men_n1254_), .Y(men_men_n1255_));
  AOI210     u1227(.A0(men_men_n1255_), .A1(men_men_n1233_), .B0(men_men_n942_), .Y(men_men_n1256_));
  INV        u1228(.A(men_men_n48_), .Y(men_men_n1257_));
  AOI220     u1229(.A0(men_men_n1257_), .A1(men_men_n1040_), .B0(men_men_n760_), .B1(men_men_n187_), .Y(men_men_n1258_));
  INV        u1230(.A(men_men_n1258_), .Y(men_men_n1259_));
  OAI220     u1231(.A0(men_men_n636_), .A1(u), .B0(men_men_n219_), .B1(c), .Y(men_men_n1260_));
  AOI210     u1232(.A0(men_men_n1227_), .A1(men_men_n40_), .B0(men_men_n1260_), .Y(men_men_n1261_));
  NO2        u1233(.A(men_men_n126_), .B(l), .Y(men_men_n1262_));
  NO2        u1234(.A(men_men_n219_), .B(k), .Y(men_men_n1263_));
  OAI210     u1235(.A0(men_men_n1263_), .A1(men_men_n1215_), .B0(men_men_n1262_), .Y(men_men_n1264_));
  OAI220     u1236(.A0(men_men_n1264_), .A1(e), .B0(men_men_n1261_), .B1(men_men_n170_), .Y(men_men_n1265_));
  NO3        u1237(.A(men_men_n1240_), .B(men_men_n454_), .C(men_men_n342_), .Y(men_men_n1266_));
  NO4        u1238(.A(men_men_n1266_), .B(men_men_n1265_), .C(men_men_n1259_), .D(men_men_n1256_), .Y(men_men_n1267_));
  NO2        u1239(.A(men_men_n48_), .B(men_men_n563_), .Y(men_men_n1268_));
  NA2        u1240(.A(men_men_n979_), .B(men_men_n1268_), .Y(men_men_n1269_));
  NO2        u1241(.A(men_men_n966_), .B(h), .Y(men_men_n1270_));
  NO2        u1242(.A(men_men_n1269_), .B(j), .Y(men_men_n1271_));
  NA3        u1243(.A(men_men_n1246_), .B(men_men_n454_), .C(f), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n1180_), .B(men_men_n41_), .Y(men_men_n1273_));
  AOI210     u1245(.A0(men_men_n108_), .A1(men_men_n39_), .B0(men_men_n1273_), .Y(men_men_n1274_));
  NO2        u1246(.A(men_men_n1274_), .B(men_men_n1272_), .Y(men_men_n1275_));
  AOI210     u1247(.A0(men_men_n514_), .A1(h), .B0(men_men_n68_), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n1276_), .B(men_men_n1213_), .Y(men_men_n1277_));
  NO2        u1249(.A(j), .B(men_men_n168_), .Y(men_men_n1278_));
  NOi21      u1250(.An(d), .B(f), .Y(men_men_n1279_));
  NO3        u1251(.A(men_men_n1220_), .B(men_men_n1279_), .C(men_men_n39_), .Y(men_men_n1280_));
  NA2        u1252(.A(men_men_n1280_), .B(men_men_n1278_), .Y(men_men_n1281_));
  NO2        u1253(.A(men_men_n1183_), .B(f), .Y(men_men_n1282_));
  NA2        u1254(.A(men_men_n1213_), .B(men_men_n1273_), .Y(men_men_n1283_));
  NO2        u1255(.A(men_men_n293_), .B(c), .Y(men_men_n1284_));
  NA2        u1256(.A(men_men_n1284_), .B(men_men_n531_), .Y(men_men_n1285_));
  NA4        u1257(.A(men_men_n1285_), .B(men_men_n1283_), .C(men_men_n1281_), .D(men_men_n1277_), .Y(men_men_n1286_));
  NO3        u1258(.A(men_men_n1286_), .B(men_men_n1275_), .C(men_men_n1271_), .Y(men_men_n1287_));
  NA4        u1259(.A(men_men_n1287_), .B(men_men_n1267_), .C(men_men_n1253_), .D(men_men_n1252_), .Y(men_men_n1288_));
  OAI220     u1260(.A0(men_men_n454_), .A1(men_men_n293_), .B0(men_men_n125_), .B1(men_men_n58_), .Y(men_men_n1289_));
  NA2        u1261(.A(men_men_n1289_), .B(men_men_n1194_), .Y(men_men_n1290_));
  INV        u1262(.A(men_men_n1290_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n1212_), .B(men_men_n1279_), .Y(men_men_n1292_));
  NO2        u1264(.A(men_men_n1292_), .B(m), .Y(men_men_n1293_));
  NA3        u1265(.A(men_men_n976_), .B(men_men_n103_), .C(men_men_n215_), .Y(men_men_n1294_));
  INV        u1266(.A(men_men_n1294_), .Y(men_men_n1295_));
  NO3        u1267(.A(men_men_n1295_), .B(men_men_n1293_), .C(men_men_n1291_), .Y(men_men_n1296_));
  NO2        u1268(.A(men_men_n1182_), .B(e), .Y(men_men_n1297_));
  NA2        u1269(.A(men_men_n1297_), .B(men_men_n392_), .Y(men_men_n1298_));
  NA2        u1270(.A(men_men_n999_), .B(men_men_n605_), .Y(men_men_n1299_));
  OR3        u1271(.A(men_men_n1263_), .B(men_men_n1079_), .C(men_men_n126_), .Y(men_men_n1300_));
  OAI220     u1272(.A0(men_men_n1300_), .A1(men_men_n1298_), .B0(men_men_n1299_), .B1(men_men_n432_), .Y(men_men_n1301_));
  NO3        u1273(.A(men_men_n1240_), .B(men_men_n342_), .C(a), .Y(men_men_n1302_));
  NO2        u1274(.A(men_men_n1302_), .B(men_men_n1301_), .Y(men_men_n1303_));
  NA2        u1275(.A(men_men_n529_), .B(u), .Y(men_men_n1304_));
  NA2        u1276(.A(men_men_n1304_), .B(men_men_n1209_), .Y(men_men_n1305_));
  NO2        u1277(.A(men_men_n1234_), .B(f), .Y(men_men_n1306_));
  NO2        u1278(.A(men_men_n1305_), .B(men_men_n207_), .Y(men_men_n1307_));
  NA2        u1279(.A(men_men_n1306_), .B(men_men_n1191_), .Y(men_men_n1308_));
  NO2        u1280(.A(men_men_n1308_), .B(men_men_n48_), .Y(men_men_n1309_));
  NO2        u1281(.A(men_men_n48_), .B(l), .Y(men_men_n1310_));
  NA2        u1282(.A(men_men_n979_), .B(men_men_n1310_), .Y(men_men_n1311_));
  NO2        u1283(.A(men_men_n242_), .B(u), .Y(men_men_n1312_));
  NO2        u1284(.A(m), .B(i), .Y(men_men_n1313_));
  AOI220     u1285(.A0(men_men_n1313_), .A1(men_men_n1211_), .B0(men_men_n958_), .B1(men_men_n1312_), .Y(men_men_n1314_));
  NA2        u1286(.A(men_men_n1314_), .B(men_men_n1311_), .Y(men_men_n1315_));
  NO3        u1287(.A(men_men_n1315_), .B(men_men_n1309_), .C(men_men_n1307_), .Y(men_men_n1316_));
  NA3        u1288(.A(men_men_n1316_), .B(men_men_n1303_), .C(men_men_n1296_), .Y(men_men_n1317_));
  NA3        u1289(.A(men_men_n859_), .B(men_men_n132_), .C(men_men_n45_), .Y(men_men_n1318_));
  AOI210     u1290(.A0(men_men_n142_), .A1(c), .B0(men_men_n1318_), .Y(men_men_n1319_));
  OAI210     u1291(.A0(men_men_n563_), .A1(u), .B0(men_men_n179_), .Y(men_men_n1320_));
  NA2        u1292(.A(men_men_n1320_), .B(men_men_n1270_), .Y(men_men_n1321_));
  NO2        u1293(.A(men_men_n71_), .B(c), .Y(men_men_n1322_));
  NO4        u1294(.A(men_men_n1199_), .B(men_men_n180_), .C(men_men_n438_), .D(men_men_n44_), .Y(men_men_n1323_));
  AOI210     u1295(.A0(men_men_n1278_), .A1(men_men_n1322_), .B0(men_men_n1323_), .Y(men_men_n1324_));
  NA2        u1296(.A(men_men_n1324_), .B(men_men_n1321_), .Y(men_men_n1325_));
  NO2        u1297(.A(men_men_n1325_), .B(men_men_n1319_), .Y(men_men_n1326_));
  NO2        u1298(.A(men_men_n1318_), .B(men_men_n105_), .Y(men_men_n1327_));
  INV        u1299(.A(men_men_n1327_), .Y(men_men_n1328_));
  AN2        u1300(.A(men_men_n976_), .B(men_men_n964_), .Y(men_men_n1329_));
  AOI220     u1301(.A0(men_men_n1313_), .A1(men_men_n614_), .B0(men_men_n1351_), .B1(men_men_n154_), .Y(men_men_n1330_));
  NOi31      u1302(.An(men_men_n30_), .B(men_men_n1330_), .C(n), .Y(men_men_n1331_));
  AOI210     u1303(.A0(men_men_n1329_), .A1(men_men_n1033_), .B0(men_men_n1331_), .Y(men_men_n1332_));
  NO2        u1304(.A(men_men_n1272_), .B(men_men_n68_), .Y(men_men_n1333_));
  NO2        u1305(.A(men_men_n1190_), .B(men_men_n112_), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n1334_), .B(men_men_n1225_), .Y(men_men_n1335_));
  NO2        u1307(.A(men_men_n1335_), .B(men_men_n1333_), .Y(men_men_n1336_));
  NA4        u1308(.A(men_men_n1336_), .B(men_men_n1332_), .C(men_men_n1328_), .D(men_men_n1326_), .Y(men_men_n1337_));
  OR4        u1309(.A(men_men_n1337_), .B(men_men_n1317_), .C(men_men_n1288_), .D(men_men_n1245_), .Y(men04));
  NOi21      u1310(.An(men_men_n1232_), .B(men_men_n937_), .Y(men_men_n1339_));
  NA2        u1311(.A(men_men_n1282_), .B(men_men_n760_), .Y(men_men_n1340_));
  NO4        u1312(.A(men_men_n1340_), .B(men_men_n1358_), .C(men_men_n473_), .D(j), .Y(men_men_n1341_));
  OR3        u1313(.A(men_men_n1341_), .B(men_men_n1339_), .C(men_men_n951_), .Y(men_men_n1342_));
  NO3        u1314(.A(men_men_n1191_), .B(men_men_n86_), .C(k), .Y(men_men_n1343_));
  AOI210     u1315(.A0(men_men_n1343_), .A1(men_men_n945_), .B0(men_men_n1053_), .Y(men_men_n1344_));
  NA2        u1316(.A(men_men_n1344_), .B(men_men_n1083_), .Y(men_men_n1345_));
  NO4        u1317(.A(men_men_n1345_), .B(men_men_n1342_), .C(men_men_n956_), .D(men_men_n941_), .Y(men_men_n1346_));
  NA4        u1318(.A(men_men_n1346_), .B(men_men_n1001_), .C(men_men_n990_), .D(men_men_n982_), .Y(men05));
  INV        u1319(.A(i), .Y(men_men_n1350_));
  INV        u1320(.A(j), .Y(men_men_n1351_));
  INV        u1321(.A(men_men_n519_), .Y(men_men_n1352_));
  INV        u1322(.A(men_men_n215_), .Y(men_men_n1353_));
  INV        u1323(.A(f), .Y(men_men_n1354_));
  INV        u1324(.A(i), .Y(men_men_n1355_));
  INV        u1325(.A(n), .Y(men_men_n1356_));
  INV        u1326(.A(c), .Y(men_men_n1357_));
  INV        u1327(.A(c), .Y(men_men_n1358_));
  INV        u1328(.A(f), .Y(men_men_n1359_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule