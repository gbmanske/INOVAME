`timescale 1 ns/10 ps

`define assert(index, dut_sum, exp_sum, dut_cout, exp_cout, message) \
	if (dut_sum !== exp_sum) begin \
		$display("ERROR in %m: %d != %d",dut_sum,exp_sum); \
		$display(message); \
	end \
	else if (dut_cout !== exp_cout) begin \
		$display("ERROR in %m: %d != %d",dut_cout,exp_cout); \
		$display(message); \
	end \
	else \
	begin \
		$display("Teste %01d correto: %d == %d",index,dut_sum,exp_sum); \
	end
	
module tb_adder;

	localparam WIDTH=16;

    logic [WIDTH-1:0] A, B;
    logic Cin;
    logic [WIDTH-1:0] S;
    logic Cout;


	cla_16bits DUT(.A(A),.B(B),.Cin(Cin),.S(S),.Cout(Cout));


	initial begin
		$dumpfile("sad.vcd");
		$dumpvars(0,tb_adder);

	//-----------------------------------------------------------Teste 1----------------------------------------------//
		
		A = 'd0;
		B = 'd0;
        Cin = 1'b0;
		#5
		`assert(1,S,'d0,Cout,1'd0,"S!=0")
		#1

	//-----------------------------------------------------------Teste 2----------------------------------------------//
		
        A = 'd500;
		B = 'd499;
        Cin = 1'b1;
		#5
		`assert(2,S,'d1000,Cout,1'd0,"S!=1000")
		#1
		
	//-----------------------------------------------------------Teste 3---------------------------------------------//
		
		A = 'd65535;
		B = 'd1;
        Cin = 1'b0;
		#5
		`assert(3,S,'d0,Cout,1'd1,"S!=0")
		#1
		
	//-----------------------------------------------------------Teste 4----------------------------------------------//'
		
		A = 'd50505;
		B = 'd5050;
        Cin = 1'b0;
		#5
		`assert(4,S,'d55555,Cout,1'd0,"S!=55555")
		#1
	
	//-----------------------------------------------------------Teste 5----------------------------------------------//
		
        A = 'd500;
		B = 'd499;
        Cin = 1'b0;
		#5
		`assert(5,S,'d999,Cout,1'd0,"S!=999")
		#1	
	//-----------------------------------------------------------Teste 6----------------------------------------------//
		
        A = 'd5050;
		B = 'd50505;
        Cin = 1'b0;
		#5
		`assert(4,S,'d55555,Cout,1'd0,"S!=55555")
		#1	
	//-----------------------------------------------------------Teste 7----------------------------------------------//
		
        A = 'd0;
		B = 'd49999;
        Cin = 1'b0;
		#5
		`assert(7,S,'d49999,Cout,1'd0,"S!=49999")
		#1	
	//-----------------------------------------------------------Teste 8----------------------------------------------//
		
        A = 'd5000;
		B = 'd499;
        Cin = 1'b0;
		#5
		`assert(8,S,'d5499,Cout,1'd0,"S!=5499")
		#1	
		
		//------------------------------------------------------Teste 9----------------------------------------------//
		
        A = 'd1;
		B = 'd0;
        Cin = 1'b0;
		#5
		`assert(9,S,'d1,Cout,1'd0,"S!=1")
		#1	

	//-----------------------------------------------------------Teste 10----------------------------------------------//
		
        A = 'd0;
		B = 'd1;
        Cin = 1'b0;
		#5
		`assert(10,S,'d1,Cout,1'd0,"S!=1")
		#1	

	//-----------------------------------------------------------Teste 11----------------------------------------------//
		
        A = 'd1;
		B = 'd1;
        Cin = 1'b0;
		#5
		`assert(11,S,'d2,Cout,1'd0,"S!=2")
		#1	

	//-----------------------------------------------------------Teste 12----------------------------------------------//
		
        A = 'd0;
		B = 'd2;
        Cin = 1'b0;
		#5
		`assert(12,S,'d2,Cout,1'd0,"S!=2")
		#1	

	//-----------------------------------------------------------Teste 13----------------------------------------------//
		
        A = 'd1;
		B = 'd2;
        Cin = 1'b0;
		#5
		`assert(13,S,'d3,Cout,1'd0,"S!=3")
		#1	

	//-----------------------------------------------------------Teste 14----------------------------------------------//
		
        A = 'd2;
		B = 'd2;
        Cin = 1'b0;
		#5
		`assert(14,S,'d4,Cout,1'd0,"S!=4")
		#1	

	//-----------------------------------------------------------Teste 15----------------------------------------------//
		
        A = 'd3;
		B = 'd0;
        Cin = 1'b0;
		#5
		`assert(15,S,'d3,Cout,1'd0,"S!=3")
		#1	

	//-----------------------------------------------------------Teste 16----------------------------------------------//
		
        A = 'd3;
		B = 'd1;
        Cin = 1'b0;
		#5
		`assert(16,S,'d4,Cout,1'd0,"S!=4")
		#1	

	//-----------------------------------------------------------Teste 17----------------------------------------------//
		
        A = 'd3;
		B = 'd3;
        Cin = 1'b0;
		#5
		`assert(17,S,'d6,Cout,1'd0,"S!=6")
		#1	

	//-----------------------------------------------------------Teste 18----------------------------------------------//
		
        A = 'd3;
		B = 'd5;
        Cin = 1'b0;
		#5
		`assert(18,S,'d8,Cout,1'd0,"S!=8")
		#1	

	//-----------------------------------------------------------Teste 19----------------------------------------------//
		
        A = 'd8;
		B = 'd7;
        Cin = 1'b0;
		#5
		`assert(19,S,'d15,Cout,1'd0,"S!=15")
		#1	

	//-----------------------------------------------------------Teste 20----------------------------------------------//
		
        A = 'd11;
		B = 'd10;
        Cin = 1'b0;
		#5
		`assert(20,S,'d21,Cout,1'd0,"S!=21")
		#1	

	//-----------------------------------------------------------Teste 21----------------------------------------------//
		
        A = 'd5;
		B = 'd2;
        Cin = 1'b0;
		#5
		`assert(21,S,'d7,Cout,1'd0,"S!=7")
		#1	

	//-----------------------------------------------------------Teste 22----------------------------------------------//
		
        A = 'd499;
		B = 'd499;
        Cin = 1'b0;
		#5
		`assert(22,S,'d998,Cout,1'd0,"S!=998")
		#1	

	$stop;

end
endmodule
