library verilog;
use verilog.vl_types.all;
entity tb_pixel_interpolator is
end tb_pixel_interpolator;
