//Benchmark atmr_alu4_1266_0.125

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n125_, ori_ori_n126_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  INV        o024(.A(i_5_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_7_), .B(i_10_), .Y(ori_ori_n48_));
  AOI210     o026(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  OAI210     o027(.A0(ori_ori_n49_), .A1(i_3_), .B0(ori_ori_n47_), .Y(ori_ori_n50_));
  NO2        o028(.A(ori_ori_n50_), .B(ori_ori_n46_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_7_), .B(i_9_), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n51_), .B(ori_ori_n45_), .Y(ori_ori_n53_));
  NO2        o031(.A(i_1_), .B(i_6_), .Y(ori_ori_n54_));
  NAi21      o032(.An(i_2_), .B(i_7_), .Y(ori_ori_n55_));
  INV        o033(.A(i_1_), .Y(ori_ori_n56_));
  NA2        o034(.A(ori_ori_n56_), .B(i_6_), .Y(ori_ori_n57_));
  NA3        o035(.A(ori_ori_n57_), .B(ori_ori_n55_), .C(ori_ori_n31_), .Y(ori_ori_n58_));
  NA2        o036(.A(i_1_), .B(i_10_), .Y(ori_ori_n59_));
  NO2        o037(.A(ori_ori_n59_), .B(i_6_), .Y(ori_ori_n60_));
  NAi21      o038(.An(ori_ori_n60_), .B(ori_ori_n58_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n49_), .B(i_2_), .Y(ori_ori_n62_));
  AOI210     o040(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n63_));
  NA2        o041(.A(i_1_), .B(i_6_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(ori_ori_n25_), .Y(ori_ori_n65_));
  INV        o043(.A(i_0_), .Y(ori_ori_n66_));
  NAi21      o044(.An(i_5_), .B(i_10_), .Y(ori_ori_n67_));
  NA2        o045(.A(i_5_), .B(i_9_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(ori_ori_n68_), .A1(ori_ori_n67_), .B0(ori_ori_n66_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n65_), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n63_), .A1(ori_ori_n62_), .B0(ori_ori_n70_), .Y(ori_ori_n71_));
  OAI210     o049(.A0(ori_ori_n71_), .A1(ori_ori_n61_), .B0(i_0_), .Y(ori_ori_n72_));
  NA2        o050(.A(i_12_), .B(i_5_), .Y(ori_ori_n73_));
  NO2        o051(.A(i_3_), .B(i_9_), .Y(ori_ori_n74_));
  NO2        o052(.A(i_3_), .B(i_7_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n74_), .B(ori_ori_n56_), .Y(ori_ori_n76_));
  INV        o054(.A(i_6_), .Y(ori_ori_n77_));
  NO2        o055(.A(i_2_), .B(i_7_), .Y(ori_ori_n78_));
  INV        o056(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NA2        o057(.A(ori_ori_n76_), .B(ori_ori_n79_), .Y(ori_ori_n80_));
  NAi21      o058(.An(i_6_), .B(i_10_), .Y(ori_ori_n81_));
  NA2        o059(.A(i_6_), .B(i_9_), .Y(ori_ori_n82_));
  AOI210     o060(.A0(ori_ori_n82_), .A1(ori_ori_n81_), .B0(ori_ori_n56_), .Y(ori_ori_n83_));
  NA2        o061(.A(i_2_), .B(i_6_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n83_), .Y(ori_ori_n85_));
  AOI210     o063(.A0(ori_ori_n85_), .A1(ori_ori_n80_), .B0(ori_ori_n73_), .Y(ori_ori_n86_));
  AN3        o064(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n87_));
  NAi21      o065(.An(i_6_), .B(i_11_), .Y(ori_ori_n88_));
  NO2        o066(.A(i_5_), .B(i_8_), .Y(ori_ori_n89_));
  NOi21      o067(.An(ori_ori_n89_), .B(ori_ori_n88_), .Y(ori_ori_n90_));
  AOI220     o068(.A0(ori_ori_n90_), .A1(ori_ori_n55_), .B0(ori_ori_n87_), .B1(ori_ori_n32_), .Y(ori_ori_n91_));
  INV        o069(.A(i_7_), .Y(ori_ori_n92_));
  NA2        o070(.A(ori_ori_n46_), .B(ori_ori_n92_), .Y(ori_ori_n93_));
  NO2        o071(.A(i_0_), .B(i_5_), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n94_), .B(ori_ori_n77_), .Y(ori_ori_n95_));
  NA2        o073(.A(i_12_), .B(i_3_), .Y(ori_ori_n96_));
  INV        o074(.A(ori_ori_n96_), .Y(ori_ori_n97_));
  NA3        o075(.A(ori_ori_n97_), .B(ori_ori_n95_), .C(ori_ori_n93_), .Y(ori_ori_n98_));
  NAi21      o076(.An(i_7_), .B(i_11_), .Y(ori_ori_n99_));
  AN2        o077(.A(i_2_), .B(i_10_), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n100_), .B(i_7_), .Y(ori_ori_n101_));
  OR2        o079(.A(ori_ori_n73_), .B(ori_ori_n54_), .Y(ori_ori_n102_));
  NO2        o080(.A(i_8_), .B(ori_ori_n92_), .Y(ori_ori_n103_));
  NO3        o081(.A(ori_ori_n103_), .B(ori_ori_n102_), .C(ori_ori_n101_), .Y(ori_ori_n104_));
  NA2        o082(.A(i_12_), .B(i_7_), .Y(ori_ori_n105_));
  NA2        o083(.A(i_11_), .B(i_12_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n507_), .B(ori_ori_n104_), .Y(ori_ori_n107_));
  NA3        o085(.A(ori_ori_n107_), .B(ori_ori_n98_), .C(ori_ori_n91_), .Y(ori_ori_n108_));
  NOi21      o086(.An(i_1_), .B(i_5_), .Y(ori_ori_n109_));
  NA2        o087(.A(ori_ori_n109_), .B(i_11_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n92_), .B(ori_ori_n37_), .Y(ori_ori_n111_));
  NA2        o089(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n112_), .B(ori_ori_n111_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n113_), .B(ori_ori_n46_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n82_), .B(ori_ori_n81_), .Y(ori_ori_n115_));
  NAi21      o093(.An(i_3_), .B(i_8_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n116_), .B(ori_ori_n55_), .Y(ori_ori_n117_));
  NOi31      o095(.An(ori_ori_n117_), .B(ori_ori_n115_), .C(ori_ori_n114_), .Y(ori_ori_n118_));
  NO2        o096(.A(i_1_), .B(ori_ori_n77_), .Y(ori_ori_n119_));
  NO2        o097(.A(i_6_), .B(i_5_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(i_3_), .Y(ori_ori_n121_));
  OAI220     o099(.A0(ori_ori_n121_), .A1(ori_ori_n99_), .B0(ori_ori_n118_), .B1(ori_ori_n110_), .Y(ori_ori_n122_));
  NO3        o100(.A(ori_ori_n122_), .B(ori_ori_n108_), .C(ori_ori_n86_), .Y(ori_ori_n123_));
  NA3        o101(.A(ori_ori_n123_), .B(ori_ori_n72_), .C(ori_ori_n53_), .Y(ori2));
  NO2        o102(.A(ori_ori_n56_), .B(ori_ori_n37_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n505_), .B(ori_ori_n125_), .Y(ori_ori_n126_));
  NA4        o104(.A(ori_ori_n126_), .B(ori_ori_n70_), .C(ori_ori_n62_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o105(.A(i_0_), .B(i_1_), .Y(ori_ori_n128_));
  NA2        o106(.A(i_2_), .B(i_3_), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n129_), .B(i_4_), .Y(ori_ori_n130_));
  NA2        o108(.A(i_1_), .B(i_5_), .Y(ori_ori_n131_));
  OR2        o109(.A(i_0_), .B(i_1_), .Y(ori_ori_n132_));
  NO3        o110(.A(ori_ori_n132_), .B(ori_ori_n73_), .C(i_13_), .Y(ori_ori_n133_));
  NAi32      o111(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n134_));
  NAi21      o112(.An(ori_ori_n134_), .B(ori_ori_n133_), .Y(ori_ori_n135_));
  NOi21      o113(.An(i_4_), .B(i_10_), .Y(ori_ori_n136_));
  NOi21      o114(.An(i_4_), .B(i_9_), .Y(ori_ori_n137_));
  NOi21      o115(.An(i_11_), .B(i_13_), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n138_), .B(ori_ori_n137_), .Y(ori_ori_n139_));
  NO2        o117(.A(ori_ori_n66_), .B(ori_ori_n56_), .Y(ori_ori_n140_));
  NO2        o118(.A(ori_ori_n66_), .B(i_5_), .Y(ori_ori_n141_));
  NO2        o119(.A(i_2_), .B(i_1_), .Y(ori_ori_n142_));
  NAi21      o120(.An(i_4_), .B(i_12_), .Y(ori_ori_n143_));
  INV        o121(.A(i_8_), .Y(ori_ori_n144_));
  NO2        o122(.A(i_3_), .B(i_8_), .Y(ori_ori_n145_));
  NO3        o123(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n146_));
  NO2        o124(.A(ori_ori_n94_), .B(ori_ori_n54_), .Y(ori_ori_n147_));
  NO2        o125(.A(i_13_), .B(i_9_), .Y(ori_ori_n148_));
  NAi21      o126(.An(i_12_), .B(i_3_), .Y(ori_ori_n149_));
  NO2        o127(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n150_));
  NA2        o128(.A(i_0_), .B(i_5_), .Y(ori_ori_n151_));
  INV        o129(.A(i_13_), .Y(ori_ori_n152_));
  NO2        o130(.A(i_12_), .B(ori_ori_n152_), .Y(ori_ori_n153_));
  NO2        o131(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n154_));
  OR2        o132(.A(i_8_), .B(i_7_), .Y(ori_ori_n155_));
  INV        o133(.A(i_12_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n44_), .B(ori_ori_n156_), .Y(ori_ori_n157_));
  NA2        o135(.A(i_2_), .B(i_1_), .Y(ori_ori_n158_));
  NO3        o136(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n159_));
  NAi21      o137(.An(i_4_), .B(i_3_), .Y(ori_ori_n160_));
  NO2        o138(.A(i_0_), .B(i_6_), .Y(ori_ori_n161_));
  NOi41      o139(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n162_));
  NO2        o140(.A(i_11_), .B(ori_ori_n152_), .Y(ori_ori_n163_));
  NOi21      o141(.An(i_1_), .B(i_6_), .Y(ori_ori_n164_));
  NAi21      o142(.An(i_3_), .B(i_7_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n156_), .B(i_9_), .Y(ori_ori_n166_));
  OR4        o144(.A(ori_ori_n166_), .B(ori_ori_n165_), .C(ori_ori_n164_), .D(ori_ori_n141_), .Y(ori_ori_n167_));
  NA2        o145(.A(ori_ori_n66_), .B(i_5_), .Y(ori_ori_n168_));
  NA2        o146(.A(i_3_), .B(i_9_), .Y(ori_ori_n169_));
  NAi21      o147(.An(i_7_), .B(i_10_), .Y(ori_ori_n170_));
  NO2        o148(.A(ori_ori_n170_), .B(ori_ori_n169_), .Y(ori_ori_n171_));
  NA3        o149(.A(ori_ori_n171_), .B(ori_ori_n168_), .C(ori_ori_n57_), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n172_), .B(ori_ori_n167_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n173_), .B(ori_ori_n163_), .Y(ori_ori_n174_));
  NA2        o152(.A(i_12_), .B(i_6_), .Y(ori_ori_n175_));
  OR2        o153(.A(i_13_), .B(i_9_), .Y(ori_ori_n176_));
  NO2        o154(.A(ori_ori_n160_), .B(i_2_), .Y(ori_ori_n177_));
  NO2        o155(.A(ori_ori_n165_), .B(i_8_), .Y(ori_ori_n178_));
  NO3        o156(.A(i_12_), .B(ori_ori_n152_), .C(ori_ori_n37_), .Y(ori_ori_n179_));
  NO2        o157(.A(i_2_), .B(ori_ori_n92_), .Y(ori_ori_n180_));
  AN2        o158(.A(i_3_), .B(i_10_), .Y(ori_ori_n181_));
  NO2        o159(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n182_));
  NO2        o160(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n183_));
  NO2        o161(.A(i_2_), .B(i_3_), .Y(ori_ori_n184_));
  NO2        o162(.A(i_12_), .B(i_10_), .Y(ori_ori_n185_));
  NOi21      o163(.An(i_5_), .B(i_0_), .Y(ori_ori_n186_));
  NOi32      o164(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n187_));
  INV        o165(.A(ori_ori_n187_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n134_), .B(ori_ori_n132_), .Y(ori_ori_n189_));
  NOi32      o167(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n190_));
  NO2        o168(.A(i_1_), .B(ori_ori_n92_), .Y(ori_ori_n191_));
  NAi21      o169(.An(i_3_), .B(i_4_), .Y(ori_ori_n192_));
  NO2        o170(.A(ori_ori_n192_), .B(i_9_), .Y(ori_ori_n193_));
  AN2        o171(.A(i_6_), .B(i_7_), .Y(ori_ori_n194_));
  OAI210     o172(.A0(ori_ori_n194_), .A1(ori_ori_n191_), .B0(ori_ori_n193_), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n192_), .B(i_10_), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n195_), .B(ori_ori_n141_), .Y(ori_ori_n197_));
  AOI210     o175(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n198_));
  OAI210     o176(.A0(ori_ori_n198_), .A1(ori_ori_n142_), .B0(ori_ori_n196_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n199_), .B(i_5_), .Y(ori_ori_n200_));
  NO3        o178(.A(ori_ori_n200_), .B(ori_ori_n197_), .C(ori_ori_n189_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n201_), .B(ori_ori_n188_), .Y(ori_ori_n202_));
  AN2        o180(.A(i_12_), .B(i_5_), .Y(ori_ori_n203_));
  NO2        o181(.A(i_11_), .B(i_6_), .Y(ori_ori_n204_));
  NO2        o182(.A(i_5_), .B(i_10_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n206_));
  NO3        o184(.A(ori_ori_n77_), .B(ori_ori_n47_), .C(i_9_), .Y(ori_ori_n207_));
  NO2        o185(.A(i_0_), .B(i_11_), .Y(ori_ori_n208_));
  NOi21      o186(.An(i_2_), .B(i_12_), .Y(ori_ori_n209_));
  NAi21      o187(.An(i_9_), .B(i_4_), .Y(ori_ori_n210_));
  OR2        o188(.A(i_13_), .B(i_10_), .Y(ori_ori_n211_));
  NO3        o189(.A(ori_ori_n211_), .B(ori_ori_n106_), .C(ori_ori_n210_), .Y(ori_ori_n212_));
  NO2        o190(.A(ori_ori_n92_), .B(ori_ori_n25_), .Y(ori_ori_n213_));
  INV        o191(.A(ori_ori_n202_), .Y(ori_ori_n214_));
  NO2        o192(.A(ori_ori_n66_), .B(i_13_), .Y(ori_ori_n215_));
  NO2        o193(.A(i_10_), .B(i_9_), .Y(ori_ori_n216_));
  NAi21      o194(.An(i_12_), .B(i_8_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n217_), .B(i_3_), .Y(ori_ori_n218_));
  NO3        o196(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n175_), .B(ori_ori_n88_), .Y(ori_ori_n220_));
  NA2        o198(.A(ori_ori_n220_), .B(ori_ori_n219_), .Y(ori_ori_n221_));
  NA2        o199(.A(i_8_), .B(i_9_), .Y(ori_ori_n222_));
  NO2        o200(.A(i_7_), .B(i_2_), .Y(ori_ori_n223_));
  OR2        o201(.A(ori_ori_n223_), .B(ori_ori_n222_), .Y(ori_ori_n224_));
  NA2        o202(.A(ori_ori_n179_), .B(ori_ori_n147_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n225_), .B(ori_ori_n224_), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n163_), .B(ori_ori_n182_), .Y(ori_ori_n227_));
  NO3        o205(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n228_));
  INV        o206(.A(ori_ori_n228_), .Y(ori_ori_n229_));
  NO2        o207(.A(ori_ori_n229_), .B(ori_ori_n227_), .Y(ori_ori_n230_));
  NO2        o208(.A(ori_ori_n230_), .B(ori_ori_n226_), .Y(ori_ori_n231_));
  NO2        o209(.A(i_11_), .B(i_1_), .Y(ori_ori_n232_));
  NOi21      o210(.An(i_2_), .B(i_7_), .Y(ori_ori_n233_));
  NA3        o211(.A(ori_ori_n162_), .B(ori_ori_n138_), .C(ori_ori_n120_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n132_), .B(i_3_), .Y(ori_ori_n236_));
  NAi31      o214(.An(ori_ori_n235_), .B(ori_ori_n236_), .C(ori_ori_n153_), .Y(ori_ori_n237_));
  NA3        o215(.A(ori_ori_n206_), .B(ori_ori_n140_), .C(ori_ori_n130_), .Y(ori_ori_n238_));
  NA3        o216(.A(ori_ori_n238_), .B(ori_ori_n237_), .C(ori_ori_n234_), .Y(ori_ori_n239_));
  INV        o217(.A(ori_ori_n239_), .Y(ori_ori_n240_));
  NA2        o218(.A(ori_ori_n219_), .B(ori_ori_n203_), .Y(ori_ori_n241_));
  NA2        o219(.A(ori_ori_n228_), .B(ori_ori_n205_), .Y(ori_ori_n242_));
  NA2        o220(.A(ori_ori_n240_), .B(ori_ori_n231_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n203_), .B(ori_ori_n152_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n194_), .B(ori_ori_n190_), .Y(ori_ori_n245_));
  OR2        o223(.A(ori_ori_n244_), .B(ori_ori_n245_), .Y(ori_ori_n246_));
  NO2        o224(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n247_));
  AOI210     o225(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n212_), .Y(ori_ori_n248_));
  NA2        o226(.A(ori_ori_n248_), .B(ori_ori_n246_), .Y(ori_ori_n249_));
  NA3        o227(.A(ori_ori_n151_), .B(ori_ori_n64_), .C(ori_ori_n44_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n179_), .B(ori_ori_n75_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n250_), .B(ori_ori_n251_), .Y(ori_ori_n252_));
  NO3        o230(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n211_), .B(i_1_), .Y(ori_ori_n254_));
  NOi31      o232(.An(ori_ori_n254_), .B(ori_ori_n220_), .C(ori_ori_n66_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n77_), .B(ori_ori_n25_), .Y(ori_ori_n256_));
  NO2        o234(.A(ori_ori_n105_), .B(ori_ori_n23_), .Y(ori_ori_n257_));
  NO2        o235(.A(i_12_), .B(ori_ori_n77_), .Y(ori_ori_n258_));
  NO3        o236(.A(ori_ori_n252_), .B(ori_ori_n249_), .C(ori_ori_n243_), .Y(ori_ori_n259_));
  NA3        o237(.A(ori_ori_n259_), .B(ori_ori_n214_), .C(ori_ori_n174_), .Y(ori7));
  NO2        o238(.A(ori_ori_n84_), .B(ori_ori_n52_), .Y(ori_ori_n261_));
  NA2        o239(.A(i_11_), .B(ori_ori_n144_), .Y(ori_ori_n262_));
  NA3        o240(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n156_), .B(i_4_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n264_), .B(i_8_), .Y(ori_ori_n265_));
  NO2        o243(.A(ori_ori_n96_), .B(ori_ori_n263_), .Y(ori_ori_n266_));
  NA2        o244(.A(i_2_), .B(ori_ori_n77_), .Y(ori_ori_n267_));
  OAI210     o245(.A0(ori_ori_n78_), .A1(ori_ori_n145_), .B0(ori_ori_n146_), .Y(ori_ori_n268_));
  NO2        o246(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n269_));
  NA2        o247(.A(i_4_), .B(i_8_), .Y(ori_ori_n270_));
  AOI210     o248(.A0(ori_ori_n270_), .A1(ori_ori_n181_), .B0(ori_ori_n269_), .Y(ori_ori_n271_));
  OAI220     o249(.A0(ori_ori_n271_), .A1(ori_ori_n267_), .B0(ori_ori_n268_), .B1(i_13_), .Y(ori_ori_n272_));
  NO3        o250(.A(ori_ori_n272_), .B(ori_ori_n266_), .C(ori_ori_n261_), .Y(ori_ori_n273_));
  AOI210     o251(.A0(ori_ori_n116_), .A1(ori_ori_n55_), .B0(i_10_), .Y(ori_ori_n274_));
  AOI210     o252(.A0(ori_ori_n274_), .A1(ori_ori_n156_), .B0(ori_ori_n136_), .Y(ori_ori_n275_));
  OR2        o253(.A(i_6_), .B(i_10_), .Y(ori_ori_n276_));
  OR3        o254(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n277_));
  OR2        o255(.A(ori_ori_n275_), .B(ori_ori_n176_), .Y(ori_ori_n278_));
  AOI210     o256(.A0(ori_ori_n278_), .A1(ori_ori_n273_), .B0(ori_ori_n56_), .Y(ori_ori_n279_));
  NOi21      o257(.An(i_11_), .B(i_7_), .Y(ori_ori_n280_));
  AO210      o258(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n281_), .B(ori_ori_n280_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n282_), .B(ori_ori_n148_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n283_), .B(ori_ori_n56_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n153_), .B(ori_ori_n56_), .Y(ori_ori_n285_));
  NO2        o263(.A(i_1_), .B(i_12_), .Y(ori_ori_n286_));
  INV        o264(.A(ori_ori_n285_), .Y(ori_ori_n287_));
  OAI210     o265(.A0(ori_ori_n287_), .A1(ori_ori_n284_), .B0(i_6_), .Y(ori_ori_n288_));
  NO2        o266(.A(i_6_), .B(i_11_), .Y(ori_ori_n289_));
  INV        o267(.A(ori_ori_n221_), .Y(ori_ori_n290_));
  NO3        o268(.A(ori_ori_n276_), .B(ori_ori_n155_), .C(ori_ori_n23_), .Y(ori_ori_n291_));
  AOI210     o269(.A0(i_1_), .A1(ori_ori_n171_), .B0(ori_ori_n291_), .Y(ori_ori_n292_));
  NO2        o270(.A(ori_ori_n292_), .B(ori_ori_n44_), .Y(ori_ori_n293_));
  INV        o271(.A(i_2_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n125_), .B(i_9_), .Y(ori_ori_n295_));
  NO2        o273(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n296_));
  NO2        o274(.A(ori_ori_n295_), .B(ori_ori_n294_), .Y(ori_ori_n297_));
  AOI210     o275(.A0(ori_ori_n232_), .A1(ori_ori_n213_), .B0(ori_ori_n159_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n298_), .B(ori_ori_n267_), .Y(ori_ori_n299_));
  NO2        o277(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n300_));
  OR2        o278(.A(ori_ori_n299_), .B(ori_ori_n297_), .Y(ori_ori_n301_));
  NO3        o279(.A(ori_ori_n301_), .B(ori_ori_n293_), .C(ori_ori_n290_), .Y(ori_ori_n302_));
  NO2        o280(.A(ori_ori_n156_), .B(ori_ori_n92_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n303_), .B(ori_ori_n280_), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n304_), .B(i_1_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n305_), .B(ori_ori_n277_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n210_), .B(ori_ori_n77_), .Y(ori_ori_n307_));
  NA2        o285(.A(ori_ori_n306_), .B(ori_ori_n46_), .Y(ori_ori_n308_));
  NO2        o286(.A(ori_ori_n155_), .B(ori_ori_n44_), .Y(ori_ori_n309_));
  NO3        o287(.A(ori_ori_n309_), .B(ori_ori_n183_), .C(ori_ori_n157_), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n106_), .B(ori_ori_n37_), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n311_), .B(i_6_), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n77_), .B(i_9_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n313_), .B(ori_ori_n56_), .Y(ori_ori_n314_));
  NO2        o292(.A(ori_ori_n314_), .B(ori_ori_n286_), .Y(ori_ori_n315_));
  NO4        o293(.A(ori_ori_n315_), .B(ori_ori_n312_), .C(ori_ori_n310_), .D(i_4_), .Y(ori_ori_n316_));
  INV        o294(.A(ori_ori_n316_), .Y(ori_ori_n317_));
  NA4        o295(.A(ori_ori_n317_), .B(ori_ori_n308_), .C(ori_ori_n302_), .D(ori_ori_n288_), .Y(ori_ori_n318_));
  AOI210     o296(.A0(ori_ori_n175_), .A1(ori_ori_n88_), .B0(i_1_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n192_), .B(i_2_), .Y(ori_ori_n320_));
  NA2        o298(.A(ori_ori_n320_), .B(ori_ori_n319_), .Y(ori_ori_n321_));
  NO2        o299(.A(ori_ori_n321_), .B(i_13_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n52_), .B(i_12_), .Y(ori_ori_n323_));
  INV        o301(.A(ori_ori_n323_), .Y(ori_ori_n324_));
  NO2        o302(.A(ori_ori_n233_), .B(ori_ori_n24_), .Y(ori_ori_n325_));
  NA2        o303(.A(ori_ori_n325_), .B(ori_ori_n307_), .Y(ori_ori_n326_));
  OAI220     o304(.A0(ori_ori_n326_), .A1(ori_ori_n41_), .B0(ori_ori_n324_), .B1(ori_ori_n84_), .Y(ori_ori_n327_));
  INV        o305(.A(ori_ori_n327_), .Y(ori_ori_n328_));
  NA2        o306(.A(ori_ori_n204_), .B(ori_ori_n296_), .Y(ori_ori_n329_));
  NO2        o307(.A(ori_ori_n329_), .B(ori_ori_n160_), .Y(ori_ori_n330_));
  NA2        o308(.A(ori_ori_n115_), .B(i_13_), .Y(ori_ori_n331_));
  NO2        o309(.A(ori_ori_n331_), .B(ori_ori_n319_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n26_), .B(ori_ori_n144_), .Y(ori_ori_n333_));
  NA2        o311(.A(ori_ori_n83_), .B(ori_ori_n93_), .Y(ori_ori_n334_));
  NO2        o312(.A(ori_ori_n334_), .B(ori_ori_n265_), .Y(ori_ori_n335_));
  NO3        o313(.A(ori_ori_n335_), .B(ori_ori_n332_), .C(ori_ori_n330_), .Y(ori_ori_n336_));
  OR2        o314(.A(i_11_), .B(i_6_), .Y(ori_ori_n337_));
  NA3        o315(.A(ori_ori_n264_), .B(ori_ori_n333_), .C(i_7_), .Y(ori_ori_n338_));
  NO2        o316(.A(ori_ori_n338_), .B(ori_ori_n337_), .Y(ori_ori_n339_));
  NA3        o317(.A(ori_ori_n209_), .B(ori_ori_n269_), .C(ori_ori_n88_), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n289_), .B(i_13_), .Y(ori_ori_n341_));
  NAi21      o319(.An(i_11_), .B(i_12_), .Y(ori_ori_n342_));
  NOi41      o320(.An(ori_ori_n101_), .B(ori_ori_n342_), .C(i_13_), .D(ori_ori_n77_), .Y(ori_ori_n343_));
  INV        o321(.A(ori_ori_n343_), .Y(ori_ori_n344_));
  NA3        o322(.A(ori_ori_n344_), .B(ori_ori_n341_), .C(ori_ori_n340_), .Y(ori_ori_n345_));
  OAI210     o323(.A0(ori_ori_n345_), .A1(ori_ori_n339_), .B0(ori_ori_n56_), .Y(ori_ori_n346_));
  NO2        o324(.A(i_2_), .B(i_12_), .Y(ori_ori_n347_));
  NA2        o325(.A(ori_ori_n191_), .B(ori_ori_n347_), .Y(ori_ori_n348_));
  INV        o326(.A(ori_ori_n348_), .Y(ori_ori_n349_));
  NA3        o327(.A(ori_ori_n349_), .B(ori_ori_n45_), .C(ori_ori_n152_), .Y(ori_ori_n350_));
  NA4        o328(.A(ori_ori_n350_), .B(ori_ori_n346_), .C(ori_ori_n336_), .D(ori_ori_n328_), .Y(ori_ori_n351_));
  OR4        o329(.A(ori_ori_n351_), .B(ori_ori_n322_), .C(ori_ori_n318_), .D(ori_ori_n279_), .Y(ori5));
  NA2        o330(.A(ori_ori_n304_), .B(ori_ori_n177_), .Y(ori_ori_n353_));
  AN2        o331(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n354_));
  NA3        o332(.A(ori_ori_n354_), .B(ori_ori_n347_), .C(ori_ori_n99_), .Y(ori_ori_n355_));
  NO2        o333(.A(ori_ori_n265_), .B(i_11_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n78_), .B(ori_ori_n356_), .Y(ori_ori_n357_));
  NA3        o335(.A(ori_ori_n357_), .B(ori_ori_n355_), .C(ori_ori_n353_), .Y(ori_ori_n358_));
  NO3        o336(.A(i_11_), .B(ori_ori_n156_), .C(i_13_), .Y(ori_ori_n359_));
  NO2        o337(.A(ori_ori_n112_), .B(ori_ori_n23_), .Y(ori_ori_n360_));
  NA2        o338(.A(i_12_), .B(i_8_), .Y(ori_ori_n361_));
  OAI210     o339(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n361_), .Y(ori_ori_n362_));
  INV        o340(.A(ori_ori_n216_), .Y(ori_ori_n363_));
  AOI220     o341(.A0(ori_ori_n184_), .A1(ori_ori_n257_), .B0(ori_ori_n362_), .B1(ori_ori_n360_), .Y(ori_ori_n364_));
  INV        o342(.A(ori_ori_n364_), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n365_), .B(ori_ori_n358_), .Y(ori_ori_n366_));
  INV        o344(.A(ori_ori_n138_), .Y(ori_ori_n367_));
  INV        o345(.A(ori_ori_n162_), .Y(ori_ori_n368_));
  OAI210     o346(.A0(ori_ori_n320_), .A1(ori_ori_n218_), .B0(ori_ori_n101_), .Y(ori_ori_n369_));
  AOI210     o347(.A0(ori_ori_n369_), .A1(ori_ori_n368_), .B0(ori_ori_n367_), .Y(ori_ori_n370_));
  NO2        o348(.A(ori_ori_n222_), .B(ori_ori_n26_), .Y(ori_ori_n371_));
  NO2        o349(.A(ori_ori_n371_), .B(ori_ori_n213_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n372_), .B(i_2_), .Y(ori_ori_n373_));
  INV        o351(.A(ori_ori_n373_), .Y(ori_ori_n374_));
  AOI210     o352(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n211_), .Y(ori_ori_n375_));
  AOI210     o353(.A0(ori_ori_n375_), .A1(ori_ori_n374_), .B0(ori_ori_n370_), .Y(ori_ori_n376_));
  NO2        o354(.A(ori_ori_n143_), .B(ori_ori_n113_), .Y(ori_ori_n377_));
  OAI210     o355(.A0(ori_ori_n377_), .A1(ori_ori_n360_), .B0(i_2_), .Y(ori_ori_n378_));
  INV        o356(.A(ori_ori_n139_), .Y(ori_ori_n379_));
  NO3        o357(.A(ori_ori_n281_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n380_));
  AOI210     o358(.A0(ori_ori_n379_), .A1(ori_ori_n78_), .B0(ori_ori_n380_), .Y(ori_ori_n381_));
  AOI210     o359(.A0(ori_ori_n381_), .A1(ori_ori_n378_), .B0(ori_ori_n144_), .Y(ori_ori_n382_));
  OA210      o360(.A0(ori_ori_n282_), .A1(ori_ori_n114_), .B0(i_13_), .Y(ori_ori_n383_));
  AOI210     o361(.A0(ori_ori_n149_), .A1(ori_ori_n129_), .B0(ori_ori_n247_), .Y(ori_ori_n384_));
  NA2        o362(.A(ori_ori_n384_), .B(ori_ori_n213_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n93_), .B(ori_ori_n44_), .Y(ori_ori_n386_));
  INV        o364(.A(ori_ori_n180_), .Y(ori_ori_n387_));
  NA4        o365(.A(ori_ori_n387_), .B(ori_ori_n181_), .C(ori_ori_n112_), .D(ori_ori_n42_), .Y(ori_ori_n388_));
  OAI210     o366(.A0(ori_ori_n388_), .A1(ori_ori_n386_), .B0(ori_ori_n385_), .Y(ori_ori_n389_));
  NO3        o367(.A(ori_ori_n389_), .B(ori_ori_n383_), .C(ori_ori_n382_), .Y(ori_ori_n390_));
  NA2        o368(.A(ori_ori_n257_), .B(ori_ori_n28_), .Y(ori_ori_n391_));
  NA2        o369(.A(ori_ori_n359_), .B(ori_ori_n178_), .Y(ori_ori_n392_));
  NA2        o370(.A(ori_ori_n392_), .B(ori_ori_n391_), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n55_), .B(i_12_), .Y(ori_ori_n394_));
  NO2        o372(.A(ori_ori_n394_), .B(ori_ori_n114_), .Y(ori_ori_n395_));
  NO2        o373(.A(ori_ori_n395_), .B(ori_ori_n262_), .Y(ori_ori_n396_));
  AOI220     o374(.A0(ori_ori_n396_), .A1(ori_ori_n36_), .B0(ori_ori_n393_), .B1(ori_ori_n46_), .Y(ori_ori_n397_));
  NA4        o375(.A(ori_ori_n397_), .B(ori_ori_n390_), .C(ori_ori_n376_), .D(ori_ori_n366_), .Y(ori6));
  OR2        o376(.A(ori_ori_n506_), .B(i_12_), .Y(ori_ori_n399_));
  NA2        o377(.A(ori_ori_n258_), .B(ori_ori_n56_), .Y(ori_ori_n400_));
  INV        o378(.A(ori_ori_n400_), .Y(ori_ori_n401_));
  NA2        o379(.A(ori_ori_n401_), .B(ori_ori_n66_), .Y(ori_ori_n402_));
  INV        o380(.A(ori_ori_n185_), .Y(ori_ori_n403_));
  NA2        o381(.A(ori_ori_n68_), .B(ori_ori_n119_), .Y(ori_ori_n404_));
  INV        o382(.A(ori_ori_n112_), .Y(ori_ori_n405_));
  NA2        o383(.A(ori_ori_n405_), .B(ori_ori_n46_), .Y(ori_ori_n406_));
  AOI210     o384(.A0(ori_ori_n406_), .A1(ori_ori_n404_), .B0(ori_ori_n403_), .Y(ori_ori_n407_));
  NO2        o385(.A(ori_ori_n164_), .B(i_9_), .Y(ori_ori_n408_));
  NA2        o386(.A(ori_ori_n408_), .B(ori_ori_n394_), .Y(ori_ori_n409_));
  AOI210     o387(.A0(ori_ori_n409_), .A1(ori_ori_n245_), .B0(ori_ori_n141_), .Y(ori_ori_n410_));
  NAi32      o388(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n411_));
  NO2        o389(.A(ori_ori_n337_), .B(ori_ori_n411_), .Y(ori_ori_n412_));
  OR3        o390(.A(ori_ori_n412_), .B(ori_ori_n410_), .C(ori_ori_n407_), .Y(ori_ori_n413_));
  BUFFER     o391(.A(ori_ori_n282_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n414_), .B(ori_ori_n128_), .Y(ori_ori_n415_));
  AO210      o393(.A0(ori_ori_n242_), .A1(ori_ori_n363_), .B0(ori_ori_n36_), .Y(ori_ori_n416_));
  NA2        o394(.A(ori_ori_n416_), .B(ori_ori_n415_), .Y(ori_ori_n417_));
  NO2        o395(.A(i_6_), .B(i_11_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n418_), .B(ori_ori_n253_), .Y(ori_ori_n419_));
  NA2        o397(.A(ori_ori_n207_), .B(ori_ori_n63_), .Y(ori_ori_n420_));
  NA3        o398(.A(ori_ori_n420_), .B(ori_ori_n419_), .C(ori_ori_n268_), .Y(ori_ori_n421_));
  NA2        o399(.A(ori_ori_n218_), .B(ori_ori_n216_), .Y(ori_ori_n422_));
  NA2        o400(.A(ori_ori_n102_), .B(ori_ori_n208_), .Y(ori_ori_n423_));
  NA2        o401(.A(ori_ori_n423_), .B(ori_ori_n422_), .Y(ori_ori_n424_));
  NO4        o402(.A(ori_ori_n424_), .B(ori_ori_n421_), .C(ori_ori_n417_), .D(ori_ori_n413_), .Y(ori_ori_n425_));
  NA4        o403(.A(ori_ori_n425_), .B(ori_ori_n402_), .C(ori_ori_n399_), .D(ori_ori_n201_), .Y(ori3));
  NA2        o404(.A(i_12_), .B(i_10_), .Y(ori_ori_n427_));
  NO2        o405(.A(i_11_), .B(ori_ori_n156_), .Y(ori_ori_n428_));
  NA2        o406(.A(ori_ori_n268_), .B(ori_ori_n195_), .Y(ori_ori_n429_));
  NA2        o407(.A(ori_ori_n429_), .B(ori_ori_n40_), .Y(ori_ori_n430_));
  NOi21      o408(.An(ori_ori_n87_), .B(ori_ori_n372_), .Y(ori_ori_n431_));
  INV        o409(.A(ori_ori_n431_), .Y(ori_ori_n432_));
  AOI210     o410(.A0(ori_ori_n432_), .A1(ori_ori_n430_), .B0(ori_ori_n47_), .Y(ori_ori_n433_));
  NO4        o411(.A(ori_ori_n198_), .B(ori_ori_n203_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n434_));
  NA2        o412(.A(ori_ori_n141_), .B(i_10_), .Y(ori_ori_n435_));
  NOi21      o413(.An(ori_ori_n435_), .B(ori_ori_n434_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n436_), .B(ori_ori_n56_), .Y(ori_ori_n437_));
  NOi21      o415(.An(i_5_), .B(i_9_), .Y(ori_ori_n438_));
  NA2        o416(.A(ori_ori_n438_), .B(ori_ori_n215_), .Y(ori_ori_n439_));
  BUFFER     o417(.A(ori_ori_n175_), .Y(ori_ori_n440_));
  NA2        o418(.A(ori_ori_n440_), .B(ori_ori_n232_), .Y(ori_ori_n441_));
  NO2        o419(.A(ori_ori_n441_), .B(ori_ori_n439_), .Y(ori_ori_n442_));
  NO3        o420(.A(ori_ori_n442_), .B(ori_ori_n437_), .C(ori_ori_n433_), .Y(ori_ori_n443_));
  NA2        o421(.A(ori_ori_n256_), .B(i_0_), .Y(ori_ori_n444_));
  NA2        o422(.A(ori_ori_n359_), .B(ori_ori_n186_), .Y(ori_ori_n445_));
  INV        o423(.A(ori_ori_n54_), .Y(ori_ori_n446_));
  NO2        o424(.A(ori_ori_n446_), .B(ori_ori_n445_), .Y(ori_ori_n447_));
  NO2        o425(.A(ori_ori_n166_), .B(ori_ori_n131_), .Y(ori_ori_n448_));
  NA2        o426(.A(i_0_), .B(i_10_), .Y(ori_ori_n449_));
  AN2        o427(.A(ori_ori_n448_), .B(i_6_), .Y(ori_ori_n450_));
  NO2        o428(.A(ori_ori_n450_), .B(ori_ori_n447_), .Y(ori_ori_n451_));
  INV        o429(.A(ori_ori_n451_), .Y(ori_ori_n452_));
  NA2        o430(.A(i_11_), .B(i_9_), .Y(ori_ori_n453_));
  NO3        o431(.A(i_12_), .B(ori_ori_n453_), .C(ori_ori_n267_), .Y(ori_ori_n454_));
  AN2        o432(.A(ori_ori_n454_), .B(i_5_), .Y(ori_ori_n455_));
  NA2        o433(.A(ori_ori_n206_), .B(ori_ori_n140_), .Y(ori_ori_n456_));
  NA2        o434(.A(ori_ori_n456_), .B(ori_ori_n135_), .Y(ori_ori_n457_));
  NO2        o435(.A(ori_ori_n453_), .B(ori_ori_n66_), .Y(ori_ori_n458_));
  NO2        o436(.A(ori_ori_n457_), .B(ori_ori_n455_), .Y(ori_ori_n459_));
  NA2        o437(.A(ori_ori_n300_), .B(ori_ori_n109_), .Y(ori_ori_n460_));
  NO2        o438(.A(i_6_), .B(ori_ori_n460_), .Y(ori_ori_n461_));
  NA2        o439(.A(ori_ori_n138_), .B(ori_ori_n94_), .Y(ori_ori_n462_));
  INV        o440(.A(ori_ori_n461_), .Y(ori_ori_n463_));
  NA2        o441(.A(ori_ori_n463_), .B(ori_ori_n459_), .Y(ori_ori_n464_));
  NO2        o442(.A(ori_ori_n427_), .B(ori_ori_n184_), .Y(ori_ori_n465_));
  NA2        o443(.A(ori_ori_n465_), .B(ori_ori_n458_), .Y(ori_ori_n466_));
  NA2        o444(.A(ori_ori_n246_), .B(ori_ori_n466_), .Y(ori_ori_n467_));
  NO3        o445(.A(ori_ori_n467_), .B(ori_ori_n464_), .C(ori_ori_n452_), .Y(ori_ori_n468_));
  NO2        o446(.A(ori_ori_n400_), .B(ori_ori_n462_), .Y(ori_ori_n469_));
  INV        o447(.A(ori_ori_n469_), .Y(ori_ori_n470_));
  NA2        o448(.A(ori_ori_n161_), .B(ori_ori_n154_), .Y(ori_ori_n471_));
  AOI210     o449(.A0(ori_ori_n471_), .A1(ori_ori_n444_), .B0(ori_ori_n131_), .Y(ori_ori_n472_));
  INV        o450(.A(ori_ori_n472_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n473_), .B(ori_ori_n470_), .Y(ori_ori_n474_));
  NO3        o452(.A(ori_ori_n449_), .B(ori_ori_n438_), .C(ori_ori_n143_), .Y(ori_ori_n475_));
  AOI220     o453(.A0(ori_ori_n475_), .A1(i_11_), .B0(ori_ori_n255_), .B1(ori_ori_n68_), .Y(ori_ori_n476_));
  NO3        o454(.A(ori_ori_n150_), .B(ori_ori_n203_), .C(i_0_), .Y(ori_ori_n477_));
  OAI210     o455(.A0(ori_ori_n477_), .A1(ori_ori_n69_), .B0(i_13_), .Y(ori_ori_n478_));
  NA2        o456(.A(ori_ori_n478_), .B(ori_ori_n476_), .Y(ori_ori_n479_));
  NA2        o457(.A(ori_ori_n241_), .B(ori_ori_n234_), .Y(ori_ori_n480_));
  INV        o458(.A(ori_ori_n480_), .Y(ori_ori_n481_));
  NA3        o459(.A(ori_ori_n205_), .B(ori_ori_n138_), .C(ori_ori_n137_), .Y(ori_ori_n482_));
  INV        o460(.A(ori_ori_n482_), .Y(ori_ori_n483_));
  NO3        o461(.A(ori_ori_n453_), .B(ori_ori_n151_), .C(ori_ori_n143_), .Y(ori_ori_n484_));
  NO2        o462(.A(ori_ori_n484_), .B(ori_ori_n483_), .Y(ori_ori_n485_));
  NA2        o463(.A(ori_ori_n485_), .B(ori_ori_n481_), .Y(ori_ori_n486_));
  NO2        o464(.A(ori_ori_n77_), .B(i_5_), .Y(ori_ori_n487_));
  NA3        o465(.A(ori_ori_n428_), .B(ori_ori_n100_), .C(ori_ori_n112_), .Y(ori_ori_n488_));
  INV        o466(.A(ori_ori_n488_), .Y(ori_ori_n489_));
  NA2        o467(.A(ori_ori_n489_), .B(ori_ori_n487_), .Y(ori_ori_n490_));
  NAi21      o468(.An(ori_ori_n159_), .B(ori_ori_n160_), .Y(ori_ori_n491_));
  NO4        o469(.A(ori_ori_n158_), .B(ori_ori_n150_), .C(i_0_), .D(i_12_), .Y(ori_ori_n492_));
  NA2        o470(.A(ori_ori_n492_), .B(ori_ori_n491_), .Y(ori_ori_n493_));
  NA2        o471(.A(ori_ori_n493_), .B(ori_ori_n490_), .Y(ori_ori_n494_));
  NO4        o472(.A(ori_ori_n494_), .B(ori_ori_n486_), .C(ori_ori_n479_), .D(ori_ori_n474_), .Y(ori_ori_n495_));
  INV        o473(.A(ori_ori_n275_), .Y(ori_ori_n496_));
  NA2        o474(.A(ori_ori_n496_), .B(ori_ori_n148_), .Y(ori_ori_n497_));
  NO2        o475(.A(ori_ori_n497_), .B(ori_ori_n66_), .Y(ori_ori_n498_));
  INV        o476(.A(ori_ori_n200_), .Y(ori_ori_n499_));
  NO2        o477(.A(ori_ori_n499_), .B(ori_ori_n367_), .Y(ori_ori_n500_));
  NO2        o478(.A(ori_ori_n500_), .B(ori_ori_n498_), .Y(ori_ori_n501_));
  NA4        o479(.A(ori_ori_n501_), .B(ori_ori_n495_), .C(ori_ori_n468_), .D(ori_ori_n443_), .Y(ori4));
  INV        o480(.A(i_6_), .Y(ori_ori_n505_));
  INV        o481(.A(ori_ori_n186_), .Y(ori_ori_n506_));
  INV        o482(.A(ori_ori_n106_), .Y(ori_ori_n507_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m0019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m0021(.A(mai_mai_n35_), .Y(mai1));
  INV        m0022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m0023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m0024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m0025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m0026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m0027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m0028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  NO2        m0029(.A(mai_mai_n48_), .B(mai_mai_n47_), .Y(mai_mai_n52_));
  NA2        m0030(.A(i_0_), .B(i_2_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_7_), .B(i_9_), .Y(mai_mai_n54_));
  NO2        m0032(.A(mai_mai_n54_), .B(mai_mai_n53_), .Y(mai_mai_n55_));
  OAI210     m0033(.A0(mai_mai_n55_), .A1(mai_mai_n52_), .B0(mai_mai_n46_), .Y(mai_mai_n56_));
  NA3        m0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n57_));
  NO2        m0035(.A(i_1_), .B(i_6_), .Y(mai_mai_n58_));
  NA2        m0036(.A(i_8_), .B(i_7_), .Y(mai_mai_n59_));
  OAI210     m0037(.A0(mai_mai_n59_), .A1(mai_mai_n58_), .B0(mai_mai_n57_), .Y(mai_mai_n60_));
  NA2        m0038(.A(mai_mai_n60_), .B(i_12_), .Y(mai_mai_n61_));
  NAi21      m0039(.An(i_2_), .B(i_7_), .Y(mai_mai_n62_));
  INV        m0040(.A(i_1_), .Y(mai_mai_n63_));
  NA2        m0041(.A(mai_mai_n63_), .B(i_6_), .Y(mai_mai_n64_));
  NA3        m0042(.A(mai_mai_n64_), .B(mai_mai_n62_), .C(mai_mai_n31_), .Y(mai_mai_n65_));
  NA2        m0043(.A(mai_mai_n65_), .B(mai_mai_n61_), .Y(mai_mai_n66_));
  NA2        m0044(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n67_));
  AOI210     m0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n68_));
  NA2        m0046(.A(i_1_), .B(i_6_), .Y(mai_mai_n69_));
  NO2        m0047(.A(mai_mai_n69_), .B(mai_mai_n25_), .Y(mai_mai_n70_));
  INV        m0048(.A(i_0_), .Y(mai_mai_n71_));
  NAi21      m0049(.An(i_5_), .B(i_10_), .Y(mai_mai_n72_));
  NA2        m0050(.A(i_5_), .B(i_9_), .Y(mai_mai_n73_));
  AOI210     m0051(.A0(mai_mai_n73_), .A1(mai_mai_n72_), .B0(mai_mai_n71_), .Y(mai_mai_n74_));
  NO2        m0052(.A(mai_mai_n74_), .B(mai_mai_n70_), .Y(mai_mai_n75_));
  OAI210     m0053(.A0(mai_mai_n68_), .A1(mai_mai_n67_), .B0(mai_mai_n75_), .Y(mai_mai_n76_));
  OAI210     m0054(.A0(mai_mai_n76_), .A1(mai_mai_n66_), .B0(i_0_), .Y(mai_mai_n77_));
  NA2        m0055(.A(i_12_), .B(i_5_), .Y(mai_mai_n78_));
  NA2        m0056(.A(i_2_), .B(i_8_), .Y(mai_mai_n79_));
  NO2        m0057(.A(mai_mai_n79_), .B(mai_mai_n58_), .Y(mai_mai_n80_));
  NO2        m0058(.A(i_3_), .B(i_9_), .Y(mai_mai_n81_));
  NO2        m0059(.A(i_3_), .B(i_7_), .Y(mai_mai_n82_));
  INV        m0060(.A(i_6_), .Y(mai_mai_n83_));
  OR4        m0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n84_));
  INV        m0062(.A(mai_mai_n84_), .Y(mai_mai_n85_));
  NO2        m0063(.A(i_2_), .B(i_7_), .Y(mai_mai_n86_));
  NA2        m0064(.A(mai_mai_n80_), .B(i_2_), .Y(mai_mai_n87_));
  NAi21      m0065(.An(i_6_), .B(i_10_), .Y(mai_mai_n88_));
  NA2        m0066(.A(i_6_), .B(i_9_), .Y(mai_mai_n89_));
  AOI210     m0067(.A0(mai_mai_n89_), .A1(mai_mai_n88_), .B0(mai_mai_n63_), .Y(mai_mai_n90_));
  NA2        m0068(.A(i_2_), .B(i_6_), .Y(mai_mai_n91_));
  NO3        m0069(.A(mai_mai_n91_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n92_));
  NO2        m0070(.A(mai_mai_n92_), .B(mai_mai_n90_), .Y(mai_mai_n93_));
  AOI210     m0071(.A0(mai_mai_n93_), .A1(mai_mai_n87_), .B0(mai_mai_n78_), .Y(mai_mai_n94_));
  AN3        m0072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n95_));
  NAi21      m0073(.An(i_6_), .B(i_11_), .Y(mai_mai_n96_));
  NO2        m0074(.A(i_5_), .B(i_8_), .Y(mai_mai_n97_));
  NOi21      m0075(.An(mai_mai_n97_), .B(mai_mai_n96_), .Y(mai_mai_n98_));
  AOI220     m0076(.A0(mai_mai_n98_), .A1(mai_mai_n62_), .B0(mai_mai_n95_), .B1(mai_mai_n32_), .Y(mai_mai_n99_));
  INV        m0077(.A(i_7_), .Y(mai_mai_n100_));
  NA2        m0078(.A(mai_mai_n47_), .B(mai_mai_n100_), .Y(mai_mai_n101_));
  NO2        m0079(.A(i_0_), .B(i_5_), .Y(mai_mai_n102_));
  NO2        m0080(.A(mai_mai_n102_), .B(mai_mai_n83_), .Y(mai_mai_n103_));
  NA2        m0081(.A(i_12_), .B(i_3_), .Y(mai_mai_n104_));
  INV        m0082(.A(mai_mai_n104_), .Y(mai_mai_n105_));
  NA3        m0083(.A(mai_mai_n105_), .B(mai_mai_n103_), .C(mai_mai_n101_), .Y(mai_mai_n106_));
  NAi21      m0084(.An(i_7_), .B(i_11_), .Y(mai_mai_n107_));
  NO3        m0085(.A(mai_mai_n107_), .B(mai_mai_n88_), .C(mai_mai_n53_), .Y(mai_mai_n108_));
  AN2        m0086(.A(i_2_), .B(i_10_), .Y(mai_mai_n109_));
  NO2        m0087(.A(mai_mai_n109_), .B(i_7_), .Y(mai_mai_n110_));
  OR2        m0088(.A(mai_mai_n78_), .B(mai_mai_n58_), .Y(mai_mai_n111_));
  NO2        m0089(.A(i_8_), .B(mai_mai_n100_), .Y(mai_mai_n112_));
  NO3        m0090(.A(mai_mai_n112_), .B(mai_mai_n111_), .C(mai_mai_n110_), .Y(mai_mai_n113_));
  NA2        m0091(.A(i_12_), .B(i_7_), .Y(mai_mai_n114_));
  NO2        m0092(.A(mai_mai_n63_), .B(mai_mai_n26_), .Y(mai_mai_n115_));
  NA2        m0093(.A(mai_mai_n115_), .B(i_0_), .Y(mai_mai_n116_));
  NA2        m0094(.A(i_11_), .B(i_12_), .Y(mai_mai_n117_));
  OAI210     m0095(.A0(mai_mai_n116_), .A1(mai_mai_n114_), .B0(mai_mai_n117_), .Y(mai_mai_n118_));
  NO2        m0096(.A(mai_mai_n118_), .B(mai_mai_n113_), .Y(mai_mai_n119_));
  NAi41      m0097(.An(mai_mai_n108_), .B(mai_mai_n119_), .C(mai_mai_n106_), .D(mai_mai_n99_), .Y(mai_mai_n120_));
  NOi21      m0098(.An(i_1_), .B(i_5_), .Y(mai_mai_n121_));
  NA2        m0099(.A(mai_mai_n121_), .B(i_11_), .Y(mai_mai_n122_));
  NA2        m0100(.A(mai_mai_n100_), .B(mai_mai_n37_), .Y(mai_mai_n123_));
  NA2        m0101(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n124_));
  NA2        m0102(.A(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n125_));
  NO2        m0103(.A(mai_mai_n125_), .B(mai_mai_n47_), .Y(mai_mai_n126_));
  NA2        m0104(.A(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n127_));
  NAi21      m0105(.An(i_3_), .B(i_8_), .Y(mai_mai_n128_));
  NA2        m0106(.A(mai_mai_n128_), .B(mai_mai_n62_), .Y(mai_mai_n129_));
  NOi21      m0107(.An(mai_mai_n129_), .B(mai_mai_n127_), .Y(mai_mai_n130_));
  NO2        m0108(.A(i_1_), .B(mai_mai_n83_), .Y(mai_mai_n131_));
  NO2        m0109(.A(i_6_), .B(i_5_), .Y(mai_mai_n132_));
  NA2        m0110(.A(mai_mai_n132_), .B(i_3_), .Y(mai_mai_n133_));
  AO210      m0111(.A0(mai_mai_n133_), .A1(mai_mai_n48_), .B0(mai_mai_n131_), .Y(mai_mai_n134_));
  OAI220     m0112(.A0(mai_mai_n134_), .A1(mai_mai_n107_), .B0(mai_mai_n130_), .B1(mai_mai_n122_), .Y(mai_mai_n135_));
  NO3        m0113(.A(mai_mai_n135_), .B(mai_mai_n120_), .C(mai_mai_n94_), .Y(mai_mai_n136_));
  NA3        m0114(.A(mai_mai_n136_), .B(mai_mai_n77_), .C(mai_mai_n56_), .Y(mai2));
  NO2        m0115(.A(mai_mai_n63_), .B(mai_mai_n37_), .Y(mai_mai_n138_));
  NA2        m0116(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n139_));
  NA2        m0117(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n140_));
  NA4        m0118(.A(mai_mai_n140_), .B(mai_mai_n75_), .C(mai_mai_n67_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0119(.A(i_8_), .B(i_7_), .Y(mai_mai_n142_));
  NA2        m0120(.A(mai_mai_n142_), .B(i_6_), .Y(mai_mai_n143_));
  NO2        m0121(.A(i_12_), .B(i_13_), .Y(mai_mai_n144_));
  NAi21      m0122(.An(i_5_), .B(i_11_), .Y(mai_mai_n145_));
  NOi21      m0123(.An(mai_mai_n144_), .B(mai_mai_n145_), .Y(mai_mai_n146_));
  NO2        m0124(.A(i_0_), .B(i_1_), .Y(mai_mai_n147_));
  NA2        m0125(.A(i_2_), .B(i_3_), .Y(mai_mai_n148_));
  NO2        m0126(.A(mai_mai_n148_), .B(i_4_), .Y(mai_mai_n149_));
  NA3        m0127(.A(mai_mai_n149_), .B(mai_mai_n147_), .C(mai_mai_n146_), .Y(mai_mai_n150_));
  AN2        m0128(.A(mai_mai_n144_), .B(mai_mai_n81_), .Y(mai_mai_n151_));
  NA2        m0129(.A(i_1_), .B(i_5_), .Y(mai_mai_n152_));
  NO2        m0130(.A(mai_mai_n71_), .B(mai_mai_n47_), .Y(mai_mai_n153_));
  NA2        m0131(.A(mai_mai_n153_), .B(mai_mai_n36_), .Y(mai_mai_n154_));
  NO3        m0132(.A(mai_mai_n154_), .B(mai_mai_n152_), .C(i_13_), .Y(mai_mai_n155_));
  OR2        m0133(.A(i_0_), .B(i_1_), .Y(mai_mai_n156_));
  NO3        m0134(.A(mai_mai_n156_), .B(mai_mai_n78_), .C(i_13_), .Y(mai_mai_n157_));
  NAi32      m0135(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n158_));
  NAi21      m0136(.An(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NOi21      m0137(.An(i_4_), .B(i_10_), .Y(mai_mai_n160_));
  NA2        m0138(.A(mai_mai_n160_), .B(mai_mai_n40_), .Y(mai_mai_n161_));
  NO2        m0139(.A(i_3_), .B(i_5_), .Y(mai_mai_n162_));
  NO3        m0140(.A(mai_mai_n71_), .B(i_2_), .C(i_1_), .Y(mai_mai_n163_));
  NA2        m0141(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  OAI210     m0142(.A0(mai_mai_n164_), .A1(mai_mai_n161_), .B0(mai_mai_n159_), .Y(mai_mai_n165_));
  NO2        m0143(.A(mai_mai_n165_), .B(mai_mai_n155_), .Y(mai_mai_n166_));
  AOI210     m0144(.A0(mai_mai_n166_), .A1(mai_mai_n150_), .B0(mai_mai_n143_), .Y(mai_mai_n167_));
  NA3        m0145(.A(mai_mai_n71_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n168_));
  NOi21      m0146(.An(i_4_), .B(i_9_), .Y(mai_mai_n169_));
  NOi21      m0147(.An(i_11_), .B(i_13_), .Y(mai_mai_n170_));
  NA2        m0148(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n171_));
  BUFFER     m0149(.A(mai_mai_n171_), .Y(mai_mai_n172_));
  NO2        m0150(.A(i_4_), .B(i_5_), .Y(mai_mai_n173_));
  NAi21      m0151(.An(i_12_), .B(i_11_), .Y(mai_mai_n174_));
  NO2        m0152(.A(mai_mai_n174_), .B(i_13_), .Y(mai_mai_n175_));
  NA2        m0153(.A(mai_mai_n175_), .B(mai_mai_n173_), .Y(mai_mai_n176_));
  AOI210     m0154(.A0(mai_mai_n176_), .A1(mai_mai_n172_), .B0(mai_mai_n168_), .Y(mai_mai_n177_));
  NO2        m0155(.A(mai_mai_n71_), .B(mai_mai_n63_), .Y(mai_mai_n178_));
  NA2        m0156(.A(mai_mai_n178_), .B(mai_mai_n47_), .Y(mai_mai_n179_));
  NA2        m0157(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n180_));
  NAi31      m0158(.An(mai_mai_n180_), .B(mai_mai_n151_), .C(i_11_), .Y(mai_mai_n181_));
  NA2        m0159(.A(i_3_), .B(i_5_), .Y(mai_mai_n182_));
  AOI210     m0160(.A0(mai_mai_n171_), .A1(mai_mai_n181_), .B0(mai_mai_n179_), .Y(mai_mai_n183_));
  NO2        m0161(.A(mai_mai_n71_), .B(i_5_), .Y(mai_mai_n184_));
  NO2        m0162(.A(i_13_), .B(i_10_), .Y(mai_mai_n185_));
  NA3        m0163(.A(mai_mai_n185_), .B(mai_mai_n184_), .C(mai_mai_n45_), .Y(mai_mai_n186_));
  NO2        m0164(.A(i_2_), .B(i_1_), .Y(mai_mai_n187_));
  NA2        m0165(.A(mai_mai_n187_), .B(i_3_), .Y(mai_mai_n188_));
  NAi21      m0166(.An(i_4_), .B(i_12_), .Y(mai_mai_n189_));
  NO4        m0167(.A(mai_mai_n189_), .B(mai_mai_n188_), .C(mai_mai_n186_), .D(mai_mai_n25_), .Y(mai_mai_n190_));
  NO3        m0168(.A(mai_mai_n190_), .B(mai_mai_n183_), .C(mai_mai_n177_), .Y(mai_mai_n191_));
  INV        m0169(.A(i_8_), .Y(mai_mai_n192_));
  NA2        m0170(.A(i_8_), .B(i_6_), .Y(mai_mai_n193_));
  NO3        m0171(.A(i_3_), .B(mai_mai_n83_), .C(mai_mai_n49_), .Y(mai_mai_n194_));
  NA2        m0172(.A(mai_mai_n194_), .B(mai_mai_n112_), .Y(mai_mai_n195_));
  NO3        m0173(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n196_));
  NA3        m0174(.A(mai_mai_n196_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n197_));
  NO3        m0175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n198_));
  OAI210     m0176(.A0(mai_mai_n95_), .A1(i_12_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  AOI210     m0177(.A0(mai_mai_n199_), .A1(mai_mai_n197_), .B0(mai_mai_n195_), .Y(mai_mai_n200_));
  NO2        m0178(.A(i_3_), .B(i_8_), .Y(mai_mai_n201_));
  NO3        m0179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n202_));
  NA3        m0180(.A(mai_mai_n202_), .B(mai_mai_n201_), .C(mai_mai_n40_), .Y(mai_mai_n203_));
  NO2        m0181(.A(i_13_), .B(i_9_), .Y(mai_mai_n204_));
  NA3        m0182(.A(mai_mai_n204_), .B(i_6_), .C(mai_mai_n192_), .Y(mai_mai_n205_));
  NAi21      m0183(.An(i_12_), .B(i_3_), .Y(mai_mai_n206_));
  NO2        m0184(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n207_));
  NO3        m0185(.A(i_0_), .B(i_2_), .C(mai_mai_n63_), .Y(mai_mai_n208_));
  NA3        m0186(.A(mai_mai_n208_), .B(mai_mai_n207_), .C(i_10_), .Y(mai_mai_n209_));
  OAI220     m0187(.A0(mai_mai_n209_), .A1(mai_mai_n205_), .B0(mai_mai_n58_), .B1(mai_mai_n203_), .Y(mai_mai_n210_));
  AOI210     m0188(.A0(mai_mai_n210_), .A1(i_7_), .B0(mai_mai_n200_), .Y(mai_mai_n211_));
  OAI220     m0189(.A0(mai_mai_n211_), .A1(i_4_), .B0(mai_mai_n193_), .B1(mai_mai_n191_), .Y(mai_mai_n212_));
  NAi21      m0190(.An(i_12_), .B(i_7_), .Y(mai_mai_n213_));
  NA3        m0191(.A(i_13_), .B(mai_mai_n192_), .C(i_10_), .Y(mai_mai_n214_));
  NO2        m0192(.A(mai_mai_n214_), .B(mai_mai_n213_), .Y(mai_mai_n215_));
  NA2        m0193(.A(i_0_), .B(i_5_), .Y(mai_mai_n216_));
  OAI220     m0194(.A0(mai_mai_n83_), .A1(mai_mai_n188_), .B0(mai_mai_n179_), .B1(mai_mai_n133_), .Y(mai_mai_n217_));
  NAi31      m0195(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n218_));
  NO2        m0196(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n219_));
  NO2        m0197(.A(mai_mai_n47_), .B(mai_mai_n63_), .Y(mai_mai_n220_));
  NA3        m0198(.A(mai_mai_n220_), .B(i_0_), .C(mai_mai_n219_), .Y(mai_mai_n221_));
  INV        m0199(.A(i_13_), .Y(mai_mai_n222_));
  NO2        m0200(.A(i_12_), .B(mai_mai_n222_), .Y(mai_mai_n223_));
  NA3        m0201(.A(mai_mai_n223_), .B(mai_mai_n196_), .C(mai_mai_n194_), .Y(mai_mai_n224_));
  OAI210     m0202(.A0(mai_mai_n221_), .A1(mai_mai_n218_), .B0(mai_mai_n224_), .Y(mai_mai_n225_));
  AOI220     m0203(.A0(mai_mai_n225_), .A1(mai_mai_n142_), .B0(mai_mai_n217_), .B1(mai_mai_n215_), .Y(mai_mai_n226_));
  NO2        m0204(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n227_));
  NO2        m0205(.A(mai_mai_n182_), .B(i_4_), .Y(mai_mai_n228_));
  NA2        m0206(.A(mai_mai_n228_), .B(mai_mai_n227_), .Y(mai_mai_n229_));
  OR2        m0207(.A(i_8_), .B(i_7_), .Y(mai_mai_n230_));
  NO2        m0208(.A(mai_mai_n230_), .B(mai_mai_n83_), .Y(mai_mai_n231_));
  NO2        m0209(.A(mai_mai_n53_), .B(i_1_), .Y(mai_mai_n232_));
  INV        m0210(.A(i_12_), .Y(mai_mai_n233_));
  NO3        m0211(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n234_));
  NA2        m0212(.A(i_2_), .B(i_1_), .Y(mai_mai_n235_));
  NO2        m0213(.A(mai_mai_n230_), .B(mai_mai_n229_), .Y(mai_mai_n236_));
  NO3        m0214(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n237_));
  NAi21      m0215(.An(i_4_), .B(i_3_), .Y(mai_mai_n238_));
  NO2        m0216(.A(mai_mai_n238_), .B(mai_mai_n73_), .Y(mai_mai_n239_));
  NO2        m0217(.A(i_0_), .B(i_6_), .Y(mai_mai_n240_));
  NOi41      m0218(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n241_));
  NA2        m0219(.A(mai_mai_n241_), .B(mai_mai_n240_), .Y(mai_mai_n242_));
  NO2        m0220(.A(mai_mai_n235_), .B(mai_mai_n182_), .Y(mai_mai_n243_));
  NAi21      m0221(.An(mai_mai_n242_), .B(mai_mai_n243_), .Y(mai_mai_n244_));
  INV        m0222(.A(mai_mai_n244_), .Y(mai_mai_n245_));
  AOI220     m0223(.A0(mai_mai_n245_), .A1(mai_mai_n40_), .B0(mai_mai_n236_), .B1(mai_mai_n204_), .Y(mai_mai_n246_));
  NO2        m0224(.A(i_11_), .B(mai_mai_n222_), .Y(mai_mai_n247_));
  NOi21      m0225(.An(i_1_), .B(i_6_), .Y(mai_mai_n248_));
  NAi21      m0226(.An(i_3_), .B(i_7_), .Y(mai_mai_n249_));
  NO2        m0227(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n250_));
  NO2        m0228(.A(i_12_), .B(i_3_), .Y(mai_mai_n251_));
  NAi21      m0229(.An(i_7_), .B(i_10_), .Y(mai_mai_n252_));
  NA3        m0230(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n253_));
  INV        m0231(.A(mai_mai_n143_), .Y(mai_mai_n254_));
  NA2        m0232(.A(mai_mai_n233_), .B(i_13_), .Y(mai_mai_n255_));
  NO2        m0233(.A(mai_mai_n255_), .B(mai_mai_n73_), .Y(mai_mai_n256_));
  NA2        m0234(.A(mai_mai_n256_), .B(mai_mai_n254_), .Y(mai_mai_n257_));
  NO2        m0235(.A(mai_mai_n230_), .B(mai_mai_n37_), .Y(mai_mai_n258_));
  NA2        m0236(.A(i_12_), .B(i_6_), .Y(mai_mai_n259_));
  OR2        m0237(.A(i_13_), .B(i_9_), .Y(mai_mai_n260_));
  NO3        m0238(.A(mai_mai_n260_), .B(mai_mai_n259_), .C(mai_mai_n49_), .Y(mai_mai_n261_));
  NO2        m0239(.A(mai_mai_n238_), .B(i_2_), .Y(mai_mai_n262_));
  NA3        m0240(.A(mai_mai_n262_), .B(mai_mai_n261_), .C(mai_mai_n45_), .Y(mai_mai_n263_));
  NA2        m0241(.A(mai_mai_n247_), .B(i_9_), .Y(mai_mai_n264_));
  OAI210     m0242(.A0(mai_mai_n63_), .A1(mai_mai_n264_), .B0(mai_mai_n263_), .Y(mai_mai_n265_));
  NA2        m0243(.A(mai_mai_n153_), .B(mai_mai_n63_), .Y(mai_mai_n266_));
  NO3        m0244(.A(i_11_), .B(mai_mai_n222_), .C(mai_mai_n25_), .Y(mai_mai_n267_));
  NO2        m0245(.A(mai_mai_n249_), .B(i_8_), .Y(mai_mai_n268_));
  NO2        m0246(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n269_));
  NA3        m0247(.A(mai_mai_n269_), .B(mai_mai_n268_), .C(mai_mai_n267_), .Y(mai_mai_n270_));
  NO3        m0248(.A(mai_mai_n26_), .B(mai_mai_n83_), .C(i_5_), .Y(mai_mai_n271_));
  NA3        m0249(.A(mai_mai_n271_), .B(mai_mai_n258_), .C(mai_mai_n223_), .Y(mai_mai_n272_));
  AOI210     m0250(.A0(mai_mai_n272_), .A1(mai_mai_n270_), .B0(mai_mai_n266_), .Y(mai_mai_n273_));
  AOI210     m0251(.A0(mai_mai_n265_), .A1(mai_mai_n258_), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  NA4        m0252(.A(mai_mai_n274_), .B(mai_mai_n257_), .C(mai_mai_n246_), .D(mai_mai_n226_), .Y(mai_mai_n275_));
  NO3        m0253(.A(i_12_), .B(mai_mai_n222_), .C(mai_mai_n37_), .Y(mai_mai_n276_));
  INV        m0254(.A(mai_mai_n276_), .Y(mai_mai_n277_));
  NA2        m0255(.A(i_8_), .B(mai_mai_n100_), .Y(mai_mai_n278_));
  NO3        m0256(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n279_));
  AOI220     m0257(.A0(mai_mai_n279_), .A1(mai_mai_n194_), .B0(mai_mai_n162_), .B1(mai_mai_n232_), .Y(mai_mai_n280_));
  NO2        m0258(.A(mai_mai_n280_), .B(mai_mai_n278_), .Y(mai_mai_n281_));
  NO2        m0259(.A(mai_mai_n235_), .B(i_0_), .Y(mai_mai_n282_));
  AOI220     m0260(.A0(mai_mai_n282_), .A1(i_8_), .B0(i_1_), .B1(mai_mai_n142_), .Y(mai_mai_n283_));
  NA2        m0261(.A(mai_mai_n269_), .B(mai_mai_n26_), .Y(mai_mai_n284_));
  NO2        m0262(.A(mai_mai_n284_), .B(mai_mai_n283_), .Y(mai_mai_n285_));
  NA2        m0263(.A(i_0_), .B(i_1_), .Y(mai_mai_n286_));
  NO2        m0264(.A(mai_mai_n286_), .B(i_2_), .Y(mai_mai_n287_));
  NO2        m0265(.A(mai_mai_n59_), .B(i_6_), .Y(mai_mai_n288_));
  NA2        m0266(.A(mai_mai_n288_), .B(mai_mai_n287_), .Y(mai_mai_n289_));
  OAI210     m0267(.A0(mai_mai_n164_), .A1(mai_mai_n143_), .B0(mai_mai_n289_), .Y(mai_mai_n290_));
  NO3        m0268(.A(mai_mai_n290_), .B(mai_mai_n285_), .C(mai_mai_n281_), .Y(mai_mai_n291_));
  NO2        m0269(.A(i_3_), .B(i_10_), .Y(mai_mai_n292_));
  NA3        m0270(.A(mai_mai_n292_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n293_));
  NO2        m0271(.A(i_2_), .B(mai_mai_n100_), .Y(mai_mai_n294_));
  NA2        m0272(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n295_));
  NA3        m0273(.A(mai_mai_n216_), .B(i_1_), .C(mai_mai_n294_), .Y(mai_mai_n296_));
  AN2        m0274(.A(i_3_), .B(i_10_), .Y(mai_mai_n297_));
  NA4        m0275(.A(mai_mai_n297_), .B(mai_mai_n196_), .C(mai_mai_n175_), .D(mai_mai_n173_), .Y(mai_mai_n298_));
  NO2        m0276(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n299_));
  NO2        m0277(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n300_));
  OR2        m0278(.A(mai_mai_n296_), .B(mai_mai_n293_), .Y(mai_mai_n301_));
  OAI220     m0279(.A0(mai_mai_n301_), .A1(i_6_), .B0(mai_mai_n291_), .B1(mai_mai_n277_), .Y(mai_mai_n302_));
  NO4        m0280(.A(mai_mai_n302_), .B(mai_mai_n275_), .C(mai_mai_n212_), .D(mai_mai_n167_), .Y(mai_mai_n303_));
  NO3        m0281(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n304_));
  NO2        m0282(.A(mai_mai_n59_), .B(mai_mai_n83_), .Y(mai_mai_n305_));
  NA2        m0283(.A(mai_mai_n282_), .B(mai_mai_n305_), .Y(mai_mai_n306_));
  NO3        m0284(.A(i_6_), .B(mai_mai_n192_), .C(i_7_), .Y(mai_mai_n307_));
  NA2        m0285(.A(mai_mai_n307_), .B(mai_mai_n196_), .Y(mai_mai_n308_));
  AOI210     m0286(.A0(mai_mai_n308_), .A1(mai_mai_n306_), .B0(i_5_), .Y(mai_mai_n309_));
  NO2        m0287(.A(i_2_), .B(i_3_), .Y(mai_mai_n310_));
  OR2        m0288(.A(i_0_), .B(i_5_), .Y(mai_mai_n311_));
  NA2        m0289(.A(mai_mai_n216_), .B(mai_mai_n311_), .Y(mai_mai_n312_));
  NA4        m0290(.A(mai_mai_n312_), .B(mai_mai_n231_), .C(mai_mai_n310_), .D(i_1_), .Y(mai_mai_n313_));
  NA3        m0291(.A(mai_mai_n282_), .B(mai_mai_n162_), .C(mai_mai_n112_), .Y(mai_mai_n314_));
  NAi21      m0292(.An(i_8_), .B(i_7_), .Y(mai_mai_n315_));
  NO2        m0293(.A(mai_mai_n315_), .B(i_6_), .Y(mai_mai_n316_));
  NO2        m0294(.A(mai_mai_n156_), .B(mai_mai_n47_), .Y(mai_mai_n317_));
  NA2        m0295(.A(mai_mai_n317_), .B(mai_mai_n316_), .Y(mai_mai_n318_));
  NA3        m0296(.A(mai_mai_n318_), .B(mai_mai_n314_), .C(mai_mai_n313_), .Y(mai_mai_n319_));
  OAI210     m0297(.A0(mai_mai_n319_), .A1(mai_mai_n309_), .B0(i_4_), .Y(mai_mai_n320_));
  NO2        m0298(.A(i_12_), .B(i_10_), .Y(mai_mai_n321_));
  NOi21      m0299(.An(i_5_), .B(i_0_), .Y(mai_mai_n322_));
  NO3        m0300(.A(mai_mai_n295_), .B(mai_mai_n322_), .C(mai_mai_n128_), .Y(mai_mai_n323_));
  NA4        m0301(.A(mai_mai_n82_), .B(mai_mai_n36_), .C(mai_mai_n83_), .D(i_8_), .Y(mai_mai_n324_));
  NA2        m0302(.A(mai_mai_n323_), .B(mai_mai_n321_), .Y(mai_mai_n325_));
  NO2        m0303(.A(i_6_), .B(i_8_), .Y(mai_mai_n326_));
  AN2        m0304(.A(i_0_), .B(mai_mai_n326_), .Y(mai_mai_n327_));
  NO2        m0305(.A(i_1_), .B(i_7_), .Y(mai_mai_n328_));
  NA3        m0306(.A(mai_mai_n326_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n329_));
  NA3        m0307(.A(mai_mai_n329_), .B(mai_mai_n325_), .C(mai_mai_n320_), .Y(mai_mai_n330_));
  NO3        m0308(.A(mai_mai_n230_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n331_));
  NO3        m0309(.A(mai_mai_n315_), .B(i_2_), .C(i_1_), .Y(mai_mai_n332_));
  OAI210     m0310(.A0(mai_mai_n332_), .A1(mai_mai_n331_), .B0(i_6_), .Y(mai_mai_n333_));
  NA3        m0311(.A(mai_mai_n248_), .B(mai_mai_n294_), .C(mai_mai_n192_), .Y(mai_mai_n334_));
  AOI210     m0312(.A0(mai_mai_n334_), .A1(mai_mai_n333_), .B0(mai_mai_n312_), .Y(mai_mai_n335_));
  NOi21      m0313(.An(mai_mai_n152_), .B(mai_mai_n103_), .Y(mai_mai_n336_));
  NO2        m0314(.A(mai_mai_n336_), .B(mai_mai_n124_), .Y(mai_mai_n337_));
  OAI210     m0315(.A0(mai_mai_n337_), .A1(mai_mai_n335_), .B0(i_3_), .Y(mai_mai_n338_));
  NO2        m0316(.A(mai_mai_n286_), .B(mai_mai_n79_), .Y(mai_mai_n339_));
  NA2        m0317(.A(mai_mai_n339_), .B(mai_mai_n132_), .Y(mai_mai_n340_));
  NO2        m0318(.A(mai_mai_n91_), .B(mai_mai_n192_), .Y(mai_mai_n341_));
  NA3        m0319(.A(mai_mai_n216_), .B(mai_mai_n341_), .C(mai_mai_n63_), .Y(mai_mai_n342_));
  AOI210     m0320(.A0(mai_mai_n342_), .A1(mai_mai_n340_), .B0(i_7_), .Y(mai_mai_n343_));
  NO2        m0321(.A(mai_mai_n192_), .B(i_9_), .Y(mai_mai_n344_));
  NA2        m0322(.A(mai_mai_n344_), .B(mai_mai_n156_), .Y(mai_mai_n345_));
  NO2        m0323(.A(mai_mai_n345_), .B(mai_mai_n47_), .Y(mai_mai_n346_));
  NO3        m0324(.A(mai_mai_n346_), .B(mai_mai_n343_), .C(mai_mai_n285_), .Y(mai_mai_n347_));
  AOI210     m0325(.A0(mai_mai_n347_), .A1(mai_mai_n338_), .B0(mai_mai_n161_), .Y(mai_mai_n348_));
  AOI210     m0326(.A0(mai_mai_n330_), .A1(mai_mai_n304_), .B0(mai_mai_n348_), .Y(mai_mai_n349_));
  NOi32      m0327(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n350_));
  INV        m0328(.A(mai_mai_n350_), .Y(mai_mai_n351_));
  NAi21      m0329(.An(i_0_), .B(i_6_), .Y(mai_mai_n352_));
  NAi21      m0330(.An(i_1_), .B(i_5_), .Y(mai_mai_n353_));
  NA2        m0331(.A(mai_mai_n353_), .B(mai_mai_n352_), .Y(mai_mai_n354_));
  NA2        m0332(.A(mai_mai_n354_), .B(mai_mai_n25_), .Y(mai_mai_n355_));
  OAI210     m0333(.A0(mai_mai_n355_), .A1(mai_mai_n158_), .B0(mai_mai_n242_), .Y(mai_mai_n356_));
  NAi41      m0334(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n357_));
  OAI220     m0335(.A0(mai_mai_n357_), .A1(mai_mai_n353_), .B0(mai_mai_n218_), .B1(mai_mai_n158_), .Y(mai_mai_n358_));
  AOI210     m0336(.A0(mai_mai_n357_), .A1(mai_mai_n158_), .B0(mai_mai_n156_), .Y(mai_mai_n359_));
  NOi32      m0337(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n360_));
  NAi21      m0338(.An(i_6_), .B(i_1_), .Y(mai_mai_n361_));
  NA3        m0339(.A(mai_mai_n361_), .B(mai_mai_n360_), .C(mai_mai_n47_), .Y(mai_mai_n362_));
  NO2        m0340(.A(mai_mai_n362_), .B(i_0_), .Y(mai_mai_n363_));
  OR3        m0341(.A(mai_mai_n363_), .B(mai_mai_n359_), .C(mai_mai_n358_), .Y(mai_mai_n364_));
  NO2        m0342(.A(i_1_), .B(mai_mai_n100_), .Y(mai_mai_n365_));
  NAi21      m0343(.An(i_3_), .B(i_4_), .Y(mai_mai_n366_));
  NO2        m0344(.A(mai_mai_n366_), .B(i_9_), .Y(mai_mai_n367_));
  NA2        m0345(.A(i_2_), .B(i_7_), .Y(mai_mai_n368_));
  NO2        m0346(.A(mai_mai_n366_), .B(i_10_), .Y(mai_mai_n369_));
  NA3        m0347(.A(mai_mai_n369_), .B(mai_mai_n368_), .C(mai_mai_n240_), .Y(mai_mai_n370_));
  NO2        m0348(.A(mai_mai_n370_), .B(mai_mai_n184_), .Y(mai_mai_n371_));
  AOI210     m0349(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n372_));
  AOI220     m0350(.A0(mai_mai_n369_), .A1(mai_mai_n328_), .B0(mai_mai_n234_), .B1(mai_mai_n187_), .Y(mai_mai_n373_));
  NO2        m0351(.A(mai_mai_n373_), .B(i_5_), .Y(mai_mai_n374_));
  NO4        m0352(.A(mai_mai_n374_), .B(mai_mai_n371_), .C(mai_mai_n364_), .D(mai_mai_n356_), .Y(mai_mai_n375_));
  NO2        m0353(.A(mai_mai_n375_), .B(mai_mai_n351_), .Y(mai_mai_n376_));
  NO2        m0354(.A(mai_mai_n59_), .B(mai_mai_n25_), .Y(mai_mai_n377_));
  AN2        m0355(.A(i_12_), .B(i_5_), .Y(mai_mai_n378_));
  NO2        m0356(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n379_));
  NA2        m0357(.A(mai_mai_n379_), .B(mai_mai_n378_), .Y(mai_mai_n380_));
  NO2        m0358(.A(i_11_), .B(i_6_), .Y(mai_mai_n381_));
  NA3        m0359(.A(mai_mai_n381_), .B(mai_mai_n317_), .C(mai_mai_n222_), .Y(mai_mai_n382_));
  NO2        m0360(.A(mai_mai_n382_), .B(mai_mai_n380_), .Y(mai_mai_n383_));
  NO2        m0361(.A(mai_mai_n238_), .B(i_5_), .Y(mai_mai_n384_));
  NO2        m0362(.A(i_5_), .B(i_10_), .Y(mai_mai_n385_));
  NA2        m0363(.A(mai_mai_n144_), .B(mai_mai_n46_), .Y(mai_mai_n386_));
  NO2        m0364(.A(mai_mai_n386_), .B(mai_mai_n238_), .Y(mai_mai_n387_));
  OAI210     m0365(.A0(mai_mai_n387_), .A1(mai_mai_n383_), .B0(mai_mai_n377_), .Y(mai_mai_n388_));
  NO2        m0366(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n389_));
  NO2        m0367(.A(mai_mai_n150_), .B(mai_mai_n83_), .Y(mai_mai_n390_));
  OAI210     m0368(.A0(mai_mai_n390_), .A1(mai_mai_n383_), .B0(mai_mai_n389_), .Y(mai_mai_n391_));
  NO3        m0369(.A(mai_mai_n83_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n392_));
  NO2        m0370(.A(i_11_), .B(i_12_), .Y(mai_mai_n393_));
  NA2        m0371(.A(mai_mai_n393_), .B(mai_mai_n36_), .Y(mai_mai_n394_));
  NO2        m0372(.A(i_9_), .B(mai_mai_n394_), .Y(mai_mai_n395_));
  NA2        m0373(.A(mai_mai_n385_), .B(mai_mai_n233_), .Y(mai_mai_n396_));
  OAI220     m0374(.A0(mai_mai_n36_), .A1(mai_mai_n218_), .B0(mai_mai_n396_), .B1(mai_mai_n324_), .Y(mai_mai_n397_));
  NAi21      m0375(.An(i_13_), .B(i_0_), .Y(mai_mai_n398_));
  NO2        m0376(.A(mai_mai_n398_), .B(mai_mai_n235_), .Y(mai_mai_n399_));
  OAI210     m0377(.A0(mai_mai_n397_), .A1(mai_mai_n395_), .B0(mai_mai_n399_), .Y(mai_mai_n400_));
  NA3        m0378(.A(mai_mai_n400_), .B(mai_mai_n391_), .C(mai_mai_n388_), .Y(mai_mai_n401_));
  NO2        m0379(.A(i_0_), .B(i_11_), .Y(mai_mai_n402_));
  AN2        m0380(.A(i_1_), .B(i_6_), .Y(mai_mai_n403_));
  NOi21      m0381(.An(i_2_), .B(i_12_), .Y(mai_mai_n404_));
  NA2        m0382(.A(mai_mai_n404_), .B(mai_mai_n403_), .Y(mai_mai_n405_));
  INV        m0383(.A(mai_mai_n405_), .Y(mai_mai_n406_));
  NA2        m0384(.A(mai_mai_n142_), .B(i_9_), .Y(mai_mai_n407_));
  NO2        m0385(.A(mai_mai_n407_), .B(i_4_), .Y(mai_mai_n408_));
  NA2        m0386(.A(mai_mai_n406_), .B(mai_mai_n408_), .Y(mai_mai_n409_));
  OR2        m0387(.A(i_13_), .B(i_10_), .Y(mai_mai_n410_));
  NO2        m0388(.A(mai_mai_n171_), .B(mai_mai_n123_), .Y(mai_mai_n411_));
  BUFFER     m0389(.A(mai_mai_n214_), .Y(mai_mai_n412_));
  NO2        m0390(.A(mai_mai_n100_), .B(mai_mai_n25_), .Y(mai_mai_n413_));
  NA2        m0391(.A(mai_mai_n276_), .B(mai_mai_n413_), .Y(mai_mai_n414_));
  NA2        m0392(.A(mai_mai_n269_), .B(mai_mai_n208_), .Y(mai_mai_n415_));
  OAI220     m0393(.A0(mai_mai_n415_), .A1(mai_mai_n412_), .B0(mai_mai_n414_), .B1(mai_mai_n336_), .Y(mai_mai_n416_));
  INV        m0394(.A(mai_mai_n416_), .Y(mai_mai_n417_));
  AOI210     m0395(.A0(mai_mai_n417_), .A1(mai_mai_n409_), .B0(mai_mai_n26_), .Y(mai_mai_n418_));
  NA2        m0396(.A(mai_mai_n314_), .B(mai_mai_n313_), .Y(mai_mai_n419_));
  AOI220     m0397(.A0(mai_mai_n288_), .A1(mai_mai_n279_), .B0(mai_mai_n282_), .B1(mai_mai_n305_), .Y(mai_mai_n420_));
  NO2        m0398(.A(mai_mai_n420_), .B(i_5_), .Y(mai_mai_n421_));
  NO2        m0399(.A(mai_mai_n182_), .B(mai_mai_n83_), .Y(mai_mai_n422_));
  AOI220     m0400(.A0(mai_mai_n422_), .A1(mai_mai_n287_), .B0(mai_mai_n271_), .B1(mai_mai_n208_), .Y(mai_mai_n423_));
  NO2        m0401(.A(mai_mai_n423_), .B(mai_mai_n278_), .Y(mai_mai_n424_));
  NO3        m0402(.A(mai_mai_n424_), .B(mai_mai_n421_), .C(mai_mai_n419_), .Y(mai_mai_n425_));
  NA2        m0403(.A(mai_mai_n194_), .B(mai_mai_n95_), .Y(mai_mai_n426_));
  NA3        m0404(.A(mai_mai_n317_), .B(mai_mai_n162_), .C(mai_mai_n83_), .Y(mai_mai_n427_));
  AOI210     m0405(.A0(mai_mai_n427_), .A1(mai_mai_n426_), .B0(mai_mai_n315_), .Y(mai_mai_n428_));
  NA2        m0406(.A(mai_mai_n192_), .B(i_10_), .Y(mai_mai_n429_));
  NA2        m0407(.A(mai_mai_n64_), .B(i_2_), .Y(mai_mai_n430_));
  NA2        m0408(.A(mai_mai_n288_), .B(mai_mai_n232_), .Y(mai_mai_n431_));
  OAI220     m0409(.A0(mai_mai_n431_), .A1(mai_mai_n182_), .B0(mai_mai_n430_), .B1(mai_mai_n429_), .Y(mai_mai_n432_));
  NO2        m0410(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n433_));
  NA3        m0411(.A(mai_mai_n328_), .B(mai_mai_n327_), .C(mai_mai_n433_), .Y(mai_mai_n434_));
  NA2        m0412(.A(mai_mai_n307_), .B(mai_mai_n312_), .Y(mai_mai_n435_));
  OAI210     m0413(.A0(mai_mai_n435_), .A1(mai_mai_n188_), .B0(mai_mai_n434_), .Y(mai_mai_n436_));
  NO3        m0414(.A(mai_mai_n436_), .B(mai_mai_n432_), .C(mai_mai_n428_), .Y(mai_mai_n437_));
  AOI210     m0415(.A0(mai_mai_n437_), .A1(mai_mai_n425_), .B0(mai_mai_n264_), .Y(mai_mai_n438_));
  NO4        m0416(.A(mai_mai_n438_), .B(mai_mai_n418_), .C(mai_mai_n401_), .D(mai_mai_n376_), .Y(mai_mai_n439_));
  NO2        m0417(.A(mai_mai_n71_), .B(i_13_), .Y(mai_mai_n440_));
  NO2        m0418(.A(i_10_), .B(i_9_), .Y(mai_mai_n441_));
  NAi21      m0419(.An(i_12_), .B(i_8_), .Y(mai_mai_n442_));
  NO2        m0420(.A(mai_mai_n442_), .B(i_3_), .Y(mai_mai_n443_));
  NA2        m0421(.A(i_2_), .B(mai_mai_n103_), .Y(mai_mai_n444_));
  NO2        m0422(.A(mai_mai_n444_), .B(mai_mai_n203_), .Y(mai_mai_n445_));
  NA2        m0423(.A(mai_mai_n300_), .B(i_0_), .Y(mai_mai_n446_));
  NO3        m0424(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n447_));
  NA2        m0425(.A(mai_mai_n259_), .B(mai_mai_n96_), .Y(mai_mai_n448_));
  NA2        m0426(.A(mai_mai_n448_), .B(mai_mai_n447_), .Y(mai_mai_n449_));
  NA2        m0427(.A(i_8_), .B(i_9_), .Y(mai_mai_n450_));
  NO2        m0428(.A(mai_mai_n449_), .B(mai_mai_n446_), .Y(mai_mai_n451_));
  NO3        m0429(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n452_));
  NA3        m0430(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n453_));
  NA4        m0431(.A(mai_mai_n145_), .B(mai_mai_n115_), .C(mai_mai_n78_), .D(mai_mai_n23_), .Y(mai_mai_n454_));
  NO2        m0432(.A(mai_mai_n454_), .B(mai_mai_n453_), .Y(mai_mai_n455_));
  NO3        m0433(.A(mai_mai_n455_), .B(mai_mai_n451_), .C(mai_mai_n445_), .Y(mai_mai_n456_));
  OA210      m0434(.A0(mai_mai_n345_), .A1(mai_mai_n100_), .B0(mai_mai_n289_), .Y(mai_mai_n457_));
  OA220      m0435(.A0(mai_mai_n457_), .A1(mai_mai_n161_), .B0(mai_mai_n205_), .B1(mai_mai_n229_), .Y(mai_mai_n458_));
  NA2        m0436(.A(mai_mai_n95_), .B(i_13_), .Y(mai_mai_n459_));
  NA2        m0437(.A(mai_mai_n422_), .B(mai_mai_n377_), .Y(mai_mai_n460_));
  NO2        m0438(.A(i_2_), .B(i_13_), .Y(mai_mai_n461_));
  NA3        m0439(.A(mai_mai_n461_), .B(mai_mai_n160_), .C(mai_mai_n98_), .Y(mai_mai_n462_));
  OAI220     m0440(.A0(mai_mai_n462_), .A1(mai_mai_n233_), .B0(mai_mai_n460_), .B1(mai_mai_n459_), .Y(mai_mai_n463_));
  NO3        m0441(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n464_));
  NO2        m0442(.A(i_6_), .B(i_7_), .Y(mai_mai_n465_));
  NA2        m0443(.A(mai_mai_n465_), .B(mai_mai_n464_), .Y(mai_mai_n466_));
  NO2        m0444(.A(i_11_), .B(i_1_), .Y(mai_mai_n467_));
  OR2        m0445(.A(i_11_), .B(i_8_), .Y(mai_mai_n468_));
  NOi21      m0446(.An(i_2_), .B(i_7_), .Y(mai_mai_n469_));
  NAi31      m0447(.An(mai_mai_n468_), .B(mai_mai_n469_), .C(i_0_), .Y(mai_mai_n470_));
  NO2        m0448(.A(mai_mai_n410_), .B(i_6_), .Y(mai_mai_n471_));
  NA3        m0449(.A(mai_mai_n471_), .B(i_1_), .C(mai_mai_n73_), .Y(mai_mai_n472_));
  NO2        m0450(.A(mai_mai_n472_), .B(mai_mai_n470_), .Y(mai_mai_n473_));
  NO2        m0451(.A(i_3_), .B(mai_mai_n192_), .Y(mai_mai_n474_));
  NO2        m0452(.A(i_6_), .B(i_10_), .Y(mai_mai_n475_));
  NA4        m0453(.A(mai_mai_n475_), .B(mai_mai_n304_), .C(mai_mai_n474_), .D(mai_mai_n233_), .Y(mai_mai_n476_));
  NO2        m0454(.A(mai_mai_n476_), .B(mai_mai_n154_), .Y(mai_mai_n477_));
  NA2        m0455(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n478_));
  NO2        m0456(.A(mai_mai_n156_), .B(i_3_), .Y(mai_mai_n479_));
  NO3        m0457(.A(mai_mai_n477_), .B(mai_mai_n473_), .C(mai_mai_n463_), .Y(mai_mai_n480_));
  NA2        m0458(.A(mai_mai_n447_), .B(mai_mai_n378_), .Y(mai_mai_n481_));
  NA2        m0459(.A(mai_mai_n452_), .B(mai_mai_n385_), .Y(mai_mai_n482_));
  NO2        m0460(.A(mai_mai_n482_), .B(mai_mai_n221_), .Y(mai_mai_n483_));
  NAi21      m0461(.An(mai_mai_n214_), .B(mai_mai_n393_), .Y(mai_mai_n484_));
  NA2        m0462(.A(mai_mai_n328_), .B(mai_mai_n216_), .Y(mai_mai_n485_));
  NO2        m0463(.A(i_0_), .B(mai_mai_n83_), .Y(mai_mai_n486_));
  NA3        m0464(.A(mai_mai_n486_), .B(mai_mai_n1030_), .C(mai_mai_n142_), .Y(mai_mai_n487_));
  OR3        m0465(.A(mai_mai_n295_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n488_));
  OAI220     m0466(.A0(mai_mai_n488_), .A1(mai_mai_n487_), .B0(mai_mai_n485_), .B1(mai_mai_n484_), .Y(mai_mai_n489_));
  NA2        m0467(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n490_));
  NA2        m0468(.A(mai_mai_n304_), .B(mai_mai_n234_), .Y(mai_mai_n491_));
  OAI220     m0469(.A0(mai_mai_n491_), .A1(mai_mai_n430_), .B0(mai_mai_n490_), .B1(mai_mai_n459_), .Y(mai_mai_n492_));
  NA4        m0470(.A(mai_mai_n297_), .B(mai_mai_n220_), .C(mai_mai_n71_), .D(mai_mai_n233_), .Y(mai_mai_n493_));
  NO2        m0471(.A(mai_mai_n493_), .B(mai_mai_n466_), .Y(mai_mai_n494_));
  NO4        m0472(.A(mai_mai_n494_), .B(mai_mai_n492_), .C(mai_mai_n489_), .D(mai_mai_n483_), .Y(mai_mai_n495_));
  NA4        m0473(.A(mai_mai_n495_), .B(mai_mai_n480_), .C(mai_mai_n458_), .D(mai_mai_n456_), .Y(mai_mai_n496_));
  NA3        m0474(.A(mai_mai_n297_), .B(mai_mai_n175_), .C(mai_mai_n173_), .Y(mai_mai_n497_));
  OAI210     m0475(.A0(mai_mai_n293_), .A1(mai_mai_n180_), .B0(mai_mai_n497_), .Y(mai_mai_n498_));
  NA2        m0476(.A(mai_mai_n231_), .B(mai_mai_n498_), .Y(mai_mai_n499_));
  NA2        m0477(.A(mai_mai_n122_), .B(mai_mai_n111_), .Y(mai_mai_n500_));
  AN2        m0478(.A(mai_mai_n500_), .B(mai_mai_n447_), .Y(mai_mai_n501_));
  INV        m0479(.A(mai_mai_n304_), .Y(mai_mai_n502_));
  OAI210     m0480(.A0(mai_mai_n502_), .A1(mai_mai_n229_), .B0(mai_mai_n298_), .Y(mai_mai_n503_));
  AOI220     m0481(.A0(mai_mai_n503_), .A1(mai_mai_n316_), .B0(mai_mai_n501_), .B1(mai_mai_n300_), .Y(mai_mai_n504_));
  NA2        m0482(.A(mai_mai_n350_), .B(mai_mai_n71_), .Y(mai_mai_n505_));
  INV        m0483(.A(mai_mai_n360_), .Y(mai_mai_n506_));
  NO2        m0484(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n507_));
  NA2        m0485(.A(mai_mai_n39_), .B(i_13_), .Y(mai_mai_n508_));
  OAI210     m0486(.A0(i_8_), .A1(mai_mai_n63_), .B0(mai_mai_n134_), .Y(mai_mai_n509_));
  NO2        m0487(.A(i_7_), .B(mai_mai_n197_), .Y(mai_mai_n510_));
  OR2        m0488(.A(mai_mai_n182_), .B(i_4_), .Y(mai_mai_n511_));
  NO2        m0489(.A(mai_mai_n511_), .B(mai_mai_n83_), .Y(mai_mai_n512_));
  AOI220     m0490(.A0(mai_mai_n512_), .A1(mai_mai_n510_), .B0(mai_mai_n509_), .B1(mai_mai_n411_), .Y(mai_mai_n513_));
  NA4        m0491(.A(mai_mai_n513_), .B(mai_mai_n508_), .C(mai_mai_n504_), .D(mai_mai_n499_), .Y(mai_mai_n514_));
  NA2        m0492(.A(mai_mai_n384_), .B(mai_mai_n287_), .Y(mai_mai_n515_));
  NA2        m0493(.A(mai_mai_n380_), .B(mai_mai_n515_), .Y(mai_mai_n516_));
  NO2        m0494(.A(i_12_), .B(mai_mai_n192_), .Y(mai_mai_n517_));
  NA2        m0495(.A(mai_mai_n517_), .B(mai_mai_n222_), .Y(mai_mai_n518_));
  NO2        m0496(.A(i_10_), .B(mai_mai_n518_), .Y(mai_mai_n519_));
  NOi31      m0497(.An(mai_mai_n307_), .B(mai_mai_n410_), .C(mai_mai_n38_), .Y(mai_mai_n520_));
  OAI210     m0498(.A0(mai_mai_n520_), .A1(mai_mai_n519_), .B0(mai_mai_n516_), .Y(mai_mai_n521_));
  NO2        m0499(.A(i_8_), .B(i_7_), .Y(mai_mai_n522_));
  OAI210     m0500(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n523_));
  NA2        m0501(.A(mai_mai_n523_), .B(mai_mai_n220_), .Y(mai_mai_n524_));
  OAI220     m0502(.A0(mai_mai_n47_), .A1(mai_mai_n511_), .B0(mai_mai_n524_), .B1(mai_mai_n238_), .Y(mai_mai_n525_));
  NA2        m0503(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n526_));
  NO2        m0504(.A(mai_mai_n526_), .B(i_6_), .Y(mai_mai_n527_));
  NA3        m0505(.A(mai_mai_n527_), .B(mai_mai_n525_), .C(mai_mai_n522_), .Y(mai_mai_n528_));
  AOI220     m0506(.A0(mai_mai_n422_), .A1(mai_mai_n317_), .B0(mai_mai_n243_), .B1(mai_mai_n240_), .Y(mai_mai_n529_));
  OAI220     m0507(.A0(mai_mai_n529_), .A1(mai_mai_n255_), .B0(mai_mai_n459_), .B1(mai_mai_n133_), .Y(mai_mai_n530_));
  NA2        m0508(.A(mai_mai_n530_), .B(mai_mai_n258_), .Y(mai_mai_n531_));
  NOi31      m0509(.An(mai_mai_n282_), .B(mai_mai_n293_), .C(mai_mai_n180_), .Y(mai_mai_n532_));
  NA3        m0510(.A(mai_mai_n297_), .B(mai_mai_n173_), .C(mai_mai_n95_), .Y(mai_mai_n533_));
  NO2        m0511(.A(mai_mai_n156_), .B(i_5_), .Y(mai_mai_n534_));
  NA2        m0512(.A(mai_mai_n534_), .B(mai_mai_n310_), .Y(mai_mai_n535_));
  NA2        m0513(.A(mai_mai_n535_), .B(mai_mai_n533_), .Y(mai_mai_n536_));
  OAI210     m0514(.A0(mai_mai_n536_), .A1(mai_mai_n532_), .B0(mai_mai_n452_), .Y(mai_mai_n537_));
  NA4        m0515(.A(mai_mai_n537_), .B(mai_mai_n531_), .C(mai_mai_n528_), .D(mai_mai_n521_), .Y(mai_mai_n538_));
  NA2        m0516(.A(mai_mai_n276_), .B(mai_mai_n82_), .Y(mai_mai_n539_));
  NO2        m0517(.A(mai_mai_n340_), .B(mai_mai_n539_), .Y(mai_mai_n540_));
  NA2        m0518(.A(mai_mai_n288_), .B(mai_mai_n279_), .Y(mai_mai_n541_));
  NO2        m0519(.A(mai_mai_n541_), .B(mai_mai_n172_), .Y(mai_mai_n542_));
  NA2        m0520(.A(mai_mai_n220_), .B(i_0_), .Y(mai_mai_n543_));
  NA2        m0521(.A(mai_mai_n441_), .B(mai_mai_n219_), .Y(mai_mai_n544_));
  NO2        m0522(.A(mai_mai_n543_), .B(mai_mai_n544_), .Y(mai_mai_n545_));
  AOI210     m0523(.A0(mai_mai_n361_), .A1(mai_mai_n47_), .B0(mai_mai_n365_), .Y(mai_mai_n546_));
  NA2        m0524(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n547_));
  NA3        m0525(.A(mai_mai_n517_), .B(mai_mai_n267_), .C(mai_mai_n547_), .Y(mai_mai_n548_));
  NO2        m0526(.A(mai_mai_n546_), .B(mai_mai_n548_), .Y(mai_mai_n549_));
  NO4        m0527(.A(mai_mai_n549_), .B(mai_mai_n545_), .C(mai_mai_n542_), .D(mai_mai_n540_), .Y(mai_mai_n550_));
  NO4        m0528(.A(mai_mai_n248_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n551_));
  NO3        m0529(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n552_));
  NO2        m0530(.A(mai_mai_n230_), .B(mai_mai_n36_), .Y(mai_mai_n553_));
  AN2        m0531(.A(mai_mai_n553_), .B(mai_mai_n552_), .Y(mai_mai_n554_));
  OA210      m0532(.A0(mai_mai_n554_), .A1(mai_mai_n551_), .B0(mai_mai_n350_), .Y(mai_mai_n555_));
  NO2        m0533(.A(mai_mai_n410_), .B(i_1_), .Y(mai_mai_n556_));
  NOi31      m0534(.An(mai_mai_n556_), .B(mai_mai_n448_), .C(mai_mai_n71_), .Y(mai_mai_n557_));
  AN3        m0535(.A(mai_mai_n557_), .B(mai_mai_n408_), .C(i_2_), .Y(mai_mai_n558_));
  NO2        m0536(.A(mai_mai_n420_), .B(mai_mai_n176_), .Y(mai_mai_n559_));
  NO3        m0537(.A(mai_mai_n559_), .B(mai_mai_n558_), .C(mai_mai_n555_), .Y(mai_mai_n560_));
  NOi21      m0538(.An(i_10_), .B(i_6_), .Y(mai_mai_n561_));
  NO2        m0539(.A(mai_mai_n83_), .B(mai_mai_n25_), .Y(mai_mai_n562_));
  AOI220     m0540(.A0(mai_mai_n276_), .A1(mai_mai_n562_), .B0(mai_mai_n267_), .B1(mai_mai_n561_), .Y(mai_mai_n563_));
  NO2        m0541(.A(mai_mai_n563_), .B(mai_mai_n446_), .Y(mai_mai_n564_));
  NO2        m0542(.A(mai_mai_n114_), .B(mai_mai_n23_), .Y(mai_mai_n565_));
  NA2        m0543(.A(mai_mai_n307_), .B(mai_mai_n163_), .Y(mai_mai_n566_));
  AOI220     m0544(.A0(mai_mai_n566_), .A1(mai_mai_n431_), .B0(mai_mai_n171_), .B1(mai_mai_n181_), .Y(mai_mai_n567_));
  NOi21      m0545(.An(mai_mai_n146_), .B(mai_mai_n324_), .Y(mai_mai_n568_));
  NO3        m0546(.A(mai_mai_n568_), .B(mai_mai_n567_), .C(mai_mai_n564_), .Y(mai_mai_n569_));
  NO2        m0547(.A(mai_mai_n505_), .B(mai_mai_n373_), .Y(mai_mai_n570_));
  INV        m0548(.A(mai_mai_n310_), .Y(mai_mai_n571_));
  NO2        m0549(.A(i_12_), .B(mai_mai_n83_), .Y(mai_mai_n572_));
  NA3        m0550(.A(mai_mai_n572_), .B(mai_mai_n267_), .C(mai_mai_n547_), .Y(mai_mai_n573_));
  NA3        m0551(.A(mai_mai_n381_), .B(mai_mai_n276_), .C(mai_mai_n216_), .Y(mai_mai_n574_));
  AOI210     m0552(.A0(mai_mai_n574_), .A1(mai_mai_n573_), .B0(mai_mai_n571_), .Y(mai_mai_n575_));
  NO3        m0553(.A(i_4_), .B(mai_mai_n333_), .C(mai_mai_n293_), .Y(mai_mai_n576_));
  OR2        m0554(.A(i_2_), .B(i_5_), .Y(mai_mai_n577_));
  OR2        m0555(.A(mai_mai_n577_), .B(mai_mai_n403_), .Y(mai_mai_n578_));
  AOI210     m0556(.A0(mai_mai_n368_), .A1(mai_mai_n240_), .B0(mai_mai_n196_), .Y(mai_mai_n579_));
  AOI210     m0557(.A0(mai_mai_n579_), .A1(mai_mai_n578_), .B0(mai_mai_n484_), .Y(mai_mai_n580_));
  NO4        m0558(.A(mai_mai_n580_), .B(mai_mai_n576_), .C(mai_mai_n575_), .D(mai_mai_n570_), .Y(mai_mai_n581_));
  NA4        m0559(.A(mai_mai_n581_), .B(mai_mai_n569_), .C(mai_mai_n560_), .D(mai_mai_n550_), .Y(mai_mai_n582_));
  NO4        m0560(.A(mai_mai_n582_), .B(mai_mai_n538_), .C(mai_mai_n514_), .D(mai_mai_n496_), .Y(mai_mai_n583_));
  NA4        m0561(.A(mai_mai_n583_), .B(mai_mai_n439_), .C(mai_mai_n349_), .D(mai_mai_n303_), .Y(mai7));
  OAI220     m0562(.A0(mai_mai_n490_), .A1(mai_mai_n117_), .B0(mai_mai_n91_), .B1(mai_mai_n54_), .Y(mai_mai_n585_));
  NO2        m0563(.A(mai_mai_n107_), .B(mai_mai_n88_), .Y(mai_mai_n586_));
  NA2        m0564(.A(mai_mai_n379_), .B(mai_mai_n586_), .Y(mai_mai_n587_));
  NA2        m0565(.A(mai_mai_n475_), .B(mai_mai_n82_), .Y(mai_mai_n588_));
  NA2        m0566(.A(i_11_), .B(mai_mai_n192_), .Y(mai_mai_n589_));
  NA2        m0567(.A(mai_mai_n144_), .B(mai_mai_n589_), .Y(mai_mai_n590_));
  OAI210     m0568(.A0(mai_mai_n590_), .A1(mai_mai_n588_), .B0(mai_mai_n587_), .Y(mai_mai_n591_));
  NA3        m0569(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n592_));
  NO2        m0570(.A(mai_mai_n233_), .B(i_4_), .Y(mai_mai_n593_));
  NA2        m0571(.A(mai_mai_n593_), .B(i_8_), .Y(mai_mai_n594_));
  NA2        m0572(.A(i_2_), .B(mai_mai_n83_), .Y(mai_mai_n595_));
  OAI210     m0573(.A0(mai_mai_n86_), .A1(mai_mai_n201_), .B0(mai_mai_n202_), .Y(mai_mai_n596_));
  NO2        m0574(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n597_));
  NA2        m0575(.A(i_4_), .B(i_8_), .Y(mai_mai_n598_));
  NO2        m0576(.A(mai_mai_n591_), .B(mai_mai_n585_), .Y(mai_mai_n599_));
  INV        m0577(.A(mai_mai_n160_), .Y(mai_mai_n600_));
  OR2        m0578(.A(i_6_), .B(i_10_), .Y(mai_mai_n601_));
  NO2        m0579(.A(mai_mai_n601_), .B(mai_mai_n23_), .Y(mai_mai_n602_));
  OR3        m0580(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n603_));
  NO3        m0581(.A(mai_mai_n603_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n604_));
  INV        m0582(.A(mai_mai_n198_), .Y(mai_mai_n605_));
  NO2        m0583(.A(mai_mai_n604_), .B(mai_mai_n602_), .Y(mai_mai_n606_));
  OA220      m0584(.A0(mai_mai_n606_), .A1(mai_mai_n571_), .B0(mai_mai_n600_), .B1(mai_mai_n260_), .Y(mai_mai_n607_));
  AOI210     m0585(.A0(mai_mai_n607_), .A1(mai_mai_n599_), .B0(mai_mai_n63_), .Y(mai_mai_n608_));
  NOi21      m0586(.An(i_11_), .B(i_7_), .Y(mai_mai_n609_));
  AO210      m0587(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n610_));
  NO2        m0588(.A(mai_mai_n610_), .B(mai_mai_n609_), .Y(mai_mai_n611_));
  NA2        m0589(.A(mai_mai_n611_), .B(mai_mai_n204_), .Y(mai_mai_n612_));
  NA3        m0590(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n613_));
  NAi31      m0591(.An(mai_mai_n613_), .B(mai_mai_n213_), .C(i_11_), .Y(mai_mai_n614_));
  AOI210     m0592(.A0(mai_mai_n614_), .A1(mai_mai_n612_), .B0(mai_mai_n63_), .Y(mai_mai_n615_));
  NA2        m0593(.A(mai_mai_n85_), .B(mai_mai_n63_), .Y(mai_mai_n616_));
  AO210      m0594(.A0(mai_mai_n616_), .A1(mai_mai_n373_), .B0(mai_mai_n41_), .Y(mai_mai_n617_));
  NO3        m0595(.A(mai_mai_n252_), .B(mai_mai_n206_), .C(mai_mai_n589_), .Y(mai_mai_n618_));
  OAI210     m0596(.A0(mai_mai_n618_), .A1(mai_mai_n223_), .B0(mai_mai_n63_), .Y(mai_mai_n619_));
  NA2        m0597(.A(mai_mai_n404_), .B(mai_mai_n31_), .Y(mai_mai_n620_));
  OR2        m0598(.A(mai_mai_n206_), .B(mai_mai_n107_), .Y(mai_mai_n621_));
  NA2        m0599(.A(mai_mai_n621_), .B(mai_mai_n620_), .Y(mai_mai_n622_));
  NO2        m0600(.A(mai_mai_n63_), .B(i_9_), .Y(mai_mai_n623_));
  NO2        m0601(.A(mai_mai_n623_), .B(i_4_), .Y(mai_mai_n624_));
  NA2        m0602(.A(mai_mai_n624_), .B(mai_mai_n622_), .Y(mai_mai_n625_));
  NO2        m0603(.A(i_1_), .B(i_12_), .Y(mai_mai_n626_));
  NA3        m0604(.A(mai_mai_n626_), .B(mai_mai_n109_), .C(mai_mai_n24_), .Y(mai_mai_n627_));
  NA4        m0605(.A(mai_mai_n627_), .B(mai_mai_n625_), .C(mai_mai_n619_), .D(mai_mai_n617_), .Y(mai_mai_n628_));
  OAI210     m0606(.A0(mai_mai_n628_), .A1(mai_mai_n615_), .B0(i_6_), .Y(mai_mai_n629_));
  OAI210     m0607(.A0(mai_mai_n613_), .A1(mai_mai_n107_), .B0(mai_mai_n453_), .Y(mai_mai_n630_));
  NA2        m0608(.A(mai_mai_n630_), .B(mai_mai_n572_), .Y(mai_mai_n631_));
  NO2        m0609(.A(mai_mai_n233_), .B(mai_mai_n83_), .Y(mai_mai_n632_));
  NO2        m0610(.A(mai_mai_n632_), .B(i_11_), .Y(mai_mai_n633_));
  NA2        m0611(.A(mai_mai_n631_), .B(mai_mai_n449_), .Y(mai_mai_n634_));
  NO4        m0612(.A(mai_mai_n213_), .B(mai_mai_n128_), .C(i_13_), .D(mai_mai_n83_), .Y(mai_mai_n635_));
  NA2        m0613(.A(mai_mai_n635_), .B(mai_mai_n623_), .Y(mai_mai_n636_));
  NO3        m0614(.A(mai_mai_n601_), .B(mai_mai_n230_), .C(mai_mai_n23_), .Y(mai_mai_n637_));
  INV        m0615(.A(mai_mai_n636_), .Y(mai_mai_n638_));
  NA3        m0616(.A(mai_mai_n522_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n639_));
  NA2        m0617(.A(mai_mai_n138_), .B(i_9_), .Y(mai_mai_n640_));
  NA3        m0618(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n641_));
  NO2        m0619(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n642_));
  NA3        m0620(.A(mai_mai_n642_), .B(mai_mai_n259_), .C(mai_mai_n45_), .Y(mai_mai_n643_));
  OAI220     m0621(.A0(mai_mai_n643_), .A1(mai_mai_n641_), .B0(mai_mai_n640_), .B1(mai_mai_n1029_), .Y(mai_mai_n644_));
  NA3        m0622(.A(mai_mai_n623_), .B(mai_mai_n310_), .C(i_6_), .Y(mai_mai_n645_));
  NO2        m0623(.A(mai_mai_n645_), .B(mai_mai_n23_), .Y(mai_mai_n646_));
  AOI210     m0624(.A0(mai_mai_n467_), .A1(mai_mai_n413_), .B0(mai_mai_n237_), .Y(mai_mai_n647_));
  NO2        m0625(.A(mai_mai_n647_), .B(mai_mai_n595_), .Y(mai_mai_n648_));
  NAi21      m0626(.An(mai_mai_n639_), .B(mai_mai_n90_), .Y(mai_mai_n649_));
  NA2        m0627(.A(mai_mai_n642_), .B(mai_mai_n259_), .Y(mai_mai_n650_));
  NO2        m0628(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n651_));
  NA2        m0629(.A(mai_mai_n651_), .B(mai_mai_n24_), .Y(mai_mai_n652_));
  OAI210     m0630(.A0(mai_mai_n652_), .A1(mai_mai_n650_), .B0(mai_mai_n649_), .Y(mai_mai_n653_));
  OR4        m0631(.A(mai_mai_n653_), .B(mai_mai_n648_), .C(mai_mai_n646_), .D(mai_mai_n644_), .Y(mai_mai_n654_));
  NO3        m0632(.A(mai_mai_n654_), .B(mai_mai_n638_), .C(mai_mai_n634_), .Y(mai_mai_n655_));
  NO2        m0633(.A(mai_mai_n233_), .B(mai_mai_n100_), .Y(mai_mai_n656_));
  NO2        m0634(.A(mai_mai_n656_), .B(mai_mai_n609_), .Y(mai_mai_n657_));
  NA2        m0635(.A(mai_mai_n657_), .B(i_1_), .Y(mai_mai_n658_));
  NO2        m0636(.A(mai_mai_n658_), .B(mai_mai_n603_), .Y(mai_mai_n659_));
  NA2        m0637(.A(mai_mai_n659_), .B(mai_mai_n47_), .Y(mai_mai_n660_));
  NA2        m0638(.A(i_3_), .B(mai_mai_n192_), .Y(mai_mai_n661_));
  NO2        m0639(.A(mai_mai_n661_), .B(mai_mai_n114_), .Y(mai_mai_n662_));
  AN2        m0640(.A(mai_mai_n662_), .B(mai_mai_n527_), .Y(mai_mai_n663_));
  NO2        m0641(.A(mai_mai_n117_), .B(mai_mai_n37_), .Y(mai_mai_n664_));
  NO2        m0642(.A(mai_mai_n83_), .B(i_9_), .Y(mai_mai_n665_));
  NA2        m0643(.A(i_1_), .B(i_3_), .Y(mai_mai_n666_));
  NO2        m0644(.A(mai_mai_n450_), .B(mai_mai_n91_), .Y(mai_mai_n667_));
  AOI210     m0645(.A0(i_11_), .A1(mai_mai_n561_), .B0(mai_mai_n667_), .Y(mai_mai_n668_));
  NO2        m0646(.A(mai_mai_n668_), .B(mai_mai_n666_), .Y(mai_mai_n669_));
  NO2        m0647(.A(mai_mai_n669_), .B(mai_mai_n663_), .Y(mai_mai_n670_));
  NA4        m0648(.A(mai_mai_n670_), .B(mai_mai_n660_), .C(mai_mai_n655_), .D(mai_mai_n629_), .Y(mai_mai_n671_));
  NO3        m0649(.A(mai_mai_n468_), .B(i_3_), .C(i_7_), .Y(mai_mai_n672_));
  NOi21      m0650(.An(mai_mai_n672_), .B(i_10_), .Y(mai_mai_n673_));
  OA210      m0651(.A0(mai_mai_n673_), .A1(mai_mai_n241_), .B0(mai_mai_n83_), .Y(mai_mai_n674_));
  NA2        m0652(.A(i_6_), .B(mai_mai_n367_), .Y(mai_mai_n675_));
  NA3        m0653(.A(mai_mai_n475_), .B(mai_mai_n507_), .C(mai_mai_n47_), .Y(mai_mai_n676_));
  NO3        m0654(.A(mai_mai_n469_), .B(mai_mai_n598_), .C(mai_mai_n83_), .Y(mai_mai_n677_));
  NA2        m0655(.A(mai_mai_n677_), .B(mai_mai_n25_), .Y(mai_mai_n678_));
  NA3        m0656(.A(mai_mai_n160_), .B(mai_mai_n82_), .C(mai_mai_n83_), .Y(mai_mai_n679_));
  NA4        m0657(.A(mai_mai_n679_), .B(mai_mai_n678_), .C(mai_mai_n676_), .D(mai_mai_n675_), .Y(mai_mai_n680_));
  OAI210     m0658(.A0(mai_mai_n680_), .A1(mai_mai_n674_), .B0(i_1_), .Y(mai_mai_n681_));
  AOI210     m0659(.A0(mai_mai_n259_), .A1(mai_mai_n96_), .B0(i_1_), .Y(mai_mai_n682_));
  NO2        m0660(.A(mai_mai_n366_), .B(i_2_), .Y(mai_mai_n683_));
  NA2        m0661(.A(mai_mai_n683_), .B(mai_mai_n682_), .Y(mai_mai_n684_));
  OAI210     m0662(.A0(mai_mai_n645_), .A1(mai_mai_n442_), .B0(mai_mai_n684_), .Y(mai_mai_n685_));
  INV        m0663(.A(mai_mai_n685_), .Y(mai_mai_n686_));
  AOI210     m0664(.A0(mai_mai_n686_), .A1(mai_mai_n681_), .B0(i_13_), .Y(mai_mai_n687_));
  OR2        m0665(.A(i_11_), .B(i_7_), .Y(mai_mai_n688_));
  NA3        m0666(.A(mai_mai_n688_), .B(mai_mai_n105_), .C(mai_mai_n138_), .Y(mai_mai_n689_));
  AOI220     m0667(.A0(mai_mai_n461_), .A1(mai_mai_n160_), .B0(i_2_), .B1(mai_mai_n138_), .Y(mai_mai_n690_));
  OAI210     m0668(.A0(mai_mai_n690_), .A1(mai_mai_n45_), .B0(mai_mai_n689_), .Y(mai_mai_n691_));
  NA2        m0669(.A(mai_mai_n241_), .B(mai_mai_n131_), .Y(mai_mai_n692_));
  NO2        m0670(.A(mai_mai_n692_), .B(mai_mai_n41_), .Y(mai_mai_n693_));
  AOI210     m0671(.A0(mai_mai_n691_), .A1(mai_mai_n326_), .B0(mai_mai_n693_), .Y(mai_mai_n694_));
  AOI220     m0672(.A0(i_12_), .A1(mai_mai_n70_), .B0(mai_mai_n381_), .B1(mai_mai_n642_), .Y(mai_mai_n695_));
  NO2        m0673(.A(mai_mai_n695_), .B(mai_mai_n238_), .Y(mai_mai_n696_));
  AOI210     m0674(.A0(mai_mai_n442_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n697_));
  NOi31      m0675(.An(mai_mai_n697_), .B(mai_mai_n588_), .C(mai_mai_n45_), .Y(mai_mai_n698_));
  NA2        m0676(.A(mai_mai_n127_), .B(i_13_), .Y(mai_mai_n699_));
  NO2        m0677(.A(mai_mai_n641_), .B(mai_mai_n114_), .Y(mai_mai_n700_));
  INV        m0678(.A(mai_mai_n700_), .Y(mai_mai_n701_));
  OAI220     m0679(.A0(mai_mai_n701_), .A1(mai_mai_n69_), .B0(mai_mai_n699_), .B1(mai_mai_n682_), .Y(mai_mai_n702_));
  NO3        m0680(.A(mai_mai_n69_), .B(mai_mai_n32_), .C(mai_mai_n100_), .Y(mai_mai_n703_));
  NA2        m0681(.A(mai_mai_n26_), .B(mai_mai_n192_), .Y(mai_mai_n704_));
  NA2        m0682(.A(mai_mai_n704_), .B(i_7_), .Y(mai_mai_n705_));
  NO3        m0683(.A(mai_mai_n469_), .B(mai_mai_n233_), .C(mai_mai_n83_), .Y(mai_mai_n706_));
  AOI210     m0684(.A0(mai_mai_n706_), .A1(mai_mai_n705_), .B0(mai_mai_n703_), .Y(mai_mai_n707_));
  AOI220     m0685(.A0(mai_mai_n381_), .A1(mai_mai_n642_), .B0(mai_mai_n90_), .B1(mai_mai_n101_), .Y(mai_mai_n708_));
  OAI220     m0686(.A0(mai_mai_n708_), .A1(mai_mai_n594_), .B0(mai_mai_n707_), .B1(mai_mai_n605_), .Y(mai_mai_n709_));
  NO4        m0687(.A(mai_mai_n709_), .B(mai_mai_n702_), .C(mai_mai_n698_), .D(mai_mai_n696_), .Y(mai_mai_n710_));
  OR2        m0688(.A(i_11_), .B(i_6_), .Y(mai_mai_n711_));
  NO2        m0689(.A(mai_mai_n701_), .B(mai_mai_n711_), .Y(mai_mai_n712_));
  NA3        m0690(.A(mai_mai_n404_), .B(mai_mai_n597_), .C(mai_mai_n96_), .Y(mai_mai_n713_));
  NA2        m0691(.A(mai_mai_n633_), .B(i_13_), .Y(mai_mai_n714_));
  NAi21      m0692(.An(i_11_), .B(i_12_), .Y(mai_mai_n715_));
  NO3        m0693(.A(mai_mai_n469_), .B(mai_mai_n572_), .C(mai_mai_n598_), .Y(mai_mai_n716_));
  NA2        m0694(.A(mai_mai_n716_), .B(mai_mai_n304_), .Y(mai_mai_n717_));
  NA3        m0695(.A(mai_mai_n717_), .B(mai_mai_n714_), .C(mai_mai_n713_), .Y(mai_mai_n718_));
  OAI210     m0696(.A0(mai_mai_n718_), .A1(mai_mai_n712_), .B0(mai_mai_n63_), .Y(mai_mai_n719_));
  OAI210     m0697(.A0(mai_mai_n233_), .A1(mai_mai_n367_), .B0(mai_mai_n365_), .Y(mai_mai_n720_));
  NO2        m0698(.A(mai_mai_n128_), .B(i_2_), .Y(mai_mai_n721_));
  NA2        m0699(.A(mai_mai_n721_), .B(mai_mai_n626_), .Y(mai_mai_n722_));
  NA2        m0700(.A(mai_mai_n722_), .B(mai_mai_n720_), .Y(mai_mai_n723_));
  NA3        m0701(.A(mai_mai_n723_), .B(mai_mai_n46_), .C(mai_mai_n222_), .Y(mai_mai_n724_));
  NA4        m0702(.A(mai_mai_n724_), .B(mai_mai_n719_), .C(mai_mai_n710_), .D(mai_mai_n694_), .Y(mai_mai_n725_));
  OR4        m0703(.A(mai_mai_n725_), .B(mai_mai_n687_), .C(mai_mai_n671_), .D(mai_mai_n608_), .Y(mai5));
  AOI210     m0704(.A0(mai_mai_n657_), .A1(mai_mai_n262_), .B0(mai_mai_n411_), .Y(mai_mai_n727_));
  NO2        m0705(.A(mai_mai_n594_), .B(i_11_), .Y(mai_mai_n728_));
  OAI210     m0706(.A0(mai_mai_n597_), .A1(mai_mai_n86_), .B0(mai_mai_n728_), .Y(mai_mai_n729_));
  NA2        m0707(.A(mai_mai_n729_), .B(mai_mai_n727_), .Y(mai_mai_n730_));
  NO3        m0708(.A(i_11_), .B(mai_mai_n233_), .C(i_13_), .Y(mai_mai_n731_));
  NO2        m0709(.A(mai_mai_n124_), .B(mai_mai_n23_), .Y(mai_mai_n732_));
  NA2        m0710(.A(i_12_), .B(i_8_), .Y(mai_mai_n733_));
  OAI210     m0711(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n733_), .Y(mai_mai_n734_));
  INV        m0712(.A(mai_mai_n441_), .Y(mai_mai_n735_));
  AOI220     m0713(.A0(mai_mai_n310_), .A1(mai_mai_n565_), .B0(mai_mai_n734_), .B1(mai_mai_n732_), .Y(mai_mai_n736_));
  INV        m0714(.A(mai_mai_n736_), .Y(mai_mai_n737_));
  NO2        m0715(.A(mai_mai_n737_), .B(mai_mai_n730_), .Y(mai_mai_n738_));
  INV        m0716(.A(mai_mai_n170_), .Y(mai_mai_n739_));
  INV        m0717(.A(mai_mai_n241_), .Y(mai_mai_n740_));
  OAI210     m0718(.A0(mai_mai_n683_), .A1(mai_mai_n443_), .B0(mai_mai_n110_), .Y(mai_mai_n741_));
  AOI210     m0719(.A0(mai_mai_n741_), .A1(mai_mai_n740_), .B0(mai_mai_n739_), .Y(mai_mai_n742_));
  NO2        m0720(.A(mai_mai_n450_), .B(mai_mai_n26_), .Y(mai_mai_n743_));
  NO2        m0721(.A(mai_mai_n743_), .B(mai_mai_n413_), .Y(mai_mai_n744_));
  NA2        m0722(.A(mai_mai_n744_), .B(i_2_), .Y(mai_mai_n745_));
  INV        m0723(.A(mai_mai_n745_), .Y(mai_mai_n746_));
  AOI210     m0724(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n410_), .Y(mai_mai_n747_));
  AOI210     m0725(.A0(mai_mai_n747_), .A1(mai_mai_n746_), .B0(mai_mai_n742_), .Y(mai_mai_n748_));
  NO2        m0726(.A(mai_mai_n189_), .B(mai_mai_n125_), .Y(mai_mai_n749_));
  OAI210     m0727(.A0(mai_mai_n749_), .A1(mai_mai_n732_), .B0(i_2_), .Y(mai_mai_n750_));
  NO2        m0728(.A(mai_mai_n750_), .B(mai_mai_n192_), .Y(mai_mai_n751_));
  OA210      m0729(.A0(mai_mai_n611_), .A1(mai_mai_n126_), .B0(i_13_), .Y(mai_mai_n752_));
  NA2        m0730(.A(mai_mai_n198_), .B(mai_mai_n201_), .Y(mai_mai_n753_));
  NA2        m0731(.A(mai_mai_n151_), .B(mai_mai_n589_), .Y(mai_mai_n754_));
  AOI210     m0732(.A0(mai_mai_n754_), .A1(mai_mai_n753_), .B0(mai_mai_n368_), .Y(mai_mai_n755_));
  AOI210     m0733(.A0(mai_mai_n206_), .A1(mai_mai_n148_), .B0(mai_mai_n507_), .Y(mai_mai_n756_));
  OAI210     m0734(.A0(mai_mai_n756_), .A1(mai_mai_n223_), .B0(mai_mai_n413_), .Y(mai_mai_n757_));
  NO2        m0735(.A(mai_mai_n101_), .B(mai_mai_n45_), .Y(mai_mai_n758_));
  INV        m0736(.A(mai_mai_n294_), .Y(mai_mai_n759_));
  NA4        m0737(.A(mai_mai_n759_), .B(mai_mai_n297_), .C(mai_mai_n124_), .D(mai_mai_n43_), .Y(mai_mai_n760_));
  OAI210     m0738(.A0(mai_mai_n760_), .A1(mai_mai_n758_), .B0(mai_mai_n757_), .Y(mai_mai_n761_));
  NO4        m0739(.A(mai_mai_n761_), .B(mai_mai_n755_), .C(mai_mai_n752_), .D(mai_mai_n751_), .Y(mai_mai_n762_));
  NA2        m0740(.A(mai_mai_n565_), .B(mai_mai_n28_), .Y(mai_mai_n763_));
  NA2        m0741(.A(mai_mai_n731_), .B(mai_mai_n268_), .Y(mai_mai_n764_));
  NA2        m0742(.A(mai_mai_n764_), .B(mai_mai_n763_), .Y(mai_mai_n765_));
  NO2        m0743(.A(mai_mai_n62_), .B(i_12_), .Y(mai_mai_n766_));
  NO2        m0744(.A(mai_mai_n766_), .B(mai_mai_n126_), .Y(mai_mai_n767_));
  NO2        m0745(.A(mai_mai_n767_), .B(mai_mai_n589_), .Y(mai_mai_n768_));
  AOI220     m0746(.A0(mai_mai_n768_), .A1(mai_mai_n36_), .B0(mai_mai_n765_), .B1(mai_mai_n47_), .Y(mai_mai_n769_));
  NA4        m0747(.A(mai_mai_n769_), .B(mai_mai_n762_), .C(mai_mai_n748_), .D(mai_mai_n738_), .Y(mai6));
  NO3        m0748(.A(mai_mai_n250_), .B(mai_mai_n299_), .C(i_1_), .Y(mai_mai_n771_));
  NO2        m0749(.A(mai_mai_n184_), .B(mai_mai_n139_), .Y(mai_mai_n772_));
  OAI210     m0750(.A0(mai_mai_n772_), .A1(mai_mai_n771_), .B0(mai_mai_n721_), .Y(mai_mai_n773_));
  NA4        m0751(.A(mai_mai_n385_), .B(mai_mai_n474_), .C(mai_mai_n69_), .D(mai_mai_n100_), .Y(mai_mai_n774_));
  INV        m0752(.A(mai_mai_n774_), .Y(mai_mai_n775_));
  NO2        m0753(.A(mai_mai_n218_), .B(mai_mai_n478_), .Y(mai_mai_n776_));
  NO2        m0754(.A(i_11_), .B(i_9_), .Y(mai_mai_n777_));
  NO3        m0755(.A(mai_mai_n776_), .B(mai_mai_n775_), .C(mai_mai_n322_), .Y(mai_mai_n778_));
  AO210      m0756(.A0(mai_mai_n778_), .A1(mai_mai_n773_), .B0(i_12_), .Y(mai_mai_n779_));
  NA2        m0757(.A(mai_mai_n369_), .B(mai_mai_n328_), .Y(mai_mai_n780_));
  NA2        m0758(.A(mai_mai_n572_), .B(mai_mai_n63_), .Y(mai_mai_n781_));
  NA2        m0759(.A(mai_mai_n673_), .B(mai_mai_n69_), .Y(mai_mai_n782_));
  NA4        m0760(.A(mai_mai_n616_), .B(mai_mai_n782_), .C(mai_mai_n781_), .D(mai_mai_n780_), .Y(mai_mai_n783_));
  INV        m0761(.A(mai_mai_n195_), .Y(mai_mai_n784_));
  AOI220     m0762(.A0(mai_mai_n784_), .A1(mai_mai_n777_), .B0(mai_mai_n783_), .B1(mai_mai_n71_), .Y(mai_mai_n785_));
  NO2        m0763(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n786_));
  NA3        m0764(.A(mai_mai_n786_), .B(mai_mai_n465_), .C(mai_mai_n385_), .Y(mai_mai_n787_));
  NAi32      m0765(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n788_));
  AOI210     m0766(.A0(mai_mai_n711_), .A1(mai_mai_n84_), .B0(mai_mai_n788_), .Y(mai_mai_n789_));
  OAI210     m0767(.A0(mai_mai_n672_), .A1(mai_mai_n553_), .B0(mai_mai_n552_), .Y(mai_mai_n790_));
  NAi31      m0768(.An(mai_mai_n789_), .B(mai_mai_n790_), .C(mai_mai_n787_), .Y(mai_mai_n791_));
  NO2        m0769(.A(mai_mai_n688_), .B(i_2_), .Y(mai_mai_n792_));
  NA2        m0770(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n793_));
  OAI210     m0771(.A0(mai_mai_n793_), .A1(mai_mai_n403_), .B0(mai_mai_n355_), .Y(mai_mai_n794_));
  NA2        m0772(.A(mai_mai_n794_), .B(mai_mai_n792_), .Y(mai_mai_n795_));
  AO220      m0773(.A0(mai_mai_n354_), .A1(mai_mai_n344_), .B0(mai_mai_n392_), .B1(mai_mai_n589_), .Y(mai_mai_n796_));
  NA3        m0774(.A(mai_mai_n796_), .B(mai_mai_n251_), .C(i_7_), .Y(mai_mai_n797_));
  NA3        m0775(.A(mai_mai_n443_), .B(mai_mai_n147_), .C(mai_mai_n67_), .Y(mai_mai_n798_));
  AO210      m0776(.A0(mai_mai_n482_), .A1(mai_mai_n735_), .B0(mai_mai_n36_), .Y(mai_mai_n799_));
  NA4        m0777(.A(mai_mai_n799_), .B(mai_mai_n798_), .C(mai_mai_n797_), .D(mai_mai_n795_), .Y(mai_mai_n800_));
  OAI210     m0778(.A0(mai_mai_n632_), .A1(i_11_), .B0(mai_mai_n84_), .Y(mai_mai_n801_));
  AOI220     m0779(.A0(mai_mai_n801_), .A1(mai_mai_n552_), .B0(mai_mai_n776_), .B1(mai_mai_n705_), .Y(mai_mai_n802_));
  NA3        m0780(.A(mai_mai_n368_), .B(mai_mai_n234_), .C(mai_mai_n147_), .Y(mai_mai_n803_));
  NA2        m0781(.A(mai_mai_n392_), .B(mai_mai_n68_), .Y(mai_mai_n804_));
  NA4        m0782(.A(mai_mai_n804_), .B(mai_mai_n803_), .C(mai_mai_n802_), .D(mai_mai_n596_), .Y(mai_mai_n805_));
  AO210      m0783(.A0(mai_mai_n507_), .A1(mai_mai_n47_), .B0(mai_mai_n85_), .Y(mai_mai_n806_));
  NA3        m0784(.A(mai_mai_n806_), .B(mai_mai_n475_), .C(mai_mai_n216_), .Y(mai_mai_n807_));
  AOI210     m0785(.A0(mai_mai_n443_), .A1(mai_mai_n441_), .B0(mai_mai_n551_), .Y(mai_mai_n808_));
  NO2        m0786(.A(mai_mai_n601_), .B(mai_mai_n101_), .Y(mai_mai_n809_));
  OAI210     m0787(.A0(mai_mai_n809_), .A1(mai_mai_n111_), .B0(mai_mai_n402_), .Y(mai_mai_n810_));
  NA2        m0788(.A(mai_mai_n240_), .B(mai_mai_n47_), .Y(mai_mai_n811_));
  NA2        m0789(.A(mai_mai_n811_), .B(mai_mai_n578_), .Y(mai_mai_n812_));
  NA3        m0790(.A(mai_mai_n812_), .B(mai_mai_n321_), .C(i_7_), .Y(mai_mai_n813_));
  NA4        m0791(.A(mai_mai_n813_), .B(mai_mai_n810_), .C(mai_mai_n808_), .D(mai_mai_n807_), .Y(mai_mai_n814_));
  NO4        m0792(.A(mai_mai_n814_), .B(mai_mai_n805_), .C(mai_mai_n800_), .D(mai_mai_n791_), .Y(mai_mai_n815_));
  NA4        m0793(.A(mai_mai_n815_), .B(mai_mai_n785_), .C(mai_mai_n779_), .D(mai_mai_n375_), .Y(mai3));
  NA2        m0794(.A(i_6_), .B(i_7_), .Y(mai_mai_n817_));
  NO2        m0795(.A(mai_mai_n817_), .B(i_0_), .Y(mai_mai_n818_));
  NO2        m0796(.A(i_11_), .B(mai_mai_n233_), .Y(mai_mai_n819_));
  OAI210     m0797(.A0(mai_mai_n818_), .A1(mai_mai_n282_), .B0(mai_mai_n819_), .Y(mai_mai_n820_));
  NO2        m0798(.A(mai_mai_n820_), .B(mai_mai_n192_), .Y(mai_mai_n821_));
  NO3        m0799(.A(mai_mai_n446_), .B(mai_mai_n88_), .C(mai_mai_n45_), .Y(mai_mai_n822_));
  OA210      m0800(.A0(mai_mai_n822_), .A1(mai_mai_n821_), .B0(mai_mai_n173_), .Y(mai_mai_n823_));
  INV        m0801(.A(mai_mai_n803_), .Y(mai_mai_n824_));
  NA2        m0802(.A(mai_mai_n824_), .B(mai_mai_n40_), .Y(mai_mai_n825_));
  NO3        m0803(.A(mai_mai_n621_), .B(mai_mai_n450_), .C(mai_mai_n131_), .Y(mai_mai_n826_));
  NA2        m0804(.A(mai_mai_n404_), .B(mai_mai_n46_), .Y(mai_mai_n827_));
  AN2        m0805(.A(mai_mai_n448_), .B(mai_mai_n55_), .Y(mai_mai_n828_));
  NO2        m0806(.A(mai_mai_n828_), .B(mai_mai_n826_), .Y(mai_mai_n829_));
  AOI210     m0807(.A0(mai_mai_n829_), .A1(mai_mai_n825_), .B0(mai_mai_n49_), .Y(mai_mai_n830_));
  NO4        m0808(.A(mai_mai_n372_), .B(mai_mai_n378_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n831_));
  NA2        m0809(.A(mai_mai_n184_), .B(mai_mai_n561_), .Y(mai_mai_n832_));
  NA2        m0810(.A(mai_mai_n697_), .B(mai_mai_n665_), .Y(mai_mai_n833_));
  NA2        m0811(.A(i_0_), .B(mai_mai_n433_), .Y(mai_mai_n834_));
  OAI220     m0812(.A0(mai_mai_n834_), .A1(mai_mai_n833_), .B0(mai_mai_n1032_), .B1(mai_mai_n63_), .Y(mai_mai_n835_));
  NOi21      m0813(.An(i_5_), .B(i_9_), .Y(mai_mai_n836_));
  NA2        m0814(.A(mai_mai_n836_), .B(mai_mai_n440_), .Y(mai_mai_n837_));
  INV        m0815(.A(mai_mai_n677_), .Y(mai_mai_n838_));
  NO3        m0816(.A(mai_mai_n407_), .B(mai_mai_n259_), .C(mai_mai_n71_), .Y(mai_mai_n839_));
  NO2        m0817(.A(mai_mai_n174_), .B(mai_mai_n148_), .Y(mai_mai_n840_));
  AOI210     m0818(.A0(mai_mai_n840_), .A1(mai_mai_n240_), .B0(mai_mai_n839_), .Y(mai_mai_n841_));
  OAI220     m0819(.A0(mai_mai_n841_), .A1(mai_mai_n180_), .B0(mai_mai_n838_), .B1(mai_mai_n837_), .Y(mai_mai_n842_));
  NO4        m0820(.A(mai_mai_n842_), .B(mai_mai_n835_), .C(mai_mai_n830_), .D(mai_mai_n823_), .Y(mai_mai_n843_));
  NOi21      m0821(.An(i_0_), .B(i_10_), .Y(mai_mai_n844_));
  NA2        m0822(.A(mai_mai_n184_), .B(mai_mai_n24_), .Y(mai_mai_n845_));
  NO2        m0823(.A(mai_mai_n664_), .B(mai_mai_n586_), .Y(mai_mai_n846_));
  NO2        m0824(.A(mai_mai_n846_), .B(mai_mai_n845_), .Y(mai_mai_n847_));
  NA2        m0825(.A(mai_mai_n304_), .B(mai_mai_n129_), .Y(mai_mai_n848_));
  NAi21      m0826(.An(mai_mai_n161_), .B(mai_mai_n433_), .Y(mai_mai_n849_));
  OAI220     m0827(.A0(mai_mai_n849_), .A1(mai_mai_n811_), .B0(mai_mai_n848_), .B1(mai_mai_n396_), .Y(mai_mai_n850_));
  NO2        m0828(.A(mai_mai_n850_), .B(mai_mai_n847_), .Y(mai_mai_n851_));
  NO2        m0829(.A(mai_mai_n385_), .B(mai_mai_n286_), .Y(mai_mai_n852_));
  NA2        m0830(.A(mai_mai_n852_), .B(mai_mai_n700_), .Y(mai_mai_n853_));
  NA2        m0831(.A(mai_mai_n562_), .B(i_0_), .Y(mai_mai_n854_));
  NO3        m0832(.A(mai_mai_n854_), .B(mai_mai_n380_), .C(mai_mai_n86_), .Y(mai_mai_n855_));
  NO4        m0833(.A(mai_mai_n577_), .B(mai_mai_n213_), .C(mai_mai_n410_), .D(mai_mai_n403_), .Y(mai_mai_n856_));
  AOI210     m0834(.A0(mai_mai_n856_), .A1(i_11_), .B0(mai_mai_n855_), .Y(mai_mai_n857_));
  AN2        m0835(.A(mai_mai_n95_), .B(mai_mai_n239_), .Y(mai_mai_n858_));
  NA2        m0836(.A(mai_mai_n731_), .B(mai_mai_n322_), .Y(mai_mai_n859_));
  AOI210     m0837(.A0(mai_mai_n475_), .A1(mai_mai_n86_), .B0(mai_mai_n58_), .Y(mai_mai_n860_));
  OAI220     m0838(.A0(mai_mai_n860_), .A1(mai_mai_n859_), .B0(mai_mai_n652_), .B1(mai_mai_n524_), .Y(mai_mai_n861_));
  INV        m0839(.A(mai_mai_n526_), .Y(mai_mai_n862_));
  NO4        m0840(.A(mai_mai_n114_), .B(mai_mai_n58_), .C(mai_mai_n661_), .D(i_5_), .Y(mai_mai_n863_));
  AN2        m0841(.A(mai_mai_n863_), .B(mai_mai_n862_), .Y(mai_mai_n864_));
  AOI210     m0842(.A0(i_0_), .A1(mai_mai_n97_), .B0(mai_mai_n184_), .Y(mai_mai_n865_));
  NA2        m0843(.A(mai_mai_n556_), .B(i_4_), .Y(mai_mai_n866_));
  NA2        m0844(.A(mai_mai_n187_), .B(mai_mai_n201_), .Y(mai_mai_n867_));
  OAI220     m0845(.A0(mai_mai_n867_), .A1(mai_mai_n859_), .B0(mai_mai_n866_), .B1(mai_mai_n865_), .Y(mai_mai_n868_));
  NO4        m0846(.A(mai_mai_n868_), .B(mai_mai_n864_), .C(mai_mai_n861_), .D(mai_mai_n858_), .Y(mai_mai_n869_));
  NA4        m0847(.A(mai_mai_n869_), .B(mai_mai_n857_), .C(mai_mai_n853_), .D(mai_mai_n851_), .Y(mai_mai_n870_));
  NO2        m0848(.A(mai_mai_n102_), .B(mai_mai_n37_), .Y(mai_mai_n871_));
  NA2        m0849(.A(i_11_), .B(i_9_), .Y(mai_mai_n872_));
  NO3        m0850(.A(i_12_), .B(mai_mai_n872_), .C(mai_mai_n595_), .Y(mai_mai_n873_));
  AO220      m0851(.A0(mai_mai_n873_), .A1(mai_mai_n871_), .B0(mai_mai_n261_), .B1(mai_mai_n85_), .Y(mai_mai_n874_));
  NA2        m0852(.A(mai_mai_n389_), .B(mai_mai_n178_), .Y(mai_mai_n875_));
  NAi31      m0853(.An(mai_mai_n256_), .B(mai_mai_n875_), .C(mai_mai_n159_), .Y(mai_mai_n876_));
  NO2        m0854(.A(mai_mai_n872_), .B(mai_mai_n71_), .Y(mai_mai_n877_));
  NO2        m0855(.A(mai_mai_n174_), .B(i_0_), .Y(mai_mai_n878_));
  INV        m0856(.A(mai_mai_n878_), .Y(mai_mai_n879_));
  NA2        m0857(.A(mai_mai_n465_), .B(mai_mai_n228_), .Y(mai_mai_n880_));
  OAI220     m0858(.A0(i_12_), .A1(mai_mai_n837_), .B0(mai_mai_n880_), .B1(mai_mai_n879_), .Y(mai_mai_n881_));
  NO3        m0859(.A(mai_mai_n881_), .B(mai_mai_n876_), .C(mai_mai_n874_), .Y(mai_mai_n882_));
  NA2        m0860(.A(mai_mai_n651_), .B(mai_mai_n121_), .Y(mai_mai_n883_));
  NO2        m0861(.A(i_6_), .B(mai_mai_n883_), .Y(mai_mai_n884_));
  AOI210     m0862(.A0(mai_mai_n442_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n885_));
  NA2        m0863(.A(mai_mai_n170_), .B(mai_mai_n102_), .Y(mai_mai_n886_));
  NOi32      m0864(.An(mai_mai_n885_), .Bn(mai_mai_n187_), .C(mai_mai_n886_), .Y(mai_mai_n887_));
  AOI210     m0865(.A0(mai_mai_n597_), .A1(mai_mai_n322_), .B0(mai_mai_n239_), .Y(mai_mai_n888_));
  NO2        m0866(.A(mai_mai_n888_), .B(mai_mai_n827_), .Y(mai_mai_n889_));
  NO3        m0867(.A(mai_mai_n889_), .B(mai_mai_n887_), .C(mai_mai_n884_), .Y(mai_mai_n890_));
  NOi21      m0868(.An(i_7_), .B(i_5_), .Y(mai_mai_n891_));
  NOi31      m0869(.An(mai_mai_n891_), .B(mai_mai_n844_), .C(mai_mai_n715_), .Y(mai_mai_n892_));
  NA3        m0870(.A(mai_mai_n892_), .B(mai_mai_n379_), .C(i_6_), .Y(mai_mai_n893_));
  OA210      m0871(.A0(mai_mai_n886_), .A1(mai_mai_n506_), .B0(mai_mai_n893_), .Y(mai_mai_n894_));
  NO3        m0872(.A(mai_mai_n398_), .B(mai_mai_n357_), .C(mai_mai_n353_), .Y(mai_mai_n895_));
  NO2        m0873(.A(mai_mai_n253_), .B(mai_mai_n311_), .Y(mai_mai_n896_));
  INV        m0874(.A(mai_mai_n715_), .Y(mai_mai_n897_));
  AOI210     m0875(.A0(mai_mai_n897_), .A1(mai_mai_n896_), .B0(mai_mai_n895_), .Y(mai_mai_n898_));
  NA4        m0876(.A(mai_mai_n898_), .B(mai_mai_n894_), .C(mai_mai_n890_), .D(mai_mai_n882_), .Y(mai_mai_n899_));
  AN2        m0877(.A(mai_mai_n326_), .B(mai_mai_n322_), .Y(mai_mai_n900_));
  AO220      m0878(.A0(mai_mai_n900_), .A1(mai_mai_n840_), .B0(mai_mai_n339_), .B1(mai_mai_n27_), .Y(mai_mai_n901_));
  NA2        m0879(.A(mai_mai_n901_), .B(i_10_), .Y(mai_mai_n902_));
  OA210      m0880(.A0(mai_mai_n465_), .A1(mai_mai_n220_), .B0(mai_mai_n464_), .Y(mai_mai_n903_));
  NA3        m0881(.A(mai_mai_n464_), .B(mai_mai_n404_), .C(mai_mai_n46_), .Y(mai_mai_n904_));
  OAI210     m0882(.A0(mai_mai_n849_), .A1(i_6_), .B0(mai_mai_n904_), .Y(mai_mai_n905_));
  NA2        m0883(.A(mai_mai_n877_), .B(mai_mai_n297_), .Y(mai_mai_n906_));
  NA2        m0884(.A(mai_mai_n186_), .B(mai_mai_n906_), .Y(mai_mai_n907_));
  AOI220     m0885(.A0(mai_mai_n907_), .A1(mai_mai_n465_), .B0(mai_mai_n905_), .B1(mai_mai_n71_), .Y(mai_mai_n908_));
  NA3        m0886(.A(mai_mai_n793_), .B(mai_mai_n377_), .C(mai_mai_n632_), .Y(mai_mai_n909_));
  NO2        m0887(.A(mai_mai_n73_), .B(mai_mai_n733_), .Y(mai_mai_n910_));
  AOI210     m0888(.A0(mai_mai_n173_), .A1(mai_mai_n586_), .B0(mai_mai_n910_), .Y(mai_mai_n911_));
  AOI210     m0889(.A0(mai_mai_n911_), .A1(mai_mai_n909_), .B0(mai_mai_n48_), .Y(mai_mai_n912_));
  NO3        m0890(.A(mai_mai_n577_), .B(mai_mai_n352_), .C(mai_mai_n24_), .Y(mai_mai_n913_));
  NO2        m0891(.A(mai_mai_n534_), .B(mai_mai_n913_), .Y(mai_mai_n914_));
  NAi21      m0892(.An(i_9_), .B(i_5_), .Y(mai_mai_n915_));
  NO2        m0893(.A(mai_mai_n915_), .B(mai_mai_n398_), .Y(mai_mai_n916_));
  NO2        m0894(.A(mai_mai_n592_), .B(mai_mai_n104_), .Y(mai_mai_n917_));
  AOI220     m0895(.A0(mai_mai_n917_), .A1(i_0_), .B0(mai_mai_n916_), .B1(mai_mai_n611_), .Y(mai_mai_n918_));
  OAI220     m0896(.A0(mai_mai_n918_), .A1(mai_mai_n83_), .B0(mai_mai_n914_), .B1(mai_mai_n171_), .Y(mai_mai_n919_));
  NO2        m0897(.A(mai_mai_n919_), .B(mai_mai_n912_), .Y(mai_mai_n920_));
  NA3        m0898(.A(mai_mai_n920_), .B(mai_mai_n908_), .C(mai_mai_n902_), .Y(mai_mai_n921_));
  NO3        m0899(.A(mai_mai_n921_), .B(mai_mai_n899_), .C(mai_mai_n870_), .Y(mai_mai_n922_));
  NO2        m0900(.A(mai_mai_n844_), .B(mai_mai_n715_), .Y(mai_mai_n923_));
  NA2        m0901(.A(mai_mai_n71_), .B(mai_mai_n45_), .Y(mai_mai_n924_));
  INV        m0902(.A(mai_mai_n924_), .Y(mai_mai_n925_));
  NO3        m0903(.A(mai_mai_n104_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n926_));
  AO220      m0904(.A0(mai_mai_n926_), .A1(mai_mai_n925_), .B0(mai_mai_n923_), .B1(mai_mai_n173_), .Y(mai_mai_n927_));
  AOI210     m0905(.A0(mai_mai_n781_), .A1(mai_mai_n675_), .B0(mai_mai_n886_), .Y(mai_mai_n928_));
  AOI210     m0906(.A0(mai_mai_n927_), .A1(mai_mai_n341_), .B0(mai_mai_n928_), .Y(mai_mai_n929_));
  NA3        m0907(.A(mai_mai_n146_), .B(mai_mai_n665_), .C(mai_mai_n71_), .Y(mai_mai_n930_));
  NO2        m0908(.A(mai_mai_n790_), .B(mai_mai_n398_), .Y(mai_mai_n931_));
  NA3        m0909(.A(mai_mai_n818_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n932_));
  NA2        m0910(.A(mai_mai_n819_), .B(i_9_), .Y(mai_mai_n933_));
  AOI210     m0911(.A0(mai_mai_n932_), .A1(mai_mai_n487_), .B0(mai_mai_n933_), .Y(mai_mai_n934_));
  OAI210     m0912(.A0(mai_mai_n240_), .A1(i_9_), .B0(mai_mai_n227_), .Y(mai_mai_n935_));
  AOI210     m0913(.A0(mai_mai_n935_), .A1(mai_mai_n854_), .B0(mai_mai_n152_), .Y(mai_mai_n936_));
  NO3        m0914(.A(mai_mai_n936_), .B(mai_mai_n934_), .C(mai_mai_n931_), .Y(mai_mai_n937_));
  NA3        m0915(.A(mai_mai_n937_), .B(mai_mai_n930_), .C(mai_mai_n929_), .Y(mai_mai_n938_));
  NA2        m0916(.A(mai_mai_n900_), .B(mai_mai_n368_), .Y(mai_mai_n939_));
  AOI210     m0917(.A0(mai_mai_n293_), .A1(mai_mai_n161_), .B0(mai_mai_n939_), .Y(mai_mai_n940_));
  NA3        m0918(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n941_));
  NA2        m0919(.A(i_5_), .B(mai_mai_n479_), .Y(mai_mai_n942_));
  AOI210     m0920(.A0(mai_mai_n941_), .A1(mai_mai_n161_), .B0(mai_mai_n942_), .Y(mai_mai_n943_));
  NO2        m0921(.A(mai_mai_n943_), .B(mai_mai_n940_), .Y(mai_mai_n944_));
  NO3        m0922(.A(mai_mai_n207_), .B(mai_mai_n378_), .C(i_0_), .Y(mai_mai_n945_));
  OAI210     m0923(.A0(mai_mai_n945_), .A1(mai_mai_n74_), .B0(i_13_), .Y(mai_mai_n946_));
  INV        m0924(.A(mai_mai_n216_), .Y(mai_mai_n947_));
  OAI220     m0925(.A0(mai_mai_n518_), .A1(mai_mai_n139_), .B0(i_12_), .B1(mai_mai_n605_), .Y(mai_mai_n948_));
  NA3        m0926(.A(mai_mai_n948_), .B(i_7_), .C(mai_mai_n947_), .Y(mai_mai_n949_));
  NA3        m0927(.A(mai_mai_n949_), .B(mai_mai_n946_), .C(mai_mai_n944_), .Y(mai_mai_n950_));
  NO2        m0928(.A(mai_mai_n238_), .B(mai_mai_n91_), .Y(mai_mai_n951_));
  AOI210     m0929(.A0(mai_mai_n951_), .A1(mai_mai_n923_), .B0(mai_mai_n108_), .Y(mai_mai_n952_));
  AOI220     m0930(.A0(mai_mai_n891_), .A1(mai_mai_n479_), .B0(mai_mai_n818_), .B1(mai_mai_n162_), .Y(mai_mai_n953_));
  NA2        m0931(.A(mai_mai_n344_), .B(mai_mai_n175_), .Y(mai_mai_n954_));
  OA220      m0932(.A0(mai_mai_n954_), .A1(mai_mai_n953_), .B0(mai_mai_n952_), .B1(i_5_), .Y(mai_mai_n955_));
  AOI210     m0933(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n174_), .Y(mai_mai_n956_));
  NA2        m0934(.A(mai_mai_n956_), .B(mai_mai_n903_), .Y(mai_mai_n957_));
  NA3        m0935(.A(mai_mai_n602_), .B(mai_mai_n184_), .C(mai_mai_n82_), .Y(mai_mai_n958_));
  NA2        m0936(.A(mai_mai_n958_), .B(mai_mai_n533_), .Y(mai_mai_n959_));
  NA2        m0937(.A(mai_mai_n481_), .B(mai_mai_n462_), .Y(mai_mai_n960_));
  NO2        m0938(.A(mai_mai_n960_), .B(mai_mai_n959_), .Y(mai_mai_n961_));
  NA3        m0939(.A(i_5_), .B(mai_mai_n282_), .C(mai_mai_n227_), .Y(mai_mai_n962_));
  INV        m0940(.A(mai_mai_n962_), .Y(mai_mai_n963_));
  NA3        m0941(.A(mai_mai_n385_), .B(mai_mai_n327_), .C(mai_mai_n219_), .Y(mai_mai_n964_));
  OAI210     m0942(.A0(mai_mai_n832_), .A1(mai_mai_n639_), .B0(mai_mai_n964_), .Y(mai_mai_n965_));
  NOi31      m0943(.An(mai_mai_n384_), .B(mai_mai_n924_), .C(mai_mai_n235_), .Y(mai_mai_n966_));
  NO3        m0944(.A(mai_mai_n966_), .B(mai_mai_n965_), .C(mai_mai_n963_), .Y(mai_mai_n967_));
  NA4        m0945(.A(mai_mai_n967_), .B(mai_mai_n961_), .C(mai_mai_n957_), .D(mai_mai_n955_), .Y(mai_mai_n968_));
  INV        m0946(.A(mai_mai_n604_), .Y(mai_mai_n969_));
  NO3        m0947(.A(mai_mai_n969_), .B(mai_mai_n547_), .C(i_7_), .Y(mai_mai_n970_));
  INV        m0948(.A(mai_mai_n970_), .Y(mai_mai_n971_));
  NA3        m0949(.A(mai_mai_n297_), .B(i_5_), .C(mai_mai_n192_), .Y(mai_mai_n972_));
  NO4        m0950(.A(mai_mai_n235_), .B(mai_mai_n207_), .C(i_0_), .D(i_12_), .Y(mai_mai_n973_));
  AOI220     m0951(.A0(mai_mai_n973_), .A1(mai_mai_n297_), .B0(mai_mai_n775_), .B1(mai_mai_n175_), .Y(mai_mai_n974_));
  BUFFER     m0952(.A(mai_mai_n152_), .Y(mai_mai_n975_));
  NO4        m0953(.A(mai_mai_n975_), .B(i_12_), .C(mai_mai_n639_), .D(mai_mai_n131_), .Y(mai_mai_n976_));
  NA2        m0954(.A(mai_mai_n976_), .B(mai_mai_n216_), .Y(mai_mai_n977_));
  NA3        m0955(.A(mai_mai_n97_), .B(mai_mai_n561_), .C(i_11_), .Y(mai_mai_n978_));
  NO2        m0956(.A(mai_mai_n978_), .B(mai_mai_n154_), .Y(mai_mai_n979_));
  NA2        m0957(.A(mai_mai_n891_), .B(mai_mai_n461_), .Y(mai_mai_n980_));
  OAI210     m0958(.A0(i_7_), .A1(mai_mai_n972_), .B0(mai_mai_n980_), .Y(mai_mai_n981_));
  AOI210     m0959(.A0(mai_mai_n981_), .A1(mai_mai_n878_), .B0(mai_mai_n979_), .Y(mai_mai_n982_));
  NA4        m0960(.A(mai_mai_n982_), .B(mai_mai_n977_), .C(mai_mai_n974_), .D(mai_mai_n971_), .Y(mai_mai_n983_));
  NO4        m0961(.A(mai_mai_n983_), .B(mai_mai_n968_), .C(mai_mai_n950_), .D(mai_mai_n938_), .Y(mai_mai_n984_));
  OAI210     m0962(.A0(mai_mai_n792_), .A1(mai_mai_n786_), .B0(mai_mai_n37_), .Y(mai_mai_n985_));
  NA3        m0963(.A(mai_mai_n885_), .B(mai_mai_n365_), .C(i_5_), .Y(mai_mai_n986_));
  NA3        m0964(.A(mai_mai_n986_), .B(mai_mai_n985_), .C(mai_mai_n600_), .Y(mai_mai_n987_));
  NA2        m0965(.A(mai_mai_n987_), .B(mai_mai_n204_), .Y(mai_mai_n988_));
  NA2        m0966(.A(mai_mai_n185_), .B(mai_mai_n187_), .Y(mai_mai_n989_));
  AO210      m0967(.A0(i_11_), .A1(mai_mai_n33_), .B0(mai_mai_n989_), .Y(mai_mai_n990_));
  OAI210     m0968(.A0(mai_mai_n604_), .A1(mai_mai_n602_), .B0(mai_mai_n310_), .Y(mai_mai_n991_));
  NAi31      m0969(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n992_));
  AOI210     m0970(.A0(mai_mai_n117_), .A1(mai_mai_n68_), .B0(mai_mai_n992_), .Y(mai_mai_n993_));
  NO2        m0971(.A(mai_mai_n993_), .B(mai_mai_n637_), .Y(mai_mai_n994_));
  NA3        m0972(.A(mai_mai_n994_), .B(mai_mai_n991_), .C(mai_mai_n990_), .Y(mai_mai_n995_));
  NO2        m0973(.A(mai_mai_n453_), .B(mai_mai_n259_), .Y(mai_mai_n996_));
  NO2        m0974(.A(mai_mai_n996_), .B(mai_mai_n856_), .Y(mai_mai_n997_));
  OAI210     m0975(.A0(mai_mai_n978_), .A1(mai_mai_n148_), .B0(mai_mai_n997_), .Y(mai_mai_n998_));
  AOI210     m0976(.A0(mai_mai_n995_), .A1(mai_mai_n49_), .B0(mai_mai_n998_), .Y(mai_mai_n999_));
  AOI210     m0977(.A0(mai_mai_n999_), .A1(mai_mai_n988_), .B0(mai_mai_n71_), .Y(mai_mai_n1000_));
  NO2        m0978(.A(mai_mai_n554_), .B(mai_mai_n374_), .Y(mai_mai_n1001_));
  NO2        m0979(.A(mai_mai_n1001_), .B(mai_mai_n739_), .Y(mai_mai_n1002_));
  NA2        m0980(.A(i_5_), .B(mai_mai_n74_), .Y(mai_mai_n1003_));
  AOI210     m0981(.A0(mai_mai_n956_), .A1(i_5_), .B0(mai_mai_n892_), .Y(mai_mai_n1004_));
  AOI210     m0982(.A0(mai_mai_n1004_), .A1(mai_mai_n1003_), .B0(mai_mai_n666_), .Y(mai_mai_n1005_));
  NA2        m0983(.A(mai_mai_n253_), .B(mai_mai_n57_), .Y(mai_mai_n1006_));
  AOI220     m0984(.A0(mai_mai_n1006_), .A1(mai_mai_n74_), .B0(mai_mai_n339_), .B1(mai_mai_n250_), .Y(mai_mai_n1007_));
  NO2        m0985(.A(mai_mai_n1007_), .B(mai_mai_n233_), .Y(mai_mai_n1008_));
  NO2        m0986(.A(mai_mai_n1008_), .B(mai_mai_n1005_), .Y(mai_mai_n1009_));
  OAI210     m0987(.A0(mai_mai_n261_), .A1(mai_mai_n157_), .B0(mai_mai_n86_), .Y(mai_mai_n1010_));
  NA3        m0988(.A(mai_mai_n743_), .B(mai_mai_n282_), .C(mai_mai_n78_), .Y(mai_mai_n1011_));
  AOI210     m0989(.A0(mai_mai_n1011_), .A1(mai_mai_n1010_), .B0(i_11_), .Y(mai_mai_n1012_));
  OAI210     m0990(.A0(mai_mai_n1031_), .A1(mai_mai_n885_), .B0(mai_mai_n204_), .Y(mai_mai_n1013_));
  NA2        m0991(.A(mai_mai_n163_), .B(i_5_), .Y(mai_mai_n1014_));
  AOI210     m0992(.A0(mai_mai_n1013_), .A1(mai_mai_n753_), .B0(mai_mai_n1014_), .Y(mai_mai_n1015_));
  NO3        m0993(.A(mai_mai_n59_), .B(mai_mai_n58_), .C(i_4_), .Y(mai_mai_n1016_));
  OAI210     m0994(.A0(mai_mai_n896_), .A1(mai_mai_n299_), .B0(mai_mai_n1016_), .Y(mai_mai_n1017_));
  NO2        m0995(.A(mai_mai_n1017_), .B(mai_mai_n715_), .Y(mai_mai_n1018_));
  NO4        m0996(.A(mai_mai_n915_), .B(mai_mai_n468_), .C(mai_mai_n249_), .D(mai_mai_n248_), .Y(mai_mai_n1019_));
  NO2        m0997(.A(mai_mai_n1019_), .B(mai_mai_n551_), .Y(mai_mai_n1020_));
  NO2        m0998(.A(mai_mai_n789_), .B(mai_mai_n358_), .Y(mai_mai_n1021_));
  AOI210     m0999(.A0(mai_mai_n1021_), .A1(mai_mai_n1020_), .B0(mai_mai_n41_), .Y(mai_mai_n1022_));
  NO4        m1000(.A(mai_mai_n1022_), .B(mai_mai_n1018_), .C(mai_mai_n1015_), .D(mai_mai_n1012_), .Y(mai_mai_n1023_));
  OAI210     m1001(.A0(mai_mai_n1009_), .A1(i_4_), .B0(mai_mai_n1023_), .Y(mai_mai_n1024_));
  NO3        m1002(.A(mai_mai_n1024_), .B(mai_mai_n1002_), .C(mai_mai_n1000_), .Y(mai_mai_n1025_));
  NA4        m1003(.A(mai_mai_n1025_), .B(mai_mai_n984_), .C(mai_mai_n922_), .D(mai_mai_n843_), .Y(mai4));
  INV        m1004(.A(i_2_), .Y(mai_mai_n1029_));
  INV        m1005(.A(i_5_), .Y(mai_mai_n1030_));
  INV        m1006(.A(i_12_), .Y(mai_mai_n1031_));
  INV        m1007(.A(mai_mai_n831_), .Y(mai_mai_n1032_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u0016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u0017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u0018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_5_), .A1(men_men_n47_), .B0(men_men_n46_), .Y(men_men_n51_));
  NA2        u0029(.A(i_0_), .B(i_2_), .Y(men_men_n52_));
  NA2        u0030(.A(i_7_), .B(i_9_), .Y(men_men_n53_));
  NO2        u0031(.A(men_men_n53_), .B(men_men_n52_), .Y(men_men_n54_));
  OAI210     u0032(.A0(men_men_n54_), .A1(men_men_n51_), .B0(men_men_n45_), .Y(men_men_n55_));
  NA3        u0033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n56_));
  NO2        u0034(.A(i_1_), .B(i_6_), .Y(men_men_n57_));
  NA2        u0035(.A(i_8_), .B(i_7_), .Y(men_men_n58_));
  OAI210     u0036(.A0(men_men_n58_), .A1(men_men_n57_), .B0(men_men_n56_), .Y(men_men_n59_));
  NA2        u0037(.A(men_men_n59_), .B(i_12_), .Y(men_men_n60_));
  NAi21      u0038(.An(i_2_), .B(i_7_), .Y(men_men_n61_));
  INV        u0039(.A(i_1_), .Y(men_men_n62_));
  NA2        u0040(.A(men_men_n62_), .B(i_6_), .Y(men_men_n63_));
  NA2        u0041(.A(i_1_), .B(i_10_), .Y(men_men_n64_));
  NO2        u0042(.A(men_men_n64_), .B(i_6_), .Y(men_men_n65_));
  NAi21      u0043(.An(men_men_n65_), .B(men_men_n60_), .Y(men_men_n66_));
  NA2        u0044(.A(men_men_n50_), .B(i_2_), .Y(men_men_n67_));
  AOI210     u0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n68_));
  NA2        u0046(.A(i_1_), .B(i_6_), .Y(men_men_n69_));
  NO2        u0047(.A(men_men_n69_), .B(men_men_n25_), .Y(men_men_n70_));
  INV        u0048(.A(i_0_), .Y(men_men_n71_));
  NAi21      u0049(.An(i_5_), .B(i_10_), .Y(men_men_n72_));
  NA2        u0050(.A(i_5_), .B(i_9_), .Y(men_men_n73_));
  AOI210     u0051(.A0(men_men_n73_), .A1(men_men_n72_), .B0(men_men_n71_), .Y(men_men_n74_));
  NO2        u0052(.A(men_men_n74_), .B(men_men_n70_), .Y(men_men_n75_));
  OAI210     u0053(.A0(men_men_n68_), .A1(men_men_n67_), .B0(men_men_n75_), .Y(men_men_n76_));
  OAI210     u0054(.A0(men_men_n76_), .A1(men_men_n66_), .B0(i_0_), .Y(men_men_n77_));
  NA2        u0055(.A(i_12_), .B(i_5_), .Y(men_men_n78_));
  NA2        u0056(.A(i_2_), .B(i_8_), .Y(men_men_n79_));
  NO2        u0057(.A(men_men_n79_), .B(men_men_n57_), .Y(men_men_n80_));
  NO2        u0058(.A(i_3_), .B(i_9_), .Y(men_men_n81_));
  NO2        u0059(.A(i_3_), .B(i_7_), .Y(men_men_n82_));
  NO2        u0060(.A(men_men_n82_), .B(men_men_n62_), .Y(men_men_n83_));
  INV        u0061(.A(i_6_), .Y(men_men_n84_));
  OR4        u0062(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n85_));
  INV        u0063(.A(men_men_n85_), .Y(men_men_n86_));
  NO2        u0064(.A(i_2_), .B(i_7_), .Y(men_men_n87_));
  OAI210     u0065(.A0(men_men_n83_), .A1(men_men_n80_), .B0(men_men_n85_), .Y(men_men_n88_));
  NAi21      u0066(.An(i_6_), .B(i_10_), .Y(men_men_n89_));
  NA2        u0067(.A(i_6_), .B(i_9_), .Y(men_men_n90_));
  AOI210     u0068(.A0(men_men_n90_), .A1(men_men_n89_), .B0(men_men_n62_), .Y(men_men_n91_));
  NA2        u0069(.A(i_2_), .B(i_6_), .Y(men_men_n92_));
  AOI210     u0070(.A0(men_men_n90_), .A1(men_men_n88_), .B0(men_men_n78_), .Y(men_men_n93_));
  AN3        u0071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n94_));
  NAi21      u0072(.An(i_6_), .B(i_11_), .Y(men_men_n95_));
  NO2        u0073(.A(i_5_), .B(i_8_), .Y(men_men_n96_));
  NA2        u0074(.A(men_men_n94_), .B(men_men_n32_), .Y(men_men_n97_));
  INV        u0075(.A(i_7_), .Y(men_men_n98_));
  NO2        u0076(.A(i_0_), .B(i_5_), .Y(men_men_n99_));
  NO2        u0077(.A(men_men_n99_), .B(men_men_n84_), .Y(men_men_n100_));
  NA2        u0078(.A(i_12_), .B(i_3_), .Y(men_men_n101_));
  INV        u0079(.A(men_men_n101_), .Y(men_men_n102_));
  NAi21      u0080(.An(i_7_), .B(i_11_), .Y(men_men_n103_));
  NO3        u0081(.A(men_men_n103_), .B(men_men_n89_), .C(men_men_n52_), .Y(men_men_n104_));
  AN2        u0082(.A(i_2_), .B(i_10_), .Y(men_men_n105_));
  NO2        u0083(.A(men_men_n105_), .B(i_7_), .Y(men_men_n106_));
  OR2        u0084(.A(men_men_n78_), .B(men_men_n57_), .Y(men_men_n107_));
  NO2        u0085(.A(i_8_), .B(men_men_n98_), .Y(men_men_n108_));
  NA2        u0086(.A(i_12_), .B(i_7_), .Y(men_men_n109_));
  NO2        u0087(.A(men_men_n62_), .B(men_men_n26_), .Y(men_men_n110_));
  NA2        u0088(.A(men_men_n110_), .B(i_0_), .Y(men_men_n111_));
  NA2        u0089(.A(i_11_), .B(i_12_), .Y(men_men_n112_));
  OAI210     u0090(.A0(men_men_n111_), .A1(men_men_n109_), .B0(men_men_n112_), .Y(men_men_n113_));
  INV        u0091(.A(men_men_n113_), .Y(men_men_n114_));
  NAi31      u0092(.An(men_men_n104_), .B(men_men_n114_), .C(men_men_n97_), .Y(men_men_n115_));
  NOi21      u0093(.An(i_1_), .B(i_5_), .Y(men_men_n116_));
  NA2        u0094(.A(men_men_n116_), .B(i_11_), .Y(men_men_n117_));
  NA2        u0095(.A(men_men_n98_), .B(men_men_n37_), .Y(men_men_n118_));
  NA2        u0096(.A(i_7_), .B(men_men_n25_), .Y(men_men_n119_));
  NA2        u0097(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NO2        u0098(.A(men_men_n120_), .B(men_men_n46_), .Y(men_men_n121_));
  NA2        u0099(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n122_));
  NAi21      u0100(.An(i_3_), .B(i_8_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n123_), .B(men_men_n61_), .Y(men_men_n124_));
  NOi31      u0102(.An(men_men_n124_), .B(men_men_n122_), .C(men_men_n121_), .Y(men_men_n125_));
  NO2        u0103(.A(i_1_), .B(men_men_n84_), .Y(men_men_n126_));
  NO2        u0104(.A(i_6_), .B(i_5_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n127_), .B(i_3_), .Y(men_men_n128_));
  AO210      u0106(.A0(men_men_n128_), .A1(men_men_n47_), .B0(men_men_n126_), .Y(men_men_n129_));
  OAI220     u0107(.A0(men_men_n129_), .A1(men_men_n103_), .B0(men_men_n125_), .B1(men_men_n117_), .Y(men_men_n130_));
  NO3        u0108(.A(men_men_n130_), .B(men_men_n115_), .C(men_men_n93_), .Y(men_men_n131_));
  NA3        u0109(.A(men_men_n131_), .B(men_men_n77_), .C(men_men_n55_), .Y(men2));
  NO2        u0110(.A(men_men_n62_), .B(men_men_n37_), .Y(men_men_n133_));
  NA2        u0111(.A(i_6_), .B(men_men_n25_), .Y(men_men_n134_));
  NA2        u0112(.A(men_men_n134_), .B(men_men_n133_), .Y(men_men_n135_));
  NA4        u0113(.A(men_men_n135_), .B(men_men_n75_), .C(men_men_n67_), .D(men_men_n30_), .Y(men0));
  AN2        u0114(.A(i_8_), .B(i_7_), .Y(men_men_n137_));
  NA2        u0115(.A(men_men_n137_), .B(i_6_), .Y(men_men_n138_));
  NO2        u0116(.A(i_12_), .B(i_13_), .Y(men_men_n139_));
  NAi21      u0117(.An(i_5_), .B(i_11_), .Y(men_men_n140_));
  NOi21      u0118(.An(men_men_n139_), .B(men_men_n140_), .Y(men_men_n141_));
  NO2        u0119(.A(i_0_), .B(i_1_), .Y(men_men_n142_));
  NA2        u0120(.A(i_2_), .B(i_3_), .Y(men_men_n143_));
  NO2        u0121(.A(men_men_n143_), .B(i_4_), .Y(men_men_n144_));
  NA3        u0122(.A(men_men_n144_), .B(men_men_n142_), .C(men_men_n141_), .Y(men_men_n145_));
  OR2        u0123(.A(men_men_n145_), .B(men_men_n25_), .Y(men_men_n146_));
  AN2        u0124(.A(men_men_n139_), .B(men_men_n81_), .Y(men_men_n147_));
  NO2        u0125(.A(men_men_n147_), .B(men_men_n27_), .Y(men_men_n148_));
  NA2        u0126(.A(i_1_), .B(i_5_), .Y(men_men_n149_));
  NO2        u0127(.A(men_men_n71_), .B(men_men_n46_), .Y(men_men_n150_));
  NA2        u0128(.A(men_men_n150_), .B(men_men_n36_), .Y(men_men_n151_));
  NO3        u0129(.A(men_men_n151_), .B(men_men_n149_), .C(men_men_n148_), .Y(men_men_n152_));
  OR2        u0130(.A(i_0_), .B(i_1_), .Y(men_men_n153_));
  NO3        u0131(.A(men_men_n153_), .B(men_men_n78_), .C(i_13_), .Y(men_men_n154_));
  NAi32      u0132(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n155_));
  NAi21      u0133(.An(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  NOi21      u0134(.An(i_4_), .B(i_10_), .Y(men_men_n157_));
  NA2        u0135(.A(men_men_n157_), .B(men_men_n39_), .Y(men_men_n158_));
  NO2        u0136(.A(i_3_), .B(i_5_), .Y(men_men_n159_));
  NO3        u0137(.A(men_men_n71_), .B(i_2_), .C(i_1_), .Y(men_men_n160_));
  NA2        u0138(.A(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  OAI210     u0139(.A0(men_men_n161_), .A1(men_men_n158_), .B0(men_men_n156_), .Y(men_men_n162_));
  NO2        u0140(.A(men_men_n162_), .B(men_men_n152_), .Y(men_men_n163_));
  AOI210     u0141(.A0(men_men_n163_), .A1(men_men_n146_), .B0(men_men_n138_), .Y(men_men_n164_));
  NA3        u0142(.A(men_men_n71_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n165_));
  NA2        u0143(.A(i_3_), .B(men_men_n48_), .Y(men_men_n166_));
  NOi21      u0144(.An(i_4_), .B(i_9_), .Y(men_men_n167_));
  NOi21      u0145(.An(i_11_), .B(i_13_), .Y(men_men_n168_));
  NA2        u0146(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  OR2        u0147(.A(men_men_n169_), .B(men_men_n166_), .Y(men_men_n170_));
  NO2        u0148(.A(i_4_), .B(i_5_), .Y(men_men_n171_));
  NAi21      u0149(.An(i_12_), .B(i_11_), .Y(men_men_n172_));
  NO2        u0150(.A(men_men_n172_), .B(i_13_), .Y(men_men_n173_));
  NA3        u0151(.A(men_men_n173_), .B(men_men_n171_), .C(men_men_n81_), .Y(men_men_n174_));
  AOI210     u0152(.A0(men_men_n174_), .A1(men_men_n170_), .B0(men_men_n165_), .Y(men_men_n175_));
  NO2        u0153(.A(men_men_n71_), .B(men_men_n62_), .Y(men_men_n176_));
  NA2        u0154(.A(men_men_n176_), .B(men_men_n46_), .Y(men_men_n177_));
  NA2        u0155(.A(men_men_n36_), .B(i_5_), .Y(men_men_n178_));
  NAi31      u0156(.An(men_men_n178_), .B(men_men_n147_), .C(i_11_), .Y(men_men_n179_));
  NA2        u0157(.A(i_3_), .B(i_5_), .Y(men_men_n180_));
  OR2        u0158(.A(men_men_n180_), .B(men_men_n169_), .Y(men_men_n181_));
  AOI210     u0159(.A0(men_men_n181_), .A1(men_men_n179_), .B0(men_men_n177_), .Y(men_men_n182_));
  NO2        u0160(.A(men_men_n71_), .B(i_5_), .Y(men_men_n183_));
  NO2        u0161(.A(i_13_), .B(i_10_), .Y(men_men_n184_));
  NA3        u0162(.A(men_men_n184_), .B(men_men_n183_), .C(men_men_n44_), .Y(men_men_n185_));
  NO2        u0163(.A(i_2_), .B(i_1_), .Y(men_men_n186_));
  NA2        u0164(.A(men_men_n186_), .B(i_3_), .Y(men_men_n187_));
  NAi21      u0165(.An(i_4_), .B(i_12_), .Y(men_men_n188_));
  NO4        u0166(.A(men_men_n188_), .B(men_men_n187_), .C(men_men_n185_), .D(men_men_n25_), .Y(men_men_n189_));
  NO3        u0167(.A(men_men_n189_), .B(men_men_n182_), .C(men_men_n175_), .Y(men_men_n190_));
  INV        u0168(.A(i_8_), .Y(men_men_n191_));
  NO2        u0169(.A(men_men_n191_), .B(i_7_), .Y(men_men_n192_));
  NA2        u0170(.A(men_men_n192_), .B(i_6_), .Y(men_men_n193_));
  NO3        u0171(.A(i_3_), .B(men_men_n84_), .C(men_men_n48_), .Y(men_men_n194_));
  NA2        u0172(.A(men_men_n194_), .B(men_men_n108_), .Y(men_men_n195_));
  NO3        u0173(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n196_));
  NA3        u0174(.A(men_men_n196_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n197_));
  NO3        u0175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n198_));
  OAI210     u0176(.A0(men_men_n94_), .A1(i_12_), .B0(men_men_n198_), .Y(men_men_n199_));
  AOI210     u0177(.A0(men_men_n199_), .A1(men_men_n197_), .B0(men_men_n195_), .Y(men_men_n200_));
  NO2        u0178(.A(i_3_), .B(i_8_), .Y(men_men_n201_));
  NO3        u0179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n202_));
  NA3        u0180(.A(men_men_n202_), .B(men_men_n201_), .C(men_men_n39_), .Y(men_men_n203_));
  NO2        u0181(.A(men_men_n99_), .B(men_men_n57_), .Y(men_men_n204_));
  NO2        u0182(.A(i_13_), .B(i_9_), .Y(men_men_n205_));
  NA3        u0183(.A(men_men_n205_), .B(i_6_), .C(men_men_n191_), .Y(men_men_n206_));
  NAi21      u0184(.An(i_12_), .B(i_3_), .Y(men_men_n207_));
  OR2        u0185(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  NO2        u0186(.A(men_men_n44_), .B(i_5_), .Y(men_men_n209_));
  NA2        u0187(.A(men_men_n209_), .B(i_10_), .Y(men_men_n210_));
  OAI220     u0188(.A0(men_men_n210_), .A1(men_men_n208_), .B0(men_men_n99_), .B1(men_men_n203_), .Y(men_men_n211_));
  AOI210     u0189(.A0(men_men_n211_), .A1(i_7_), .B0(men_men_n200_), .Y(men_men_n212_));
  OAI220     u0190(.A0(men_men_n212_), .A1(i_4_), .B0(men_men_n193_), .B1(men_men_n190_), .Y(men_men_n213_));
  NAi21      u0191(.An(i_12_), .B(i_7_), .Y(men_men_n214_));
  NA3        u0192(.A(i_13_), .B(men_men_n191_), .C(i_10_), .Y(men_men_n215_));
  NO2        u0193(.A(men_men_n215_), .B(men_men_n214_), .Y(men_men_n216_));
  NA2        u0194(.A(i_0_), .B(i_5_), .Y(men_men_n217_));
  NA2        u0195(.A(men_men_n217_), .B(men_men_n100_), .Y(men_men_n218_));
  OAI220     u0196(.A0(men_men_n218_), .A1(men_men_n187_), .B0(men_men_n177_), .B1(men_men_n128_), .Y(men_men_n219_));
  NAi31      u0197(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n220_));
  NO2        u0198(.A(men_men_n36_), .B(i_13_), .Y(men_men_n221_));
  NO2        u0199(.A(men_men_n71_), .B(men_men_n26_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n46_), .B(men_men_n62_), .Y(men_men_n223_));
  NA3        u0201(.A(men_men_n223_), .B(men_men_n222_), .C(men_men_n221_), .Y(men_men_n224_));
  INV        u0202(.A(i_13_), .Y(men_men_n225_));
  NO2        u0203(.A(i_12_), .B(men_men_n225_), .Y(men_men_n226_));
  NA3        u0204(.A(men_men_n226_), .B(men_men_n196_), .C(men_men_n194_), .Y(men_men_n227_));
  OAI210     u0205(.A0(men_men_n224_), .A1(men_men_n220_), .B0(men_men_n227_), .Y(men_men_n228_));
  AOI220     u0206(.A0(men_men_n228_), .A1(men_men_n137_), .B0(men_men_n219_), .B1(men_men_n216_), .Y(men_men_n229_));
  NO2        u0207(.A(i_12_), .B(men_men_n37_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n180_), .B(i_4_), .Y(men_men_n231_));
  OR2        u0209(.A(i_8_), .B(i_7_), .Y(men_men_n232_));
  NO2        u0210(.A(men_men_n232_), .B(men_men_n84_), .Y(men_men_n233_));
  NO2        u0211(.A(men_men_n52_), .B(i_1_), .Y(men_men_n234_));
  NA2        u0212(.A(men_men_n234_), .B(men_men_n233_), .Y(men_men_n235_));
  INV        u0213(.A(i_12_), .Y(men_men_n236_));
  NO2        u0214(.A(men_men_n44_), .B(men_men_n236_), .Y(men_men_n237_));
  NO3        u0215(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n238_));
  NA2        u0216(.A(i_2_), .B(i_1_), .Y(men_men_n239_));
  NO2        u0217(.A(men_men_n235_), .B(men_men_n180_), .Y(men_men_n240_));
  NO3        u0218(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n241_));
  NAi21      u0219(.An(i_4_), .B(i_3_), .Y(men_men_n242_));
  NO2        u0220(.A(men_men_n242_), .B(men_men_n73_), .Y(men_men_n243_));
  NO2        u0221(.A(i_0_), .B(i_6_), .Y(men_men_n244_));
  NOi41      u0222(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n245_));
  NA2        u0223(.A(men_men_n245_), .B(men_men_n244_), .Y(men_men_n246_));
  NO2        u0224(.A(men_men_n239_), .B(men_men_n180_), .Y(men_men_n247_));
  NAi21      u0225(.An(men_men_n246_), .B(men_men_n247_), .Y(men_men_n248_));
  INV        u0226(.A(men_men_n248_), .Y(men_men_n249_));
  AOI220     u0227(.A0(men_men_n249_), .A1(men_men_n39_), .B0(men_men_n240_), .B1(men_men_n205_), .Y(men_men_n250_));
  NO2        u0228(.A(i_11_), .B(men_men_n225_), .Y(men_men_n251_));
  NOi21      u0229(.An(i_1_), .B(i_6_), .Y(men_men_n252_));
  NAi21      u0230(.An(i_3_), .B(i_7_), .Y(men_men_n253_));
  NA2        u0231(.A(men_men_n236_), .B(i_9_), .Y(men_men_n254_));
  OR4        u0232(.A(men_men_n254_), .B(men_men_n253_), .C(men_men_n252_), .D(men_men_n183_), .Y(men_men_n255_));
  NO2        u0233(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n256_));
  NO2        u0234(.A(i_12_), .B(i_3_), .Y(men_men_n257_));
  NA2        u0235(.A(men_men_n71_), .B(i_5_), .Y(men_men_n258_));
  NA2        u0236(.A(i_3_), .B(i_9_), .Y(men_men_n259_));
  NAi21      u0237(.An(i_7_), .B(i_10_), .Y(men_men_n260_));
  NO2        u0238(.A(men_men_n260_), .B(men_men_n259_), .Y(men_men_n261_));
  NA3        u0239(.A(men_men_n261_), .B(men_men_n258_), .C(men_men_n63_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n262_), .B(men_men_n255_), .Y(men_men_n263_));
  NA3        u0241(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n264_));
  INV        u0242(.A(men_men_n138_), .Y(men_men_n265_));
  NA2        u0243(.A(men_men_n236_), .B(i_13_), .Y(men_men_n266_));
  NO2        u0244(.A(men_men_n266_), .B(men_men_n73_), .Y(men_men_n267_));
  AOI220     u0245(.A0(men_men_n267_), .A1(men_men_n265_), .B0(men_men_n263_), .B1(men_men_n251_), .Y(men_men_n268_));
  NO2        u0246(.A(men_men_n232_), .B(men_men_n37_), .Y(men_men_n269_));
  NA2        u0247(.A(i_12_), .B(i_6_), .Y(men_men_n270_));
  OR2        u0248(.A(i_13_), .B(i_9_), .Y(men_men_n271_));
  NO3        u0249(.A(men_men_n271_), .B(men_men_n270_), .C(men_men_n48_), .Y(men_men_n272_));
  NO2        u0250(.A(men_men_n242_), .B(i_2_), .Y(men_men_n273_));
  NA3        u0251(.A(men_men_n273_), .B(men_men_n272_), .C(men_men_n44_), .Y(men_men_n274_));
  NA2        u0252(.A(men_men_n251_), .B(i_9_), .Y(men_men_n275_));
  OAI210     u0253(.A0(men_men_n71_), .A1(men_men_n275_), .B0(men_men_n274_), .Y(men_men_n276_));
  NA2        u0254(.A(men_men_n150_), .B(men_men_n62_), .Y(men_men_n277_));
  NO3        u0255(.A(i_11_), .B(men_men_n225_), .C(men_men_n25_), .Y(men_men_n278_));
  NO2        u0256(.A(i_6_), .B(men_men_n48_), .Y(men_men_n279_));
  NA3        u0257(.A(men_men_n279_), .B(i_7_), .C(men_men_n278_), .Y(men_men_n280_));
  NO3        u0258(.A(men_men_n26_), .B(men_men_n84_), .C(i_5_), .Y(men_men_n281_));
  NA3        u0259(.A(men_men_n281_), .B(men_men_n269_), .C(men_men_n226_), .Y(men_men_n282_));
  AOI210     u0260(.A0(men_men_n282_), .A1(men_men_n280_), .B0(men_men_n277_), .Y(men_men_n283_));
  AOI210     u0261(.A0(men_men_n276_), .A1(men_men_n269_), .B0(men_men_n283_), .Y(men_men_n284_));
  NA4        u0262(.A(men_men_n284_), .B(men_men_n268_), .C(men_men_n250_), .D(men_men_n229_), .Y(men_men_n285_));
  NO3        u0263(.A(i_12_), .B(men_men_n225_), .C(men_men_n37_), .Y(men_men_n286_));
  INV        u0264(.A(men_men_n286_), .Y(men_men_n287_));
  NOi21      u0265(.An(men_men_n159_), .B(men_men_n84_), .Y(men_men_n288_));
  NO3        u0266(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n289_));
  AOI220     u0267(.A0(men_men_n289_), .A1(men_men_n194_), .B0(men_men_n288_), .B1(men_men_n234_), .Y(men_men_n290_));
  NO2        u0268(.A(men_men_n290_), .B(i_7_), .Y(men_men_n291_));
  NO3        u0269(.A(i_0_), .B(i_2_), .C(men_men_n62_), .Y(men_men_n292_));
  NO2        u0270(.A(men_men_n239_), .B(i_0_), .Y(men_men_n293_));
  AOI220     u0271(.A0(men_men_n293_), .A1(men_men_n192_), .B0(men_men_n292_), .B1(men_men_n137_), .Y(men_men_n294_));
  NA2        u0272(.A(men_men_n279_), .B(men_men_n26_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n295_), .B(men_men_n294_), .Y(men_men_n296_));
  NA2        u0274(.A(i_0_), .B(i_1_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n297_), .B(i_2_), .Y(men_men_n298_));
  NO2        u0276(.A(men_men_n58_), .B(i_6_), .Y(men_men_n299_));
  NA3        u0277(.A(men_men_n299_), .B(men_men_n298_), .C(men_men_n159_), .Y(men_men_n300_));
  OAI210     u0278(.A0(men_men_n161_), .A1(men_men_n138_), .B0(men_men_n300_), .Y(men_men_n301_));
  NO3        u0279(.A(men_men_n301_), .B(men_men_n296_), .C(men_men_n291_), .Y(men_men_n302_));
  NO2        u0280(.A(i_3_), .B(i_10_), .Y(men_men_n303_));
  NA3        u0281(.A(men_men_n303_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n304_));
  NO2        u0282(.A(i_4_), .B(i_8_), .Y(men_men_n305_));
  NOi21      u0283(.An(men_men_n217_), .B(men_men_n99_), .Y(men_men_n306_));
  NA3        u0284(.A(men_men_n306_), .B(men_men_n305_), .C(i_7_), .Y(men_men_n307_));
  AN2        u0285(.A(i_3_), .B(i_10_), .Y(men_men_n308_));
  NA4        u0286(.A(men_men_n308_), .B(men_men_n196_), .C(men_men_n173_), .D(men_men_n171_), .Y(men_men_n309_));
  NO2        u0287(.A(i_5_), .B(men_men_n37_), .Y(men_men_n310_));
  NO2        u0288(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n311_));
  OR2        u0289(.A(men_men_n307_), .B(men_men_n304_), .Y(men_men_n312_));
  OAI220     u0290(.A0(men_men_n312_), .A1(i_6_), .B0(men_men_n302_), .B1(men_men_n287_), .Y(men_men_n313_));
  NO4        u0291(.A(men_men_n313_), .B(men_men_n285_), .C(men_men_n213_), .D(men_men_n164_), .Y(men_men_n314_));
  NO3        u0292(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n315_));
  NO3        u0293(.A(i_6_), .B(men_men_n191_), .C(i_7_), .Y(men_men_n316_));
  AOI210     u0294(.A0(men_men_n1104_), .A1(men_men_n239_), .B0(men_men_n166_), .Y(men_men_n317_));
  NO2        u0295(.A(i_2_), .B(i_3_), .Y(men_men_n318_));
  OR2        u0296(.A(i_0_), .B(i_5_), .Y(men_men_n319_));
  NA2        u0297(.A(men_men_n217_), .B(men_men_n319_), .Y(men_men_n320_));
  NA4        u0298(.A(men_men_n320_), .B(men_men_n233_), .C(men_men_n318_), .D(i_1_), .Y(men_men_n321_));
  NA3        u0299(.A(men_men_n293_), .B(men_men_n288_), .C(men_men_n108_), .Y(men_men_n322_));
  NAi21      u0300(.An(i_8_), .B(i_7_), .Y(men_men_n323_));
  NO2        u0301(.A(men_men_n323_), .B(i_6_), .Y(men_men_n324_));
  NO2        u0302(.A(men_men_n153_), .B(men_men_n46_), .Y(men_men_n325_));
  NA3        u0303(.A(men_men_n325_), .B(men_men_n324_), .C(men_men_n159_), .Y(men_men_n326_));
  NA3        u0304(.A(men_men_n326_), .B(men_men_n322_), .C(men_men_n321_), .Y(men_men_n327_));
  OAI210     u0305(.A0(men_men_n327_), .A1(men_men_n317_), .B0(i_4_), .Y(men_men_n328_));
  NO2        u0306(.A(i_12_), .B(i_10_), .Y(men_men_n329_));
  NOi21      u0307(.An(i_5_), .B(i_0_), .Y(men_men_n330_));
  AOI210     u0308(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n98_), .Y(men_men_n331_));
  NO4        u0309(.A(men_men_n331_), .B(i_4_), .C(men_men_n330_), .D(men_men_n123_), .Y(men_men_n332_));
  NA4        u0310(.A(men_men_n82_), .B(men_men_n36_), .C(men_men_n84_), .D(i_8_), .Y(men_men_n333_));
  NA2        u0311(.A(men_men_n332_), .B(men_men_n329_), .Y(men_men_n334_));
  NO2        u0312(.A(i_6_), .B(i_8_), .Y(men_men_n335_));
  NOi21      u0313(.An(i_0_), .B(i_2_), .Y(men_men_n336_));
  AN2        u0314(.A(men_men_n336_), .B(men_men_n335_), .Y(men_men_n337_));
  NO2        u0315(.A(i_1_), .B(i_7_), .Y(men_men_n338_));
  AO220      u0316(.A0(men_men_n338_), .A1(men_men_n337_), .B0(men_men_n324_), .B1(men_men_n234_), .Y(men_men_n339_));
  NA3        u0317(.A(men_men_n339_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n340_));
  NA3        u0318(.A(men_men_n340_), .B(men_men_n334_), .C(men_men_n328_), .Y(men_men_n341_));
  AOI210     u0319(.A0(i_8_), .A1(i_8_), .B0(men_men_n320_), .Y(men_men_n342_));
  NOi21      u0320(.An(men_men_n149_), .B(men_men_n100_), .Y(men_men_n343_));
  NO2        u0321(.A(men_men_n343_), .B(men_men_n119_), .Y(men_men_n344_));
  OAI210     u0322(.A0(men_men_n344_), .A1(men_men_n342_), .B0(i_3_), .Y(men_men_n345_));
  INV        u0323(.A(men_men_n82_), .Y(men_men_n346_));
  NO2        u0324(.A(men_men_n297_), .B(men_men_n79_), .Y(men_men_n347_));
  NA2        u0325(.A(men_men_n347_), .B(men_men_n127_), .Y(men_men_n348_));
  NO2        u0326(.A(men_men_n92_), .B(men_men_n191_), .Y(men_men_n349_));
  NA3        u0327(.A(men_men_n306_), .B(men_men_n349_), .C(men_men_n62_), .Y(men_men_n350_));
  AOI210     u0328(.A0(men_men_n350_), .A1(men_men_n348_), .B0(men_men_n346_), .Y(men_men_n351_));
  NO2        u0329(.A(men_men_n191_), .B(i_9_), .Y(men_men_n352_));
  NA3        u0330(.A(men_men_n352_), .B(men_men_n204_), .C(men_men_n153_), .Y(men_men_n353_));
  NO2        u0331(.A(men_men_n353_), .B(men_men_n46_), .Y(men_men_n354_));
  NO3        u0332(.A(men_men_n354_), .B(men_men_n351_), .C(men_men_n296_), .Y(men_men_n355_));
  AOI210     u0333(.A0(men_men_n355_), .A1(men_men_n345_), .B0(men_men_n158_), .Y(men_men_n356_));
  AOI210     u0334(.A0(men_men_n341_), .A1(men_men_n315_), .B0(men_men_n356_), .Y(men_men_n357_));
  NOi32      u0335(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n358_));
  INV        u0336(.A(men_men_n358_), .Y(men_men_n359_));
  NAi21      u0337(.An(i_0_), .B(i_6_), .Y(men_men_n360_));
  NAi21      u0338(.An(i_1_), .B(i_5_), .Y(men_men_n361_));
  NA2        u0339(.A(men_men_n361_), .B(men_men_n360_), .Y(men_men_n362_));
  NA2        u0340(.A(men_men_n362_), .B(men_men_n25_), .Y(men_men_n363_));
  OAI210     u0341(.A0(men_men_n363_), .A1(men_men_n155_), .B0(men_men_n246_), .Y(men_men_n364_));
  NAi41      u0342(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n365_));
  OAI220     u0343(.A0(men_men_n365_), .A1(men_men_n361_), .B0(men_men_n220_), .B1(men_men_n155_), .Y(men_men_n366_));
  AOI210     u0344(.A0(men_men_n365_), .A1(men_men_n155_), .B0(men_men_n153_), .Y(men_men_n367_));
  NOi32      u0345(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n368_));
  NAi21      u0346(.An(i_6_), .B(i_1_), .Y(men_men_n369_));
  NA3        u0347(.A(men_men_n369_), .B(men_men_n368_), .C(men_men_n46_), .Y(men_men_n370_));
  NO2        u0348(.A(men_men_n370_), .B(i_0_), .Y(men_men_n371_));
  OR3        u0349(.A(men_men_n371_), .B(men_men_n367_), .C(men_men_n366_), .Y(men_men_n372_));
  NO2        u0350(.A(i_1_), .B(men_men_n98_), .Y(men_men_n373_));
  NAi21      u0351(.An(i_3_), .B(i_4_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n374_), .B(i_9_), .Y(men_men_n375_));
  AN2        u0353(.A(i_6_), .B(i_7_), .Y(men_men_n376_));
  OAI210     u0354(.A0(men_men_n376_), .A1(men_men_n373_), .B0(men_men_n375_), .Y(men_men_n377_));
  NA2        u0355(.A(i_2_), .B(i_7_), .Y(men_men_n378_));
  NO2        u0356(.A(men_men_n374_), .B(i_10_), .Y(men_men_n379_));
  NA3        u0357(.A(men_men_n379_), .B(men_men_n378_), .C(men_men_n244_), .Y(men_men_n380_));
  AOI210     u0358(.A0(men_men_n380_), .A1(men_men_n377_), .B0(men_men_n183_), .Y(men_men_n381_));
  AOI210     u0359(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n382_));
  OAI210     u0360(.A0(men_men_n382_), .A1(men_men_n186_), .B0(men_men_n379_), .Y(men_men_n383_));
  AOI220     u0361(.A0(men_men_n379_), .A1(men_men_n338_), .B0(men_men_n238_), .B1(men_men_n186_), .Y(men_men_n384_));
  AOI210     u0362(.A0(men_men_n384_), .A1(men_men_n383_), .B0(i_5_), .Y(men_men_n385_));
  NO4        u0363(.A(men_men_n385_), .B(men_men_n381_), .C(men_men_n372_), .D(men_men_n364_), .Y(men_men_n386_));
  NO2        u0364(.A(men_men_n386_), .B(men_men_n359_), .Y(men_men_n387_));
  NO2        u0365(.A(men_men_n58_), .B(men_men_n25_), .Y(men_men_n388_));
  AN2        u0366(.A(i_12_), .B(i_5_), .Y(men_men_n389_));
  NO2        u0367(.A(i_4_), .B(men_men_n26_), .Y(men_men_n390_));
  NA2        u0368(.A(men_men_n390_), .B(men_men_n389_), .Y(men_men_n391_));
  NO2        u0369(.A(i_11_), .B(i_6_), .Y(men_men_n392_));
  NA3        u0370(.A(men_men_n392_), .B(men_men_n325_), .C(men_men_n225_), .Y(men_men_n393_));
  NO2        u0371(.A(men_men_n393_), .B(men_men_n391_), .Y(men_men_n394_));
  NO2        u0372(.A(men_men_n242_), .B(i_5_), .Y(men_men_n395_));
  NO2        u0373(.A(i_5_), .B(i_10_), .Y(men_men_n396_));
  AOI220     u0374(.A0(men_men_n396_), .A1(men_men_n273_), .B0(men_men_n395_), .B1(men_men_n196_), .Y(men_men_n397_));
  NO2        u0375(.A(i_6_), .B(men_men_n397_), .Y(men_men_n398_));
  OAI210     u0376(.A0(men_men_n398_), .A1(men_men_n394_), .B0(men_men_n388_), .Y(men_men_n399_));
  NO2        u0377(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n400_));
  NO2        u0378(.A(men_men_n145_), .B(men_men_n84_), .Y(men_men_n401_));
  OAI210     u0379(.A0(men_men_n401_), .A1(men_men_n394_), .B0(men_men_n400_), .Y(men_men_n402_));
  NO3        u0380(.A(men_men_n84_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n403_));
  NO2        u0381(.A(i_3_), .B(men_men_n98_), .Y(men_men_n404_));
  NA4        u0382(.A(men_men_n303_), .B(men_men_n90_), .C(men_men_n73_), .D(men_men_n53_), .Y(men_men_n405_));
  NO2        u0383(.A(i_11_), .B(i_12_), .Y(men_men_n406_));
  NA2        u0384(.A(men_men_n406_), .B(men_men_n36_), .Y(men_men_n407_));
  NO2        u0385(.A(men_men_n405_), .B(men_men_n407_), .Y(men_men_n408_));
  NA2        u0386(.A(men_men_n396_), .B(men_men_n236_), .Y(men_men_n409_));
  NA3        u0387(.A(men_men_n108_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n410_));
  OAI220     u0388(.A0(men_men_n410_), .A1(men_men_n220_), .B0(men_men_n409_), .B1(men_men_n333_), .Y(men_men_n411_));
  NAi21      u0389(.An(i_13_), .B(i_0_), .Y(men_men_n412_));
  NO2        u0390(.A(men_men_n412_), .B(men_men_n239_), .Y(men_men_n413_));
  OAI210     u0391(.A0(men_men_n411_), .A1(men_men_n408_), .B0(men_men_n413_), .Y(men_men_n414_));
  NA3        u0392(.A(men_men_n414_), .B(men_men_n402_), .C(men_men_n399_), .Y(men_men_n415_));
  NA2        u0393(.A(men_men_n44_), .B(men_men_n225_), .Y(men_men_n416_));
  NO3        u0394(.A(i_1_), .B(i_12_), .C(men_men_n84_), .Y(men_men_n417_));
  NO2        u0395(.A(i_0_), .B(i_11_), .Y(men_men_n418_));
  AN2        u0396(.A(i_1_), .B(i_6_), .Y(men_men_n419_));
  NOi21      u0397(.An(i_2_), .B(i_12_), .Y(men_men_n420_));
  NA2        u0398(.A(men_men_n420_), .B(men_men_n419_), .Y(men_men_n421_));
  NO2        u0399(.A(men_men_n421_), .B(men_men_n1095_), .Y(men_men_n422_));
  NA2        u0400(.A(men_men_n137_), .B(i_9_), .Y(men_men_n423_));
  NO2        u0401(.A(men_men_n423_), .B(i_4_), .Y(men_men_n424_));
  NA2        u0402(.A(men_men_n422_), .B(men_men_n424_), .Y(men_men_n425_));
  NAi21      u0403(.An(i_9_), .B(i_4_), .Y(men_men_n426_));
  OR2        u0404(.A(i_13_), .B(i_10_), .Y(men_men_n427_));
  NO3        u0405(.A(men_men_n427_), .B(men_men_n112_), .C(men_men_n426_), .Y(men_men_n428_));
  NO2        u0406(.A(men_men_n169_), .B(men_men_n118_), .Y(men_men_n429_));
  OR2        u0407(.A(men_men_n215_), .B(men_men_n214_), .Y(men_men_n430_));
  NO2        u0408(.A(men_men_n98_), .B(men_men_n25_), .Y(men_men_n431_));
  NA2        u0409(.A(men_men_n286_), .B(men_men_n431_), .Y(men_men_n432_));
  NA2        u0410(.A(men_men_n279_), .B(i_1_), .Y(men_men_n433_));
  OAI220     u0411(.A0(men_men_n433_), .A1(men_men_n430_), .B0(men_men_n432_), .B1(men_men_n343_), .Y(men_men_n434_));
  INV        u0412(.A(men_men_n434_), .Y(men_men_n435_));
  AOI210     u0413(.A0(men_men_n435_), .A1(men_men_n425_), .B0(men_men_n26_), .Y(men_men_n436_));
  NA2        u0414(.A(men_men_n322_), .B(men_men_n321_), .Y(men_men_n437_));
  AOI220     u0415(.A0(men_men_n299_), .A1(men_men_n289_), .B0(men_men_n293_), .B1(i_6_), .Y(men_men_n438_));
  NO2        u0416(.A(men_men_n438_), .B(men_men_n166_), .Y(men_men_n439_));
  NO2        u0417(.A(men_men_n180_), .B(men_men_n84_), .Y(men_men_n440_));
  AOI220     u0418(.A0(men_men_n440_), .A1(men_men_n298_), .B0(men_men_n281_), .B1(i_1_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n441_), .B(i_7_), .Y(men_men_n442_));
  NO3        u0420(.A(men_men_n442_), .B(men_men_n439_), .C(men_men_n437_), .Y(men_men_n443_));
  NA2        u0421(.A(men_men_n194_), .B(men_men_n94_), .Y(men_men_n444_));
  NA3        u0422(.A(men_men_n325_), .B(men_men_n159_), .C(men_men_n84_), .Y(men_men_n445_));
  AOI210     u0423(.A0(men_men_n445_), .A1(men_men_n444_), .B0(men_men_n323_), .Y(men_men_n446_));
  NA2        u0424(.A(men_men_n191_), .B(i_10_), .Y(men_men_n447_));
  NA3        u0425(.A(men_men_n258_), .B(men_men_n63_), .C(i_2_), .Y(men_men_n448_));
  NA2        u0426(.A(men_men_n299_), .B(men_men_n234_), .Y(men_men_n449_));
  OAI220     u0427(.A0(men_men_n449_), .A1(men_men_n180_), .B0(men_men_n448_), .B1(men_men_n447_), .Y(men_men_n450_));
  NO2        u0428(.A(i_3_), .B(men_men_n48_), .Y(men_men_n451_));
  NA3        u0429(.A(men_men_n338_), .B(men_men_n337_), .C(men_men_n451_), .Y(men_men_n452_));
  NA2        u0430(.A(men_men_n316_), .B(men_men_n320_), .Y(men_men_n453_));
  OAI210     u0431(.A0(men_men_n453_), .A1(men_men_n187_), .B0(men_men_n452_), .Y(men_men_n454_));
  NO3        u0432(.A(men_men_n454_), .B(men_men_n450_), .C(men_men_n446_), .Y(men_men_n455_));
  AOI210     u0433(.A0(men_men_n455_), .A1(men_men_n443_), .B0(men_men_n275_), .Y(men_men_n456_));
  NO4        u0434(.A(men_men_n456_), .B(men_men_n436_), .C(men_men_n415_), .D(men_men_n387_), .Y(men_men_n457_));
  NO2        u0435(.A(men_men_n71_), .B(i_13_), .Y(men_men_n458_));
  NO2        u0436(.A(i_10_), .B(i_9_), .Y(men_men_n459_));
  NAi21      u0437(.An(i_12_), .B(i_8_), .Y(men_men_n460_));
  NO2        u0438(.A(men_men_n460_), .B(i_3_), .Y(men_men_n461_));
  NO2        u0439(.A(men_men_n46_), .B(i_4_), .Y(men_men_n462_));
  NA2        u0440(.A(men_men_n462_), .B(men_men_n100_), .Y(men_men_n463_));
  NO2        u0441(.A(men_men_n463_), .B(men_men_n203_), .Y(men_men_n464_));
  NA2        u0442(.A(men_men_n311_), .B(i_0_), .Y(men_men_n465_));
  NO3        u0443(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n466_));
  NA2        u0444(.A(men_men_n270_), .B(men_men_n95_), .Y(men_men_n467_));
  NA2        u0445(.A(men_men_n467_), .B(men_men_n466_), .Y(men_men_n468_));
  NA2        u0446(.A(i_8_), .B(i_9_), .Y(men_men_n469_));
  NA2        u0447(.A(men_men_n286_), .B(men_men_n204_), .Y(men_men_n470_));
  OAI220     u0448(.A0(men_men_n470_), .A1(men_men_n469_), .B0(men_men_n468_), .B1(men_men_n465_), .Y(men_men_n471_));
  NA2        u0449(.A(men_men_n251_), .B(men_men_n310_), .Y(men_men_n472_));
  NO3        u0450(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n473_));
  AOI210     u0451(.A0(men_men_n257_), .A1(men_men_n186_), .B0(men_men_n473_), .Y(men_men_n474_));
  NA3        u0452(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n475_));
  NA4        u0453(.A(men_men_n140_), .B(men_men_n110_), .C(men_men_n78_), .D(men_men_n23_), .Y(men_men_n476_));
  OAI220     u0454(.A0(men_men_n476_), .A1(men_men_n475_), .B0(men_men_n474_), .B1(men_men_n472_), .Y(men_men_n477_));
  NO3        u0455(.A(men_men_n477_), .B(men_men_n471_), .C(men_men_n464_), .Y(men_men_n478_));
  NA2        u0456(.A(men_men_n298_), .B(men_men_n103_), .Y(men_men_n479_));
  OR2        u0457(.A(men_men_n479_), .B(men_men_n206_), .Y(men_men_n480_));
  OA210      u0458(.A0(men_men_n353_), .A1(men_men_n98_), .B0(men_men_n300_), .Y(men_men_n481_));
  OA220      u0459(.A0(men_men_n481_), .A1(men_men_n158_), .B0(men_men_n480_), .B1(men_men_n180_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n94_), .B(i_13_), .Y(men_men_n483_));
  NA2        u0461(.A(men_men_n440_), .B(men_men_n388_), .Y(men_men_n484_));
  NO2        u0462(.A(i_2_), .B(i_13_), .Y(men_men_n485_));
  NO2        u0463(.A(men_men_n484_), .B(men_men_n483_), .Y(men_men_n486_));
  NO3        u0464(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n487_));
  NO2        u0465(.A(i_6_), .B(i_7_), .Y(men_men_n488_));
  NA2        u0466(.A(men_men_n488_), .B(men_men_n487_), .Y(men_men_n489_));
  OR2        u0467(.A(i_11_), .B(i_8_), .Y(men_men_n490_));
  NOi21      u0468(.An(i_2_), .B(i_7_), .Y(men_men_n491_));
  NAi31      u0469(.An(men_men_n490_), .B(men_men_n491_), .C(men_men_n1097_), .Y(men_men_n492_));
  NO2        u0470(.A(men_men_n427_), .B(i_6_), .Y(men_men_n493_));
  NA3        u0471(.A(men_men_n493_), .B(men_men_n1100_), .C(men_men_n73_), .Y(men_men_n494_));
  NO2        u0472(.A(men_men_n494_), .B(men_men_n492_), .Y(men_men_n495_));
  NO2        u0473(.A(i_3_), .B(men_men_n191_), .Y(men_men_n496_));
  NO2        u0474(.A(i_6_), .B(i_10_), .Y(men_men_n497_));
  NA4        u0475(.A(men_men_n497_), .B(men_men_n315_), .C(men_men_n496_), .D(men_men_n236_), .Y(men_men_n498_));
  NO2        u0476(.A(men_men_n498_), .B(men_men_n151_), .Y(men_men_n499_));
  NA3        u0477(.A(men_men_n245_), .B(men_men_n168_), .C(men_men_n127_), .Y(men_men_n500_));
  NA2        u0478(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n501_));
  NO2        u0479(.A(men_men_n153_), .B(i_3_), .Y(men_men_n502_));
  NAi31      u0480(.An(men_men_n501_), .B(men_men_n502_), .C(men_men_n226_), .Y(men_men_n503_));
  NA3        u0481(.A(men_men_n400_), .B(men_men_n176_), .C(men_men_n144_), .Y(men_men_n504_));
  NA3        u0482(.A(men_men_n504_), .B(men_men_n503_), .C(men_men_n500_), .Y(men_men_n505_));
  NO4        u0483(.A(men_men_n505_), .B(men_men_n499_), .C(men_men_n495_), .D(men_men_n486_), .Y(men_men_n506_));
  NA2        u0484(.A(men_men_n473_), .B(men_men_n396_), .Y(men_men_n507_));
  NO2        u0485(.A(men_men_n507_), .B(men_men_n224_), .Y(men_men_n508_));
  NAi21      u0486(.An(men_men_n215_), .B(men_men_n406_), .Y(men_men_n509_));
  NO2        u0487(.A(men_men_n26_), .B(i_5_), .Y(men_men_n510_));
  NO2        u0488(.A(i_0_), .B(men_men_n84_), .Y(men_men_n511_));
  NA3        u0489(.A(men_men_n511_), .B(men_men_n510_), .C(men_men_n137_), .Y(men_men_n512_));
  OAI220     u0490(.A0(men_men_n38_), .A1(men_men_n512_), .B0(i_0_), .B1(men_men_n509_), .Y(men_men_n513_));
  NA2        u0491(.A(men_men_n27_), .B(i_10_), .Y(men_men_n514_));
  NA2        u0492(.A(men_men_n315_), .B(men_men_n238_), .Y(men_men_n515_));
  OAI220     u0493(.A0(men_men_n515_), .A1(men_men_n448_), .B0(men_men_n514_), .B1(men_men_n483_), .Y(men_men_n516_));
  NA4        u0494(.A(men_men_n308_), .B(men_men_n223_), .C(men_men_n71_), .D(men_men_n236_), .Y(men_men_n517_));
  NO2        u0495(.A(men_men_n517_), .B(men_men_n489_), .Y(men_men_n518_));
  NO4        u0496(.A(men_men_n518_), .B(men_men_n516_), .C(men_men_n513_), .D(men_men_n508_), .Y(men_men_n519_));
  NA4        u0497(.A(men_men_n519_), .B(men_men_n506_), .C(men_men_n482_), .D(men_men_n478_), .Y(men_men_n520_));
  NA3        u0498(.A(men_men_n308_), .B(men_men_n173_), .C(men_men_n171_), .Y(men_men_n521_));
  OAI210     u0499(.A0(men_men_n304_), .A1(men_men_n178_), .B0(men_men_n521_), .Y(men_men_n522_));
  AN2        u0500(.A(men_men_n289_), .B(men_men_n233_), .Y(men_men_n523_));
  NA2        u0501(.A(men_men_n523_), .B(men_men_n522_), .Y(men_men_n524_));
  NA2        u0502(.A(men_men_n117_), .B(men_men_n107_), .Y(men_men_n525_));
  AO220      u0503(.A0(men_men_n525_), .A1(men_men_n466_), .B0(men_men_n428_), .B1(i_6_), .Y(men_men_n526_));
  NA2        u0504(.A(men_men_n315_), .B(men_men_n160_), .Y(men_men_n527_));
  OAI210     u0505(.A0(men_men_n527_), .A1(men_men_n180_), .B0(men_men_n309_), .Y(men_men_n528_));
  AOI220     u0506(.A0(men_men_n528_), .A1(men_men_n324_), .B0(men_men_n526_), .B1(men_men_n311_), .Y(men_men_n529_));
  NA2        u0507(.A(men_men_n389_), .B(men_men_n225_), .Y(men_men_n530_));
  NA2        u0508(.A(men_men_n358_), .B(men_men_n71_), .Y(men_men_n531_));
  NA2        u0509(.A(men_men_n376_), .B(men_men_n368_), .Y(men_men_n532_));
  AO210      u0510(.A0(men_men_n531_), .A1(men_men_n530_), .B0(men_men_n532_), .Y(men_men_n533_));
  NO2        u0511(.A(men_men_n36_), .B(i_8_), .Y(men_men_n534_));
  NAi41      u0512(.An(men_men_n531_), .B(men_men_n497_), .C(men_men_n534_), .D(men_men_n46_), .Y(men_men_n535_));
  INV        u0513(.A(men_men_n428_), .Y(men_men_n536_));
  NA3        u0514(.A(men_men_n536_), .B(men_men_n535_), .C(men_men_n533_), .Y(men_men_n537_));
  INV        u0515(.A(men_men_n537_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n258_), .B(men_men_n63_), .Y(men_men_n539_));
  OAI210     u0517(.A0(i_8_), .A1(men_men_n539_), .B0(men_men_n129_), .Y(men_men_n540_));
  AOI210     u0518(.A0(men_men_n192_), .A1(i_9_), .B0(men_men_n269_), .Y(men_men_n541_));
  NO2        u0519(.A(men_men_n541_), .B(men_men_n197_), .Y(men_men_n542_));
  AOI220     u0520(.A0(i_6_), .A1(men_men_n542_), .B0(men_men_n540_), .B1(men_men_n429_), .Y(men_men_n543_));
  NA4        u0521(.A(men_men_n543_), .B(men_men_n538_), .C(men_men_n529_), .D(men_men_n524_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n395_), .B(men_men_n298_), .Y(men_men_n545_));
  OAI210     u0523(.A0(men_men_n391_), .A1(men_men_n165_), .B0(men_men_n545_), .Y(men_men_n546_));
  NO2        u0524(.A(i_12_), .B(men_men_n191_), .Y(men_men_n547_));
  NA2        u0525(.A(men_men_n547_), .B(men_men_n225_), .Y(men_men_n548_));
  NA3        u0526(.A(men_men_n497_), .B(men_men_n171_), .C(men_men_n27_), .Y(men_men_n549_));
  NO3        u0527(.A(men_men_n549_), .B(men_men_n548_), .C(men_men_n479_), .Y(men_men_n550_));
  NOi31      u0528(.An(men_men_n316_), .B(men_men_n427_), .C(men_men_n38_), .Y(men_men_n551_));
  OAI210     u0529(.A0(men_men_n551_), .A1(men_men_n550_), .B0(men_men_n546_), .Y(men_men_n552_));
  NO2        u0530(.A(i_8_), .B(i_7_), .Y(men_men_n553_));
  OAI210     u0531(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n554_), .B(men_men_n223_), .Y(men_men_n555_));
  AOI220     u0533(.A0(men_men_n325_), .A1(men_men_n39_), .B0(men_men_n234_), .B1(men_men_n205_), .Y(men_men_n556_));
  OAI220     u0534(.A0(men_men_n556_), .A1(men_men_n180_), .B0(men_men_n555_), .B1(men_men_n242_), .Y(men_men_n557_));
  NA2        u0535(.A(men_men_n44_), .B(i_10_), .Y(men_men_n558_));
  NO2        u0536(.A(men_men_n558_), .B(i_6_), .Y(men_men_n559_));
  NA3        u0537(.A(men_men_n559_), .B(men_men_n557_), .C(men_men_n553_), .Y(men_men_n560_));
  AOI220     u0538(.A0(men_men_n440_), .A1(men_men_n325_), .B0(men_men_n247_), .B1(men_men_n244_), .Y(men_men_n561_));
  OAI220     u0539(.A0(men_men_n561_), .A1(men_men_n266_), .B0(men_men_n483_), .B1(men_men_n128_), .Y(men_men_n562_));
  NA2        u0540(.A(men_men_n562_), .B(men_men_n269_), .Y(men_men_n563_));
  NOi31      u0541(.An(men_men_n293_), .B(men_men_n304_), .C(men_men_n178_), .Y(men_men_n564_));
  NA3        u0542(.A(men_men_n308_), .B(men_men_n171_), .C(men_men_n94_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n221_), .B(men_men_n44_), .Y(men_men_n566_));
  NO2        u0544(.A(men_men_n153_), .B(i_5_), .Y(men_men_n567_));
  NA3        u0545(.A(men_men_n567_), .B(men_men_n416_), .C(men_men_n318_), .Y(men_men_n568_));
  OAI210     u0546(.A0(men_men_n568_), .A1(men_men_n566_), .B0(men_men_n565_), .Y(men_men_n569_));
  OAI210     u0547(.A0(men_men_n569_), .A1(men_men_n564_), .B0(men_men_n473_), .Y(men_men_n570_));
  NA4        u0548(.A(men_men_n570_), .B(men_men_n563_), .C(men_men_n560_), .D(men_men_n552_), .Y(men_men_n571_));
  NA2        u0549(.A(men_men_n286_), .B(men_men_n82_), .Y(men_men_n572_));
  AOI210     u0550(.A0(i_11_), .A1(men_men_n348_), .B0(men_men_n572_), .Y(men_men_n573_));
  NA2        u0551(.A(men_men_n299_), .B(men_men_n289_), .Y(men_men_n574_));
  NO2        u0552(.A(men_men_n574_), .B(men_men_n170_), .Y(men_men_n575_));
  NA2        u0553(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n576_));
  NA2        u0554(.A(men_men_n459_), .B(men_men_n221_), .Y(men_men_n577_));
  NO2        u0555(.A(men_men_n576_), .B(men_men_n577_), .Y(men_men_n578_));
  NA2        u0556(.A(i_0_), .B(men_men_n48_), .Y(men_men_n579_));
  NA3        u0557(.A(men_men_n547_), .B(men_men_n278_), .C(men_men_n579_), .Y(men_men_n580_));
  NO2        u0558(.A(men_men_n1101_), .B(men_men_n580_), .Y(men_men_n581_));
  NO4        u0559(.A(men_men_n581_), .B(men_men_n578_), .C(men_men_n575_), .D(men_men_n573_), .Y(men_men_n582_));
  NO4        u0560(.A(men_men_n252_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n583_));
  NO3        u0561(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n584_));
  NO2        u0562(.A(men_men_n232_), .B(men_men_n36_), .Y(men_men_n585_));
  AN2        u0563(.A(men_men_n585_), .B(men_men_n584_), .Y(men_men_n586_));
  OA210      u0564(.A0(men_men_n586_), .A1(men_men_n583_), .B0(men_men_n358_), .Y(men_men_n587_));
  NO2        u0565(.A(men_men_n427_), .B(i_1_), .Y(men_men_n588_));
  NOi31      u0566(.An(men_men_n588_), .B(men_men_n467_), .C(men_men_n71_), .Y(men_men_n589_));
  AN4        u0567(.A(men_men_n589_), .B(men_men_n424_), .C(men_men_n510_), .D(i_2_), .Y(men_men_n590_));
  NO2        u0568(.A(men_men_n438_), .B(men_men_n174_), .Y(men_men_n591_));
  NO3        u0569(.A(men_men_n591_), .B(men_men_n590_), .C(men_men_n587_), .Y(men_men_n592_));
  NOi21      u0570(.An(i_10_), .B(i_6_), .Y(men_men_n593_));
  NO2        u0571(.A(men_men_n84_), .B(men_men_n25_), .Y(men_men_n594_));
  AOI220     u0572(.A0(men_men_n286_), .A1(men_men_n594_), .B0(men_men_n278_), .B1(men_men_n593_), .Y(men_men_n595_));
  NO2        u0573(.A(men_men_n595_), .B(men_men_n465_), .Y(men_men_n596_));
  NO2        u0574(.A(men_men_n109_), .B(men_men_n23_), .Y(men_men_n597_));
  NA2        u0575(.A(men_men_n316_), .B(men_men_n160_), .Y(men_men_n598_));
  AOI220     u0576(.A0(men_men_n598_), .A1(men_men_n449_), .B0(men_men_n181_), .B1(men_men_n179_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n196_), .B(men_men_n37_), .Y(men_men_n600_));
  NOi31      u0578(.An(men_men_n141_), .B(men_men_n600_), .C(men_men_n333_), .Y(men_men_n601_));
  NO3        u0579(.A(men_men_n601_), .B(men_men_n599_), .C(men_men_n596_), .Y(men_men_n602_));
  NO2        u0580(.A(men_men_n531_), .B(men_men_n384_), .Y(men_men_n603_));
  INV        u0581(.A(men_men_n318_), .Y(men_men_n604_));
  NO2        u0582(.A(i_12_), .B(men_men_n84_), .Y(men_men_n605_));
  NA3        u0583(.A(men_men_n605_), .B(men_men_n278_), .C(men_men_n579_), .Y(men_men_n606_));
  NA3        u0584(.A(men_men_n392_), .B(men_men_n286_), .C(men_men_n217_), .Y(men_men_n607_));
  AOI210     u0585(.A0(men_men_n607_), .A1(men_men_n606_), .B0(men_men_n604_), .Y(men_men_n608_));
  NA2        u0586(.A(men_men_n171_), .B(i_0_), .Y(men_men_n609_));
  NO3        u0587(.A(men_men_n609_), .B(i_8_), .C(men_men_n304_), .Y(men_men_n610_));
  OR2        u0588(.A(i_2_), .B(i_5_), .Y(men_men_n611_));
  OR2        u0589(.A(men_men_n611_), .B(men_men_n419_), .Y(men_men_n612_));
  AOI210     u0590(.A0(i_0_), .A1(men_men_n612_), .B0(men_men_n509_), .Y(men_men_n613_));
  NO4        u0591(.A(men_men_n613_), .B(men_men_n610_), .C(men_men_n608_), .D(men_men_n603_), .Y(men_men_n614_));
  NA4        u0592(.A(men_men_n614_), .B(men_men_n602_), .C(men_men_n592_), .D(men_men_n582_), .Y(men_men_n615_));
  NO4        u0593(.A(men_men_n615_), .B(men_men_n571_), .C(men_men_n544_), .D(men_men_n520_), .Y(men_men_n616_));
  NA4        u0594(.A(men_men_n616_), .B(men_men_n457_), .C(men_men_n357_), .D(men_men_n314_), .Y(men7));
  NO2        u0595(.A(men_men_n103_), .B(men_men_n89_), .Y(men_men_n618_));
  NA2        u0596(.A(men_men_n390_), .B(men_men_n618_), .Y(men_men_n619_));
  NA2        u0597(.A(men_men_n497_), .B(men_men_n82_), .Y(men_men_n620_));
  NA2        u0598(.A(i_11_), .B(men_men_n191_), .Y(men_men_n621_));
  OAI210     u0599(.A0(men_men_n1102_), .A1(men_men_n620_), .B0(men_men_n619_), .Y(men_men_n622_));
  NA3        u0600(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n623_));
  NO2        u0601(.A(men_men_n236_), .B(i_4_), .Y(men_men_n624_));
  NA2        u0602(.A(men_men_n624_), .B(i_8_), .Y(men_men_n625_));
  AOI210     u0603(.A0(men_men_n625_), .A1(men_men_n101_), .B0(men_men_n623_), .Y(men_men_n626_));
  NA2        u0604(.A(i_2_), .B(men_men_n84_), .Y(men_men_n627_));
  OAI210     u0605(.A0(men_men_n87_), .A1(men_men_n201_), .B0(men_men_n202_), .Y(men_men_n628_));
  NO2        u0606(.A(i_7_), .B(men_men_n37_), .Y(men_men_n629_));
  NA2        u0607(.A(i_4_), .B(i_8_), .Y(men_men_n630_));
  AOI210     u0608(.A0(men_men_n630_), .A1(men_men_n308_), .B0(men_men_n629_), .Y(men_men_n631_));
  OAI220     u0609(.A0(men_men_n631_), .A1(men_men_n627_), .B0(men_men_n628_), .B1(i_13_), .Y(men_men_n632_));
  NO3        u0610(.A(men_men_n632_), .B(men_men_n626_), .C(men_men_n622_), .Y(men_men_n633_));
  AOI210     u0611(.A0(men_men_n123_), .A1(men_men_n61_), .B0(i_10_), .Y(men_men_n634_));
  AOI210     u0612(.A0(men_men_n634_), .A1(men_men_n236_), .B0(men_men_n157_), .Y(men_men_n635_));
  OR2        u0613(.A(i_6_), .B(i_10_), .Y(men_men_n636_));
  NO2        u0614(.A(men_men_n636_), .B(men_men_n23_), .Y(men_men_n637_));
  OR3        u0615(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n638_));
  NO3        u0616(.A(men_men_n638_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n639_));
  INV        u0617(.A(men_men_n198_), .Y(men_men_n640_));
  NO2        u0618(.A(men_men_n639_), .B(men_men_n637_), .Y(men_men_n641_));
  OA220      u0619(.A0(men_men_n641_), .A1(men_men_n604_), .B0(men_men_n635_), .B1(men_men_n271_), .Y(men_men_n642_));
  AOI210     u0620(.A0(men_men_n642_), .A1(men_men_n633_), .B0(men_men_n62_), .Y(men_men_n643_));
  NOi21      u0621(.An(i_11_), .B(i_7_), .Y(men_men_n644_));
  AO210      u0622(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n645_));
  NO2        u0623(.A(men_men_n645_), .B(men_men_n644_), .Y(men_men_n646_));
  NA3        u0624(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n647_));
  NAi31      u0625(.An(men_men_n647_), .B(men_men_n214_), .C(i_11_), .Y(men_men_n648_));
  NO2        u0626(.A(men_men_n648_), .B(men_men_n62_), .Y(men_men_n649_));
  AO210      u0627(.A0(men_men_n85_), .A1(men_men_n384_), .B0(men_men_n40_), .Y(men_men_n650_));
  NO3        u0628(.A(men_men_n260_), .B(men_men_n207_), .C(men_men_n621_), .Y(men_men_n651_));
  OAI210     u0629(.A0(men_men_n651_), .A1(men_men_n226_), .B0(men_men_n62_), .Y(men_men_n652_));
  NA2        u0630(.A(men_men_n420_), .B(men_men_n31_), .Y(men_men_n653_));
  OR2        u0631(.A(men_men_n207_), .B(men_men_n103_), .Y(men_men_n654_));
  NA2        u0632(.A(men_men_n654_), .B(men_men_n653_), .Y(men_men_n655_));
  NO2        u0633(.A(men_men_n62_), .B(i_9_), .Y(men_men_n656_));
  NA2        u0634(.A(men_men_n62_), .B(men_men_n655_), .Y(men_men_n657_));
  NO2        u0635(.A(i_1_), .B(i_12_), .Y(men_men_n658_));
  NA3        u0636(.A(men_men_n658_), .B(men_men_n105_), .C(men_men_n24_), .Y(men_men_n659_));
  NA4        u0637(.A(men_men_n659_), .B(men_men_n657_), .C(men_men_n652_), .D(men_men_n650_), .Y(men_men_n660_));
  OAI210     u0638(.A0(men_men_n660_), .A1(men_men_n649_), .B0(i_6_), .Y(men_men_n661_));
  OAI210     u0639(.A0(men_men_n647_), .A1(men_men_n103_), .B0(men_men_n475_), .Y(men_men_n662_));
  NA2        u0640(.A(men_men_n662_), .B(men_men_n605_), .Y(men_men_n663_));
  NO2        u0641(.A(i_6_), .B(i_11_), .Y(men_men_n664_));
  NA3        u0642(.A(men_men_n663_), .B(men_men_n536_), .C(men_men_n468_), .Y(men_men_n665_));
  NO4        u0643(.A(men_men_n214_), .B(men_men_n123_), .C(i_13_), .D(men_men_n84_), .Y(men_men_n666_));
  NA2        u0644(.A(men_men_n666_), .B(men_men_n656_), .Y(men_men_n667_));
  NO3        u0645(.A(men_men_n636_), .B(men_men_n232_), .C(men_men_n23_), .Y(men_men_n668_));
  AOI210     u0646(.A0(i_1_), .A1(men_men_n261_), .B0(men_men_n668_), .Y(men_men_n669_));
  OAI210     u0647(.A0(men_men_n669_), .A1(men_men_n44_), .B0(men_men_n667_), .Y(men_men_n670_));
  NA3        u0648(.A(men_men_n553_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n671_));
  NA2        u0649(.A(men_men_n133_), .B(i_9_), .Y(men_men_n672_));
  NA3        u0650(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n673_));
  NO2        u0651(.A(men_men_n46_), .B(i_1_), .Y(men_men_n674_));
  NA3        u0652(.A(men_men_n674_), .B(men_men_n270_), .C(men_men_n44_), .Y(men_men_n675_));
  OAI220     u0653(.A0(men_men_n675_), .A1(men_men_n673_), .B0(men_men_n672_), .B1(men_men_n1094_), .Y(men_men_n676_));
  NA3        u0654(.A(men_men_n656_), .B(men_men_n318_), .C(i_6_), .Y(men_men_n677_));
  NO2        u0655(.A(men_men_n677_), .B(men_men_n23_), .Y(men_men_n678_));
  NAi21      u0656(.An(men_men_n671_), .B(men_men_n91_), .Y(men_men_n679_));
  NA2        u0657(.A(men_men_n674_), .B(men_men_n270_), .Y(men_men_n680_));
  NO2        u0658(.A(i_11_), .B(men_men_n37_), .Y(men_men_n681_));
  NA2        u0659(.A(men_men_n681_), .B(men_men_n24_), .Y(men_men_n682_));
  OAI210     u0660(.A0(men_men_n682_), .A1(men_men_n680_), .B0(men_men_n679_), .Y(men_men_n683_));
  OR3        u0661(.A(men_men_n683_), .B(men_men_n678_), .C(men_men_n676_), .Y(men_men_n684_));
  NO3        u0662(.A(men_men_n684_), .B(men_men_n670_), .C(men_men_n665_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n236_), .B(men_men_n98_), .Y(men_men_n686_));
  NO2        u0664(.A(men_men_n686_), .B(men_men_n644_), .Y(men_men_n687_));
  NO2        u0665(.A(men_men_n426_), .B(men_men_n84_), .Y(men_men_n688_));
  NA2        u0666(.A(i_3_), .B(men_men_n191_), .Y(men_men_n689_));
  AN2        u0667(.A(men_men_n1105_), .B(men_men_n559_), .Y(men_men_n690_));
  NO2        u0668(.A(men_men_n232_), .B(men_men_n44_), .Y(men_men_n691_));
  NO3        u0669(.A(men_men_n691_), .B(men_men_n311_), .C(men_men_n237_), .Y(men_men_n692_));
  NO2        u0670(.A(men_men_n112_), .B(men_men_n37_), .Y(men_men_n693_));
  NO2        u0671(.A(men_men_n693_), .B(i_6_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n84_), .B(i_9_), .Y(men_men_n695_));
  NO2        u0673(.A(men_men_n695_), .B(men_men_n62_), .Y(men_men_n696_));
  NO2        u0674(.A(men_men_n696_), .B(men_men_n658_), .Y(men_men_n697_));
  NO4        u0675(.A(men_men_n697_), .B(men_men_n694_), .C(men_men_n692_), .D(i_4_), .Y(men_men_n698_));
  NA2        u0676(.A(i_1_), .B(i_3_), .Y(men_men_n699_));
  NO2        u0677(.A(men_men_n469_), .B(men_men_n92_), .Y(men_men_n700_));
  AOI210     u0678(.A0(men_men_n691_), .A1(men_men_n593_), .B0(men_men_n700_), .Y(men_men_n701_));
  NO2        u0679(.A(men_men_n701_), .B(men_men_n699_), .Y(men_men_n702_));
  NO3        u0680(.A(men_men_n702_), .B(men_men_n698_), .C(men_men_n690_), .Y(men_men_n703_));
  NA3        u0681(.A(men_men_n703_), .B(men_men_n685_), .C(men_men_n661_), .Y(men_men_n704_));
  NO3        u0682(.A(men_men_n490_), .B(i_3_), .C(i_7_), .Y(men_men_n705_));
  OA210      u0683(.A0(men_men_n705_), .A1(men_men_n245_), .B0(men_men_n84_), .Y(men_men_n706_));
  NA2        u0684(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n707_));
  NA3        u0685(.A(men_men_n497_), .B(men_men_n534_), .C(men_men_n46_), .Y(men_men_n708_));
  NO3        u0686(.A(men_men_n491_), .B(men_men_n630_), .C(men_men_n84_), .Y(men_men_n709_));
  NA2        u0687(.A(men_men_n709_), .B(men_men_n25_), .Y(men_men_n710_));
  NA3        u0688(.A(men_men_n157_), .B(men_men_n82_), .C(men_men_n84_), .Y(men_men_n711_));
  NA4        u0689(.A(men_men_n711_), .B(men_men_n710_), .C(men_men_n708_), .D(men_men_n707_), .Y(men_men_n712_));
  OAI210     u0690(.A0(men_men_n712_), .A1(men_men_n706_), .B0(i_1_), .Y(men_men_n713_));
  NO2        u0691(.A(men_men_n374_), .B(i_2_), .Y(men_men_n714_));
  AOI210     u0692(.A0(men_men_n677_), .A1(men_men_n713_), .B0(i_13_), .Y(men_men_n715_));
  OR2        u0693(.A(i_11_), .B(i_7_), .Y(men_men_n716_));
  NA3        u0694(.A(men_men_n716_), .B(men_men_n102_), .C(men_men_n133_), .Y(men_men_n717_));
  AOI220     u0695(.A0(men_men_n485_), .A1(men_men_n157_), .B0(men_men_n462_), .B1(men_men_n133_), .Y(men_men_n718_));
  OAI210     u0696(.A0(men_men_n718_), .A1(men_men_n44_), .B0(men_men_n717_), .Y(men_men_n719_));
  AOI210     u0697(.A0(men_men_n673_), .A1(men_men_n53_), .B0(i_12_), .Y(men_men_n720_));
  NO2        u0698(.A(men_men_n491_), .B(men_men_n24_), .Y(men_men_n721_));
  AOI220     u0699(.A0(men_men_n721_), .A1(men_men_n688_), .B0(men_men_n245_), .B1(men_men_n126_), .Y(men_men_n722_));
  OAI220     u0700(.A0(men_men_n722_), .A1(men_men_n40_), .B0(men_men_n1093_), .B1(men_men_n92_), .Y(men_men_n723_));
  AOI210     u0701(.A0(men_men_n719_), .A1(men_men_n335_), .B0(men_men_n723_), .Y(men_men_n724_));
  NA2        u0702(.A(men_men_n109_), .B(men_men_n103_), .Y(men_men_n725_));
  AOI220     u0703(.A0(men_men_n725_), .A1(men_men_n70_), .B0(men_men_n392_), .B1(men_men_n674_), .Y(men_men_n726_));
  NO2        u0704(.A(men_men_n726_), .B(men_men_n242_), .Y(men_men_n727_));
  AOI210     u0705(.A0(men_men_n460_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n728_));
  NOi31      u0706(.An(men_men_n728_), .B(men_men_n620_), .C(men_men_n44_), .Y(men_men_n729_));
  NA2        u0707(.A(men_men_n122_), .B(i_13_), .Y(men_men_n730_));
  NO2        u0708(.A(men_men_n673_), .B(men_men_n109_), .Y(men_men_n731_));
  INV        u0709(.A(men_men_n731_), .Y(men_men_n732_));
  OAI220     u0710(.A0(men_men_n732_), .A1(men_men_n69_), .B0(men_men_n730_), .B1(men_men_n1099_), .Y(men_men_n733_));
  NO3        u0711(.A(men_men_n69_), .B(men_men_n32_), .C(men_men_n98_), .Y(men_men_n734_));
  NA2        u0712(.A(men_men_n26_), .B(men_men_n191_), .Y(men_men_n735_));
  NA2        u0713(.A(men_men_n735_), .B(i_7_), .Y(men_men_n736_));
  NO3        u0714(.A(men_men_n491_), .B(men_men_n236_), .C(men_men_n84_), .Y(men_men_n737_));
  AOI210     u0715(.A0(men_men_n737_), .A1(men_men_n736_), .B0(men_men_n734_), .Y(men_men_n738_));
  AOI220     u0716(.A0(men_men_n392_), .A1(men_men_n674_), .B0(men_men_n91_), .B1(i_2_), .Y(men_men_n739_));
  OAI220     u0717(.A0(men_men_n739_), .A1(men_men_n625_), .B0(men_men_n738_), .B1(men_men_n640_), .Y(men_men_n740_));
  NO4        u0718(.A(men_men_n740_), .B(men_men_n733_), .C(men_men_n729_), .D(men_men_n727_), .Y(men_men_n741_));
  OR2        u0719(.A(i_11_), .B(i_6_), .Y(men_men_n742_));
  NA3        u0720(.A(men_men_n624_), .B(men_men_n735_), .C(i_7_), .Y(men_men_n743_));
  AOI210     u0721(.A0(men_men_n743_), .A1(men_men_n732_), .B0(men_men_n742_), .Y(men_men_n744_));
  NA2        u0722(.A(men_men_n664_), .B(i_13_), .Y(men_men_n745_));
  NA2        u0723(.A(i_2_), .B(men_men_n735_), .Y(men_men_n746_));
  NAi21      u0724(.An(i_11_), .B(i_12_), .Y(men_men_n747_));
  NOi41      u0725(.An(men_men_n106_), .B(men_men_n747_), .C(i_13_), .D(men_men_n84_), .Y(men_men_n748_));
  NO3        u0726(.A(men_men_n491_), .B(men_men_n605_), .C(men_men_n630_), .Y(men_men_n749_));
  AOI220     u0727(.A0(men_men_n749_), .A1(men_men_n315_), .B0(men_men_n748_), .B1(men_men_n746_), .Y(men_men_n750_));
  NA2        u0728(.A(men_men_n750_), .B(men_men_n745_), .Y(men_men_n751_));
  OAI210     u0729(.A0(men_men_n751_), .A1(men_men_n744_), .B0(men_men_n62_), .Y(men_men_n752_));
  NO2        u0730(.A(i_2_), .B(i_12_), .Y(men_men_n753_));
  OAI210     u0731(.A0(men_men_n634_), .A1(men_men_n373_), .B0(men_men_n753_), .Y(men_men_n754_));
  NA2        u0732(.A(i_8_), .B(men_men_n25_), .Y(men_men_n755_));
  NO3        u0733(.A(men_men_n755_), .B(men_men_n390_), .C(men_men_n624_), .Y(men_men_n756_));
  OAI210     u0734(.A0(men_men_n756_), .A1(men_men_n375_), .B0(men_men_n373_), .Y(men_men_n757_));
  NO2        u0735(.A(men_men_n123_), .B(i_2_), .Y(men_men_n758_));
  NA2        u0736(.A(men_men_n758_), .B(men_men_n658_), .Y(men_men_n759_));
  NA3        u0737(.A(men_men_n759_), .B(men_men_n757_), .C(men_men_n754_), .Y(men_men_n760_));
  NA3        u0738(.A(men_men_n760_), .B(men_men_n45_), .C(men_men_n225_), .Y(men_men_n761_));
  NA4        u0739(.A(men_men_n761_), .B(men_men_n752_), .C(men_men_n741_), .D(men_men_n724_), .Y(men_men_n762_));
  OR4        u0740(.A(men_men_n762_), .B(men_men_n715_), .C(men_men_n704_), .D(men_men_n643_), .Y(men5));
  AOI210     u0741(.A0(men_men_n687_), .A1(men_men_n273_), .B0(men_men_n429_), .Y(men_men_n764_));
  AO210      u0742(.A0(men_men_n24_), .A1(i_10_), .B0(men_men_n251_), .Y(men_men_n765_));
  NA3        u0743(.A(men_men_n765_), .B(men_men_n753_), .C(men_men_n103_), .Y(men_men_n766_));
  NA3        u0744(.A(men_men_n766_), .B(men_men_n764_), .C(men_men_n536_), .Y(men_men_n767_));
  NO3        u0745(.A(i_11_), .B(men_men_n236_), .C(i_13_), .Y(men_men_n768_));
  NO2        u0746(.A(men_men_n119_), .B(men_men_n23_), .Y(men_men_n769_));
  NA2        u0747(.A(i_12_), .B(i_8_), .Y(men_men_n770_));
  INV        u0748(.A(men_men_n459_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n318_), .B(men_men_n597_), .Y(men_men_n772_));
  INV        u0750(.A(men_men_n772_), .Y(men_men_n773_));
  NO2        u0751(.A(men_men_n773_), .B(men_men_n767_), .Y(men_men_n774_));
  INV        u0752(.A(men_men_n168_), .Y(men_men_n775_));
  OAI210     u0753(.A0(men_men_n714_), .A1(men_men_n461_), .B0(men_men_n106_), .Y(men_men_n776_));
  NO2        u0754(.A(men_men_n776_), .B(men_men_n775_), .Y(men_men_n777_));
  NO2        u0755(.A(men_men_n469_), .B(men_men_n26_), .Y(men_men_n778_));
  NO2        u0756(.A(men_men_n778_), .B(men_men_n431_), .Y(men_men_n779_));
  NA2        u0757(.A(men_men_n779_), .B(i_2_), .Y(men_men_n780_));
  INV        u0758(.A(men_men_n780_), .Y(men_men_n781_));
  AOI210     u0759(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n427_), .Y(men_men_n782_));
  AOI210     u0760(.A0(men_men_n782_), .A1(men_men_n781_), .B0(men_men_n777_), .Y(men_men_n783_));
  NO2        u0761(.A(men_men_n188_), .B(men_men_n120_), .Y(men_men_n784_));
  OAI210     u0762(.A0(men_men_n784_), .A1(men_men_n769_), .B0(i_2_), .Y(men_men_n785_));
  INV        u0763(.A(men_men_n169_), .Y(men_men_n786_));
  NO3        u0764(.A(men_men_n645_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n787_));
  AOI210     u0765(.A0(men_men_n786_), .A1(men_men_n87_), .B0(men_men_n787_), .Y(men_men_n788_));
  AOI210     u0766(.A0(men_men_n788_), .A1(men_men_n785_), .B0(men_men_n191_), .Y(men_men_n789_));
  OA210      u0767(.A0(men_men_n646_), .A1(men_men_n121_), .B0(i_13_), .Y(men_men_n790_));
  NA2        u0768(.A(men_men_n198_), .B(men_men_n201_), .Y(men_men_n791_));
  NA2        u0769(.A(men_men_n147_), .B(men_men_n621_), .Y(men_men_n792_));
  AOI210     u0770(.A0(men_men_n792_), .A1(men_men_n791_), .B0(men_men_n378_), .Y(men_men_n793_));
  AOI210     u0771(.A0(men_men_n207_), .A1(men_men_n143_), .B0(men_men_n534_), .Y(men_men_n794_));
  OAI210     u0772(.A0(men_men_n794_), .A1(men_men_n226_), .B0(men_men_n431_), .Y(men_men_n795_));
  NA3        u0773(.A(men_men_n308_), .B(men_men_n119_), .C(men_men_n42_), .Y(men_men_n796_));
  OAI210     u0774(.A0(men_men_n796_), .A1(men_men_n46_), .B0(men_men_n795_), .Y(men_men_n797_));
  NO4        u0775(.A(men_men_n797_), .B(men_men_n793_), .C(men_men_n790_), .D(men_men_n789_), .Y(men_men_n798_));
  NO2        u0776(.A(men_men_n61_), .B(i_12_), .Y(men_men_n799_));
  NO2        u0777(.A(men_men_n799_), .B(men_men_n121_), .Y(men_men_n800_));
  NO2        u0778(.A(men_men_n800_), .B(men_men_n621_), .Y(men_men_n801_));
  NA2        u0779(.A(men_men_n801_), .B(men_men_n36_), .Y(men_men_n802_));
  NA4        u0780(.A(men_men_n802_), .B(men_men_n798_), .C(men_men_n783_), .D(men_men_n774_), .Y(men6));
  NO3        u0781(.A(men_men_n256_), .B(men_men_n310_), .C(i_1_), .Y(men_men_n804_));
  NO2        u0782(.A(men_men_n183_), .B(men_men_n134_), .Y(men_men_n805_));
  OAI210     u0783(.A0(men_men_n805_), .A1(men_men_n804_), .B0(men_men_n758_), .Y(men_men_n806_));
  NA4        u0784(.A(men_men_n396_), .B(men_men_n496_), .C(men_men_n69_), .D(men_men_n98_), .Y(men_men_n807_));
  INV        u0785(.A(men_men_n807_), .Y(men_men_n808_));
  NO2        u0786(.A(men_men_n220_), .B(men_men_n501_), .Y(men_men_n809_));
  NO2        u0787(.A(i_11_), .B(i_9_), .Y(men_men_n810_));
  NO3        u0788(.A(men_men_n809_), .B(men_men_n808_), .C(men_men_n330_), .Y(men_men_n811_));
  AO210      u0789(.A0(men_men_n811_), .A1(men_men_n806_), .B0(i_12_), .Y(men_men_n812_));
  NA2        u0790(.A(men_men_n379_), .B(men_men_n338_), .Y(men_men_n813_));
  NA2        u0791(.A(men_men_n605_), .B(men_men_n62_), .Y(men_men_n814_));
  NA2        u0792(.A(men_men_n705_), .B(men_men_n69_), .Y(men_men_n815_));
  NA4        u0793(.A(men_men_n85_), .B(men_men_n815_), .C(men_men_n814_), .D(men_men_n813_), .Y(men_men_n816_));
  INV        u0794(.A(men_men_n195_), .Y(men_men_n817_));
  AOI220     u0795(.A0(men_men_n817_), .A1(men_men_n810_), .B0(men_men_n816_), .B1(men_men_n71_), .Y(men_men_n818_));
  INV        u0796(.A(men_men_n329_), .Y(men_men_n819_));
  NA2        u0797(.A(men_men_n73_), .B(men_men_n126_), .Y(men_men_n820_));
  INV        u0798(.A(men_men_n119_), .Y(men_men_n821_));
  NA2        u0799(.A(men_men_n821_), .B(men_men_n46_), .Y(men_men_n822_));
  AOI210     u0800(.A0(men_men_n822_), .A1(men_men_n820_), .B0(men_men_n819_), .Y(men_men_n823_));
  NO3        u0801(.A(men_men_n252_), .B(men_men_n127_), .C(i_9_), .Y(men_men_n824_));
  NA2        u0802(.A(men_men_n824_), .B(men_men_n799_), .Y(men_men_n825_));
  AOI210     u0803(.A0(men_men_n825_), .A1(men_men_n532_), .B0(men_men_n183_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n32_), .B(i_11_), .Y(men_men_n827_));
  NA3        u0805(.A(men_men_n827_), .B(men_men_n488_), .C(men_men_n396_), .Y(men_men_n828_));
  OAI210     u0806(.A0(men_men_n705_), .A1(men_men_n585_), .B0(men_men_n584_), .Y(men_men_n829_));
  NA2        u0807(.A(men_men_n829_), .B(men_men_n828_), .Y(men_men_n830_));
  OR3        u0808(.A(men_men_n830_), .B(men_men_n826_), .C(men_men_n823_), .Y(men_men_n831_));
  NO2        u0809(.A(men_men_n716_), .B(i_2_), .Y(men_men_n832_));
  NA2        u0810(.A(men_men_n48_), .B(men_men_n37_), .Y(men_men_n833_));
  NA2        u0811(.A(men_men_n1103_), .B(men_men_n832_), .Y(men_men_n834_));
  AO220      u0812(.A0(men_men_n362_), .A1(men_men_n352_), .B0(men_men_n403_), .B1(men_men_n621_), .Y(men_men_n835_));
  NA3        u0813(.A(men_men_n835_), .B(men_men_n257_), .C(i_7_), .Y(men_men_n836_));
  OR2        u0814(.A(men_men_n646_), .B(men_men_n461_), .Y(men_men_n837_));
  NA3        u0815(.A(men_men_n837_), .B(men_men_n142_), .C(men_men_n67_), .Y(men_men_n838_));
  AO210      u0816(.A0(men_men_n507_), .A1(men_men_n771_), .B0(men_men_n36_), .Y(men_men_n839_));
  NA4        u0817(.A(men_men_n839_), .B(men_men_n838_), .C(men_men_n836_), .D(men_men_n834_), .Y(men_men_n840_));
  OAI210     u0818(.A0(i_6_), .A1(i_11_), .B0(men_men_n85_), .Y(men_men_n841_));
  AOI220     u0819(.A0(men_men_n841_), .A1(men_men_n584_), .B0(men_men_n809_), .B1(men_men_n736_), .Y(men_men_n842_));
  NA3        u0820(.A(men_men_n378_), .B(men_men_n238_), .C(men_men_n142_), .Y(men_men_n843_));
  OAI210     u0821(.A0(men_men_n403_), .A1(men_men_n202_), .B0(men_men_n68_), .Y(men_men_n844_));
  NA4        u0822(.A(men_men_n844_), .B(men_men_n843_), .C(men_men_n842_), .D(men_men_n628_), .Y(men_men_n845_));
  AO210      u0823(.A0(men_men_n534_), .A1(men_men_n46_), .B0(men_men_n86_), .Y(men_men_n846_));
  NA3        u0824(.A(men_men_n846_), .B(men_men_n497_), .C(men_men_n217_), .Y(men_men_n847_));
  AOI210     u0825(.A0(men_men_n461_), .A1(men_men_n459_), .B0(men_men_n583_), .Y(men_men_n848_));
  NO2        u0826(.A(men_men_n636_), .B(i_2_), .Y(men_men_n849_));
  OAI210     u0827(.A0(men_men_n849_), .A1(men_men_n107_), .B0(men_men_n418_), .Y(men_men_n850_));
  NA2        u0828(.A(men_men_n244_), .B(men_men_n46_), .Y(men_men_n851_));
  NA2        u0829(.A(men_men_n851_), .B(men_men_n612_), .Y(men_men_n852_));
  NA3        u0830(.A(men_men_n852_), .B(men_men_n329_), .C(i_7_), .Y(men_men_n853_));
  NA4        u0831(.A(men_men_n853_), .B(men_men_n850_), .C(men_men_n848_), .D(men_men_n847_), .Y(men_men_n854_));
  NO4        u0832(.A(men_men_n854_), .B(men_men_n845_), .C(men_men_n840_), .D(men_men_n831_), .Y(men_men_n855_));
  NA4        u0833(.A(men_men_n855_), .B(men_men_n818_), .C(men_men_n812_), .D(men_men_n386_), .Y(men3));
  NA2        u0834(.A(i_12_), .B(i_10_), .Y(men_men_n857_));
  NA2        u0835(.A(i_6_), .B(i_7_), .Y(men_men_n858_));
  NO2        u0836(.A(men_men_n858_), .B(i_0_), .Y(men_men_n859_));
  NO2        u0837(.A(i_11_), .B(men_men_n236_), .Y(men_men_n860_));
  OAI210     u0838(.A0(men_men_n859_), .A1(men_men_n293_), .B0(men_men_n860_), .Y(men_men_n861_));
  NO2        u0839(.A(men_men_n861_), .B(men_men_n191_), .Y(men_men_n862_));
  NO3        u0840(.A(men_men_n465_), .B(men_men_n89_), .C(men_men_n44_), .Y(men_men_n863_));
  OA210      u0841(.A0(men_men_n863_), .A1(men_men_n862_), .B0(men_men_n171_), .Y(men_men_n864_));
  NA3        u0842(.A(men_men_n843_), .B(men_men_n628_), .C(men_men_n377_), .Y(men_men_n865_));
  NA2        u0843(.A(men_men_n865_), .B(men_men_n39_), .Y(men_men_n866_));
  NOi21      u0844(.An(men_men_n94_), .B(men_men_n779_), .Y(men_men_n867_));
  NO3        u0845(.A(men_men_n654_), .B(men_men_n469_), .C(men_men_n126_), .Y(men_men_n868_));
  NA2        u0846(.A(men_men_n420_), .B(men_men_n45_), .Y(men_men_n869_));
  AN2        u0847(.A(men_men_n467_), .B(men_men_n54_), .Y(men_men_n870_));
  NO3        u0848(.A(men_men_n870_), .B(men_men_n868_), .C(men_men_n867_), .Y(men_men_n871_));
  AOI210     u0849(.A0(men_men_n871_), .A1(men_men_n866_), .B0(men_men_n48_), .Y(men_men_n872_));
  NA2        u0850(.A(men_men_n183_), .B(men_men_n593_), .Y(men_men_n873_));
  NA2        u0851(.A(men_men_n728_), .B(men_men_n695_), .Y(men_men_n874_));
  NA2        u0852(.A(men_men_n336_), .B(men_men_n451_), .Y(men_men_n875_));
  OAI220     u0853(.A0(men_men_n875_), .A1(men_men_n874_), .B0(men_men_n873_), .B1(men_men_n62_), .Y(men_men_n876_));
  NOi21      u0854(.An(i_5_), .B(i_9_), .Y(men_men_n877_));
  NA2        u0855(.A(men_men_n877_), .B(men_men_n458_), .Y(men_men_n878_));
  INV        u0856(.A(men_men_n709_), .Y(men_men_n879_));
  NO3        u0857(.A(men_men_n423_), .B(men_men_n270_), .C(men_men_n71_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n172_), .B(men_men_n143_), .Y(men_men_n881_));
  AOI210     u0859(.A0(men_men_n881_), .A1(men_men_n244_), .B0(men_men_n880_), .Y(men_men_n882_));
  OAI220     u0860(.A0(men_men_n882_), .A1(men_men_n178_), .B0(men_men_n879_), .B1(men_men_n878_), .Y(men_men_n883_));
  NO4        u0861(.A(men_men_n883_), .B(men_men_n876_), .C(men_men_n872_), .D(men_men_n864_), .Y(men_men_n884_));
  NOi21      u0862(.An(i_0_), .B(i_10_), .Y(men_men_n885_));
  NA2        u0863(.A(men_men_n183_), .B(men_men_n24_), .Y(men_men_n886_));
  NO2        u0864(.A(men_men_n693_), .B(men_men_n618_), .Y(men_men_n887_));
  NO2        u0865(.A(men_men_n887_), .B(men_men_n886_), .Y(men_men_n888_));
  NA2        u0866(.A(men_men_n315_), .B(men_men_n124_), .Y(men_men_n889_));
  NAi21      u0867(.An(men_men_n158_), .B(men_men_n451_), .Y(men_men_n890_));
  OAI220     u0868(.A0(men_men_n890_), .A1(men_men_n851_), .B0(men_men_n889_), .B1(men_men_n409_), .Y(men_men_n891_));
  NO2        u0869(.A(men_men_n891_), .B(men_men_n888_), .Y(men_men_n892_));
  NO2        u0870(.A(men_men_n396_), .B(men_men_n297_), .Y(men_men_n893_));
  NA2        u0871(.A(men_men_n893_), .B(men_men_n731_), .Y(men_men_n894_));
  NA2        u0872(.A(men_men_n594_), .B(i_0_), .Y(men_men_n895_));
  NO3        u0873(.A(men_men_n895_), .B(men_men_n391_), .C(men_men_n87_), .Y(men_men_n896_));
  NO4        u0874(.A(men_men_n611_), .B(men_men_n214_), .C(men_men_n427_), .D(men_men_n419_), .Y(men_men_n897_));
  AOI210     u0875(.A0(men_men_n897_), .A1(i_11_), .B0(men_men_n896_), .Y(men_men_n898_));
  INV        u0876(.A(men_men_n488_), .Y(men_men_n899_));
  AN2        u0877(.A(men_men_n94_), .B(men_men_n243_), .Y(men_men_n900_));
  NA2        u0878(.A(men_men_n768_), .B(men_men_n330_), .Y(men_men_n901_));
  AOI210     u0879(.A0(men_men_n497_), .A1(men_men_n87_), .B0(men_men_n57_), .Y(men_men_n902_));
  OAI220     u0880(.A0(men_men_n902_), .A1(men_men_n901_), .B0(men_men_n682_), .B1(men_men_n555_), .Y(men_men_n903_));
  NO2        u0881(.A(men_men_n254_), .B(men_men_n149_), .Y(men_men_n904_));
  NA2        u0882(.A(i_0_), .B(i_10_), .Y(men_men_n905_));
  OAI210     u0883(.A0(men_men_n905_), .A1(men_men_n84_), .B0(men_men_n558_), .Y(men_men_n906_));
  NO4        u0884(.A(men_men_n109_), .B(men_men_n57_), .C(men_men_n689_), .D(i_5_), .Y(men_men_n907_));
  AO220      u0885(.A0(men_men_n907_), .A1(men_men_n906_), .B0(men_men_n904_), .B1(i_6_), .Y(men_men_n908_));
  AOI220     u0886(.A0(men_men_n336_), .A1(men_men_n96_), .B0(men_men_n183_), .B1(men_men_n82_), .Y(men_men_n909_));
  NA2        u0887(.A(men_men_n588_), .B(i_4_), .Y(men_men_n910_));
  NA2        u0888(.A(men_men_n186_), .B(men_men_n201_), .Y(men_men_n911_));
  OAI220     u0889(.A0(men_men_n911_), .A1(men_men_n901_), .B0(men_men_n910_), .B1(men_men_n909_), .Y(men_men_n912_));
  NO4        u0890(.A(men_men_n912_), .B(men_men_n908_), .C(men_men_n903_), .D(men_men_n900_), .Y(men_men_n913_));
  NA4        u0891(.A(men_men_n913_), .B(men_men_n898_), .C(men_men_n894_), .D(men_men_n892_), .Y(men_men_n914_));
  NO2        u0892(.A(men_men_n99_), .B(men_men_n37_), .Y(men_men_n915_));
  NA2        u0893(.A(i_11_), .B(i_9_), .Y(men_men_n916_));
  NO3        u0894(.A(i_12_), .B(men_men_n916_), .C(men_men_n627_), .Y(men_men_n917_));
  AO220      u0895(.A0(men_men_n917_), .A1(men_men_n915_), .B0(men_men_n272_), .B1(men_men_n86_), .Y(men_men_n918_));
  NO2        u0896(.A(men_men_n48_), .B(i_7_), .Y(men_men_n919_));
  NO2        u0897(.A(men_men_n916_), .B(men_men_n71_), .Y(men_men_n920_));
  NO2        u0898(.A(men_men_n172_), .B(i_0_), .Y(men_men_n921_));
  INV        u0899(.A(men_men_n921_), .Y(men_men_n922_));
  NA2        u0900(.A(men_men_n488_), .B(men_men_n231_), .Y(men_men_n923_));
  AOI210     u0901(.A0(men_men_n376_), .A1(men_men_n41_), .B0(men_men_n417_), .Y(men_men_n924_));
  OAI220     u0902(.A0(men_men_n924_), .A1(men_men_n878_), .B0(men_men_n923_), .B1(men_men_n922_), .Y(men_men_n925_));
  NO2        u0903(.A(men_men_n925_), .B(men_men_n918_), .Y(men_men_n926_));
  AOI210     u0904(.A0(men_men_n460_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n927_));
  NA2        u0905(.A(men_men_n168_), .B(men_men_n99_), .Y(men_men_n928_));
  NOi32      u0906(.An(men_men_n927_), .Bn(men_men_n186_), .C(men_men_n928_), .Y(men_men_n929_));
  AOI210     u0907(.A0(men_men_n629_), .A1(men_men_n330_), .B0(men_men_n243_), .Y(men_men_n930_));
  NO2        u0908(.A(men_men_n930_), .B(men_men_n869_), .Y(men_men_n931_));
  NO2        u0909(.A(men_men_n931_), .B(men_men_n929_), .Y(men_men_n932_));
  NOi21      u0910(.An(i_7_), .B(i_5_), .Y(men_men_n933_));
  NOi31      u0911(.An(men_men_n933_), .B(men_men_n885_), .C(men_men_n747_), .Y(men_men_n934_));
  NA3        u0912(.A(men_men_n934_), .B(men_men_n390_), .C(i_6_), .Y(men_men_n935_));
  OA210      u0913(.A0(men_men_n928_), .A1(men_men_n532_), .B0(men_men_n935_), .Y(men_men_n936_));
  NO3        u0914(.A(men_men_n412_), .B(men_men_n365_), .C(men_men_n361_), .Y(men_men_n937_));
  INV        u0915(.A(men_men_n319_), .Y(men_men_n938_));
  NO2        u0916(.A(men_men_n747_), .B(men_men_n259_), .Y(men_men_n939_));
  AOI210     u0917(.A0(men_men_n939_), .A1(men_men_n938_), .B0(men_men_n937_), .Y(men_men_n940_));
  NA4        u0918(.A(men_men_n940_), .B(men_men_n936_), .C(men_men_n932_), .D(men_men_n926_), .Y(men_men_n941_));
  NO2        u0919(.A(men_men_n886_), .B(men_men_n239_), .Y(men_men_n942_));
  AN2        u0920(.A(men_men_n335_), .B(men_men_n330_), .Y(men_men_n943_));
  AO220      u0921(.A0(men_men_n943_), .A1(men_men_n881_), .B0(men_men_n347_), .B1(men_men_n27_), .Y(men_men_n944_));
  OAI210     u0922(.A0(men_men_n944_), .A1(men_men_n942_), .B0(i_10_), .Y(men_men_n945_));
  INV        u0923(.A(men_men_n857_), .Y(men_men_n946_));
  OA210      u0924(.A0(men_men_n488_), .A1(men_men_n223_), .B0(men_men_n487_), .Y(men_men_n947_));
  OAI210     u0925(.A0(men_men_n947_), .A1(men_men_n946_), .B0(men_men_n920_), .Y(men_men_n948_));
  NA3        u0926(.A(men_men_n487_), .B(men_men_n420_), .C(men_men_n45_), .Y(men_men_n949_));
  OAI210     u0927(.A0(men_men_n890_), .A1(men_men_n899_), .B0(men_men_n949_), .Y(men_men_n950_));
  NO2        u0928(.A(men_men_n257_), .B(men_men_n46_), .Y(men_men_n951_));
  NA2        u0929(.A(men_men_n920_), .B(men_men_n308_), .Y(men_men_n952_));
  OAI210     u0930(.A0(men_men_n951_), .A1(men_men_n185_), .B0(men_men_n952_), .Y(men_men_n953_));
  AOI220     u0931(.A0(men_men_n953_), .A1(men_men_n488_), .B0(men_men_n950_), .B1(men_men_n71_), .Y(men_men_n954_));
  NA3        u0932(.A(men_men_n833_), .B(men_men_n388_), .C(i_6_), .Y(men_men_n955_));
  NA2        u0933(.A(men_men_n92_), .B(men_men_n44_), .Y(men_men_n956_));
  NO2        u0934(.A(men_men_n73_), .B(men_men_n770_), .Y(men_men_n957_));
  AOI220     u0935(.A0(men_men_n957_), .A1(men_men_n956_), .B0(men_men_n171_), .B1(men_men_n618_), .Y(men_men_n958_));
  AOI210     u0936(.A0(men_men_n958_), .A1(men_men_n955_), .B0(men_men_n47_), .Y(men_men_n959_));
  NO3        u0937(.A(men_men_n611_), .B(men_men_n360_), .C(men_men_n24_), .Y(men_men_n960_));
  AOI210     u0938(.A0(men_men_n721_), .A1(men_men_n567_), .B0(men_men_n960_), .Y(men_men_n961_));
  NAi21      u0939(.An(i_9_), .B(i_5_), .Y(men_men_n962_));
  NO2        u0940(.A(men_men_n962_), .B(men_men_n412_), .Y(men_men_n963_));
  NO2        u0941(.A(men_men_n623_), .B(men_men_n101_), .Y(men_men_n964_));
  AOI220     u0942(.A0(men_men_n964_), .A1(i_0_), .B0(men_men_n963_), .B1(men_men_n646_), .Y(men_men_n965_));
  OAI220     u0943(.A0(men_men_n965_), .A1(men_men_n84_), .B0(men_men_n961_), .B1(men_men_n169_), .Y(men_men_n966_));
  NO3        u0944(.A(men_men_n966_), .B(men_men_n959_), .C(men_men_n537_), .Y(men_men_n967_));
  NA4        u0945(.A(men_men_n967_), .B(men_men_n954_), .C(men_men_n948_), .D(men_men_n945_), .Y(men_men_n968_));
  NO3        u0946(.A(men_men_n968_), .B(men_men_n941_), .C(men_men_n914_), .Y(men_men_n969_));
  NO2        u0947(.A(men_men_n885_), .B(men_men_n747_), .Y(men_men_n970_));
  NA2        u0948(.A(men_men_n71_), .B(men_men_n44_), .Y(men_men_n971_));
  NA2        u0949(.A(men_men_n905_), .B(men_men_n971_), .Y(men_men_n972_));
  NO3        u0950(.A(men_men_n101_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n973_));
  AO220      u0951(.A0(men_men_n973_), .A1(men_men_n972_), .B0(men_men_n970_), .B1(men_men_n171_), .Y(men_men_n974_));
  AOI210     u0952(.A0(men_men_n814_), .A1(men_men_n707_), .B0(men_men_n928_), .Y(men_men_n975_));
  AOI210     u0953(.A0(men_men_n974_), .A1(men_men_n349_), .B0(men_men_n975_), .Y(men_men_n976_));
  NA2        u0954(.A(men_men_n758_), .B(men_men_n141_), .Y(men_men_n977_));
  INV        u0955(.A(men_men_n977_), .Y(men_men_n978_));
  NA3        u0956(.A(men_men_n978_), .B(men_men_n695_), .C(men_men_n71_), .Y(men_men_n979_));
  NO2        u0957(.A(men_men_n829_), .B(men_men_n412_), .Y(men_men_n980_));
  NA3        u0958(.A(men_men_n859_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n981_));
  NA2        u0959(.A(men_men_n860_), .B(i_9_), .Y(men_men_n982_));
  AOI210     u0960(.A0(men_men_n981_), .A1(men_men_n512_), .B0(men_men_n982_), .Y(men_men_n983_));
  OAI210     u0961(.A0(men_men_n244_), .A1(i_9_), .B0(men_men_n230_), .Y(men_men_n984_));
  AOI210     u0962(.A0(men_men_n984_), .A1(men_men_n895_), .B0(men_men_n149_), .Y(men_men_n985_));
  NO3        u0963(.A(men_men_n985_), .B(men_men_n983_), .C(men_men_n980_), .Y(men_men_n986_));
  NA3        u0964(.A(men_men_n986_), .B(men_men_n979_), .C(men_men_n976_), .Y(men_men_n987_));
  NA2        u0965(.A(men_men_n943_), .B(men_men_n378_), .Y(men_men_n988_));
  AOI210     u0966(.A0(men_men_n304_), .A1(men_men_n158_), .B0(men_men_n988_), .Y(men_men_n989_));
  NA2        u0967(.A(men_men_n39_), .B(men_men_n44_), .Y(men_men_n990_));
  NA2        u0968(.A(men_men_n919_), .B(men_men_n502_), .Y(men_men_n991_));
  AOI210     u0969(.A0(men_men_n990_), .A1(men_men_n158_), .B0(men_men_n991_), .Y(men_men_n992_));
  NO2        u0970(.A(men_men_n992_), .B(men_men_n989_), .Y(men_men_n993_));
  NO3        u0971(.A(men_men_n905_), .B(men_men_n877_), .C(men_men_n188_), .Y(men_men_n994_));
  AOI220     u0972(.A0(men_men_n994_), .A1(i_11_), .B0(men_men_n589_), .B1(men_men_n73_), .Y(men_men_n995_));
  NO3        u0973(.A(men_men_n209_), .B(men_men_n389_), .C(i_0_), .Y(men_men_n996_));
  OAI210     u0974(.A0(men_men_n996_), .A1(men_men_n74_), .B0(i_13_), .Y(men_men_n997_));
  INV        u0975(.A(men_men_n217_), .Y(men_men_n998_));
  OAI220     u0976(.A0(men_men_n548_), .A1(men_men_n134_), .B0(men_men_n1098_), .B1(men_men_n640_), .Y(men_men_n999_));
  NA3        u0977(.A(men_men_n999_), .B(men_men_n404_), .C(men_men_n998_), .Y(men_men_n1000_));
  NA4        u0978(.A(men_men_n1000_), .B(men_men_n997_), .C(men_men_n995_), .D(men_men_n993_), .Y(men_men_n1001_));
  NO2        u0979(.A(men_men_n242_), .B(men_men_n92_), .Y(men_men_n1002_));
  AOI210     u0980(.A0(men_men_n1002_), .A1(men_men_n970_), .B0(men_men_n104_), .Y(men_men_n1003_));
  AOI220     u0981(.A0(men_men_n933_), .A1(men_men_n502_), .B0(men_men_n859_), .B1(men_men_n159_), .Y(men_men_n1004_));
  NA2        u0982(.A(men_men_n352_), .B(men_men_n173_), .Y(men_men_n1005_));
  OA220      u0983(.A0(men_men_n1005_), .A1(men_men_n1004_), .B0(men_men_n1003_), .B1(i_5_), .Y(men_men_n1006_));
  AOI210     u0984(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n172_), .Y(men_men_n1007_));
  NA2        u0985(.A(men_men_n1007_), .B(men_men_n947_), .Y(men_men_n1008_));
  NA3        u0986(.A(men_men_n637_), .B(men_men_n183_), .C(men_men_n82_), .Y(men_men_n1009_));
  NA2        u0987(.A(men_men_n1009_), .B(men_men_n565_), .Y(men_men_n1010_));
  NO3        u0988(.A(men_men_n869_), .B(men_men_n53_), .C(men_men_n48_), .Y(men_men_n1011_));
  NO3        u0989(.A(men_men_n1096_), .B(men_men_n1011_), .C(men_men_n1010_), .Y(men_men_n1012_));
  NA3        u0990(.A(men_men_n396_), .B(men_men_n168_), .C(men_men_n167_), .Y(men_men_n1013_));
  NA3        u0991(.A(men_men_n919_), .B(men_men_n293_), .C(men_men_n230_), .Y(men_men_n1014_));
  NA2        u0992(.A(men_men_n1014_), .B(men_men_n1013_), .Y(men_men_n1015_));
  NA3        u0993(.A(men_men_n396_), .B(men_men_n337_), .C(men_men_n221_), .Y(men_men_n1016_));
  OAI210     u0994(.A0(men_men_n873_), .A1(men_men_n671_), .B0(men_men_n1016_), .Y(men_men_n1017_));
  NOi31      u0995(.An(men_men_n395_), .B(men_men_n971_), .C(men_men_n239_), .Y(men_men_n1018_));
  NO3        u0996(.A(men_men_n916_), .B(men_men_n217_), .C(men_men_n188_), .Y(men_men_n1019_));
  NO4        u0997(.A(men_men_n1019_), .B(men_men_n1018_), .C(men_men_n1017_), .D(men_men_n1015_), .Y(men_men_n1020_));
  NA4        u0998(.A(men_men_n1020_), .B(men_men_n1012_), .C(men_men_n1008_), .D(men_men_n1006_), .Y(men_men_n1021_));
  AOI210     u0999(.A0(men_men_n588_), .A1(men_men_n547_), .B0(men_men_n639_), .Y(men_men_n1022_));
  NO3        u1000(.A(men_men_n1022_), .B(men_men_n579_), .C(men_men_n346_), .Y(men_men_n1023_));
  NO2        u1001(.A(men_men_n84_), .B(i_5_), .Y(men_men_n1024_));
  NA3        u1002(.A(men_men_n860_), .B(men_men_n105_), .C(men_men_n119_), .Y(men_men_n1025_));
  INV        u1003(.A(men_men_n1025_), .Y(men_men_n1026_));
  AOI210     u1004(.A0(men_men_n1026_), .A1(men_men_n1024_), .B0(men_men_n1023_), .Y(men_men_n1027_));
  NA3        u1005(.A(men_men_n308_), .B(i_5_), .C(men_men_n191_), .Y(men_men_n1028_));
  NAi31      u1006(.An(men_men_n241_), .B(men_men_n1028_), .C(men_men_n242_), .Y(men_men_n1029_));
  NO4        u1007(.A(men_men_n239_), .B(men_men_n209_), .C(i_0_), .D(i_12_), .Y(men_men_n1030_));
  AOI220     u1008(.A0(men_men_n1030_), .A1(men_men_n1029_), .B0(men_men_n808_), .B1(men_men_n173_), .Y(men_men_n1031_));
  AN2        u1009(.A(men_men_n905_), .B(men_men_n149_), .Y(men_men_n1032_));
  NO4        u1010(.A(men_men_n1032_), .B(i_12_), .C(men_men_n671_), .D(men_men_n126_), .Y(men_men_n1033_));
  NA2        u1011(.A(men_men_n1033_), .B(men_men_n217_), .Y(men_men_n1034_));
  NA3        u1012(.A(men_men_n96_), .B(men_men_n593_), .C(i_11_), .Y(men_men_n1035_));
  NO2        u1013(.A(men_men_n1035_), .B(men_men_n151_), .Y(men_men_n1036_));
  NA2        u1014(.A(men_men_n933_), .B(men_men_n485_), .Y(men_men_n1037_));
  NA2        u1015(.A(men_men_n63_), .B(men_men_n98_), .Y(men_men_n1038_));
  OAI220     u1016(.A0(men_men_n1038_), .A1(men_men_n1028_), .B0(men_men_n1037_), .B1(men_men_n696_), .Y(men_men_n1039_));
  AOI210     u1017(.A0(men_men_n1039_), .A1(men_men_n921_), .B0(men_men_n1036_), .Y(men_men_n1040_));
  NA4        u1018(.A(men_men_n1040_), .B(men_men_n1034_), .C(men_men_n1031_), .D(men_men_n1027_), .Y(men_men_n1041_));
  NO4        u1019(.A(men_men_n1041_), .B(men_men_n1021_), .C(men_men_n1001_), .D(men_men_n987_), .Y(men_men_n1042_));
  OAI210     u1020(.A0(men_men_n832_), .A1(men_men_n827_), .B0(men_men_n37_), .Y(men_men_n1043_));
  NA3        u1021(.A(men_men_n927_), .B(men_men_n373_), .C(i_5_), .Y(men_men_n1044_));
  NA3        u1022(.A(men_men_n1044_), .B(men_men_n1043_), .C(men_men_n635_), .Y(men_men_n1045_));
  NA2        u1023(.A(men_men_n1045_), .B(men_men_n205_), .Y(men_men_n1046_));
  AN2        u1024(.A(men_men_n716_), .B(men_men_n374_), .Y(men_men_n1047_));
  NA2        u1025(.A(men_men_n184_), .B(men_men_n186_), .Y(men_men_n1048_));
  AO210      u1026(.A0(men_men_n1047_), .A1(men_men_n33_), .B0(men_men_n1048_), .Y(men_men_n1049_));
  OAI210     u1027(.A0(men_men_n639_), .A1(men_men_n637_), .B0(men_men_n318_), .Y(men_men_n1050_));
  NAi31      u1028(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1051_));
  AOI210     u1029(.A0(men_men_n112_), .A1(men_men_n68_), .B0(men_men_n1051_), .Y(men_men_n1052_));
  NO2        u1030(.A(men_men_n1052_), .B(men_men_n668_), .Y(men_men_n1053_));
  NA3        u1031(.A(men_men_n1053_), .B(men_men_n1050_), .C(men_men_n1049_), .Y(men_men_n1054_));
  NO2        u1032(.A(men_men_n475_), .B(men_men_n270_), .Y(men_men_n1055_));
  NO4        u1033(.A(men_men_n232_), .B(men_men_n140_), .C(men_men_n699_), .D(men_men_n37_), .Y(men_men_n1056_));
  NO3        u1034(.A(men_men_n1056_), .B(men_men_n1055_), .C(men_men_n897_), .Y(men_men_n1057_));
  OAI210     u1035(.A0(men_men_n1035_), .A1(men_men_n143_), .B0(men_men_n1057_), .Y(men_men_n1058_));
  AOI210     u1036(.A0(men_men_n1054_), .A1(men_men_n48_), .B0(men_men_n1058_), .Y(men_men_n1059_));
  AOI210     u1037(.A0(men_men_n1059_), .A1(men_men_n1046_), .B0(men_men_n71_), .Y(men_men_n1060_));
  NO2        u1038(.A(men_men_n586_), .B(men_men_n385_), .Y(men_men_n1061_));
  NO2        u1039(.A(men_men_n1061_), .B(men_men_n775_), .Y(men_men_n1062_));
  OAI210     u1040(.A0(men_men_n78_), .A1(men_men_n53_), .B0(men_men_n103_), .Y(men_men_n1063_));
  NA2        u1041(.A(men_men_n1063_), .B(men_men_n74_), .Y(men_men_n1064_));
  AOI210     u1042(.A0(men_men_n1007_), .A1(men_men_n919_), .B0(men_men_n934_), .Y(men_men_n1065_));
  AOI210     u1043(.A0(men_men_n1065_), .A1(men_men_n1064_), .B0(men_men_n699_), .Y(men_men_n1066_));
  NA2        u1044(.A(men_men_n264_), .B(men_men_n56_), .Y(men_men_n1067_));
  AOI220     u1045(.A0(men_men_n1067_), .A1(men_men_n74_), .B0(men_men_n347_), .B1(men_men_n256_), .Y(men_men_n1068_));
  NO2        u1046(.A(men_men_n1068_), .B(men_men_n236_), .Y(men_men_n1069_));
  NA3        u1047(.A(men_men_n94_), .B(men_men_n310_), .C(men_men_n31_), .Y(men_men_n1070_));
  INV        u1048(.A(men_men_n1070_), .Y(men_men_n1071_));
  NO3        u1049(.A(men_men_n1071_), .B(men_men_n1069_), .C(men_men_n1066_), .Y(men_men_n1072_));
  OAI210     u1050(.A0(men_men_n272_), .A1(men_men_n154_), .B0(men_men_n87_), .Y(men_men_n1073_));
  NA3        u1051(.A(men_men_n778_), .B(men_men_n293_), .C(men_men_n78_), .Y(men_men_n1074_));
  AOI210     u1052(.A0(men_men_n1074_), .A1(men_men_n1073_), .B0(i_11_), .Y(men_men_n1075_));
  NA2        u1053(.A(men_men_n630_), .B(men_men_n214_), .Y(men_men_n1076_));
  OAI210     u1054(.A0(men_men_n1076_), .A1(men_men_n927_), .B0(men_men_n205_), .Y(men_men_n1077_));
  NA2        u1055(.A(men_men_n160_), .B(i_5_), .Y(men_men_n1078_));
  AOI210     u1056(.A0(men_men_n1077_), .A1(men_men_n791_), .B0(men_men_n1078_), .Y(men_men_n1079_));
  NO3        u1057(.A(men_men_n58_), .B(men_men_n57_), .C(i_4_), .Y(men_men_n1080_));
  OAI210     u1058(.A0(men_men_n938_), .A1(men_men_n310_), .B0(men_men_n1080_), .Y(men_men_n1081_));
  NO2        u1059(.A(men_men_n1081_), .B(men_men_n747_), .Y(men_men_n1082_));
  NO4        u1060(.A(men_men_n962_), .B(men_men_n490_), .C(men_men_n253_), .D(men_men_n252_), .Y(men_men_n1083_));
  NO2        u1061(.A(men_men_n1083_), .B(men_men_n583_), .Y(men_men_n1084_));
  INV        u1062(.A(men_men_n366_), .Y(men_men_n1085_));
  AOI210     u1063(.A0(men_men_n1085_), .A1(men_men_n1084_), .B0(men_men_n40_), .Y(men_men_n1086_));
  NO4        u1064(.A(men_men_n1086_), .B(men_men_n1082_), .C(men_men_n1079_), .D(men_men_n1075_), .Y(men_men_n1087_));
  OAI210     u1065(.A0(men_men_n1072_), .A1(i_4_), .B0(men_men_n1087_), .Y(men_men_n1088_));
  NO3        u1066(.A(men_men_n1088_), .B(men_men_n1062_), .C(men_men_n1060_), .Y(men_men_n1089_));
  NA4        u1067(.A(men_men_n1089_), .B(men_men_n1042_), .C(men_men_n969_), .D(men_men_n884_), .Y(men4));
  INV        u1068(.A(men_men_n720_), .Y(men_men_n1093_));
  INV        u1069(.A(i_2_), .Y(men_men_n1094_));
  INV        u1070(.A(i_5_), .Y(men_men_n1095_));
  INV        u1071(.A(men_men_n500_), .Y(men_men_n1096_));
  INV        u1072(.A(i_3_), .Y(men_men_n1097_));
  INV        u1073(.A(i_6_), .Y(men_men_n1098_));
  INV        u1074(.A(i_1_), .Y(men_men_n1099_));
  INV        u1075(.A(i_4_), .Y(men_men_n1100_));
  INV        u1076(.A(men_men_n369_), .Y(men_men_n1101_));
  INV        u1077(.A(men_men_n139_), .Y(men_men_n1102_));
  INV        u1078(.A(men_men_n833_), .Y(men_men_n1103_));
  INV        u1079(.A(men_men_n196_), .Y(men_men_n1104_));
  INV        u1080(.A(men_men_n109_), .Y(men_men_n1105_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule