library verilog;
use verilog.vl_types.all;
entity testevirg_vlg_vec_tst is
end testevirg_vlg_vec_tst;
