// Benchmark "top" written by ABC on Thu Jun 20 14:00:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n140_, new_new_n141_, new_new_n142_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1072_, new_new_n1073_, new_new_n1074_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(zz01));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  OAI210     g0034(.A0(new_new_n56_), .A1(new_new_n53_), .B0(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  NO2        g0065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  OAI210     g0067(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n89_), .Y(new_new_n90_));
  NAi21      g0068(.An(i_6_), .B(i_10_), .Y(new_new_n91_));
  NA2        g0069(.A(i_6_), .B(i_9_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n92_), .A1(new_new_n91_), .B0(new_new_n64_), .Y(new_new_n93_));
  NA2        g0071(.A(i_2_), .B(i_6_), .Y(new_new_n94_));
  NO3        g0072(.A(new_new_n94_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n95_));
  NO2        g0073(.A(new_new_n95_), .B(new_new_n93_), .Y(new_new_n96_));
  AOI210     g0074(.A0(new_new_n96_), .A1(new_new_n90_), .B0(new_new_n81_), .Y(new_new_n97_));
  AN3        g0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g0076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g0077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NOi21      g0078(.An(new_new_n100_), .B(new_new_n99_), .Y(new_new_n101_));
  AOI220     g0079(.A0(new_new_n101_), .A1(new_new_n63_), .B0(new_new_n98_), .B1(new_new_n32_), .Y(new_new_n102_));
  INV        g0080(.A(i_7_), .Y(new_new_n103_));
  NA2        g0081(.A(new_new_n47_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g0082(.A(i_0_), .B(i_5_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(new_new_n87_), .Y(new_new_n106_));
  NA2        g0084(.A(i_12_), .B(i_3_), .Y(new_new_n107_));
  INV        g0085(.A(new_new_n107_), .Y(new_new_n108_));
  NA3        g0086(.A(new_new_n108_), .B(new_new_n106_), .C(new_new_n104_), .Y(new_new_n109_));
  NAi21      g0087(.An(i_7_), .B(i_11_), .Y(new_new_n110_));
  AN2        g0088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g0089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g0090(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n113_));
  NO2        g0091(.A(i_8_), .B(new_new_n103_), .Y(new_new_n114_));
  NO3        g0092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g0093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NO2        g0094(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n117_));
  NA2        g0095(.A(new_new_n117_), .B(i_0_), .Y(new_new_n118_));
  NA2        g0096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  OAI210     g0097(.A0(new_new_n118_), .A1(new_new_n116_), .B0(new_new_n119_), .Y(new_new_n120_));
  NO2        g0098(.A(new_new_n120_), .B(new_new_n115_), .Y(new_new_n121_));
  NA3        g0099(.A(new_new_n121_), .B(new_new_n109_), .C(new_new_n102_), .Y(new_new_n122_));
  NOi21      g0100(.An(i_1_), .B(i_5_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n123_), .B(i_11_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n125_));
  NA2        g0103(.A(i_7_), .B(new_new_n25_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(new_new_n125_), .Y(new_new_n127_));
  NO2        g0105(.A(new_new_n127_), .B(new_new_n47_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n92_), .B(new_new_n91_), .Y(new_new_n129_));
  NAi21      g0107(.An(i_3_), .B(i_8_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n130_), .B(new_new_n63_), .Y(new_new_n131_));
  NOi31      g0109(.An(new_new_n131_), .B(new_new_n129_), .C(new_new_n128_), .Y(new_new_n132_));
  NO2        g0110(.A(i_1_), .B(new_new_n87_), .Y(new_new_n133_));
  NO2        g0111(.A(i_6_), .B(i_5_), .Y(new_new_n134_));
  NA2        g0112(.A(new_new_n134_), .B(i_3_), .Y(new_new_n135_));
  AO210      g0113(.A0(new_new_n135_), .A1(new_new_n48_), .B0(new_new_n133_), .Y(new_new_n136_));
  OAI220     g0114(.A0(new_new_n136_), .A1(new_new_n110_), .B0(new_new_n132_), .B1(new_new_n124_), .Y(new_new_n137_));
  NO3        g0115(.A(new_new_n137_), .B(new_new_n122_), .C(new_new_n97_), .Y(new_new_n138_));
  NA3        g0116(.A(new_new_n138_), .B(new_new_n80_), .C(new_new_n57_), .Y(zz02));
  NO2        g0117(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n140_));
  NA2        g0118(.A(i_6_), .B(new_new_n25_), .Y(new_new_n141_));
  NA2        g0119(.A(new_new_n141_), .B(new_new_n140_), .Y(new_new_n142_));
  NA4        g0120(.A(new_new_n142_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(zz00));
  AN2        g0121(.A(i_8_), .B(i_7_), .Y(new_new_n144_));
  NA2        g0122(.A(new_new_n144_), .B(i_6_), .Y(new_new_n145_));
  NO2        g0123(.A(i_12_), .B(i_13_), .Y(new_new_n146_));
  NAi21      g0124(.An(i_5_), .B(i_11_), .Y(new_new_n147_));
  NOi21      g0125(.An(new_new_n146_), .B(new_new_n147_), .Y(new_new_n148_));
  NO2        g0126(.A(i_0_), .B(i_1_), .Y(new_new_n149_));
  NA2        g0127(.A(i_2_), .B(i_3_), .Y(new_new_n150_));
  NO2        g0128(.A(new_new_n150_), .B(i_4_), .Y(new_new_n151_));
  NA3        g0129(.A(new_new_n151_), .B(new_new_n149_), .C(new_new_n148_), .Y(new_new_n152_));
  AN2        g0130(.A(new_new_n146_), .B(new_new_n84_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n153_), .B(new_new_n27_), .Y(new_new_n154_));
  NA2        g0132(.A(i_1_), .B(i_5_), .Y(new_new_n155_));
  NO2        g0133(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n156_));
  NA2        g0134(.A(new_new_n156_), .B(new_new_n36_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n155_), .C(new_new_n154_), .Y(new_new_n158_));
  OR2        g0136(.A(i_0_), .B(i_1_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n159_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n160_));
  NAi32      g0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n161_));
  NAi21      g0139(.An(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  NOi21      g0140(.An(i_4_), .B(i_10_), .Y(new_new_n163_));
  NA2        g0141(.A(new_new_n163_), .B(new_new_n40_), .Y(new_new_n164_));
  NO2        g0142(.A(i_3_), .B(i_5_), .Y(new_new_n165_));
  NO3        g0143(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n166_));
  NA2        g0144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  OAI210     g0145(.A0(new_new_n167_), .A1(new_new_n164_), .B0(new_new_n162_), .Y(new_new_n168_));
  NO2        g0146(.A(new_new_n168_), .B(new_new_n158_), .Y(new_new_n169_));
  AOI210     g0147(.A0(new_new_n169_), .A1(new_new_n152_), .B0(new_new_n145_), .Y(new_new_n170_));
  NA3        g0148(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n171_));
  NA2        g0149(.A(i_3_), .B(new_new_n49_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_4_), .B(i_9_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_11_), .B(i_13_), .Y(new_new_n174_));
  NA2        g0152(.A(new_new_n174_), .B(new_new_n173_), .Y(new_new_n175_));
  OR2        g0153(.A(new_new_n175_), .B(new_new_n172_), .Y(new_new_n176_));
  NO2        g0154(.A(i_4_), .B(i_5_), .Y(new_new_n177_));
  NAi21      g0155(.An(i_12_), .B(i_11_), .Y(new_new_n178_));
  NO2        g0156(.A(new_new_n178_), .B(i_13_), .Y(new_new_n179_));
  NA3        g0157(.A(new_new_n179_), .B(new_new_n177_), .C(new_new_n84_), .Y(new_new_n180_));
  AOI210     g0158(.A0(new_new_n180_), .A1(new_new_n176_), .B0(new_new_n171_), .Y(new_new_n181_));
  NO2        g0159(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n182_), .B(new_new_n47_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n36_), .B(i_5_), .Y(new_new_n184_));
  NAi31      g0162(.An(new_new_n184_), .B(new_new_n153_), .C(i_11_), .Y(new_new_n185_));
  NA2        g0163(.A(i_3_), .B(i_5_), .Y(new_new_n186_));
  OR2        g0164(.A(new_new_n186_), .B(new_new_n175_), .Y(new_new_n187_));
  AOI210     g0165(.A0(new_new_n187_), .A1(new_new_n185_), .B0(new_new_n183_), .Y(new_new_n188_));
  NO2        g0166(.A(new_new_n74_), .B(i_5_), .Y(new_new_n189_));
  NO2        g0167(.A(i_13_), .B(i_10_), .Y(new_new_n190_));
  NA3        g0168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n45_), .Y(new_new_n191_));
  NO2        g0169(.A(i_2_), .B(i_1_), .Y(new_new_n192_));
  NA2        g0170(.A(new_new_n192_), .B(i_3_), .Y(new_new_n193_));
  NAi21      g0171(.An(i_4_), .B(i_12_), .Y(new_new_n194_));
  NO4        g0172(.A(new_new_n194_), .B(new_new_n193_), .C(new_new_n191_), .D(new_new_n25_), .Y(new_new_n195_));
  NO3        g0173(.A(new_new_n195_), .B(new_new_n188_), .C(new_new_n181_), .Y(new_new_n196_));
  INV        g0174(.A(i_8_), .Y(new_new_n197_));
  NO2        g0175(.A(new_new_n197_), .B(i_7_), .Y(new_new_n198_));
  NA2        g0176(.A(new_new_n198_), .B(i_6_), .Y(new_new_n199_));
  NO3        g0177(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n200_));
  NA2        g0178(.A(new_new_n200_), .B(new_new_n114_), .Y(new_new_n201_));
  NO3        g0179(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n202_));
  NA3        g0180(.A(new_new_n202_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n203_));
  NO3        g0181(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n204_));
  OAI210     g0182(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n204_), .Y(new_new_n205_));
  AOI210     g0183(.A0(new_new_n205_), .A1(new_new_n203_), .B0(new_new_n201_), .Y(new_new_n206_));
  NO2        g0184(.A(i_3_), .B(i_8_), .Y(new_new_n207_));
  NO3        g0185(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n208_));
  NO2        g0186(.A(new_new_n105_), .B(new_new_n59_), .Y(new_new_n209_));
  NO2        g0187(.A(i_13_), .B(i_9_), .Y(new_new_n210_));
  NA3        g0188(.A(new_new_n210_), .B(i_6_), .C(new_new_n197_), .Y(new_new_n211_));
  NAi21      g0189(.An(i_12_), .B(i_3_), .Y(new_new_n212_));
  NO2        g0190(.A(new_new_n45_), .B(i_5_), .Y(new_new_n213_));
  NO3        g0191(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n214_));
  NA3        g0192(.A(new_new_n214_), .B(new_new_n213_), .C(i_10_), .Y(new_new_n215_));
  NO2        g0193(.A(new_new_n215_), .B(new_new_n211_), .Y(new_new_n216_));
  AOI210     g0194(.A0(new_new_n216_), .A1(i_7_), .B0(new_new_n206_), .Y(new_new_n217_));
  OAI220     g0195(.A0(new_new_n217_), .A1(i_4_), .B0(new_new_n199_), .B1(new_new_n196_), .Y(new_new_n218_));
  NAi21      g0196(.An(i_12_), .B(i_7_), .Y(new_new_n219_));
  NA3        g0197(.A(i_13_), .B(new_new_n197_), .C(i_10_), .Y(new_new_n220_));
  NA2        g0198(.A(i_0_), .B(i_5_), .Y(new_new_n221_));
  NAi31      g0199(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n36_), .B(i_13_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n225_));
  NA3        g0203(.A(new_new_n225_), .B(new_new_n224_), .C(new_new_n223_), .Y(new_new_n226_));
  INV        g0204(.A(i_13_), .Y(new_new_n227_));
  NO2        g0205(.A(i_12_), .B(new_new_n227_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n226_), .B(new_new_n222_), .Y(new_new_n229_));
  NA2        g0207(.A(new_new_n229_), .B(new_new_n144_), .Y(new_new_n230_));
  NO2        g0208(.A(i_12_), .B(new_new_n37_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n186_), .B(i_4_), .Y(new_new_n232_));
  NA2        g0210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  OR2        g0211(.A(i_8_), .B(i_7_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n234_), .B(new_new_n87_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n54_), .B(i_1_), .Y(new_new_n236_));
  NA2        g0214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  INV        g0215(.A(i_12_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n45_), .B(new_new_n238_), .Y(new_new_n239_));
  NO3        g0217(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n240_));
  NA2        g0218(.A(i_2_), .B(i_1_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n237_), .B(new_new_n233_), .Y(new_new_n242_));
  NO3        g0220(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n243_));
  NAi21      g0221(.An(i_4_), .B(i_3_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n244_), .B(new_new_n76_), .Y(new_new_n245_));
  NO2        g0223(.A(i_0_), .B(i_6_), .Y(new_new_n246_));
  NOi41      g0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n247_));
  NA2        g0225(.A(new_new_n247_), .B(new_new_n246_), .Y(new_new_n248_));
  NO2        g0226(.A(new_new_n241_), .B(new_new_n186_), .Y(new_new_n249_));
  NAi21      g0227(.An(new_new_n248_), .B(new_new_n249_), .Y(new_new_n250_));
  INV        g0228(.A(new_new_n250_), .Y(new_new_n251_));
  AOI220     g0229(.A0(new_new_n251_), .A1(new_new_n40_), .B0(new_new_n242_), .B1(new_new_n210_), .Y(new_new_n252_));
  NO2        g0230(.A(i_11_), .B(new_new_n227_), .Y(new_new_n253_));
  NOi21      g0231(.An(i_1_), .B(i_6_), .Y(new_new_n254_));
  NAi21      g0232(.An(i_3_), .B(i_7_), .Y(new_new_n255_));
  NA2        g0233(.A(new_new_n238_), .B(i_9_), .Y(new_new_n256_));
  OR4        g0234(.A(new_new_n256_), .B(new_new_n255_), .C(new_new_n254_), .D(new_new_n189_), .Y(new_new_n257_));
  NO2        g0235(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n258_));
  NO2        g0236(.A(i_12_), .B(i_3_), .Y(new_new_n259_));
  NA2        g0237(.A(new_new_n74_), .B(i_5_), .Y(new_new_n260_));
  NA2        g0238(.A(i_3_), .B(i_9_), .Y(new_new_n261_));
  NAi21      g0239(.An(i_7_), .B(i_10_), .Y(new_new_n262_));
  NO2        g0240(.A(new_new_n262_), .B(new_new_n261_), .Y(new_new_n263_));
  NA3        g0241(.A(new_new_n263_), .B(new_new_n260_), .C(new_new_n65_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n264_), .B(new_new_n257_), .Y(new_new_n265_));
  NA3        g0243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n266_));
  INV        g0244(.A(new_new_n145_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n238_), .B(i_13_), .Y(new_new_n268_));
  NO2        g0246(.A(new_new_n268_), .B(new_new_n76_), .Y(new_new_n269_));
  AOI220     g0247(.A0(new_new_n269_), .A1(new_new_n267_), .B0(new_new_n265_), .B1(new_new_n253_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n234_), .B(new_new_n37_), .Y(new_new_n271_));
  NA2        g0249(.A(i_12_), .B(i_6_), .Y(new_new_n272_));
  OR2        g0250(.A(i_13_), .B(i_9_), .Y(new_new_n273_));
  NO3        g0251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n49_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n244_), .B(i_2_), .Y(new_new_n275_));
  NA2        g0253(.A(new_new_n253_), .B(i_9_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n156_), .B(new_new_n64_), .Y(new_new_n277_));
  NO3        g0255(.A(i_11_), .B(new_new_n227_), .C(new_new_n25_), .Y(new_new_n278_));
  NO2        g0256(.A(new_new_n255_), .B(i_8_), .Y(new_new_n279_));
  NO2        g0257(.A(i_6_), .B(new_new_n49_), .Y(new_new_n280_));
  NA3        g0258(.A(new_new_n280_), .B(new_new_n279_), .C(new_new_n278_), .Y(new_new_n281_));
  NO3        g0259(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n282_));
  NA3        g0260(.A(new_new_n282_), .B(new_new_n271_), .C(new_new_n228_), .Y(new_new_n283_));
  AOI210     g0261(.A0(new_new_n283_), .A1(new_new_n281_), .B0(new_new_n277_), .Y(new_new_n284_));
  INV        g0262(.A(new_new_n284_), .Y(new_new_n285_));
  NA4        g0263(.A(new_new_n285_), .B(new_new_n270_), .C(new_new_n252_), .D(new_new_n230_), .Y(new_new_n286_));
  NO3        g0264(.A(i_12_), .B(new_new_n227_), .C(new_new_n37_), .Y(new_new_n287_));
  INV        g0265(.A(new_new_n287_), .Y(new_new_n288_));
  NA2        g0266(.A(i_8_), .B(new_new_n103_), .Y(new_new_n289_));
  NOi21      g0267(.An(new_new_n165_), .B(new_new_n87_), .Y(new_new_n290_));
  NO3        g0268(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n291_));
  AOI220     g0269(.A0(new_new_n291_), .A1(new_new_n200_), .B0(new_new_n290_), .B1(new_new_n236_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n292_), .B(new_new_n289_), .Y(new_new_n293_));
  NO3        g0271(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n241_), .B(i_0_), .Y(new_new_n295_));
  AOI220     g0273(.A0(new_new_n295_), .A1(new_new_n198_), .B0(new_new_n294_), .B1(new_new_n144_), .Y(new_new_n296_));
  NA2        g0274(.A(new_new_n280_), .B(new_new_n26_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(new_new_n296_), .Y(new_new_n298_));
  NA2        g0276(.A(i_0_), .B(i_1_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n299_), .B(i_2_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n60_), .B(i_6_), .Y(new_new_n301_));
  NA3        g0279(.A(new_new_n301_), .B(new_new_n300_), .C(new_new_n165_), .Y(new_new_n302_));
  OAI210     g0280(.A0(new_new_n167_), .A1(new_new_n145_), .B0(new_new_n302_), .Y(new_new_n303_));
  NO3        g0281(.A(new_new_n303_), .B(new_new_n298_), .C(new_new_n293_), .Y(new_new_n304_));
  NO2        g0282(.A(i_3_), .B(i_10_), .Y(new_new_n305_));
  NA3        g0283(.A(new_new_n305_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n306_));
  NO2        g0284(.A(i_2_), .B(new_new_n103_), .Y(new_new_n307_));
  NA2        g0285(.A(i_1_), .B(new_new_n36_), .Y(new_new_n308_));
  NO2        g0286(.A(new_new_n308_), .B(i_8_), .Y(new_new_n309_));
  NA2        g0287(.A(new_new_n309_), .B(new_new_n307_), .Y(new_new_n310_));
  AN2        g0288(.A(i_3_), .B(i_10_), .Y(new_new_n311_));
  NA4        g0289(.A(new_new_n311_), .B(new_new_n202_), .C(new_new_n179_), .D(new_new_n177_), .Y(new_new_n312_));
  NO2        g0290(.A(i_5_), .B(new_new_n37_), .Y(new_new_n313_));
  NO2        g0291(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n314_));
  OR2        g0292(.A(new_new_n310_), .B(new_new_n306_), .Y(new_new_n315_));
  OAI220     g0293(.A0(new_new_n315_), .A1(i_6_), .B0(new_new_n304_), .B1(new_new_n288_), .Y(new_new_n316_));
  NO4        g0294(.A(new_new_n316_), .B(new_new_n286_), .C(new_new_n218_), .D(new_new_n170_), .Y(new_new_n317_));
  NO3        g0295(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n318_));
  NO2        g0296(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n319_));
  NA2        g0297(.A(new_new_n295_), .B(new_new_n319_), .Y(new_new_n320_));
  NO3        g0298(.A(i_6_), .B(new_new_n197_), .C(i_7_), .Y(new_new_n321_));
  NA2        g0299(.A(new_new_n321_), .B(new_new_n202_), .Y(new_new_n322_));
  AOI210     g0300(.A0(new_new_n322_), .A1(new_new_n320_), .B0(new_new_n172_), .Y(new_new_n323_));
  NO2        g0301(.A(i_2_), .B(i_3_), .Y(new_new_n324_));
  OR2        g0302(.A(i_0_), .B(i_5_), .Y(new_new_n325_));
  NA2        g0303(.A(new_new_n221_), .B(new_new_n325_), .Y(new_new_n326_));
  NA4        g0304(.A(new_new_n326_), .B(new_new_n235_), .C(new_new_n324_), .D(i_1_), .Y(new_new_n327_));
  NA3        g0305(.A(new_new_n295_), .B(new_new_n290_), .C(new_new_n114_), .Y(new_new_n328_));
  NAi21      g0306(.An(i_8_), .B(i_7_), .Y(new_new_n329_));
  NO2        g0307(.A(new_new_n329_), .B(i_6_), .Y(new_new_n330_));
  NO2        g0308(.A(new_new_n159_), .B(new_new_n47_), .Y(new_new_n331_));
  NA3        g0309(.A(new_new_n331_), .B(new_new_n330_), .C(new_new_n165_), .Y(new_new_n332_));
  NA3        g0310(.A(new_new_n332_), .B(new_new_n328_), .C(new_new_n327_), .Y(new_new_n333_));
  OAI210     g0311(.A0(new_new_n333_), .A1(new_new_n323_), .B0(i_4_), .Y(new_new_n334_));
  NO2        g0312(.A(i_12_), .B(i_10_), .Y(new_new_n335_));
  NOi21      g0313(.An(i_5_), .B(i_0_), .Y(new_new_n336_));
  AOI210     g0314(.A0(i_2_), .A1(new_new_n49_), .B0(new_new_n103_), .Y(new_new_n337_));
  NO4        g0315(.A(new_new_n337_), .B(new_new_n308_), .C(new_new_n336_), .D(new_new_n130_), .Y(new_new_n338_));
  NA4        g0316(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n339_));
  NA2        g0317(.A(new_new_n338_), .B(new_new_n335_), .Y(new_new_n340_));
  NO2        g0318(.A(i_6_), .B(i_8_), .Y(new_new_n341_));
  NOi21      g0319(.An(i_0_), .B(i_2_), .Y(new_new_n342_));
  AN2        g0320(.A(new_new_n342_), .B(new_new_n341_), .Y(new_new_n343_));
  NO2        g0321(.A(i_1_), .B(i_7_), .Y(new_new_n344_));
  AO220      g0322(.A0(new_new_n344_), .A1(new_new_n343_), .B0(new_new_n330_), .B1(new_new_n236_), .Y(new_new_n345_));
  NA3        g0323(.A(new_new_n345_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n346_));
  NA3        g0324(.A(new_new_n346_), .B(new_new_n340_), .C(new_new_n334_), .Y(new_new_n347_));
  NO3        g0325(.A(new_new_n234_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n348_));
  NO3        g0326(.A(new_new_n329_), .B(i_2_), .C(i_1_), .Y(new_new_n349_));
  OAI210     g0327(.A0(new_new_n349_), .A1(new_new_n348_), .B0(i_6_), .Y(new_new_n350_));
  NA3        g0328(.A(new_new_n254_), .B(new_new_n307_), .C(new_new_n197_), .Y(new_new_n351_));
  AOI210     g0329(.A0(new_new_n351_), .A1(new_new_n350_), .B0(new_new_n326_), .Y(new_new_n352_));
  NOi21      g0330(.An(new_new_n155_), .B(new_new_n106_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n353_), .B(new_new_n126_), .Y(new_new_n354_));
  OAI210     g0332(.A0(new_new_n354_), .A1(new_new_n352_), .B0(i_3_), .Y(new_new_n355_));
  INV        g0333(.A(new_new_n85_), .Y(new_new_n356_));
  NO2        g0334(.A(new_new_n299_), .B(new_new_n82_), .Y(new_new_n357_));
  NA2        g0335(.A(new_new_n357_), .B(new_new_n134_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n94_), .B(new_new_n197_), .Y(new_new_n359_));
  NA2        g0337(.A(new_new_n359_), .B(new_new_n64_), .Y(new_new_n360_));
  AOI210     g0338(.A0(new_new_n360_), .A1(new_new_n358_), .B0(new_new_n356_), .Y(new_new_n361_));
  NO2        g0339(.A(new_new_n197_), .B(i_9_), .Y(new_new_n362_));
  NA3        g0340(.A(new_new_n362_), .B(new_new_n209_), .C(new_new_n159_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n363_), .B(new_new_n47_), .Y(new_new_n364_));
  NO3        g0342(.A(new_new_n364_), .B(new_new_n361_), .C(new_new_n298_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n365_), .A1(new_new_n355_), .B0(new_new_n164_), .Y(new_new_n366_));
  AOI210     g0344(.A0(new_new_n347_), .A1(new_new_n318_), .B0(new_new_n366_), .Y(new_new_n367_));
  NOi32      g0345(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n368_));
  INV        g0346(.A(new_new_n368_), .Y(new_new_n369_));
  NAi21      g0347(.An(i_0_), .B(i_6_), .Y(new_new_n370_));
  NAi21      g0348(.An(i_1_), .B(i_5_), .Y(new_new_n371_));
  NA2        g0349(.A(new_new_n371_), .B(new_new_n370_), .Y(new_new_n372_));
  INV        g0350(.A(new_new_n248_), .Y(new_new_n373_));
  NAi41      g0351(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n374_));
  OAI220     g0352(.A0(new_new_n374_), .A1(new_new_n371_), .B0(new_new_n222_), .B1(new_new_n161_), .Y(new_new_n375_));
  AOI210     g0353(.A0(new_new_n374_), .A1(new_new_n161_), .B0(new_new_n159_), .Y(new_new_n376_));
  NOi32      g0354(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n377_));
  NAi21      g0355(.An(i_6_), .B(i_1_), .Y(new_new_n378_));
  NA3        g0356(.A(new_new_n378_), .B(new_new_n377_), .C(new_new_n47_), .Y(new_new_n379_));
  NO2        g0357(.A(new_new_n379_), .B(i_0_), .Y(new_new_n380_));
  OR3        g0358(.A(new_new_n380_), .B(new_new_n376_), .C(new_new_n375_), .Y(new_new_n381_));
  NO2        g0359(.A(i_1_), .B(new_new_n103_), .Y(new_new_n382_));
  NAi21      g0360(.An(i_3_), .B(i_4_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n383_), .B(i_9_), .Y(new_new_n384_));
  AN2        g0362(.A(i_6_), .B(i_7_), .Y(new_new_n385_));
  OAI210     g0363(.A0(new_new_n385_), .A1(new_new_n382_), .B0(new_new_n384_), .Y(new_new_n386_));
  NA2        g0364(.A(i_2_), .B(i_7_), .Y(new_new_n387_));
  NO2        g0365(.A(new_new_n383_), .B(i_10_), .Y(new_new_n388_));
  NA3        g0366(.A(new_new_n388_), .B(new_new_n387_), .C(new_new_n246_), .Y(new_new_n389_));
  AOI210     g0367(.A0(new_new_n389_), .A1(new_new_n386_), .B0(new_new_n189_), .Y(new_new_n390_));
  AOI210     g0368(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n391_));
  OAI210     g0369(.A0(new_new_n391_), .A1(new_new_n192_), .B0(new_new_n388_), .Y(new_new_n392_));
  AOI220     g0370(.A0(new_new_n388_), .A1(new_new_n344_), .B0(new_new_n240_), .B1(new_new_n192_), .Y(new_new_n393_));
  AOI210     g0371(.A0(new_new_n393_), .A1(new_new_n392_), .B0(i_5_), .Y(new_new_n394_));
  NO4        g0372(.A(new_new_n394_), .B(new_new_n390_), .C(new_new_n381_), .D(new_new_n373_), .Y(new_new_n395_));
  NO2        g0373(.A(new_new_n395_), .B(new_new_n369_), .Y(new_new_n396_));
  NO2        g0374(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n397_));
  AN2        g0375(.A(i_12_), .B(i_5_), .Y(new_new_n398_));
  NA2        g0376(.A(i_3_), .B(new_new_n398_), .Y(new_new_n399_));
  NO2        g0377(.A(i_11_), .B(i_6_), .Y(new_new_n400_));
  NA3        g0378(.A(new_new_n400_), .B(new_new_n331_), .C(new_new_n227_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n401_), .B(new_new_n399_), .Y(new_new_n402_));
  NO2        g0380(.A(new_new_n244_), .B(i_5_), .Y(new_new_n403_));
  NO2        g0381(.A(i_5_), .B(i_10_), .Y(new_new_n404_));
  AOI220     g0382(.A0(new_new_n404_), .A1(new_new_n275_), .B0(new_new_n403_), .B1(new_new_n202_), .Y(new_new_n405_));
  NA2        g0383(.A(new_new_n146_), .B(new_new_n46_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n406_), .B(new_new_n405_), .Y(new_new_n407_));
  OAI210     g0385(.A0(new_new_n407_), .A1(new_new_n402_), .B0(new_new_n397_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n409_));
  NO3        g0387(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n410_));
  NO2        g0388(.A(i_3_), .B(new_new_n103_), .Y(new_new_n411_));
  NO2        g0389(.A(i_11_), .B(i_12_), .Y(new_new_n412_));
  NA2        g0390(.A(new_new_n404_), .B(new_new_n238_), .Y(new_new_n413_));
  NA3        g0391(.A(new_new_n114_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n414_));
  OAI220     g0392(.A0(new_new_n414_), .A1(new_new_n222_), .B0(new_new_n413_), .B1(new_new_n339_), .Y(new_new_n415_));
  NAi21      g0393(.An(i_13_), .B(i_0_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n416_), .B(new_new_n241_), .Y(new_new_n417_));
  NA2        g0395(.A(new_new_n415_), .B(new_new_n417_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n418_), .B(new_new_n408_), .Y(new_new_n419_));
  NO3        g0397(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n420_));
  NO2        g0398(.A(i_0_), .B(i_11_), .Y(new_new_n421_));
  INV        g0399(.A(i_5_), .Y(new_new_n422_));
  AN2        g0400(.A(i_1_), .B(i_6_), .Y(new_new_n423_));
  NOi21      g0401(.An(i_2_), .B(i_12_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n424_), .B(new_new_n423_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n425_), .B(new_new_n422_), .Y(new_new_n426_));
  NA2        g0404(.A(new_new_n144_), .B(i_9_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n427_), .B(i_4_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n426_), .B(new_new_n428_), .Y(new_new_n429_));
  NAi21      g0407(.An(i_9_), .B(i_4_), .Y(new_new_n430_));
  OR2        g0408(.A(i_13_), .B(i_10_), .Y(new_new_n431_));
  NO3        g0409(.A(new_new_n431_), .B(new_new_n119_), .C(new_new_n430_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n175_), .B(new_new_n125_), .Y(new_new_n433_));
  OR2        g0411(.A(new_new_n220_), .B(new_new_n219_), .Y(new_new_n434_));
  NO2        g0412(.A(new_new_n103_), .B(new_new_n25_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n287_), .B(new_new_n435_), .Y(new_new_n436_));
  NA2        g0414(.A(new_new_n280_), .B(new_new_n214_), .Y(new_new_n437_));
  OAI220     g0415(.A0(new_new_n437_), .A1(new_new_n434_), .B0(new_new_n436_), .B1(new_new_n353_), .Y(new_new_n438_));
  INV        g0416(.A(new_new_n438_), .Y(new_new_n439_));
  AOI210     g0417(.A0(new_new_n439_), .A1(new_new_n429_), .B0(new_new_n26_), .Y(new_new_n440_));
  NA2        g0418(.A(new_new_n328_), .B(new_new_n327_), .Y(new_new_n441_));
  AOI220     g0419(.A0(new_new_n301_), .A1(new_new_n291_), .B0(new_new_n295_), .B1(new_new_n319_), .Y(new_new_n442_));
  NO2        g0420(.A(new_new_n442_), .B(new_new_n172_), .Y(new_new_n443_));
  NO2        g0421(.A(new_new_n186_), .B(new_new_n87_), .Y(new_new_n444_));
  AOI220     g0422(.A0(new_new_n444_), .A1(new_new_n300_), .B0(new_new_n282_), .B1(new_new_n214_), .Y(new_new_n445_));
  NO2        g0423(.A(new_new_n445_), .B(new_new_n289_), .Y(new_new_n446_));
  NO3        g0424(.A(new_new_n446_), .B(new_new_n443_), .C(new_new_n441_), .Y(new_new_n447_));
  NA2        g0425(.A(new_new_n200_), .B(new_new_n98_), .Y(new_new_n448_));
  NA3        g0426(.A(new_new_n331_), .B(new_new_n165_), .C(new_new_n87_), .Y(new_new_n449_));
  AOI210     g0427(.A0(new_new_n449_), .A1(new_new_n448_), .B0(new_new_n329_), .Y(new_new_n450_));
  NA2        g0428(.A(new_new_n197_), .B(i_10_), .Y(new_new_n451_));
  NA3        g0429(.A(new_new_n260_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n452_));
  NA2        g0430(.A(new_new_n301_), .B(new_new_n236_), .Y(new_new_n453_));
  OAI220     g0431(.A0(new_new_n453_), .A1(new_new_n186_), .B0(new_new_n452_), .B1(new_new_n451_), .Y(new_new_n454_));
  NO2        g0432(.A(i_3_), .B(new_new_n49_), .Y(new_new_n455_));
  NA3        g0433(.A(new_new_n344_), .B(new_new_n343_), .C(new_new_n455_), .Y(new_new_n456_));
  NA2        g0434(.A(new_new_n321_), .B(new_new_n326_), .Y(new_new_n457_));
  OAI210     g0435(.A0(new_new_n457_), .A1(new_new_n193_), .B0(new_new_n456_), .Y(new_new_n458_));
  NO3        g0436(.A(new_new_n458_), .B(new_new_n454_), .C(new_new_n450_), .Y(new_new_n459_));
  AOI210     g0437(.A0(new_new_n459_), .A1(new_new_n447_), .B0(new_new_n276_), .Y(new_new_n460_));
  NO4        g0438(.A(new_new_n460_), .B(new_new_n440_), .C(new_new_n419_), .D(new_new_n396_), .Y(new_new_n461_));
  NO2        g0439(.A(new_new_n64_), .B(i_4_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n74_), .B(i_13_), .Y(new_new_n463_));
  NO2        g0441(.A(i_10_), .B(i_9_), .Y(new_new_n464_));
  NAi21      g0442(.An(i_12_), .B(i_8_), .Y(new_new_n465_));
  NO2        g0443(.A(new_new_n465_), .B(i_3_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n314_), .B(i_0_), .Y(new_new_n467_));
  NO3        g0445(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n272_), .B(new_new_n99_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n469_), .B(new_new_n468_), .Y(new_new_n470_));
  NA2        g0448(.A(i_8_), .B(i_9_), .Y(new_new_n471_));
  AOI210     g0449(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n472_));
  OR2        g0450(.A(new_new_n472_), .B(new_new_n471_), .Y(new_new_n473_));
  NA2        g0451(.A(new_new_n287_), .B(new_new_n209_), .Y(new_new_n474_));
  NO2        g0452(.A(new_new_n474_), .B(new_new_n473_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n253_), .B(new_new_n313_), .Y(new_new_n476_));
  NO3        g0454(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n477_));
  AOI210     g0455(.A0(new_new_n259_), .A1(new_new_n192_), .B0(new_new_n477_), .Y(new_new_n478_));
  NA3        g0456(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n479_));
  NA4        g0457(.A(new_new_n147_), .B(new_new_n117_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n480_));
  OAI220     g0458(.A0(new_new_n480_), .A1(new_new_n479_), .B0(new_new_n478_), .B1(new_new_n476_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n481_), .B(new_new_n475_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n300_), .B(new_new_n110_), .Y(new_new_n483_));
  OR2        g0461(.A(new_new_n483_), .B(new_new_n211_), .Y(new_new_n484_));
  OA220      g0462(.A0(new_new_n302_), .A1(new_new_n164_), .B0(new_new_n484_), .B1(new_new_n233_), .Y(new_new_n485_));
  NA2        g0463(.A(new_new_n98_), .B(i_13_), .Y(new_new_n486_));
  NO2        g0464(.A(i_2_), .B(i_13_), .Y(new_new_n487_));
  NO3        g0465(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n488_));
  NO2        g0466(.A(i_6_), .B(i_7_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n490_));
  NO2        g0468(.A(i_11_), .B(i_1_), .Y(new_new_n491_));
  NO2        g0469(.A(new_new_n74_), .B(i_3_), .Y(new_new_n492_));
  OR2        g0470(.A(i_11_), .B(i_8_), .Y(new_new_n493_));
  NOi21      g0471(.An(i_2_), .B(i_7_), .Y(new_new_n494_));
  NAi31      g0472(.An(new_new_n493_), .B(new_new_n494_), .C(new_new_n492_), .Y(new_new_n495_));
  NO2        g0473(.A(new_new_n431_), .B(i_6_), .Y(new_new_n496_));
  NA3        g0474(.A(new_new_n496_), .B(new_new_n462_), .C(new_new_n76_), .Y(new_new_n497_));
  NO2        g0475(.A(new_new_n497_), .B(new_new_n495_), .Y(new_new_n498_));
  NO2        g0476(.A(i_3_), .B(new_new_n197_), .Y(new_new_n499_));
  NO2        g0477(.A(i_6_), .B(i_10_), .Y(new_new_n500_));
  NA4        g0478(.A(new_new_n500_), .B(new_new_n318_), .C(new_new_n499_), .D(new_new_n238_), .Y(new_new_n501_));
  NO2        g0479(.A(new_new_n501_), .B(new_new_n157_), .Y(new_new_n502_));
  NA3        g0480(.A(new_new_n247_), .B(new_new_n174_), .C(new_new_n134_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n504_));
  NO2        g0482(.A(new_new_n159_), .B(i_3_), .Y(new_new_n505_));
  NAi31      g0483(.An(new_new_n504_), .B(new_new_n505_), .C(new_new_n228_), .Y(new_new_n506_));
  NA3        g0484(.A(new_new_n409_), .B(new_new_n182_), .C(new_new_n151_), .Y(new_new_n507_));
  NA3        g0485(.A(new_new_n507_), .B(new_new_n506_), .C(new_new_n503_), .Y(new_new_n508_));
  NO3        g0486(.A(new_new_n508_), .B(new_new_n502_), .C(new_new_n498_), .Y(new_new_n509_));
  NA2        g0487(.A(new_new_n468_), .B(new_new_n398_), .Y(new_new_n510_));
  NA2        g0488(.A(new_new_n477_), .B(new_new_n404_), .Y(new_new_n511_));
  NO2        g0489(.A(new_new_n511_), .B(new_new_n226_), .Y(new_new_n512_));
  NAi21      g0490(.An(new_new_n220_), .B(new_new_n412_), .Y(new_new_n513_));
  NO2        g0491(.A(new_new_n26_), .B(i_5_), .Y(new_new_n514_));
  NO2        g0492(.A(i_0_), .B(new_new_n87_), .Y(new_new_n515_));
  NA3        g0493(.A(new_new_n515_), .B(new_new_n514_), .C(new_new_n144_), .Y(new_new_n516_));
  OR3        g0494(.A(new_new_n308_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n517_));
  NO2        g0495(.A(new_new_n517_), .B(new_new_n516_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n27_), .B(i_10_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n318_), .B(new_new_n240_), .Y(new_new_n520_));
  OAI220     g0498(.A0(new_new_n520_), .A1(new_new_n452_), .B0(new_new_n519_), .B1(new_new_n486_), .Y(new_new_n521_));
  NA4        g0499(.A(new_new_n311_), .B(new_new_n225_), .C(new_new_n74_), .D(new_new_n238_), .Y(new_new_n522_));
  NO2        g0500(.A(new_new_n522_), .B(new_new_n490_), .Y(new_new_n523_));
  NO4        g0501(.A(new_new_n523_), .B(new_new_n521_), .C(new_new_n518_), .D(new_new_n512_), .Y(new_new_n524_));
  NA4        g0502(.A(new_new_n524_), .B(new_new_n509_), .C(new_new_n485_), .D(new_new_n482_), .Y(new_new_n525_));
  NA3        g0503(.A(new_new_n311_), .B(new_new_n179_), .C(new_new_n177_), .Y(new_new_n526_));
  OAI210     g0504(.A0(new_new_n306_), .A1(new_new_n184_), .B0(new_new_n526_), .Y(new_new_n527_));
  AN2        g0505(.A(new_new_n291_), .B(new_new_n235_), .Y(new_new_n528_));
  NA2        g0506(.A(new_new_n528_), .B(new_new_n527_), .Y(new_new_n529_));
  NA2        g0507(.A(new_new_n318_), .B(new_new_n166_), .Y(new_new_n530_));
  OAI210     g0508(.A0(new_new_n530_), .A1(new_new_n233_), .B0(new_new_n312_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n531_), .B(new_new_n330_), .Y(new_new_n532_));
  NA4        g0510(.A(new_new_n463_), .B(new_new_n462_), .C(new_new_n207_), .D(i_2_), .Y(new_new_n533_));
  INV        g0511(.A(new_new_n533_), .Y(new_new_n534_));
  NA2        g0512(.A(new_new_n398_), .B(new_new_n227_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n368_), .B(new_new_n74_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n385_), .B(new_new_n377_), .Y(new_new_n537_));
  AO210      g0515(.A0(new_new_n536_), .A1(new_new_n535_), .B0(new_new_n537_), .Y(new_new_n538_));
  NO2        g0516(.A(new_new_n36_), .B(i_8_), .Y(new_new_n539_));
  NAi41      g0517(.An(new_new_n536_), .B(new_new_n500_), .C(new_new_n539_), .D(new_new_n47_), .Y(new_new_n540_));
  AOI210     g0518(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n432_), .Y(new_new_n541_));
  NA3        g0519(.A(new_new_n541_), .B(new_new_n540_), .C(new_new_n538_), .Y(new_new_n542_));
  AOI210     g0520(.A0(new_new_n534_), .A1(new_new_n208_), .B0(new_new_n542_), .Y(new_new_n543_));
  INV        g0521(.A(new_new_n136_), .Y(new_new_n544_));
  AOI210     g0522(.A0(new_new_n198_), .A1(i_9_), .B0(new_new_n271_), .Y(new_new_n545_));
  NO2        g0523(.A(new_new_n545_), .B(new_new_n203_), .Y(new_new_n546_));
  OR2        g0524(.A(new_new_n186_), .B(i_4_), .Y(new_new_n547_));
  NO2        g0525(.A(new_new_n547_), .B(new_new_n87_), .Y(new_new_n548_));
  AOI220     g0526(.A0(new_new_n548_), .A1(new_new_n546_), .B0(new_new_n544_), .B1(new_new_n433_), .Y(new_new_n549_));
  NA4        g0527(.A(new_new_n549_), .B(new_new_n543_), .C(new_new_n532_), .D(new_new_n529_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n403_), .B(new_new_n300_), .Y(new_new_n551_));
  OAI210     g0529(.A0(new_new_n399_), .A1(new_new_n171_), .B0(new_new_n551_), .Y(new_new_n552_));
  NO2        g0530(.A(i_12_), .B(new_new_n197_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n553_), .B(new_new_n227_), .Y(new_new_n554_));
  NA3        g0532(.A(new_new_n500_), .B(new_new_n177_), .C(new_new_n27_), .Y(new_new_n555_));
  NO2        g0533(.A(new_new_n555_), .B(new_new_n554_), .Y(new_new_n556_));
  NOi31      g0534(.An(new_new_n321_), .B(new_new_n431_), .C(new_new_n38_), .Y(new_new_n557_));
  OAI210     g0535(.A0(new_new_n557_), .A1(new_new_n556_), .B0(new_new_n552_), .Y(new_new_n558_));
  NO2        g0536(.A(i_8_), .B(i_7_), .Y(new_new_n559_));
  OAI210     g0537(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n560_));
  NA2        g0538(.A(new_new_n560_), .B(new_new_n225_), .Y(new_new_n561_));
  AOI220     g0539(.A0(new_new_n331_), .A1(new_new_n40_), .B0(new_new_n236_), .B1(new_new_n210_), .Y(new_new_n562_));
  OAI220     g0540(.A0(new_new_n562_), .A1(new_new_n547_), .B0(new_new_n561_), .B1(new_new_n244_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n45_), .B(i_10_), .Y(new_new_n564_));
  NO2        g0542(.A(new_new_n564_), .B(i_6_), .Y(new_new_n565_));
  NA3        g0543(.A(new_new_n565_), .B(new_new_n563_), .C(new_new_n559_), .Y(new_new_n566_));
  NOi31      g0544(.An(new_new_n295_), .B(new_new_n306_), .C(new_new_n184_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n159_), .B(i_5_), .Y(new_new_n568_));
  NA2        g0546(.A(new_new_n567_), .B(new_new_n477_), .Y(new_new_n569_));
  NA3        g0547(.A(new_new_n569_), .B(new_new_n566_), .C(new_new_n558_), .Y(new_new_n570_));
  NA3        g0548(.A(new_new_n221_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n571_));
  NA2        g0549(.A(new_new_n287_), .B(new_new_n85_), .Y(new_new_n572_));
  AOI210     g0550(.A0(new_new_n571_), .A1(new_new_n358_), .B0(new_new_n572_), .Y(new_new_n573_));
  NA2        g0551(.A(new_new_n301_), .B(new_new_n291_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n574_), .B(new_new_n176_), .Y(new_new_n575_));
  NA2        g0553(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n464_), .B(new_new_n223_), .Y(new_new_n577_));
  NO2        g0555(.A(new_new_n576_), .B(new_new_n577_), .Y(new_new_n578_));
  AOI210     g0556(.A0(new_new_n378_), .A1(new_new_n47_), .B0(new_new_n382_), .Y(new_new_n579_));
  NA2        g0557(.A(i_0_), .B(new_new_n49_), .Y(new_new_n580_));
  NA3        g0558(.A(new_new_n553_), .B(new_new_n278_), .C(new_new_n580_), .Y(new_new_n581_));
  NO2        g0559(.A(new_new_n579_), .B(new_new_n581_), .Y(new_new_n582_));
  NO4        g0560(.A(new_new_n582_), .B(new_new_n578_), .C(new_new_n575_), .D(new_new_n573_), .Y(new_new_n583_));
  NO4        g0561(.A(new_new_n254_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n584_));
  NO3        g0562(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n234_), .B(new_new_n36_), .Y(new_new_n586_));
  AN2        g0564(.A(new_new_n586_), .B(new_new_n585_), .Y(new_new_n587_));
  OA210      g0565(.A0(new_new_n587_), .A1(new_new_n584_), .B0(new_new_n368_), .Y(new_new_n588_));
  NO2        g0566(.A(new_new_n431_), .B(i_1_), .Y(new_new_n589_));
  NOi31      g0567(.An(new_new_n589_), .B(new_new_n469_), .C(new_new_n74_), .Y(new_new_n590_));
  AN4        g0568(.A(new_new_n590_), .B(new_new_n428_), .C(new_new_n514_), .D(i_2_), .Y(new_new_n591_));
  NO2        g0569(.A(new_new_n442_), .B(new_new_n180_), .Y(new_new_n592_));
  NO3        g0570(.A(new_new_n592_), .B(new_new_n591_), .C(new_new_n588_), .Y(new_new_n593_));
  NOi21      g0571(.An(i_10_), .B(i_6_), .Y(new_new_n594_));
  NO2        g0572(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n596_));
  NA2        g0574(.A(new_new_n321_), .B(new_new_n166_), .Y(new_new_n597_));
  AOI220     g0575(.A0(new_new_n597_), .A1(new_new_n453_), .B0(new_new_n187_), .B1(new_new_n185_), .Y(new_new_n598_));
  NOi31      g0576(.An(new_new_n148_), .B(i_10_), .C(new_new_n339_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n599_), .B(new_new_n598_), .Y(new_new_n600_));
  NO2        g0578(.A(i_12_), .B(new_new_n87_), .Y(new_new_n601_));
  NA2        g0579(.A(new_new_n177_), .B(i_0_), .Y(new_new_n602_));
  NO3        g0580(.A(new_new_n602_), .B(new_new_n350_), .C(new_new_n306_), .Y(new_new_n603_));
  OR2        g0581(.A(i_2_), .B(i_5_), .Y(new_new_n604_));
  OR2        g0582(.A(new_new_n604_), .B(new_new_n423_), .Y(new_new_n605_));
  AOI210     g0583(.A0(new_new_n387_), .A1(new_new_n246_), .B0(new_new_n202_), .Y(new_new_n606_));
  AOI210     g0584(.A0(new_new_n606_), .A1(new_new_n605_), .B0(new_new_n513_), .Y(new_new_n607_));
  NO2        g0585(.A(new_new_n607_), .B(new_new_n603_), .Y(new_new_n608_));
  NA4        g0586(.A(new_new_n608_), .B(new_new_n600_), .C(new_new_n593_), .D(new_new_n583_), .Y(new_new_n609_));
  NO4        g0587(.A(new_new_n609_), .B(new_new_n570_), .C(new_new_n550_), .D(new_new_n525_), .Y(new_new_n610_));
  NA4        g0588(.A(new_new_n610_), .B(new_new_n461_), .C(new_new_n367_), .D(new_new_n317_), .Y(zz07));
  NO2        g0589(.A(new_new_n94_), .B(new_new_n55_), .Y(new_new_n612_));
  NA2        g0590(.A(new_new_n500_), .B(new_new_n85_), .Y(new_new_n613_));
  NA2        g0591(.A(i_11_), .B(new_new_n197_), .Y(new_new_n614_));
  NA2        g0592(.A(new_new_n146_), .B(new_new_n614_), .Y(new_new_n615_));
  NO2        g0593(.A(new_new_n615_), .B(new_new_n613_), .Y(new_new_n616_));
  NA3        g0594(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n617_));
  NO2        g0595(.A(new_new_n238_), .B(i_4_), .Y(new_new_n618_));
  NA2        g0596(.A(new_new_n618_), .B(i_8_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n107_), .B(new_new_n617_), .Y(new_new_n620_));
  NA2        g0598(.A(i_2_), .B(new_new_n87_), .Y(new_new_n621_));
  OAI210     g0599(.A0(new_new_n88_), .A1(new_new_n207_), .B0(new_new_n208_), .Y(new_new_n622_));
  NO2        g0600(.A(i_7_), .B(new_new_n37_), .Y(new_new_n623_));
  NA2        g0601(.A(i_4_), .B(i_8_), .Y(new_new_n624_));
  AOI210     g0602(.A0(new_new_n624_), .A1(new_new_n311_), .B0(new_new_n623_), .Y(new_new_n625_));
  OAI220     g0603(.A0(new_new_n625_), .A1(new_new_n621_), .B0(new_new_n622_), .B1(i_13_), .Y(new_new_n626_));
  NO4        g0604(.A(new_new_n626_), .B(new_new_n620_), .C(new_new_n616_), .D(new_new_n612_), .Y(new_new_n627_));
  AOI210     g0605(.A0(new_new_n130_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n628_));
  AOI210     g0606(.A0(new_new_n628_), .A1(new_new_n238_), .B0(new_new_n163_), .Y(new_new_n629_));
  OR2        g0607(.A(i_6_), .B(i_10_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n630_), .B(new_new_n23_), .Y(new_new_n631_));
  OR3        g0609(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n632_));
  NO3        g0610(.A(new_new_n632_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n633_));
  INV        g0611(.A(new_new_n204_), .Y(new_new_n634_));
  OR2        g0612(.A(new_new_n629_), .B(new_new_n273_), .Y(new_new_n635_));
  AOI210     g0613(.A0(new_new_n635_), .A1(new_new_n627_), .B0(new_new_n64_), .Y(new_new_n636_));
  NOi21      g0614(.An(i_11_), .B(i_7_), .Y(new_new_n637_));
  AO210      g0615(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n638_));
  NO2        g0616(.A(new_new_n638_), .B(new_new_n637_), .Y(new_new_n639_));
  NA2        g0617(.A(new_new_n639_), .B(new_new_n210_), .Y(new_new_n640_));
  NA3        g0618(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n641_));
  NO2        g0619(.A(new_new_n640_), .B(new_new_n64_), .Y(new_new_n642_));
  OR2        g0620(.A(new_new_n393_), .B(new_new_n41_), .Y(new_new_n643_));
  NO3        g0621(.A(new_new_n262_), .B(new_new_n212_), .C(new_new_n614_), .Y(new_new_n644_));
  OAI210     g0622(.A0(new_new_n644_), .A1(new_new_n228_), .B0(new_new_n64_), .Y(new_new_n645_));
  NA2        g0623(.A(new_new_n424_), .B(new_new_n31_), .Y(new_new_n646_));
  OR2        g0624(.A(new_new_n212_), .B(new_new_n110_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n647_), .B(new_new_n646_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n64_), .B(i_9_), .Y(new_new_n649_));
  NO2        g0627(.A(new_new_n649_), .B(i_4_), .Y(new_new_n650_));
  NA2        g0628(.A(new_new_n650_), .B(new_new_n648_), .Y(new_new_n651_));
  NO2        g0629(.A(i_1_), .B(i_12_), .Y(new_new_n652_));
  NA3        g0630(.A(new_new_n651_), .B(new_new_n645_), .C(new_new_n643_), .Y(new_new_n653_));
  OAI210     g0631(.A0(new_new_n653_), .A1(new_new_n642_), .B0(i_6_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n641_), .B(new_new_n110_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n655_), .B(new_new_n601_), .Y(new_new_n656_));
  NO2        g0634(.A(i_6_), .B(i_11_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n656_), .B(new_new_n470_), .Y(new_new_n658_));
  NO4        g0636(.A(new_new_n219_), .B(new_new_n130_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n659_));
  NA2        g0637(.A(new_new_n659_), .B(new_new_n649_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n238_), .B(i_6_), .Y(new_new_n661_));
  NO3        g0639(.A(new_new_n630_), .B(new_new_n234_), .C(new_new_n23_), .Y(new_new_n662_));
  AOI210     g0640(.A0(i_1_), .A1(new_new_n263_), .B0(new_new_n662_), .Y(new_new_n663_));
  OAI210     g0641(.A0(new_new_n663_), .A1(new_new_n45_), .B0(new_new_n660_), .Y(new_new_n664_));
  NA3        g0642(.A(new_new_n559_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n140_), .B(i_9_), .Y(new_new_n666_));
  NA3        g0644(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n47_), .B(i_1_), .Y(new_new_n668_));
  NA3        g0646(.A(new_new_n668_), .B(new_new_n272_), .C(new_new_n45_), .Y(new_new_n669_));
  OAI220     g0647(.A0(new_new_n669_), .A1(new_new_n667_), .B0(new_new_n666_), .B1(new_new_n1073_), .Y(new_new_n670_));
  NA3        g0648(.A(new_new_n649_), .B(new_new_n324_), .C(i_6_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n671_), .B(new_new_n23_), .Y(new_new_n672_));
  AOI210     g0650(.A0(new_new_n491_), .A1(new_new_n435_), .B0(new_new_n243_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n673_), .B(new_new_n621_), .Y(new_new_n674_));
  NAi21      g0652(.An(new_new_n665_), .B(new_new_n93_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n668_), .B(new_new_n272_), .Y(new_new_n676_));
  NO2        g0654(.A(i_11_), .B(new_new_n37_), .Y(new_new_n677_));
  NA2        g0655(.A(new_new_n677_), .B(new_new_n24_), .Y(new_new_n678_));
  OAI210     g0656(.A0(new_new_n678_), .A1(new_new_n676_), .B0(new_new_n675_), .Y(new_new_n679_));
  OR4        g0657(.A(new_new_n679_), .B(new_new_n674_), .C(new_new_n672_), .D(new_new_n670_), .Y(new_new_n680_));
  NO3        g0658(.A(new_new_n680_), .B(new_new_n664_), .C(new_new_n658_), .Y(new_new_n681_));
  NO2        g0659(.A(new_new_n238_), .B(new_new_n103_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n682_), .B(new_new_n637_), .Y(new_new_n683_));
  NA2        g0661(.A(new_new_n683_), .B(i_1_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n684_), .B(new_new_n632_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n430_), .B(new_new_n87_), .Y(new_new_n686_));
  NA2        g0664(.A(new_new_n685_), .B(new_new_n47_), .Y(new_new_n687_));
  NA2        g0665(.A(i_3_), .B(new_new_n197_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n688_), .B(new_new_n116_), .Y(new_new_n689_));
  AN2        g0667(.A(new_new_n689_), .B(new_new_n565_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n234_), .B(new_new_n45_), .Y(new_new_n691_));
  NO3        g0669(.A(new_new_n691_), .B(new_new_n314_), .C(new_new_n239_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n119_), .B(new_new_n37_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n693_), .B(i_6_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n87_), .B(i_9_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n695_), .B(new_new_n64_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n696_), .B(new_new_n652_), .Y(new_new_n697_));
  NO4        g0675(.A(new_new_n697_), .B(new_new_n694_), .C(new_new_n692_), .D(i_4_), .Y(new_new_n698_));
  NA2        g0676(.A(i_1_), .B(i_3_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n471_), .B(new_new_n94_), .Y(new_new_n700_));
  AOI210     g0678(.A0(new_new_n691_), .A1(new_new_n594_), .B0(new_new_n700_), .Y(new_new_n701_));
  NO2        g0679(.A(new_new_n701_), .B(new_new_n699_), .Y(new_new_n702_));
  NO3        g0680(.A(new_new_n702_), .B(new_new_n698_), .C(new_new_n690_), .Y(new_new_n703_));
  NA4        g0681(.A(new_new_n703_), .B(new_new_n687_), .C(new_new_n681_), .D(new_new_n654_), .Y(new_new_n704_));
  NO3        g0682(.A(new_new_n493_), .B(i_3_), .C(i_7_), .Y(new_new_n705_));
  NOi21      g0683(.An(new_new_n705_), .B(i_10_), .Y(new_new_n706_));
  OA210      g0684(.A0(new_new_n706_), .A1(new_new_n247_), .B0(new_new_n87_), .Y(new_new_n707_));
  NA2        g0685(.A(new_new_n385_), .B(new_new_n384_), .Y(new_new_n708_));
  NA3        g0686(.A(new_new_n500_), .B(new_new_n539_), .C(new_new_n47_), .Y(new_new_n709_));
  NO3        g0687(.A(new_new_n494_), .B(new_new_n624_), .C(new_new_n87_), .Y(new_new_n710_));
  NA2        g0688(.A(new_new_n710_), .B(new_new_n25_), .Y(new_new_n711_));
  NA3        g0689(.A(new_new_n711_), .B(new_new_n709_), .C(new_new_n708_), .Y(new_new_n712_));
  OAI210     g0690(.A0(new_new_n712_), .A1(new_new_n707_), .B0(i_1_), .Y(new_new_n713_));
  AOI210     g0691(.A0(new_new_n272_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n714_));
  NO2        g0692(.A(new_new_n383_), .B(i_2_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n715_), .B(new_new_n714_), .Y(new_new_n716_));
  OAI210     g0694(.A0(new_new_n671_), .A1(new_new_n465_), .B0(new_new_n716_), .Y(new_new_n717_));
  INV        g0695(.A(new_new_n717_), .Y(new_new_n718_));
  AOI210     g0696(.A0(new_new_n718_), .A1(new_new_n713_), .B0(i_13_), .Y(new_new_n719_));
  OR2        g0697(.A(i_11_), .B(i_7_), .Y(new_new_n720_));
  AOI210     g0698(.A0(new_new_n667_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n721_));
  NO2        g0699(.A(new_new_n494_), .B(new_new_n24_), .Y(new_new_n722_));
  AOI220     g0700(.A0(new_new_n722_), .A1(new_new_n686_), .B0(new_new_n247_), .B1(new_new_n133_), .Y(new_new_n723_));
  OAI220     g0701(.A0(new_new_n723_), .A1(new_new_n41_), .B0(new_new_n1072_), .B1(new_new_n94_), .Y(new_new_n724_));
  INV        g0702(.A(new_new_n724_), .Y(new_new_n725_));
  INV        g0703(.A(new_new_n116_), .Y(new_new_n726_));
  AOI220     g0704(.A0(new_new_n726_), .A1(new_new_n73_), .B0(new_new_n400_), .B1(new_new_n668_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n727_), .B(new_new_n244_), .Y(new_new_n728_));
  AOI210     g0706(.A0(new_new_n465_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n729_));
  NOi31      g0707(.An(new_new_n729_), .B(new_new_n613_), .C(new_new_n45_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n129_), .B(i_13_), .Y(new_new_n731_));
  NO2        g0709(.A(new_new_n667_), .B(new_new_n116_), .Y(new_new_n732_));
  INV        g0710(.A(new_new_n732_), .Y(new_new_n733_));
  OAI220     g0711(.A0(new_new_n733_), .A1(new_new_n72_), .B0(new_new_n731_), .B1(new_new_n714_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n26_), .B(new_new_n197_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n735_), .B(i_7_), .Y(new_new_n736_));
  NO3        g0714(.A(new_new_n494_), .B(new_new_n238_), .C(new_new_n87_), .Y(new_new_n737_));
  NA2        g0715(.A(new_new_n737_), .B(new_new_n736_), .Y(new_new_n738_));
  AOI220     g0716(.A0(new_new_n400_), .A1(new_new_n668_), .B0(new_new_n93_), .B1(new_new_n104_), .Y(new_new_n739_));
  OAI220     g0717(.A0(new_new_n739_), .A1(new_new_n619_), .B0(new_new_n738_), .B1(new_new_n634_), .Y(new_new_n740_));
  NO4        g0718(.A(new_new_n740_), .B(new_new_n734_), .C(new_new_n730_), .D(new_new_n728_), .Y(new_new_n741_));
  OR2        g0719(.A(i_11_), .B(i_6_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n618_), .B(new_new_n735_), .C(i_7_), .Y(new_new_n743_));
  AOI210     g0721(.A0(new_new_n743_), .A1(new_new_n733_), .B0(new_new_n742_), .Y(new_new_n744_));
  NA3        g0722(.A(new_new_n424_), .B(new_new_n623_), .C(new_new_n99_), .Y(new_new_n745_));
  NA2        g0723(.A(new_new_n657_), .B(i_13_), .Y(new_new_n746_));
  NA2        g0724(.A(new_new_n104_), .B(new_new_n735_), .Y(new_new_n747_));
  NAi21      g0725(.An(i_11_), .B(i_12_), .Y(new_new_n748_));
  NOi41      g0726(.An(new_new_n112_), .B(new_new_n748_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n749_));
  NO3        g0727(.A(new_new_n494_), .B(new_new_n601_), .C(new_new_n624_), .Y(new_new_n750_));
  AOI220     g0728(.A0(new_new_n750_), .A1(new_new_n318_), .B0(new_new_n749_), .B1(new_new_n747_), .Y(new_new_n751_));
  NA3        g0729(.A(new_new_n751_), .B(new_new_n746_), .C(new_new_n745_), .Y(new_new_n752_));
  OAI210     g0730(.A0(new_new_n752_), .A1(new_new_n744_), .B0(new_new_n64_), .Y(new_new_n753_));
  NO2        g0731(.A(i_2_), .B(i_12_), .Y(new_new_n754_));
  NA2        g0732(.A(new_new_n382_), .B(new_new_n754_), .Y(new_new_n755_));
  NA2        g0733(.A(new_new_n384_), .B(new_new_n382_), .Y(new_new_n756_));
  NO2        g0734(.A(new_new_n130_), .B(i_2_), .Y(new_new_n757_));
  NA2        g0735(.A(new_new_n757_), .B(new_new_n652_), .Y(new_new_n758_));
  NA3        g0736(.A(new_new_n758_), .B(new_new_n756_), .C(new_new_n755_), .Y(new_new_n759_));
  NA3        g0737(.A(new_new_n759_), .B(new_new_n46_), .C(new_new_n227_), .Y(new_new_n760_));
  NA4        g0738(.A(new_new_n760_), .B(new_new_n753_), .C(new_new_n741_), .D(new_new_n725_), .Y(new_new_n761_));
  OR4        g0739(.A(new_new_n761_), .B(new_new_n719_), .C(new_new_n704_), .D(new_new_n636_), .Y(zz05));
  NA2        g0740(.A(new_new_n683_), .B(new_new_n275_), .Y(new_new_n763_));
  AN2        g0741(.A(new_new_n24_), .B(i_10_), .Y(new_new_n764_));
  NA3        g0742(.A(new_new_n764_), .B(new_new_n754_), .C(new_new_n110_), .Y(new_new_n765_));
  NO2        g0743(.A(new_new_n619_), .B(i_11_), .Y(new_new_n766_));
  OAI210     g0744(.A0(new_new_n623_), .A1(new_new_n88_), .B0(new_new_n766_), .Y(new_new_n767_));
  NA3        g0745(.A(new_new_n767_), .B(new_new_n765_), .C(new_new_n763_), .Y(new_new_n768_));
  NO3        g0746(.A(i_11_), .B(new_new_n238_), .C(i_13_), .Y(new_new_n769_));
  NO2        g0747(.A(new_new_n126_), .B(new_new_n23_), .Y(new_new_n770_));
  NA2        g0748(.A(i_12_), .B(i_8_), .Y(new_new_n771_));
  OAI210     g0749(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n771_), .Y(new_new_n772_));
  INV        g0750(.A(new_new_n464_), .Y(new_new_n773_));
  AOI220     g0751(.A0(new_new_n324_), .A1(new_new_n596_), .B0(new_new_n772_), .B1(new_new_n770_), .Y(new_new_n774_));
  INV        g0752(.A(new_new_n774_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n775_), .B(new_new_n768_), .Y(new_new_n776_));
  INV        g0754(.A(new_new_n174_), .Y(new_new_n777_));
  INV        g0755(.A(new_new_n247_), .Y(new_new_n778_));
  OAI210     g0756(.A0(new_new_n715_), .A1(new_new_n466_), .B0(new_new_n112_), .Y(new_new_n779_));
  AOI210     g0757(.A0(new_new_n779_), .A1(new_new_n778_), .B0(new_new_n777_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n471_), .B(new_new_n26_), .Y(new_new_n781_));
  NO2        g0759(.A(new_new_n781_), .B(new_new_n435_), .Y(new_new_n782_));
  NA2        g0760(.A(new_new_n782_), .B(i_2_), .Y(new_new_n783_));
  INV        g0761(.A(new_new_n783_), .Y(new_new_n784_));
  AOI210     g0762(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n431_), .Y(new_new_n785_));
  AOI210     g0763(.A0(new_new_n785_), .A1(new_new_n784_), .B0(new_new_n780_), .Y(new_new_n786_));
  NO2        g0764(.A(new_new_n194_), .B(new_new_n127_), .Y(new_new_n787_));
  OAI210     g0765(.A0(new_new_n787_), .A1(new_new_n770_), .B0(i_2_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n175_), .Y(new_new_n789_));
  NO3        g0767(.A(new_new_n638_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n790_));
  AOI210     g0768(.A0(new_new_n789_), .A1(new_new_n88_), .B0(new_new_n790_), .Y(new_new_n791_));
  AOI210     g0769(.A0(new_new_n791_), .A1(new_new_n788_), .B0(new_new_n197_), .Y(new_new_n792_));
  OA210      g0770(.A0(new_new_n639_), .A1(new_new_n128_), .B0(i_13_), .Y(new_new_n793_));
  NA2        g0771(.A(new_new_n204_), .B(new_new_n207_), .Y(new_new_n794_));
  NA2        g0772(.A(new_new_n153_), .B(new_new_n614_), .Y(new_new_n795_));
  AOI210     g0773(.A0(new_new_n795_), .A1(new_new_n794_), .B0(new_new_n387_), .Y(new_new_n796_));
  AOI210     g0774(.A0(new_new_n212_), .A1(new_new_n150_), .B0(new_new_n539_), .Y(new_new_n797_));
  OAI210     g0775(.A0(new_new_n797_), .A1(new_new_n228_), .B0(new_new_n435_), .Y(new_new_n798_));
  NO2        g0776(.A(new_new_n104_), .B(new_new_n45_), .Y(new_new_n799_));
  INV        g0777(.A(new_new_n307_), .Y(new_new_n800_));
  NA4        g0778(.A(new_new_n800_), .B(new_new_n311_), .C(new_new_n126_), .D(new_new_n43_), .Y(new_new_n801_));
  OAI210     g0779(.A0(new_new_n801_), .A1(new_new_n799_), .B0(new_new_n798_), .Y(new_new_n802_));
  NO4        g0780(.A(new_new_n802_), .B(new_new_n796_), .C(new_new_n793_), .D(new_new_n792_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n596_), .B(new_new_n28_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n769_), .B(new_new_n279_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n805_), .B(new_new_n804_), .Y(new_new_n806_));
  NO2        g0784(.A(new_new_n63_), .B(i_12_), .Y(new_new_n807_));
  NO2        g0785(.A(new_new_n807_), .B(new_new_n128_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n808_), .B(new_new_n614_), .Y(new_new_n809_));
  AOI220     g0787(.A0(new_new_n809_), .A1(new_new_n36_), .B0(new_new_n806_), .B1(new_new_n47_), .Y(new_new_n810_));
  NA4        g0788(.A(new_new_n810_), .B(new_new_n803_), .C(new_new_n786_), .D(new_new_n776_), .Y(zz06));
  NO3        g0789(.A(new_new_n258_), .B(new_new_n313_), .C(i_1_), .Y(new_new_n812_));
  NO2        g0790(.A(new_new_n189_), .B(new_new_n141_), .Y(new_new_n813_));
  OAI210     g0791(.A0(new_new_n813_), .A1(new_new_n812_), .B0(new_new_n757_), .Y(new_new_n814_));
  NA4        g0792(.A(new_new_n404_), .B(new_new_n499_), .C(new_new_n72_), .D(new_new_n103_), .Y(new_new_n815_));
  INV        g0793(.A(new_new_n815_), .Y(new_new_n816_));
  NO2        g0794(.A(new_new_n222_), .B(new_new_n504_), .Y(new_new_n817_));
  NO2        g0795(.A(i_11_), .B(i_9_), .Y(new_new_n818_));
  NO2        g0796(.A(new_new_n816_), .B(new_new_n336_), .Y(new_new_n819_));
  AO210      g0797(.A0(new_new_n819_), .A1(new_new_n814_), .B0(i_12_), .Y(new_new_n820_));
  NA2        g0798(.A(new_new_n388_), .B(new_new_n344_), .Y(new_new_n821_));
  NA2        g0799(.A(new_new_n601_), .B(new_new_n64_), .Y(new_new_n822_));
  NA2        g0800(.A(new_new_n706_), .B(new_new_n72_), .Y(new_new_n823_));
  NA3        g0801(.A(new_new_n823_), .B(new_new_n822_), .C(new_new_n821_), .Y(new_new_n824_));
  INV        g0802(.A(new_new_n201_), .Y(new_new_n825_));
  AOI220     g0803(.A0(new_new_n825_), .A1(new_new_n818_), .B0(new_new_n824_), .B1(new_new_n74_), .Y(new_new_n826_));
  INV        g0804(.A(new_new_n335_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n76_), .B(new_new_n133_), .Y(new_new_n828_));
  INV        g0806(.A(new_new_n126_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n829_), .B(new_new_n47_), .Y(new_new_n830_));
  AOI210     g0808(.A0(new_new_n830_), .A1(new_new_n828_), .B0(new_new_n827_), .Y(new_new_n831_));
  NO3        g0809(.A(new_new_n254_), .B(new_new_n134_), .C(i_9_), .Y(new_new_n832_));
  NA2        g0810(.A(new_new_n832_), .B(new_new_n807_), .Y(new_new_n833_));
  AOI210     g0811(.A0(new_new_n833_), .A1(new_new_n537_), .B0(new_new_n189_), .Y(new_new_n834_));
  NO2        g0812(.A(new_new_n32_), .B(i_11_), .Y(new_new_n835_));
  NA3        g0813(.A(new_new_n835_), .B(new_new_n489_), .C(new_new_n404_), .Y(new_new_n836_));
  NAi32      g0814(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n837_));
  NO2        g0815(.A(new_new_n742_), .B(new_new_n837_), .Y(new_new_n838_));
  OAI210     g0816(.A0(new_new_n705_), .A1(new_new_n586_), .B0(new_new_n585_), .Y(new_new_n839_));
  NAi31      g0817(.An(new_new_n838_), .B(new_new_n839_), .C(new_new_n836_), .Y(new_new_n840_));
  OR3        g0818(.A(new_new_n840_), .B(new_new_n834_), .C(new_new_n831_), .Y(new_new_n841_));
  NO2        g0819(.A(new_new_n720_), .B(i_2_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n843_));
  NO2        g0821(.A(new_new_n843_), .B(new_new_n423_), .Y(new_new_n844_));
  NA2        g0822(.A(new_new_n844_), .B(new_new_n842_), .Y(new_new_n845_));
  AO220      g0823(.A0(new_new_n372_), .A1(new_new_n362_), .B0(new_new_n410_), .B1(new_new_n614_), .Y(new_new_n846_));
  NA3        g0824(.A(new_new_n846_), .B(new_new_n259_), .C(i_7_), .Y(new_new_n847_));
  NA3        g0825(.A(new_new_n639_), .B(new_new_n149_), .C(new_new_n70_), .Y(new_new_n848_));
  AO210      g0826(.A0(new_new_n511_), .A1(new_new_n773_), .B0(new_new_n36_), .Y(new_new_n849_));
  NA4        g0827(.A(new_new_n849_), .B(new_new_n848_), .C(new_new_n847_), .D(new_new_n845_), .Y(new_new_n850_));
  NO2        g0828(.A(i_6_), .B(i_11_), .Y(new_new_n851_));
  AOI220     g0829(.A0(new_new_n851_), .A1(new_new_n585_), .B0(new_new_n817_), .B1(new_new_n736_), .Y(new_new_n852_));
  NA3        g0830(.A(new_new_n387_), .B(new_new_n240_), .C(new_new_n149_), .Y(new_new_n853_));
  NA2        g0831(.A(new_new_n410_), .B(new_new_n71_), .Y(new_new_n854_));
  NA4        g0832(.A(new_new_n854_), .B(new_new_n853_), .C(new_new_n852_), .D(new_new_n622_), .Y(new_new_n855_));
  AN2        g0833(.A(new_new_n539_), .B(new_new_n47_), .Y(new_new_n856_));
  NA3        g0834(.A(new_new_n856_), .B(new_new_n500_), .C(new_new_n221_), .Y(new_new_n857_));
  AOI210     g0835(.A0(new_new_n466_), .A1(new_new_n464_), .B0(new_new_n584_), .Y(new_new_n858_));
  NO2        g0836(.A(new_new_n630_), .B(new_new_n104_), .Y(new_new_n859_));
  OAI210     g0837(.A0(new_new_n859_), .A1(new_new_n113_), .B0(new_new_n421_), .Y(new_new_n860_));
  INV        g0838(.A(new_new_n605_), .Y(new_new_n861_));
  NA3        g0839(.A(new_new_n861_), .B(new_new_n335_), .C(i_7_), .Y(new_new_n862_));
  NA4        g0840(.A(new_new_n862_), .B(new_new_n860_), .C(new_new_n858_), .D(new_new_n857_), .Y(new_new_n863_));
  NO4        g0841(.A(new_new_n863_), .B(new_new_n855_), .C(new_new_n850_), .D(new_new_n841_), .Y(new_new_n864_));
  NA4        g0842(.A(new_new_n864_), .B(new_new_n826_), .C(new_new_n820_), .D(new_new_n395_), .Y(zz03));
  NA2        g0843(.A(i_12_), .B(i_10_), .Y(new_new_n866_));
  NA2        g0844(.A(i_6_), .B(i_7_), .Y(new_new_n867_));
  NO2        g0845(.A(new_new_n867_), .B(i_0_), .Y(new_new_n868_));
  NO2        g0846(.A(i_11_), .B(new_new_n238_), .Y(new_new_n869_));
  OAI210     g0847(.A0(new_new_n868_), .A1(new_new_n295_), .B0(new_new_n869_), .Y(new_new_n870_));
  NO2        g0848(.A(new_new_n870_), .B(new_new_n197_), .Y(new_new_n871_));
  NO3        g0849(.A(new_new_n467_), .B(new_new_n91_), .C(new_new_n45_), .Y(new_new_n872_));
  OA210      g0850(.A0(new_new_n872_), .A1(new_new_n871_), .B0(new_new_n177_), .Y(new_new_n873_));
  NA2        g0851(.A(new_new_n853_), .B(new_new_n386_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n874_), .B(new_new_n40_), .Y(new_new_n875_));
  NOi21      g0853(.An(new_new_n98_), .B(new_new_n782_), .Y(new_new_n876_));
  NO3        g0854(.A(new_new_n647_), .B(new_new_n471_), .C(new_new_n133_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n424_), .B(new_new_n46_), .Y(new_new_n878_));
  AN2        g0856(.A(new_new_n469_), .B(new_new_n56_), .Y(new_new_n879_));
  NO3        g0857(.A(new_new_n879_), .B(new_new_n877_), .C(new_new_n876_), .Y(new_new_n880_));
  AOI210     g0858(.A0(new_new_n880_), .A1(new_new_n875_), .B0(new_new_n49_), .Y(new_new_n881_));
  NO4        g0859(.A(new_new_n391_), .B(new_new_n398_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n882_));
  NA2        g0860(.A(new_new_n189_), .B(new_new_n594_), .Y(new_new_n883_));
  NOi31      g0861(.An(new_new_n883_), .B(new_new_n882_), .C(new_new_n39_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n729_), .B(new_new_n695_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n342_), .B(new_new_n455_), .Y(new_new_n886_));
  OAI220     g0864(.A0(new_new_n886_), .A1(new_new_n885_), .B0(new_new_n884_), .B1(new_new_n64_), .Y(new_new_n887_));
  NOi21      g0865(.An(i_5_), .B(i_9_), .Y(new_new_n888_));
  NA2        g0866(.A(new_new_n888_), .B(new_new_n463_), .Y(new_new_n889_));
  BUFFER     g0867(.A(new_new_n272_), .Y(new_new_n890_));
  AOI210     g0868(.A0(new_new_n890_), .A1(new_new_n491_), .B0(new_new_n710_), .Y(new_new_n891_));
  NO3        g0869(.A(new_new_n427_), .B(new_new_n272_), .C(new_new_n74_), .Y(new_new_n892_));
  NO2        g0870(.A(new_new_n178_), .B(new_new_n150_), .Y(new_new_n893_));
  AOI210     g0871(.A0(new_new_n893_), .A1(new_new_n246_), .B0(new_new_n892_), .Y(new_new_n894_));
  OAI220     g0872(.A0(new_new_n894_), .A1(new_new_n184_), .B0(new_new_n891_), .B1(new_new_n889_), .Y(new_new_n895_));
  NO4        g0873(.A(new_new_n895_), .B(new_new_n887_), .C(new_new_n881_), .D(new_new_n873_), .Y(new_new_n896_));
  NA2        g0874(.A(new_new_n189_), .B(new_new_n24_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n318_), .B(new_new_n131_), .Y(new_new_n898_));
  NO2        g0876(.A(new_new_n898_), .B(new_new_n413_), .Y(new_new_n899_));
  INV        g0877(.A(new_new_n899_), .Y(new_new_n900_));
  NO2        g0878(.A(new_new_n404_), .B(new_new_n299_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n901_), .B(new_new_n732_), .Y(new_new_n902_));
  NA2        g0880(.A(new_new_n595_), .B(i_0_), .Y(new_new_n903_));
  NO4        g0881(.A(new_new_n604_), .B(new_new_n219_), .C(new_new_n431_), .D(new_new_n423_), .Y(new_new_n904_));
  NA2        g0882(.A(new_new_n904_), .B(i_11_), .Y(new_new_n905_));
  AN2        g0883(.A(new_new_n98_), .B(new_new_n245_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n769_), .B(new_new_n336_), .Y(new_new_n907_));
  AOI210     g0885(.A0(new_new_n500_), .A1(new_new_n88_), .B0(new_new_n59_), .Y(new_new_n908_));
  OAI220     g0886(.A0(new_new_n908_), .A1(new_new_n907_), .B0(new_new_n678_), .B1(new_new_n561_), .Y(new_new_n909_));
  NO2        g0887(.A(new_new_n256_), .B(new_new_n155_), .Y(new_new_n910_));
  NA2        g0888(.A(i_0_), .B(i_10_), .Y(new_new_n911_));
  OAI210     g0889(.A0(new_new_n911_), .A1(new_new_n87_), .B0(new_new_n564_), .Y(new_new_n912_));
  NO4        g0890(.A(new_new_n116_), .B(new_new_n59_), .C(new_new_n688_), .D(i_5_), .Y(new_new_n913_));
  AO220      g0891(.A0(new_new_n913_), .A1(new_new_n912_), .B0(new_new_n910_), .B1(i_6_), .Y(new_new_n914_));
  AOI220     g0892(.A0(new_new_n342_), .A1(new_new_n100_), .B0(new_new_n189_), .B1(new_new_n85_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n589_), .B(i_4_), .Y(new_new_n916_));
  NA2        g0894(.A(new_new_n192_), .B(new_new_n207_), .Y(new_new_n917_));
  OAI220     g0895(.A0(new_new_n917_), .A1(new_new_n907_), .B0(new_new_n916_), .B1(new_new_n915_), .Y(new_new_n918_));
  NO4        g0896(.A(new_new_n918_), .B(new_new_n914_), .C(new_new_n909_), .D(new_new_n906_), .Y(new_new_n919_));
  NA4        g0897(.A(new_new_n919_), .B(new_new_n905_), .C(new_new_n902_), .D(new_new_n900_), .Y(new_new_n920_));
  NO2        g0898(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n921_));
  NA2        g0899(.A(i_11_), .B(i_9_), .Y(new_new_n922_));
  NO3        g0900(.A(i_12_), .B(new_new_n922_), .C(new_new_n621_), .Y(new_new_n923_));
  AN2        g0901(.A(new_new_n923_), .B(new_new_n921_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n49_), .B(i_7_), .Y(new_new_n925_));
  NA2        g0903(.A(new_new_n409_), .B(new_new_n182_), .Y(new_new_n926_));
  NA3        g0904(.A(new_new_n926_), .B(new_new_n476_), .C(new_new_n162_), .Y(new_new_n927_));
  NO2        g0905(.A(new_new_n922_), .B(new_new_n74_), .Y(new_new_n928_));
  NO2        g0906(.A(new_new_n178_), .B(i_0_), .Y(new_new_n929_));
  INV        g0907(.A(new_new_n929_), .Y(new_new_n930_));
  NA2        g0908(.A(new_new_n489_), .B(new_new_n232_), .Y(new_new_n931_));
  AOI210     g0909(.A0(new_new_n385_), .A1(new_new_n42_), .B0(new_new_n420_), .Y(new_new_n932_));
  OAI220     g0910(.A0(new_new_n932_), .A1(new_new_n889_), .B0(new_new_n931_), .B1(new_new_n930_), .Y(new_new_n933_));
  NO3        g0911(.A(new_new_n933_), .B(new_new_n927_), .C(new_new_n924_), .Y(new_new_n934_));
  NA2        g0912(.A(new_new_n677_), .B(new_new_n123_), .Y(new_new_n935_));
  NO2        g0913(.A(i_6_), .B(new_new_n935_), .Y(new_new_n936_));
  AOI210     g0914(.A0(new_new_n465_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n174_), .B(new_new_n105_), .Y(new_new_n938_));
  NOi32      g0916(.An(new_new_n937_), .Bn(new_new_n192_), .C(new_new_n938_), .Y(new_new_n939_));
  NO2        g0917(.A(new_new_n939_), .B(new_new_n936_), .Y(new_new_n940_));
  NOi21      g0918(.An(i_7_), .B(i_5_), .Y(new_new_n941_));
  OR2        g0919(.A(new_new_n938_), .B(new_new_n537_), .Y(new_new_n942_));
  NO3        g0920(.A(new_new_n416_), .B(new_new_n374_), .C(new_new_n371_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n266_), .B(new_new_n325_), .Y(new_new_n944_));
  NO2        g0922(.A(new_new_n748_), .B(new_new_n261_), .Y(new_new_n945_));
  AOI210     g0923(.A0(new_new_n945_), .A1(new_new_n944_), .B0(new_new_n943_), .Y(new_new_n946_));
  NA4        g0924(.A(new_new_n946_), .B(new_new_n942_), .C(new_new_n940_), .D(new_new_n934_), .Y(new_new_n947_));
  NO2        g0925(.A(new_new_n897_), .B(new_new_n241_), .Y(new_new_n948_));
  AN2        g0926(.A(new_new_n341_), .B(new_new_n336_), .Y(new_new_n949_));
  AO220      g0927(.A0(new_new_n949_), .A1(new_new_n893_), .B0(new_new_n357_), .B1(new_new_n27_), .Y(new_new_n950_));
  OAI210     g0928(.A0(new_new_n950_), .A1(new_new_n948_), .B0(i_10_), .Y(new_new_n951_));
  NO2        g0929(.A(new_new_n866_), .B(new_new_n324_), .Y(new_new_n952_));
  OA210      g0930(.A0(new_new_n489_), .A1(new_new_n225_), .B0(new_new_n488_), .Y(new_new_n953_));
  NA2        g0931(.A(new_new_n952_), .B(new_new_n928_), .Y(new_new_n954_));
  NO2        g0932(.A(new_new_n259_), .B(new_new_n47_), .Y(new_new_n955_));
  NO2        g0933(.A(new_new_n955_), .B(new_new_n191_), .Y(new_new_n956_));
  NA2        g0934(.A(new_new_n956_), .B(new_new_n489_), .Y(new_new_n957_));
  NA2        g0935(.A(new_new_n722_), .B(new_new_n568_), .Y(new_new_n958_));
  NAi21      g0936(.An(i_9_), .B(i_5_), .Y(new_new_n959_));
  NO2        g0937(.A(new_new_n959_), .B(new_new_n416_), .Y(new_new_n960_));
  NO2        g0938(.A(new_new_n617_), .B(new_new_n107_), .Y(new_new_n961_));
  AOI220     g0939(.A0(new_new_n961_), .A1(i_0_), .B0(new_new_n960_), .B1(new_new_n639_), .Y(new_new_n962_));
  OAI220     g0940(.A0(new_new_n962_), .A1(new_new_n87_), .B0(new_new_n958_), .B1(new_new_n175_), .Y(new_new_n963_));
  NO2        g0941(.A(new_new_n963_), .B(new_new_n542_), .Y(new_new_n964_));
  NA4        g0942(.A(new_new_n964_), .B(new_new_n957_), .C(new_new_n954_), .D(new_new_n951_), .Y(new_new_n965_));
  NO3        g0943(.A(new_new_n965_), .B(new_new_n947_), .C(new_new_n920_), .Y(new_new_n966_));
  NO2        g0944(.A(i_0_), .B(new_new_n748_), .Y(new_new_n967_));
  NA2        g0945(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n968_));
  NA2        g0946(.A(new_new_n911_), .B(new_new_n968_), .Y(new_new_n969_));
  NO3        g0947(.A(new_new_n107_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n970_));
  AO220      g0948(.A0(new_new_n970_), .A1(new_new_n969_), .B0(new_new_n967_), .B1(new_new_n177_), .Y(new_new_n971_));
  AOI210     g0949(.A0(new_new_n822_), .A1(new_new_n708_), .B0(new_new_n938_), .Y(new_new_n972_));
  AOI210     g0950(.A0(new_new_n971_), .A1(new_new_n359_), .B0(new_new_n972_), .Y(new_new_n973_));
  NA2        g0951(.A(new_new_n757_), .B(new_new_n148_), .Y(new_new_n974_));
  INV        g0952(.A(new_new_n974_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n975_), .B(new_new_n695_), .C(new_new_n74_), .Y(new_new_n976_));
  NO2        g0954(.A(new_new_n839_), .B(new_new_n416_), .Y(new_new_n977_));
  NA3        g0955(.A(new_new_n868_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n978_));
  NA2        g0956(.A(new_new_n869_), .B(i_9_), .Y(new_new_n979_));
  AOI210     g0957(.A0(new_new_n978_), .A1(new_new_n516_), .B0(new_new_n979_), .Y(new_new_n980_));
  OAI210     g0958(.A0(new_new_n246_), .A1(i_9_), .B0(new_new_n231_), .Y(new_new_n981_));
  AOI210     g0959(.A0(new_new_n981_), .A1(new_new_n903_), .B0(new_new_n155_), .Y(new_new_n982_));
  NO3        g0960(.A(new_new_n982_), .B(new_new_n980_), .C(new_new_n977_), .Y(new_new_n983_));
  NA3        g0961(.A(new_new_n983_), .B(new_new_n976_), .C(new_new_n973_), .Y(new_new_n984_));
  NA2        g0962(.A(new_new_n949_), .B(new_new_n387_), .Y(new_new_n985_));
  AOI210     g0963(.A0(new_new_n306_), .A1(new_new_n164_), .B0(new_new_n985_), .Y(new_new_n986_));
  NA3        g0964(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n987_));
  NA2        g0965(.A(new_new_n925_), .B(new_new_n505_), .Y(new_new_n988_));
  AOI210     g0966(.A0(new_new_n987_), .A1(new_new_n164_), .B0(new_new_n988_), .Y(new_new_n989_));
  NO2        g0967(.A(new_new_n989_), .B(new_new_n986_), .Y(new_new_n990_));
  NO3        g0968(.A(new_new_n911_), .B(new_new_n888_), .C(new_new_n194_), .Y(new_new_n991_));
  AOI220     g0969(.A0(new_new_n991_), .A1(i_11_), .B0(new_new_n590_), .B1(new_new_n76_), .Y(new_new_n992_));
  NO3        g0970(.A(new_new_n213_), .B(new_new_n398_), .C(i_0_), .Y(new_new_n993_));
  OAI210     g0971(.A0(new_new_n993_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n994_));
  INV        g0972(.A(new_new_n221_), .Y(new_new_n995_));
  OAI220     g0973(.A0(new_new_n554_), .A1(new_new_n141_), .B0(new_new_n661_), .B1(new_new_n634_), .Y(new_new_n996_));
  NA3        g0974(.A(new_new_n996_), .B(new_new_n411_), .C(new_new_n995_), .Y(new_new_n997_));
  NA4        g0975(.A(new_new_n997_), .B(new_new_n994_), .C(new_new_n992_), .D(new_new_n990_), .Y(new_new_n998_));
  AOI220     g0976(.A0(new_new_n941_), .A1(new_new_n505_), .B0(new_new_n868_), .B1(new_new_n165_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n362_), .B(new_new_n179_), .Y(new_new_n1000_));
  OR2        g0978(.A(new_new_n1000_), .B(new_new_n999_), .Y(new_new_n1001_));
  AOI210     g0979(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n178_), .Y(new_new_n1002_));
  NA2        g0980(.A(new_new_n1002_), .B(new_new_n953_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n631_), .B(new_new_n189_), .C(new_new_n85_), .Y(new_new_n1004_));
  INV        g0982(.A(new_new_n1004_), .Y(new_new_n1005_));
  NO3        g0983(.A(new_new_n878_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n1006_));
  NA2        g0984(.A(new_new_n510_), .B(new_new_n503_), .Y(new_new_n1007_));
  NO3        g0985(.A(new_new_n1007_), .B(new_new_n1006_), .C(new_new_n1005_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n404_), .B(new_new_n174_), .C(new_new_n173_), .Y(new_new_n1009_));
  NA3        g0987(.A(new_new_n404_), .B(new_new_n343_), .C(new_new_n223_), .Y(new_new_n1010_));
  OAI210     g0988(.A0(new_new_n883_), .A1(new_new_n665_), .B0(new_new_n1010_), .Y(new_new_n1011_));
  NOi31      g0989(.An(new_new_n403_), .B(new_new_n968_), .C(new_new_n241_), .Y(new_new_n1012_));
  NO3        g0990(.A(new_new_n922_), .B(new_new_n221_), .C(new_new_n194_), .Y(new_new_n1013_));
  NO4        g0991(.A(new_new_n1013_), .B(new_new_n1012_), .C(new_new_n1011_), .D(new_new_n1074_), .Y(new_new_n1014_));
  NA4        g0992(.A(new_new_n1014_), .B(new_new_n1008_), .C(new_new_n1003_), .D(new_new_n1001_), .Y(new_new_n1015_));
  INV        g0993(.A(new_new_n633_), .Y(new_new_n1016_));
  NO3        g0994(.A(new_new_n1016_), .B(new_new_n580_), .C(new_new_n356_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n87_), .B(i_5_), .Y(new_new_n1018_));
  NA3        g0996(.A(new_new_n869_), .B(new_new_n111_), .C(new_new_n126_), .Y(new_new_n1019_));
  INV        g0997(.A(new_new_n1019_), .Y(new_new_n1020_));
  AOI210     g0998(.A0(new_new_n1020_), .A1(new_new_n1018_), .B0(new_new_n1017_), .Y(new_new_n1021_));
  NAi21      g0999(.An(new_new_n243_), .B(new_new_n244_), .Y(new_new_n1022_));
  NO4        g1000(.A(new_new_n241_), .B(new_new_n213_), .C(i_0_), .D(i_12_), .Y(new_new_n1023_));
  AOI220     g1001(.A0(new_new_n1023_), .A1(new_new_n1022_), .B0(new_new_n816_), .B1(new_new_n179_), .Y(new_new_n1024_));
  AN2        g1002(.A(new_new_n911_), .B(new_new_n155_), .Y(new_new_n1025_));
  NO4        g1003(.A(new_new_n1025_), .B(i_12_), .C(new_new_n665_), .D(new_new_n133_), .Y(new_new_n1026_));
  NA2        g1004(.A(new_new_n1026_), .B(new_new_n221_), .Y(new_new_n1027_));
  NA3        g1005(.A(new_new_n100_), .B(new_new_n594_), .C(i_11_), .Y(new_new_n1028_));
  NO2        g1006(.A(new_new_n1028_), .B(new_new_n157_), .Y(new_new_n1029_));
  NA2        g1007(.A(new_new_n941_), .B(new_new_n487_), .Y(new_new_n1030_));
  NO2        g1008(.A(new_new_n1030_), .B(new_new_n696_), .Y(new_new_n1031_));
  AOI210     g1009(.A0(new_new_n1031_), .A1(new_new_n929_), .B0(new_new_n1029_), .Y(new_new_n1032_));
  NA4        g1010(.A(new_new_n1032_), .B(new_new_n1027_), .C(new_new_n1024_), .D(new_new_n1021_), .Y(new_new_n1033_));
  NO4        g1011(.A(new_new_n1033_), .B(new_new_n1015_), .C(new_new_n998_), .D(new_new_n984_), .Y(new_new_n1034_));
  OAI210     g1012(.A0(new_new_n842_), .A1(new_new_n835_), .B0(new_new_n37_), .Y(new_new_n1035_));
  NA3        g1013(.A(new_new_n937_), .B(new_new_n382_), .C(i_5_), .Y(new_new_n1036_));
  NA3        g1014(.A(new_new_n1036_), .B(new_new_n1035_), .C(new_new_n629_), .Y(new_new_n1037_));
  NA2        g1015(.A(new_new_n1037_), .B(new_new_n210_), .Y(new_new_n1038_));
  AN2        g1016(.A(new_new_n720_), .B(new_new_n383_), .Y(new_new_n1039_));
  NA2        g1017(.A(new_new_n190_), .B(new_new_n192_), .Y(new_new_n1040_));
  AO210      g1018(.A0(new_new_n1039_), .A1(new_new_n33_), .B0(new_new_n1040_), .Y(new_new_n1041_));
  OAI210     g1019(.A0(new_new_n633_), .A1(new_new_n631_), .B0(new_new_n324_), .Y(new_new_n1042_));
  NAi31      g1020(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1043_));
  AOI210     g1021(.A0(new_new_n119_), .A1(new_new_n71_), .B0(new_new_n1043_), .Y(new_new_n1044_));
  NO2        g1022(.A(new_new_n1044_), .B(new_new_n662_), .Y(new_new_n1045_));
  NA3        g1023(.A(new_new_n1045_), .B(new_new_n1042_), .C(new_new_n1041_), .Y(new_new_n1046_));
  NO2        g1024(.A(new_new_n479_), .B(new_new_n272_), .Y(new_new_n1047_));
  NO4        g1025(.A(new_new_n234_), .B(new_new_n147_), .C(new_new_n699_), .D(new_new_n37_), .Y(new_new_n1048_));
  NO3        g1026(.A(new_new_n1048_), .B(new_new_n1047_), .C(new_new_n904_), .Y(new_new_n1049_));
  OAI210     g1027(.A0(new_new_n1028_), .A1(new_new_n150_), .B0(new_new_n1049_), .Y(new_new_n1050_));
  AOI210     g1028(.A0(new_new_n1046_), .A1(new_new_n49_), .B0(new_new_n1050_), .Y(new_new_n1051_));
  AOI210     g1029(.A0(new_new_n1051_), .A1(new_new_n1038_), .B0(new_new_n74_), .Y(new_new_n1052_));
  NO2        g1030(.A(new_new_n587_), .B(new_new_n394_), .Y(new_new_n1053_));
  NO2        g1031(.A(new_new_n1053_), .B(new_new_n777_), .Y(new_new_n1054_));
  NA2        g1032(.A(new_new_n266_), .B(new_new_n58_), .Y(new_new_n1055_));
  AOI220     g1033(.A0(new_new_n1055_), .A1(new_new_n77_), .B0(new_new_n357_), .B1(new_new_n258_), .Y(new_new_n1056_));
  NO2        g1034(.A(new_new_n1056_), .B(new_new_n238_), .Y(new_new_n1057_));
  NA3        g1035(.A(new_new_n98_), .B(new_new_n313_), .C(new_new_n31_), .Y(new_new_n1058_));
  INV        g1036(.A(new_new_n1058_), .Y(new_new_n1059_));
  NO2        g1037(.A(new_new_n1059_), .B(new_new_n1057_), .Y(new_new_n1060_));
  OAI210     g1038(.A0(new_new_n274_), .A1(new_new_n160_), .B0(new_new_n88_), .Y(new_new_n1061_));
  NO2        g1039(.A(new_new_n1061_), .B(i_11_), .Y(new_new_n1062_));
  NO4        g1040(.A(new_new_n959_), .B(new_new_n493_), .C(new_new_n255_), .D(new_new_n254_), .Y(new_new_n1063_));
  NO2        g1041(.A(new_new_n1063_), .B(new_new_n584_), .Y(new_new_n1064_));
  NO2        g1042(.A(new_new_n1064_), .B(new_new_n41_), .Y(new_new_n1065_));
  NO2        g1043(.A(new_new_n1065_), .B(new_new_n1062_), .Y(new_new_n1066_));
  OAI210     g1044(.A0(new_new_n1060_), .A1(i_4_), .B0(new_new_n1066_), .Y(new_new_n1067_));
  NO3        g1045(.A(new_new_n1067_), .B(new_new_n1054_), .C(new_new_n1052_), .Y(new_new_n1068_));
  NA4        g1046(.A(new_new_n1068_), .B(new_new_n1034_), .C(new_new_n966_), .D(new_new_n896_), .Y(zz04));
  INV        g1047(.A(new_new_n721_), .Y(new_new_n1072_));
  INV        g1048(.A(i_2_), .Y(new_new_n1073_));
  INV        g1049(.A(new_new_n1009_), .Y(new_new_n1074_));
endmodule


