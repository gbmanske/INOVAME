//Benchmark atmr_intb_466_0.5

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n89_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n180_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n478_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o00(.A(x11), .Y(ori_ori_n23_));
  NA2        o01(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o02(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o03(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o04(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o05(.A(x02), .Y(ori_ori_n28_));
  INV        o06(.A(x10), .Y(ori_ori_n29_));
  NA2        o07(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o08(.A(x03), .Y(ori_ori_n31_));
  NA2        o09(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o10(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o11(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o12(.A(x04), .Y(ori_ori_n35_));
  INV        o13(.A(x08), .Y(ori_ori_n36_));
  NA2        o14(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o15(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o16(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o17(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o18(.A(x05), .Y(ori_ori_n41_));
  NO2        o19(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o20(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o21(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o22(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o23(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o24(.A(x01), .Y(ori_ori_n47_));
  INV        o25(.A(x06), .Y(ori_ori_n48_));
  INV        o26(.A(x09), .Y(ori_ori_n49_));
  NO2        o27(.A(x10), .B(x02), .Y(ori_ori_n50_));
  INV        o28(.A(x00), .Y(ori_ori_n51_));
  INV        o29(.A(x07), .Y(ori_ori_n52_));
  NO2        o30(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n53_));
  NO2        o31(.A(x08), .B(x01), .Y(ori_ori_n54_));
  OAI210     o32(.A0(ori_ori_n54_), .A1(ori_ori_n53_), .B0(ori_ori_n35_), .Y(ori_ori_n55_));
  INV        o33(.A(ori_ori_n55_), .Y(ori_ori_n56_));
  NA2        o34(.A(x11), .B(x00), .Y(ori_ori_n57_));
  NO2        o35(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n58_));
  NOi21      o36(.An(ori_ori_n57_), .B(ori_ori_n58_), .Y(ori_ori_n59_));
  INV        o37(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  NO2        o38(.A(ori_ori_n60_), .B(x07), .Y(ori_ori_n61_));
  INV        o39(.A(ori_ori_n61_), .Y(ori01));
  INV        o40(.A(x12), .Y(ori_ori_n63_));
  NA2        o41(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n64_));
  NA2        o42(.A(x10), .B(ori_ori_n51_), .Y(ori_ori_n65_));
  NA2        o43(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  NO2        o44(.A(x09), .B(x05), .Y(ori_ori_n67_));
  NA2        o45(.A(ori_ori_n67_), .B(ori_ori_n47_), .Y(ori_ori_n68_));
  NO2        o46(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n69_));
  NA2        o47(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n70_));
  INV        o48(.A(ori_ori_n70_), .Y(ori_ori_n71_));
  NO2        o49(.A(ori_ori_n49_), .B(x03), .Y(ori_ori_n72_));
  NA2        o50(.A(x13), .B(ori_ori_n63_), .Y(ori_ori_n73_));
  INV        o51(.A(ori_ori_n59_), .Y(ori_ori_n74_));
  NO2        o52(.A(ori_ori_n74_), .B(x07), .Y(ori_ori_n75_));
  INV        o53(.A(ori_ori_n75_), .Y(ori_ori_n76_));
  OAI210     o54(.A0(ori_ori_n71_), .A1(ori_ori_n52_), .B0(ori_ori_n76_), .Y(ori02));
  INV        o55(.A(ori_ori_n66_), .Y(ori_ori_n78_));
  NA2        o56(.A(ori_ori_n78_), .B(ori_ori_n48_), .Y(ori_ori_n79_));
  NO2        o57(.A(ori_ori_n69_), .B(ori_ori_n50_), .Y(ori_ori_n80_));
  INV        o58(.A(ori_ori_n80_), .Y(ori_ori_n81_));
  NA2        o59(.A(ori_ori_n81_), .B(x06), .Y(ori_ori_n82_));
  NA2        o60(.A(ori_ori_n82_), .B(ori_ori_n79_), .Y(ori_ori_n83_));
  INV        o61(.A(ori_ori_n83_), .Y(ori03));
  OR2        o62(.A(ori_ori_n42_), .B(ori_ori_n72_), .Y(ori_ori_n85_));
  AOI210     o63(.A0(ori_ori_n35_), .A1(ori_ori_n63_), .B0(ori_ori_n85_), .Y(ori_ori_n86_));
  NA2        o64(.A(ori_ori_n86_), .B(x05), .Y(ori_ori_n87_));
  NA2        o65(.A(ori_ori_n68_), .B(ori_ori_n87_), .Y(ori04));
  NO2        o66(.A(ori_ori_n56_), .B(ori_ori_n39_), .Y(ori_ori_n89_));
  XO2        o67(.A(ori_ori_n89_), .B(ori_ori_n73_), .Y(ori05));
  ZERO       o68(.Y(ori06));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  INV        m017(.A(x05), .Y(mai_mai_n40_));
  NO2        m018(.A(x09), .B(x02), .Y(mai_mai_n41_));
  NO2        m019(.A(mai_mai_n39_), .B(mai_mai_n34_), .Y(mai00));
  INV        m020(.A(x01), .Y(mai_mai_n43_));
  INV        m021(.A(x06), .Y(mai_mai_n44_));
  NO3        m022(.A(x02), .B(x11), .C(x09), .Y(mai_mai_n45_));
  INV        m023(.A(x09), .Y(mai_mai_n46_));
  NO2        m024(.A(x10), .B(x02), .Y(mai_mai_n47_));
  NO2        m025(.A(x02), .B(x07), .Y(mai_mai_n48_));
  OAI210     m026(.A0(mai_mai_n48_), .A1(mai_mai_n45_), .B0(mai_mai_n43_), .Y(mai_mai_n49_));
  NOi21      m027(.An(x01), .B(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x00), .Y(mai_mai_n51_));
  NO2        m029(.A(mai_mai_n46_), .B(mai_mai_n51_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(mai_mai_n50_), .Y(mai_mai_n53_));
  NA2        m031(.A(x09), .B(mai_mai_n51_), .Y(mai_mai_n54_));
  INV        m032(.A(x07), .Y(mai_mai_n55_));
  NA2        m033(.A(mai_mai_n55_), .B(mai_mai_n44_), .Y(mai_mai_n56_));
  OAI210     m034(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n56_), .Y(mai_mai_n57_));
  AOI220     m035(.A0(mai_mai_n57_), .A1(mai_mai_n53_), .B0(mai_mai_n53_), .B1(mai_mai_n31_), .Y(mai_mai_n58_));
  AOI210     m036(.A0(mai_mai_n58_), .A1(mai_mai_n49_), .B0(x05), .Y(mai_mai_n59_));
  NO2        m037(.A(mai_mai_n55_), .B(mai_mai_n23_), .Y(mai_mai_n60_));
  OAI210     m038(.A0(x02), .A1(mai_mai_n60_), .B0(x03), .Y(mai_mai_n61_));
  NO2        m039(.A(x09), .B(mai_mai_n40_), .Y(mai_mai_n62_));
  NO2        m040(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n63_));
  NO2        m041(.A(x08), .B(x01), .Y(mai_mai_n64_));
  OAI210     m042(.A0(mai_mai_n64_), .A1(mai_mai_n63_), .B0(mai_mai_n35_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n46_), .B(mai_mai_n36_), .Y(mai_mai_n66_));
  INV        m044(.A(mai_mai_n65_), .Y(mai_mai_n67_));
  AN2        m045(.A(mai_mai_n67_), .B(mai_mai_n61_), .Y(mai_mai_n68_));
  INV        m046(.A(mai_mai_n65_), .Y(mai_mai_n69_));
  NO2        m047(.A(x06), .B(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x11), .B(x00), .Y(mai_mai_n71_));
  NO2        m049(.A(x11), .B(mai_mai_n43_), .Y(mai_mai_n72_));
  NOi21      m050(.An(mai_mai_n71_), .B(mai_mai_n72_), .Y(mai_mai_n73_));
  AOI210     m051(.A0(mai_mai_n70_), .A1(mai_mai_n69_), .B0(mai_mai_n73_), .Y(mai_mai_n74_));
  NO2        m052(.A(x02), .B(x11), .Y(mai_mai_n75_));
  NOi21      m053(.An(x01), .B(x10), .Y(mai_mai_n76_));
  NO2        m054(.A(mai_mai_n29_), .B(mai_mai_n51_), .Y(mai_mai_n77_));
  NO3        m055(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(x06), .Y(mai_mai_n78_));
  AOI220     m056(.A0(mai_mai_n78_), .A1(mai_mai_n27_), .B0(mai_mai_n75_), .B1(mai_mai_n69_), .Y(mai_mai_n79_));
  OAI210     m057(.A0(mai_mai_n74_), .A1(x07), .B0(mai_mai_n79_), .Y(mai_mai_n80_));
  NO3        m058(.A(mai_mai_n80_), .B(mai_mai_n68_), .C(mai_mai_n59_), .Y(mai01));
  INV        m059(.A(x12), .Y(mai_mai_n82_));
  INV        m060(.A(x13), .Y(mai_mai_n83_));
  NA2        m061(.A(mai_mai_n76_), .B(mai_mai_n28_), .Y(mai_mai_n84_));
  NO2        m062(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n85_));
  NA2        m063(.A(mai_mai_n29_), .B(mai_mai_n43_), .Y(mai_mai_n86_));
  NA2        m064(.A(x10), .B(mai_mai_n51_), .Y(mai_mai_n87_));
  NA2        m065(.A(mai_mai_n87_), .B(mai_mai_n86_), .Y(mai_mai_n88_));
  NA2        m066(.A(mai_mai_n46_), .B(x05), .Y(mai_mai_n89_));
  NO2        m067(.A(mai_mai_n54_), .B(x05), .Y(mai_mai_n90_));
  NO2        m068(.A(mai_mai_n46_), .B(mai_mai_n40_), .Y(mai_mai_n91_));
  NA2        m069(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n92_));
  NO2        m070(.A(x09), .B(x05), .Y(mai_mai_n93_));
  NA2        m071(.A(mai_mai_n93_), .B(mai_mai_n43_), .Y(mai_mai_n94_));
  NA2        m072(.A(x09), .B(x00), .Y(mai_mai_n95_));
  NA2        m073(.A(mai_mai_n85_), .B(mai_mai_n95_), .Y(mai_mai_n96_));
  NO2        m074(.A(x03), .B(x02), .Y(mai_mai_n97_));
  NA2        m075(.A(mai_mai_n65_), .B(mai_mai_n83_), .Y(mai_mai_n98_));
  OA210      m076(.A0(x02), .A1(x11), .B0(mai_mai_n191_), .Y(mai_mai_n99_));
  OAI210     m077(.A0(x03), .A1(mai_mai_n23_), .B0(mai_mai_n99_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n101_));
  NA2        m079(.A(x10), .B(x05), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n83_), .B(x12), .Y(mai_mai_n103_));
  AOI210     m081(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n103_), .Y(mai_mai_n104_));
  NA2        m082(.A(mai_mai_n104_), .B(x12), .Y(mai_mai_n105_));
  INV        m083(.A(mai_mai_n105_), .Y(mai_mai_n106_));
  AOI210     m084(.A0(mai_mai_n100_), .A1(mai_mai_n82_), .B0(mai_mai_n106_), .Y(mai_mai_n107_));
  INV        m085(.A(x12), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n51_), .B(mai_mai_n23_), .Y(mai_mai_n109_));
  OAI210     m087(.A0(mai_mai_n108_), .A1(mai_mai_n51_), .B0(mai_mai_n109_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n46_), .B(x03), .Y(mai_mai_n111_));
  INV        m089(.A(mai_mai_n72_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n112_), .B(x12), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n46_), .B(mai_mai_n36_), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n29_), .B(mai_mai_n44_), .Y(mai_mai_n115_));
  NA2        m093(.A(x13), .B(mai_mai_n82_), .Y(mai_mai_n116_));
  NA3        m094(.A(mai_mai_n116_), .B(x12), .C(mai_mai_n73_), .Y(mai_mai_n117_));
  INV        m095(.A(mai_mai_n117_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n113_), .B(mai_mai_n118_), .Y(mai_mai_n119_));
  AOI210     m097(.A0(mai_mai_n119_), .A1(mai_mai_n110_), .B0(x07), .Y(mai_mai_n120_));
  NO2        m098(.A(x08), .B(x05), .Y(mai_mai_n121_));
  NO2        m099(.A(x12), .B(x02), .Y(mai_mai_n122_));
  INV        m100(.A(mai_mai_n122_), .Y(mai_mai_n123_));
  NO2        m101(.A(mai_mai_n123_), .B(mai_mai_n112_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n46_), .B(mai_mai_n40_), .Y(mai_mai_n125_));
  NO2        m103(.A(mai_mai_n125_), .B(x01), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n83_), .B(x04), .Y(mai_mai_n127_));
  NO3        m105(.A(mai_mai_n71_), .B(x12), .C(x03), .Y(mai_mai_n128_));
  NO3        m106(.A(mai_mai_n128_), .B(mai_mai_n124_), .C(mai_mai_n120_), .Y(mai_mai_n129_));
  OAI210     m107(.A0(mai_mai_n107_), .A1(mai_mai_n55_), .B0(mai_mai_n129_), .Y(mai02));
  INV        m108(.A(mai_mai_n89_), .Y(mai_mai_n131_));
  OAI210     m109(.A0(mai_mai_n190_), .A1(mai_mai_n131_), .B0(mai_mai_n102_), .Y(mai_mai_n132_));
  INV        m110(.A(mai_mai_n102_), .Y(mai_mai_n133_));
  AOI220     m111(.A0(x09), .A1(mai_mai_n133_), .B0(mai_mai_n98_), .B1(mai_mai_n97_), .Y(mai_mai_n134_));
  AOI210     m112(.A0(mai_mai_n134_), .A1(mai_mai_n132_), .B0(mai_mai_n44_), .Y(mai_mai_n135_));
  AOI220     m113(.A0(mai_mai_n121_), .A1(mai_mai_n52_), .B0(mai_mai_n50_), .B1(mai_mai_n36_), .Y(mai_mai_n136_));
  NOi21      m114(.An(x04), .B(mai_mai_n136_), .Y(mai_mai_n137_));
  AOI210     m115(.A0(x13), .A1(mai_mai_n62_), .B0(mai_mai_n137_), .Y(mai_mai_n138_));
  AOI210     m116(.A0(mai_mai_n138_), .A1(x02), .B0(mai_mai_n92_), .Y(mai_mai_n139_));
  NO2        m117(.A(mai_mai_n115_), .B(mai_mai_n43_), .Y(mai_mai_n140_));
  INV        m118(.A(mai_mai_n140_), .Y(mai_mai_n141_));
  OAI210     m119(.A0(mai_mai_n44_), .A1(mai_mai_n192_), .B0(mai_mai_n77_), .Y(mai_mai_n142_));
  NA3        m120(.A(mai_mai_n77_), .B(mai_mai_n64_), .C(mai_mai_n111_), .Y(mai_mai_n143_));
  NA3        m121(.A(mai_mai_n76_), .B(mai_mai_n63_), .C(mai_mai_n41_), .Y(mai_mai_n144_));
  AOI210     m122(.A0(mai_mai_n144_), .A1(mai_mai_n143_), .B0(x04), .Y(mai_mai_n145_));
  INV        m123(.A(mai_mai_n97_), .Y(mai_mai_n146_));
  OAI210     m124(.A0(mai_mai_n146_), .A1(mai_mai_n88_), .B0(mai_mai_n84_), .Y(mai_mai_n147_));
  AOI210     m125(.A0(mai_mai_n147_), .A1(x13), .B0(mai_mai_n145_), .Y(mai_mai_n148_));
  NA3        m126(.A(mai_mai_n148_), .B(mai_mai_n142_), .C(mai_mai_n141_), .Y(mai_mai_n149_));
  NO3        m127(.A(mai_mai_n149_), .B(mai_mai_n139_), .C(mai_mai_n135_), .Y(mai_mai_n150_));
  NA2        m128(.A(mai_mai_n91_), .B(x03), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n127_), .B(mai_mai_n82_), .Y(mai_mai_n152_));
  NA2        m130(.A(mai_mai_n82_), .B(mai_mai_n40_), .Y(mai_mai_n153_));
  NA3        m131(.A(mai_mai_n153_), .B(mai_mai_n152_), .C(mai_mai_n88_), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n154_), .B(mai_mai_n44_), .Y(mai_mai_n155_));
  INV        m133(.A(mai_mai_n114_), .Y(mai_mai_n156_));
  NA2        m134(.A(mai_mai_n103_), .B(x04), .Y(mai_mai_n157_));
  NO3        m135(.A(mai_mai_n103_), .B(mai_mai_n101_), .C(mai_mai_n47_), .Y(mai_mai_n158_));
  NA2        m136(.A(x12), .B(mai_mai_n158_), .Y(mai_mai_n159_));
  NA2        m137(.A(mai_mai_n159_), .B(x06), .Y(mai_mai_n160_));
  NA2        m138(.A(mai_mai_n160_), .B(mai_mai_n155_), .Y(mai_mai_n161_));
  OAI210     m139(.A0(mai_mai_n150_), .A1(x12), .B0(mai_mai_n161_), .Y(mai03));
  OR2        m140(.A(mai_mai_n41_), .B(mai_mai_n111_), .Y(mai_mai_n163_));
  AOI210     m141(.A0(mai_mai_n98_), .A1(mai_mai_n82_), .B0(mai_mai_n163_), .Y(mai_mai_n164_));
  AO210      m142(.A0(mai_mai_n156_), .A1(mai_mai_n66_), .B0(mai_mai_n157_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n103_), .B(mai_mai_n97_), .Y(mai_mai_n166_));
  NA2        m144(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  OAI210     m145(.A0(mai_mai_n167_), .A1(mai_mai_n164_), .B0(x05), .Y(mai_mai_n168_));
  NA2        m146(.A(mai_mai_n163_), .B(x05), .Y(mai_mai_n169_));
  NO2        m147(.A(x04), .B(mai_mai_n169_), .Y(mai_mai_n170_));
  OAI220     m148(.A0(x05), .A1(mai_mai_n53_), .B0(x02), .B1(mai_mai_n136_), .Y(mai_mai_n171_));
  OAI210     m149(.A0(mai_mai_n171_), .A1(mai_mai_n170_), .B0(mai_mai_n82_), .Y(mai_mai_n172_));
  AOI210     m150(.A0(mai_mai_n94_), .A1(mai_mai_n54_), .B0(mai_mai_n38_), .Y(mai_mai_n173_));
  OAI220     m151(.A0(mai_mai_n54_), .A1(mai_mai_n37_), .B0(mai_mai_n96_), .B1(x13), .Y(mai_mai_n174_));
  OAI210     m152(.A0(mai_mai_n174_), .A1(mai_mai_n173_), .B0(x04), .Y(mai_mai_n175_));
  NO3        m153(.A(mai_mai_n153_), .B(mai_mai_n65_), .C(mai_mai_n53_), .Y(mai_mai_n176_));
  NO2        m154(.A(mai_mai_n82_), .B(mai_mai_n94_), .Y(mai_mai_n177_));
  NO3        m155(.A(mai_mai_n90_), .B(mai_mai_n177_), .C(mai_mai_n176_), .Y(mai_mai_n178_));
  NA4        m156(.A(mai_mai_n178_), .B(mai_mai_n175_), .C(mai_mai_n172_), .D(mai_mai_n168_), .Y(mai04));
  NO2        m157(.A(mai_mai_n69_), .B(mai_mai_n39_), .Y(mai_mai_n180_));
  XO2        m158(.A(mai_mai_n180_), .B(mai_mai_n116_), .Y(mai05));
  NOi21      m159(.An(mai_mai_n151_), .B(mai_mai_n90_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n89_), .B(mai_mai_n28_), .Y(mai_mai_n183_));
  NO2        m161(.A(mai_mai_n183_), .B(mai_mai_n126_), .Y(mai_mai_n184_));
  NA3        m162(.A(mai_mai_n184_), .B(mai_mai_n182_), .C(mai_mai_n152_), .Y(mai_mai_n185_));
  NA2        m163(.A(x14), .B(mai_mai_n185_), .Y(mai_mai_n186_));
  INV        m164(.A(mai_mai_n186_), .Y(mai06));
  INV        m165(.A(mai_mai_n32_), .Y(mai_mai_n190_));
  INV        m166(.A(mai_mai_n97_), .Y(mai_mai_n191_));
  INV        m167(.A(x03), .Y(mai_mai_n192_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men05));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men05), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  AOI220     u039(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n61_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  OAI220     u042(.A0(men_men_n64_), .A1(men_men_n58_), .B0(men_men_n62_), .B1(men_men_n60_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n30_), .A1(x11), .B0(men_men_n66_), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n59_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  NA2        u048(.A(x09), .B(x05), .Y(men_men_n71_));
  NA2        u049(.A(x10), .B(x06), .Y(men_men_n72_));
  NA3        u050(.A(men_men_n72_), .B(men_men_n71_), .C(men_men_n28_), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n74_));
  NA2        u052(.A(men_men_n73_), .B(x03), .Y(men_men_n75_));
  NOi31      u053(.An(x08), .B(x04), .C(x00), .Y(men_men_n76_));
  NO2        u054(.A(x10), .B(x09), .Y(men_men_n77_));
  AOI210     u055(.A0(men_men_n478_), .A1(men_men_n76_), .B0(men_men_n24_), .Y(men_men_n78_));
  NO2        u056(.A(x09), .B(men_men_n41_), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n79_), .B(men_men_n36_), .Y(men_men_n80_));
  OAI210     u058(.A0(men_men_n79_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n81_));
  AOI210     u059(.A0(men_men_n80_), .A1(men_men_n48_), .B0(men_men_n81_), .Y(men_men_n82_));
  NO2        u060(.A(men_men_n36_), .B(x00), .Y(men_men_n83_));
  NO2        u061(.A(x08), .B(x01), .Y(men_men_n84_));
  OAI210     u062(.A0(men_men_n84_), .A1(men_men_n83_), .B0(men_men_n35_), .Y(men_men_n85_));
  NA2        u063(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n86_));
  NO3        u064(.A(men_men_n85_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n87_));
  AN2        u065(.A(men_men_n87_), .B(men_men_n75_), .Y(men_men_n88_));
  INV        u066(.A(men_men_n85_), .Y(men_men_n89_));
  NO2        u067(.A(x06), .B(x05), .Y(men_men_n90_));
  NA2        u068(.A(x11), .B(x00), .Y(men_men_n91_));
  NO2        u069(.A(x11), .B(men_men_n47_), .Y(men_men_n92_));
  NOi21      u070(.An(men_men_n91_), .B(men_men_n92_), .Y(men_men_n93_));
  AOI210     u071(.A0(men_men_n90_), .A1(men_men_n89_), .B0(men_men_n93_), .Y(men_men_n94_));
  NO2        u072(.A(men_men_n53_), .B(x11), .Y(men_men_n95_));
  NOi21      u073(.An(x01), .B(x10), .Y(men_men_n96_));
  NO2        u074(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n97_));
  NO3        u075(.A(men_men_n97_), .B(men_men_n96_), .C(x06), .Y(men_men_n98_));
  AOI220     u076(.A0(men_men_n98_), .A1(men_men_n27_), .B0(men_men_n95_), .B1(men_men_n89_), .Y(men_men_n99_));
  OAI210     u077(.A0(men_men_n94_), .A1(x07), .B0(men_men_n99_), .Y(men_men_n100_));
  NO3        u078(.A(men_men_n100_), .B(men_men_n88_), .C(men_men_n69_), .Y(men01));
  INV        u079(.A(x12), .Y(men_men_n102_));
  INV        u080(.A(x13), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n90_), .B(x01), .Y(men_men_n104_));
  NA2        u082(.A(men_men_n104_), .B(men_men_n70_), .Y(men_men_n105_));
  NA2        u083(.A(x08), .B(x04), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n57_), .Y(men_men_n107_));
  NA2        u085(.A(men_men_n107_), .B(men_men_n105_), .Y(men_men_n108_));
  NA2        u086(.A(men_men_n96_), .B(men_men_n28_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(men_men_n71_), .Y(men_men_n110_));
  NO2        u088(.A(x10), .B(x01), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n29_), .B(x00), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n112_), .B(men_men_n111_), .Y(men_men_n113_));
  NA2        u091(.A(x04), .B(men_men_n28_), .Y(men_men_n114_));
  NO3        u092(.A(men_men_n114_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n115_));
  AOI210     u093(.A0(men_men_n115_), .A1(men_men_n113_), .B0(men_men_n110_), .Y(men_men_n116_));
  AOI210     u094(.A0(men_men_n116_), .A1(men_men_n108_), .B0(men_men_n103_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n56_), .B(x05), .Y(men_men_n118_));
  NOi21      u096(.An(men_men_n118_), .B(men_men_n58_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n35_), .B(x02), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n103_), .B(men_men_n36_), .Y(men_men_n121_));
  NA3        u099(.A(men_men_n121_), .B(men_men_n120_), .C(x06), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n122_), .B(men_men_n119_), .Y(men_men_n123_));
  NO2        u101(.A(men_men_n84_), .B(x13), .Y(men_men_n124_));
  NA2        u102(.A(x09), .B(men_men_n35_), .Y(men_men_n125_));
  NO2        u103(.A(men_men_n125_), .B(men_men_n124_), .Y(men_men_n126_));
  NA2        u104(.A(x13), .B(men_men_n35_), .Y(men_men_n127_));
  NO2        u105(.A(men_men_n127_), .B(x05), .Y(men_men_n128_));
  NO2        u106(.A(men_men_n128_), .B(men_men_n126_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n130_), .B(men_men_n103_), .Y(men_men_n131_));
  AOI210     u109(.A0(men_men_n131_), .A1(men_men_n80_), .B0(men_men_n119_), .Y(men_men_n132_));
  AOI210     u110(.A0(men_men_n132_), .A1(men_men_n129_), .B0(men_men_n72_), .Y(men_men_n133_));
  NA2        u111(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n134_));
  NA2        u112(.A(x10), .B(men_men_n57_), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n135_), .B(men_men_n134_), .Y(men_men_n136_));
  NA2        u114(.A(men_men_n51_), .B(x05), .Y(men_men_n137_));
  NA2        u115(.A(men_men_n36_), .B(x04), .Y(men_men_n138_));
  NA3        u116(.A(men_men_n138_), .B(men_men_n137_), .C(x13), .Y(men_men_n139_));
  NO3        u117(.A(men_men_n130_), .B(men_men_n79_), .C(men_men_n36_), .Y(men_men_n140_));
  NO2        u118(.A(men_men_n60_), .B(x05), .Y(men_men_n141_));
  NOi41      u119(.An(men_men_n139_), .B(men_men_n141_), .C(men_men_n140_), .D(men_men_n136_), .Y(men_men_n142_));
  NO3        u120(.A(men_men_n142_), .B(x06), .C(x03), .Y(men_men_n143_));
  NO4        u121(.A(men_men_n143_), .B(men_men_n133_), .C(men_men_n123_), .D(men_men_n117_), .Y(men_men_n144_));
  NA2        u122(.A(x13), .B(men_men_n36_), .Y(men_men_n145_));
  OAI210     u123(.A0(men_men_n84_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n146_), .B(men_men_n145_), .Y(men_men_n147_));
  NOi21      u125(.An(men_men_n90_), .B(men_men_n57_), .Y(men_men_n148_));
  NO2        u126(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n149_));
  OA210      u127(.A0(men_men_n148_), .A1(men_men_n77_), .B0(men_men_n149_), .Y(men_men_n150_));
  NO2        u128(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n29_), .B(x06), .Y(men_men_n152_));
  AOI210     u130(.A0(men_men_n152_), .A1(men_men_n49_), .B0(men_men_n151_), .Y(men_men_n153_));
  OA210      u131(.A0(men_men_n153_), .A1(men_men_n150_), .B0(men_men_n147_), .Y(men_men_n154_));
  NO2        u132(.A(x09), .B(x05), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n155_), .B(men_men_n47_), .Y(men_men_n156_));
  AOI210     u134(.A0(men_men_n156_), .A1(men_men_n113_), .B0(men_men_n49_), .Y(men_men_n157_));
  NA2        u135(.A(x09), .B(x00), .Y(men_men_n158_));
  NA2        u136(.A(men_men_n118_), .B(men_men_n158_), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n76_), .B(men_men_n51_), .Y(men_men_n160_));
  AOI210     u138(.A0(men_men_n160_), .A1(men_men_n159_), .B0(men_men_n152_), .Y(men_men_n161_));
  NO3        u139(.A(men_men_n161_), .B(men_men_n157_), .C(men_men_n154_), .Y(men_men_n162_));
  NO2        u140(.A(x03), .B(x02), .Y(men_men_n163_));
  NA2        u141(.A(men_men_n85_), .B(men_men_n103_), .Y(men_men_n164_));
  OAI210     u142(.A0(men_men_n164_), .A1(men_men_n119_), .B0(men_men_n163_), .Y(men_men_n165_));
  OA210      u143(.A0(men_men_n162_), .A1(x11), .B0(men_men_n165_), .Y(men_men_n166_));
  OAI210     u144(.A0(men_men_n144_), .A1(men_men_n23_), .B0(men_men_n166_), .Y(men_men_n167_));
  NA2        u145(.A(men_men_n113_), .B(men_men_n40_), .Y(men_men_n168_));
  NA2        u146(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n169_));
  NAi21      u147(.An(x06), .B(x10), .Y(men_men_n170_));
  NOi21      u148(.An(x01), .B(x13), .Y(men_men_n171_));
  NA2        u149(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  OR2        u150(.A(men_men_n172_), .B(men_men_n169_), .Y(men_men_n173_));
  AOI210     u151(.A0(men_men_n173_), .A1(men_men_n168_), .B0(men_men_n41_), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n29_), .B(x03), .Y(men_men_n175_));
  NA2        u153(.A(men_men_n103_), .B(x01), .Y(men_men_n176_));
  NO2        u154(.A(men_men_n176_), .B(x08), .Y(men_men_n177_));
  OAI210     u155(.A0(x05), .A1(men_men_n177_), .B0(men_men_n51_), .Y(men_men_n178_));
  AOI210     u156(.A0(men_men_n178_), .A1(men_men_n175_), .B0(men_men_n48_), .Y(men_men_n179_));
  AOI210     u157(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n180_));
  OAI210     u158(.A0(men_men_n179_), .A1(men_men_n174_), .B0(men_men_n180_), .Y(men_men_n181_));
  NA2        u159(.A(x04), .B(x02), .Y(men_men_n182_));
  NA2        u160(.A(x10), .B(x05), .Y(men_men_n183_));
  NA2        u161(.A(x09), .B(x06), .Y(men_men_n184_));
  AOI210     u162(.A0(men_men_n184_), .A1(men_men_n183_), .B0(men_men_n169_), .Y(men_men_n185_));
  NO2        u163(.A(x09), .B(x01), .Y(men_men_n186_));
  NO3        u164(.A(men_men_n186_), .B(men_men_n111_), .C(men_men_n31_), .Y(men_men_n187_));
  OAI210     u165(.A0(men_men_n187_), .A1(men_men_n185_), .B0(x00), .Y(men_men_n188_));
  NO2        u166(.A(men_men_n118_), .B(x08), .Y(men_men_n189_));
  NA3        u167(.A(men_men_n171_), .B(men_men_n170_), .C(men_men_n51_), .Y(men_men_n190_));
  NA2        u168(.A(men_men_n96_), .B(x05), .Y(men_men_n191_));
  OAI210     u169(.A0(men_men_n191_), .A1(men_men_n121_), .B0(men_men_n190_), .Y(men_men_n192_));
  AOI210     u170(.A0(men_men_n189_), .A1(x06), .B0(men_men_n192_), .Y(men_men_n193_));
  OAI210     u171(.A0(men_men_n193_), .A1(x11), .B0(men_men_n188_), .Y(men_men_n194_));
  NAi21      u172(.An(men_men_n182_), .B(men_men_n194_), .Y(men_men_n195_));
  INV        u173(.A(men_men_n25_), .Y(men_men_n196_));
  NAi21      u174(.An(x13), .B(x00), .Y(men_men_n197_));
  AOI210     u175(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n197_), .Y(men_men_n198_));
  AOI220     u176(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n199_));
  OAI210     u177(.A0(men_men_n183_), .A1(men_men_n35_), .B0(men_men_n199_), .Y(men_men_n200_));
  AN2        u178(.A(men_men_n200_), .B(men_men_n198_), .Y(men_men_n201_));
  AN2        u179(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n97_), .B(x06), .Y(men_men_n203_));
  NO2        u181(.A(men_men_n197_), .B(men_men_n36_), .Y(men_men_n204_));
  INV        u182(.A(men_men_n204_), .Y(men_men_n205_));
  OAI220     u183(.A0(men_men_n205_), .A1(men_men_n184_), .B0(men_men_n203_), .B1(men_men_n202_), .Y(men_men_n206_));
  OAI210     u184(.A0(men_men_n206_), .A1(men_men_n201_), .B0(men_men_n196_), .Y(men_men_n207_));
  NOi21      u185(.An(x09), .B(x00), .Y(men_men_n208_));
  NO3        u186(.A(men_men_n83_), .B(men_men_n208_), .C(men_men_n47_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n209_), .B(men_men_n135_), .Y(men_men_n210_));
  NA2        u188(.A(x10), .B(x08), .Y(men_men_n211_));
  INV        u189(.A(men_men_n211_), .Y(men_men_n212_));
  NA2        u190(.A(x06), .B(x05), .Y(men_men_n213_));
  OAI210     u191(.A0(men_men_n213_), .A1(men_men_n35_), .B0(men_men_n102_), .Y(men_men_n214_));
  AOI210     u192(.A0(men_men_n212_), .A1(men_men_n58_), .B0(men_men_n214_), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n215_), .B(men_men_n210_), .Y(men_men_n216_));
  NO2        u194(.A(men_men_n103_), .B(x12), .Y(men_men_n217_));
  AOI210     u195(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n217_), .Y(men_men_n218_));
  NA2        u196(.A(men_men_n96_), .B(men_men_n51_), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n220_));
  NA2        u198(.A(men_men_n220_), .B(x02), .Y(men_men_n221_));
  NO2        u199(.A(men_men_n221_), .B(men_men_n219_), .Y(men_men_n222_));
  AOI210     u200(.A0(men_men_n218_), .A1(men_men_n216_), .B0(men_men_n222_), .Y(men_men_n223_));
  NA4        u201(.A(men_men_n223_), .B(men_men_n207_), .C(men_men_n195_), .D(men_men_n181_), .Y(men_men_n224_));
  AOI210     u202(.A0(men_men_n167_), .A1(men_men_n102_), .B0(men_men_n224_), .Y(men_men_n225_));
  AOI210     u203(.A0(men_men_n145_), .A1(x09), .B0(men_men_n73_), .Y(men_men_n226_));
  NA2        u204(.A(men_men_n226_), .B(men_men_n147_), .Y(men_men_n227_));
  NA2        u205(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n228_));
  NA2        u206(.A(men_men_n228_), .B(men_men_n146_), .Y(men_men_n229_));
  AOI210     u207(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n230_));
  NO2        u208(.A(men_men_n134_), .B(x06), .Y(men_men_n231_));
  AOI210     u209(.A0(men_men_n230_), .A1(men_men_n229_), .B0(men_men_n231_), .Y(men_men_n232_));
  AOI210     u210(.A0(men_men_n232_), .A1(men_men_n227_), .B0(x12), .Y(men_men_n233_));
  INV        u211(.A(men_men_n76_), .Y(men_men_n234_));
  AOI210     u212(.A0(men_men_n211_), .A1(x05), .B0(men_men_n51_), .Y(men_men_n235_));
  OAI210     u213(.A0(men_men_n235_), .A1(men_men_n172_), .B0(men_men_n57_), .Y(men_men_n236_));
  NA2        u214(.A(men_men_n236_), .B(men_men_n234_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n96_), .B(x06), .Y(men_men_n238_));
  AOI210     u216(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n239_));
  NO3        u217(.A(men_men_n239_), .B(men_men_n238_), .C(men_men_n41_), .Y(men_men_n240_));
  NA4        u218(.A(men_men_n170_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n241_));
  NA2        u219(.A(men_men_n241_), .B(men_men_n152_), .Y(men_men_n242_));
  OAI210     u220(.A0(men_men_n242_), .A1(men_men_n240_), .B0(x02), .Y(men_men_n243_));
  AOI210     u221(.A0(men_men_n243_), .A1(men_men_n237_), .B0(men_men_n23_), .Y(men_men_n244_));
  OAI210     u222(.A0(men_men_n233_), .A1(men_men_n57_), .B0(men_men_n244_), .Y(men_men_n245_));
  INV        u223(.A(men_men_n152_), .Y(men_men_n246_));
  NO2        u224(.A(men_men_n51_), .B(x03), .Y(men_men_n247_));
  OAI210     u225(.A0(men_men_n79_), .A1(men_men_n36_), .B0(men_men_n125_), .Y(men_men_n248_));
  NO2        u226(.A(men_men_n103_), .B(x03), .Y(men_men_n249_));
  AOI220     u227(.A0(men_men_n249_), .A1(men_men_n248_), .B0(men_men_n76_), .B1(men_men_n247_), .Y(men_men_n250_));
  NA2        u228(.A(men_men_n32_), .B(x06), .Y(men_men_n251_));
  INV        u229(.A(men_men_n170_), .Y(men_men_n252_));
  NOi21      u230(.An(x13), .B(x04), .Y(men_men_n253_));
  NO3        u231(.A(men_men_n253_), .B(men_men_n76_), .C(men_men_n208_), .Y(men_men_n254_));
  NO2        u232(.A(men_men_n254_), .B(x05), .Y(men_men_n255_));
  AOI220     u233(.A0(men_men_n255_), .A1(men_men_n251_), .B0(men_men_n252_), .B1(men_men_n57_), .Y(men_men_n256_));
  OAI210     u234(.A0(men_men_n250_), .A1(men_men_n246_), .B0(men_men_n256_), .Y(men_men_n257_));
  INV        u235(.A(men_men_n92_), .Y(men_men_n258_));
  NA2        u236(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n259_));
  NO2        u237(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n260_));
  OAI210     u238(.A0(men_men_n260_), .A1(men_men_n200_), .B0(men_men_n198_), .Y(men_men_n261_));
  AOI210     u239(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n262_));
  NO2        u240(.A(x06), .B(x00), .Y(men_men_n263_));
  NO3        u241(.A(men_men_n263_), .B(men_men_n262_), .C(men_men_n41_), .Y(men_men_n264_));
  OAI210     u242(.A0(men_men_n106_), .A1(men_men_n158_), .B0(men_men_n72_), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n265_), .B(men_men_n264_), .Y(men_men_n266_));
  NA2        u244(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n267_));
  NA2        u245(.A(men_men_n267_), .B(x03), .Y(men_men_n268_));
  OA210      u246(.A0(men_men_n268_), .A1(men_men_n266_), .B0(men_men_n261_), .Y(men_men_n269_));
  NA2        u247(.A(x13), .B(men_men_n102_), .Y(men_men_n270_));
  NA3        u248(.A(men_men_n270_), .B(men_men_n214_), .C(men_men_n93_), .Y(men_men_n271_));
  OAI210     u249(.A0(men_men_n269_), .A1(men_men_n259_), .B0(men_men_n271_), .Y(men_men_n272_));
  AOI210     u250(.A0(men_men_n92_), .A1(men_men_n257_), .B0(men_men_n272_), .Y(men_men_n273_));
  AOI210     u251(.A0(men_men_n273_), .A1(men_men_n245_), .B0(x07), .Y(men_men_n274_));
  NA2        u252(.A(men_men_n71_), .B(men_men_n29_), .Y(men_men_n275_));
  NOi31      u253(.An(men_men_n145_), .B(men_men_n253_), .C(men_men_n208_), .Y(men_men_n276_));
  AOI210     u254(.A0(men_men_n276_), .A1(men_men_n160_), .B0(men_men_n275_), .Y(men_men_n277_));
  NO2        u255(.A(men_men_n103_), .B(x06), .Y(men_men_n278_));
  INV        u256(.A(men_men_n278_), .Y(men_men_n279_));
  NO2        u257(.A(x08), .B(x05), .Y(men_men_n280_));
  NO2        u258(.A(men_men_n280_), .B(men_men_n262_), .Y(men_men_n281_));
  OAI210     u259(.A0(men_men_n76_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n282_));
  OAI210     u260(.A0(men_men_n281_), .A1(men_men_n279_), .B0(men_men_n282_), .Y(men_men_n283_));
  NO2        u261(.A(x12), .B(x02), .Y(men_men_n284_));
  INV        u262(.A(men_men_n284_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n285_), .B(men_men_n258_), .Y(men_men_n286_));
  OA210      u264(.A0(men_men_n283_), .A1(men_men_n277_), .B0(men_men_n286_), .Y(men_men_n287_));
  NA2        u265(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n288_));
  NO2        u266(.A(men_men_n288_), .B(x01), .Y(men_men_n289_));
  NOi21      u267(.An(men_men_n84_), .B(men_men_n125_), .Y(men_men_n290_));
  NO2        u268(.A(men_men_n290_), .B(men_men_n289_), .Y(men_men_n291_));
  AOI210     u269(.A0(men_men_n291_), .A1(men_men_n139_), .B0(men_men_n29_), .Y(men_men_n292_));
  NA2        u270(.A(men_men_n278_), .B(men_men_n248_), .Y(men_men_n293_));
  NA2        u271(.A(men_men_n103_), .B(x04), .Y(men_men_n294_));
  NA2        u272(.A(men_men_n294_), .B(men_men_n28_), .Y(men_men_n295_));
  OAI210     u273(.A0(men_men_n295_), .A1(men_men_n124_), .B0(men_men_n293_), .Y(men_men_n296_));
  NO3        u274(.A(men_men_n91_), .B(x12), .C(x03), .Y(men_men_n297_));
  OAI210     u275(.A0(men_men_n296_), .A1(men_men_n292_), .B0(men_men_n297_), .Y(men_men_n298_));
  AOI210     u276(.A0(men_men_n219_), .A1(men_men_n213_), .B0(men_men_n106_), .Y(men_men_n299_));
  NOi21      u277(.An(men_men_n275_), .B(men_men_n238_), .Y(men_men_n300_));
  NO2        u278(.A(men_men_n25_), .B(x00), .Y(men_men_n301_));
  OAI210     u279(.A0(men_men_n300_), .A1(men_men_n299_), .B0(men_men_n301_), .Y(men_men_n302_));
  NO2        u280(.A(men_men_n58_), .B(x05), .Y(men_men_n303_));
  NO3        u281(.A(men_men_n303_), .B(men_men_n239_), .C(men_men_n203_), .Y(men_men_n304_));
  NO2        u282(.A(men_men_n259_), .B(men_men_n28_), .Y(men_men_n305_));
  OAI210     u283(.A0(men_men_n304_), .A1(men_men_n246_), .B0(men_men_n305_), .Y(men_men_n306_));
  NA3        u284(.A(men_men_n306_), .B(men_men_n302_), .C(men_men_n298_), .Y(men_men_n307_));
  NO3        u285(.A(men_men_n307_), .B(men_men_n287_), .C(men_men_n274_), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n225_), .A1(men_men_n61_), .B0(men_men_n308_), .Y(men02));
  AOI210     u287(.A0(men_men_n145_), .A1(men_men_n85_), .B0(men_men_n137_), .Y(men_men_n310_));
  NOi21      u288(.An(men_men_n254_), .B(men_men_n186_), .Y(men_men_n311_));
  NO2        u289(.A(men_men_n103_), .B(men_men_n35_), .Y(men_men_n312_));
  NA3        u290(.A(men_men_n312_), .B(men_men_n212_), .C(men_men_n56_), .Y(men_men_n313_));
  OAI210     u291(.A0(men_men_n311_), .A1(men_men_n32_), .B0(men_men_n313_), .Y(men_men_n314_));
  OAI210     u292(.A0(men_men_n314_), .A1(men_men_n310_), .B0(men_men_n183_), .Y(men_men_n315_));
  INV        u293(.A(men_men_n183_), .Y(men_men_n316_));
  AOI210     u294(.A0(men_men_n120_), .A1(men_men_n86_), .B0(men_men_n239_), .Y(men_men_n317_));
  OAI220     u295(.A0(men_men_n317_), .A1(men_men_n103_), .B0(men_men_n85_), .B1(men_men_n51_), .Y(men_men_n318_));
  AOI220     u296(.A0(men_men_n318_), .A1(men_men_n316_), .B0(men_men_n164_), .B1(men_men_n163_), .Y(men_men_n319_));
  AOI210     u297(.A0(men_men_n319_), .A1(men_men_n315_), .B0(men_men_n48_), .Y(men_men_n320_));
  NO2        u298(.A(x05), .B(x02), .Y(men_men_n321_));
  OAI210     u299(.A0(men_men_n229_), .A1(men_men_n208_), .B0(men_men_n321_), .Y(men_men_n322_));
  AOI220     u300(.A0(men_men_n280_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n323_));
  NOi21      u301(.An(men_men_n312_), .B(men_men_n323_), .Y(men_men_n324_));
  AOI210     u302(.A0(men_men_n253_), .A1(men_men_n79_), .B0(men_men_n324_), .Y(men_men_n325_));
  AOI210     u303(.A0(men_men_n325_), .A1(men_men_n322_), .B0(men_men_n152_), .Y(men_men_n326_));
  NAi21      u304(.An(men_men_n255_), .B(men_men_n250_), .Y(men_men_n327_));
  NO2        u305(.A(men_men_n267_), .B(men_men_n47_), .Y(men_men_n328_));
  NA2        u306(.A(men_men_n328_), .B(men_men_n327_), .Y(men_men_n329_));
  AN2        u307(.A(men_men_n249_), .B(men_men_n248_), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n331_));
  NA2        u309(.A(x13), .B(men_men_n28_), .Y(men_men_n332_));
  OA210      u310(.A0(men_men_n332_), .A1(x08), .B0(men_men_n156_), .Y(men_men_n333_));
  AOI210     u311(.A0(men_men_n333_), .A1(men_men_n146_), .B0(men_men_n331_), .Y(men_men_n334_));
  OAI210     u312(.A0(men_men_n334_), .A1(men_men_n330_), .B0(men_men_n97_), .Y(men_men_n335_));
  NA3        u313(.A(men_men_n97_), .B(men_men_n84_), .C(men_men_n247_), .Y(men_men_n336_));
  NA3        u314(.A(men_men_n96_), .B(men_men_n83_), .C(men_men_n42_), .Y(men_men_n337_));
  AOI210     u315(.A0(men_men_n337_), .A1(men_men_n336_), .B0(x04), .Y(men_men_n338_));
  INV        u316(.A(men_men_n163_), .Y(men_men_n339_));
  OAI220     u317(.A0(men_men_n281_), .A1(men_men_n109_), .B0(men_men_n339_), .B1(men_men_n136_), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n340_), .A1(x13), .B0(men_men_n338_), .Y(men_men_n341_));
  NA3        u319(.A(men_men_n341_), .B(men_men_n335_), .C(men_men_n329_), .Y(men_men_n342_));
  NO3        u320(.A(men_men_n342_), .B(men_men_n326_), .C(men_men_n320_), .Y(men_men_n343_));
  NA2        u321(.A(men_men_n151_), .B(x03), .Y(men_men_n344_));
  INV        u322(.A(men_men_n197_), .Y(men_men_n345_));
  OAI210     u323(.A0(men_men_n51_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n346_));
  AOI220     u324(.A0(men_men_n346_), .A1(men_men_n345_), .B0(men_men_n220_), .B1(x08), .Y(men_men_n347_));
  OAI210     u325(.A0(men_men_n347_), .A1(men_men_n303_), .B0(men_men_n344_), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n348_), .B(men_men_n111_), .Y(men_men_n349_));
  NA2        u327(.A(men_men_n182_), .B(men_men_n176_), .Y(men_men_n350_));
  AN2        u328(.A(men_men_n350_), .B(men_men_n189_), .Y(men_men_n351_));
  INV        u329(.A(men_men_n56_), .Y(men_men_n352_));
  OAI220     u330(.A0(men_men_n294_), .A1(men_men_n352_), .B0(men_men_n137_), .B1(men_men_n28_), .Y(men_men_n353_));
  OAI210     u331(.A0(men_men_n353_), .A1(men_men_n351_), .B0(men_men_n112_), .Y(men_men_n354_));
  NA2        u332(.A(men_men_n102_), .B(men_men_n41_), .Y(men_men_n355_));
  NA3        u333(.A(men_men_n354_), .B(men_men_n349_), .C(men_men_n48_), .Y(men_men_n356_));
  INV        u334(.A(men_men_n220_), .Y(men_men_n357_));
  NO2        u335(.A(men_men_n177_), .B(men_men_n40_), .Y(men_men_n358_));
  NA2        u336(.A(men_men_n32_), .B(x05), .Y(men_men_n359_));
  OAI220     u337(.A0(men_men_n359_), .A1(men_men_n358_), .B0(men_men_n357_), .B1(men_men_n59_), .Y(men_men_n360_));
  NA2        u338(.A(men_men_n360_), .B(x02), .Y(men_men_n361_));
  INV        u339(.A(men_men_n260_), .Y(men_men_n362_));
  NA2        u340(.A(men_men_n217_), .B(x04), .Y(men_men_n363_));
  NO2        u341(.A(men_men_n363_), .B(men_men_n362_), .Y(men_men_n364_));
  NO3        u342(.A(men_men_n199_), .B(x13), .C(men_men_n31_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n365_), .A1(men_men_n364_), .B0(men_men_n97_), .Y(men_men_n366_));
  NO3        u344(.A(men_men_n217_), .B(men_men_n175_), .C(men_men_n52_), .Y(men_men_n367_));
  OAI210     u345(.A0(men_men_n158_), .A1(men_men_n36_), .B0(men_men_n102_), .Y(men_men_n368_));
  OAI210     u346(.A0(men_men_n368_), .A1(men_men_n209_), .B0(men_men_n367_), .Y(men_men_n369_));
  NA4        u347(.A(men_men_n369_), .B(men_men_n366_), .C(men_men_n361_), .D(x06), .Y(men_men_n370_));
  NA2        u348(.A(x09), .B(x03), .Y(men_men_n371_));
  OAI220     u349(.A0(men_men_n371_), .A1(men_men_n135_), .B0(men_men_n228_), .B1(men_men_n63_), .Y(men_men_n372_));
  OAI220     u350(.A0(men_men_n176_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n373_));
  NO3        u351(.A(men_men_n303_), .B(men_men_n134_), .C(x08), .Y(men_men_n374_));
  AOI210     u352(.A0(men_men_n373_), .A1(men_men_n246_), .B0(men_men_n374_), .Y(men_men_n375_));
  NO2        u353(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n376_));
  NO3        u354(.A(men_men_n118_), .B(men_men_n135_), .C(men_men_n38_), .Y(men_men_n377_));
  AOI210     u355(.A0(men_men_n367_), .A1(men_men_n376_), .B0(men_men_n377_), .Y(men_men_n378_));
  OAI210     u356(.A0(men_men_n375_), .A1(men_men_n28_), .B0(men_men_n378_), .Y(men_men_n379_));
  AO220      u357(.A0(men_men_n379_), .A1(x04), .B0(men_men_n372_), .B1(x05), .Y(men_men_n380_));
  AOI210     u358(.A0(men_men_n370_), .A1(men_men_n356_), .B0(men_men_n380_), .Y(men_men_n381_));
  OAI210     u359(.A0(men_men_n343_), .A1(x12), .B0(men_men_n381_), .Y(men03));
  OR2        u360(.A(men_men_n42_), .B(men_men_n247_), .Y(men_men_n383_));
  AOI210     u361(.A0(men_men_n164_), .A1(men_men_n102_), .B0(men_men_n383_), .Y(men_men_n384_));
  AO210      u362(.A0(men_men_n362_), .A1(men_men_n86_), .B0(men_men_n363_), .Y(men_men_n385_));
  NA2        u363(.A(men_men_n217_), .B(men_men_n163_), .Y(men_men_n386_));
  NA3        u364(.A(men_men_n386_), .B(men_men_n385_), .C(men_men_n221_), .Y(men_men_n387_));
  OAI210     u365(.A0(men_men_n387_), .A1(men_men_n384_), .B0(x05), .Y(men_men_n388_));
  INV        u366(.A(x05), .Y(men_men_n389_));
  AOI210     u367(.A0(men_men_n146_), .A1(men_men_n234_), .B0(men_men_n389_), .Y(men_men_n390_));
  AOI210     u368(.A0(men_men_n249_), .A1(men_men_n80_), .B0(men_men_n128_), .Y(men_men_n391_));
  OAI220     u369(.A0(men_men_n391_), .A1(men_men_n59_), .B0(men_men_n332_), .B1(men_men_n323_), .Y(men_men_n392_));
  OAI210     u370(.A0(men_men_n392_), .A1(men_men_n390_), .B0(men_men_n102_), .Y(men_men_n393_));
  AOI210     u371(.A0(men_men_n156_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n394_));
  NO2        u372(.A(men_men_n186_), .B(men_men_n141_), .Y(men_men_n395_));
  OAI220     u373(.A0(men_men_n395_), .A1(men_men_n37_), .B0(men_men_n159_), .B1(x13), .Y(men_men_n396_));
  OAI210     u374(.A0(men_men_n396_), .A1(men_men_n394_), .B0(x04), .Y(men_men_n397_));
  NO3        u375(.A(men_men_n355_), .B(men_men_n85_), .C(men_men_n59_), .Y(men_men_n398_));
  AOI210     u376(.A0(men_men_n205_), .A1(men_men_n102_), .B0(men_men_n156_), .Y(men_men_n399_));
  OA210      u377(.A0(men_men_n177_), .A1(x12), .B0(men_men_n141_), .Y(men_men_n400_));
  NO3        u378(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n398_), .Y(men_men_n401_));
  NA4        u379(.A(men_men_n401_), .B(men_men_n397_), .C(men_men_n393_), .D(men_men_n388_), .Y(men04));
  AOI210     u380(.A0(men_men_n71_), .A1(men_men_n52_), .B0(men_men_n231_), .Y(men_men_n403_));
  AOI210     u381(.A0(men_men_n403_), .A1(men_men_n331_), .B0(men_men_n25_), .Y(men_men_n404_));
  NAi41      u382(.An(men_men_n77_), .B(men_men_n152_), .C(men_men_n137_), .D(men_men_n31_), .Y(men_men_n405_));
  AOI210     u383(.A0(men_men_n252_), .A1(men_men_n57_), .B0(men_men_n90_), .Y(men_men_n406_));
  AOI210     u384(.A0(men_men_n406_), .A1(men_men_n405_), .B0(men_men_n24_), .Y(men_men_n407_));
  OAI210     u385(.A0(men_men_n407_), .A1(men_men_n404_), .B0(men_men_n102_), .Y(men_men_n408_));
  NA2        u386(.A(x11), .B(men_men_n31_), .Y(men_men_n409_));
  NA2        u387(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n410_));
  NA2        u388(.A(men_men_n275_), .B(x03), .Y(men_men_n411_));
  OAI220     u389(.A0(men_men_n411_), .A1(men_men_n410_), .B0(men_men_n409_), .B1(men_men_n81_), .Y(men_men_n412_));
  OAI210     u390(.A0(men_men_n26_), .A1(men_men_n102_), .B0(x07), .Y(men_men_n413_));
  AOI210     u391(.A0(men_men_n412_), .A1(x06), .B0(men_men_n413_), .Y(men_men_n414_));
  AOI220     u392(.A0(men_men_n81_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n415_));
  NO3        u393(.A(men_men_n415_), .B(men_men_n23_), .C(x00), .Y(men_men_n416_));
  NA2        u394(.A(men_men_n70_), .B(x02), .Y(men_men_n417_));
  AOI210     u395(.A0(men_men_n417_), .A1(men_men_n411_), .B0(men_men_n278_), .Y(men_men_n418_));
  OR2        u396(.A(men_men_n418_), .B(men_men_n259_), .Y(men_men_n419_));
  NA2        u397(.A(men_men_n171_), .B(x05), .Y(men_men_n420_));
  NA3        u398(.A(men_men_n420_), .B(men_men_n263_), .C(men_men_n258_), .Y(men_men_n421_));
  NO2        u399(.A(men_men_n23_), .B(x10), .Y(men_men_n422_));
  OAI210     u400(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n423_));
  OR3        u401(.A(men_men_n423_), .B(men_men_n422_), .C(men_men_n44_), .Y(men_men_n424_));
  NA3        u402(.A(men_men_n424_), .B(men_men_n421_), .C(men_men_n419_), .Y(men_men_n425_));
  OAI210     u403(.A0(men_men_n425_), .A1(men_men_n416_), .B0(men_men_n102_), .Y(men_men_n426_));
  NA2        u404(.A(men_men_n33_), .B(men_men_n102_), .Y(men_men_n427_));
  AOI210     u405(.A0(men_men_n427_), .A1(men_men_n92_), .B0(x07), .Y(men_men_n428_));
  AOI220     u406(.A0(men_men_n428_), .A1(men_men_n426_), .B0(men_men_n414_), .B1(men_men_n408_), .Y(men_men_n429_));
  NA3        u407(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n430_));
  AO210      u408(.A0(men_men_n430_), .A1(men_men_n288_), .B0(men_men_n285_), .Y(men_men_n431_));
  AOI210     u409(.A0(men_men_n422_), .A1(men_men_n74_), .B0(men_men_n151_), .Y(men_men_n432_));
  OR2        u410(.A(men_men_n432_), .B(x03), .Y(men_men_n433_));
  NA2        u411(.A(men_men_n376_), .B(men_men_n61_), .Y(men_men_n434_));
  NO2        u412(.A(men_men_n434_), .B(x11), .Y(men_men_n435_));
  NO3        u413(.A(men_men_n435_), .B(men_men_n155_), .C(men_men_n28_), .Y(men_men_n436_));
  AOI220     u414(.A0(men_men_n436_), .A1(men_men_n433_), .B0(men_men_n431_), .B1(men_men_n47_), .Y(men_men_n437_));
  NO4        u415(.A(men_men_n355_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n438_));
  OAI210     u416(.A0(men_men_n438_), .A1(men_men_n437_), .B0(men_men_n103_), .Y(men_men_n439_));
  AOI210     u417(.A0(men_men_n363_), .A1(men_men_n114_), .B0(men_men_n284_), .Y(men_men_n440_));
  NOi21      u418(.An(men_men_n344_), .B(men_men_n141_), .Y(men_men_n441_));
  NO2        u419(.A(men_men_n441_), .B(men_men_n285_), .Y(men_men_n442_));
  OAI210     u420(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n443_));
  AOI210     u421(.A0(men_men_n270_), .A1(men_men_n47_), .B0(men_men_n443_), .Y(men_men_n444_));
  NO4        u422(.A(men_men_n444_), .B(men_men_n442_), .C(men_men_n440_), .D(x08), .Y(men_men_n445_));
  AOI210     u423(.A0(men_men_n422_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n446_));
  NA2        u424(.A(x09), .B(men_men_n41_), .Y(men_men_n447_));
  OAI220     u425(.A0(men_men_n447_), .A1(men_men_n446_), .B0(men_men_n409_), .B1(men_men_n66_), .Y(men_men_n448_));
  NO2        u426(.A(x13), .B(x12), .Y(men_men_n449_));
  NO2        u427(.A(men_men_n137_), .B(men_men_n28_), .Y(men_men_n450_));
  NO2        u428(.A(men_men_n450_), .B(men_men_n289_), .Y(men_men_n451_));
  OR3        u429(.A(men_men_n451_), .B(x12), .C(x03), .Y(men_men_n452_));
  NA3        u430(.A(men_men_n357_), .B(men_men_n130_), .C(x12), .Y(men_men_n453_));
  AO210      u431(.A0(men_men_n357_), .A1(men_men_n130_), .B0(men_men_n270_), .Y(men_men_n454_));
  NA4        u432(.A(men_men_n454_), .B(men_men_n453_), .C(men_men_n452_), .D(x08), .Y(men_men_n455_));
  AOI210     u433(.A0(men_men_n449_), .A1(men_men_n448_), .B0(men_men_n455_), .Y(men_men_n456_));
  AOI210     u434(.A0(men_men_n445_), .A1(men_men_n439_), .B0(men_men_n456_), .Y(men_men_n457_));
  OAI210     u435(.A0(men_men_n434_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n458_));
  NA2        u436(.A(men_men_n316_), .B(x07), .Y(men_men_n459_));
  OAI220     u437(.A0(men_men_n459_), .A1(men_men_n410_), .B0(men_men_n155_), .B1(men_men_n43_), .Y(men_men_n460_));
  OAI210     u438(.A0(men_men_n460_), .A1(men_men_n458_), .B0(men_men_n204_), .Y(men_men_n461_));
  INV        u439(.A(x14), .Y(men_men_n462_));
  NO3        u440(.A(men_men_n344_), .B(men_men_n109_), .C(x11), .Y(men_men_n463_));
  NO3        u441(.A(men_men_n176_), .B(men_men_n74_), .C(men_men_n57_), .Y(men_men_n464_));
  NO3        u442(.A(men_men_n430_), .B(men_men_n355_), .C(men_men_n197_), .Y(men_men_n465_));
  NO4        u443(.A(men_men_n465_), .B(men_men_n464_), .C(men_men_n463_), .D(men_men_n462_), .Y(men_men_n466_));
  NA2        u444(.A(men_men_n466_), .B(men_men_n461_), .Y(men_men_n467_));
  AOI220     u445(.A0(men_men_n427_), .A1(men_men_n61_), .B0(men_men_n450_), .B1(men_men_n175_), .Y(men_men_n468_));
  NOi21      u446(.An(men_men_n294_), .B(men_men_n159_), .Y(men_men_n469_));
  NO3        u447(.A(men_men_n134_), .B(men_men_n24_), .C(x06), .Y(men_men_n470_));
  AOI210     u448(.A0(men_men_n301_), .A1(men_men_n252_), .B0(men_men_n470_), .Y(men_men_n471_));
  OAI210     u449(.A0(men_men_n44_), .A1(x04), .B0(men_men_n471_), .Y(men_men_n472_));
  OAI210     u450(.A0(men_men_n472_), .A1(men_men_n469_), .B0(men_men_n102_), .Y(men_men_n473_));
  OAI210     u451(.A0(men_men_n468_), .A1(men_men_n91_), .B0(men_men_n473_), .Y(men_men_n474_));
  NO4        u452(.A(men_men_n474_), .B(men_men_n467_), .C(men_men_n457_), .D(men_men_n429_), .Y(men06));
  INV        u453(.A(x07), .Y(men_men_n478_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule