//Benchmark atmr_alu4_1266_0.5

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n115_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n83_, mai_mai_n84_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n141_, men_men_n142_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1146_, men_men_n1147_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o00(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o01(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o02(.A(i_9_), .Y(ori_ori_n25_));
  INV        o03(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o04(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o05(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o06(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o07(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o08(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o09(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o10(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o11(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o12(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o13(.A(i_4_), .Y(ori_ori_n36_));
  INV        o14(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o15(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o16(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori7));
  INV        o17(.A(ori_ori_n35_), .Y(ori1));
  INV        o18(.A(i_2_), .Y(ori_ori_n41_));
  INV        o19(.A(i_5_), .Y(ori_ori_n42_));
  NO2        o20(.A(i_7_), .B(i_10_), .Y(ori_ori_n43_));
  AOI210     o21(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n43_), .Y(ori_ori_n44_));
  INV        o22(.A(i_5_), .Y(ori_ori_n45_));
  NA2        o23(.A(ori_ori_n45_), .B(i_11_), .Y(ori_ori_n46_));
  INV        o24(.A(i_1_), .Y(ori_ori_n47_));
  NA2        o25(.A(ori_ori_n44_), .B(i_2_), .Y(ori_ori_n48_));
  NA2        o26(.A(i_1_), .B(i_6_), .Y(ori_ori_n49_));
  NO2        o27(.A(ori_ori_n49_), .B(ori_ori_n25_), .Y(ori_ori_n50_));
  INV        o28(.A(i_0_), .Y(ori_ori_n51_));
  NAi21      o29(.An(i_5_), .B(i_10_), .Y(ori_ori_n52_));
  NA2        o30(.A(i_5_), .B(i_9_), .Y(ori_ori_n53_));
  AOI210     o31(.A0(ori_ori_n53_), .A1(ori_ori_n52_), .B0(ori_ori_n51_), .Y(ori_ori_n54_));
  NO2        o32(.A(ori_ori_n54_), .B(ori_ori_n50_), .Y(ori_ori_n55_));
  NA2        o33(.A(i_12_), .B(i_5_), .Y(ori_ori_n56_));
  NA2        o34(.A(i_6_), .B(i_9_), .Y(ori_ori_n57_));
  NA2        o35(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n58_));
  NA2        o36(.A(ori_ori_n58_), .B(i_7_), .Y(ori_ori_n59_));
  NO2        o37(.A(ori_ori_n59_), .B(ori_ori_n41_), .Y(ori_ori_n60_));
  NA3        o38(.A(ori_ori_n56_), .B(ori_ori_n51_), .C(ori_ori_n46_), .Y(ori2));
  NO2        o39(.A(ori_ori_n47_), .B(ori_ori_n37_), .Y(ori_ori_n62_));
  INV        o40(.A(i_6_), .Y(ori_ori_n63_));
  NA2        o41(.A(ori_ori_n63_), .B(ori_ori_n62_), .Y(ori_ori_n64_));
  NA4        o42(.A(ori_ori_n64_), .B(ori_ori_n55_), .C(ori_ori_n48_), .D(ori_ori_n30_), .Y(ori0));
  INV        o43(.A(i_5_), .Y(ori_ori_n66_));
  INV        o44(.A(i_12_), .Y(ori_ori_n67_));
  INV        o45(.A(i_0_), .Y(ori_ori_n68_));
  NOi21      o46(.An(i_5_), .B(i_0_), .Y(ori_ori_n69_));
  NO2        o47(.A(i_0_), .B(i_11_), .Y(ori_ori_n70_));
  NO2        o48(.A(i_10_), .B(i_9_), .Y(ori_ori_n71_));
  NO2        o49(.A(ori_ori_n37_), .B(i_6_), .Y(ori_ori_n72_));
  INV        o50(.A(ori_ori_n72_), .Y(ori_ori_n73_));
  NO2        o51(.A(ori_ori_n73_), .B(ori_ori_n47_), .Y(ori_ori_n74_));
  NOi21      o52(.An(i_11_), .B(i_7_), .Y(ori_ori_n75_));
  AO210      o53(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n76_));
  NO2        o54(.A(ori_ori_n76_), .B(ori_ori_n75_), .Y(ori_ori_n77_));
  NA2        o55(.A(ori_ori_n115_), .B(ori_ori_n47_), .Y(ori_ori_n78_));
  INV        o56(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NA2        o57(.A(ori_ori_n79_), .B(i_6_), .Y(ori_ori_n80_));
  NO2        o58(.A(i_6_), .B(i_11_), .Y(ori_ori_n81_));
  INV        o59(.A(ori_ori_n80_), .Y(ori_ori_n82_));
  INV        o60(.A(i_1_), .Y(ori_ori_n83_));
  NO2        o61(.A(ori_ori_n57_), .B(ori_ori_n83_), .Y(ori_ori_n84_));
  INV        o62(.A(ori_ori_n84_), .Y(ori_ori_n85_));
  NA2        o63(.A(ori_ori_n81_), .B(ori_ori_n47_), .Y(ori_ori_n86_));
  NA2        o64(.A(ori_ori_n86_), .B(ori_ori_n85_), .Y(ori_ori_n87_));
  OR3        o65(.A(ori_ori_n87_), .B(ori_ori_n82_), .C(ori_ori_n74_), .Y(ori5));
  INV        o66(.A(ori_ori_n71_), .Y(ori_ori_n89_));
  OA210      o67(.A0(ori_ori_n77_), .A1(ori_ori_n60_), .B0(i_13_), .Y(ori_ori_n90_));
  INV        o68(.A(i_2_), .Y(ori_ori_n91_));
  NA2        o69(.A(i_10_), .B(ori_ori_n58_), .Y(ori_ori_n92_));
  NO2        o70(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  NO2        o71(.A(ori_ori_n93_), .B(ori_ori_n90_), .Y(ori_ori_n94_));
  INV        o72(.A(ori_ori_n69_), .Y(ori_ori_n95_));
  OR2        o73(.A(ori_ori_n95_), .B(i_12_), .Y(ori_ori_n96_));
  OR2        o74(.A(ori_ori_n89_), .B(ori_ori_n36_), .Y(ori_ori_n97_));
  INV        o75(.A(ori_ori_n97_), .Y(ori_ori_n98_));
  NA2        o76(.A(ori_ori_n56_), .B(ori_ori_n70_), .Y(ori_ori_n99_));
  INV        o77(.A(ori_ori_n99_), .Y(ori_ori_n100_));
  NO2        o78(.A(ori_ori_n100_), .B(ori_ori_n98_), .Y(ori_ori_n101_));
  NA2        o79(.A(ori_ori_n101_), .B(ori_ori_n96_), .Y(ori3));
  NA2        o80(.A(i_9_), .B(i_0_), .Y(ori_ori_n103_));
  NA2        o81(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n104_));
  AOI210     o82(.A0(ori_ori_n104_), .A1(ori_ori_n103_), .B0(ori_ori_n66_), .Y(ori_ori_n105_));
  NO3        o83(.A(i_11_), .B(i_5_), .C(i_0_), .Y(ori_ori_n106_));
  NO2        o84(.A(ori_ori_n106_), .B(ori_ori_n105_), .Y(ori_ori_n107_));
  NA2        o85(.A(i_10_), .B(ori_ori_n42_), .Y(ori_ori_n108_));
  NO2        o86(.A(ori_ori_n108_), .B(ori_ori_n51_), .Y(ori_ori_n109_));
  INV        o87(.A(ori_ori_n109_), .Y(ori_ori_n110_));
  NA2        o88(.A(ori_ori_n110_), .B(ori_ori_n107_), .Y(ori4));
  INV        o89(.A(ori_ori_n94_), .Y(ori6));
  INV        o90(.A(i_12_), .Y(ori_ori_n115_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NOi21      m016(.An(i_12_), .B(i_13_), .Y(mai_mai_n39_));
  INV        m017(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NAi31      m018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n41_));
  INV        m019(.A(mai_mai_n35_), .Y(mai1));
  INV        m020(.A(i_11_), .Y(mai_mai_n43_));
  NO2        m021(.A(mai_mai_n43_), .B(i_6_), .Y(mai_mai_n44_));
  INV        m022(.A(i_2_), .Y(mai_mai_n45_));
  INV        m023(.A(i_5_), .Y(mai_mai_n46_));
  NO2        m024(.A(i_7_), .B(i_10_), .Y(mai_mai_n47_));
  AOI210     m025(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n47_), .Y(mai_mai_n48_));
  INV        m026(.A(i_1_), .Y(mai_mai_n49_));
  NA2        m027(.A(mai_mai_n48_), .B(i_2_), .Y(mai_mai_n50_));
  AOI210     m028(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_1_), .B(i_6_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(mai_mai_n25_), .Y(mai_mai_n53_));
  INV        m031(.A(i_0_), .Y(mai_mai_n54_));
  NAi21      m032(.An(i_5_), .B(i_10_), .Y(mai_mai_n55_));
  NA2        m033(.A(i_5_), .B(i_9_), .Y(mai_mai_n56_));
  AOI210     m034(.A0(mai_mai_n56_), .A1(mai_mai_n55_), .B0(mai_mai_n54_), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n58_));
  NA2        m036(.A(i_12_), .B(i_5_), .Y(mai_mai_n59_));
  NO2        m037(.A(i_3_), .B(i_9_), .Y(mai_mai_n60_));
  INV        m038(.A(i_6_), .Y(mai_mai_n61_));
  INV        m039(.A(i_11_), .Y(mai_mai_n62_));
  NO2        m040(.A(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  NAi21      m041(.An(i_6_), .B(i_10_), .Y(mai_mai_n64_));
  NA2        m042(.A(i_6_), .B(i_9_), .Y(mai_mai_n65_));
  AN3        m043(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n66_));
  NAi21      m044(.An(i_6_), .B(i_11_), .Y(mai_mai_n67_));
  NA2        m045(.A(mai_mai_n66_), .B(mai_mai_n32_), .Y(mai_mai_n68_));
  INV        m046(.A(i_7_), .Y(mai_mai_n69_));
  NO2        m047(.A(i_0_), .B(i_5_), .Y(mai_mai_n70_));
  NO2        m048(.A(i_2_), .B(i_7_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_12_), .B(i_7_), .Y(mai_mai_n72_));
  NO2        m050(.A(mai_mai_n49_), .B(mai_mai_n26_), .Y(mai_mai_n73_));
  NA2        m051(.A(i_11_), .B(i_12_), .Y(mai_mai_n74_));
  NA2        m052(.A(mai_mai_n74_), .B(mai_mai_n68_), .Y(mai_mai_n75_));
  NA2        m053(.A(mai_mai_n69_), .B(mai_mai_n37_), .Y(mai_mai_n76_));
  NA2        m054(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n77_));
  NA2        m055(.A(mai_mai_n77_), .B(mai_mai_n76_), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n78_), .B(mai_mai_n45_), .Y(mai_mai_n79_));
  NA2        m057(.A(mai_mai_n65_), .B(mai_mai_n64_), .Y(mai_mai_n80_));
  INV        m058(.A(mai_mai_n75_), .Y(mai_mai_n81_));
  NA2        m059(.A(mai_mai_n81_), .B(mai_mai_n436_), .Y(mai2));
  NO2        m060(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n83_));
  NA2        m061(.A(mai_mai_n432_), .B(mai_mai_n83_), .Y(mai_mai_n84_));
  NA4        m062(.A(mai_mai_n84_), .B(mai_mai_n58_), .C(mai_mai_n50_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m063(.A(i_8_), .B(i_7_), .Y(mai_mai_n86_));
  NO2        m064(.A(i_12_), .B(i_13_), .Y(mai_mai_n87_));
  NAi21      m065(.An(i_5_), .B(i_11_), .Y(mai_mai_n88_));
  NOi21      m066(.An(mai_mai_n87_), .B(mai_mai_n88_), .Y(mai_mai_n89_));
  NO2        m067(.A(i_0_), .B(i_1_), .Y(mai_mai_n90_));
  NA2        m068(.A(i_2_), .B(i_3_), .Y(mai_mai_n91_));
  NO2        m069(.A(mai_mai_n91_), .B(i_4_), .Y(mai_mai_n92_));
  AN2        m070(.A(mai_mai_n87_), .B(mai_mai_n60_), .Y(mai_mai_n93_));
  OR2        m071(.A(i_0_), .B(i_1_), .Y(mai_mai_n94_));
  NO3        m072(.A(mai_mai_n94_), .B(mai_mai_n59_), .C(i_13_), .Y(mai_mai_n95_));
  NAi32      m073(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n96_));
  NAi21      m074(.An(mai_mai_n96_), .B(mai_mai_n95_), .Y(mai_mai_n97_));
  NOi21      m075(.An(i_4_), .B(i_10_), .Y(mai_mai_n98_));
  NA2        m076(.A(mai_mai_n98_), .B(mai_mai_n39_), .Y(mai_mai_n99_));
  NOi21      m077(.An(i_11_), .B(i_13_), .Y(mai_mai_n100_));
  NA2        m078(.A(mai_mai_n100_), .B(i_4_), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n54_), .B(mai_mai_n49_), .Y(mai_mai_n102_));
  NA2        m080(.A(i_3_), .B(i_5_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n54_), .B(i_5_), .Y(mai_mai_n104_));
  NO2        m082(.A(i_13_), .B(i_10_), .Y(mai_mai_n105_));
  NA3        m083(.A(mai_mai_n105_), .B(mai_mai_n104_), .C(mai_mai_n43_), .Y(mai_mai_n106_));
  NAi21      m084(.An(i_4_), .B(i_12_), .Y(mai_mai_n107_));
  INV        m085(.A(i_8_), .Y(mai_mai_n108_));
  NO3        m086(.A(i_3_), .B(mai_mai_n61_), .C(mai_mai_n46_), .Y(mai_mai_n109_));
  INV        m087(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NO2        m088(.A(i_0_), .B(i_1_), .Y(mai_mai_n111_));
  NA3        m089(.A(mai_mai_n111_), .B(mai_mai_n39_), .C(mai_mai_n43_), .Y(mai_mai_n112_));
  NO3        m090(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n113_));
  NA2        m091(.A(i_12_), .B(mai_mai_n113_), .Y(mai_mai_n114_));
  AOI210     m092(.A0(mai_mai_n114_), .A1(mai_mai_n112_), .B0(mai_mai_n110_), .Y(mai_mai_n115_));
  NO3        m093(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n116_));
  NO2        m094(.A(i_13_), .B(i_9_), .Y(mai_mai_n117_));
  NAi21      m095(.An(i_12_), .B(i_3_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n43_), .B(i_5_), .Y(mai_mai_n119_));
  NA3        m097(.A(i_13_), .B(mai_mai_n108_), .C(i_10_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n120_), .B(i_12_), .Y(mai_mai_n121_));
  NA2        m099(.A(i_0_), .B(i_5_), .Y(mai_mai_n122_));
  NAi31      m100(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n123_));
  NO2        m101(.A(mai_mai_n45_), .B(mai_mai_n49_), .Y(mai_mai_n124_));
  INV        m102(.A(i_13_), .Y(mai_mai_n125_));
  NO2        m103(.A(i_12_), .B(mai_mai_n125_), .Y(mai_mai_n126_));
  NA3        m104(.A(mai_mai_n126_), .B(mai_mai_n111_), .C(mai_mai_n109_), .Y(mai_mai_n127_));
  INV        m105(.A(mai_mai_n127_), .Y(mai_mai_n128_));
  AOI220     m106(.A0(mai_mai_n128_), .A1(mai_mai_n86_), .B0(i_3_), .B1(mai_mai_n121_), .Y(mai_mai_n129_));
  INV        m107(.A(i_12_), .Y(mai_mai_n130_));
  NO3        m108(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n131_));
  NA2        m109(.A(i_2_), .B(i_1_), .Y(mai_mai_n132_));
  NO3        m110(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n133_));
  NAi21      m111(.An(i_4_), .B(i_3_), .Y(mai_mai_n134_));
  NOi41      m112(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n135_));
  NO2        m113(.A(i_11_), .B(mai_mai_n125_), .Y(mai_mai_n136_));
  NO2        m114(.A(i_12_), .B(i_3_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n130_), .B(i_13_), .Y(mai_mai_n138_));
  NO2        m116(.A(mai_mai_n138_), .B(mai_mai_n56_), .Y(mai_mai_n139_));
  NA2        m117(.A(mai_mai_n139_), .B(mai_mai_n86_), .Y(mai_mai_n140_));
  NO2        m118(.A(i_8_), .B(mai_mai_n37_), .Y(mai_mai_n141_));
  NA2        m119(.A(i_12_), .B(i_6_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n134_), .B(i_2_), .Y(mai_mai_n143_));
  NA3        m121(.A(mai_mai_n143_), .B(mai_mai_n434_), .C(mai_mai_n43_), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n136_), .B(i_9_), .Y(mai_mai_n145_));
  INV        m123(.A(mai_mai_n144_), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n146_), .B(mai_mai_n141_), .Y(mai_mai_n147_));
  NA3        m125(.A(mai_mai_n147_), .B(mai_mai_n140_), .C(mai_mai_n129_), .Y(mai_mai_n148_));
  NO3        m126(.A(i_12_), .B(mai_mai_n125_), .C(mai_mai_n37_), .Y(mai_mai_n149_));
  INV        m127(.A(mai_mai_n149_), .Y(mai_mai_n150_));
  NO2        m128(.A(i_3_), .B(i_10_), .Y(mai_mai_n151_));
  NA3        m129(.A(mai_mai_n151_), .B(mai_mai_n39_), .C(mai_mai_n43_), .Y(mai_mai_n152_));
  AN2        m130(.A(i_3_), .B(i_10_), .Y(mai_mai_n153_));
  NO2        m131(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n154_));
  OAI220     m132(.A0(mai_mai_n152_), .A1(i_6_), .B0(mai_mai_n442_), .B1(mai_mai_n150_), .Y(mai_mai_n155_));
  NO3        m133(.A(mai_mai_n155_), .B(mai_mai_n148_), .C(mai_mai_n115_), .Y(mai_mai_n156_));
  NO3        m134(.A(mai_mai_n43_), .B(i_13_), .C(i_9_), .Y(mai_mai_n157_));
  NOi21      m135(.An(i_5_), .B(i_0_), .Y(mai_mai_n158_));
  INV        m136(.A(mai_mai_n99_), .Y(mai_mai_n159_));
  AOI210     m137(.A0(i_4_), .A1(mai_mai_n157_), .B0(mai_mai_n159_), .Y(mai_mai_n160_));
  NOi32      m138(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n161_));
  INV        m139(.A(mai_mai_n161_), .Y(mai_mai_n162_));
  NO2        m140(.A(i_9_), .B(mai_mai_n96_), .Y(mai_mai_n163_));
  NO2        m141(.A(mai_mai_n96_), .B(mai_mai_n94_), .Y(mai_mai_n164_));
  NOi32      m142(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n45_), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n166_), .B(i_0_), .Y(mai_mai_n167_));
  OR2        m145(.A(mai_mai_n167_), .B(mai_mai_n164_), .Y(mai_mai_n168_));
  NAi21      m146(.An(i_3_), .B(i_4_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n169_), .B(i_9_), .Y(mai_mai_n170_));
  NA2        m148(.A(i_7_), .B(mai_mai_n170_), .Y(mai_mai_n171_));
  NA2        m149(.A(i_2_), .B(i_7_), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n169_), .B(i_10_), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n171_), .B(mai_mai_n104_), .Y(mai_mai_n174_));
  INV        m152(.A(mai_mai_n173_), .Y(mai_mai_n175_));
  NO2        m153(.A(mai_mai_n175_), .B(i_5_), .Y(mai_mai_n176_));
  NO4        m154(.A(mai_mai_n176_), .B(mai_mai_n174_), .C(mai_mai_n168_), .D(mai_mai_n163_), .Y(mai_mai_n177_));
  NO2        m155(.A(mai_mai_n177_), .B(mai_mai_n162_), .Y(mai_mai_n178_));
  AN2        m156(.A(i_12_), .B(i_5_), .Y(mai_mai_n179_));
  NA2        m157(.A(i_3_), .B(mai_mai_n179_), .Y(mai_mai_n180_));
  NO2        m158(.A(i_11_), .B(i_6_), .Y(mai_mai_n181_));
  NA3        m159(.A(mai_mai_n181_), .B(i_2_), .C(mai_mai_n125_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n182_), .B(mai_mai_n180_), .Y(mai_mai_n183_));
  NO2        m161(.A(i_5_), .B(i_10_), .Y(mai_mai_n184_));
  INV        m162(.A(mai_mai_n183_), .Y(mai_mai_n185_));
  NO2        m163(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n186_));
  NO3        m164(.A(mai_mai_n61_), .B(mai_mai_n46_), .C(i_9_), .Y(mai_mai_n187_));
  INV        m165(.A(mai_mai_n123_), .Y(mai_mai_n188_));
  NAi21      m166(.An(i_13_), .B(i_0_), .Y(mai_mai_n189_));
  NO2        m167(.A(mai_mai_n189_), .B(mai_mai_n132_), .Y(mai_mai_n190_));
  NA2        m168(.A(mai_mai_n188_), .B(mai_mai_n190_), .Y(mai_mai_n191_));
  NA2        m169(.A(mai_mai_n191_), .B(mai_mai_n185_), .Y(mai_mai_n192_));
  NA2        m170(.A(mai_mai_n43_), .B(mai_mai_n125_), .Y(mai_mai_n193_));
  NO2        m171(.A(i_0_), .B(i_11_), .Y(mai_mai_n194_));
  AN2        m172(.A(i_1_), .B(i_6_), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n86_), .B(i_9_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n196_), .B(i_4_), .Y(mai_mai_n197_));
  OR2        m175(.A(i_13_), .B(i_10_), .Y(mai_mai_n198_));
  NO2        m176(.A(mai_mai_n69_), .B(mai_mai_n25_), .Y(mai_mai_n199_));
  INV        m177(.A(mai_mai_n145_), .Y(mai_mai_n200_));
  NO3        m178(.A(mai_mai_n200_), .B(mai_mai_n192_), .C(mai_mai_n178_), .Y(mai_mai_n201_));
  NO2        m179(.A(mai_mai_n54_), .B(i_13_), .Y(mai_mai_n202_));
  NO2        m180(.A(i_10_), .B(i_9_), .Y(mai_mai_n203_));
  NO2        m181(.A(i_12_), .B(i_3_), .Y(mai_mai_n204_));
  NA2        m182(.A(i_8_), .B(i_9_), .Y(mai_mai_n205_));
  INV        m183(.A(mai_mai_n149_), .Y(mai_mai_n206_));
  NO2        m184(.A(mai_mai_n206_), .B(mai_mai_n205_), .Y(mai_mai_n207_));
  NA2        m185(.A(mai_mai_n136_), .B(mai_mai_n154_), .Y(mai_mai_n208_));
  NO3        m186(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n209_));
  INV        m187(.A(mai_mai_n209_), .Y(mai_mai_n210_));
  NA3        m188(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n211_));
  NA3        m189(.A(mai_mai_n88_), .B(mai_mai_n73_), .C(mai_mai_n23_), .Y(mai_mai_n212_));
  OAI220     m190(.A0(mai_mai_n212_), .A1(mai_mai_n211_), .B0(mai_mai_n210_), .B1(mai_mai_n208_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n213_), .B(mai_mai_n207_), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n66_), .B(i_13_), .Y(mai_mai_n215_));
  NA2        m193(.A(i_3_), .B(i_9_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n217_));
  NO2        m195(.A(i_11_), .B(i_1_), .Y(mai_mai_n218_));
  NA2        m196(.A(i_2_), .B(i_0_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n198_), .B(i_6_), .Y(mai_mai_n220_));
  NA2        m198(.A(mai_mai_n220_), .B(i_1_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n221_), .B(mai_mai_n219_), .Y(mai_mai_n222_));
  NO2        m200(.A(i_6_), .B(i_10_), .Y(mai_mai_n223_));
  NA2        m201(.A(mai_mai_n135_), .B(mai_mai_n100_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n94_), .B(i_3_), .Y(mai_mai_n225_));
  NAi31      m203(.An(i_11_), .B(mai_mai_n225_), .C(mai_mai_n126_), .Y(mai_mai_n226_));
  NA3        m204(.A(mai_mai_n186_), .B(mai_mai_n102_), .C(mai_mai_n92_), .Y(mai_mai_n227_));
  NA3        m205(.A(mai_mai_n227_), .B(mai_mai_n226_), .C(mai_mai_n224_), .Y(mai_mai_n228_));
  NO3        m206(.A(mai_mai_n228_), .B(mai_mai_n222_), .C(mai_mai_n217_), .Y(mai_mai_n229_));
  NA2        m207(.A(mai_mai_n229_), .B(mai_mai_n214_), .Y(mai_mai_n230_));
  INV        m208(.A(mai_mai_n157_), .Y(mai_mai_n231_));
  NO2        m209(.A(mai_mai_n231_), .B(i_12_), .Y(mai_mai_n232_));
  INV        m210(.A(mai_mai_n232_), .Y(mai_mai_n233_));
  NA3        m211(.A(mai_mai_n202_), .B(i_1_), .C(i_2_), .Y(mai_mai_n234_));
  INV        m212(.A(mai_mai_n234_), .Y(mai_mai_n235_));
  NA2        m213(.A(mai_mai_n179_), .B(mai_mai_n125_), .Y(mai_mai_n236_));
  NA2        m214(.A(i_7_), .B(mai_mai_n165_), .Y(mai_mai_n237_));
  OR2        m215(.A(mai_mai_n236_), .B(mai_mai_n237_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n239_));
  INV        m217(.A(mai_mai_n238_), .Y(mai_mai_n240_));
  AOI210     m218(.A0(mai_mai_n235_), .A1(mai_mai_n116_), .B0(mai_mai_n240_), .Y(mai_mai_n241_));
  NO2        m219(.A(i_7_), .B(mai_mai_n112_), .Y(mai_mai_n242_));
  NA2        m220(.A(i_5_), .B(mai_mai_n242_), .Y(mai_mai_n243_));
  NA3        m221(.A(mai_mai_n243_), .B(mai_mai_n241_), .C(mai_mai_n233_), .Y(mai_mai_n244_));
  NOi31      m222(.An(i_8_), .B(mai_mai_n198_), .C(mai_mai_n38_), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n245_), .B(mai_mai_n437_), .Y(mai_mai_n246_));
  NO2        m224(.A(i_8_), .B(i_7_), .Y(mai_mai_n247_));
  INV        m225(.A(mai_mai_n124_), .Y(mai_mai_n248_));
  OAI220     m226(.A0(i_9_), .A1(mai_mai_n103_), .B0(mai_mai_n248_), .B1(mai_mai_n134_), .Y(mai_mai_n249_));
  NA3        m227(.A(i_10_), .B(mai_mai_n249_), .C(mai_mai_n247_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n215_), .B(i_6_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n251_), .B(mai_mai_n141_), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n94_), .B(i_5_), .Y(mai_mai_n253_));
  NA2        m231(.A(mai_mai_n253_), .B(mai_mai_n193_), .Y(mai_mai_n254_));
  INV        m232(.A(mai_mai_n254_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n255_), .B(mai_mai_n209_), .Y(mai_mai_n256_));
  NA4        m234(.A(mai_mai_n256_), .B(mai_mai_n252_), .C(mai_mai_n250_), .D(mai_mai_n246_), .Y(mai_mai_n257_));
  NO3        m235(.A(mai_mai_n41_), .B(i_2_), .C(mai_mai_n46_), .Y(mai_mai_n258_));
  NO3        m236(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n259_));
  AN4        m237(.A(mai_mai_n435_), .B(mai_mai_n197_), .C(i_3_), .D(i_2_), .Y(mai_mai_n260_));
  INV        m238(.A(mai_mai_n260_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n72_), .B(mai_mai_n23_), .Y(mai_mai_n262_));
  NOi21      m240(.An(mai_mai_n89_), .B(i_4_), .Y(mai_mai_n263_));
  NA3        m241(.A(mai_mai_n152_), .B(mai_mai_n438_), .C(mai_mai_n261_), .Y(mai_mai_n264_));
  NO4        m242(.A(mai_mai_n264_), .B(mai_mai_n257_), .C(mai_mai_n244_), .D(mai_mai_n230_), .Y(mai_mai_n265_));
  NA4        m243(.A(mai_mai_n265_), .B(mai_mai_n201_), .C(mai_mai_n160_), .D(mai_mai_n156_), .Y(mai7));
  NA2        m244(.A(i_11_), .B(mai_mai_n108_), .Y(mai_mai_n267_));
  NA2        m245(.A(i_12_), .B(i_8_), .Y(mai_mai_n268_));
  INV        m246(.A(mai_mai_n116_), .Y(mai_mai_n269_));
  OR3        m247(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n270_));
  INV        m248(.A(mai_mai_n113_), .Y(mai_mai_n271_));
  NO2        m249(.A(mai_mai_n270_), .B(mai_mai_n49_), .Y(mai_mai_n272_));
  NOi21      m250(.An(i_11_), .B(i_7_), .Y(mai_mai_n273_));
  AO210      m251(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n274_), .B(mai_mai_n273_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n62_), .B(mai_mai_n49_), .Y(mai_mai_n276_));
  OR2        m254(.A(mai_mai_n276_), .B(mai_mai_n40_), .Y(mai_mai_n277_));
  NA2        m255(.A(mai_mai_n126_), .B(mai_mai_n49_), .Y(mai_mai_n278_));
  NO2        m256(.A(mai_mai_n49_), .B(i_9_), .Y(mai_mai_n279_));
  NO2        m257(.A(i_1_), .B(i_12_), .Y(mai_mai_n280_));
  NA2        m258(.A(mai_mai_n278_), .B(mai_mai_n277_), .Y(mai_mai_n281_));
  NA2        m259(.A(mai_mai_n281_), .B(i_6_), .Y(mai_mai_n282_));
  NO2        m260(.A(i_6_), .B(i_11_), .Y(mai_mai_n283_));
  NO3        m261(.A(i_12_), .B(i_13_), .C(mai_mai_n61_), .Y(mai_mai_n284_));
  NA2        m262(.A(mai_mai_n284_), .B(mai_mai_n279_), .Y(mai_mai_n285_));
  INV        m263(.A(mai_mai_n285_), .Y(mai_mai_n286_));
  INV        m264(.A(i_2_), .Y(mai_mai_n287_));
  NA2        m265(.A(mai_mai_n83_), .B(i_9_), .Y(mai_mai_n288_));
  NO2        m266(.A(mai_mai_n288_), .B(mai_mai_n287_), .Y(mai_mai_n289_));
  NA2        m267(.A(mai_mai_n279_), .B(i_6_), .Y(mai_mai_n290_));
  NO2        m268(.A(mai_mai_n290_), .B(mai_mai_n23_), .Y(mai_mai_n291_));
  AOI210     m269(.A0(mai_mai_n218_), .A1(mai_mai_n199_), .B0(mai_mai_n133_), .Y(mai_mai_n292_));
  NO2        m270(.A(mai_mai_n292_), .B(mai_mai_n440_), .Y(mai_mai_n293_));
  NO2        m271(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n294_));
  OR3        m272(.A(mai_mai_n293_), .B(mai_mai_n291_), .C(mai_mai_n289_), .Y(mai_mai_n295_));
  NO2        m273(.A(mai_mai_n295_), .B(mai_mai_n286_), .Y(mai_mai_n296_));
  NO2        m274(.A(mai_mai_n130_), .B(mai_mai_n69_), .Y(mai_mai_n297_));
  NO2        m275(.A(mai_mai_n297_), .B(mai_mai_n273_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n296_), .B(mai_mai_n282_), .Y(mai_mai_n299_));
  AOI210     m277(.A0(mai_mai_n142_), .A1(mai_mai_n67_), .B0(i_1_), .Y(mai_mai_n300_));
  NA2        m278(.A(i_4_), .B(mai_mai_n300_), .Y(mai_mai_n301_));
  NO2        m279(.A(mai_mai_n301_), .B(i_13_), .Y(mai_mai_n302_));
  NA2        m280(.A(mai_mai_n80_), .B(i_13_), .Y(mai_mai_n303_));
  NO2        m281(.A(mai_mai_n303_), .B(mai_mai_n300_), .Y(mai_mai_n304_));
  NO2        m282(.A(mai_mai_n130_), .B(mai_mai_n61_), .Y(mai_mai_n305_));
  NO2        m283(.A(mai_mai_n431_), .B(mai_mai_n271_), .Y(mai_mai_n306_));
  NO2        m284(.A(mai_mai_n306_), .B(mai_mai_n304_), .Y(mai_mai_n307_));
  NA2        m285(.A(mai_mai_n283_), .B(i_13_), .Y(mai_mai_n308_));
  INV        m286(.A(mai_mai_n308_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n309_), .B(mai_mai_n49_), .Y(mai_mai_n310_));
  NO2        m288(.A(i_2_), .B(i_12_), .Y(mai_mai_n311_));
  NA3        m289(.A(mai_mai_n280_), .B(mai_mai_n44_), .C(mai_mai_n125_), .Y(mai_mai_n312_));
  NA3        m290(.A(mai_mai_n312_), .B(mai_mai_n310_), .C(mai_mai_n307_), .Y(mai_mai_n313_));
  OR4        m291(.A(mai_mai_n313_), .B(mai_mai_n302_), .C(mai_mai_n299_), .D(mai_mai_n272_), .Y(mai5));
  NA2        m292(.A(mai_mai_n298_), .B(mai_mai_n143_), .Y(mai_mai_n315_));
  AN2        m293(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n316_), .B(mai_mai_n311_), .Y(mai_mai_n317_));
  NO2        m295(.A(mai_mai_n268_), .B(i_11_), .Y(mai_mai_n318_));
  NA2        m296(.A(mai_mai_n63_), .B(mai_mai_n318_), .Y(mai_mai_n319_));
  NA3        m297(.A(mai_mai_n319_), .B(mai_mai_n317_), .C(mai_mai_n315_), .Y(mai_mai_n320_));
  NO3        m298(.A(i_11_), .B(mai_mai_n130_), .C(i_13_), .Y(mai_mai_n321_));
  NO2        m299(.A(mai_mai_n77_), .B(mai_mai_n23_), .Y(mai_mai_n322_));
  INV        m300(.A(mai_mai_n203_), .Y(mai_mai_n323_));
  NA2        m301(.A(i_12_), .B(mai_mai_n322_), .Y(mai_mai_n324_));
  INV        m302(.A(mai_mai_n324_), .Y(mai_mai_n325_));
  NO2        m303(.A(mai_mai_n325_), .B(mai_mai_n320_), .Y(mai_mai_n326_));
  INV        m304(.A(mai_mai_n100_), .Y(mai_mai_n327_));
  OAI210     m305(.A0(i_4_), .A1(mai_mai_n204_), .B0(mai_mai_n71_), .Y(mai_mai_n328_));
  NO2        m306(.A(mai_mai_n328_), .B(mai_mai_n327_), .Y(mai_mai_n329_));
  AOI210     m307(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n198_), .Y(mai_mai_n330_));
  AOI210     m308(.A0(mai_mai_n330_), .A1(i_2_), .B0(mai_mai_n329_), .Y(mai_mai_n331_));
  NO2        m309(.A(mai_mai_n107_), .B(mai_mai_n78_), .Y(mai_mai_n332_));
  OAI210     m310(.A0(mai_mai_n332_), .A1(mai_mai_n322_), .B0(i_2_), .Y(mai_mai_n333_));
  NO3        m311(.A(mai_mai_n274_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n334_));
  INV        m312(.A(mai_mai_n334_), .Y(mai_mai_n335_));
  AOI210     m313(.A0(mai_mai_n335_), .A1(mai_mai_n333_), .B0(mai_mai_n108_), .Y(mai_mai_n336_));
  OA210      m314(.A0(mai_mai_n275_), .A1(mai_mai_n79_), .B0(i_13_), .Y(mai_mai_n337_));
  INV        m315(.A(mai_mai_n113_), .Y(mai_mai_n338_));
  INV        m316(.A(mai_mai_n93_), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(mai_mai_n172_), .Y(mai_mai_n340_));
  AOI210     m318(.A0(mai_mai_n118_), .A1(mai_mai_n91_), .B0(mai_mai_n239_), .Y(mai_mai_n341_));
  NA2        m319(.A(mai_mai_n341_), .B(mai_mai_n199_), .Y(mai_mai_n342_));
  NO2        m320(.A(i_2_), .B(mai_mai_n43_), .Y(mai_mai_n343_));
  NA3        m321(.A(mai_mai_n153_), .B(mai_mai_n77_), .C(mai_mai_n41_), .Y(mai_mai_n344_));
  OAI210     m322(.A0(mai_mai_n344_), .A1(mai_mai_n343_), .B0(mai_mai_n342_), .Y(mai_mai_n345_));
  NO4        m323(.A(mai_mai_n345_), .B(mai_mai_n340_), .C(mai_mai_n337_), .D(mai_mai_n336_), .Y(mai_mai_n346_));
  INV        m324(.A(mai_mai_n262_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n321_), .B(i_7_), .Y(mai_mai_n348_));
  NA2        m326(.A(mai_mai_n348_), .B(mai_mai_n347_), .Y(mai_mai_n349_));
  NO2        m327(.A(i_2_), .B(i_12_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n350_), .B(mai_mai_n79_), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n351_), .B(mai_mai_n267_), .Y(mai_mai_n352_));
  AOI220     m330(.A0(mai_mai_n352_), .A1(mai_mai_n36_), .B0(mai_mai_n349_), .B1(mai_mai_n45_), .Y(mai_mai_n353_));
  NA4        m331(.A(mai_mai_n353_), .B(mai_mai_n346_), .C(mai_mai_n331_), .D(mai_mai_n326_), .Y(mai6));
  NO2        m332(.A(mai_mai_n123_), .B(i_11_), .Y(mai_mai_n355_));
  NO2        m333(.A(i_11_), .B(i_9_), .Y(mai_mai_n356_));
  NO2        m334(.A(mai_mai_n184_), .B(mai_mai_n158_), .Y(mai_mai_n357_));
  OR2        m335(.A(mai_mai_n357_), .B(i_12_), .Y(mai_mai_n358_));
  AOI220     m336(.A0(mai_mai_n109_), .A1(mai_mai_n356_), .B0(mai_mai_n173_), .B1(mai_mai_n54_), .Y(mai_mai_n359_));
  NA2        m337(.A(mai_mai_n430_), .B(mai_mai_n350_), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n360_), .A1(mai_mai_n237_), .B0(mai_mai_n104_), .Y(mai_mai_n361_));
  INV        m339(.A(i_11_), .Y(mai_mai_n362_));
  NA2        m340(.A(mai_mai_n362_), .B(mai_mai_n184_), .Y(mai_mai_n363_));
  NAi32      m341(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n364_));
  AOI210     m342(.A0(i_11_), .A1(i_11_), .B0(mai_mai_n364_), .Y(mai_mai_n365_));
  NA2        m343(.A(i_4_), .B(mai_mai_n259_), .Y(mai_mai_n366_));
  NAi31      m344(.An(mai_mai_n365_), .B(mai_mai_n366_), .C(mai_mai_n363_), .Y(mai_mai_n367_));
  OR2        m345(.A(mai_mai_n367_), .B(mai_mai_n361_), .Y(mai_mai_n368_));
  NA3        m346(.A(mai_mai_n439_), .B(mai_mai_n137_), .C(i_7_), .Y(mai_mai_n369_));
  NA2        m347(.A(mai_mai_n433_), .B(mai_mai_n90_), .Y(mai_mai_n370_));
  OR2        m348(.A(mai_mai_n323_), .B(mai_mai_n36_), .Y(mai_mai_n371_));
  NA3        m349(.A(mai_mai_n371_), .B(mai_mai_n370_), .C(mai_mai_n369_), .Y(mai_mai_n372_));
  INV        m350(.A(mai_mai_n355_), .Y(mai_mai_n373_));
  NA2        m351(.A(mai_mai_n131_), .B(mai_mai_n90_), .Y(mai_mai_n374_));
  OAI210     m352(.A0(mai_mai_n187_), .A1(mai_mai_n116_), .B0(mai_mai_n51_), .Y(mai_mai_n375_));
  NA4        m353(.A(mai_mai_n375_), .B(mai_mai_n374_), .C(mai_mai_n373_), .D(mai_mai_n269_), .Y(mai_mai_n376_));
  NA3        m354(.A(mai_mai_n239_), .B(mai_mai_n223_), .C(mai_mai_n122_), .Y(mai_mai_n377_));
  AOI210     m355(.A0(mai_mai_n204_), .A1(mai_mai_n203_), .B0(mai_mai_n258_), .Y(mai_mai_n378_));
  INV        m356(.A(mai_mai_n194_), .Y(mai_mai_n379_));
  NA3        m357(.A(mai_mai_n379_), .B(mai_mai_n378_), .C(mai_mai_n377_), .Y(mai_mai_n380_));
  NO4        m358(.A(mai_mai_n380_), .B(mai_mai_n376_), .C(mai_mai_n372_), .D(mai_mai_n368_), .Y(mai_mai_n381_));
  NA4        m359(.A(mai_mai_n381_), .B(mai_mai_n359_), .C(mai_mai_n358_), .D(mai_mai_n177_), .Y(mai3));
  NA2        m360(.A(mai_mai_n170_), .B(mai_mai_n39_), .Y(mai_mai_n383_));
  NO2        m361(.A(mai_mai_n383_), .B(mai_mai_n46_), .Y(mai_mai_n384_));
  NOi21      m362(.An(i_5_), .B(i_9_), .Y(mai_mai_n385_));
  NA2        m363(.A(mai_mai_n385_), .B(mai_mai_n202_), .Y(mai_mai_n386_));
  INV        m364(.A(mai_mai_n384_), .Y(mai_mai_n387_));
  NO4        m365(.A(i_5_), .B(i_12_), .C(mai_mai_n198_), .D(mai_mai_n195_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n388_), .B(i_11_), .Y(mai_mai_n389_));
  NA2        m367(.A(mai_mai_n321_), .B(mai_mai_n158_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n390_), .B(mai_mai_n389_), .Y(mai_mai_n391_));
  NA2        m369(.A(mai_mai_n186_), .B(mai_mai_n102_), .Y(mai_mai_n392_));
  NA3        m370(.A(mai_mai_n392_), .B(mai_mai_n208_), .C(mai_mai_n97_), .Y(mai_mai_n393_));
  NO2        m371(.A(i_12_), .B(mai_mai_n386_), .Y(mai_mai_n394_));
  NO2        m372(.A(mai_mai_n394_), .B(mai_mai_n393_), .Y(mai_mai_n395_));
  NA2        m373(.A(mai_mai_n294_), .B(i_1_), .Y(mai_mai_n396_));
  NO2        m374(.A(i_6_), .B(mai_mai_n396_), .Y(mai_mai_n397_));
  NA2        m375(.A(mai_mai_n100_), .B(mai_mai_n70_), .Y(mai_mai_n398_));
  INV        m376(.A(mai_mai_n397_), .Y(mai_mai_n399_));
  NA2        m377(.A(mai_mai_n399_), .B(mai_mai_n395_), .Y(mai_mai_n400_));
  NO3        m378(.A(i_5_), .B(i_0_), .C(mai_mai_n24_), .Y(mai_mai_n401_));
  INV        m379(.A(mai_mai_n401_), .Y(mai_mai_n402_));
  NAi21      m380(.An(i_9_), .B(i_5_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n403_), .B(mai_mai_n189_), .Y(mai_mai_n404_));
  NA2        m382(.A(mai_mai_n404_), .B(mai_mai_n275_), .Y(mai_mai_n405_));
  OAI220     m383(.A0(mai_mai_n405_), .A1(mai_mai_n61_), .B0(mai_mai_n402_), .B1(mai_mai_n101_), .Y(mai_mai_n406_));
  NO2        m384(.A(mai_mai_n406_), .B(mai_mai_n240_), .Y(mai_mai_n407_));
  NA2        m385(.A(mai_mai_n407_), .B(mai_mai_n106_), .Y(mai_mai_n408_));
  NO3        m386(.A(mai_mai_n408_), .B(mai_mai_n400_), .C(mai_mai_n391_), .Y(mai_mai_n409_));
  NO2        m387(.A(i_12_), .B(mai_mai_n398_), .Y(mai_mai_n410_));
  INV        m388(.A(mai_mai_n158_), .Y(mai_mai_n411_));
  NO2        m389(.A(mai_mai_n99_), .B(mai_mai_n411_), .Y(mai_mai_n412_));
  NO3        m390(.A(mai_mai_n119_), .B(mai_mai_n179_), .C(i_0_), .Y(mai_mai_n413_));
  OAI210     m391(.A0(mai_mai_n413_), .A1(mai_mai_n57_), .B0(i_13_), .Y(mai_mai_n414_));
  INV        m392(.A(mai_mai_n122_), .Y(mai_mai_n415_));
  NA3        m393(.A(mai_mai_n113_), .B(i_7_), .C(mai_mai_n415_), .Y(mai_mai_n416_));
  NA3        m394(.A(mai_mai_n416_), .B(mai_mai_n414_), .C(mai_mai_n429_), .Y(mai_mai_n417_));
  NA3        m395(.A(mai_mai_n184_), .B(mai_mai_n100_), .C(i_4_), .Y(mai_mai_n418_));
  NO3        m396(.A(mai_mai_n441_), .B(mai_mai_n417_), .C(mai_mai_n410_), .Y(mai_mai_n419_));
  NA2        m397(.A(mai_mai_n37_), .B(mai_mai_n117_), .Y(mai_mai_n420_));
  NO2        m398(.A(mai_mai_n420_), .B(mai_mai_n54_), .Y(mai_mai_n421_));
  INV        m399(.A(mai_mai_n258_), .Y(mai_mai_n422_));
  INV        m400(.A(mai_mai_n365_), .Y(mai_mai_n423_));
  AOI210     m401(.A0(mai_mai_n423_), .A1(mai_mai_n422_), .B0(mai_mai_n40_), .Y(mai_mai_n424_));
  NO2        m402(.A(mai_mai_n424_), .B(mai_mai_n421_), .Y(mai_mai_n425_));
  NA4        m403(.A(mai_mai_n425_), .B(mai_mai_n419_), .C(mai_mai_n409_), .D(mai_mai_n387_), .Y(mai4));
  INV        m404(.A(mai_mai_n412_), .Y(mai_mai_n429_));
  INV        m405(.A(i_9_), .Y(mai_mai_n430_));
  INV        m406(.A(mai_mai_n305_), .Y(mai_mai_n431_));
  INV        m407(.A(i_6_), .Y(mai_mai_n432_));
  INV        m408(.A(i_12_), .Y(mai_mai_n433_));
  INV        m409(.A(i_9_), .Y(mai_mai_n434_));
  INV        m410(.A(i_10_), .Y(mai_mai_n435_));
  INV        m411(.A(mai_mai_n57_), .Y(mai_mai_n436_));
  INV        m412(.A(mai_mai_n134_), .Y(mai_mai_n437_));
  INV        m413(.A(mai_mai_n263_), .Y(mai_mai_n438_));
  INV        m414(.A(i_9_), .Y(mai_mai_n439_));
  INV        m415(.A(i_2_), .Y(mai_mai_n440_));
  INV        m416(.A(mai_mai_n418_), .Y(mai_mai_n441_));
  INV        m417(.A(mai_mai_n26_), .Y(mai_mai_n442_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u0016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u0017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u0018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  NO2        u0028(.A(men_men_n50_), .B(i_3_), .Y(men_men_n51_));
  AOI210     u0029(.A0(men_men_n51_), .A1(men_men_n47_), .B0(men_men_n46_), .Y(men_men_n52_));
  NA2        u0030(.A(i_0_), .B(i_2_), .Y(men_men_n53_));
  NA2        u0031(.A(i_7_), .B(i_9_), .Y(men_men_n54_));
  NO2        u0032(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n52_), .B(men_men_n45_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n50_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(men_men_n81_), .B(men_men_n58_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_9_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_7_), .Y(men_men_n84_));
  NO3        u0062(.A(men_men_n84_), .B(men_men_n83_), .C(men_men_n63_), .Y(men_men_n85_));
  INV        u0063(.A(i_6_), .Y(men_men_n86_));
  OR4        u0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n87_));
  INV        u0065(.A(men_men_n87_), .Y(men_men_n88_));
  NO2        u0066(.A(i_2_), .B(i_7_), .Y(men_men_n89_));
  OAI210     u0067(.A0(men_men_n85_), .A1(men_men_n82_), .B0(i_2_), .Y(men_men_n90_));
  NAi21      u0068(.An(i_6_), .B(i_10_), .Y(men_men_n91_));
  NA2        u0069(.A(i_6_), .B(i_9_), .Y(men_men_n92_));
  AOI210     u0070(.A0(men_men_n92_), .A1(men_men_n91_), .B0(men_men_n63_), .Y(men_men_n93_));
  NA2        u0071(.A(i_2_), .B(i_6_), .Y(men_men_n94_));
  NO3        u0072(.A(men_men_n94_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n95_));
  NO2        u0073(.A(men_men_n95_), .B(men_men_n93_), .Y(men_men_n96_));
  AOI210     u0074(.A0(men_men_n96_), .A1(men_men_n90_), .B0(men_men_n80_), .Y(men_men_n97_));
  AN3        u0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n98_));
  NAi21      u0076(.An(i_6_), .B(i_11_), .Y(men_men_n99_));
  NO2        u0077(.A(i_5_), .B(i_8_), .Y(men_men_n100_));
  NOi21      u0078(.An(men_men_n100_), .B(men_men_n99_), .Y(men_men_n101_));
  NA2        u0079(.A(men_men_n101_), .B(men_men_n62_), .Y(men_men_n102_));
  INV        u0080(.A(i_7_), .Y(men_men_n103_));
  NA2        u0081(.A(men_men_n46_), .B(men_men_n103_), .Y(men_men_n104_));
  NO2        u0082(.A(i_0_), .B(i_5_), .Y(men_men_n105_));
  NO2        u0083(.A(men_men_n105_), .B(men_men_n86_), .Y(men_men_n106_));
  NA2        u0084(.A(i_12_), .B(i_3_), .Y(men_men_n107_));
  INV        u0085(.A(men_men_n107_), .Y(men_men_n108_));
  NA3        u0086(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n104_), .Y(men_men_n109_));
  NAi21      u0087(.An(i_7_), .B(i_11_), .Y(men_men_n110_));
  NO3        u0088(.A(men_men_n110_), .B(men_men_n91_), .C(men_men_n53_), .Y(men_men_n111_));
  AN2        u0089(.A(i_2_), .B(i_10_), .Y(men_men_n112_));
  NO2        u0090(.A(men_men_n112_), .B(i_7_), .Y(men_men_n113_));
  OR2        u0091(.A(men_men_n80_), .B(men_men_n58_), .Y(men_men_n114_));
  NO2        u0092(.A(i_8_), .B(men_men_n103_), .Y(men_men_n115_));
  NO3        u0093(.A(men_men_n115_), .B(men_men_n114_), .C(men_men_n113_), .Y(men_men_n116_));
  NA2        u0094(.A(i_12_), .B(i_7_), .Y(men_men_n117_));
  NO2        u0095(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n118_));
  INV        u0096(.A(men_men_n118_), .Y(men_men_n119_));
  NA2        u0097(.A(i_11_), .B(i_12_), .Y(men_men_n120_));
  OAI210     u0098(.A0(men_men_n119_), .A1(men_men_n117_), .B0(men_men_n120_), .Y(men_men_n121_));
  NO2        u0099(.A(men_men_n121_), .B(men_men_n116_), .Y(men_men_n122_));
  NA3        u0100(.A(men_men_n122_), .B(men_men_n109_), .C(men_men_n102_), .Y(men_men_n123_));
  NOi21      u0101(.An(i_1_), .B(i_5_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(i_11_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n103_), .B(men_men_n37_), .Y(men_men_n126_));
  NA2        u0104(.A(i_7_), .B(men_men_n25_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n128_));
  NO2        u0106(.A(men_men_n128_), .B(men_men_n46_), .Y(men_men_n129_));
  NA2        u0107(.A(men_men_n92_), .B(men_men_n91_), .Y(men_men_n130_));
  NAi21      u0108(.An(i_3_), .B(i_8_), .Y(men_men_n131_));
  NA2        u0109(.A(men_men_n131_), .B(men_men_n62_), .Y(men_men_n132_));
  NOi31      u0110(.An(men_men_n132_), .B(men_men_n130_), .C(men_men_n129_), .Y(men_men_n133_));
  NO2        u0111(.A(i_1_), .B(men_men_n86_), .Y(men_men_n134_));
  NO2        u0112(.A(i_6_), .B(i_5_), .Y(men_men_n135_));
  NA2        u0113(.A(men_men_n135_), .B(i_3_), .Y(men_men_n136_));
  AO210      u0114(.A0(men_men_n136_), .A1(men_men_n47_), .B0(men_men_n134_), .Y(men_men_n137_));
  OAI220     u0115(.A0(men_men_n137_), .A1(men_men_n110_), .B0(men_men_n133_), .B1(men_men_n125_), .Y(men_men_n138_));
  NO3        u0116(.A(men_men_n138_), .B(men_men_n123_), .C(men_men_n97_), .Y(men_men_n139_));
  NA3        u0117(.A(men_men_n139_), .B(men_men_n79_), .C(men_men_n56_), .Y(men2));
  NO2        u0118(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n141_));
  NA2        u0119(.A(i_6_), .B(men_men_n25_), .Y(men_men_n142_));
  NA3        u0120(.A(men_men_n77_), .B(men_men_n69_), .C(men_men_n30_), .Y(men0));
  AN2        u0121(.A(i_8_), .B(i_7_), .Y(men_men_n144_));
  NA2        u0122(.A(men_men_n144_), .B(i_6_), .Y(men_men_n145_));
  NO2        u0123(.A(i_12_), .B(i_13_), .Y(men_men_n146_));
  NAi21      u0124(.An(i_5_), .B(i_11_), .Y(men_men_n147_));
  NOi21      u0125(.An(men_men_n146_), .B(men_men_n147_), .Y(men_men_n148_));
  NO2        u0126(.A(i_0_), .B(i_1_), .Y(men_men_n149_));
  NA2        u0127(.A(i_2_), .B(i_3_), .Y(men_men_n150_));
  NO2        u0128(.A(men_men_n150_), .B(i_4_), .Y(men_men_n151_));
  NA3        u0129(.A(men_men_n151_), .B(men_men_n149_), .C(men_men_n148_), .Y(men_men_n152_));
  OR2        u0130(.A(men_men_n152_), .B(men_men_n25_), .Y(men_men_n153_));
  AN2        u0131(.A(men_men_n146_), .B(men_men_n83_), .Y(men_men_n154_));
  NO2        u0132(.A(men_men_n154_), .B(men_men_n27_), .Y(men_men_n155_));
  NA2        u0133(.A(i_1_), .B(i_5_), .Y(men_men_n156_));
  NO2        u0134(.A(men_men_n73_), .B(men_men_n46_), .Y(men_men_n157_));
  NA2        u0135(.A(men_men_n157_), .B(men_men_n36_), .Y(men_men_n158_));
  NO3        u0136(.A(men_men_n158_), .B(men_men_n156_), .C(men_men_n155_), .Y(men_men_n159_));
  OR2        u0137(.A(i_0_), .B(i_1_), .Y(men_men_n160_));
  NO3        u0138(.A(men_men_n160_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n161_));
  NAi32      u0139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n162_));
  NAi21      u0140(.An(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  NOi21      u0141(.An(i_4_), .B(i_10_), .Y(men_men_n164_));
  NA2        u0142(.A(men_men_n164_), .B(men_men_n39_), .Y(men_men_n165_));
  NO2        u0143(.A(i_3_), .B(i_5_), .Y(men_men_n166_));
  NO3        u0144(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n167_));
  NA2        u0145(.A(men_men_n167_), .B(men_men_n166_), .Y(men_men_n168_));
  OAI210     u0146(.A0(men_men_n168_), .A1(men_men_n165_), .B0(men_men_n163_), .Y(men_men_n169_));
  NO2        u0147(.A(men_men_n169_), .B(men_men_n159_), .Y(men_men_n170_));
  AOI210     u0148(.A0(men_men_n170_), .A1(men_men_n153_), .B0(men_men_n145_), .Y(men_men_n171_));
  NA3        u0149(.A(men_men_n73_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n172_));
  NA2        u0150(.A(i_3_), .B(men_men_n48_), .Y(men_men_n173_));
  NOi21      u0151(.An(i_4_), .B(i_9_), .Y(men_men_n174_));
  NOi21      u0152(.An(i_11_), .B(i_13_), .Y(men_men_n175_));
  NA2        u0153(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  OR2        u0154(.A(men_men_n176_), .B(men_men_n173_), .Y(men_men_n177_));
  NO2        u0155(.A(i_4_), .B(i_5_), .Y(men_men_n178_));
  NAi21      u0156(.An(i_12_), .B(i_11_), .Y(men_men_n179_));
  NO2        u0157(.A(men_men_n179_), .B(i_13_), .Y(men_men_n180_));
  NA3        u0158(.A(men_men_n180_), .B(men_men_n178_), .C(men_men_n83_), .Y(men_men_n181_));
  AOI210     u0159(.A0(men_men_n181_), .A1(men_men_n177_), .B0(men_men_n172_), .Y(men_men_n182_));
  NO2        u0160(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n183_));
  NA2        u0161(.A(men_men_n183_), .B(men_men_n46_), .Y(men_men_n184_));
  NA2        u0162(.A(men_men_n36_), .B(i_5_), .Y(men_men_n185_));
  NAi31      u0163(.An(men_men_n185_), .B(men_men_n154_), .C(i_11_), .Y(men_men_n186_));
  NA2        u0164(.A(i_3_), .B(i_5_), .Y(men_men_n187_));
  OR2        u0165(.A(men_men_n187_), .B(men_men_n176_), .Y(men_men_n188_));
  AOI210     u0166(.A0(men_men_n188_), .A1(men_men_n186_), .B0(men_men_n184_), .Y(men_men_n189_));
  NO2        u0167(.A(men_men_n73_), .B(i_5_), .Y(men_men_n190_));
  NO2        u0168(.A(i_13_), .B(i_10_), .Y(men_men_n191_));
  NA3        u0169(.A(men_men_n191_), .B(men_men_n190_), .C(men_men_n44_), .Y(men_men_n192_));
  NO2        u0170(.A(i_2_), .B(i_1_), .Y(men_men_n193_));
  NA2        u0171(.A(men_men_n193_), .B(i_3_), .Y(men_men_n194_));
  NAi21      u0172(.An(i_4_), .B(i_12_), .Y(men_men_n195_));
  NO4        u0173(.A(men_men_n195_), .B(men_men_n194_), .C(men_men_n192_), .D(men_men_n25_), .Y(men_men_n196_));
  NO3        u0174(.A(men_men_n196_), .B(men_men_n189_), .C(men_men_n182_), .Y(men_men_n197_));
  INV        u0175(.A(i_8_), .Y(men_men_n198_));
  NO2        u0176(.A(men_men_n198_), .B(i_7_), .Y(men_men_n199_));
  NA2        u0177(.A(men_men_n199_), .B(i_6_), .Y(men_men_n200_));
  NO3        u0178(.A(i_3_), .B(men_men_n86_), .C(men_men_n48_), .Y(men_men_n201_));
  NA2        u0179(.A(men_men_n201_), .B(men_men_n115_), .Y(men_men_n202_));
  NO3        u0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n203_));
  NA3        u0181(.A(men_men_n203_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n204_));
  NO3        u0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n205_));
  OAI210     u0183(.A0(men_men_n98_), .A1(i_12_), .B0(men_men_n205_), .Y(men_men_n206_));
  AOI210     u0184(.A0(men_men_n206_), .A1(men_men_n204_), .B0(men_men_n202_), .Y(men_men_n207_));
  NO2        u0185(.A(i_3_), .B(i_8_), .Y(men_men_n208_));
  NO3        u0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n209_));
  NA3        u0187(.A(men_men_n209_), .B(men_men_n208_), .C(men_men_n39_), .Y(men_men_n210_));
  NO2        u0188(.A(men_men_n105_), .B(men_men_n58_), .Y(men_men_n211_));
  INV        u0189(.A(men_men_n211_), .Y(men_men_n212_));
  NO2        u0190(.A(i_13_), .B(i_9_), .Y(men_men_n213_));
  NA3        u0191(.A(men_men_n213_), .B(i_6_), .C(men_men_n198_), .Y(men_men_n214_));
  NAi21      u0192(.An(i_12_), .B(i_3_), .Y(men_men_n215_));
  OR2        u0193(.A(men_men_n215_), .B(men_men_n214_), .Y(men_men_n216_));
  NO2        u0194(.A(men_men_n44_), .B(i_5_), .Y(men_men_n217_));
  NO3        u0195(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n218_));
  NA3        u0196(.A(men_men_n218_), .B(men_men_n217_), .C(i_10_), .Y(men_men_n219_));
  OAI220     u0197(.A0(men_men_n219_), .A1(men_men_n216_), .B0(men_men_n212_), .B1(men_men_n210_), .Y(men_men_n220_));
  AOI210     u0198(.A0(men_men_n220_), .A1(i_7_), .B0(men_men_n207_), .Y(men_men_n221_));
  OAI220     u0199(.A0(men_men_n221_), .A1(i_4_), .B0(men_men_n200_), .B1(men_men_n197_), .Y(men_men_n222_));
  NAi21      u0200(.An(i_12_), .B(i_7_), .Y(men_men_n223_));
  NA3        u0201(.A(i_13_), .B(men_men_n198_), .C(i_10_), .Y(men_men_n224_));
  NO2        u0202(.A(men_men_n224_), .B(men_men_n223_), .Y(men_men_n225_));
  NA2        u0203(.A(i_0_), .B(i_5_), .Y(men_men_n226_));
  NA2        u0204(.A(men_men_n226_), .B(men_men_n106_), .Y(men_men_n227_));
  OAI220     u0205(.A0(men_men_n227_), .A1(men_men_n194_), .B0(men_men_n184_), .B1(men_men_n136_), .Y(men_men_n228_));
  NAi31      u0206(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n229_));
  NO2        u0207(.A(men_men_n36_), .B(i_13_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n73_), .B(men_men_n26_), .Y(men_men_n231_));
  NO2        u0209(.A(men_men_n46_), .B(men_men_n63_), .Y(men_men_n232_));
  NA3        u0210(.A(men_men_n232_), .B(men_men_n231_), .C(men_men_n230_), .Y(men_men_n233_));
  INV        u0211(.A(i_13_), .Y(men_men_n234_));
  NO2        u0212(.A(i_12_), .B(men_men_n234_), .Y(men_men_n235_));
  NA3        u0213(.A(men_men_n235_), .B(men_men_n203_), .C(men_men_n201_), .Y(men_men_n236_));
  OAI210     u0214(.A0(men_men_n233_), .A1(men_men_n229_), .B0(men_men_n236_), .Y(men_men_n237_));
  AOI220     u0215(.A0(men_men_n237_), .A1(men_men_n144_), .B0(men_men_n228_), .B1(men_men_n225_), .Y(men_men_n238_));
  NO2        u0216(.A(i_12_), .B(men_men_n37_), .Y(men_men_n239_));
  NO2        u0217(.A(men_men_n187_), .B(i_4_), .Y(men_men_n240_));
  NA2        u0218(.A(men_men_n240_), .B(men_men_n239_), .Y(men_men_n241_));
  OR2        u0219(.A(i_8_), .B(i_7_), .Y(men_men_n242_));
  NO2        u0220(.A(men_men_n242_), .B(men_men_n86_), .Y(men_men_n243_));
  NO2        u0221(.A(men_men_n53_), .B(i_1_), .Y(men_men_n244_));
  NA2        u0222(.A(men_men_n244_), .B(men_men_n243_), .Y(men_men_n245_));
  INV        u0223(.A(i_12_), .Y(men_men_n246_));
  NO2        u0224(.A(men_men_n44_), .B(men_men_n246_), .Y(men_men_n247_));
  NO3        u0225(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n248_));
  NA2        u0226(.A(i_2_), .B(i_1_), .Y(men_men_n249_));
  NO2        u0227(.A(men_men_n245_), .B(men_men_n241_), .Y(men_men_n250_));
  NO3        u0228(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n251_));
  NAi21      u0229(.An(i_4_), .B(i_3_), .Y(men_men_n252_));
  NO2        u0230(.A(men_men_n252_), .B(men_men_n75_), .Y(men_men_n253_));
  NO2        u0231(.A(i_0_), .B(i_6_), .Y(men_men_n254_));
  NOi41      u0232(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n255_));
  NA2        u0233(.A(men_men_n255_), .B(men_men_n254_), .Y(men_men_n256_));
  NO2        u0234(.A(men_men_n249_), .B(men_men_n187_), .Y(men_men_n257_));
  NAi21      u0235(.An(men_men_n256_), .B(men_men_n257_), .Y(men_men_n258_));
  INV        u0236(.A(men_men_n258_), .Y(men_men_n259_));
  AOI220     u0237(.A0(men_men_n259_), .A1(men_men_n39_), .B0(men_men_n250_), .B1(men_men_n213_), .Y(men_men_n260_));
  NO2        u0238(.A(i_11_), .B(men_men_n234_), .Y(men_men_n261_));
  NOi21      u0239(.An(i_1_), .B(i_6_), .Y(men_men_n262_));
  NAi21      u0240(.An(i_3_), .B(i_7_), .Y(men_men_n263_));
  NA2        u0241(.A(men_men_n246_), .B(i_9_), .Y(men_men_n264_));
  OR4        u0242(.A(men_men_n264_), .B(men_men_n263_), .C(men_men_n262_), .D(men_men_n190_), .Y(men_men_n265_));
  NO2        u0243(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n266_));
  NO2        u0244(.A(i_12_), .B(i_3_), .Y(men_men_n267_));
  NA2        u0245(.A(men_men_n73_), .B(i_5_), .Y(men_men_n268_));
  NA2        u0246(.A(i_3_), .B(i_9_), .Y(men_men_n269_));
  NAi21      u0247(.An(i_7_), .B(i_10_), .Y(men_men_n270_));
  NO2        u0248(.A(men_men_n270_), .B(men_men_n269_), .Y(men_men_n271_));
  NA3        u0249(.A(men_men_n271_), .B(men_men_n268_), .C(men_men_n64_), .Y(men_men_n272_));
  NA2        u0250(.A(men_men_n272_), .B(men_men_n265_), .Y(men_men_n273_));
  NA3        u0251(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n274_));
  INV        u0252(.A(men_men_n145_), .Y(men_men_n275_));
  NA2        u0253(.A(men_men_n246_), .B(i_13_), .Y(men_men_n276_));
  NO2        u0254(.A(men_men_n276_), .B(men_men_n75_), .Y(men_men_n277_));
  AOI220     u0255(.A0(men_men_n277_), .A1(men_men_n275_), .B0(men_men_n273_), .B1(men_men_n261_), .Y(men_men_n278_));
  NO2        u0256(.A(men_men_n242_), .B(men_men_n37_), .Y(men_men_n279_));
  NA2        u0257(.A(i_12_), .B(i_6_), .Y(men_men_n280_));
  OR2        u0258(.A(i_13_), .B(i_9_), .Y(men_men_n281_));
  NO3        u0259(.A(men_men_n281_), .B(men_men_n280_), .C(men_men_n48_), .Y(men_men_n282_));
  NO2        u0260(.A(men_men_n252_), .B(i_2_), .Y(men_men_n283_));
  NA3        u0261(.A(men_men_n283_), .B(men_men_n282_), .C(men_men_n44_), .Y(men_men_n284_));
  NA2        u0262(.A(men_men_n261_), .B(i_9_), .Y(men_men_n285_));
  NA2        u0263(.A(men_men_n268_), .B(men_men_n64_), .Y(men_men_n286_));
  OAI210     u0264(.A0(men_men_n286_), .A1(men_men_n285_), .B0(men_men_n284_), .Y(men_men_n287_));
  NA2        u0265(.A(men_men_n157_), .B(men_men_n63_), .Y(men_men_n288_));
  NO3        u0266(.A(i_11_), .B(men_men_n234_), .C(men_men_n25_), .Y(men_men_n289_));
  NO2        u0267(.A(men_men_n263_), .B(i_8_), .Y(men_men_n290_));
  NO2        u0268(.A(i_6_), .B(men_men_n48_), .Y(men_men_n291_));
  NA3        u0269(.A(men_men_n291_), .B(men_men_n290_), .C(men_men_n289_), .Y(men_men_n292_));
  NO3        u0270(.A(men_men_n26_), .B(men_men_n86_), .C(i_5_), .Y(men_men_n293_));
  NA3        u0271(.A(men_men_n293_), .B(men_men_n279_), .C(men_men_n235_), .Y(men_men_n294_));
  AOI210     u0272(.A0(men_men_n294_), .A1(men_men_n292_), .B0(men_men_n288_), .Y(men_men_n295_));
  AOI210     u0273(.A0(men_men_n287_), .A1(men_men_n279_), .B0(men_men_n295_), .Y(men_men_n296_));
  NA4        u0274(.A(men_men_n296_), .B(men_men_n278_), .C(men_men_n260_), .D(men_men_n238_), .Y(men_men_n297_));
  NO3        u0275(.A(i_12_), .B(men_men_n234_), .C(men_men_n37_), .Y(men_men_n298_));
  INV        u0276(.A(men_men_n298_), .Y(men_men_n299_));
  NA2        u0277(.A(i_8_), .B(men_men_n103_), .Y(men_men_n300_));
  NOi21      u0278(.An(men_men_n166_), .B(men_men_n86_), .Y(men_men_n301_));
  NO3        u0279(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n302_));
  AOI220     u0280(.A0(men_men_n302_), .A1(men_men_n201_), .B0(men_men_n301_), .B1(men_men_n244_), .Y(men_men_n303_));
  NO2        u0281(.A(men_men_n303_), .B(men_men_n300_), .Y(men_men_n304_));
  NO3        u0282(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n305_));
  NO2        u0283(.A(men_men_n249_), .B(i_0_), .Y(men_men_n306_));
  AOI220     u0284(.A0(men_men_n306_), .A1(men_men_n199_), .B0(men_men_n305_), .B1(men_men_n144_), .Y(men_men_n307_));
  NA2        u0285(.A(men_men_n291_), .B(men_men_n26_), .Y(men_men_n308_));
  NO2        u0286(.A(men_men_n308_), .B(men_men_n307_), .Y(men_men_n309_));
  NA2        u0287(.A(i_0_), .B(i_1_), .Y(men_men_n310_));
  NO2        u0288(.A(men_men_n310_), .B(i_2_), .Y(men_men_n311_));
  NO2        u0289(.A(men_men_n59_), .B(i_6_), .Y(men_men_n312_));
  NA3        u0290(.A(men_men_n312_), .B(men_men_n311_), .C(men_men_n166_), .Y(men_men_n313_));
  OAI210     u0291(.A0(men_men_n168_), .A1(men_men_n145_), .B0(men_men_n313_), .Y(men_men_n314_));
  NO3        u0292(.A(men_men_n314_), .B(men_men_n309_), .C(men_men_n304_), .Y(men_men_n315_));
  NO2        u0293(.A(i_3_), .B(i_10_), .Y(men_men_n316_));
  NA3        u0294(.A(men_men_n316_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n317_));
  NO2        u0295(.A(i_2_), .B(men_men_n103_), .Y(men_men_n318_));
  NA2        u0296(.A(i_1_), .B(men_men_n36_), .Y(men_men_n319_));
  NO2        u0297(.A(men_men_n319_), .B(i_8_), .Y(men_men_n320_));
  NOi21      u0298(.An(men_men_n226_), .B(men_men_n105_), .Y(men_men_n321_));
  NA3        u0299(.A(men_men_n321_), .B(men_men_n320_), .C(men_men_n318_), .Y(men_men_n322_));
  AN2        u0300(.A(i_3_), .B(i_10_), .Y(men_men_n323_));
  NA4        u0301(.A(men_men_n323_), .B(men_men_n203_), .C(men_men_n180_), .D(men_men_n178_), .Y(men_men_n324_));
  NO2        u0302(.A(i_5_), .B(men_men_n37_), .Y(men_men_n325_));
  NO2        u0303(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n326_));
  OR2        u0304(.A(men_men_n322_), .B(men_men_n317_), .Y(men_men_n327_));
  OAI220     u0305(.A0(men_men_n327_), .A1(i_6_), .B0(men_men_n315_), .B1(men_men_n299_), .Y(men_men_n328_));
  NO4        u0306(.A(men_men_n328_), .B(men_men_n297_), .C(men_men_n222_), .D(men_men_n171_), .Y(men_men_n329_));
  NO3        u0307(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n330_));
  NO2        u0308(.A(men_men_n59_), .B(men_men_n86_), .Y(men_men_n331_));
  NA2        u0309(.A(men_men_n306_), .B(men_men_n331_), .Y(men_men_n332_));
  NO3        u0310(.A(i_6_), .B(men_men_n198_), .C(i_7_), .Y(men_men_n333_));
  NA2        u0311(.A(men_men_n333_), .B(men_men_n203_), .Y(men_men_n334_));
  AOI210     u0312(.A0(men_men_n334_), .A1(men_men_n332_), .B0(men_men_n173_), .Y(men_men_n335_));
  NO2        u0313(.A(i_2_), .B(i_3_), .Y(men_men_n336_));
  OR2        u0314(.A(i_0_), .B(i_5_), .Y(men_men_n337_));
  NA2        u0315(.A(men_men_n226_), .B(men_men_n337_), .Y(men_men_n338_));
  NA4        u0316(.A(men_men_n338_), .B(men_men_n243_), .C(men_men_n336_), .D(i_1_), .Y(men_men_n339_));
  NA3        u0317(.A(men_men_n306_), .B(men_men_n301_), .C(men_men_n115_), .Y(men_men_n340_));
  NAi21      u0318(.An(i_8_), .B(i_7_), .Y(men_men_n341_));
  NO2        u0319(.A(men_men_n341_), .B(i_6_), .Y(men_men_n342_));
  NO2        u0320(.A(men_men_n160_), .B(men_men_n46_), .Y(men_men_n343_));
  NA3        u0321(.A(men_men_n343_), .B(men_men_n342_), .C(men_men_n166_), .Y(men_men_n344_));
  NA3        u0322(.A(men_men_n344_), .B(men_men_n340_), .C(men_men_n339_), .Y(men_men_n345_));
  OAI210     u0323(.A0(men_men_n345_), .A1(men_men_n335_), .B0(i_4_), .Y(men_men_n346_));
  NO2        u0324(.A(i_12_), .B(i_10_), .Y(men_men_n347_));
  NOi21      u0325(.An(i_5_), .B(i_0_), .Y(men_men_n348_));
  AOI210     u0326(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n103_), .Y(men_men_n349_));
  NO4        u0327(.A(men_men_n349_), .B(men_men_n319_), .C(men_men_n348_), .D(men_men_n131_), .Y(men_men_n350_));
  NA4        u0328(.A(men_men_n84_), .B(men_men_n36_), .C(men_men_n86_), .D(i_8_), .Y(men_men_n351_));
  NA2        u0329(.A(men_men_n350_), .B(men_men_n347_), .Y(men_men_n352_));
  NO2        u0330(.A(i_6_), .B(i_8_), .Y(men_men_n353_));
  NOi21      u0331(.An(i_0_), .B(i_2_), .Y(men_men_n354_));
  AN2        u0332(.A(men_men_n354_), .B(men_men_n353_), .Y(men_men_n355_));
  NO2        u0333(.A(i_1_), .B(i_7_), .Y(men_men_n356_));
  AO220      u0334(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n342_), .B1(men_men_n244_), .Y(men_men_n357_));
  NA3        u0335(.A(men_men_n357_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n358_));
  NA3        u0336(.A(men_men_n358_), .B(men_men_n352_), .C(men_men_n346_), .Y(men_men_n359_));
  NO3        u0337(.A(men_men_n242_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n360_));
  NO3        u0338(.A(men_men_n341_), .B(i_2_), .C(i_1_), .Y(men_men_n361_));
  OAI210     u0339(.A0(men_men_n361_), .A1(men_men_n360_), .B0(i_6_), .Y(men_men_n362_));
  NA3        u0340(.A(men_men_n262_), .B(men_men_n318_), .C(men_men_n198_), .Y(men_men_n363_));
  AOI210     u0341(.A0(men_men_n363_), .A1(men_men_n362_), .B0(men_men_n338_), .Y(men_men_n364_));
  NOi21      u0342(.An(men_men_n156_), .B(men_men_n106_), .Y(men_men_n365_));
  NO2        u0343(.A(men_men_n365_), .B(men_men_n127_), .Y(men_men_n366_));
  OAI210     u0344(.A0(men_men_n366_), .A1(men_men_n364_), .B0(i_3_), .Y(men_men_n367_));
  INV        u0345(.A(men_men_n84_), .Y(men_men_n368_));
  NO2        u0346(.A(men_men_n310_), .B(men_men_n81_), .Y(men_men_n369_));
  NA2        u0347(.A(men_men_n369_), .B(men_men_n135_), .Y(men_men_n370_));
  NO2        u0348(.A(men_men_n94_), .B(men_men_n198_), .Y(men_men_n371_));
  NA3        u0349(.A(men_men_n321_), .B(men_men_n371_), .C(men_men_n63_), .Y(men_men_n372_));
  AOI210     u0350(.A0(men_men_n372_), .A1(men_men_n370_), .B0(men_men_n368_), .Y(men_men_n373_));
  NO2        u0351(.A(men_men_n198_), .B(i_9_), .Y(men_men_n374_));
  NA2        u0352(.A(men_men_n374_), .B(men_men_n211_), .Y(men_men_n375_));
  NO2        u0353(.A(men_men_n375_), .B(men_men_n46_), .Y(men_men_n376_));
  NO3        u0354(.A(men_men_n376_), .B(men_men_n373_), .C(men_men_n309_), .Y(men_men_n377_));
  AOI210     u0355(.A0(men_men_n377_), .A1(men_men_n367_), .B0(men_men_n165_), .Y(men_men_n378_));
  AOI210     u0356(.A0(men_men_n359_), .A1(men_men_n330_), .B0(men_men_n378_), .Y(men_men_n379_));
  NOi32      u0357(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n380_));
  INV        u0358(.A(men_men_n380_), .Y(men_men_n381_));
  NAi21      u0359(.An(i_0_), .B(i_6_), .Y(men_men_n382_));
  NAi21      u0360(.An(i_1_), .B(i_5_), .Y(men_men_n383_));
  NA2        u0361(.A(men_men_n383_), .B(men_men_n382_), .Y(men_men_n384_));
  NA2        u0362(.A(men_men_n384_), .B(men_men_n25_), .Y(men_men_n385_));
  OAI210     u0363(.A0(men_men_n385_), .A1(men_men_n162_), .B0(men_men_n256_), .Y(men_men_n386_));
  NAi41      u0364(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n387_));
  OAI220     u0365(.A0(men_men_n387_), .A1(men_men_n383_), .B0(men_men_n229_), .B1(men_men_n162_), .Y(men_men_n388_));
  AOI210     u0366(.A0(men_men_n387_), .A1(men_men_n162_), .B0(men_men_n160_), .Y(men_men_n389_));
  NOi32      u0367(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n390_));
  NAi21      u0368(.An(i_6_), .B(i_1_), .Y(men_men_n391_));
  NA3        u0369(.A(men_men_n391_), .B(men_men_n390_), .C(men_men_n46_), .Y(men_men_n392_));
  NO2        u0370(.A(men_men_n392_), .B(i_0_), .Y(men_men_n393_));
  OR3        u0371(.A(men_men_n393_), .B(men_men_n389_), .C(men_men_n388_), .Y(men_men_n394_));
  NO2        u0372(.A(i_1_), .B(men_men_n103_), .Y(men_men_n395_));
  NAi21      u0373(.An(i_3_), .B(i_4_), .Y(men_men_n396_));
  NO2        u0374(.A(men_men_n396_), .B(i_9_), .Y(men_men_n397_));
  AN2        u0375(.A(i_6_), .B(i_7_), .Y(men_men_n398_));
  OAI210     u0376(.A0(men_men_n398_), .A1(men_men_n395_), .B0(men_men_n397_), .Y(men_men_n399_));
  NA2        u0377(.A(i_2_), .B(i_7_), .Y(men_men_n400_));
  NO2        u0378(.A(men_men_n396_), .B(i_10_), .Y(men_men_n401_));
  NA3        u0379(.A(men_men_n401_), .B(men_men_n400_), .C(men_men_n254_), .Y(men_men_n402_));
  AOI210     u0380(.A0(men_men_n402_), .A1(men_men_n399_), .B0(men_men_n190_), .Y(men_men_n403_));
  AOI210     u0381(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n404_));
  OAI210     u0382(.A0(men_men_n404_), .A1(men_men_n193_), .B0(men_men_n401_), .Y(men_men_n405_));
  AOI220     u0383(.A0(men_men_n401_), .A1(men_men_n356_), .B0(men_men_n248_), .B1(men_men_n193_), .Y(men_men_n406_));
  AOI210     u0384(.A0(men_men_n406_), .A1(men_men_n405_), .B0(i_5_), .Y(men_men_n407_));
  NO4        u0385(.A(men_men_n407_), .B(men_men_n403_), .C(men_men_n394_), .D(men_men_n386_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n408_), .B(men_men_n381_), .Y(men_men_n409_));
  NO2        u0387(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n410_));
  AN2        u0388(.A(i_12_), .B(i_5_), .Y(men_men_n411_));
  NO2        u0389(.A(i_4_), .B(men_men_n26_), .Y(men_men_n412_));
  NA2        u0390(.A(men_men_n412_), .B(men_men_n411_), .Y(men_men_n413_));
  NO2        u0391(.A(i_11_), .B(i_6_), .Y(men_men_n414_));
  NA3        u0392(.A(men_men_n414_), .B(men_men_n343_), .C(men_men_n234_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n415_), .B(men_men_n413_), .Y(men_men_n416_));
  NO2        u0394(.A(men_men_n252_), .B(i_5_), .Y(men_men_n417_));
  NO2        u0395(.A(i_5_), .B(i_10_), .Y(men_men_n418_));
  AOI220     u0396(.A0(men_men_n418_), .A1(men_men_n283_), .B0(men_men_n417_), .B1(men_men_n203_), .Y(men_men_n419_));
  NA2        u0397(.A(men_men_n146_), .B(men_men_n45_), .Y(men_men_n420_));
  NO2        u0398(.A(men_men_n420_), .B(men_men_n419_), .Y(men_men_n421_));
  OAI210     u0399(.A0(men_men_n421_), .A1(men_men_n416_), .B0(men_men_n410_), .Y(men_men_n422_));
  NO2        u0400(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n423_));
  NO2        u0401(.A(men_men_n152_), .B(men_men_n86_), .Y(men_men_n424_));
  OAI210     u0402(.A0(men_men_n424_), .A1(men_men_n416_), .B0(men_men_n423_), .Y(men_men_n425_));
  NO3        u0403(.A(men_men_n86_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n426_));
  NO2        u0404(.A(i_3_), .B(men_men_n103_), .Y(men_men_n427_));
  NA3        u0405(.A(men_men_n316_), .B(men_men_n75_), .C(men_men_n54_), .Y(men_men_n428_));
  NO2        u0406(.A(i_11_), .B(i_12_), .Y(men_men_n429_));
  NA2        u0407(.A(men_men_n429_), .B(men_men_n36_), .Y(men_men_n430_));
  NO2        u0408(.A(men_men_n428_), .B(men_men_n430_), .Y(men_men_n431_));
  NA2        u0409(.A(men_men_n418_), .B(men_men_n246_), .Y(men_men_n432_));
  NA3        u0410(.A(men_men_n115_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n433_));
  NO2        u0411(.A(men_men_n433_), .B(men_men_n229_), .Y(men_men_n434_));
  NAi21      u0412(.An(i_13_), .B(i_0_), .Y(men_men_n435_));
  NO2        u0413(.A(men_men_n435_), .B(men_men_n249_), .Y(men_men_n436_));
  OAI210     u0414(.A0(men_men_n434_), .A1(men_men_n431_), .B0(men_men_n436_), .Y(men_men_n437_));
  NA3        u0415(.A(men_men_n437_), .B(men_men_n425_), .C(men_men_n422_), .Y(men_men_n438_));
  NA2        u0416(.A(men_men_n44_), .B(men_men_n234_), .Y(men_men_n439_));
  NO3        u0417(.A(i_1_), .B(i_12_), .C(men_men_n86_), .Y(men_men_n440_));
  NO2        u0418(.A(i_0_), .B(i_11_), .Y(men_men_n441_));
  AN2        u0419(.A(i_1_), .B(i_6_), .Y(men_men_n442_));
  NOi21      u0420(.An(i_2_), .B(i_12_), .Y(men_men_n443_));
  NA2        u0421(.A(men_men_n443_), .B(men_men_n442_), .Y(men_men_n444_));
  NO2        u0422(.A(men_men_n444_), .B(men_men_n1147_), .Y(men_men_n445_));
  NA2        u0423(.A(men_men_n144_), .B(i_9_), .Y(men_men_n446_));
  NO2        u0424(.A(men_men_n446_), .B(i_4_), .Y(men_men_n447_));
  NA2        u0425(.A(men_men_n445_), .B(men_men_n447_), .Y(men_men_n448_));
  NAi21      u0426(.An(i_9_), .B(i_4_), .Y(men_men_n449_));
  OR2        u0427(.A(i_13_), .B(i_10_), .Y(men_men_n450_));
  NO3        u0428(.A(men_men_n450_), .B(men_men_n120_), .C(men_men_n449_), .Y(men_men_n451_));
  NO2        u0429(.A(men_men_n176_), .B(men_men_n126_), .Y(men_men_n452_));
  OR2        u0430(.A(men_men_n224_), .B(men_men_n223_), .Y(men_men_n453_));
  NO2        u0431(.A(men_men_n103_), .B(men_men_n25_), .Y(men_men_n454_));
  NA2        u0432(.A(men_men_n298_), .B(men_men_n454_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n291_), .B(men_men_n218_), .Y(men_men_n456_));
  OAI220     u0434(.A0(men_men_n456_), .A1(men_men_n453_), .B0(men_men_n455_), .B1(men_men_n365_), .Y(men_men_n457_));
  INV        u0435(.A(men_men_n457_), .Y(men_men_n458_));
  AOI210     u0436(.A0(men_men_n458_), .A1(men_men_n448_), .B0(men_men_n26_), .Y(men_men_n459_));
  NA2        u0437(.A(men_men_n340_), .B(men_men_n339_), .Y(men_men_n460_));
  AOI220     u0438(.A0(men_men_n312_), .A1(men_men_n302_), .B0(men_men_n306_), .B1(men_men_n331_), .Y(men_men_n461_));
  NO2        u0439(.A(men_men_n461_), .B(men_men_n173_), .Y(men_men_n462_));
  NO2        u0440(.A(men_men_n187_), .B(men_men_n86_), .Y(men_men_n463_));
  AOI220     u0441(.A0(men_men_n463_), .A1(men_men_n311_), .B0(men_men_n293_), .B1(men_men_n218_), .Y(men_men_n464_));
  NO2        u0442(.A(men_men_n464_), .B(men_men_n300_), .Y(men_men_n465_));
  NO3        u0443(.A(men_men_n465_), .B(men_men_n462_), .C(men_men_n460_), .Y(men_men_n466_));
  NA2        u0444(.A(men_men_n201_), .B(men_men_n98_), .Y(men_men_n467_));
  NA3        u0445(.A(men_men_n343_), .B(men_men_n166_), .C(men_men_n86_), .Y(men_men_n468_));
  AOI210     u0446(.A0(men_men_n468_), .A1(men_men_n467_), .B0(men_men_n341_), .Y(men_men_n469_));
  NA2        u0447(.A(men_men_n198_), .B(i_10_), .Y(men_men_n470_));
  NA3        u0448(.A(men_men_n268_), .B(men_men_n64_), .C(i_2_), .Y(men_men_n471_));
  NA2        u0449(.A(men_men_n312_), .B(men_men_n244_), .Y(men_men_n472_));
  OAI220     u0450(.A0(men_men_n472_), .A1(men_men_n187_), .B0(men_men_n471_), .B1(men_men_n470_), .Y(men_men_n473_));
  NO2        u0451(.A(i_3_), .B(men_men_n48_), .Y(men_men_n474_));
  NA3        u0452(.A(men_men_n356_), .B(men_men_n355_), .C(men_men_n474_), .Y(men_men_n475_));
  NA2        u0453(.A(men_men_n333_), .B(men_men_n338_), .Y(men_men_n476_));
  OAI210     u0454(.A0(men_men_n476_), .A1(men_men_n194_), .B0(men_men_n475_), .Y(men_men_n477_));
  NO3        u0455(.A(men_men_n477_), .B(men_men_n473_), .C(men_men_n469_), .Y(men_men_n478_));
  AOI210     u0456(.A0(men_men_n478_), .A1(men_men_n466_), .B0(men_men_n285_), .Y(men_men_n479_));
  NO4        u0457(.A(men_men_n479_), .B(men_men_n459_), .C(men_men_n438_), .D(men_men_n409_), .Y(men_men_n480_));
  NO2        u0458(.A(men_men_n63_), .B(i_4_), .Y(men_men_n481_));
  NO2        u0459(.A(i_10_), .B(i_9_), .Y(men_men_n482_));
  NAi21      u0460(.An(i_12_), .B(i_8_), .Y(men_men_n483_));
  NO2        u0461(.A(men_men_n483_), .B(i_3_), .Y(men_men_n484_));
  NO2        u0462(.A(men_men_n46_), .B(i_4_), .Y(men_men_n485_));
  NA2        u0463(.A(men_men_n485_), .B(men_men_n106_), .Y(men_men_n486_));
  NO2        u0464(.A(men_men_n486_), .B(men_men_n210_), .Y(men_men_n487_));
  NA2        u0465(.A(men_men_n326_), .B(i_0_), .Y(men_men_n488_));
  NO3        u0466(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n280_), .B(men_men_n99_), .Y(men_men_n490_));
  NA2        u0468(.A(men_men_n490_), .B(men_men_n489_), .Y(men_men_n491_));
  NA2        u0469(.A(i_8_), .B(i_9_), .Y(men_men_n492_));
  AOI210     u0470(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n493_));
  OR2        u0471(.A(men_men_n493_), .B(men_men_n492_), .Y(men_men_n494_));
  NA2        u0472(.A(men_men_n298_), .B(men_men_n211_), .Y(men_men_n495_));
  OAI220     u0473(.A0(men_men_n495_), .A1(men_men_n494_), .B0(men_men_n491_), .B1(men_men_n488_), .Y(men_men_n496_));
  NA2        u0474(.A(men_men_n261_), .B(men_men_n325_), .Y(men_men_n497_));
  NO3        u0475(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n498_));
  INV        u0476(.A(men_men_n498_), .Y(men_men_n499_));
  NA3        u0477(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n500_));
  NA4        u0478(.A(men_men_n147_), .B(men_men_n118_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n501_));
  OAI220     u0479(.A0(men_men_n501_), .A1(men_men_n500_), .B0(men_men_n499_), .B1(men_men_n497_), .Y(men_men_n502_));
  NO3        u0480(.A(men_men_n502_), .B(men_men_n496_), .C(men_men_n487_), .Y(men_men_n503_));
  NA2        u0481(.A(men_men_n311_), .B(men_men_n110_), .Y(men_men_n504_));
  OR2        u0482(.A(men_men_n504_), .B(men_men_n214_), .Y(men_men_n505_));
  OA210      u0483(.A0(men_men_n375_), .A1(men_men_n103_), .B0(men_men_n313_), .Y(men_men_n506_));
  OA220      u0484(.A0(men_men_n506_), .A1(men_men_n165_), .B0(men_men_n505_), .B1(men_men_n241_), .Y(men_men_n507_));
  NA2        u0485(.A(men_men_n98_), .B(i_13_), .Y(men_men_n508_));
  NA2        u0486(.A(men_men_n463_), .B(men_men_n410_), .Y(men_men_n509_));
  NO2        u0487(.A(i_2_), .B(i_13_), .Y(men_men_n510_));
  NA3        u0488(.A(men_men_n510_), .B(men_men_n164_), .C(men_men_n101_), .Y(men_men_n511_));
  OAI220     u0489(.A0(men_men_n511_), .A1(men_men_n246_), .B0(men_men_n509_), .B1(men_men_n508_), .Y(men_men_n512_));
  NO3        u0490(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n513_));
  NO2        u0491(.A(i_6_), .B(i_7_), .Y(men_men_n514_));
  NA2        u0492(.A(men_men_n514_), .B(men_men_n513_), .Y(men_men_n515_));
  NO2        u0493(.A(i_11_), .B(i_1_), .Y(men_men_n516_));
  NO2        u0494(.A(men_men_n73_), .B(i_3_), .Y(men_men_n517_));
  OR2        u0495(.A(i_11_), .B(i_8_), .Y(men_men_n518_));
  NOi21      u0496(.An(i_2_), .B(i_7_), .Y(men_men_n519_));
  NAi31      u0497(.An(men_men_n518_), .B(men_men_n519_), .C(men_men_n517_), .Y(men_men_n520_));
  NO2        u0498(.A(men_men_n450_), .B(i_6_), .Y(men_men_n521_));
  NA3        u0499(.A(men_men_n521_), .B(men_men_n481_), .C(men_men_n75_), .Y(men_men_n522_));
  NO2        u0500(.A(men_men_n522_), .B(men_men_n520_), .Y(men_men_n523_));
  NO2        u0501(.A(i_3_), .B(men_men_n198_), .Y(men_men_n524_));
  NO2        u0502(.A(i_6_), .B(i_10_), .Y(men_men_n525_));
  NA4        u0503(.A(men_men_n525_), .B(men_men_n330_), .C(men_men_n524_), .D(men_men_n246_), .Y(men_men_n526_));
  NO2        u0504(.A(men_men_n526_), .B(men_men_n158_), .Y(men_men_n527_));
  NA3        u0505(.A(men_men_n255_), .B(men_men_n175_), .C(men_men_n135_), .Y(men_men_n528_));
  NA2        u0506(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n529_));
  NO2        u0507(.A(men_men_n160_), .B(i_3_), .Y(men_men_n530_));
  NAi31      u0508(.An(men_men_n529_), .B(men_men_n530_), .C(men_men_n235_), .Y(men_men_n531_));
  NA3        u0509(.A(men_men_n423_), .B(men_men_n183_), .C(men_men_n151_), .Y(men_men_n532_));
  NA3        u0510(.A(men_men_n532_), .B(men_men_n531_), .C(men_men_n528_), .Y(men_men_n533_));
  NO4        u0511(.A(men_men_n533_), .B(men_men_n527_), .C(men_men_n523_), .D(men_men_n512_), .Y(men_men_n534_));
  NA2        u0512(.A(men_men_n489_), .B(men_men_n411_), .Y(men_men_n535_));
  NA2        u0513(.A(men_men_n498_), .B(men_men_n418_), .Y(men_men_n536_));
  NO2        u0514(.A(men_men_n536_), .B(men_men_n233_), .Y(men_men_n537_));
  NAi21      u0515(.An(men_men_n224_), .B(men_men_n429_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n356_), .B(men_men_n226_), .Y(men_men_n539_));
  NO2        u0517(.A(men_men_n26_), .B(i_5_), .Y(men_men_n540_));
  NO2        u0518(.A(i_0_), .B(men_men_n86_), .Y(men_men_n541_));
  NA3        u0519(.A(men_men_n541_), .B(men_men_n540_), .C(men_men_n144_), .Y(men_men_n542_));
  OR3        u0520(.A(men_men_n319_), .B(men_men_n38_), .C(men_men_n46_), .Y(men_men_n543_));
  OAI220     u0521(.A0(men_men_n543_), .A1(men_men_n542_), .B0(men_men_n539_), .B1(men_men_n538_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n27_), .B(i_10_), .Y(men_men_n545_));
  NA2        u0523(.A(men_men_n330_), .B(men_men_n248_), .Y(men_men_n546_));
  OAI220     u0524(.A0(men_men_n546_), .A1(men_men_n471_), .B0(men_men_n545_), .B1(men_men_n508_), .Y(men_men_n547_));
  NA4        u0525(.A(men_men_n323_), .B(men_men_n232_), .C(men_men_n73_), .D(men_men_n246_), .Y(men_men_n548_));
  NO2        u0526(.A(men_men_n548_), .B(men_men_n515_), .Y(men_men_n549_));
  NO4        u0527(.A(men_men_n549_), .B(men_men_n547_), .C(men_men_n544_), .D(men_men_n537_), .Y(men_men_n550_));
  NA4        u0528(.A(men_men_n550_), .B(men_men_n534_), .C(men_men_n507_), .D(men_men_n503_), .Y(men_men_n551_));
  NA3        u0529(.A(men_men_n323_), .B(men_men_n180_), .C(men_men_n178_), .Y(men_men_n552_));
  OAI210     u0530(.A0(men_men_n317_), .A1(men_men_n185_), .B0(men_men_n552_), .Y(men_men_n553_));
  AN2        u0531(.A(men_men_n302_), .B(men_men_n243_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n554_), .B(men_men_n553_), .Y(men_men_n555_));
  NA2        u0533(.A(men_men_n125_), .B(men_men_n114_), .Y(men_men_n556_));
  AO220      u0534(.A0(men_men_n556_), .A1(men_men_n489_), .B0(men_men_n451_), .B1(i_6_), .Y(men_men_n557_));
  NA2        u0535(.A(men_men_n330_), .B(men_men_n167_), .Y(men_men_n558_));
  OAI210     u0536(.A0(men_men_n558_), .A1(men_men_n241_), .B0(men_men_n324_), .Y(men_men_n559_));
  AOI220     u0537(.A0(men_men_n559_), .A1(men_men_n342_), .B0(men_men_n557_), .B1(men_men_n326_), .Y(men_men_n560_));
  NA2        u0538(.A(men_men_n411_), .B(men_men_n234_), .Y(men_men_n561_));
  NA2        u0539(.A(men_men_n380_), .B(men_men_n73_), .Y(men_men_n562_));
  NA2        u0540(.A(men_men_n398_), .B(men_men_n390_), .Y(men_men_n563_));
  AO210      u0541(.A0(men_men_n562_), .A1(men_men_n561_), .B0(men_men_n563_), .Y(men_men_n564_));
  NO2        u0542(.A(men_men_n36_), .B(i_8_), .Y(men_men_n565_));
  INV        u0543(.A(men_men_n451_), .Y(men_men_n566_));
  NA2        u0544(.A(men_men_n566_), .B(men_men_n564_), .Y(men_men_n567_));
  INV        u0545(.A(men_men_n567_), .Y(men_men_n568_));
  NA2        u0546(.A(men_men_n268_), .B(men_men_n64_), .Y(men_men_n569_));
  OAI210     u0547(.A0(i_8_), .A1(men_men_n569_), .B0(men_men_n137_), .Y(men_men_n570_));
  AOI210     u0548(.A0(men_men_n199_), .A1(i_9_), .B0(men_men_n279_), .Y(men_men_n571_));
  NO2        u0549(.A(men_men_n571_), .B(men_men_n204_), .Y(men_men_n572_));
  OR2        u0550(.A(men_men_n187_), .B(i_4_), .Y(men_men_n573_));
  NO2        u0551(.A(men_men_n573_), .B(men_men_n86_), .Y(men_men_n574_));
  AOI220     u0552(.A0(men_men_n574_), .A1(men_men_n572_), .B0(men_men_n570_), .B1(men_men_n452_), .Y(men_men_n575_));
  NA4        u0553(.A(men_men_n575_), .B(men_men_n568_), .C(men_men_n560_), .D(men_men_n555_), .Y(men_men_n576_));
  NA2        u0554(.A(men_men_n417_), .B(men_men_n311_), .Y(men_men_n577_));
  OAI210     u0555(.A0(men_men_n413_), .A1(men_men_n172_), .B0(men_men_n577_), .Y(men_men_n578_));
  NO2        u0556(.A(i_12_), .B(men_men_n198_), .Y(men_men_n579_));
  NA2        u0557(.A(men_men_n579_), .B(men_men_n234_), .Y(men_men_n580_));
  NA3        u0558(.A(men_men_n525_), .B(men_men_n178_), .C(men_men_n27_), .Y(men_men_n581_));
  NO3        u0559(.A(men_men_n581_), .B(men_men_n580_), .C(men_men_n504_), .Y(men_men_n582_));
  NOi31      u0560(.An(men_men_n333_), .B(men_men_n450_), .C(men_men_n38_), .Y(men_men_n583_));
  OAI210     u0561(.A0(men_men_n583_), .A1(men_men_n582_), .B0(men_men_n578_), .Y(men_men_n584_));
  NO2        u0562(.A(i_8_), .B(i_7_), .Y(men_men_n585_));
  OAI210     u0563(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n586_));
  NA2        u0564(.A(men_men_n586_), .B(men_men_n232_), .Y(men_men_n587_));
  AOI220     u0565(.A0(men_men_n343_), .A1(men_men_n39_), .B0(men_men_n244_), .B1(men_men_n213_), .Y(men_men_n588_));
  OAI220     u0566(.A0(men_men_n588_), .A1(men_men_n573_), .B0(men_men_n587_), .B1(men_men_n252_), .Y(men_men_n589_));
  NA2        u0567(.A(men_men_n44_), .B(i_10_), .Y(men_men_n590_));
  NO2        u0568(.A(men_men_n590_), .B(i_6_), .Y(men_men_n591_));
  NA3        u0569(.A(men_men_n591_), .B(men_men_n589_), .C(men_men_n585_), .Y(men_men_n592_));
  AOI220     u0570(.A0(men_men_n463_), .A1(men_men_n343_), .B0(men_men_n257_), .B1(men_men_n254_), .Y(men_men_n593_));
  OAI220     u0571(.A0(men_men_n593_), .A1(men_men_n276_), .B0(men_men_n508_), .B1(men_men_n136_), .Y(men_men_n594_));
  NA2        u0572(.A(men_men_n594_), .B(men_men_n279_), .Y(men_men_n595_));
  NOi31      u0573(.An(men_men_n306_), .B(men_men_n317_), .C(men_men_n185_), .Y(men_men_n596_));
  NA3        u0574(.A(men_men_n323_), .B(men_men_n178_), .C(men_men_n98_), .Y(men_men_n597_));
  NO2        u0575(.A(men_men_n230_), .B(men_men_n44_), .Y(men_men_n598_));
  NO2        u0576(.A(men_men_n160_), .B(i_5_), .Y(men_men_n599_));
  NA3        u0577(.A(men_men_n599_), .B(men_men_n439_), .C(men_men_n336_), .Y(men_men_n600_));
  OAI210     u0578(.A0(men_men_n600_), .A1(men_men_n598_), .B0(men_men_n597_), .Y(men_men_n601_));
  OAI210     u0579(.A0(men_men_n601_), .A1(men_men_n596_), .B0(men_men_n498_), .Y(men_men_n602_));
  NA4        u0580(.A(men_men_n602_), .B(men_men_n595_), .C(men_men_n592_), .D(men_men_n584_), .Y(men_men_n603_));
  NA3        u0581(.A(men_men_n226_), .B(men_men_n71_), .C(men_men_n44_), .Y(men_men_n604_));
  NA2        u0582(.A(men_men_n298_), .B(men_men_n84_), .Y(men_men_n605_));
  AOI210     u0583(.A0(men_men_n604_), .A1(men_men_n370_), .B0(men_men_n605_), .Y(men_men_n606_));
  NA2        u0584(.A(men_men_n312_), .B(men_men_n302_), .Y(men_men_n607_));
  NO2        u0585(.A(men_men_n607_), .B(men_men_n177_), .Y(men_men_n608_));
  NA2        u0586(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n609_));
  NA2        u0587(.A(men_men_n482_), .B(men_men_n230_), .Y(men_men_n610_));
  NO2        u0588(.A(men_men_n609_), .B(men_men_n610_), .Y(men_men_n611_));
  AOI210     u0589(.A0(men_men_n391_), .A1(men_men_n46_), .B0(men_men_n395_), .Y(men_men_n612_));
  NA2        u0590(.A(i_0_), .B(men_men_n48_), .Y(men_men_n613_));
  NA3        u0591(.A(men_men_n579_), .B(men_men_n289_), .C(men_men_n613_), .Y(men_men_n614_));
  NO2        u0592(.A(men_men_n612_), .B(men_men_n614_), .Y(men_men_n615_));
  NO4        u0593(.A(men_men_n615_), .B(men_men_n611_), .C(men_men_n608_), .D(men_men_n606_), .Y(men_men_n616_));
  NO4        u0594(.A(men_men_n262_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n617_));
  NO3        u0595(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n618_));
  NO2        u0596(.A(men_men_n242_), .B(men_men_n36_), .Y(men_men_n619_));
  AN2        u0597(.A(men_men_n619_), .B(men_men_n618_), .Y(men_men_n620_));
  OA210      u0598(.A0(men_men_n620_), .A1(men_men_n617_), .B0(men_men_n380_), .Y(men_men_n621_));
  NO2        u0599(.A(men_men_n450_), .B(i_1_), .Y(men_men_n622_));
  NOi31      u0600(.An(men_men_n622_), .B(men_men_n490_), .C(men_men_n73_), .Y(men_men_n623_));
  AN4        u0601(.A(men_men_n623_), .B(men_men_n447_), .C(men_men_n540_), .D(i_2_), .Y(men_men_n624_));
  NO2        u0602(.A(men_men_n461_), .B(men_men_n181_), .Y(men_men_n625_));
  NO3        u0603(.A(men_men_n625_), .B(men_men_n624_), .C(men_men_n621_), .Y(men_men_n626_));
  NOi21      u0604(.An(i_10_), .B(i_6_), .Y(men_men_n627_));
  NO2        u0605(.A(men_men_n86_), .B(men_men_n25_), .Y(men_men_n628_));
  AOI220     u0606(.A0(men_men_n298_), .A1(men_men_n628_), .B0(men_men_n289_), .B1(men_men_n627_), .Y(men_men_n629_));
  NO2        u0607(.A(men_men_n629_), .B(men_men_n488_), .Y(men_men_n630_));
  NO2        u0608(.A(men_men_n117_), .B(men_men_n23_), .Y(men_men_n631_));
  NA2        u0609(.A(men_men_n333_), .B(men_men_n167_), .Y(men_men_n632_));
  AOI220     u0610(.A0(men_men_n632_), .A1(men_men_n472_), .B0(men_men_n188_), .B1(men_men_n186_), .Y(men_men_n633_));
  NO2        u0611(.A(men_men_n203_), .B(men_men_n37_), .Y(men_men_n634_));
  NOi31      u0612(.An(men_men_n148_), .B(men_men_n634_), .C(men_men_n351_), .Y(men_men_n635_));
  NO3        u0613(.A(men_men_n635_), .B(men_men_n633_), .C(men_men_n630_), .Y(men_men_n636_));
  NO2        u0614(.A(men_men_n562_), .B(men_men_n406_), .Y(men_men_n637_));
  INV        u0615(.A(men_men_n336_), .Y(men_men_n638_));
  NO2        u0616(.A(i_12_), .B(men_men_n86_), .Y(men_men_n639_));
  NA3        u0617(.A(men_men_n639_), .B(men_men_n289_), .C(men_men_n613_), .Y(men_men_n640_));
  NA3        u0618(.A(men_men_n414_), .B(men_men_n298_), .C(men_men_n226_), .Y(men_men_n641_));
  AOI210     u0619(.A0(men_men_n641_), .A1(men_men_n640_), .B0(men_men_n638_), .Y(men_men_n642_));
  NA2        u0620(.A(men_men_n178_), .B(i_0_), .Y(men_men_n643_));
  NO3        u0621(.A(men_men_n643_), .B(men_men_n362_), .C(men_men_n317_), .Y(men_men_n644_));
  OR2        u0622(.A(i_2_), .B(i_5_), .Y(men_men_n645_));
  OR2        u0623(.A(men_men_n645_), .B(men_men_n442_), .Y(men_men_n646_));
  AOI210     u0624(.A0(men_men_n400_), .A1(men_men_n254_), .B0(men_men_n203_), .Y(men_men_n647_));
  AOI210     u0625(.A0(men_men_n647_), .A1(men_men_n646_), .B0(men_men_n538_), .Y(men_men_n648_));
  NO4        u0626(.A(men_men_n648_), .B(men_men_n644_), .C(men_men_n642_), .D(men_men_n637_), .Y(men_men_n649_));
  NA4        u0627(.A(men_men_n649_), .B(men_men_n636_), .C(men_men_n626_), .D(men_men_n616_), .Y(men_men_n650_));
  NO4        u0628(.A(men_men_n650_), .B(men_men_n603_), .C(men_men_n576_), .D(men_men_n551_), .Y(men_men_n651_));
  NA4        u0629(.A(men_men_n651_), .B(men_men_n480_), .C(men_men_n379_), .D(men_men_n329_), .Y(men7));
  NO2        u0630(.A(men_men_n94_), .B(men_men_n54_), .Y(men_men_n653_));
  NO2        u0631(.A(men_men_n110_), .B(men_men_n91_), .Y(men_men_n654_));
  NA2        u0632(.A(men_men_n412_), .B(men_men_n654_), .Y(men_men_n655_));
  NA2        u0633(.A(men_men_n525_), .B(men_men_n84_), .Y(men_men_n656_));
  NA2        u0634(.A(i_11_), .B(men_men_n198_), .Y(men_men_n657_));
  NA2        u0635(.A(men_men_n146_), .B(men_men_n657_), .Y(men_men_n658_));
  OAI210     u0636(.A0(men_men_n658_), .A1(men_men_n656_), .B0(men_men_n655_), .Y(men_men_n659_));
  NA3        u0637(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n660_));
  NO2        u0638(.A(men_men_n246_), .B(i_4_), .Y(men_men_n661_));
  NA2        u0639(.A(men_men_n661_), .B(i_8_), .Y(men_men_n662_));
  AOI210     u0640(.A0(men_men_n662_), .A1(men_men_n107_), .B0(men_men_n660_), .Y(men_men_n663_));
  NA2        u0641(.A(i_2_), .B(men_men_n86_), .Y(men_men_n664_));
  OAI210     u0642(.A0(men_men_n89_), .A1(men_men_n208_), .B0(men_men_n209_), .Y(men_men_n665_));
  NO2        u0643(.A(i_7_), .B(men_men_n37_), .Y(men_men_n666_));
  NA2        u0644(.A(i_4_), .B(i_8_), .Y(men_men_n667_));
  AOI210     u0645(.A0(men_men_n667_), .A1(men_men_n323_), .B0(men_men_n666_), .Y(men_men_n668_));
  OAI220     u0646(.A0(men_men_n668_), .A1(men_men_n664_), .B0(men_men_n665_), .B1(i_13_), .Y(men_men_n669_));
  NO4        u0647(.A(men_men_n669_), .B(men_men_n663_), .C(men_men_n659_), .D(men_men_n653_), .Y(men_men_n670_));
  AOI210     u0648(.A0(men_men_n131_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n671_));
  AOI210     u0649(.A0(men_men_n671_), .A1(men_men_n246_), .B0(men_men_n164_), .Y(men_men_n672_));
  OR2        u0650(.A(i_6_), .B(i_10_), .Y(men_men_n673_));
  NO2        u0651(.A(men_men_n673_), .B(men_men_n23_), .Y(men_men_n674_));
  OR3        u0652(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n675_));
  NO3        u0653(.A(men_men_n675_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n676_));
  INV        u0654(.A(men_men_n205_), .Y(men_men_n677_));
  NO2        u0655(.A(men_men_n676_), .B(men_men_n674_), .Y(men_men_n678_));
  OA220      u0656(.A0(men_men_n678_), .A1(men_men_n638_), .B0(men_men_n672_), .B1(men_men_n281_), .Y(men_men_n679_));
  AOI210     u0657(.A0(men_men_n679_), .A1(men_men_n670_), .B0(men_men_n63_), .Y(men_men_n680_));
  NOi21      u0658(.An(i_11_), .B(i_7_), .Y(men_men_n681_));
  AO210      u0659(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n682_));
  NO2        u0660(.A(men_men_n682_), .B(men_men_n681_), .Y(men_men_n683_));
  NA2        u0661(.A(men_men_n683_), .B(men_men_n213_), .Y(men_men_n684_));
  NA3        u0662(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n685_));
  NAi31      u0663(.An(men_men_n685_), .B(men_men_n223_), .C(i_11_), .Y(men_men_n686_));
  AOI210     u0664(.A0(men_men_n686_), .A1(men_men_n684_), .B0(men_men_n63_), .Y(men_men_n687_));
  NA2        u0665(.A(men_men_n88_), .B(men_men_n63_), .Y(men_men_n688_));
  AO210      u0666(.A0(men_men_n688_), .A1(men_men_n406_), .B0(men_men_n40_), .Y(men_men_n689_));
  NO3        u0667(.A(men_men_n270_), .B(men_men_n215_), .C(men_men_n657_), .Y(men_men_n690_));
  NA2        u0668(.A(men_men_n690_), .B(men_men_n63_), .Y(men_men_n691_));
  NA2        u0669(.A(men_men_n443_), .B(men_men_n31_), .Y(men_men_n692_));
  OR2        u0670(.A(men_men_n215_), .B(men_men_n110_), .Y(men_men_n693_));
  NA2        u0671(.A(men_men_n693_), .B(men_men_n692_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n63_), .B(i_9_), .Y(men_men_n695_));
  NO2        u0673(.A(men_men_n695_), .B(i_4_), .Y(men_men_n696_));
  NA2        u0674(.A(men_men_n696_), .B(men_men_n694_), .Y(men_men_n697_));
  NO2        u0675(.A(i_1_), .B(i_12_), .Y(men_men_n698_));
  NA3        u0676(.A(men_men_n698_), .B(men_men_n112_), .C(men_men_n24_), .Y(men_men_n699_));
  NA4        u0677(.A(men_men_n699_), .B(men_men_n697_), .C(men_men_n691_), .D(men_men_n689_), .Y(men_men_n700_));
  OAI210     u0678(.A0(men_men_n700_), .A1(men_men_n687_), .B0(i_6_), .Y(men_men_n701_));
  OAI210     u0679(.A0(men_men_n685_), .A1(men_men_n110_), .B0(men_men_n500_), .Y(men_men_n702_));
  NA2        u0680(.A(men_men_n702_), .B(men_men_n639_), .Y(men_men_n703_));
  NO2        u0681(.A(men_men_n246_), .B(men_men_n86_), .Y(men_men_n704_));
  NA2        u0682(.A(men_men_n703_), .B(men_men_n491_), .Y(men_men_n705_));
  NO4        u0683(.A(men_men_n223_), .B(men_men_n131_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n706_));
  NA2        u0684(.A(men_men_n706_), .B(men_men_n695_), .Y(men_men_n707_));
  NA2        u0685(.A(men_men_n246_), .B(i_6_), .Y(men_men_n708_));
  NO3        u0686(.A(men_men_n673_), .B(men_men_n242_), .C(men_men_n23_), .Y(men_men_n709_));
  AOI210     u0687(.A0(i_1_), .A1(men_men_n271_), .B0(men_men_n709_), .Y(men_men_n710_));
  OAI210     u0688(.A0(men_men_n710_), .A1(men_men_n44_), .B0(men_men_n707_), .Y(men_men_n711_));
  NA3        u0689(.A(men_men_n585_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n712_));
  NA3        u0690(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n713_));
  NO2        u0691(.A(men_men_n46_), .B(i_1_), .Y(men_men_n714_));
  NA3        u0692(.A(men_men_n714_), .B(men_men_n280_), .C(men_men_n44_), .Y(men_men_n715_));
  NO2        u0693(.A(men_men_n715_), .B(men_men_n713_), .Y(men_men_n716_));
  NA3        u0694(.A(men_men_n695_), .B(men_men_n336_), .C(i_6_), .Y(men_men_n717_));
  NO2        u0695(.A(men_men_n717_), .B(men_men_n23_), .Y(men_men_n718_));
  NAi21      u0696(.An(men_men_n712_), .B(men_men_n93_), .Y(men_men_n719_));
  NA2        u0697(.A(men_men_n714_), .B(men_men_n280_), .Y(men_men_n720_));
  NO2        u0698(.A(i_11_), .B(men_men_n37_), .Y(men_men_n721_));
  NA2        u0699(.A(men_men_n721_), .B(men_men_n24_), .Y(men_men_n722_));
  OAI210     u0700(.A0(men_men_n722_), .A1(men_men_n720_), .B0(men_men_n719_), .Y(men_men_n723_));
  OR3        u0701(.A(men_men_n723_), .B(men_men_n718_), .C(men_men_n716_), .Y(men_men_n724_));
  NO3        u0702(.A(men_men_n724_), .B(men_men_n711_), .C(men_men_n705_), .Y(men_men_n725_));
  NO2        u0703(.A(men_men_n246_), .B(men_men_n103_), .Y(men_men_n726_));
  NO2        u0704(.A(men_men_n726_), .B(men_men_n681_), .Y(men_men_n727_));
  NA2        u0705(.A(men_men_n727_), .B(i_1_), .Y(men_men_n728_));
  NO2        u0706(.A(men_men_n728_), .B(men_men_n675_), .Y(men_men_n729_));
  NO2        u0707(.A(men_men_n449_), .B(men_men_n86_), .Y(men_men_n730_));
  NA2        u0708(.A(men_men_n729_), .B(men_men_n46_), .Y(men_men_n731_));
  NA2        u0709(.A(i_3_), .B(men_men_n198_), .Y(men_men_n732_));
  NO2        u0710(.A(men_men_n732_), .B(men_men_n117_), .Y(men_men_n733_));
  AN2        u0711(.A(men_men_n733_), .B(men_men_n591_), .Y(men_men_n734_));
  NO2        u0712(.A(men_men_n242_), .B(men_men_n44_), .Y(men_men_n735_));
  NO3        u0713(.A(men_men_n735_), .B(men_men_n326_), .C(men_men_n247_), .Y(men_men_n736_));
  NO2        u0714(.A(men_men_n120_), .B(men_men_n37_), .Y(men_men_n737_));
  NO2        u0715(.A(men_men_n737_), .B(i_6_), .Y(men_men_n738_));
  NO2        u0716(.A(men_men_n86_), .B(i_9_), .Y(men_men_n739_));
  NO2        u0717(.A(men_men_n739_), .B(men_men_n63_), .Y(men_men_n740_));
  NO2        u0718(.A(men_men_n740_), .B(men_men_n698_), .Y(men_men_n741_));
  NO4        u0719(.A(men_men_n741_), .B(men_men_n738_), .C(men_men_n736_), .D(i_4_), .Y(men_men_n742_));
  NA2        u0720(.A(i_1_), .B(i_3_), .Y(men_men_n743_));
  NO2        u0721(.A(men_men_n492_), .B(men_men_n94_), .Y(men_men_n744_));
  AOI210     u0722(.A0(men_men_n735_), .A1(men_men_n627_), .B0(men_men_n744_), .Y(men_men_n745_));
  NO2        u0723(.A(men_men_n745_), .B(men_men_n743_), .Y(men_men_n746_));
  NO3        u0724(.A(men_men_n746_), .B(men_men_n742_), .C(men_men_n734_), .Y(men_men_n747_));
  NA4        u0725(.A(men_men_n747_), .B(men_men_n731_), .C(men_men_n725_), .D(men_men_n701_), .Y(men_men_n748_));
  NO3        u0726(.A(men_men_n518_), .B(i_3_), .C(i_7_), .Y(men_men_n749_));
  NOi21      u0727(.An(men_men_n749_), .B(i_10_), .Y(men_men_n750_));
  OA210      u0728(.A0(men_men_n750_), .A1(men_men_n255_), .B0(men_men_n86_), .Y(men_men_n751_));
  NA2        u0729(.A(men_men_n398_), .B(men_men_n397_), .Y(men_men_n752_));
  NA3        u0730(.A(men_men_n525_), .B(men_men_n565_), .C(men_men_n46_), .Y(men_men_n753_));
  NO3        u0731(.A(men_men_n519_), .B(men_men_n667_), .C(men_men_n86_), .Y(men_men_n754_));
  NA2        u0732(.A(men_men_n754_), .B(men_men_n25_), .Y(men_men_n755_));
  NA3        u0733(.A(men_men_n164_), .B(men_men_n84_), .C(men_men_n86_), .Y(men_men_n756_));
  NA4        u0734(.A(men_men_n756_), .B(men_men_n755_), .C(men_men_n753_), .D(men_men_n752_), .Y(men_men_n757_));
  OAI210     u0735(.A0(men_men_n757_), .A1(men_men_n751_), .B0(i_1_), .Y(men_men_n758_));
  AOI210     u0736(.A0(men_men_n280_), .A1(men_men_n99_), .B0(i_1_), .Y(men_men_n759_));
  NO2        u0737(.A(men_men_n396_), .B(i_2_), .Y(men_men_n760_));
  NA2        u0738(.A(men_men_n760_), .B(men_men_n759_), .Y(men_men_n761_));
  OAI210     u0739(.A0(men_men_n717_), .A1(men_men_n483_), .B0(men_men_n761_), .Y(men_men_n762_));
  INV        u0740(.A(men_men_n762_), .Y(men_men_n763_));
  NA2        u0741(.A(men_men_n763_), .B(men_men_n758_), .Y(men_men_n764_));
  OR2        u0742(.A(i_11_), .B(i_7_), .Y(men_men_n765_));
  NA3        u0743(.A(men_men_n765_), .B(men_men_n108_), .C(men_men_n141_), .Y(men_men_n766_));
  AOI220     u0744(.A0(men_men_n510_), .A1(men_men_n164_), .B0(men_men_n485_), .B1(men_men_n141_), .Y(men_men_n767_));
  OAI210     u0745(.A0(men_men_n767_), .A1(men_men_n44_), .B0(men_men_n766_), .Y(men_men_n768_));
  AOI210     u0746(.A0(men_men_n713_), .A1(men_men_n54_), .B0(i_12_), .Y(men_men_n769_));
  NO2        u0747(.A(men_men_n519_), .B(men_men_n24_), .Y(men_men_n770_));
  AOI220     u0748(.A0(men_men_n770_), .A1(men_men_n730_), .B0(men_men_n255_), .B1(men_men_n134_), .Y(men_men_n771_));
  OAI220     u0749(.A0(men_men_n771_), .A1(men_men_n40_), .B0(men_men_n1146_), .B1(men_men_n94_), .Y(men_men_n772_));
  AOI210     u0750(.A0(men_men_n768_), .A1(men_men_n353_), .B0(men_men_n772_), .Y(men_men_n773_));
  NA2        u0751(.A(men_men_n117_), .B(men_men_n110_), .Y(men_men_n774_));
  AOI220     u0752(.A0(men_men_n774_), .A1(men_men_n72_), .B0(men_men_n414_), .B1(men_men_n714_), .Y(men_men_n775_));
  NO2        u0753(.A(men_men_n775_), .B(men_men_n252_), .Y(men_men_n776_));
  AOI210     u0754(.A0(men_men_n483_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n777_));
  NOi31      u0755(.An(men_men_n777_), .B(men_men_n656_), .C(men_men_n44_), .Y(men_men_n778_));
  NO2        u0756(.A(men_men_n713_), .B(men_men_n117_), .Y(men_men_n779_));
  INV        u0757(.A(men_men_n779_), .Y(men_men_n780_));
  NO2        u0758(.A(men_men_n780_), .B(men_men_n71_), .Y(men_men_n781_));
  NO3        u0759(.A(men_men_n71_), .B(men_men_n32_), .C(men_men_n103_), .Y(men_men_n782_));
  NA2        u0760(.A(men_men_n26_), .B(men_men_n198_), .Y(men_men_n783_));
  NA2        u0761(.A(men_men_n783_), .B(i_7_), .Y(men_men_n784_));
  NO3        u0762(.A(men_men_n519_), .B(men_men_n246_), .C(men_men_n86_), .Y(men_men_n785_));
  AOI210     u0763(.A0(men_men_n785_), .A1(men_men_n784_), .B0(men_men_n782_), .Y(men_men_n786_));
  AOI220     u0764(.A0(men_men_n414_), .A1(men_men_n714_), .B0(men_men_n93_), .B1(men_men_n104_), .Y(men_men_n787_));
  OAI220     u0765(.A0(men_men_n787_), .A1(men_men_n662_), .B0(men_men_n786_), .B1(men_men_n677_), .Y(men_men_n788_));
  NO4        u0766(.A(men_men_n788_), .B(men_men_n781_), .C(men_men_n778_), .D(men_men_n776_), .Y(men_men_n789_));
  OR2        u0767(.A(i_11_), .B(i_6_), .Y(men_men_n790_));
  NA3        u0768(.A(men_men_n661_), .B(men_men_n783_), .C(i_7_), .Y(men_men_n791_));
  AOI210     u0769(.A0(men_men_n791_), .A1(men_men_n780_), .B0(men_men_n790_), .Y(men_men_n792_));
  NA3        u0770(.A(men_men_n443_), .B(men_men_n666_), .C(men_men_n99_), .Y(men_men_n793_));
  NA2        u0771(.A(men_men_n104_), .B(men_men_n783_), .Y(men_men_n794_));
  NAi21      u0772(.An(i_11_), .B(i_12_), .Y(men_men_n795_));
  NOi41      u0773(.An(men_men_n113_), .B(men_men_n795_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n796_));
  NO3        u0774(.A(men_men_n519_), .B(men_men_n639_), .C(men_men_n667_), .Y(men_men_n797_));
  AOI220     u0775(.A0(men_men_n797_), .A1(men_men_n330_), .B0(men_men_n796_), .B1(men_men_n794_), .Y(men_men_n798_));
  NA2        u0776(.A(men_men_n798_), .B(men_men_n793_), .Y(men_men_n799_));
  OAI210     u0777(.A0(men_men_n799_), .A1(men_men_n792_), .B0(men_men_n63_), .Y(men_men_n800_));
  NO2        u0778(.A(i_2_), .B(i_12_), .Y(men_men_n801_));
  NA2        u0779(.A(men_men_n395_), .B(men_men_n801_), .Y(men_men_n802_));
  NA2        u0780(.A(i_8_), .B(men_men_n25_), .Y(men_men_n803_));
  NO3        u0781(.A(men_men_n803_), .B(men_men_n412_), .C(men_men_n661_), .Y(men_men_n804_));
  OAI210     u0782(.A0(men_men_n804_), .A1(men_men_n397_), .B0(men_men_n395_), .Y(men_men_n805_));
  NO2        u0783(.A(men_men_n131_), .B(i_2_), .Y(men_men_n806_));
  NA2        u0784(.A(men_men_n806_), .B(men_men_n698_), .Y(men_men_n807_));
  NA3        u0785(.A(men_men_n807_), .B(men_men_n805_), .C(men_men_n802_), .Y(men_men_n808_));
  NA2        u0786(.A(men_men_n808_), .B(men_men_n45_), .Y(men_men_n809_));
  NA4        u0787(.A(men_men_n809_), .B(men_men_n800_), .C(men_men_n789_), .D(men_men_n773_), .Y(men_men_n810_));
  OR4        u0788(.A(men_men_n810_), .B(men_men_n764_), .C(men_men_n748_), .D(men_men_n680_), .Y(men5));
  AOI210     u0789(.A0(men_men_n727_), .A1(men_men_n283_), .B0(men_men_n452_), .Y(men_men_n812_));
  NA3        u0790(.A(men_men_n24_), .B(men_men_n801_), .C(men_men_n110_), .Y(men_men_n813_));
  NA2        u0791(.A(men_men_n89_), .B(men_men_n661_), .Y(men_men_n814_));
  NA3        u0792(.A(men_men_n814_), .B(men_men_n813_), .C(men_men_n812_), .Y(men_men_n815_));
  NO3        u0793(.A(i_11_), .B(men_men_n246_), .C(i_13_), .Y(men_men_n816_));
  NO2        u0794(.A(men_men_n127_), .B(men_men_n23_), .Y(men_men_n817_));
  NA2        u0795(.A(i_12_), .B(i_8_), .Y(men_men_n818_));
  OAI210     u0796(.A0(men_men_n46_), .A1(i_3_), .B0(men_men_n818_), .Y(men_men_n819_));
  AOI220     u0797(.A0(men_men_n336_), .A1(men_men_n631_), .B0(men_men_n819_), .B1(men_men_n817_), .Y(men_men_n820_));
  INV        u0798(.A(men_men_n820_), .Y(men_men_n821_));
  NO2        u0799(.A(men_men_n821_), .B(men_men_n815_), .Y(men_men_n822_));
  INV        u0800(.A(men_men_n175_), .Y(men_men_n823_));
  INV        u0801(.A(men_men_n255_), .Y(men_men_n824_));
  OAI210     u0802(.A0(men_men_n760_), .A1(men_men_n484_), .B0(men_men_n113_), .Y(men_men_n825_));
  AOI210     u0803(.A0(men_men_n825_), .A1(men_men_n824_), .B0(men_men_n823_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n492_), .B(men_men_n26_), .Y(men_men_n827_));
  NO2        u0805(.A(men_men_n827_), .B(men_men_n454_), .Y(men_men_n828_));
  NA2        u0806(.A(men_men_n828_), .B(i_2_), .Y(men_men_n829_));
  INV        u0807(.A(men_men_n829_), .Y(men_men_n830_));
  AOI210     u0808(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n450_), .Y(men_men_n831_));
  AOI210     u0809(.A0(men_men_n831_), .A1(men_men_n830_), .B0(men_men_n826_), .Y(men_men_n832_));
  NO2        u0810(.A(men_men_n195_), .B(men_men_n128_), .Y(men_men_n833_));
  OAI210     u0811(.A0(men_men_n833_), .A1(men_men_n817_), .B0(i_2_), .Y(men_men_n834_));
  INV        u0812(.A(men_men_n176_), .Y(men_men_n835_));
  NO3        u0813(.A(men_men_n682_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n836_));
  AOI210     u0814(.A0(men_men_n835_), .A1(men_men_n89_), .B0(men_men_n836_), .Y(men_men_n837_));
  AOI210     u0815(.A0(men_men_n837_), .A1(men_men_n834_), .B0(men_men_n198_), .Y(men_men_n838_));
  NA2        u0816(.A(men_men_n205_), .B(men_men_n208_), .Y(men_men_n839_));
  NA2        u0817(.A(men_men_n154_), .B(men_men_n657_), .Y(men_men_n840_));
  AOI210     u0818(.A0(men_men_n840_), .A1(men_men_n839_), .B0(men_men_n400_), .Y(men_men_n841_));
  AOI210     u0819(.A0(men_men_n215_), .A1(men_men_n150_), .B0(men_men_n565_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n842_), .B(men_men_n454_), .Y(men_men_n843_));
  NA3        u0821(.A(men_men_n103_), .B(men_men_n323_), .C(men_men_n42_), .Y(men_men_n844_));
  OAI210     u0822(.A0(men_men_n844_), .A1(i_11_), .B0(men_men_n843_), .Y(men_men_n845_));
  NO3        u0823(.A(men_men_n845_), .B(men_men_n841_), .C(men_men_n838_), .Y(men_men_n846_));
  NA2        u0824(.A(men_men_n631_), .B(men_men_n28_), .Y(men_men_n847_));
  INV        u0825(.A(men_men_n290_), .Y(men_men_n848_));
  NA2        u0826(.A(men_men_n848_), .B(men_men_n847_), .Y(men_men_n849_));
  NO2        u0827(.A(men_men_n62_), .B(i_12_), .Y(men_men_n850_));
  INV        u0828(.A(men_men_n129_), .Y(men_men_n851_));
  NO2        u0829(.A(men_men_n851_), .B(men_men_n657_), .Y(men_men_n852_));
  AOI220     u0830(.A0(men_men_n852_), .A1(men_men_n36_), .B0(men_men_n849_), .B1(men_men_n46_), .Y(men_men_n853_));
  NA4        u0831(.A(men_men_n853_), .B(men_men_n846_), .C(men_men_n832_), .D(men_men_n822_), .Y(men6));
  NO2        u0832(.A(men_men_n325_), .B(i_1_), .Y(men_men_n855_));
  NO2        u0833(.A(men_men_n190_), .B(men_men_n142_), .Y(men_men_n856_));
  OAI210     u0834(.A0(men_men_n856_), .A1(men_men_n855_), .B0(men_men_n806_), .Y(men_men_n857_));
  NA4        u0835(.A(men_men_n418_), .B(men_men_n524_), .C(men_men_n71_), .D(men_men_n103_), .Y(men_men_n858_));
  INV        u0836(.A(men_men_n858_), .Y(men_men_n859_));
  NO2        u0837(.A(men_men_n229_), .B(men_men_n529_), .Y(men_men_n860_));
  NO2        u0838(.A(i_11_), .B(i_9_), .Y(men_men_n861_));
  AO210      u0839(.A0(men_men_n858_), .A1(men_men_n857_), .B0(i_12_), .Y(men_men_n862_));
  NA2        u0840(.A(men_men_n401_), .B(men_men_n356_), .Y(men_men_n863_));
  NA2        u0841(.A(men_men_n639_), .B(men_men_n63_), .Y(men_men_n864_));
  NA2        u0842(.A(men_men_n750_), .B(men_men_n71_), .Y(men_men_n865_));
  NA4        u0843(.A(men_men_n688_), .B(men_men_n865_), .C(men_men_n864_), .D(men_men_n863_), .Y(men_men_n866_));
  INV        u0844(.A(men_men_n202_), .Y(men_men_n867_));
  AOI220     u0845(.A0(men_men_n867_), .A1(men_men_n861_), .B0(men_men_n866_), .B1(men_men_n73_), .Y(men_men_n868_));
  INV        u0846(.A(men_men_n347_), .Y(men_men_n869_));
  NA2        u0847(.A(men_men_n75_), .B(men_men_n134_), .Y(men_men_n870_));
  INV        u0848(.A(men_men_n127_), .Y(men_men_n871_));
  NA2        u0849(.A(men_men_n871_), .B(men_men_n46_), .Y(men_men_n872_));
  AOI210     u0850(.A0(men_men_n872_), .A1(men_men_n870_), .B0(men_men_n869_), .Y(men_men_n873_));
  NO3        u0851(.A(men_men_n262_), .B(men_men_n135_), .C(i_9_), .Y(men_men_n874_));
  NA2        u0852(.A(men_men_n874_), .B(men_men_n850_), .Y(men_men_n875_));
  AOI210     u0853(.A0(men_men_n875_), .A1(men_men_n563_), .B0(men_men_n190_), .Y(men_men_n876_));
  NO2        u0854(.A(men_men_n32_), .B(i_11_), .Y(men_men_n877_));
  NA3        u0855(.A(men_men_n877_), .B(men_men_n514_), .C(men_men_n418_), .Y(men_men_n878_));
  NAi32      u0856(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n879_));
  AOI210     u0857(.A0(men_men_n790_), .A1(men_men_n87_), .B0(men_men_n879_), .Y(men_men_n880_));
  OAI210     u0858(.A0(men_men_n749_), .A1(men_men_n619_), .B0(men_men_n618_), .Y(men_men_n881_));
  NAi31      u0859(.An(men_men_n880_), .B(men_men_n881_), .C(men_men_n878_), .Y(men_men_n882_));
  OR3        u0860(.A(men_men_n882_), .B(men_men_n876_), .C(men_men_n873_), .Y(men_men_n883_));
  NO2        u0861(.A(men_men_n765_), .B(i_2_), .Y(men_men_n884_));
  NA2        u0862(.A(men_men_n48_), .B(men_men_n37_), .Y(men_men_n885_));
  OAI210     u0863(.A0(men_men_n885_), .A1(men_men_n442_), .B0(men_men_n385_), .Y(men_men_n886_));
  NA2        u0864(.A(men_men_n886_), .B(men_men_n884_), .Y(men_men_n887_));
  AO220      u0865(.A0(men_men_n384_), .A1(men_men_n374_), .B0(men_men_n426_), .B1(men_men_n657_), .Y(men_men_n888_));
  NA3        u0866(.A(men_men_n888_), .B(men_men_n267_), .C(i_7_), .Y(men_men_n889_));
  OR2        u0867(.A(men_men_n683_), .B(men_men_n484_), .Y(men_men_n890_));
  NA3        u0868(.A(men_men_n890_), .B(men_men_n149_), .C(men_men_n69_), .Y(men_men_n891_));
  OR2        u0869(.A(men_men_n536_), .B(men_men_n36_), .Y(men_men_n892_));
  NA4        u0870(.A(men_men_n892_), .B(men_men_n891_), .C(men_men_n889_), .D(men_men_n887_), .Y(men_men_n893_));
  OAI210     u0871(.A0(men_men_n704_), .A1(i_11_), .B0(men_men_n87_), .Y(men_men_n894_));
  AOI220     u0872(.A0(men_men_n894_), .A1(men_men_n618_), .B0(men_men_n860_), .B1(men_men_n784_), .Y(men_men_n895_));
  NA3        u0873(.A(men_men_n400_), .B(men_men_n248_), .C(men_men_n149_), .Y(men_men_n896_));
  NA2        u0874(.A(men_men_n426_), .B(men_men_n70_), .Y(men_men_n897_));
  NA4        u0875(.A(men_men_n897_), .B(men_men_n896_), .C(men_men_n895_), .D(men_men_n665_), .Y(men_men_n898_));
  AO210      u0876(.A0(men_men_n565_), .A1(men_men_n46_), .B0(men_men_n88_), .Y(men_men_n899_));
  NA2        u0877(.A(men_men_n899_), .B(men_men_n525_), .Y(men_men_n900_));
  AOI210     u0878(.A0(men_men_n484_), .A1(men_men_n482_), .B0(men_men_n617_), .Y(men_men_n901_));
  NO2        u0879(.A(men_men_n673_), .B(men_men_n104_), .Y(men_men_n902_));
  OAI210     u0880(.A0(men_men_n902_), .A1(men_men_n114_), .B0(men_men_n441_), .Y(men_men_n903_));
  NA2        u0881(.A(men_men_n254_), .B(men_men_n46_), .Y(men_men_n904_));
  INV        u0882(.A(men_men_n646_), .Y(men_men_n905_));
  NA3        u0883(.A(men_men_n905_), .B(men_men_n347_), .C(i_7_), .Y(men_men_n906_));
  NA4        u0884(.A(men_men_n906_), .B(men_men_n903_), .C(men_men_n901_), .D(men_men_n900_), .Y(men_men_n907_));
  NO4        u0885(.A(men_men_n907_), .B(men_men_n898_), .C(men_men_n893_), .D(men_men_n883_), .Y(men_men_n908_));
  NA4        u0886(.A(men_men_n908_), .B(men_men_n868_), .C(men_men_n862_), .D(men_men_n408_), .Y(men3));
  NA2        u0887(.A(i_12_), .B(i_10_), .Y(men_men_n910_));
  NA2        u0888(.A(i_6_), .B(i_7_), .Y(men_men_n911_));
  NO2        u0889(.A(men_men_n911_), .B(i_0_), .Y(men_men_n912_));
  NO2        u0890(.A(i_11_), .B(men_men_n246_), .Y(men_men_n913_));
  OAI210     u0891(.A0(men_men_n912_), .A1(men_men_n306_), .B0(men_men_n913_), .Y(men_men_n914_));
  NO2        u0892(.A(men_men_n914_), .B(men_men_n198_), .Y(men_men_n915_));
  NO3        u0893(.A(men_men_n488_), .B(men_men_n91_), .C(men_men_n44_), .Y(men_men_n916_));
  OA210      u0894(.A0(men_men_n916_), .A1(men_men_n915_), .B0(men_men_n178_), .Y(men_men_n917_));
  NA3        u0895(.A(men_men_n896_), .B(men_men_n665_), .C(men_men_n399_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n918_), .B(men_men_n39_), .Y(men_men_n919_));
  NOi21      u0897(.An(men_men_n98_), .B(men_men_n828_), .Y(men_men_n920_));
  NO3        u0898(.A(men_men_n693_), .B(men_men_n492_), .C(men_men_n134_), .Y(men_men_n921_));
  NA2        u0899(.A(men_men_n443_), .B(men_men_n45_), .Y(men_men_n922_));
  AN2        u0900(.A(men_men_n490_), .B(men_men_n55_), .Y(men_men_n923_));
  NO3        u0901(.A(men_men_n923_), .B(men_men_n921_), .C(men_men_n920_), .Y(men_men_n924_));
  AOI210     u0902(.A0(men_men_n924_), .A1(men_men_n919_), .B0(men_men_n48_), .Y(men_men_n925_));
  NO4        u0903(.A(men_men_n404_), .B(men_men_n411_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n926_));
  NA2        u0904(.A(men_men_n190_), .B(men_men_n627_), .Y(men_men_n927_));
  NOi21      u0905(.An(men_men_n927_), .B(men_men_n926_), .Y(men_men_n928_));
  NA2        u0906(.A(men_men_n777_), .B(men_men_n739_), .Y(men_men_n929_));
  NA2        u0907(.A(men_men_n354_), .B(men_men_n474_), .Y(men_men_n930_));
  OAI220     u0908(.A0(men_men_n930_), .A1(men_men_n929_), .B0(men_men_n928_), .B1(men_men_n63_), .Y(men_men_n931_));
  NOi21      u0909(.An(i_5_), .B(i_9_), .Y(men_men_n932_));
  NA2        u0910(.A(men_men_n932_), .B(i_0_), .Y(men_men_n933_));
  AOI210     u0911(.A0(men_men_n280_), .A1(men_men_n516_), .B0(men_men_n754_), .Y(men_men_n934_));
  NO3        u0912(.A(men_men_n446_), .B(men_men_n280_), .C(men_men_n73_), .Y(men_men_n935_));
  NO2        u0913(.A(men_men_n179_), .B(men_men_n150_), .Y(men_men_n936_));
  AOI210     u0914(.A0(men_men_n936_), .A1(men_men_n254_), .B0(men_men_n935_), .Y(men_men_n937_));
  OAI220     u0915(.A0(men_men_n937_), .A1(men_men_n185_), .B0(men_men_n934_), .B1(men_men_n933_), .Y(men_men_n938_));
  NO4        u0916(.A(men_men_n938_), .B(men_men_n931_), .C(men_men_n925_), .D(men_men_n917_), .Y(men_men_n939_));
  NA2        u0917(.A(men_men_n190_), .B(men_men_n24_), .Y(men_men_n940_));
  NO2        u0918(.A(men_men_n737_), .B(men_men_n654_), .Y(men_men_n941_));
  NO2        u0919(.A(men_men_n941_), .B(men_men_n940_), .Y(men_men_n942_));
  NA2        u0920(.A(men_men_n330_), .B(men_men_n132_), .Y(men_men_n943_));
  NAi21      u0921(.An(men_men_n165_), .B(men_men_n474_), .Y(men_men_n944_));
  OAI220     u0922(.A0(men_men_n944_), .A1(men_men_n904_), .B0(men_men_n943_), .B1(men_men_n432_), .Y(men_men_n945_));
  NO2        u0923(.A(men_men_n945_), .B(men_men_n942_), .Y(men_men_n946_));
  NO2        u0924(.A(men_men_n418_), .B(men_men_n310_), .Y(men_men_n947_));
  NA2        u0925(.A(men_men_n947_), .B(men_men_n779_), .Y(men_men_n948_));
  NA2        u0926(.A(men_men_n628_), .B(i_0_), .Y(men_men_n949_));
  NO3        u0927(.A(men_men_n949_), .B(men_men_n413_), .C(men_men_n89_), .Y(men_men_n950_));
  NO4        u0928(.A(men_men_n645_), .B(men_men_n223_), .C(men_men_n450_), .D(men_men_n442_), .Y(men_men_n951_));
  AOI210     u0929(.A0(men_men_n951_), .A1(i_11_), .B0(men_men_n950_), .Y(men_men_n952_));
  INV        u0930(.A(men_men_n514_), .Y(men_men_n953_));
  AN2        u0931(.A(men_men_n98_), .B(men_men_n253_), .Y(men_men_n954_));
  NA2        u0932(.A(men_men_n816_), .B(men_men_n348_), .Y(men_men_n955_));
  AOI210     u0933(.A0(men_men_n525_), .A1(men_men_n89_), .B0(men_men_n58_), .Y(men_men_n956_));
  OAI220     u0934(.A0(men_men_n956_), .A1(men_men_n955_), .B0(men_men_n722_), .B1(men_men_n587_), .Y(men_men_n957_));
  NO2        u0935(.A(men_men_n264_), .B(men_men_n156_), .Y(men_men_n958_));
  NA2        u0936(.A(i_0_), .B(i_10_), .Y(men_men_n959_));
  NO4        u0937(.A(men_men_n117_), .B(men_men_n58_), .C(men_men_n732_), .D(i_5_), .Y(men_men_n960_));
  AO220      u0938(.A0(men_men_n960_), .A1(i_10_), .B0(men_men_n958_), .B1(i_6_), .Y(men_men_n961_));
  AOI220     u0939(.A0(men_men_n354_), .A1(men_men_n100_), .B0(men_men_n190_), .B1(men_men_n84_), .Y(men_men_n962_));
  NA2        u0940(.A(men_men_n622_), .B(i_4_), .Y(men_men_n963_));
  NA2        u0941(.A(men_men_n193_), .B(men_men_n208_), .Y(men_men_n964_));
  OAI220     u0942(.A0(men_men_n964_), .A1(men_men_n955_), .B0(men_men_n963_), .B1(men_men_n962_), .Y(men_men_n965_));
  NO4        u0943(.A(men_men_n965_), .B(men_men_n961_), .C(men_men_n957_), .D(men_men_n954_), .Y(men_men_n966_));
  NA4        u0944(.A(men_men_n966_), .B(men_men_n952_), .C(men_men_n948_), .D(men_men_n946_), .Y(men_men_n967_));
  NO2        u0945(.A(men_men_n105_), .B(men_men_n37_), .Y(men_men_n968_));
  NA2        u0946(.A(i_11_), .B(i_9_), .Y(men_men_n969_));
  NO3        u0947(.A(i_12_), .B(men_men_n969_), .C(men_men_n664_), .Y(men_men_n970_));
  AO220      u0948(.A0(men_men_n970_), .A1(men_men_n968_), .B0(men_men_n282_), .B1(men_men_n88_), .Y(men_men_n971_));
  NO2        u0949(.A(men_men_n48_), .B(i_7_), .Y(men_men_n972_));
  NAi31      u0950(.An(men_men_n277_), .B(men_men_n497_), .C(men_men_n163_), .Y(men_men_n973_));
  NO2        u0951(.A(men_men_n969_), .B(men_men_n73_), .Y(men_men_n974_));
  NO2        u0952(.A(men_men_n179_), .B(i_0_), .Y(men_men_n975_));
  INV        u0953(.A(men_men_n975_), .Y(men_men_n976_));
  NA2        u0954(.A(men_men_n514_), .B(men_men_n240_), .Y(men_men_n977_));
  AOI210     u0955(.A0(men_men_n398_), .A1(men_men_n41_), .B0(men_men_n440_), .Y(men_men_n978_));
  OAI220     u0956(.A0(men_men_n978_), .A1(men_men_n933_), .B0(men_men_n977_), .B1(men_men_n976_), .Y(men_men_n979_));
  NO3        u0957(.A(men_men_n979_), .B(men_men_n973_), .C(men_men_n971_), .Y(men_men_n980_));
  AOI210     u0958(.A0(men_men_n483_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n981_));
  NA2        u0959(.A(men_men_n175_), .B(men_men_n105_), .Y(men_men_n982_));
  NOi32      u0960(.An(men_men_n981_), .Bn(men_men_n193_), .C(men_men_n982_), .Y(men_men_n983_));
  AOI210     u0961(.A0(men_men_n666_), .A1(men_men_n348_), .B0(men_men_n253_), .Y(men_men_n984_));
  NO2        u0962(.A(men_men_n984_), .B(men_men_n922_), .Y(men_men_n985_));
  NO2        u0963(.A(men_men_n985_), .B(men_men_n983_), .Y(men_men_n986_));
  NOi21      u0964(.An(i_7_), .B(i_5_), .Y(men_men_n987_));
  NOi31      u0965(.An(men_men_n987_), .B(i_0_), .C(men_men_n795_), .Y(men_men_n988_));
  NA3        u0966(.A(men_men_n988_), .B(men_men_n412_), .C(i_6_), .Y(men_men_n989_));
  OA210      u0967(.A0(men_men_n982_), .A1(men_men_n563_), .B0(men_men_n989_), .Y(men_men_n990_));
  NO3        u0968(.A(men_men_n435_), .B(men_men_n387_), .C(men_men_n383_), .Y(men_men_n991_));
  NO2        u0969(.A(men_men_n274_), .B(men_men_n337_), .Y(men_men_n992_));
  NO2        u0970(.A(men_men_n795_), .B(men_men_n269_), .Y(men_men_n993_));
  AOI210     u0971(.A0(men_men_n993_), .A1(men_men_n992_), .B0(men_men_n991_), .Y(men_men_n994_));
  NA4        u0972(.A(men_men_n994_), .B(men_men_n990_), .C(men_men_n986_), .D(men_men_n980_), .Y(men_men_n995_));
  NO2        u0973(.A(men_men_n940_), .B(men_men_n249_), .Y(men_men_n996_));
  AN2        u0974(.A(men_men_n353_), .B(men_men_n348_), .Y(men_men_n997_));
  AO220      u0975(.A0(men_men_n997_), .A1(men_men_n936_), .B0(men_men_n369_), .B1(men_men_n27_), .Y(men_men_n998_));
  OAI210     u0976(.A0(men_men_n998_), .A1(men_men_n996_), .B0(i_10_), .Y(men_men_n999_));
  NO2        u0977(.A(men_men_n910_), .B(men_men_n336_), .Y(men_men_n1000_));
  OA210      u0978(.A0(men_men_n514_), .A1(men_men_n232_), .B0(men_men_n513_), .Y(men_men_n1001_));
  NA2        u0979(.A(men_men_n1000_), .B(men_men_n974_), .Y(men_men_n1002_));
  NA3        u0980(.A(men_men_n513_), .B(men_men_n443_), .C(men_men_n45_), .Y(men_men_n1003_));
  OAI210     u0981(.A0(men_men_n944_), .A1(men_men_n953_), .B0(men_men_n1003_), .Y(men_men_n1004_));
  NO2        u0982(.A(men_men_n267_), .B(men_men_n46_), .Y(men_men_n1005_));
  NA2        u0983(.A(men_men_n974_), .B(men_men_n323_), .Y(men_men_n1006_));
  OAI210     u0984(.A0(men_men_n1005_), .A1(men_men_n192_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  AOI220     u0985(.A0(men_men_n1007_), .A1(men_men_n514_), .B0(men_men_n1004_), .B1(men_men_n73_), .Y(men_men_n1008_));
  NA3        u0986(.A(men_men_n885_), .B(men_men_n410_), .C(men_men_n704_), .Y(men_men_n1009_));
  NA2        u0987(.A(men_men_n94_), .B(men_men_n44_), .Y(men_men_n1010_));
  NO2        u0988(.A(men_men_n75_), .B(men_men_n818_), .Y(men_men_n1011_));
  AOI220     u0989(.A0(men_men_n1011_), .A1(men_men_n1010_), .B0(men_men_n178_), .B1(men_men_n654_), .Y(men_men_n1012_));
  AOI210     u0990(.A0(men_men_n1012_), .A1(men_men_n1009_), .B0(men_men_n47_), .Y(men_men_n1013_));
  NO3        u0991(.A(men_men_n645_), .B(men_men_n382_), .C(men_men_n24_), .Y(men_men_n1014_));
  AOI210     u0992(.A0(men_men_n770_), .A1(men_men_n599_), .B0(men_men_n1014_), .Y(men_men_n1015_));
  NAi21      u0993(.An(i_9_), .B(i_5_), .Y(men_men_n1016_));
  NO2        u0994(.A(men_men_n1016_), .B(men_men_n435_), .Y(men_men_n1017_));
  NO2        u0995(.A(men_men_n660_), .B(men_men_n107_), .Y(men_men_n1018_));
  AOI220     u0996(.A0(men_men_n1018_), .A1(i_0_), .B0(men_men_n1017_), .B1(men_men_n683_), .Y(men_men_n1019_));
  OAI220     u0997(.A0(men_men_n1019_), .A1(men_men_n86_), .B0(men_men_n1015_), .B1(men_men_n176_), .Y(men_men_n1020_));
  NO3        u0998(.A(men_men_n1020_), .B(men_men_n1013_), .C(men_men_n567_), .Y(men_men_n1021_));
  NA4        u0999(.A(men_men_n1021_), .B(men_men_n1008_), .C(men_men_n1002_), .D(men_men_n999_), .Y(men_men_n1022_));
  NO3        u1000(.A(men_men_n1022_), .B(men_men_n995_), .C(men_men_n967_), .Y(men_men_n1023_));
  NO2        u1001(.A(i_0_), .B(men_men_n795_), .Y(men_men_n1024_));
  NA2        u1002(.A(men_men_n73_), .B(men_men_n44_), .Y(men_men_n1025_));
  NA2        u1003(.A(men_men_n959_), .B(men_men_n1025_), .Y(men_men_n1026_));
  NO3        u1004(.A(men_men_n107_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n1027_));
  AO220      u1005(.A0(men_men_n1027_), .A1(men_men_n1026_), .B0(men_men_n1024_), .B1(men_men_n178_), .Y(men_men_n1028_));
  AOI210     u1006(.A0(men_men_n864_), .A1(men_men_n752_), .B0(men_men_n982_), .Y(men_men_n1029_));
  AOI210     u1007(.A0(men_men_n1028_), .A1(men_men_n371_), .B0(men_men_n1029_), .Y(men_men_n1030_));
  NA2        u1008(.A(men_men_n806_), .B(men_men_n148_), .Y(men_men_n1031_));
  INV        u1009(.A(men_men_n1031_), .Y(men_men_n1032_));
  NA3        u1010(.A(men_men_n1032_), .B(men_men_n739_), .C(men_men_n73_), .Y(men_men_n1033_));
  NO2        u1011(.A(men_men_n881_), .B(men_men_n435_), .Y(men_men_n1034_));
  NA3        u1012(.A(men_men_n912_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n1035_));
  NA2        u1013(.A(men_men_n913_), .B(i_9_), .Y(men_men_n1036_));
  AOI210     u1014(.A0(men_men_n1035_), .A1(men_men_n542_), .B0(men_men_n1036_), .Y(men_men_n1037_));
  OAI210     u1015(.A0(men_men_n254_), .A1(i_9_), .B0(men_men_n239_), .Y(men_men_n1038_));
  AOI210     u1016(.A0(men_men_n1038_), .A1(men_men_n949_), .B0(men_men_n156_), .Y(men_men_n1039_));
  NO3        u1017(.A(men_men_n1039_), .B(men_men_n1037_), .C(men_men_n1034_), .Y(men_men_n1040_));
  NA3        u1018(.A(men_men_n1040_), .B(men_men_n1033_), .C(men_men_n1030_), .Y(men_men_n1041_));
  NA2        u1019(.A(men_men_n997_), .B(men_men_n400_), .Y(men_men_n1042_));
  AOI210     u1020(.A0(men_men_n317_), .A1(men_men_n165_), .B0(men_men_n1042_), .Y(men_men_n1043_));
  NA3        u1021(.A(men_men_n39_), .B(men_men_n28_), .C(men_men_n44_), .Y(men_men_n1044_));
  NA2        u1022(.A(men_men_n972_), .B(men_men_n530_), .Y(men_men_n1045_));
  AOI210     u1023(.A0(men_men_n1044_), .A1(men_men_n165_), .B0(men_men_n1045_), .Y(men_men_n1046_));
  NO2        u1024(.A(men_men_n1046_), .B(men_men_n1043_), .Y(men_men_n1047_));
  NO2        u1025(.A(men_men_n959_), .B(men_men_n195_), .Y(men_men_n1048_));
  AOI220     u1026(.A0(men_men_n1048_), .A1(i_11_), .B0(men_men_n623_), .B1(men_men_n75_), .Y(men_men_n1049_));
  INV        u1027(.A(men_men_n226_), .Y(men_men_n1050_));
  OAI220     u1028(.A0(men_men_n580_), .A1(men_men_n142_), .B0(men_men_n708_), .B1(men_men_n677_), .Y(men_men_n1051_));
  NA3        u1029(.A(men_men_n1051_), .B(men_men_n427_), .C(men_men_n1050_), .Y(men_men_n1052_));
  NA3        u1030(.A(men_men_n1052_), .B(men_men_n1049_), .C(men_men_n1047_), .Y(men_men_n1053_));
  NO2        u1031(.A(men_men_n252_), .B(men_men_n94_), .Y(men_men_n1054_));
  AOI210     u1032(.A0(men_men_n1054_), .A1(men_men_n1024_), .B0(men_men_n111_), .Y(men_men_n1055_));
  AOI220     u1033(.A0(men_men_n987_), .A1(men_men_n530_), .B0(men_men_n912_), .B1(men_men_n166_), .Y(men_men_n1056_));
  NA2        u1034(.A(men_men_n374_), .B(men_men_n180_), .Y(men_men_n1057_));
  OA220      u1035(.A0(men_men_n1057_), .A1(men_men_n1056_), .B0(men_men_n1055_), .B1(i_5_), .Y(men_men_n1058_));
  AOI210     u1036(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n179_), .Y(men_men_n1059_));
  NA2        u1037(.A(men_men_n1059_), .B(men_men_n1001_), .Y(men_men_n1060_));
  NA3        u1038(.A(men_men_n674_), .B(men_men_n190_), .C(men_men_n84_), .Y(men_men_n1061_));
  NA2        u1039(.A(men_men_n1061_), .B(men_men_n597_), .Y(men_men_n1062_));
  NO3        u1040(.A(men_men_n922_), .B(men_men_n54_), .C(men_men_n48_), .Y(men_men_n1063_));
  NA3        u1041(.A(men_men_n535_), .B(men_men_n528_), .C(men_men_n511_), .Y(men_men_n1064_));
  NO3        u1042(.A(men_men_n1064_), .B(men_men_n1063_), .C(men_men_n1062_), .Y(men_men_n1065_));
  NA3        u1043(.A(men_men_n418_), .B(men_men_n175_), .C(men_men_n174_), .Y(men_men_n1066_));
  NA3        u1044(.A(men_men_n972_), .B(men_men_n306_), .C(men_men_n239_), .Y(men_men_n1067_));
  NA2        u1045(.A(men_men_n1067_), .B(men_men_n1066_), .Y(men_men_n1068_));
  NA3        u1046(.A(men_men_n418_), .B(men_men_n355_), .C(men_men_n230_), .Y(men_men_n1069_));
  INV        u1047(.A(men_men_n1069_), .Y(men_men_n1070_));
  NOi31      u1048(.An(men_men_n417_), .B(men_men_n1025_), .C(men_men_n249_), .Y(men_men_n1071_));
  NO2        u1049(.A(men_men_n969_), .B(men_men_n195_), .Y(men_men_n1072_));
  NO4        u1050(.A(men_men_n1072_), .B(men_men_n1071_), .C(men_men_n1070_), .D(men_men_n1068_), .Y(men_men_n1073_));
  NA4        u1051(.A(men_men_n1073_), .B(men_men_n1065_), .C(men_men_n1060_), .D(men_men_n1058_), .Y(men_men_n1074_));
  AOI210     u1052(.A0(men_men_n622_), .A1(men_men_n579_), .B0(men_men_n676_), .Y(men_men_n1075_));
  NO3        u1053(.A(men_men_n1075_), .B(men_men_n613_), .C(men_men_n368_), .Y(men_men_n1076_));
  NO2        u1054(.A(men_men_n86_), .B(i_5_), .Y(men_men_n1077_));
  NA3        u1055(.A(men_men_n913_), .B(men_men_n112_), .C(men_men_n127_), .Y(men_men_n1078_));
  INV        u1056(.A(men_men_n1078_), .Y(men_men_n1079_));
  AOI210     u1057(.A0(men_men_n1079_), .A1(men_men_n1077_), .B0(men_men_n1076_), .Y(men_men_n1080_));
  NA3        u1058(.A(men_men_n323_), .B(i_5_), .C(men_men_n198_), .Y(men_men_n1081_));
  NAi31      u1059(.An(men_men_n251_), .B(men_men_n1081_), .C(men_men_n252_), .Y(men_men_n1082_));
  NO4        u1060(.A(men_men_n249_), .B(men_men_n217_), .C(i_0_), .D(i_12_), .Y(men_men_n1083_));
  AOI220     u1061(.A0(men_men_n1083_), .A1(men_men_n1082_), .B0(men_men_n859_), .B1(men_men_n180_), .Y(men_men_n1084_));
  AN2        u1062(.A(men_men_n959_), .B(men_men_n156_), .Y(men_men_n1085_));
  NO4        u1063(.A(men_men_n1085_), .B(i_12_), .C(men_men_n712_), .D(men_men_n134_), .Y(men_men_n1086_));
  NA2        u1064(.A(men_men_n1086_), .B(men_men_n226_), .Y(men_men_n1087_));
  NA3        u1065(.A(men_men_n100_), .B(men_men_n627_), .C(i_11_), .Y(men_men_n1088_));
  NO2        u1066(.A(men_men_n1088_), .B(men_men_n158_), .Y(men_men_n1089_));
  NA2        u1067(.A(men_men_n987_), .B(men_men_n510_), .Y(men_men_n1090_));
  NA2        u1068(.A(men_men_n64_), .B(men_men_n103_), .Y(men_men_n1091_));
  OAI220     u1069(.A0(men_men_n1091_), .A1(men_men_n1081_), .B0(men_men_n1090_), .B1(men_men_n740_), .Y(men_men_n1092_));
  AOI210     u1070(.A0(men_men_n1092_), .A1(men_men_n975_), .B0(men_men_n1089_), .Y(men_men_n1093_));
  NA4        u1071(.A(men_men_n1093_), .B(men_men_n1087_), .C(men_men_n1084_), .D(men_men_n1080_), .Y(men_men_n1094_));
  NO4        u1072(.A(men_men_n1094_), .B(men_men_n1074_), .C(men_men_n1053_), .D(men_men_n1041_), .Y(men_men_n1095_));
  OAI210     u1073(.A0(men_men_n884_), .A1(men_men_n877_), .B0(men_men_n37_), .Y(men_men_n1096_));
  NA3        u1074(.A(men_men_n981_), .B(men_men_n395_), .C(i_5_), .Y(men_men_n1097_));
  NA3        u1075(.A(men_men_n1097_), .B(men_men_n1096_), .C(men_men_n672_), .Y(men_men_n1098_));
  NA2        u1076(.A(men_men_n1098_), .B(men_men_n213_), .Y(men_men_n1099_));
  AN2        u1077(.A(men_men_n765_), .B(men_men_n396_), .Y(men_men_n1100_));
  NA2        u1078(.A(men_men_n191_), .B(men_men_n193_), .Y(men_men_n1101_));
  AO210      u1079(.A0(men_men_n1100_), .A1(men_men_n33_), .B0(men_men_n1101_), .Y(men_men_n1102_));
  OAI210     u1080(.A0(men_men_n676_), .A1(men_men_n674_), .B0(men_men_n336_), .Y(men_men_n1103_));
  NAi31      u1081(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1104_));
  NO2        u1082(.A(men_men_n70_), .B(men_men_n1104_), .Y(men_men_n1105_));
  NO2        u1083(.A(men_men_n1105_), .B(men_men_n709_), .Y(men_men_n1106_));
  NA3        u1084(.A(men_men_n1106_), .B(men_men_n1103_), .C(men_men_n1102_), .Y(men_men_n1107_));
  NO2        u1085(.A(men_men_n500_), .B(men_men_n280_), .Y(men_men_n1108_));
  NO4        u1086(.A(men_men_n242_), .B(men_men_n147_), .C(men_men_n743_), .D(men_men_n37_), .Y(men_men_n1109_));
  NO3        u1087(.A(men_men_n1109_), .B(men_men_n1108_), .C(men_men_n951_), .Y(men_men_n1110_));
  OAI210     u1088(.A0(men_men_n1088_), .A1(men_men_n150_), .B0(men_men_n1110_), .Y(men_men_n1111_));
  AOI210     u1089(.A0(men_men_n1107_), .A1(men_men_n48_), .B0(men_men_n1111_), .Y(men_men_n1112_));
  AOI210     u1090(.A0(men_men_n1112_), .A1(men_men_n1099_), .B0(men_men_n73_), .Y(men_men_n1113_));
  NO2        u1091(.A(men_men_n620_), .B(men_men_n407_), .Y(men_men_n1114_));
  NO2        u1092(.A(men_men_n1114_), .B(men_men_n823_), .Y(men_men_n1115_));
  OAI210     u1093(.A0(men_men_n80_), .A1(men_men_n54_), .B0(men_men_n110_), .Y(men_men_n1116_));
  NA2        u1094(.A(men_men_n1116_), .B(men_men_n76_), .Y(men_men_n1117_));
  AOI210     u1095(.A0(men_men_n1059_), .A1(men_men_n972_), .B0(men_men_n988_), .Y(men_men_n1118_));
  AOI210     u1096(.A0(men_men_n1118_), .A1(men_men_n1117_), .B0(men_men_n743_), .Y(men_men_n1119_));
  NA2        u1097(.A(men_men_n274_), .B(men_men_n57_), .Y(men_men_n1120_));
  AOI220     u1098(.A0(men_men_n1120_), .A1(men_men_n76_), .B0(men_men_n369_), .B1(men_men_n266_), .Y(men_men_n1121_));
  NO2        u1099(.A(men_men_n1121_), .B(men_men_n246_), .Y(men_men_n1122_));
  NA3        u1100(.A(men_men_n98_), .B(men_men_n325_), .C(men_men_n31_), .Y(men_men_n1123_));
  INV        u1101(.A(men_men_n1123_), .Y(men_men_n1124_));
  NO3        u1102(.A(men_men_n1124_), .B(men_men_n1122_), .C(men_men_n1119_), .Y(men_men_n1125_));
  OAI210     u1103(.A0(men_men_n282_), .A1(men_men_n161_), .B0(men_men_n89_), .Y(men_men_n1126_));
  NA3        u1104(.A(men_men_n827_), .B(men_men_n306_), .C(men_men_n80_), .Y(men_men_n1127_));
  AOI210     u1105(.A0(men_men_n1127_), .A1(men_men_n1126_), .B0(i_11_), .Y(men_men_n1128_));
  NA2        u1106(.A(men_men_n667_), .B(men_men_n223_), .Y(men_men_n1129_));
  OAI210     u1107(.A0(men_men_n1129_), .A1(men_men_n981_), .B0(men_men_n213_), .Y(men_men_n1130_));
  NA2        u1108(.A(men_men_n167_), .B(i_5_), .Y(men_men_n1131_));
  AOI210     u1109(.A0(men_men_n1130_), .A1(men_men_n839_), .B0(men_men_n1131_), .Y(men_men_n1132_));
  NO3        u1110(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1133_));
  OAI210     u1111(.A0(men_men_n992_), .A1(men_men_n325_), .B0(men_men_n1133_), .Y(men_men_n1134_));
  NO2        u1112(.A(men_men_n1134_), .B(men_men_n795_), .Y(men_men_n1135_));
  NO4        u1113(.A(men_men_n1016_), .B(men_men_n518_), .C(men_men_n263_), .D(men_men_n262_), .Y(men_men_n1136_));
  NO2        u1114(.A(men_men_n1136_), .B(men_men_n617_), .Y(men_men_n1137_));
  NO2        u1115(.A(men_men_n880_), .B(men_men_n388_), .Y(men_men_n1138_));
  AOI210     u1116(.A0(men_men_n1138_), .A1(men_men_n1137_), .B0(men_men_n40_), .Y(men_men_n1139_));
  NO4        u1117(.A(men_men_n1139_), .B(men_men_n1135_), .C(men_men_n1132_), .D(men_men_n1128_), .Y(men_men_n1140_));
  OAI210     u1118(.A0(men_men_n1125_), .A1(i_4_), .B0(men_men_n1140_), .Y(men_men_n1141_));
  NO3        u1119(.A(men_men_n1141_), .B(men_men_n1115_), .C(men_men_n1113_), .Y(men_men_n1142_));
  NA4        u1120(.A(men_men_n1142_), .B(men_men_n1095_), .C(men_men_n1023_), .D(men_men_n939_), .Y(men4));
  INV        u1121(.A(men_men_n769_), .Y(men_men_n1146_));
  INV        u1122(.A(i_5_), .Y(men_men_n1147_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule