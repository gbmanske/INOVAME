//Benchmark atmr_prom1_2672_0.25

module atmr_prom1(x0, x1, x2, x3, x4, x5, x6, x7, x8, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27, z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27, z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39;
 wire ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1374_, ori_ori_n1376_, ori_ori_n1377_, ori_ori_n1378_, ori_ori_n1379_, ori_ori_n1380_, ori_ori_n1381_, ori_ori_n1382_, ori_ori_n1383_, ori_ori_n1384_, ori_ori_n1385_, ori_ori_n1386_, ori_ori_n1387_, ori_ori_n1388_, ori_ori_n1389_, ori_ori_n1390_, ori_ori_n1391_, ori_ori_n1392_, ori_ori_n1393_, ori_ori_n1394_, ori_ori_n1395_, ori_ori_n1396_, ori_ori_n1397_, ori_ori_n1398_, ori_ori_n1399_, ori_ori_n1400_, ori_ori_n1401_, ori_ori_n1402_, ori_ori_n1403_, ori_ori_n1404_, ori_ori_n1405_, ori_ori_n1406_, ori_ori_n1407_, ori_ori_n1408_, ori_ori_n1409_, ori_ori_n1410_, ori_ori_n1411_, ori_ori_n1412_, ori_ori_n1413_, ori_ori_n1414_, ori_ori_n1415_, ori_ori_n1416_, ori_ori_n1417_, ori_ori_n1418_, ori_ori_n1419_, ori_ori_n1420_, ori_ori_n1421_, ori_ori_n1422_, ori_ori_n1423_, ori_ori_n1424_, ori_ori_n1425_, ori_ori_n1426_, ori_ori_n1427_, ori_ori_n1428_, ori_ori_n1429_, ori_ori_n1430_, ori_ori_n1431_, ori_ori_n1432_, ori_ori_n1433_, ori_ori_n1434_, ori_ori_n1435_, ori_ori_n1436_, ori_ori_n1437_, ori_ori_n1438_, ori_ori_n1439_, ori_ori_n1441_, ori_ori_n1442_, ori_ori_n1443_, ori_ori_n1444_, ori_ori_n1445_, ori_ori_n1446_, ori_ori_n1447_, ori_ori_n1448_, ori_ori_n1449_, ori_ori_n1450_, ori_ori_n1451_, ori_ori_n1452_, ori_ori_n1453_, ori_ori_n1454_, ori_ori_n1455_, ori_ori_n1456_, ori_ori_n1457_, ori_ori_n1458_, ori_ori_n1459_, ori_ori_n1460_, ori_ori_n1461_, ori_ori_n1462_, ori_ori_n1463_, ori_ori_n1464_, ori_ori_n1465_, ori_ori_n1466_, ori_ori_n1467_, ori_ori_n1468_, ori_ori_n1469_, ori_ori_n1470_, ori_ori_n1471_, ori_ori_n1472_, ori_ori_n1473_, ori_ori_n1474_, ori_ori_n1475_, ori_ori_n1476_, ori_ori_n1477_, ori_ori_n1478_, ori_ori_n1479_, ori_ori_n1480_, ori_ori_n1481_, ori_ori_n1482_, ori_ori_n1483_, ori_ori_n1484_, ori_ori_n1485_, ori_ori_n1486_, ori_ori_n1487_, ori_ori_n1488_, ori_ori_n1489_, ori_ori_n1490_, ori_ori_n1491_, ori_ori_n1492_, ori_ori_n1493_, ori_ori_n1494_, ori_ori_n1495_, ori_ori_n1497_, ori_ori_n1498_, ori_ori_n1499_, ori_ori_n1500_, ori_ori_n1501_, ori_ori_n1502_, ori_ori_n1503_, ori_ori_n1504_, ori_ori_n1505_, ori_ori_n1506_, ori_ori_n1507_, ori_ori_n1508_, ori_ori_n1509_, ori_ori_n1510_, ori_ori_n1511_, ori_ori_n1512_, ori_ori_n1513_, ori_ori_n1514_, ori_ori_n1515_, ori_ori_n1516_, ori_ori_n1517_, ori_ori_n1518_, ori_ori_n1519_, ori_ori_n1520_, ori_ori_n1522_, ori_ori_n1523_, ori_ori_n1524_, ori_ori_n1525_, ori_ori_n1526_, ori_ori_n1527_, ori_ori_n1528_, ori_ori_n1529_, ori_ori_n1530_, ori_ori_n1531_, ori_ori_n1532_, ori_ori_n1533_, ori_ori_n1534_, ori_ori_n1535_, ori_ori_n1536_, ori_ori_n1537_, ori_ori_n1538_, ori_ori_n1539_, ori_ori_n1540_, ori_ori_n1541_, ori_ori_n1542_, ori_ori_n1543_, ori_ori_n1544_, ori_ori_n1545_, ori_ori_n1546_, ori_ori_n1547_, ori_ori_n1548_, ori_ori_n1549_, ori_ori_n1550_, ori_ori_n1551_, ori_ori_n1552_, ori_ori_n1553_, ori_ori_n1554_, ori_ori_n1555_, ori_ori_n1556_, ori_ori_n1557_, ori_ori_n1558_, ori_ori_n1559_, ori_ori_n1560_, ori_ori_n1561_, ori_ori_n1562_, ori_ori_n1563_, ori_ori_n1564_, ori_ori_n1565_, ori_ori_n1566_, ori_ori_n1567_, ori_ori_n1568_, ori_ori_n1569_, ori_ori_n1570_, ori_ori_n1571_, ori_ori_n1572_, ori_ori_n1573_, ori_ori_n1574_, ori_ori_n1575_, ori_ori_n1576_, ori_ori_n1577_, ori_ori_n1578_, ori_ori_n1579_, ori_ori_n1580_, ori_ori_n1581_, ori_ori_n1582_, ori_ori_n1583_, ori_ori_n1584_, ori_ori_n1585_, ori_ori_n1586_, ori_ori_n1587_, ori_ori_n1588_, ori_ori_n1589_, ori_ori_n1590_, ori_ori_n1591_, ori_ori_n1592_, ori_ori_n1593_, ori_ori_n1594_, ori_ori_n1595_, ori_ori_n1596_, ori_ori_n1597_, ori_ori_n1598_, ori_ori_n1599_, ori_ori_n1600_, ori_ori_n1601_, ori_ori_n1602_, ori_ori_n1603_, ori_ori_n1605_, ori_ori_n1606_, ori_ori_n1607_, ori_ori_n1608_, ori_ori_n1609_, ori_ori_n1610_, ori_ori_n1611_, ori_ori_n1612_, ori_ori_n1613_, ori_ori_n1614_, ori_ori_n1615_, ori_ori_n1616_, ori_ori_n1617_, ori_ori_n1618_, ori_ori_n1619_, ori_ori_n1620_, ori_ori_n1621_, ori_ori_n1622_, ori_ori_n1623_, ori_ori_n1624_, ori_ori_n1625_, ori_ori_n1626_, ori_ori_n1627_, ori_ori_n1628_, ori_ori_n1629_, ori_ori_n1630_, ori_ori_n1631_, ori_ori_n1632_, ori_ori_n1633_, ori_ori_n1634_, ori_ori_n1635_, ori_ori_n1636_, ori_ori_n1637_, ori_ori_n1638_, ori_ori_n1639_, ori_ori_n1640_, ori_ori_n1641_, ori_ori_n1642_, ori_ori_n1643_, ori_ori_n1644_, ori_ori_n1645_, ori_ori_n1646_, ori_ori_n1647_, ori_ori_n1648_, ori_ori_n1649_, ori_ori_n1650_, ori_ori_n1651_, ori_ori_n1652_, ori_ori_n1653_, ori_ori_n1654_, ori_ori_n1656_, ori_ori_n1657_, ori_ori_n1658_, ori_ori_n1659_, ori_ori_n1660_, ori_ori_n1661_, ori_ori_n1662_, ori_ori_n1663_, ori_ori_n1664_, ori_ori_n1665_, ori_ori_n1666_, ori_ori_n1667_, ori_ori_n1668_, ori_ori_n1669_, ori_ori_n1670_, ori_ori_n1671_, ori_ori_n1673_, ori_ori_n1674_, ori_ori_n1675_, ori_ori_n1676_, ori_ori_n1677_, ori_ori_n1678_, ori_ori_n1679_, ori_ori_n1680_, ori_ori_n1681_, ori_ori_n1682_, ori_ori_n1683_, ori_ori_n1685_, ori_ori_n1686_, ori_ori_n1687_, ori_ori_n1688_, ori_ori_n1689_, ori_ori_n1690_, ori_ori_n1691_, ori_ori_n1692_, ori_ori_n1694_, ori_ori_n1695_, ori_ori_n1696_, ori_ori_n1697_, ori_ori_n1698_, ori_ori_n1699_, ori_ori_n1700_, ori_ori_n1701_, ori_ori_n1702_, ori_ori_n1703_, ori_ori_n1704_, ori_ori_n1705_, ori_ori_n1706_, ori_ori_n1707_, ori_ori_n1708_, ori_ori_n1709_, ori_ori_n1710_, ori_ori_n1711_, ori_ori_n1712_, ori_ori_n1713_, ori_ori_n1714_, ori_ori_n1715_, ori_ori_n1716_, ori_ori_n1717_, ori_ori_n1718_, ori_ori_n1719_, ori_ori_n1720_, ori_ori_n1721_, ori_ori_n1722_, ori_ori_n1723_, ori_ori_n1724_, ori_ori_n1725_, ori_ori_n1726_, ori_ori_n1727_, ori_ori_n1729_, ori_ori_n1730_, ori_ori_n1731_, ori_ori_n1732_, ori_ori_n1733_, ori_ori_n1734_, ori_ori_n1735_, ori_ori_n1736_, ori_ori_n1737_, ori_ori_n1738_, ori_ori_n1739_, ori_ori_n1740_, ori_ori_n1741_, ori_ori_n1743_, ori_ori_n1744_, ori_ori_n1745_, ori_ori_n1746_, ori_ori_n1747_, ori_ori_n1748_, ori_ori_n1749_, ori_ori_n1750_, ori_ori_n1751_, ori_ori_n1752_, ori_ori_n1753_, ori_ori_n1754_, ori_ori_n1755_, ori_ori_n1756_, ori_ori_n1757_, ori_ori_n1758_, ori_ori_n1759_, ori_ori_n1760_, ori_ori_n1761_, ori_ori_n1762_, ori_ori_n1763_, ori_ori_n1764_, ori_ori_n1765_, ori_ori_n1766_, ori_ori_n1767_, ori_ori_n1768_, ori_ori_n1769_, ori_ori_n1770_, ori_ori_n1771_, ori_ori_n1772_, ori_ori_n1773_, ori_ori_n1774_, ori_ori_n1775_, ori_ori_n1776_, ori_ori_n1777_, ori_ori_n1778_, ori_ori_n1779_, ori_ori_n1780_, ori_ori_n1781_, ori_ori_n1782_, ori_ori_n1783_, ori_ori_n1784_, ori_ori_n1785_, ori_ori_n1786_, ori_ori_n1787_, ori_ori_n1788_, ori_ori_n1790_, ori_ori_n1791_, ori_ori_n1792_, ori_ori_n1793_, ori_ori_n1794_, ori_ori_n1795_, ori_ori_n1796_, ori_ori_n1797_, ori_ori_n1798_, ori_ori_n1799_, ori_ori_n1800_, ori_ori_n1801_, ori_ori_n1802_, ori_ori_n1803_, ori_ori_n1804_, ori_ori_n1805_, ori_ori_n1806_, ori_ori_n1807_, ori_ori_n1808_, ori_ori_n1809_, ori_ori_n1810_, ori_ori_n1811_, ori_ori_n1812_, ori_ori_n1813_, ori_ori_n1814_, ori_ori_n1815_, ori_ori_n1816_, ori_ori_n1817_, ori_ori_n1818_, ori_ori_n1819_, ori_ori_n1820_, ori_ori_n1821_, ori_ori_n1822_, ori_ori_n1823_, ori_ori_n1824_, ori_ori_n1825_, ori_ori_n1826_, ori_ori_n1827_, ori_ori_n1828_, ori_ori_n1829_, ori_ori_n1830_, ori_ori_n1831_, ori_ori_n1832_, ori_ori_n1833_, ori_ori_n1834_, ori_ori_n1835_, ori_ori_n1836_, ori_ori_n1837_, ori_ori_n1838_, ori_ori_n1839_, ori_ori_n1840_, ori_ori_n1841_, ori_ori_n1842_, ori_ori_n1843_, ori_ori_n1844_, ori_ori_n1845_, ori_ori_n1846_, ori_ori_n1847_, ori_ori_n1848_, ori_ori_n1849_, ori_ori_n1850_, ori_ori_n1851_, ori_ori_n1852_, ori_ori_n1853_, ori_ori_n1854_, ori_ori_n1856_, ori_ori_n1857_, ori_ori_n1858_, ori_ori_n1859_, ori_ori_n1860_, ori_ori_n1861_, ori_ori_n1862_, ori_ori_n1863_, ori_ori_n1864_, ori_ori_n1865_, ori_ori_n1866_, ori_ori_n1867_, ori_ori_n1868_, ori_ori_n1869_, ori_ori_n1870_, ori_ori_n1871_, ori_ori_n1872_, ori_ori_n1873_, ori_ori_n1874_, ori_ori_n1875_, ori_ori_n1876_, ori_ori_n1877_, ori_ori_n1878_, ori_ori_n1879_, ori_ori_n1880_, ori_ori_n1881_, ori_ori_n1882_, ori_ori_n1883_, ori_ori_n1884_, ori_ori_n1885_, ori_ori_n1886_, ori_ori_n1887_, ori_ori_n1888_, ori_ori_n1889_, ori_ori_n1890_, ori_ori_n1891_, ori_ori_n1892_, ori_ori_n1893_, ori_ori_n1894_, ori_ori_n1895_, ori_ori_n1896_, ori_ori_n1897_, ori_ori_n1898_, ori_ori_n1899_, ori_ori_n1900_, ori_ori_n1901_, ori_ori_n1902_, ori_ori_n1903_, ori_ori_n1904_, ori_ori_n1905_, ori_ori_n1906_, ori_ori_n1907_, ori_ori_n1908_, ori_ori_n1909_, ori_ori_n1910_, ori_ori_n1911_, ori_ori_n1912_, ori_ori_n1913_, ori_ori_n1914_, ori_ori_n1915_, ori_ori_n1916_, ori_ori_n1917_, ori_ori_n1918_, ori_ori_n1919_, ori_ori_n1920_, ori_ori_n1921_, ori_ori_n1922_, ori_ori_n1923_, ori_ori_n1924_, ori_ori_n1925_, ori_ori_n1926_, ori_ori_n1927_, ori_ori_n1928_, ori_ori_n1929_, ori_ori_n1930_, ori_ori_n1931_, ori_ori_n1933_, ori_ori_n1934_, ori_ori_n1935_, ori_ori_n1936_, ori_ori_n1937_, ori_ori_n1938_, ori_ori_n1939_, ori_ori_n1940_, ori_ori_n1941_, ori_ori_n1942_, ori_ori_n1943_, ori_ori_n1944_, ori_ori_n1945_, ori_ori_n1946_, ori_ori_n1947_, ori_ori_n1948_, ori_ori_n1949_, ori_ori_n1950_, ori_ori_n1951_, ori_ori_n1952_, ori_ori_n1953_, ori_ori_n1954_, ori_ori_n1955_, ori_ori_n1956_, ori_ori_n1957_, ori_ori_n1958_, ori_ori_n1959_, ori_ori_n1960_, ori_ori_n1961_, ori_ori_n1962_, ori_ori_n1963_, ori_ori_n1964_, ori_ori_n1965_, ori_ori_n1966_, ori_ori_n1967_, ori_ori_n1968_, ori_ori_n1969_, ori_ori_n1970_, ori_ori_n1971_, ori_ori_n1972_, ori_ori_n1973_, ori_ori_n1974_, ori_ori_n1975_, ori_ori_n1976_, ori_ori_n1977_, ori_ori_n1978_, ori_ori_n1979_, ori_ori_n1980_, ori_ori_n1981_, ori_ori_n1982_, ori_ori_n1983_, ori_ori_n1984_, ori_ori_n1985_, ori_ori_n1986_, ori_ori_n1987_, ori_ori_n1988_, ori_ori_n1989_, ori_ori_n1990_, ori_ori_n1991_, ori_ori_n1992_, ori_ori_n1993_, ori_ori_n1994_, ori_ori_n1995_, ori_ori_n1996_, ori_ori_n1997_, ori_ori_n1998_, ori_ori_n1999_, ori_ori_n2000_, ori_ori_n2001_, ori_ori_n2002_, ori_ori_n2004_, ori_ori_n2005_, ori_ori_n2006_, ori_ori_n2007_, ori_ori_n2008_, ori_ori_n2009_, ori_ori_n2010_, ori_ori_n2011_, ori_ori_n2012_, ori_ori_n2013_, ori_ori_n2014_, ori_ori_n2015_, ori_ori_n2016_, ori_ori_n2017_, ori_ori_n2018_, ori_ori_n2019_, ori_ori_n2020_, ori_ori_n2021_, ori_ori_n2022_, ori_ori_n2023_, ori_ori_n2024_, ori_ori_n2025_, ori_ori_n2026_, ori_ori_n2027_, ori_ori_n2028_, ori_ori_n2029_, ori_ori_n2030_, ori_ori_n2031_, ori_ori_n2032_, ori_ori_n2033_, ori_ori_n2034_, ori_ori_n2035_, ori_ori_n2036_, ori_ori_n2037_, ori_ori_n2038_, ori_ori_n2039_, ori_ori_n2040_, ori_ori_n2041_, ori_ori_n2042_, ori_ori_n2043_, ori_ori_n2044_, ori_ori_n2045_, ori_ori_n2046_, ori_ori_n2047_, ori_ori_n2048_, ori_ori_n2049_, ori_ori_n2050_, ori_ori_n2051_, ori_ori_n2052_, ori_ori_n2053_, ori_ori_n2054_, ori_ori_n2055_, ori_ori_n2056_, ori_ori_n2057_, ori_ori_n2058_, ori_ori_n2059_, ori_ori_n2060_, ori_ori_n2061_, ori_ori_n2062_, ori_ori_n2063_, ori_ori_n2064_, ori_ori_n2065_, ori_ori_n2066_, ori_ori_n2067_, ori_ori_n2068_, ori_ori_n2069_, ori_ori_n2070_, ori_ori_n2071_, ori_ori_n2072_, ori_ori_n2073_, ori_ori_n2074_, ori_ori_n2075_, ori_ori_n2076_, ori_ori_n2077_, ori_ori_n2078_, ori_ori_n2079_, ori_ori_n2081_, ori_ori_n2082_, ori_ori_n2083_, ori_ori_n2084_, ori_ori_n2085_, ori_ori_n2086_, ori_ori_n2087_, ori_ori_n2088_, ori_ori_n2089_, ori_ori_n2090_, ori_ori_n2091_, ori_ori_n2092_, ori_ori_n2093_, ori_ori_n2094_, ori_ori_n2095_, ori_ori_n2096_, ori_ori_n2097_, ori_ori_n2098_, ori_ori_n2099_, ori_ori_n2100_, ori_ori_n2101_, ori_ori_n2102_, ori_ori_n2103_, ori_ori_n2104_, ori_ori_n2105_, ori_ori_n2106_, ori_ori_n2107_, ori_ori_n2108_, ori_ori_n2109_, ori_ori_n2110_, ori_ori_n2111_, ori_ori_n2112_, ori_ori_n2113_, ori_ori_n2114_, ori_ori_n2115_, ori_ori_n2116_, ori_ori_n2117_, ori_ori_n2118_, ori_ori_n2119_, ori_ori_n2120_, ori_ori_n2121_, ori_ori_n2122_, ori_ori_n2123_, ori_ori_n2124_, ori_ori_n2125_, ori_ori_n2126_, ori_ori_n2127_, ori_ori_n2128_, ori_ori_n2129_, ori_ori_n2130_, ori_ori_n2131_, ori_ori_n2132_, ori_ori_n2133_, ori_ori_n2134_, ori_ori_n2135_, ori_ori_n2136_, ori_ori_n2137_, ori_ori_n2138_, ori_ori_n2139_, ori_ori_n2140_, ori_ori_n2141_, ori_ori_n2142_, ori_ori_n2143_, ori_ori_n2144_, ori_ori_n2146_, ori_ori_n2147_, ori_ori_n2148_, ori_ori_n2149_, ori_ori_n2150_, ori_ori_n2151_, ori_ori_n2152_, ori_ori_n2153_, ori_ori_n2154_, ori_ori_n2155_, ori_ori_n2156_, ori_ori_n2157_, ori_ori_n2158_, ori_ori_n2159_, ori_ori_n2160_, ori_ori_n2161_, ori_ori_n2162_, ori_ori_n2163_, ori_ori_n2164_, ori_ori_n2165_, ori_ori_n2166_, ori_ori_n2167_, ori_ori_n2168_, ori_ori_n2169_, ori_ori_n2170_, ori_ori_n2171_, ori_ori_n2172_, ori_ori_n2173_, ori_ori_n2174_, ori_ori_n2175_, ori_ori_n2176_, ori_ori_n2177_, ori_ori_n2178_, ori_ori_n2179_, ori_ori_n2180_, ori_ori_n2181_, ori_ori_n2182_, ori_ori_n2183_, ori_ori_n2184_, ori_ori_n2185_, ori_ori_n2186_, ori_ori_n2187_, ori_ori_n2188_, ori_ori_n2189_, ori_ori_n2190_, ori_ori_n2191_, ori_ori_n2192_, ori_ori_n2193_, ori_ori_n2194_, ori_ori_n2195_, ori_ori_n2196_, ori_ori_n2197_, ori_ori_n2198_, ori_ori_n2199_, ori_ori_n2200_, ori_ori_n2201_, ori_ori_n2202_, ori_ori_n2203_, ori_ori_n2204_, ori_ori_n2206_, ori_ori_n2207_, ori_ori_n2208_, ori_ori_n2209_, ori_ori_n2210_, ori_ori_n2211_, ori_ori_n2212_, ori_ori_n2213_, ori_ori_n2214_, ori_ori_n2215_, ori_ori_n2216_, ori_ori_n2217_, ori_ori_n2218_, ori_ori_n2219_, ori_ori_n2220_, ori_ori_n2221_, ori_ori_n2222_, ori_ori_n2223_, ori_ori_n2224_, ori_ori_n2225_, ori_ori_n2226_, ori_ori_n2227_, ori_ori_n2228_, ori_ori_n2229_, ori_ori_n2230_, ori_ori_n2231_, ori_ori_n2232_, ori_ori_n2233_, ori_ori_n2234_, ori_ori_n2235_, ori_ori_n2236_, ori_ori_n2237_, ori_ori_n2238_, ori_ori_n2239_, ori_ori_n2240_, ori_ori_n2241_, ori_ori_n2242_, ori_ori_n2243_, ori_ori_n2244_, ori_ori_n2245_, ori_ori_n2246_, ori_ori_n2247_, ori_ori_n2248_, ori_ori_n2249_, ori_ori_n2250_, ori_ori_n2251_, ori_ori_n2252_, ori_ori_n2253_, ori_ori_n2254_, ori_ori_n2255_, ori_ori_n2256_, ori_ori_n2257_, ori_ori_n2258_, ori_ori_n2259_, ori_ori_n2260_, ori_ori_n2261_, ori_ori_n2262_, ori_ori_n2263_, ori_ori_n2264_, ori_ori_n2265_, ori_ori_n2266_, ori_ori_n2267_, ori_ori_n2268_, ori_ori_n2269_, ori_ori_n2270_, ori_ori_n2271_, ori_ori_n2272_, ori_ori_n2273_, ori_ori_n2274_, ori_ori_n2276_, ori_ori_n2277_, ori_ori_n2278_, ori_ori_n2279_, ori_ori_n2280_, ori_ori_n2281_, ori_ori_n2282_, ori_ori_n2283_, ori_ori_n2284_, ori_ori_n2285_, ori_ori_n2286_, ori_ori_n2287_, ori_ori_n2288_, ori_ori_n2289_, ori_ori_n2290_, ori_ori_n2291_, ori_ori_n2292_, ori_ori_n2293_, ori_ori_n2294_, ori_ori_n2295_, ori_ori_n2296_, ori_ori_n2297_, ori_ori_n2298_, ori_ori_n2299_, ori_ori_n2300_, ori_ori_n2301_, ori_ori_n2302_, ori_ori_n2303_, ori_ori_n2304_, ori_ori_n2305_, ori_ori_n2306_, ori_ori_n2307_, ori_ori_n2308_, ori_ori_n2309_, ori_ori_n2310_, ori_ori_n2311_, ori_ori_n2312_, ori_ori_n2313_, ori_ori_n2314_, ori_ori_n2315_, ori_ori_n2316_, ori_ori_n2317_, ori_ori_n2318_, ori_ori_n2319_, ori_ori_n2320_, ori_ori_n2321_, ori_ori_n2322_, ori_ori_n2323_, ori_ori_n2324_, ori_ori_n2325_, ori_ori_n2326_, ori_ori_n2327_, ori_ori_n2328_, ori_ori_n2329_, ori_ori_n2330_, ori_ori_n2331_, ori_ori_n2332_, ori_ori_n2333_, ori_ori_n2334_, ori_ori_n2336_, ori_ori_n2337_, ori_ori_n2338_, ori_ori_n2339_, ori_ori_n2340_, ori_ori_n2341_, ori_ori_n2342_, ori_ori_n2343_, ori_ori_n2344_, ori_ori_n2345_, ori_ori_n2346_, ori_ori_n2347_, ori_ori_n2348_, ori_ori_n2349_, ori_ori_n2350_, ori_ori_n2351_, ori_ori_n2352_, ori_ori_n2353_, ori_ori_n2354_, ori_ori_n2355_, ori_ori_n2356_, ori_ori_n2357_, ori_ori_n2358_, ori_ori_n2359_, ori_ori_n2360_, ori_ori_n2361_, ori_ori_n2362_, ori_ori_n2363_, ori_ori_n2364_, ori_ori_n2365_, ori_ori_n2366_, ori_ori_n2367_, ori_ori_n2368_, ori_ori_n2369_, ori_ori_n2370_, ori_ori_n2371_, ori_ori_n2372_, ori_ori_n2373_, ori_ori_n2374_, ori_ori_n2375_, ori_ori_n2376_, ori_ori_n2377_, ori_ori_n2378_, ori_ori_n2379_, ori_ori_n2380_, ori_ori_n2381_, ori_ori_n2382_, ori_ori_n2383_, ori_ori_n2384_, ori_ori_n2385_, ori_ori_n2386_, ori_ori_n2387_, ori_ori_n2388_, ori_ori_n2389_, ori_ori_n2390_, ori_ori_n2391_, ori_ori_n2392_, ori_ori_n2393_, ori_ori_n2394_, ori_ori_n2395_, ori_ori_n2396_, ori_ori_n2397_, ori_ori_n2398_, ori_ori_n2399_, ori_ori_n2401_, ori_ori_n2402_, ori_ori_n2403_, ori_ori_n2404_, ori_ori_n2405_, ori_ori_n2406_, ori_ori_n2407_, ori_ori_n2408_, ori_ori_n2409_, ori_ori_n2410_, ori_ori_n2411_, ori_ori_n2412_, ori_ori_n2413_, ori_ori_n2414_, ori_ori_n2415_, ori_ori_n2416_, ori_ori_n2417_, ori_ori_n2418_, ori_ori_n2419_, ori_ori_n2420_, ori_ori_n2421_, ori_ori_n2422_, ori_ori_n2423_, ori_ori_n2424_, ori_ori_n2425_, ori_ori_n2426_, ori_ori_n2427_, ori_ori_n2428_, ori_ori_n2429_, ori_ori_n2430_, ori_ori_n2431_, ori_ori_n2432_, ori_ori_n2433_, ori_ori_n2434_, ori_ori_n2435_, ori_ori_n2436_, ori_ori_n2437_, ori_ori_n2438_, ori_ori_n2439_, ori_ori_n2440_, ori_ori_n2441_, ori_ori_n2442_, ori_ori_n2443_, ori_ori_n2444_, ori_ori_n2445_, ori_ori_n2446_, ori_ori_n2447_, ori_ori_n2448_, ori_ori_n2449_, ori_ori_n2450_, ori_ori_n2451_, ori_ori_n2452_, ori_ori_n2453_, ori_ori_n2454_, ori_ori_n2455_, ori_ori_n2456_, ori_ori_n2457_, ori_ori_n2458_, ori_ori_n2459_, ori_ori_n2460_, ori_ori_n2461_, ori_ori_n2462_, ori_ori_n2466_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1540_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1543_, mai_mai_n1544_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1549_, mai_mai_n1550_, mai_mai_n1551_, mai_mai_n1552_, mai_mai_n1553_, mai_mai_n1554_, mai_mai_n1555_, mai_mai_n1556_, mai_mai_n1557_, mai_mai_n1559_, mai_mai_n1560_, mai_mai_n1561_, mai_mai_n1562_, mai_mai_n1563_, mai_mai_n1564_, mai_mai_n1565_, mai_mai_n1566_, mai_mai_n1567_, mai_mai_n1568_, mai_mai_n1569_, mai_mai_n1570_, mai_mai_n1571_, mai_mai_n1572_, mai_mai_n1573_, mai_mai_n1574_, mai_mai_n1575_, mai_mai_n1576_, mai_mai_n1577_, mai_mai_n1578_, mai_mai_n1579_, mai_mai_n1580_, mai_mai_n1581_, mai_mai_n1582_, mai_mai_n1583_, mai_mai_n1584_, mai_mai_n1585_, mai_mai_n1586_, mai_mai_n1587_, mai_mai_n1588_, mai_mai_n1589_, mai_mai_n1590_, mai_mai_n1591_, mai_mai_n1592_, mai_mai_n1593_, mai_mai_n1594_, mai_mai_n1595_, mai_mai_n1596_, mai_mai_n1597_, mai_mai_n1598_, mai_mai_n1599_, mai_mai_n1600_, mai_mai_n1601_, mai_mai_n1602_, mai_mai_n1603_, mai_mai_n1604_, mai_mai_n1605_, mai_mai_n1606_, mai_mai_n1607_, mai_mai_n1608_, mai_mai_n1609_, mai_mai_n1610_, mai_mai_n1611_, mai_mai_n1612_, mai_mai_n1613_, mai_mai_n1614_, mai_mai_n1615_, mai_mai_n1616_, mai_mai_n1617_, mai_mai_n1618_, mai_mai_n1619_, mai_mai_n1620_, mai_mai_n1621_, mai_mai_n1622_, mai_mai_n1623_, mai_mai_n1624_, mai_mai_n1625_, mai_mai_n1626_, mai_mai_n1627_, mai_mai_n1628_, mai_mai_n1629_, mai_mai_n1630_, mai_mai_n1631_, mai_mai_n1632_, mai_mai_n1633_, mai_mai_n1634_, mai_mai_n1635_, mai_mai_n1636_, mai_mai_n1637_, mai_mai_n1638_, mai_mai_n1639_, mai_mai_n1640_, mai_mai_n1641_, mai_mai_n1642_, mai_mai_n1644_, mai_mai_n1645_, mai_mai_n1646_, mai_mai_n1647_, mai_mai_n1648_, mai_mai_n1649_, mai_mai_n1650_, mai_mai_n1651_, mai_mai_n1652_, mai_mai_n1653_, mai_mai_n1654_, mai_mai_n1655_, mai_mai_n1656_, mai_mai_n1657_, mai_mai_n1658_, mai_mai_n1659_, mai_mai_n1660_, mai_mai_n1661_, mai_mai_n1662_, mai_mai_n1663_, mai_mai_n1664_, mai_mai_n1665_, mai_mai_n1666_, mai_mai_n1667_, mai_mai_n1668_, mai_mai_n1669_, mai_mai_n1670_, mai_mai_n1671_, mai_mai_n1672_, mai_mai_n1673_, mai_mai_n1674_, mai_mai_n1675_, mai_mai_n1676_, mai_mai_n1677_, mai_mai_n1678_, mai_mai_n1679_, mai_mai_n1680_, mai_mai_n1681_, mai_mai_n1682_, mai_mai_n1683_, mai_mai_n1684_, mai_mai_n1685_, mai_mai_n1686_, mai_mai_n1687_, mai_mai_n1688_, mai_mai_n1689_, mai_mai_n1690_, mai_mai_n1691_, mai_mai_n1692_, mai_mai_n1693_, mai_mai_n1695_, mai_mai_n1696_, mai_mai_n1697_, mai_mai_n1698_, mai_mai_n1699_, mai_mai_n1700_, mai_mai_n1701_, mai_mai_n1702_, mai_mai_n1703_, mai_mai_n1704_, mai_mai_n1705_, mai_mai_n1706_, mai_mai_n1707_, mai_mai_n1708_, mai_mai_n1709_, mai_mai_n1710_, mai_mai_n1711_, mai_mai_n1712_, mai_mai_n1714_, mai_mai_n1715_, mai_mai_n1716_, mai_mai_n1717_, mai_mai_n1718_, mai_mai_n1719_, mai_mai_n1720_, mai_mai_n1721_, mai_mai_n1722_, mai_mai_n1723_, mai_mai_n1724_, mai_mai_n1725_, mai_mai_n1727_, mai_mai_n1728_, mai_mai_n1729_, mai_mai_n1730_, mai_mai_n1731_, mai_mai_n1732_, mai_mai_n1733_, mai_mai_n1734_, mai_mai_n1735_, mai_mai_n1736_, mai_mai_n1737_, mai_mai_n1738_, mai_mai_n1739_, mai_mai_n1740_, mai_mai_n1742_, mai_mai_n1743_, mai_mai_n1744_, mai_mai_n1745_, mai_mai_n1746_, mai_mai_n1747_, mai_mai_n1748_, mai_mai_n1749_, mai_mai_n1750_, mai_mai_n1751_, mai_mai_n1752_, mai_mai_n1753_, mai_mai_n1754_, mai_mai_n1755_, mai_mai_n1756_, mai_mai_n1757_, mai_mai_n1758_, mai_mai_n1759_, mai_mai_n1760_, mai_mai_n1761_, mai_mai_n1762_, mai_mai_n1763_, mai_mai_n1764_, mai_mai_n1765_, mai_mai_n1766_, mai_mai_n1767_, mai_mai_n1768_, mai_mai_n1769_, mai_mai_n1770_, mai_mai_n1771_, mai_mai_n1772_, mai_mai_n1773_, mai_mai_n1774_, mai_mai_n1775_, mai_mai_n1776_, mai_mai_n1777_, mai_mai_n1778_, mai_mai_n1779_, mai_mai_n1780_, mai_mai_n1781_, mai_mai_n1782_, mai_mai_n1783_, mai_mai_n1785_, mai_mai_n1786_, mai_mai_n1787_, mai_mai_n1788_, mai_mai_n1789_, mai_mai_n1790_, mai_mai_n1791_, mai_mai_n1792_, mai_mai_n1793_, mai_mai_n1794_, mai_mai_n1795_, mai_mai_n1796_, mai_mai_n1797_, mai_mai_n1799_, mai_mai_n1800_, mai_mai_n1801_, mai_mai_n1802_, mai_mai_n1803_, mai_mai_n1804_, mai_mai_n1805_, mai_mai_n1806_, mai_mai_n1807_, mai_mai_n1808_, mai_mai_n1809_, mai_mai_n1810_, mai_mai_n1811_, mai_mai_n1812_, mai_mai_n1813_, mai_mai_n1814_, mai_mai_n1815_, mai_mai_n1816_, mai_mai_n1817_, mai_mai_n1818_, mai_mai_n1819_, mai_mai_n1820_, mai_mai_n1821_, mai_mai_n1822_, mai_mai_n1823_, mai_mai_n1824_, mai_mai_n1825_, mai_mai_n1826_, mai_mai_n1827_, mai_mai_n1828_, mai_mai_n1829_, mai_mai_n1830_, mai_mai_n1831_, mai_mai_n1832_, mai_mai_n1833_, mai_mai_n1834_, mai_mai_n1835_, mai_mai_n1836_, mai_mai_n1837_, mai_mai_n1838_, mai_mai_n1839_, mai_mai_n1840_, mai_mai_n1841_, mai_mai_n1842_, mai_mai_n1843_, mai_mai_n1844_, mai_mai_n1846_, mai_mai_n1847_, mai_mai_n1848_, mai_mai_n1849_, mai_mai_n1850_, mai_mai_n1851_, mai_mai_n1852_, mai_mai_n1853_, mai_mai_n1854_, mai_mai_n1855_, mai_mai_n1856_, mai_mai_n1857_, mai_mai_n1858_, mai_mai_n1859_, mai_mai_n1860_, mai_mai_n1861_, mai_mai_n1862_, mai_mai_n1863_, mai_mai_n1864_, mai_mai_n1865_, mai_mai_n1866_, mai_mai_n1867_, mai_mai_n1868_, mai_mai_n1869_, mai_mai_n1870_, mai_mai_n1871_, mai_mai_n1872_, mai_mai_n1873_, mai_mai_n1874_, mai_mai_n1875_, mai_mai_n1876_, mai_mai_n1877_, mai_mai_n1878_, mai_mai_n1879_, mai_mai_n1880_, mai_mai_n1881_, mai_mai_n1882_, mai_mai_n1883_, mai_mai_n1884_, mai_mai_n1885_, mai_mai_n1886_, mai_mai_n1887_, mai_mai_n1888_, mai_mai_n1889_, mai_mai_n1890_, mai_mai_n1891_, mai_mai_n1892_, mai_mai_n1893_, mai_mai_n1894_, mai_mai_n1895_, mai_mai_n1896_, mai_mai_n1897_, mai_mai_n1898_, mai_mai_n1899_, mai_mai_n1900_, mai_mai_n1901_, mai_mai_n1902_, mai_mai_n1903_, mai_mai_n1904_, mai_mai_n1906_, mai_mai_n1907_, mai_mai_n1908_, mai_mai_n1909_, mai_mai_n1910_, mai_mai_n1911_, mai_mai_n1912_, mai_mai_n1913_, mai_mai_n1914_, mai_mai_n1915_, mai_mai_n1916_, mai_mai_n1917_, mai_mai_n1918_, mai_mai_n1919_, mai_mai_n1920_, mai_mai_n1921_, mai_mai_n1922_, mai_mai_n1923_, mai_mai_n1924_, mai_mai_n1925_, mai_mai_n1926_, mai_mai_n1927_, mai_mai_n1928_, mai_mai_n1929_, mai_mai_n1930_, mai_mai_n1931_, mai_mai_n1932_, mai_mai_n1933_, mai_mai_n1934_, mai_mai_n1935_, mai_mai_n1936_, mai_mai_n1937_, mai_mai_n1938_, mai_mai_n1939_, mai_mai_n1940_, mai_mai_n1941_, mai_mai_n1942_, mai_mai_n1943_, mai_mai_n1944_, mai_mai_n1945_, mai_mai_n1946_, mai_mai_n1947_, mai_mai_n1948_, mai_mai_n1949_, mai_mai_n1950_, mai_mai_n1951_, mai_mai_n1952_, mai_mai_n1953_, mai_mai_n1954_, mai_mai_n1955_, mai_mai_n1956_, mai_mai_n1957_, mai_mai_n1958_, mai_mai_n1959_, mai_mai_n1960_, mai_mai_n1961_, mai_mai_n1962_, mai_mai_n1963_, mai_mai_n1964_, mai_mai_n1965_, mai_mai_n1966_, mai_mai_n1967_, mai_mai_n1968_, mai_mai_n1969_, mai_mai_n1970_, mai_mai_n1971_, mai_mai_n1972_, mai_mai_n1973_, mai_mai_n1974_, mai_mai_n1975_, mai_mai_n1976_, mai_mai_n1978_, mai_mai_n1979_, mai_mai_n1980_, mai_mai_n1981_, mai_mai_n1982_, mai_mai_n1983_, mai_mai_n1984_, mai_mai_n1985_, mai_mai_n1986_, mai_mai_n1987_, mai_mai_n1988_, mai_mai_n1989_, mai_mai_n1990_, mai_mai_n1991_, mai_mai_n1992_, mai_mai_n1993_, mai_mai_n1994_, mai_mai_n1995_, mai_mai_n1996_, mai_mai_n1997_, mai_mai_n1998_, mai_mai_n1999_, mai_mai_n2000_, mai_mai_n2001_, mai_mai_n2002_, mai_mai_n2003_, mai_mai_n2004_, mai_mai_n2005_, mai_mai_n2006_, mai_mai_n2007_, mai_mai_n2008_, mai_mai_n2009_, mai_mai_n2010_, mai_mai_n2011_, mai_mai_n2012_, mai_mai_n2013_, mai_mai_n2014_, mai_mai_n2015_, mai_mai_n2016_, mai_mai_n2017_, mai_mai_n2018_, mai_mai_n2019_, mai_mai_n2020_, mai_mai_n2021_, mai_mai_n2022_, mai_mai_n2023_, mai_mai_n2024_, mai_mai_n2025_, mai_mai_n2026_, mai_mai_n2027_, mai_mai_n2028_, mai_mai_n2029_, mai_mai_n2030_, mai_mai_n2031_, mai_mai_n2032_, mai_mai_n2033_, mai_mai_n2034_, mai_mai_n2035_, mai_mai_n2036_, mai_mai_n2037_, mai_mai_n2038_, mai_mai_n2039_, mai_mai_n2040_, mai_mai_n2041_, mai_mai_n2042_, mai_mai_n2043_, mai_mai_n2044_, mai_mai_n2045_, mai_mai_n2047_, mai_mai_n2048_, mai_mai_n2049_, mai_mai_n2050_, mai_mai_n2051_, mai_mai_n2052_, mai_mai_n2053_, mai_mai_n2054_, mai_mai_n2055_, mai_mai_n2056_, mai_mai_n2057_, mai_mai_n2058_, mai_mai_n2059_, mai_mai_n2060_, mai_mai_n2061_, mai_mai_n2062_, mai_mai_n2063_, mai_mai_n2064_, mai_mai_n2065_, mai_mai_n2066_, mai_mai_n2067_, mai_mai_n2068_, mai_mai_n2069_, mai_mai_n2070_, mai_mai_n2071_, mai_mai_n2072_, mai_mai_n2073_, mai_mai_n2074_, mai_mai_n2075_, mai_mai_n2076_, mai_mai_n2077_, mai_mai_n2078_, mai_mai_n2079_, mai_mai_n2080_, mai_mai_n2081_, mai_mai_n2082_, mai_mai_n2083_, mai_mai_n2084_, mai_mai_n2085_, mai_mai_n2086_, mai_mai_n2087_, mai_mai_n2088_, mai_mai_n2089_, mai_mai_n2090_, mai_mai_n2091_, mai_mai_n2092_, mai_mai_n2093_, mai_mai_n2094_, mai_mai_n2095_, mai_mai_n2096_, mai_mai_n2097_, mai_mai_n2098_, mai_mai_n2099_, mai_mai_n2100_, mai_mai_n2101_, mai_mai_n2102_, mai_mai_n2103_, mai_mai_n2104_, mai_mai_n2105_, mai_mai_n2106_, mai_mai_n2107_, mai_mai_n2108_, mai_mai_n2109_, mai_mai_n2110_, mai_mai_n2111_, mai_mai_n2112_, mai_mai_n2113_, mai_mai_n2114_, mai_mai_n2115_, mai_mai_n2116_, mai_mai_n2117_, mai_mai_n2118_, mai_mai_n2120_, mai_mai_n2121_, mai_mai_n2122_, mai_mai_n2123_, mai_mai_n2124_, mai_mai_n2125_, mai_mai_n2126_, mai_mai_n2127_, mai_mai_n2128_, mai_mai_n2129_, mai_mai_n2130_, mai_mai_n2131_, mai_mai_n2132_, mai_mai_n2133_, mai_mai_n2134_, mai_mai_n2135_, mai_mai_n2136_, mai_mai_n2137_, mai_mai_n2138_, mai_mai_n2139_, mai_mai_n2140_, mai_mai_n2141_, mai_mai_n2142_, mai_mai_n2143_, mai_mai_n2144_, mai_mai_n2145_, mai_mai_n2146_, mai_mai_n2147_, mai_mai_n2148_, mai_mai_n2149_, mai_mai_n2150_, mai_mai_n2151_, mai_mai_n2152_, mai_mai_n2153_, mai_mai_n2154_, mai_mai_n2155_, mai_mai_n2156_, mai_mai_n2157_, mai_mai_n2158_, mai_mai_n2159_, mai_mai_n2160_, mai_mai_n2161_, mai_mai_n2162_, mai_mai_n2163_, mai_mai_n2164_, mai_mai_n2165_, mai_mai_n2166_, mai_mai_n2167_, mai_mai_n2168_, mai_mai_n2169_, mai_mai_n2170_, mai_mai_n2171_, mai_mai_n2172_, mai_mai_n2173_, mai_mai_n2174_, mai_mai_n2175_, mai_mai_n2176_, mai_mai_n2177_, mai_mai_n2178_, mai_mai_n2179_, mai_mai_n2180_, mai_mai_n2181_, mai_mai_n2182_, mai_mai_n2184_, mai_mai_n2185_, mai_mai_n2186_, mai_mai_n2187_, mai_mai_n2188_, mai_mai_n2189_, mai_mai_n2190_, mai_mai_n2191_, mai_mai_n2192_, mai_mai_n2193_, mai_mai_n2194_, mai_mai_n2195_, mai_mai_n2196_, mai_mai_n2197_, mai_mai_n2198_, mai_mai_n2199_, mai_mai_n2200_, mai_mai_n2201_, mai_mai_n2202_, mai_mai_n2203_, mai_mai_n2204_, mai_mai_n2205_, mai_mai_n2206_, mai_mai_n2207_, mai_mai_n2208_, mai_mai_n2209_, mai_mai_n2210_, mai_mai_n2211_, mai_mai_n2212_, mai_mai_n2213_, mai_mai_n2214_, mai_mai_n2215_, mai_mai_n2216_, mai_mai_n2217_, mai_mai_n2218_, mai_mai_n2219_, mai_mai_n2220_, mai_mai_n2221_, mai_mai_n2222_, mai_mai_n2223_, mai_mai_n2224_, mai_mai_n2225_, mai_mai_n2226_, mai_mai_n2227_, mai_mai_n2228_, mai_mai_n2229_, mai_mai_n2230_, mai_mai_n2231_, mai_mai_n2232_, mai_mai_n2233_, mai_mai_n2234_, mai_mai_n2235_, mai_mai_n2236_, mai_mai_n2237_, mai_mai_n2238_, mai_mai_n2239_, mai_mai_n2241_, mai_mai_n2242_, mai_mai_n2243_, mai_mai_n2244_, mai_mai_n2245_, mai_mai_n2246_, mai_mai_n2247_, mai_mai_n2248_, mai_mai_n2249_, mai_mai_n2250_, mai_mai_n2251_, mai_mai_n2252_, mai_mai_n2253_, mai_mai_n2254_, mai_mai_n2255_, mai_mai_n2256_, mai_mai_n2257_, mai_mai_n2258_, mai_mai_n2259_, mai_mai_n2260_, mai_mai_n2261_, mai_mai_n2262_, mai_mai_n2263_, mai_mai_n2264_, mai_mai_n2265_, mai_mai_n2266_, mai_mai_n2267_, mai_mai_n2268_, mai_mai_n2269_, mai_mai_n2270_, mai_mai_n2271_, mai_mai_n2272_, mai_mai_n2273_, mai_mai_n2274_, mai_mai_n2275_, mai_mai_n2276_, mai_mai_n2277_, mai_mai_n2278_, mai_mai_n2279_, mai_mai_n2280_, mai_mai_n2281_, mai_mai_n2282_, mai_mai_n2283_, mai_mai_n2284_, mai_mai_n2285_, mai_mai_n2286_, mai_mai_n2287_, mai_mai_n2288_, mai_mai_n2289_, mai_mai_n2290_, mai_mai_n2291_, mai_mai_n2292_, mai_mai_n2293_, mai_mai_n2294_, mai_mai_n2295_, mai_mai_n2296_, mai_mai_n2297_, mai_mai_n2298_, mai_mai_n2299_, mai_mai_n2300_, mai_mai_n2301_, mai_mai_n2302_, mai_mai_n2303_, mai_mai_n2304_, mai_mai_n2305_, mai_mai_n2306_, mai_mai_n2307_, mai_mai_n2308_, mai_mai_n2309_, mai_mai_n2310_, mai_mai_n2311_, mai_mai_n2312_, mai_mai_n2313_, mai_mai_n2315_, mai_mai_n2316_, mai_mai_n2317_, mai_mai_n2318_, mai_mai_n2319_, mai_mai_n2320_, mai_mai_n2321_, mai_mai_n2322_, mai_mai_n2323_, mai_mai_n2324_, mai_mai_n2325_, mai_mai_n2326_, mai_mai_n2327_, mai_mai_n2328_, mai_mai_n2329_, mai_mai_n2330_, mai_mai_n2331_, mai_mai_n2332_, mai_mai_n2333_, mai_mai_n2334_, mai_mai_n2335_, mai_mai_n2336_, mai_mai_n2337_, mai_mai_n2338_, mai_mai_n2339_, mai_mai_n2340_, mai_mai_n2341_, mai_mai_n2342_, mai_mai_n2343_, mai_mai_n2344_, mai_mai_n2345_, mai_mai_n2346_, mai_mai_n2347_, mai_mai_n2348_, mai_mai_n2349_, mai_mai_n2350_, mai_mai_n2351_, mai_mai_n2352_, mai_mai_n2353_, mai_mai_n2354_, mai_mai_n2355_, mai_mai_n2356_, mai_mai_n2357_, mai_mai_n2358_, mai_mai_n2359_, mai_mai_n2360_, mai_mai_n2361_, mai_mai_n2362_, mai_mai_n2363_, mai_mai_n2364_, mai_mai_n2365_, mai_mai_n2366_, mai_mai_n2367_, mai_mai_n2368_, mai_mai_n2369_, mai_mai_n2370_, mai_mai_n2371_, mai_mai_n2372_, mai_mai_n2373_, mai_mai_n2374_, mai_mai_n2375_, mai_mai_n2376_, mai_mai_n2377_, mai_mai_n2379_, mai_mai_n2380_, mai_mai_n2381_, mai_mai_n2382_, mai_mai_n2383_, mai_mai_n2384_, mai_mai_n2385_, mai_mai_n2386_, mai_mai_n2387_, mai_mai_n2388_, mai_mai_n2389_, mai_mai_n2390_, mai_mai_n2391_, mai_mai_n2392_, mai_mai_n2393_, mai_mai_n2394_, mai_mai_n2395_, mai_mai_n2396_, mai_mai_n2397_, mai_mai_n2398_, mai_mai_n2399_, mai_mai_n2400_, mai_mai_n2401_, mai_mai_n2402_, mai_mai_n2403_, mai_mai_n2404_, mai_mai_n2405_, mai_mai_n2406_, mai_mai_n2407_, mai_mai_n2408_, mai_mai_n2409_, mai_mai_n2410_, mai_mai_n2411_, mai_mai_n2412_, mai_mai_n2413_, mai_mai_n2414_, mai_mai_n2415_, mai_mai_n2416_, mai_mai_n2417_, mai_mai_n2418_, mai_mai_n2419_, mai_mai_n2420_, mai_mai_n2421_, mai_mai_n2422_, mai_mai_n2423_, mai_mai_n2424_, mai_mai_n2425_, mai_mai_n2426_, mai_mai_n2427_, mai_mai_n2428_, mai_mai_n2429_, mai_mai_n2430_, mai_mai_n2431_, mai_mai_n2432_, mai_mai_n2433_, mai_mai_n2434_, mai_mai_n2435_, mai_mai_n2436_, mai_mai_n2437_, mai_mai_n2438_, mai_mai_n2439_, mai_mai_n2440_, mai_mai_n2441_, mai_mai_n2442_, mai_mai_n2444_, mai_mai_n2445_, mai_mai_n2446_, mai_mai_n2447_, mai_mai_n2448_, mai_mai_n2449_, mai_mai_n2450_, mai_mai_n2451_, mai_mai_n2452_, mai_mai_n2453_, mai_mai_n2454_, mai_mai_n2455_, mai_mai_n2456_, mai_mai_n2457_, mai_mai_n2458_, mai_mai_n2459_, mai_mai_n2460_, mai_mai_n2461_, mai_mai_n2462_, mai_mai_n2463_, mai_mai_n2464_, mai_mai_n2465_, mai_mai_n2466_, mai_mai_n2467_, mai_mai_n2468_, mai_mai_n2469_, mai_mai_n2470_, mai_mai_n2471_, mai_mai_n2472_, mai_mai_n2473_, mai_mai_n2474_, mai_mai_n2475_, mai_mai_n2476_, mai_mai_n2477_, mai_mai_n2478_, mai_mai_n2479_, mai_mai_n2480_, mai_mai_n2481_, mai_mai_n2482_, mai_mai_n2483_, mai_mai_n2484_, mai_mai_n2485_, mai_mai_n2486_, mai_mai_n2487_, mai_mai_n2488_, mai_mai_n2489_, mai_mai_n2490_, mai_mai_n2491_, mai_mai_n2492_, mai_mai_n2493_, mai_mai_n2494_, mai_mai_n2495_, mai_mai_n2496_, mai_mai_n2497_, mai_mai_n2498_, mai_mai_n2499_, mai_mai_n2500_, mai_mai_n2501_, mai_mai_n2502_, mai_mai_n2503_, mai_mai_n2504_, mai_mai_n2505_, mai_mai_n2506_, mai_mai_n2510_, mai_mai_n2511_, mai_mai_n2512_, mai_mai_n2513_, mai_mai_n2514_, mai_mai_n2515_, mai_mai_n2516_, mai_mai_n2517_, mai_mai_n2518_, mai_mai_n2519_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1606_, men_men_n1607_, men_men_n1608_, men_men_n1609_, men_men_n1610_, men_men_n1611_, men_men_n1612_, men_men_n1613_, men_men_n1614_, men_men_n1615_, men_men_n1616_, men_men_n1617_, men_men_n1618_, men_men_n1619_, men_men_n1620_, men_men_n1621_, men_men_n1622_, men_men_n1623_, men_men_n1624_, men_men_n1625_, men_men_n1626_, men_men_n1627_, men_men_n1628_, men_men_n1629_, men_men_n1630_, men_men_n1631_, men_men_n1632_, men_men_n1633_, men_men_n1634_, men_men_n1635_, men_men_n1636_, men_men_n1637_, men_men_n1638_, men_men_n1639_, men_men_n1640_, men_men_n1641_, men_men_n1642_, men_men_n1643_, men_men_n1644_, men_men_n1645_, men_men_n1646_, men_men_n1647_, men_men_n1648_, men_men_n1649_, men_men_n1650_, men_men_n1651_, men_men_n1652_, men_men_n1653_, men_men_n1654_, men_men_n1655_, men_men_n1656_, men_men_n1657_, men_men_n1658_, men_men_n1659_, men_men_n1660_, men_men_n1661_, men_men_n1662_, men_men_n1663_, men_men_n1664_, men_men_n1665_, men_men_n1666_, men_men_n1667_, men_men_n1668_, men_men_n1669_, men_men_n1670_, men_men_n1671_, men_men_n1672_, men_men_n1674_, men_men_n1675_, men_men_n1676_, men_men_n1677_, men_men_n1678_, men_men_n1679_, men_men_n1680_, men_men_n1681_, men_men_n1682_, men_men_n1683_, men_men_n1684_, men_men_n1685_, men_men_n1686_, men_men_n1687_, men_men_n1688_, men_men_n1689_, men_men_n1690_, men_men_n1691_, men_men_n1692_, men_men_n1693_, men_men_n1694_, men_men_n1695_, men_men_n1696_, men_men_n1697_, men_men_n1698_, men_men_n1699_, men_men_n1700_, men_men_n1701_, men_men_n1702_, men_men_n1703_, men_men_n1704_, men_men_n1705_, men_men_n1706_, men_men_n1707_, men_men_n1708_, men_men_n1709_, men_men_n1710_, men_men_n1711_, men_men_n1712_, men_men_n1713_, men_men_n1714_, men_men_n1715_, men_men_n1716_, men_men_n1717_, men_men_n1718_, men_men_n1719_, men_men_n1720_, men_men_n1721_, men_men_n1722_, men_men_n1723_, men_men_n1724_, men_men_n1725_, men_men_n1726_, men_men_n1727_, men_men_n1728_, men_men_n1729_, men_men_n1731_, men_men_n1732_, men_men_n1733_, men_men_n1734_, men_men_n1735_, men_men_n1736_, men_men_n1737_, men_men_n1738_, men_men_n1739_, men_men_n1740_, men_men_n1741_, men_men_n1742_, men_men_n1743_, men_men_n1744_, men_men_n1745_, men_men_n1746_, men_men_n1747_, men_men_n1748_, men_men_n1750_, men_men_n1751_, men_men_n1752_, men_men_n1753_, men_men_n1754_, men_men_n1755_, men_men_n1756_, men_men_n1757_, men_men_n1758_, men_men_n1759_, men_men_n1760_, men_men_n1761_, men_men_n1762_, men_men_n1764_, men_men_n1765_, men_men_n1766_, men_men_n1767_, men_men_n1768_, men_men_n1769_, men_men_n1770_, men_men_n1771_, men_men_n1772_, men_men_n1773_, men_men_n1774_, men_men_n1775_, men_men_n1776_, men_men_n1777_, men_men_n1778_, men_men_n1779_, men_men_n1780_, men_men_n1782_, men_men_n1783_, men_men_n1784_, men_men_n1785_, men_men_n1786_, men_men_n1787_, men_men_n1788_, men_men_n1789_, men_men_n1790_, men_men_n1791_, men_men_n1792_, men_men_n1793_, men_men_n1794_, men_men_n1795_, men_men_n1796_, men_men_n1797_, men_men_n1798_, men_men_n1799_, men_men_n1800_, men_men_n1801_, men_men_n1802_, men_men_n1803_, men_men_n1804_, men_men_n1805_, men_men_n1806_, men_men_n1807_, men_men_n1808_, men_men_n1809_, men_men_n1810_, men_men_n1811_, men_men_n1812_, men_men_n1813_, men_men_n1814_, men_men_n1815_, men_men_n1816_, men_men_n1817_, men_men_n1818_, men_men_n1819_, men_men_n1820_, men_men_n1821_, men_men_n1822_, men_men_n1823_, men_men_n1824_, men_men_n1825_, men_men_n1827_, men_men_n1828_, men_men_n1829_, men_men_n1830_, men_men_n1831_, men_men_n1832_, men_men_n1833_, men_men_n1834_, men_men_n1835_, men_men_n1836_, men_men_n1837_, men_men_n1838_, men_men_n1839_, men_men_n1840_, men_men_n1842_, men_men_n1843_, men_men_n1844_, men_men_n1845_, men_men_n1846_, men_men_n1847_, men_men_n1848_, men_men_n1849_, men_men_n1850_, men_men_n1851_, men_men_n1852_, men_men_n1853_, men_men_n1854_, men_men_n1855_, men_men_n1856_, men_men_n1857_, men_men_n1858_, men_men_n1859_, men_men_n1860_, men_men_n1861_, men_men_n1862_, men_men_n1863_, men_men_n1864_, men_men_n1865_, men_men_n1866_, men_men_n1867_, men_men_n1868_, men_men_n1869_, men_men_n1870_, men_men_n1871_, men_men_n1872_, men_men_n1873_, men_men_n1874_, men_men_n1875_, men_men_n1876_, men_men_n1877_, men_men_n1878_, men_men_n1879_, men_men_n1880_, men_men_n1881_, men_men_n1882_, men_men_n1883_, men_men_n1884_, men_men_n1885_, men_men_n1886_, men_men_n1887_, men_men_n1888_, men_men_n1889_, men_men_n1890_, men_men_n1892_, men_men_n1893_, men_men_n1894_, men_men_n1895_, men_men_n1896_, men_men_n1897_, men_men_n1898_, men_men_n1899_, men_men_n1900_, men_men_n1901_, men_men_n1902_, men_men_n1903_, men_men_n1904_, men_men_n1905_, men_men_n1906_, men_men_n1907_, men_men_n1908_, men_men_n1909_, men_men_n1910_, men_men_n1911_, men_men_n1912_, men_men_n1913_, men_men_n1914_, men_men_n1915_, men_men_n1916_, men_men_n1917_, men_men_n1918_, men_men_n1919_, men_men_n1920_, men_men_n1921_, men_men_n1922_, men_men_n1923_, men_men_n1924_, men_men_n1925_, men_men_n1926_, men_men_n1927_, men_men_n1928_, men_men_n1929_, men_men_n1930_, men_men_n1931_, men_men_n1932_, men_men_n1933_, men_men_n1934_, men_men_n1935_, men_men_n1936_, men_men_n1937_, men_men_n1938_, men_men_n1939_, men_men_n1940_, men_men_n1941_, men_men_n1942_, men_men_n1943_, men_men_n1944_, men_men_n1945_, men_men_n1946_, men_men_n1947_, men_men_n1948_, men_men_n1949_, men_men_n1950_, men_men_n1951_, men_men_n1953_, men_men_n1954_, men_men_n1955_, men_men_n1956_, men_men_n1957_, men_men_n1958_, men_men_n1959_, men_men_n1960_, men_men_n1961_, men_men_n1962_, men_men_n1963_, men_men_n1964_, men_men_n1965_, men_men_n1966_, men_men_n1967_, men_men_n1968_, men_men_n1969_, men_men_n1970_, men_men_n1971_, men_men_n1972_, men_men_n1973_, men_men_n1974_, men_men_n1975_, men_men_n1976_, men_men_n1977_, men_men_n1978_, men_men_n1979_, men_men_n1980_, men_men_n1981_, men_men_n1982_, men_men_n1983_, men_men_n1984_, men_men_n1985_, men_men_n1986_, men_men_n1987_, men_men_n1988_, men_men_n1989_, men_men_n1990_, men_men_n1991_, men_men_n1992_, men_men_n1993_, men_men_n1994_, men_men_n1995_, men_men_n1996_, men_men_n1997_, men_men_n1998_, men_men_n1999_, men_men_n2000_, men_men_n2001_, men_men_n2002_, men_men_n2003_, men_men_n2004_, men_men_n2005_, men_men_n2006_, men_men_n2007_, men_men_n2008_, men_men_n2009_, men_men_n2010_, men_men_n2011_, men_men_n2012_, men_men_n2013_, men_men_n2014_, men_men_n2015_, men_men_n2016_, men_men_n2017_, men_men_n2018_, men_men_n2019_, men_men_n2020_, men_men_n2021_, men_men_n2022_, men_men_n2023_, men_men_n2024_, men_men_n2025_, men_men_n2026_, men_men_n2027_, men_men_n2029_, men_men_n2030_, men_men_n2031_, men_men_n2032_, men_men_n2033_, men_men_n2034_, men_men_n2035_, men_men_n2036_, men_men_n2037_, men_men_n2038_, men_men_n2039_, men_men_n2040_, men_men_n2041_, men_men_n2042_, men_men_n2043_, men_men_n2044_, men_men_n2045_, men_men_n2046_, men_men_n2047_, men_men_n2048_, men_men_n2049_, men_men_n2050_, men_men_n2051_, men_men_n2052_, men_men_n2053_, men_men_n2054_, men_men_n2055_, men_men_n2056_, men_men_n2057_, men_men_n2058_, men_men_n2059_, men_men_n2060_, men_men_n2061_, men_men_n2062_, men_men_n2063_, men_men_n2064_, men_men_n2065_, men_men_n2066_, men_men_n2067_, men_men_n2068_, men_men_n2069_, men_men_n2070_, men_men_n2071_, men_men_n2072_, men_men_n2073_, men_men_n2074_, men_men_n2075_, men_men_n2076_, men_men_n2077_, men_men_n2078_, men_men_n2079_, men_men_n2080_, men_men_n2081_, men_men_n2082_, men_men_n2083_, men_men_n2084_, men_men_n2085_, men_men_n2086_, men_men_n2087_, men_men_n2088_, men_men_n2089_, men_men_n2090_, men_men_n2091_, men_men_n2092_, men_men_n2093_, men_men_n2094_, men_men_n2095_, men_men_n2096_, men_men_n2097_, men_men_n2098_, men_men_n2100_, men_men_n2101_, men_men_n2102_, men_men_n2103_, men_men_n2104_, men_men_n2105_, men_men_n2106_, men_men_n2107_, men_men_n2108_, men_men_n2109_, men_men_n2110_, men_men_n2111_, men_men_n2112_, men_men_n2113_, men_men_n2114_, men_men_n2115_, men_men_n2116_, men_men_n2117_, men_men_n2118_, men_men_n2119_, men_men_n2120_, men_men_n2121_, men_men_n2122_, men_men_n2123_, men_men_n2124_, men_men_n2125_, men_men_n2126_, men_men_n2127_, men_men_n2128_, men_men_n2129_, men_men_n2130_, men_men_n2131_, men_men_n2132_, men_men_n2133_, men_men_n2134_, men_men_n2135_, men_men_n2136_, men_men_n2137_, men_men_n2138_, men_men_n2139_, men_men_n2140_, men_men_n2141_, men_men_n2142_, men_men_n2143_, men_men_n2144_, men_men_n2145_, men_men_n2146_, men_men_n2147_, men_men_n2148_, men_men_n2149_, men_men_n2150_, men_men_n2151_, men_men_n2152_, men_men_n2153_, men_men_n2154_, men_men_n2155_, men_men_n2156_, men_men_n2157_, men_men_n2158_, men_men_n2159_, men_men_n2160_, men_men_n2161_, men_men_n2162_, men_men_n2163_, men_men_n2164_, men_men_n2165_, men_men_n2166_, men_men_n2167_, men_men_n2168_, men_men_n2169_, men_men_n2171_, men_men_n2172_, men_men_n2173_, men_men_n2174_, men_men_n2175_, men_men_n2176_, men_men_n2177_, men_men_n2178_, men_men_n2179_, men_men_n2180_, men_men_n2181_, men_men_n2182_, men_men_n2183_, men_men_n2184_, men_men_n2185_, men_men_n2186_, men_men_n2187_, men_men_n2188_, men_men_n2189_, men_men_n2190_, men_men_n2191_, men_men_n2192_, men_men_n2193_, men_men_n2194_, men_men_n2195_, men_men_n2196_, men_men_n2197_, men_men_n2198_, men_men_n2199_, men_men_n2200_, men_men_n2201_, men_men_n2202_, men_men_n2203_, men_men_n2204_, men_men_n2205_, men_men_n2206_, men_men_n2207_, men_men_n2208_, men_men_n2209_, men_men_n2210_, men_men_n2211_, men_men_n2212_, men_men_n2213_, men_men_n2214_, men_men_n2215_, men_men_n2216_, men_men_n2217_, men_men_n2218_, men_men_n2219_, men_men_n2220_, men_men_n2221_, men_men_n2222_, men_men_n2223_, men_men_n2224_, men_men_n2225_, men_men_n2226_, men_men_n2227_, men_men_n2228_, men_men_n2229_, men_men_n2230_, men_men_n2231_, men_men_n2232_, men_men_n2233_, men_men_n2234_, men_men_n2235_, men_men_n2237_, men_men_n2238_, men_men_n2239_, men_men_n2240_, men_men_n2241_, men_men_n2242_, men_men_n2243_, men_men_n2244_, men_men_n2245_, men_men_n2246_, men_men_n2247_, men_men_n2248_, men_men_n2249_, men_men_n2250_, men_men_n2251_, men_men_n2252_, men_men_n2253_, men_men_n2254_, men_men_n2255_, men_men_n2256_, men_men_n2257_, men_men_n2258_, men_men_n2259_, men_men_n2260_, men_men_n2261_, men_men_n2262_, men_men_n2263_, men_men_n2264_, men_men_n2265_, men_men_n2266_, men_men_n2267_, men_men_n2268_, men_men_n2269_, men_men_n2270_, men_men_n2271_, men_men_n2272_, men_men_n2273_, men_men_n2274_, men_men_n2275_, men_men_n2276_, men_men_n2277_, men_men_n2278_, men_men_n2279_, men_men_n2280_, men_men_n2281_, men_men_n2282_, men_men_n2283_, men_men_n2284_, men_men_n2285_, men_men_n2286_, men_men_n2287_, men_men_n2288_, men_men_n2289_, men_men_n2290_, men_men_n2292_, men_men_n2293_, men_men_n2294_, men_men_n2295_, men_men_n2296_, men_men_n2297_, men_men_n2298_, men_men_n2299_, men_men_n2300_, men_men_n2301_, men_men_n2302_, men_men_n2303_, men_men_n2304_, men_men_n2305_, men_men_n2306_, men_men_n2307_, men_men_n2308_, men_men_n2309_, men_men_n2310_, men_men_n2311_, men_men_n2312_, men_men_n2313_, men_men_n2314_, men_men_n2315_, men_men_n2316_, men_men_n2317_, men_men_n2318_, men_men_n2319_, men_men_n2320_, men_men_n2321_, men_men_n2322_, men_men_n2323_, men_men_n2324_, men_men_n2325_, men_men_n2326_, men_men_n2327_, men_men_n2328_, men_men_n2329_, men_men_n2330_, men_men_n2331_, men_men_n2332_, men_men_n2333_, men_men_n2334_, men_men_n2335_, men_men_n2336_, men_men_n2337_, men_men_n2338_, men_men_n2339_, men_men_n2340_, men_men_n2341_, men_men_n2342_, men_men_n2343_, men_men_n2344_, men_men_n2345_, men_men_n2346_, men_men_n2347_, men_men_n2348_, men_men_n2349_, men_men_n2350_, men_men_n2351_, men_men_n2352_, men_men_n2353_, men_men_n2354_, men_men_n2355_, men_men_n2356_, men_men_n2357_, men_men_n2358_, men_men_n2359_, men_men_n2360_, men_men_n2361_, men_men_n2362_, men_men_n2363_, men_men_n2364_, men_men_n2366_, men_men_n2367_, men_men_n2368_, men_men_n2369_, men_men_n2370_, men_men_n2371_, men_men_n2372_, men_men_n2373_, men_men_n2374_, men_men_n2375_, men_men_n2376_, men_men_n2377_, men_men_n2378_, men_men_n2379_, men_men_n2380_, men_men_n2381_, men_men_n2382_, men_men_n2383_, men_men_n2384_, men_men_n2385_, men_men_n2386_, men_men_n2387_, men_men_n2388_, men_men_n2389_, men_men_n2390_, men_men_n2391_, men_men_n2392_, men_men_n2393_, men_men_n2394_, men_men_n2395_, men_men_n2396_, men_men_n2397_, men_men_n2398_, men_men_n2399_, men_men_n2400_, men_men_n2401_, men_men_n2402_, men_men_n2403_, men_men_n2404_, men_men_n2405_, men_men_n2406_, men_men_n2407_, men_men_n2408_, men_men_n2409_, men_men_n2410_, men_men_n2411_, men_men_n2412_, men_men_n2413_, men_men_n2414_, men_men_n2415_, men_men_n2416_, men_men_n2417_, men_men_n2418_, men_men_n2419_, men_men_n2420_, men_men_n2422_, men_men_n2423_, men_men_n2424_, men_men_n2425_, men_men_n2426_, men_men_n2427_, men_men_n2428_, men_men_n2429_, men_men_n2430_, men_men_n2431_, men_men_n2432_, men_men_n2433_, men_men_n2434_, men_men_n2435_, men_men_n2436_, men_men_n2437_, men_men_n2438_, men_men_n2439_, men_men_n2440_, men_men_n2441_, men_men_n2442_, men_men_n2443_, men_men_n2444_, men_men_n2445_, men_men_n2446_, men_men_n2447_, men_men_n2448_, men_men_n2449_, men_men_n2450_, men_men_n2451_, men_men_n2452_, men_men_n2453_, men_men_n2454_, men_men_n2455_, men_men_n2456_, men_men_n2457_, men_men_n2458_, men_men_n2459_, men_men_n2460_, men_men_n2461_, men_men_n2462_, men_men_n2463_, men_men_n2464_, men_men_n2465_, men_men_n2466_, men_men_n2467_, men_men_n2468_, men_men_n2469_, men_men_n2470_, men_men_n2471_, men_men_n2472_, men_men_n2473_, men_men_n2474_, men_men_n2475_, men_men_n2476_, men_men_n2477_, men_men_n2478_, men_men_n2479_, men_men_n2481_, men_men_n2482_, men_men_n2483_, men_men_n2484_, men_men_n2485_, men_men_n2486_, men_men_n2487_, men_men_n2488_, men_men_n2489_, men_men_n2490_, men_men_n2491_, men_men_n2492_, men_men_n2493_, men_men_n2494_, men_men_n2495_, men_men_n2496_, men_men_n2497_, men_men_n2498_, men_men_n2499_, men_men_n2500_, men_men_n2501_, men_men_n2502_, men_men_n2503_, men_men_n2504_, men_men_n2505_, men_men_n2506_, men_men_n2507_, men_men_n2508_, men_men_n2509_, men_men_n2510_, men_men_n2511_, men_men_n2512_, men_men_n2513_, men_men_n2514_, men_men_n2515_, men_men_n2516_, men_men_n2517_, men_men_n2518_, men_men_n2519_, men_men_n2520_, men_men_n2521_, men_men_n2522_, men_men_n2523_, men_men_n2524_, men_men_n2525_, men_men_n2526_, men_men_n2527_, men_men_n2528_, men_men_n2529_, men_men_n2530_, men_men_n2531_, men_men_n2532_, men_men_n2533_, men_men_n2534_, men_men_n2535_, men_men_n2536_, men_men_n2537_, men_men_n2538_, men_men_n2539_, men_men_n2540_, men_men_n2541_, men_men_n2542_, men_men_n2543_, men_men_n2544_, men_men_n2545_, men_men_n2546_, men_men_n2550_, men_men_n2551_, men_men_n2552_, men_men_n2553_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13, ori14, mai14, men14, ori15, mai15, men15, ori16, mai16, men16, ori17, mai17, men17, ori18, mai18, men18, ori19, mai19, men19, ori20, mai20, men20, ori21, mai21, men21, ori22, mai22, men22, ori23, mai23, men23, ori24, mai24, men24, ori25, mai25, men25, ori26, mai26, men26, ori27, mai27, men27, ori28, mai28, men28, ori29, mai29, men29, ori30, mai30, men30, ori31, mai31, men31, ori32, mai32, men32, ori33, mai33, men33, ori34, mai34, men34, ori35, mai35, men35, ori36, mai36, men36, ori37, mai37, men37, ori38, mai38, men38, ori39, mai39, men39;
  INV        o0000(.A(x3), .Y(ori_ori_n50_));
  NA2        o0001(.A(ori_ori_n50_), .B(x2), .Y(ori_ori_n51_));
  NA2        o0002(.A(x7), .B(x0), .Y(ori_ori_n52_));
  INV        o0003(.A(x1), .Y(ori_ori_n53_));
  NA2        o0004(.A(x5), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  INV        o0005(.A(x8), .Y(ori_ori_n55_));
  INV        o0006(.A(x4), .Y(ori_ori_n56_));
  INV        o0007(.A(x7), .Y(ori_ori_n57_));
  NA2        o0008(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0009(.A(x0), .Y(ori_ori_n59_));
  NA2        o0010(.A(x4), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NA4        o0011(.A(ori_ori_n60_), .B(ori_ori_n58_), .C(ori_ori_n55_), .D(x6), .Y(ori_ori_n61_));
  NA2        o0012(.A(ori_ori_n56_), .B(ori_ori_n59_), .Y(ori_ori_n62_));
  NO2        o0013(.A(ori_ori_n55_), .B(x6), .Y(ori_ori_n63_));
  NA2        o0014(.A(ori_ori_n57_), .B(x4), .Y(ori_ori_n64_));
  NA3        o0015(.A(ori_ori_n64_), .B(ori_ori_n63_), .C(ori_ori_n62_), .Y(ori_ori_n65_));
  AOI210     o0016(.A0(ori_ori_n65_), .A1(ori_ori_n61_), .B0(ori_ori_n54_), .Y(ori_ori_n66_));
  NO2        o0017(.A(x8), .B(ori_ori_n57_), .Y(ori_ori_n67_));
  NO2        o0018(.A(x7), .B(ori_ori_n59_), .Y(ori_ori_n68_));
  NO2        o0019(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  NAi21      o0020(.An(x5), .B(x1), .Y(ori_ori_n70_));
  INV        o0021(.A(x6), .Y(ori_ori_n71_));
  NA2        o0022(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n72_));
  NO3        o0023(.A(ori_ori_n72_), .B(ori_ori_n70_), .C(ori_ori_n69_), .Y(ori_ori_n73_));
  OAI210     o0024(.A0(ori_ori_n73_), .A1(ori_ori_n66_), .B0(ori_ori_n52_), .Y(ori_ori_n74_));
  NA2        o0025(.A(x7), .B(x4), .Y(ori_ori_n75_));
  NO2        o0026(.A(ori_ori_n75_), .B(x1), .Y(ori_ori_n76_));
  NO2        o0027(.A(ori_ori_n71_), .B(x5), .Y(ori_ori_n77_));
  NO2        o0028(.A(x8), .B(ori_ori_n59_), .Y(ori_ori_n78_));
  NA3        o0029(.A(ori_ori_n78_), .B(ori_ori_n77_), .C(ori_ori_n76_), .Y(ori_ori_n79_));
  AOI210     o0030(.A0(ori_ori_n79_), .A1(ori_ori_n74_), .B0(ori_ori_n51_), .Y(ori_ori_n80_));
  NA2        o0031(.A(x5), .B(x3), .Y(ori_ori_n81_));
  NO2        o0032(.A(x6), .B(x0), .Y(ori_ori_n82_));
  NO2        o0033(.A(ori_ori_n82_), .B(x4), .Y(ori_ori_n83_));
  NO2        o0034(.A(x4), .B(x2), .Y(ori_ori_n84_));
  NO2        o0035(.A(ori_ori_n71_), .B(ori_ori_n59_), .Y(ori_ori_n85_));
  NO2        o0036(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n86_));
  NA2        o0037(.A(x8), .B(x1), .Y(ori_ori_n87_));
  NO2        o0038(.A(ori_ori_n87_), .B(x7), .Y(ori_ori_n88_));
  NO3        o0039(.A(x8), .B(ori_ori_n57_), .C(x6), .Y(ori_ori_n89_));
  NO2        o0040(.A(x1), .B(ori_ori_n59_), .Y(ori_ori_n90_));
  NO2        o0041(.A(ori_ori_n56_), .B(x2), .Y(ori_ori_n91_));
  XO2        o0042(.A(x7), .B(x1), .Y(ori_ori_n92_));
  INV        o0043(.A(ori_ori_n92_), .Y(ori_ori_n93_));
  NO2        o0044(.A(ori_ori_n93_), .B(x6), .Y(ori_ori_n94_));
  NO2        o0045(.A(ori_ori_n50_), .B(x0), .Y(ori_ori_n95_));
  NA2        o0046(.A(ori_ori_n95_), .B(ori_ori_n55_), .Y(ori_ori_n96_));
  NO2        o0047(.A(x6), .B(x5), .Y(ori_ori_n97_));
  NO2        o0048(.A(ori_ori_n57_), .B(x5), .Y(ori_ori_n98_));
  NO2        o0049(.A(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  NA2        o0050(.A(x6), .B(x1), .Y(ori_ori_n100_));
  NA2        o0051(.A(ori_ori_n100_), .B(ori_ori_n84_), .Y(ori_ori_n101_));
  NO4        o0052(.A(ori_ori_n101_), .B(ori_ori_n99_), .C(ori_ori_n96_), .D(ori_ori_n94_), .Y(ori_ori_n102_));
  NA2        o0053(.A(x3), .B(x0), .Y(ori_ori_n103_));
  INV        o0054(.A(x5), .Y(ori_ori_n104_));
  NA2        o0055(.A(ori_ori_n71_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  INV        o0056(.A(x2), .Y(ori_ori_n106_));
  NO2        o0057(.A(ori_ori_n56_), .B(ori_ori_n106_), .Y(ori_ori_n107_));
  NA2        o0058(.A(ori_ori_n57_), .B(ori_ori_n104_), .Y(ori_ori_n108_));
  NA3        o0059(.A(ori_ori_n108_), .B(ori_ori_n107_), .C(ori_ori_n105_), .Y(ori_ori_n109_));
  NO3        o0060(.A(ori_ori_n109_), .B(ori_ori_n103_), .C(ori_ori_n53_), .Y(ori_ori_n110_));
  NO3        o0061(.A(ori_ori_n110_), .B(ori_ori_n102_), .C(ori_ori_n80_), .Y(ori00));
  NO2        o0062(.A(x7), .B(x6), .Y(ori_ori_n112_));
  INV        o0063(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  NO2        o0064(.A(ori_ori_n55_), .B(ori_ori_n53_), .Y(ori_ori_n114_));
  NA2        o0065(.A(ori_ori_n114_), .B(ori_ori_n56_), .Y(ori_ori_n115_));
  XN2        o0066(.A(x6), .B(x1), .Y(ori_ori_n116_));
  INV        o0067(.A(ori_ori_n116_), .Y(ori_ori_n117_));
  NO2        o0068(.A(x6), .B(x4), .Y(ori_ori_n118_));
  NA2        o0069(.A(x6), .B(x4), .Y(ori_ori_n119_));
  NAi21      o0070(.An(ori_ori_n118_), .B(ori_ori_n119_), .Y(ori_ori_n120_));
  XN2        o0071(.A(x7), .B(x6), .Y(ori_ori_n121_));
  NO2        o0072(.A(x3), .B(ori_ori_n106_), .Y(ori_ori_n122_));
  NA2        o0073(.A(ori_ori_n122_), .B(ori_ori_n104_), .Y(ori_ori_n123_));
  NA2        o0074(.A(x3), .B(ori_ori_n106_), .Y(ori_ori_n124_));
  NO2        o0075(.A(ori_ori_n55_), .B(ori_ori_n57_), .Y(ori_ori_n125_));
  NA2        o0076(.A(ori_ori_n125_), .B(ori_ori_n56_), .Y(ori_ori_n126_));
  NA2        o0077(.A(ori_ori_n55_), .B(ori_ori_n57_), .Y(ori_ori_n127_));
  NA2        o0078(.A(ori_ori_n127_), .B(x2), .Y(ori_ori_n128_));
  NA2        o0079(.A(x8), .B(x3), .Y(ori_ori_n129_));
  NO2        o0080(.A(x5), .B(x0), .Y(ori_ori_n130_));
  NO2        o0081(.A(x6), .B(x1), .Y(ori_ori_n131_));
  NA2        o0082(.A(x8), .B(ori_ori_n104_), .Y(ori_ori_n132_));
  NA2        o0083(.A(x4), .B(ori_ori_n50_), .Y(ori_ori_n133_));
  NAi21      o0084(.An(x7), .B(x2), .Y(ori_ori_n134_));
  XO2        o0085(.A(x8), .B(x7), .Y(ori_ori_n135_));
  NA2        o0086(.A(ori_ori_n135_), .B(ori_ori_n106_), .Y(ori_ori_n136_));
  NA2        o0087(.A(x6), .B(x5), .Y(ori_ori_n137_));
  NO2        o0088(.A(ori_ori_n56_), .B(x0), .Y(ori_ori_n138_));
  NO2        o0089(.A(ori_ori_n50_), .B(x1), .Y(ori_ori_n139_));
  NA2        o0090(.A(ori_ori_n139_), .B(ori_ori_n138_), .Y(ori_ori_n140_));
  NO3        o0091(.A(ori_ori_n140_), .B(ori_ori_n137_), .C(ori_ori_n136_), .Y(ori01));
  NA2        o0092(.A(ori_ori_n57_), .B(ori_ori_n59_), .Y(ori_ori_n142_));
  NO2        o0093(.A(x2), .B(x1), .Y(ori_ori_n143_));
  NA2        o0094(.A(x2), .B(x1), .Y(ori_ori_n144_));
  NOi21      o0095(.An(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n145_));
  NA2        o0096(.A(ori_ori_n104_), .B(ori_ori_n53_), .Y(ori_ori_n146_));
  INV        o0097(.A(ori_ori_n146_), .Y(ori_ori_n147_));
  NAi21      o0098(.An(x8), .B(x1), .Y(ori_ori_n148_));
  NO2        o0099(.A(ori_ori_n148_), .B(x3), .Y(ori_ori_n149_));
  OAI210     o0100(.A0(ori_ori_n149_), .A1(ori_ori_n147_), .B0(ori_ori_n145_), .Y(ori_ori_n150_));
  NO2        o0101(.A(x5), .B(ori_ori_n50_), .Y(ori_ori_n151_));
  NO2        o0102(.A(ori_ori_n106_), .B(x1), .Y(ori_ori_n152_));
  NO2        o0103(.A(ori_ori_n150_), .B(ori_ori_n142_), .Y(ori_ori_n153_));
  NAi21      o0104(.An(x7), .B(x0), .Y(ori_ori_n154_));
  NO2        o0105(.A(ori_ori_n55_), .B(x2), .Y(ori_ori_n155_));
  NO2        o0106(.A(ori_ori_n81_), .B(x1), .Y(ori_ori_n156_));
  NA2        o0107(.A(x5), .B(ori_ori_n50_), .Y(ori_ori_n157_));
  NO2        o0108(.A(ori_ori_n157_), .B(ori_ori_n148_), .Y(ori_ori_n158_));
  NA2        o0109(.A(x8), .B(x5), .Y(ori_ori_n159_));
  NO3        o0110(.A(x3), .B(ori_ori_n106_), .C(ori_ori_n53_), .Y(ori_ori_n160_));
  NO2        o0111(.A(ori_ori_n160_), .B(ori_ori_n158_), .Y(ori_ori_n161_));
  NO2        o0112(.A(ori_ori_n161_), .B(ori_ori_n154_), .Y(ori_ori_n162_));
  NO2        o0113(.A(ori_ori_n57_), .B(x3), .Y(ori_ori_n163_));
  NO2        o0114(.A(ori_ori_n55_), .B(x0), .Y(ori_ori_n164_));
  NA3        o0115(.A(ori_ori_n104_), .B(ori_ori_n106_), .C(x1), .Y(ori_ori_n165_));
  NO2        o0116(.A(ori_ori_n165_), .B(ori_ori_n164_), .Y(ori_ori_n166_));
  NO2        o0117(.A(ori_ori_n87_), .B(ori_ori_n50_), .Y(ori_ori_n167_));
  NA2        o0118(.A(ori_ori_n104_), .B(x0), .Y(ori_ori_n168_));
  NA2        o0119(.A(ori_ori_n166_), .B(ori_ori_n163_), .Y(ori_ori_n169_));
  NA2        o0120(.A(x7), .B(ori_ori_n106_), .Y(ori_ori_n170_));
  NA2        o0121(.A(ori_ori_n151_), .B(x8), .Y(ori_ori_n171_));
  NA4        o0122(.A(x5), .B(x3), .C(x1), .D(x0), .Y(ori_ori_n172_));
  AO210      o0123(.A0(ori_ori_n172_), .A1(ori_ori_n171_), .B0(ori_ori_n170_), .Y(ori_ori_n173_));
  NO2        o0124(.A(ori_ori_n144_), .B(ori_ori_n50_), .Y(ori_ori_n174_));
  NAi21      o0125(.An(x1), .B(x2), .Y(ori_ori_n175_));
  NO2        o0126(.A(ori_ori_n157_), .B(ori_ori_n175_), .Y(ori_ori_n176_));
  NA2        o0127(.A(x8), .B(x7), .Y(ori_ori_n177_));
  NO2        o0128(.A(ori_ori_n177_), .B(x0), .Y(ori_ori_n178_));
  NA2        o0129(.A(ori_ori_n174_), .B(ori_ori_n178_), .Y(ori_ori_n179_));
  NA3        o0130(.A(ori_ori_n179_), .B(ori_ori_n173_), .C(ori_ori_n169_), .Y(ori_ori_n180_));
  NO3        o0131(.A(ori_ori_n180_), .B(ori_ori_n162_), .C(ori_ori_n153_), .Y(ori_ori_n181_));
  NA2        o0132(.A(x3), .B(x1), .Y(ori_ori_n182_));
  NA2        o0133(.A(ori_ori_n50_), .B(ori_ori_n106_), .Y(ori_ori_n183_));
  NA2        o0134(.A(ori_ori_n176_), .B(ori_ori_n67_), .Y(ori_ori_n184_));
  NA2        o0135(.A(ori_ori_n125_), .B(ori_ori_n106_), .Y(ori_ori_n185_));
  OAI210     o0136(.A0(ori_ori_n185_), .A1(ori_ori_n182_), .B0(ori_ori_n184_), .Y(ori_ori_n186_));
  XO2        o0137(.A(x5), .B(x3), .Y(ori_ori_n187_));
  NA2        o0138(.A(ori_ori_n187_), .B(x8), .Y(ori_ori_n188_));
  NA2        o0139(.A(x8), .B(ori_ori_n59_), .Y(ori_ori_n189_));
  NA2        o0140(.A(x7), .B(ori_ori_n71_), .Y(ori_ori_n190_));
  NO2        o0141(.A(ori_ori_n175_), .B(ori_ori_n190_), .Y(ori_ori_n191_));
  NA2        o0142(.A(ori_ori_n186_), .B(x0), .Y(ori_ori_n192_));
  OAI210     o0143(.A0(ori_ori_n181_), .A1(ori_ori_n71_), .B0(ori_ori_n192_), .Y(ori_ori_n193_));
  NO2        o0144(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n194_));
  NA4        o0145(.A(ori_ori_n55_), .B(x5), .C(x3), .D(x2), .Y(ori_ori_n195_));
  NA2        o0146(.A(x8), .B(ori_ori_n50_), .Y(ori_ori_n196_));
  INV        o0147(.A(x2), .Y(ori_ori_n197_));
  NA2        o0148(.A(ori_ori_n55_), .B(x3), .Y(ori_ori_n198_));
  NO2        o0149(.A(ori_ori_n195_), .B(ori_ori_n53_), .Y(ori_ori_n199_));
  NO2        o0150(.A(ori_ori_n106_), .B(ori_ori_n59_), .Y(ori_ori_n200_));
  NA2        o0151(.A(x5), .B(x1), .Y(ori_ori_n201_));
  NO2        o0152(.A(ori_ori_n201_), .B(x6), .Y(ori_ori_n202_));
  NO2        o0153(.A(x3), .B(x1), .Y(ori_ori_n203_));
  AOI210     o0154(.A0(ori_ori_n203_), .A1(ori_ori_n77_), .B0(ori_ori_n202_), .Y(ori_ori_n204_));
  NO2        o0155(.A(ori_ori_n81_), .B(ori_ori_n55_), .Y(ori_ori_n205_));
  NO2        o0156(.A(ori_ori_n100_), .B(ori_ori_n50_), .Y(ori_ori_n206_));
  NO2        o0157(.A(ori_ori_n206_), .B(ori_ori_n205_), .Y(ori_ori_n207_));
  OAI210     o0158(.A0(ori_ori_n204_), .A1(x8), .B0(ori_ori_n207_), .Y(ori_ori_n208_));
  NO2        o0159(.A(ori_ori_n55_), .B(x5), .Y(ori_ori_n209_));
  NA2        o0160(.A(ori_ori_n209_), .B(ori_ori_n71_), .Y(ori_ori_n210_));
  NAi21      o0161(.An(x2), .B(x5), .Y(ori_ori_n211_));
  NA2        o0162(.A(x8), .B(x6), .Y(ori_ori_n212_));
  NA2        o0163(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n213_));
  AN2        o0164(.A(ori_ori_n208_), .B(ori_ori_n200_), .Y(ori_ori_n214_));
  OAI210     o0165(.A0(ori_ori_n214_), .A1(ori_ori_n199_), .B0(ori_ori_n194_), .Y(ori_ori_n215_));
  NA2        o0166(.A(ori_ori_n71_), .B(ori_ori_n56_), .Y(ori_ori_n216_));
  NO2        o0167(.A(ori_ori_n216_), .B(x7), .Y(ori_ori_n217_));
  NO2        o0168(.A(ori_ori_n104_), .B(ori_ori_n53_), .Y(ori_ori_n218_));
  NA2        o0169(.A(ori_ori_n218_), .B(ori_ori_n106_), .Y(ori_ori_n219_));
  NA2        o0170(.A(x3), .B(ori_ori_n59_), .Y(ori_ori_n220_));
  NO2        o0171(.A(ori_ori_n165_), .B(ori_ori_n220_), .Y(ori_ori_n221_));
  NO2        o0172(.A(x1), .B(x0), .Y(ori_ori_n222_));
  NA2        o0173(.A(ori_ori_n222_), .B(ori_ori_n106_), .Y(ori_ori_n223_));
  NA2        o0174(.A(ori_ori_n104_), .B(ori_ori_n50_), .Y(ori_ori_n224_));
  XN2        o0175(.A(x3), .B(x2), .Y(ori_ori_n225_));
  NO2        o0176(.A(ori_ori_n104_), .B(x0), .Y(ori_ori_n226_));
  NA2        o0177(.A(x8), .B(ori_ori_n53_), .Y(ori_ori_n227_));
  NO2        o0178(.A(ori_ori_n224_), .B(ori_ori_n223_), .Y(ori_ori_n228_));
  NA2        o0179(.A(ori_ori_n228_), .B(ori_ori_n217_), .Y(ori_ori_n229_));
  NO2        o0180(.A(x7), .B(x1), .Y(ori_ori_n230_));
  NOi21      o0181(.An(x8), .B(x3), .Y(ori_ori_n231_));
  NA2        o0182(.A(ori_ori_n231_), .B(ori_ori_n59_), .Y(ori_ori_n232_));
  NA2        o0183(.A(x5), .B(x0), .Y(ori_ori_n233_));
  NAi21      o0184(.An(ori_ori_n130_), .B(ori_ori_n233_), .Y(ori_ori_n234_));
  NA2        o0185(.A(ori_ori_n71_), .B(ori_ori_n50_), .Y(ori_ori_n235_));
  OAI210     o0186(.A0(ori_ori_n235_), .A1(ori_ori_n234_), .B0(ori_ori_n232_), .Y(ori_ori_n236_));
  NA3        o0187(.A(ori_ori_n236_), .B(ori_ori_n132_), .C(ori_ori_n230_), .Y(ori_ori_n237_));
  NA2        o0188(.A(x8), .B(ori_ori_n57_), .Y(ori_ori_n238_));
  NO2        o0189(.A(ori_ori_n238_), .B(x5), .Y(ori_ori_n239_));
  NO2        o0190(.A(ori_ori_n139_), .B(ori_ori_n71_), .Y(ori_ori_n240_));
  NA2        o0191(.A(x1), .B(x0), .Y(ori_ori_n241_));
  NA2        o0192(.A(ori_ori_n50_), .B(ori_ori_n59_), .Y(ori_ori_n242_));
  NA2        o0193(.A(ori_ori_n237_), .B(ori_ori_n172_), .Y(ori_ori_n243_));
  NO2        o0194(.A(ori_ori_n104_), .B(x3), .Y(ori_ori_n244_));
  NO2        o0195(.A(ori_ori_n106_), .B(x0), .Y(ori_ori_n245_));
  NO2        o0196(.A(ori_ori_n55_), .B(x7), .Y(ori_ori_n246_));
  NO3        o0197(.A(x8), .B(ori_ori_n50_), .C(x0), .Y(ori_ori_n247_));
  NAi21      o0198(.An(x8), .B(x0), .Y(ori_ori_n248_));
  NAi21      o0199(.An(x1), .B(x3), .Y(ori_ori_n249_));
  NO2        o0200(.A(ori_ori_n249_), .B(ori_ori_n248_), .Y(ori_ori_n250_));
  NO2        o0201(.A(x2), .B(ori_ori_n53_), .Y(ori_ori_n251_));
  AOI210     o0202(.A0(ori_ori_n251_), .A1(ori_ori_n247_), .B0(ori_ori_n250_), .Y(ori_ori_n252_));
  NOi21      o0203(.An(x5), .B(x6), .Y(ori_ori_n253_));
  NO2        o0204(.A(ori_ori_n57_), .B(x4), .Y(ori_ori_n254_));
  NA2        o0205(.A(ori_ori_n254_), .B(ori_ori_n253_), .Y(ori_ori_n255_));
  NO2        o0206(.A(ori_ori_n255_), .B(ori_ori_n252_), .Y(ori_ori_n256_));
  AOI210     o0207(.A0(ori_ori_n243_), .A1(ori_ori_n107_), .B0(ori_ori_n256_), .Y(ori_ori_n257_));
  NA3        o0208(.A(ori_ori_n257_), .B(ori_ori_n229_), .C(ori_ori_n215_), .Y(ori_ori_n258_));
  AOI210     o0209(.A0(ori_ori_n193_), .A1(ori_ori_n56_), .B0(ori_ori_n258_), .Y(ori02));
  NO2        o0210(.A(x8), .B(ori_ori_n104_), .Y(ori_ori_n260_));
  XN2        o0211(.A(x7), .B(x3), .Y(ori_ori_n261_));
  INV        o0212(.A(ori_ori_n261_), .Y(ori_ori_n262_));
  NO2        o0213(.A(x2), .B(x0), .Y(ori_ori_n263_));
  NA2        o0214(.A(ori_ori_n263_), .B(ori_ori_n71_), .Y(ori_ori_n264_));
  NO2        o0215(.A(ori_ori_n57_), .B(x1), .Y(ori_ori_n265_));
  NO3        o0216(.A(ori_ori_n265_), .B(ori_ori_n264_), .C(ori_ori_n262_), .Y(ori_ori_n266_));
  NA2        o0217(.A(ori_ori_n53_), .B(x0), .Y(ori_ori_n267_));
  NO2        o0218(.A(ori_ori_n249_), .B(x6), .Y(ori_ori_n268_));
  XO2        o0219(.A(x7), .B(x0), .Y(ori_ori_n269_));
  NO2        o0220(.A(ori_ori_n269_), .B(ori_ori_n263_), .Y(ori_ori_n270_));
  NA2        o0221(.A(ori_ori_n270_), .B(ori_ori_n268_), .Y(ori_ori_n271_));
  AN2        o0222(.A(x7), .B(x2), .Y(ori_ori_n272_));
  NA2        o0223(.A(ori_ori_n272_), .B(ori_ori_n50_), .Y(ori_ori_n273_));
  OAI210     o0224(.A0(ori_ori_n273_), .A1(ori_ori_n267_), .B0(ori_ori_n271_), .Y(ori_ori_n274_));
  OAI210     o0225(.A0(ori_ori_n274_), .A1(ori_ori_n266_), .B0(ori_ori_n260_), .Y(ori_ori_n275_));
  NAi21      o0226(.An(x8), .B(x6), .Y(ori_ori_n276_));
  NO2        o0227(.A(ori_ori_n104_), .B(ori_ori_n59_), .Y(ori_ori_n277_));
  NA2        o0228(.A(x7), .B(x3), .Y(ori_ori_n278_));
  NO2        o0229(.A(ori_ori_n278_), .B(x2), .Y(ori_ori_n279_));
  NA2        o0230(.A(x2), .B(x0), .Y(ori_ori_n280_));
  NA2        o0231(.A(ori_ori_n106_), .B(ori_ori_n59_), .Y(ori_ori_n281_));
  NA2        o0232(.A(ori_ori_n281_), .B(ori_ori_n280_), .Y(ori_ori_n282_));
  NAi21      o0233(.An(x7), .B(x1), .Y(ori_ori_n283_));
  NO2        o0234(.A(ori_ori_n283_), .B(x3), .Y(ori_ori_n284_));
  AOI220     o0235(.A0(ori_ori_n284_), .A1(ori_ori_n282_), .B0(ori_ori_n279_), .B1(ori_ori_n277_), .Y(ori_ori_n285_));
  NA2        o0236(.A(ori_ori_n251_), .B(ori_ori_n50_), .Y(ori_ori_n286_));
  NA3        o0237(.A(x7), .B(ori_ori_n104_), .C(x0), .Y(ori_ori_n287_));
  NA2        o0238(.A(ori_ori_n151_), .B(ori_ori_n57_), .Y(ori_ori_n288_));
  NO2        o0239(.A(ori_ori_n285_), .B(ori_ori_n276_), .Y(ori_ori_n289_));
  INV        o0240(.A(ori_ori_n269_), .Y(ori_ori_n290_));
  NO2        o0241(.A(x7), .B(ori_ori_n71_), .Y(ori_ori_n291_));
  NA2        o0242(.A(ori_ori_n104_), .B(x3), .Y(ori_ori_n292_));
  NO2        o0243(.A(ori_ori_n292_), .B(ori_ori_n291_), .Y(ori_ori_n293_));
  NA2        o0244(.A(ori_ori_n293_), .B(ori_ori_n290_), .Y(ori_ori_n294_));
  NA2        o0245(.A(ori_ori_n50_), .B(x0), .Y(ori_ori_n295_));
  NO2        o0246(.A(ori_ori_n295_), .B(x7), .Y(ori_ori_n296_));
  NA2        o0247(.A(ori_ori_n155_), .B(x1), .Y(ori_ori_n297_));
  NO2        o0248(.A(ori_ori_n294_), .B(ori_ori_n297_), .Y(ori_ori_n298_));
  NO2        o0249(.A(ori_ori_n57_), .B(ori_ori_n50_), .Y(ori_ori_n299_));
  NO2        o0250(.A(ori_ori_n55_), .B(ori_ori_n106_), .Y(ori_ori_n300_));
  NA3        o0251(.A(ori_ori_n300_), .B(ori_ori_n299_), .C(ori_ori_n59_), .Y(ori_ori_n301_));
  NO2        o0252(.A(ori_ori_n146_), .B(x6), .Y(ori_ori_n302_));
  NO2        o0253(.A(ori_ori_n100_), .B(ori_ori_n104_), .Y(ori_ori_n303_));
  NA2        o0254(.A(ori_ori_n57_), .B(ori_ori_n106_), .Y(ori_ori_n304_));
  NO2        o0255(.A(ori_ori_n304_), .B(ori_ori_n242_), .Y(ori_ori_n305_));
  OAI210     o0256(.A0(ori_ori_n303_), .A1(ori_ori_n302_), .B0(ori_ori_n305_), .Y(ori_ori_n306_));
  OAI210     o0257(.A0(ori_ori_n301_), .A1(ori_ori_n100_), .B0(ori_ori_n306_), .Y(ori_ori_n307_));
  NO3        o0258(.A(ori_ori_n307_), .B(ori_ori_n298_), .C(ori_ori_n289_), .Y(ori_ori_n308_));
  AOI210     o0259(.A0(ori_ori_n308_), .A1(ori_ori_n275_), .B0(x4), .Y(ori_ori_n309_));
  NA2        o0260(.A(x8), .B(ori_ori_n71_), .Y(ori_ori_n310_));
  NO2        o0261(.A(x3), .B(ori_ori_n59_), .Y(ori_ori_n311_));
  NO2        o0262(.A(x3), .B(x0), .Y(ori_ori_n312_));
  NAi21      o0263(.An(ori_ori_n312_), .B(ori_ori_n103_), .Y(ori_ori_n313_));
  NA2        o0264(.A(x5), .B(x2), .Y(ori_ori_n314_));
  INV        o0265(.A(ori_ori_n314_), .Y(ori_ori_n315_));
  NO2        o0266(.A(ori_ori_n106_), .B(ori_ori_n53_), .Y(ori_ori_n316_));
  NA2        o0267(.A(ori_ori_n316_), .B(x3), .Y(ori_ori_n317_));
  NO2        o0268(.A(ori_ori_n55_), .B(x1), .Y(ori_ori_n318_));
  NA2        o0269(.A(ori_ori_n318_), .B(ori_ori_n106_), .Y(ori_ori_n319_));
  INV        o0270(.A(ori_ori_n317_), .Y(ori_ori_n320_));
  NAi32      o0271(.An(x3), .Bn(x0), .C(x2), .Y(ori_ori_n321_));
  NO2        o0272(.A(ori_ori_n50_), .B(x2), .Y(ori_ori_n322_));
  NAi21      o0273(.An(x6), .B(x5), .Y(ori_ori_n323_));
  NO2        o0274(.A(x2), .B(ori_ori_n59_), .Y(ori_ori_n324_));
  NO4        o0275(.A(ori_ori_n324_), .B(ori_ori_n323_), .C(ori_ori_n148_), .D(ori_ori_n322_), .Y(ori_ori_n325_));
  AOI220     o0276(.A0(ori_ori_n325_), .A1(ori_ori_n321_), .B0(ori_ori_n320_), .B1(ori_ori_n85_), .Y(ori_ori_n326_));
  NO2        o0277(.A(ori_ori_n326_), .B(ori_ori_n75_), .Y(ori_ori_n327_));
  NO2        o0278(.A(ori_ori_n104_), .B(ori_ori_n50_), .Y(ori_ori_n328_));
  NO2        o0279(.A(ori_ori_n263_), .B(ori_ori_n200_), .Y(ori_ori_n329_));
  XO2        o0280(.A(x7), .B(x2), .Y(ori_ori_n330_));
  INV        o0281(.A(ori_ori_n330_), .Y(ori_ori_n331_));
  XO2        o0282(.A(x6), .B(x2), .Y(ori_ori_n332_));
  NAi21      o0283(.An(x0), .B(x6), .Y(ori_ori_n333_));
  XN2        o0284(.A(x7), .B(x5), .Y(ori_ori_n334_));
  NA2        o0285(.A(x7), .B(x5), .Y(ori_ori_n335_));
  NO2        o0286(.A(x8), .B(x6), .Y(ori_ori_n336_));
  NAi21      o0287(.An(ori_ori_n336_), .B(ori_ori_n212_), .Y(ori_ori_n337_));
  NA2        o0288(.A(ori_ori_n104_), .B(x2), .Y(ori_ori_n338_));
  NO2        o0289(.A(ori_ori_n338_), .B(ori_ori_n64_), .Y(ori_ori_n339_));
  NA2        o0290(.A(x1), .B(ori_ori_n59_), .Y(ori_ori_n340_));
  NA2        o0291(.A(x4), .B(x2), .Y(ori_ori_n341_));
  NO2        o0292(.A(ori_ori_n341_), .B(ori_ori_n104_), .Y(ori_ori_n342_));
  NAi21      o0293(.An(x1), .B(x6), .Y(ori_ori_n343_));
  NA2        o0294(.A(ori_ori_n312_), .B(ori_ori_n246_), .Y(ori_ori_n344_));
  OAI220     o0295(.A0(ori_ori_n344_), .A1(ori_ori_n343_), .B0(ori_ori_n103_), .B1(ori_ori_n53_), .Y(ori_ori_n345_));
  NA2        o0296(.A(x8), .B(x2), .Y(ori_ori_n346_));
  NO2        o0297(.A(ori_ori_n346_), .B(ori_ori_n50_), .Y(ori_ori_n347_));
  NA2        o0298(.A(ori_ori_n345_), .B(ori_ori_n342_), .Y(ori_ori_n348_));
  INV        o0299(.A(ori_ori_n348_), .Y(ori_ori_n349_));
  NO3        o0300(.A(ori_ori_n349_), .B(ori_ori_n327_), .C(ori_ori_n309_), .Y(ori03));
  NAi21      o0301(.An(x2), .B(x0), .Y(ori_ori_n351_));
  NO3        o0302(.A(x8), .B(x6), .C(x4), .Y(ori_ori_n352_));
  INV        o0303(.A(ori_ori_n352_), .Y(ori_ori_n353_));
  NA2        o0304(.A(ori_ori_n107_), .B(ori_ori_n59_), .Y(ori_ori_n354_));
  NO2        o0305(.A(ori_ori_n354_), .B(ori_ori_n55_), .Y(ori_ori_n355_));
  NA2        o0306(.A(ori_ori_n355_), .B(ori_ori_n151_), .Y(ori_ori_n356_));
  NA2        o0307(.A(x3), .B(x2), .Y(ori_ori_n357_));
  NO2        o0308(.A(ori_ori_n148_), .B(x0), .Y(ori_ori_n358_));
  NA2        o0309(.A(x8), .B(x0), .Y(ori_ori_n359_));
  NO2        o0310(.A(ori_ori_n359_), .B(x6), .Y(ori_ori_n360_));
  AOI210     o0311(.A0(ori_ori_n360_), .A1(x5), .B0(ori_ori_n358_), .Y(ori_ori_n361_));
  NO2        o0312(.A(ori_ori_n361_), .B(ori_ori_n357_), .Y(ori_ori_n362_));
  NO2        o0313(.A(x5), .B(ori_ori_n59_), .Y(ori_ori_n363_));
  NO2        o0314(.A(x3), .B(x2), .Y(ori_ori_n364_));
  NA2        o0315(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n365_));
  NO2        o0316(.A(ori_ori_n53_), .B(x0), .Y(ori_ori_n366_));
  NA2        o0317(.A(ori_ori_n366_), .B(x5), .Y(ori_ori_n367_));
  AOI210     o0318(.A0(ori_ori_n367_), .A1(ori_ori_n365_), .B0(ori_ori_n276_), .Y(ori_ori_n368_));
  NA2        o0319(.A(ori_ori_n232_), .B(ori_ori_n159_), .Y(ori_ori_n369_));
  NO2        o0320(.A(ori_ori_n50_), .B(ori_ori_n59_), .Y(ori_ori_n370_));
  NO2        o0321(.A(ori_ori_n71_), .B(x0), .Y(ori_ori_n371_));
  NO4        o0322(.A(ori_ori_n371_), .B(ori_ori_n370_), .C(x2), .D(ori_ori_n53_), .Y(ori_ori_n372_));
  AO210      o0323(.A0(ori_ori_n372_), .A1(ori_ori_n369_), .B0(ori_ori_n368_), .Y(ori_ori_n373_));
  OAI210     o0324(.A0(ori_ori_n373_), .A1(ori_ori_n362_), .B0(x4), .Y(ori_ori_n374_));
  NO2        o0325(.A(x4), .B(ori_ori_n53_), .Y(ori_ori_n375_));
  NA2        o0326(.A(ori_ori_n375_), .B(ori_ori_n59_), .Y(ori_ori_n376_));
  NO3        o0327(.A(ori_ori_n376_), .B(ori_ori_n212_), .C(x5), .Y(ori_ori_n377_));
  NA2        o0328(.A(x7), .B(ori_ori_n104_), .Y(ori_ori_n378_));
  NO3        o0329(.A(x5), .B(ori_ori_n53_), .C(x0), .Y(ori_ori_n379_));
  INV        o0330(.A(ori_ori_n379_), .Y(ori_ori_n380_));
  NO2        o0331(.A(x6), .B(ori_ori_n56_), .Y(ori_ori_n381_));
  NO2        o0332(.A(x8), .B(ori_ori_n50_), .Y(ori_ori_n382_));
  NA2        o0333(.A(ori_ori_n382_), .B(ori_ori_n381_), .Y(ori_ori_n383_));
  OAI210     o0334(.A0(ori_ori_n383_), .A1(ori_ori_n380_), .B0(ori_ori_n378_), .Y(ori_ori_n384_));
  AOI210     o0335(.A0(ori_ori_n377_), .A1(x2), .B0(ori_ori_n384_), .Y(ori_ori_n385_));
  AOI220     o0336(.A0(ori_ori_n385_), .A1(ori_ori_n374_), .B0(ori_ori_n356_), .B1(x7), .Y(ori_ori_n386_));
  NA2        o0337(.A(x7), .B(ori_ori_n53_), .Y(ori_ori_n387_));
  NO2        o0338(.A(ori_ori_n231_), .B(ori_ori_n106_), .Y(ori_ori_n388_));
  NO2        o0339(.A(ori_ori_n55_), .B(ori_ori_n59_), .Y(ori_ori_n389_));
  NO3        o0340(.A(ori_ori_n389_), .B(ori_ori_n388_), .C(ori_ori_n137_), .Y(ori_ori_n390_));
  AOI210     o0341(.A0(x8), .A1(ori_ori_n97_), .B0(ori_ori_n390_), .Y(ori_ori_n391_));
  NO2        o0342(.A(x5), .B(x2), .Y(ori_ori_n392_));
  NO2        o0343(.A(x8), .B(x3), .Y(ori_ori_n393_));
  NA2        o0344(.A(ori_ori_n393_), .B(ori_ori_n392_), .Y(ori_ori_n394_));
  NA2        o0345(.A(ori_ori_n189_), .B(x2), .Y(ori_ori_n395_));
  NO3        o0346(.A(ori_ori_n393_), .B(ori_ori_n313_), .C(ori_ori_n323_), .Y(ori_ori_n396_));
  NA2        o0347(.A(ori_ori_n396_), .B(ori_ori_n395_), .Y(ori_ori_n397_));
  OAI210     o0348(.A0(ori_ori_n391_), .A1(ori_ori_n263_), .B0(ori_ori_n397_), .Y(ori_ori_n398_));
  NA2        o0349(.A(ori_ori_n398_), .B(x4), .Y(ori_ori_n399_));
  NA2        o0350(.A(ori_ori_n55_), .B(ori_ori_n59_), .Y(ori_ori_n400_));
  NO2        o0351(.A(ori_ori_n400_), .B(x5), .Y(ori_ori_n401_));
  NAi21      o0352(.An(x4), .B(x6), .Y(ori_ori_n402_));
  NO2        o0353(.A(ori_ori_n402_), .B(ori_ori_n51_), .Y(ori_ori_n403_));
  NO2        o0354(.A(ori_ori_n55_), .B(ori_ori_n71_), .Y(ori_ori_n404_));
  NO2        o0355(.A(ori_ori_n50_), .B(ori_ori_n106_), .Y(ori_ori_n405_));
  NO2        o0356(.A(ori_ori_n212_), .B(x0), .Y(ori_ori_n406_));
  NO2        o0357(.A(ori_ori_n323_), .B(x8), .Y(ori_ori_n407_));
  OAI210     o0358(.A0(ori_ori_n407_), .A1(ori_ori_n406_), .B0(ori_ori_n405_), .Y(ori_ori_n408_));
  NA2        o0359(.A(ori_ori_n365_), .B(ori_ori_n408_), .Y(ori_ori_n409_));
  AOI220     o0360(.A0(ori_ori_n409_), .A1(ori_ori_n56_), .B0(ori_ori_n403_), .B1(ori_ori_n401_), .Y(ori_ori_n410_));
  AOI210     o0361(.A0(ori_ori_n410_), .A1(ori_ori_n399_), .B0(ori_ori_n387_), .Y(ori_ori_n411_));
  NA2        o0362(.A(ori_ori_n57_), .B(ori_ori_n53_), .Y(ori_ori_n412_));
  NO2        o0363(.A(ori_ori_n71_), .B(ori_ori_n56_), .Y(ori_ori_n413_));
  NA2        o0364(.A(ori_ori_n322_), .B(ori_ori_n59_), .Y(ori_ori_n414_));
  NO3        o0365(.A(x6), .B(x4), .C(ori_ori_n50_), .Y(ori_ori_n415_));
  NA2        o0366(.A(ori_ori_n389_), .B(x5), .Y(ori_ori_n416_));
  NO2        o0367(.A(x8), .B(x5), .Y(ori_ori_n417_));
  NAi21      o0368(.An(ori_ori_n417_), .B(ori_ori_n159_), .Y(ori_ori_n418_));
  OAI210     o0369(.A0(ori_ori_n418_), .A1(ori_ori_n281_), .B0(ori_ori_n416_), .Y(ori_ori_n419_));
  NA2        o0370(.A(ori_ori_n329_), .B(ori_ori_n77_), .Y(ori_ori_n420_));
  NOi21      o0371(.An(x3), .B(x4), .Y(ori_ori_n421_));
  NA2        o0372(.A(ori_ori_n55_), .B(ori_ori_n106_), .Y(ori_ori_n422_));
  NA2        o0373(.A(ori_ori_n422_), .B(ori_ori_n421_), .Y(ori_ori_n423_));
  NO2        o0374(.A(ori_ori_n51_), .B(x6), .Y(ori_ori_n424_));
  NO2        o0375(.A(ori_ori_n137_), .B(ori_ori_n55_), .Y(ori_ori_n425_));
  NO3        o0376(.A(ori_ori_n56_), .B(x2), .C(x0), .Y(ori_ori_n426_));
  AOI220     o0377(.A0(ori_ori_n426_), .A1(ori_ori_n425_), .B0(ori_ori_n424_), .B1(ori_ori_n401_), .Y(ori_ori_n427_));
  OAI210     o0378(.A0(ori_ori_n423_), .A1(ori_ori_n420_), .B0(ori_ori_n427_), .Y(ori_ori_n428_));
  AOI210     o0379(.A0(ori_ori_n419_), .A1(ori_ori_n415_), .B0(ori_ori_n428_), .Y(ori_ori_n429_));
  NO2        o0380(.A(ori_ori_n429_), .B(ori_ori_n412_), .Y(ori_ori_n430_));
  NA2        o0381(.A(x7), .B(x1), .Y(ori_ori_n431_));
  NO3        o0382(.A(x5), .B(x4), .C(x2), .Y(ori_ori_n432_));
  NO2        o0383(.A(x4), .B(ori_ori_n106_), .Y(ori_ori_n433_));
  NA2        o0384(.A(ori_ori_n433_), .B(x6), .Y(ori_ori_n434_));
  NA3        o0385(.A(ori_ori_n104_), .B(x4), .C(ori_ori_n106_), .Y(ori_ori_n435_));
  AOI210     o0386(.A0(ori_ori_n435_), .A1(ori_ori_n434_), .B0(ori_ori_n96_), .Y(ori_ori_n436_));
  NA2        o0387(.A(ori_ori_n421_), .B(ori_ori_n71_), .Y(ori_ori_n437_));
  NA2        o0388(.A(ori_ori_n155_), .B(ori_ori_n59_), .Y(ori_ori_n438_));
  NO2        o0389(.A(ori_ori_n438_), .B(ori_ori_n437_), .Y(ori_ori_n439_));
  NA2        o0390(.A(ori_ori_n405_), .B(x4), .Y(ori_ori_n440_));
  NO3        o0391(.A(ori_ori_n440_), .B(ori_ori_n336_), .C(ori_ori_n371_), .Y(ori_ori_n441_));
  NO3        o0392(.A(ori_ori_n441_), .B(ori_ori_n439_), .C(ori_ori_n436_), .Y(ori_ori_n442_));
  NA2        o0393(.A(x5), .B(x4), .Y(ori_ori_n443_));
  NO2        o0394(.A(ori_ori_n71_), .B(ori_ori_n53_), .Y(ori_ori_n444_));
  NO3        o0395(.A(x8), .B(x3), .C(x2), .Y(ori_ori_n445_));
  NA3        o0396(.A(ori_ori_n445_), .B(ori_ori_n444_), .C(ori_ori_n59_), .Y(ori_ori_n446_));
  NO3        o0397(.A(x6), .B(x5), .C(x2), .Y(ori_ori_n447_));
  NA3        o0398(.A(ori_ori_n447_), .B(ori_ori_n265_), .C(ori_ori_n78_), .Y(ori_ori_n448_));
  OAI210     o0399(.A0(ori_ori_n446_), .A1(ori_ori_n443_), .B0(ori_ori_n448_), .Y(ori_ori_n449_));
  NA2        o0400(.A(ori_ori_n71_), .B(x2), .Y(ori_ori_n450_));
  NO3        o0401(.A(x4), .B(x3), .C(ori_ori_n59_), .Y(ori_ori_n451_));
  NA2        o0402(.A(ori_ori_n451_), .B(ori_ori_n209_), .Y(ori_ori_n452_));
  NO3        o0403(.A(ori_ori_n452_), .B(ori_ori_n450_), .C(ori_ori_n92_), .Y(ori_ori_n453_));
  XO2        o0404(.A(x4), .B(x0), .Y(ori_ori_n454_));
  NA2        o0405(.A(ori_ori_n242_), .B(x5), .Y(ori_ori_n455_));
  NO2        o0406(.A(ori_ori_n56_), .B(ori_ori_n50_), .Y(ori_ori_n456_));
  NO2        o0407(.A(ori_ori_n456_), .B(ori_ori_n63_), .Y(ori_ori_n457_));
  NO4        o0408(.A(ori_ori_n457_), .B(ori_ori_n455_), .C(ori_ori_n454_), .D(ori_ori_n144_), .Y(ori_ori_n458_));
  NO3        o0409(.A(ori_ori_n458_), .B(ori_ori_n453_), .C(ori_ori_n449_), .Y(ori_ori_n459_));
  OAI210     o0410(.A0(ori_ori_n442_), .A1(ori_ori_n431_), .B0(ori_ori_n459_), .Y(ori_ori_n460_));
  NO4        o0411(.A(ori_ori_n460_), .B(ori_ori_n430_), .C(ori_ori_n411_), .D(ori_ori_n386_), .Y(ori04));
  NO2        o0412(.A(x7), .B(x2), .Y(ori_ori_n462_));
  NO2        o0413(.A(x3), .B(ori_ori_n53_), .Y(ori_ori_n463_));
  NO2        o0414(.A(ori_ori_n463_), .B(ori_ori_n139_), .Y(ori_ori_n464_));
  XN2        o0415(.A(x8), .B(x1), .Y(ori_ori_n465_));
  NO2        o0416(.A(ori_ori_n465_), .B(ori_ori_n137_), .Y(ori_ori_n466_));
  NA2        o0417(.A(ori_ori_n466_), .B(ori_ori_n464_), .Y(ori_ori_n467_));
  NA2        o0418(.A(x6), .B(x3), .Y(ori_ori_n468_));
  NO2        o0419(.A(ori_ori_n468_), .B(x5), .Y(ori_ori_n469_));
  NA2        o0420(.A(ori_ori_n71_), .B(x1), .Y(ori_ori_n470_));
  NO2        o0421(.A(ori_ori_n417_), .B(ori_ori_n231_), .Y(ori_ori_n471_));
  NO3        o0422(.A(ori_ori_n471_), .B(ori_ori_n393_), .C(ori_ori_n470_), .Y(ori_ori_n472_));
  INV        o0423(.A(ori_ori_n472_), .Y(ori_ori_n473_));
  AOI210     o0424(.A0(ori_ori_n473_), .A1(ori_ori_n467_), .B0(x0), .Y(ori_ori_n474_));
  NOi21      o0425(.An(ori_ori_n159_), .B(ori_ori_n417_), .Y(ori_ori_n475_));
  NA2        o0426(.A(ori_ori_n105_), .B(x1), .Y(ori_ori_n476_));
  NO3        o0427(.A(ori_ori_n476_), .B(ori_ori_n475_), .C(ori_ori_n295_), .Y(ori_ori_n477_));
  OAI210     o0428(.A0(ori_ori_n477_), .A1(ori_ori_n474_), .B0(ori_ori_n462_), .Y(ori_ori_n478_));
  NA2        o0429(.A(ori_ori_n129_), .B(ori_ori_n220_), .Y(ori_ori_n479_));
  OR3        o0430(.A(ori_ori_n479_), .B(ori_ori_n337_), .C(ori_ori_n54_), .Y(ori_ori_n480_));
  OR2        o0431(.A(x6), .B(x0), .Y(ori_ori_n481_));
  NO3        o0432(.A(ori_ori_n481_), .B(x3), .C(x1), .Y(ori_ori_n482_));
  AOI220     o0433(.A0(ori_ori_n482_), .A1(ori_ori_n104_), .B0(ori_ori_n253_), .B1(ori_ori_n247_), .Y(ori_ori_n483_));
  AOI210     o0434(.A0(ori_ori_n483_), .A1(ori_ori_n480_), .B0(ori_ori_n170_), .Y(ori_ori_n484_));
  NA2        o0435(.A(x7), .B(x2), .Y(ori_ori_n485_));
  INV        o0436(.A(ori_ori_n129_), .Y(ori_ori_n486_));
  NA2        o0437(.A(ori_ori_n486_), .B(ori_ori_n82_), .Y(ori_ori_n487_));
  NO2        o0438(.A(ori_ori_n292_), .B(ori_ori_n55_), .Y(ori_ori_n488_));
  NO3        o0439(.A(x3), .B(x1), .C(x0), .Y(ori_ori_n489_));
  OR2        o0440(.A(x6), .B(x1), .Y(ori_ori_n490_));
  NA2        o0441(.A(ori_ori_n490_), .B(x0), .Y(ori_ori_n491_));
  AOI220     o0442(.A0(ori_ori_n491_), .A1(ori_ori_n488_), .B0(ori_ori_n489_), .B1(ori_ori_n425_), .Y(ori_ori_n492_));
  AOI210     o0443(.A0(ori_ori_n492_), .A1(ori_ori_n487_), .B0(ori_ori_n485_), .Y(ori_ori_n493_));
  NA2        o0444(.A(ori_ori_n71_), .B(x0), .Y(ori_ori_n494_));
  NOi31      o0445(.An(ori_ori_n315_), .B(ori_ori_n494_), .C(ori_ori_n238_), .Y(ori_ori_n495_));
  NO4        o0446(.A(ori_ori_n495_), .B(ori_ori_n493_), .C(ori_ori_n484_), .D(ori_ori_n56_), .Y(ori_ori_n496_));
  NA2        o0447(.A(ori_ori_n496_), .B(ori_ori_n478_), .Y(ori_ori_n497_));
  NA3        o0448(.A(x8), .B(x7), .C(x0), .Y(ori_ori_n498_));
  INV        o0449(.A(ori_ori_n498_), .Y(ori_ori_n499_));
  NA2        o0450(.A(ori_ori_n389_), .B(ori_ori_n57_), .Y(ori_ori_n500_));
  NO2        o0451(.A(x8), .B(x0), .Y(ori_ori_n501_));
  NA2        o0452(.A(ori_ori_n501_), .B(ori_ori_n331_), .Y(ori_ori_n502_));
  AOI210     o0453(.A0(ori_ori_n502_), .A1(ori_ori_n500_), .B0(ori_ori_n249_), .Y(ori_ori_n503_));
  NA2        o0454(.A(ori_ori_n503_), .B(ori_ori_n253_), .Y(ori_ori_n504_));
  NO2        o0455(.A(ori_ori_n71_), .B(ori_ori_n106_), .Y(ori_ori_n505_));
  NO2        o0456(.A(ori_ori_n335_), .B(x8), .Y(ori_ori_n506_));
  NO2        o0457(.A(ori_ori_n506_), .B(ori_ori_n239_), .Y(ori_ori_n507_));
  NO3        o0458(.A(ori_ori_n507_), .B(ori_ori_n340_), .C(ori_ori_n244_), .Y(ori_ori_n508_));
  NO2        o0459(.A(ori_ori_n262_), .B(x8), .Y(ori_ori_n509_));
  OAI210     o0460(.A0(ori_ori_n417_), .A1(ori_ori_n299_), .B0(ori_ori_n222_), .Y(ori_ori_n510_));
  NA2        o0461(.A(ori_ori_n318_), .B(ori_ori_n163_), .Y(ori_ori_n511_));
  OAI220     o0462(.A0(ori_ori_n511_), .A1(ori_ori_n59_), .B0(ori_ori_n510_), .B1(ori_ori_n509_), .Y(ori_ori_n512_));
  OAI210     o0463(.A0(ori_ori_n512_), .A1(ori_ori_n508_), .B0(ori_ori_n505_), .Y(ori_ori_n513_));
  NO2        o0464(.A(x8), .B(x2), .Y(ori_ori_n514_));
  NA2        o0465(.A(ori_ori_n296_), .B(ori_ori_n152_), .Y(ori_ori_n515_));
  NO2        o0466(.A(ori_ori_n515_), .B(ori_ori_n105_), .Y(ori_ori_n516_));
  NA2        o0467(.A(ori_ori_n311_), .B(x2), .Y(ori_ori_n517_));
  NO2        o0468(.A(ori_ori_n57_), .B(ori_ori_n53_), .Y(ori_ori_n518_));
  NA2        o0469(.A(ori_ori_n518_), .B(ori_ori_n63_), .Y(ori_ori_n519_));
  AOI210     o0470(.A0(ori_ori_n517_), .A1(ori_ori_n414_), .B0(ori_ori_n519_), .Y(ori_ori_n520_));
  NA2        o0471(.A(ori_ori_n106_), .B(ori_ori_n53_), .Y(ori_ori_n521_));
  NO2        o0472(.A(ori_ori_n521_), .B(x8), .Y(ori_ori_n522_));
  NA2        o0473(.A(x7), .B(ori_ori_n50_), .Y(ori_ori_n523_));
  NO2        o0474(.A(ori_ori_n168_), .B(ori_ori_n523_), .Y(ori_ori_n524_));
  AN2        o0475(.A(ori_ori_n524_), .B(ori_ori_n522_), .Y(ori_ori_n525_));
  NA2        o0476(.A(ori_ori_n363_), .B(ori_ori_n139_), .Y(ori_ori_n526_));
  NO2        o0477(.A(ori_ori_n71_), .B(x2), .Y(ori_ori_n527_));
  NA2        o0478(.A(ori_ori_n527_), .B(ori_ori_n246_), .Y(ori_ori_n528_));
  OAI210     o0479(.A0(ori_ori_n528_), .A1(ori_ori_n526_), .B0(ori_ori_n56_), .Y(ori_ori_n529_));
  NO4        o0480(.A(ori_ori_n529_), .B(ori_ori_n525_), .C(ori_ori_n520_), .D(ori_ori_n516_), .Y(ori_ori_n530_));
  NA3        o0481(.A(ori_ori_n530_), .B(ori_ori_n513_), .C(ori_ori_n504_), .Y(ori_ori_n531_));
  NA2        o0482(.A(ori_ori_n53_), .B(ori_ori_n59_), .Y(ori_ori_n532_));
  NOi21      o0483(.An(x2), .B(x7), .Y(ori_ori_n533_));
  NO2        o0484(.A(x6), .B(x3), .Y(ori_ori_n534_));
  NA2        o0485(.A(ori_ori_n534_), .B(ori_ori_n533_), .Y(ori_ori_n535_));
  NO2        o0486(.A(x6), .B(ori_ori_n59_), .Y(ori_ori_n536_));
  NO3        o0487(.A(ori_ori_n57_), .B(x2), .C(x1), .Y(ori_ori_n537_));
  NO3        o0488(.A(ori_ori_n57_), .B(x2), .C(x0), .Y(ori_ori_n538_));
  AOI220     o0489(.A0(ori_ori_n538_), .A1(ori_ori_n206_), .B0(ori_ori_n537_), .B1(ori_ori_n536_), .Y(ori_ori_n539_));
  OAI210     o0490(.A0(ori_ori_n535_), .A1(ori_ori_n532_), .B0(ori_ori_n539_), .Y(ori_ori_n540_));
  NO2        o0491(.A(ori_ori_n97_), .B(ori_ori_n53_), .Y(ori_ori_n541_));
  NA2        o0492(.A(ori_ori_n201_), .B(ori_ori_n57_), .Y(ori_ori_n542_));
  NA2        o0493(.A(ori_ori_n541_), .B(ori_ori_n542_), .Y(ori_ori_n543_));
  NO3        o0494(.A(ori_ori_n543_), .B(ori_ori_n440_), .C(ori_ori_n59_), .Y(ori_ori_n544_));
  AO210      o0495(.A0(ori_ori_n540_), .A1(ori_ori_n417_), .B0(ori_ori_n544_), .Y(ori_ori_n545_));
  AOI210     o0496(.A0(ori_ori_n531_), .A1(ori_ori_n497_), .B0(ori_ori_n545_), .Y(ori05));
  AOI210     o0497(.A0(ori_ori_n151_), .A1(ori_ori_n55_), .B0(ori_ori_n456_), .Y(ori_ori_n547_));
  OR2        o0498(.A(ori_ori_n547_), .B(ori_ori_n57_), .Y(ori_ori_n548_));
  NO2        o0499(.A(x7), .B(ori_ori_n104_), .Y(ori_ori_n549_));
  NO2        o0500(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n550_));
  NA2        o0501(.A(x5), .B(ori_ori_n56_), .Y(ori_ori_n551_));
  NO2        o0502(.A(ori_ori_n551_), .B(ori_ori_n523_), .Y(ori_ori_n552_));
  AOI210     o0503(.A0(ori_ori_n550_), .A1(ori_ori_n549_), .B0(ori_ori_n552_), .Y(ori_ori_n553_));
  AOI210     o0504(.A0(ori_ori_n553_), .A1(ori_ori_n548_), .B0(ori_ori_n106_), .Y(ori_ori_n554_));
  NO2        o0505(.A(x7), .B(x4), .Y(ori_ori_n555_));
  NO2        o0506(.A(ori_ori_n64_), .B(ori_ori_n55_), .Y(ori_ori_n556_));
  NO2        o0507(.A(ori_ori_n183_), .B(x5), .Y(ori_ori_n557_));
  NA2        o0508(.A(ori_ori_n104_), .B(ori_ori_n106_), .Y(ori_ori_n558_));
  AN2        o0509(.A(ori_ori_n557_), .B(ori_ori_n556_), .Y(ori_ori_n559_));
  OAI210     o0510(.A0(ori_ori_n559_), .A1(ori_ori_n554_), .B0(ori_ori_n444_), .Y(ori_ori_n560_));
  NO2        o0511(.A(x6), .B(ori_ori_n50_), .Y(ori_ori_n561_));
  NA2        o0512(.A(ori_ori_n55_), .B(x4), .Y(ori_ori_n562_));
  NO2        o0513(.A(ori_ori_n104_), .B(ori_ori_n106_), .Y(ori_ori_n563_));
  NA2        o0514(.A(ori_ori_n563_), .B(x7), .Y(ori_ori_n564_));
  NA2        o0515(.A(ori_ori_n392_), .B(ori_ori_n230_), .Y(ori_ori_n565_));
  NO2        o0516(.A(ori_ori_n565_), .B(ori_ori_n562_), .Y(ori_ori_n566_));
  NA2        o0517(.A(ori_ori_n104_), .B(x4), .Y(ori_ori_n567_));
  XO2        o0518(.A(x7), .B(x5), .Y(ori_ori_n568_));
  NO2        o0519(.A(ori_ori_n568_), .B(ori_ori_n53_), .Y(ori_ori_n569_));
  NO2        o0520(.A(ori_ori_n104_), .B(x2), .Y(ori_ori_n570_));
  NO2        o0521(.A(ori_ori_n75_), .B(ori_ori_n55_), .Y(ori_ori_n571_));
  NA2        o0522(.A(ori_ori_n571_), .B(ori_ori_n570_), .Y(ori_ori_n572_));
  INV        o0523(.A(ori_ori_n572_), .Y(ori_ori_n573_));
  OAI210     o0524(.A0(ori_ori_n573_), .A1(ori_ori_n566_), .B0(ori_ori_n561_), .Y(ori_ori_n574_));
  NO2        o0525(.A(ori_ori_n71_), .B(ori_ori_n50_), .Y(ori_ori_n575_));
  NO2        o0526(.A(x5), .B(ori_ori_n56_), .Y(ori_ori_n576_));
  XO2        o0527(.A(x5), .B(x2), .Y(ori_ori_n577_));
  NO3        o0528(.A(x8), .B(x7), .C(ori_ori_n106_), .Y(ori_ori_n578_));
  NA2        o0529(.A(ori_ori_n244_), .B(ori_ori_n533_), .Y(ori_ori_n579_));
  NOi21      o0530(.An(x4), .B(x1), .Y(ori_ori_n580_));
  NA2        o0531(.A(x4), .B(x1), .Y(ori_ori_n581_));
  NO2        o0532(.A(ori_ori_n581_), .B(ori_ori_n50_), .Y(ori_ori_n582_));
  AOI210     o0533(.A0(ori_ori_n582_), .A1(ori_ori_n563_), .B0(ori_ori_n59_), .Y(ori_ori_n583_));
  NA3        o0534(.A(ori_ori_n583_), .B(ori_ori_n574_), .C(ori_ori_n560_), .Y(ori_ori_n584_));
  NA2        o0535(.A(ori_ori_n575_), .B(ori_ori_n56_), .Y(ori_ori_n585_));
  NA2        o0536(.A(ori_ori_n514_), .B(ori_ori_n549_), .Y(ori_ori_n586_));
  NO2        o0537(.A(ori_ori_n586_), .B(ori_ori_n585_), .Y(ori_ori_n587_));
  NA2        o0538(.A(ori_ori_n57_), .B(x6), .Y(ori_ori_n588_));
  INV        o0539(.A(x3), .Y(ori_ori_n589_));
  NA2        o0540(.A(ori_ori_n576_), .B(ori_ori_n143_), .Y(ori_ori_n590_));
  NO3        o0541(.A(ori_ori_n590_), .B(ori_ori_n589_), .C(ori_ori_n382_), .Y(ori_ori_n591_));
  NA2        o0542(.A(ori_ori_n254_), .B(ori_ori_n71_), .Y(ori_ori_n592_));
  NO2        o0543(.A(ori_ori_n346_), .B(x3), .Y(ori_ori_n593_));
  NA2        o0544(.A(ori_ori_n593_), .B(ori_ori_n218_), .Y(ori_ori_n594_));
  INV        o0545(.A(ori_ori_n382_), .Y(ori_ori_n595_));
  NO2        o0546(.A(ori_ori_n421_), .B(ori_ori_n104_), .Y(ori_ori_n596_));
  NO2        o0547(.A(ori_ori_n521_), .B(x6), .Y(ori_ori_n597_));
  NA2        o0548(.A(ori_ori_n597_), .B(ori_ori_n596_), .Y(ori_ori_n598_));
  OAI220     o0549(.A0(ori_ori_n598_), .A1(ori_ori_n595_), .B0(ori_ori_n594_), .B1(ori_ori_n592_), .Y(ori_ori_n599_));
  NO4        o0550(.A(ori_ori_n599_), .B(ori_ori_n591_), .C(x0), .D(ori_ori_n587_), .Y(ori_ori_n600_));
  NA2        o0551(.A(ori_ori_n57_), .B(x5), .Y(ori_ori_n601_));
  NO2        o0552(.A(ori_ori_n601_), .B(x1), .Y(ori_ori_n602_));
  NA2        o0553(.A(x8), .B(ori_ori_n56_), .Y(ori_ori_n603_));
  NO2        o0554(.A(ori_ori_n603_), .B(ori_ori_n124_), .Y(ori_ori_n604_));
  NA2        o0555(.A(x8), .B(x4), .Y(ori_ori_n605_));
  NO2        o0556(.A(x8), .B(x4), .Y(ori_ori_n606_));
  NAi21      o0557(.An(ori_ori_n606_), .B(ori_ori_n605_), .Y(ori_ori_n607_));
  NAi21      o0558(.An(ori_ori_n514_), .B(ori_ori_n346_), .Y(ori_ori_n608_));
  NO4        o0559(.A(ori_ori_n608_), .B(ori_ori_n607_), .C(ori_ori_n382_), .D(ori_ori_n71_), .Y(ori_ori_n609_));
  OAI210     o0560(.A0(ori_ori_n609_), .A1(ori_ori_n604_), .B0(ori_ori_n602_), .Y(ori_ori_n610_));
  NO3        o0561(.A(x8), .B(ori_ori_n104_), .C(x4), .Y(ori_ori_n611_));
  INV        o0562(.A(ori_ori_n611_), .Y(ori_ori_n612_));
  NO2        o0563(.A(ori_ori_n612_), .B(ori_ori_n106_), .Y(ori_ori_n613_));
  NO2        o0564(.A(x5), .B(x4), .Y(ori_ori_n614_));
  NA3        o0565(.A(ori_ori_n614_), .B(ori_ori_n63_), .C(ori_ori_n106_), .Y(ori_ori_n615_));
  NO2        o0566(.A(x6), .B(ori_ori_n106_), .Y(ori_ori_n616_));
  NA2        o0567(.A(ori_ori_n603_), .B(ori_ori_n616_), .Y(ori_ori_n617_));
  OAI210     o0568(.A0(ori_ori_n617_), .A1(ori_ori_n475_), .B0(ori_ori_n615_), .Y(ori_ori_n618_));
  OAI210     o0569(.A0(ori_ori_n618_), .A1(ori_ori_n613_), .B0(ori_ori_n284_), .Y(ori_ori_n619_));
  NA3        o0570(.A(ori_ori_n619_), .B(ori_ori_n610_), .C(ori_ori_n600_), .Y(ori_ori_n620_));
  OR2        o0571(.A(x4), .B(x1), .Y(ori_ori_n621_));
  NO2        o0572(.A(ori_ori_n621_), .B(x3), .Y(ori_ori_n622_));
  NA2        o0573(.A(ori_ori_n55_), .B(x2), .Y(ori_ori_n623_));
  NO3        o0574(.A(ori_ori_n334_), .B(ori_ori_n623_), .C(x6), .Y(ori_ori_n624_));
  AOI220     o0575(.A0(ori_ori_n624_), .A1(ori_ori_n622_), .B0(ori_ori_n620_), .B1(ori_ori_n584_), .Y(ori06));
  NA2        o0576(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n626_));
  NA2        o0577(.A(x6), .B(ori_ori_n106_), .Y(ori_ori_n627_));
  NA2        o0578(.A(ori_ori_n627_), .B(ori_ori_n55_), .Y(ori_ori_n628_));
  NA2        o0579(.A(x5), .B(ori_ori_n59_), .Y(ori_ori_n629_));
  NO2        o0580(.A(ori_ori_n629_), .B(ori_ori_n114_), .Y(ori_ori_n630_));
  NA3        o0581(.A(ori_ori_n630_), .B(ori_ori_n628_), .C(ori_ori_n450_), .Y(ori_ori_n631_));
  NO2        o0582(.A(ori_ori_n346_), .B(x0), .Y(ori_ori_n632_));
  NA2        o0583(.A(ori_ori_n310_), .B(x2), .Y(ori_ori_n633_));
  NOi21      o0584(.An(x6), .B(x8), .Y(ori_ori_n634_));
  NO2        o0585(.A(ori_ori_n631_), .B(ori_ori_n626_), .Y(ori_ori_n635_));
  NA2        o0586(.A(ori_ori_n56_), .B(ori_ori_n50_), .Y(ori_ori_n636_));
  NA2        o0587(.A(ori_ori_n333_), .B(ori_ori_n323_), .Y(ori_ori_n637_));
  NO2        o0588(.A(ori_ori_n71_), .B(ori_ori_n104_), .Y(ori_ori_n638_));
  NO2        o0589(.A(ori_ori_n53_), .B(ori_ori_n59_), .Y(ori_ori_n639_));
  NO4        o0590(.A(ori_ori_n639_), .B(ori_ori_n623_), .C(ori_ori_n638_), .D(ori_ori_n444_), .Y(ori_ori_n640_));
  AOI220     o0591(.A0(ori_ori_n640_), .A1(ori_ori_n637_), .B0(ori_ori_n379_), .B1(ori_ori_n63_), .Y(ori_ori_n641_));
  NO2        o0592(.A(ori_ori_n641_), .B(ori_ori_n636_), .Y(ori_ori_n642_));
  NO2        o0593(.A(ori_ori_n54_), .B(x0), .Y(ori_ori_n643_));
  NA2        o0594(.A(x4), .B(x3), .Y(ori_ori_n644_));
  OAI210     o0595(.A0(ori_ori_n644_), .A1(x8), .B0(ori_ori_n468_), .Y(ori_ori_n645_));
  NA2        o0596(.A(ori_ori_n645_), .B(ori_ori_n643_), .Y(ori_ori_n646_));
  NO2        o0597(.A(ori_ori_n100_), .B(ori_ori_n56_), .Y(ori_ori_n647_));
  NA3        o0598(.A(ori_ori_n647_), .B(ori_ori_n231_), .C(ori_ori_n363_), .Y(ori_ori_n648_));
  AOI210     o0599(.A0(ori_ori_n648_), .A1(ori_ori_n646_), .B0(x2), .Y(ori_ori_n649_));
  INV        o0600(.A(ori_ori_n342_), .Y(ori_ori_n650_));
  NO2        o0601(.A(ori_ori_n366_), .B(x8), .Y(ori_ori_n651_));
  NO2        o0602(.A(ori_ori_n232_), .B(ori_ori_n470_), .Y(ori_ori_n652_));
  AOI210     o0603(.A0(ori_ori_n651_), .A1(ori_ori_n240_), .B0(ori_ori_n652_), .Y(ori_ori_n653_));
  NO2        o0604(.A(x5), .B(x3), .Y(ori_ori_n654_));
  NA3        o0605(.A(ori_ori_n501_), .B(ori_ori_n654_), .C(x1), .Y(ori_ori_n655_));
  OR2        o0606(.A(ori_ori_n655_), .B(ori_ori_n450_), .Y(ori_ori_n656_));
  OAI210     o0607(.A0(ori_ori_n653_), .A1(ori_ori_n650_), .B0(ori_ori_n656_), .Y(ori_ori_n657_));
  OR4        o0608(.A(ori_ori_n657_), .B(ori_ori_n649_), .C(ori_ori_n642_), .D(ori_ori_n635_), .Y(ori_ori_n658_));
  NA2        o0609(.A(x7), .B(ori_ori_n56_), .Y(ori_ori_n659_));
  NO2        o0610(.A(ori_ori_n563_), .B(ori_ori_n59_), .Y(ori_ori_n660_));
  NO2        o0611(.A(ori_ori_n157_), .B(x6), .Y(ori_ori_n661_));
  AN2        o0612(.A(ori_ori_n426_), .B(ori_ori_n293_), .Y(ori_ori_n662_));
  NA2        o0613(.A(ori_ori_n662_), .B(ori_ori_n318_), .Y(ori_ori_n663_));
  NO2        o0614(.A(ori_ori_n280_), .B(ori_ori_n104_), .Y(ori_ori_n664_));
  NO2        o0615(.A(ori_ori_n56_), .B(x3), .Y(ori_ori_n665_));
  NA2        o0616(.A(ori_ori_n665_), .B(ori_ori_n71_), .Y(ori_ori_n666_));
  NO2        o0617(.A(ori_ori_n666_), .B(ori_ori_n227_), .Y(ori_ori_n667_));
  NO2        o0618(.A(ori_ori_n71_), .B(x3), .Y(ori_ori_n668_));
  NA3        o0619(.A(ori_ori_n668_), .B(ori_ori_n518_), .C(ori_ori_n56_), .Y(ori_ori_n669_));
  NO2        o0620(.A(ori_ori_n57_), .B(x6), .Y(ori_ori_n670_));
  INV        o0621(.A(ori_ori_n669_), .Y(ori_ori_n671_));
  OR3        o0622(.A(ori_ori_n671_), .B(ori_ori_n667_), .C(ori_ori_n582_), .Y(ori_ori_n672_));
  NA2        o0623(.A(ori_ori_n672_), .B(ori_ori_n664_), .Y(ori_ori_n673_));
  NA2        o0624(.A(x7), .B(x6), .Y(ori_ori_n674_));
  NA3        o0625(.A(x2), .B(x1), .C(x0), .Y(ori_ori_n675_));
  NO3        o0626(.A(ori_ori_n675_), .B(ori_ori_n674_), .C(ori_ori_n547_), .Y(ori_ori_n676_));
  NA2        o0627(.A(ori_ori_n445_), .B(ori_ori_n138_), .Y(ori_ori_n677_));
  NO2        o0628(.A(x5), .B(x1), .Y(ori_ori_n678_));
  NA2        o0629(.A(ori_ori_n678_), .B(ori_ori_n670_), .Y(ori_ori_n679_));
  NA2        o0630(.A(x4), .B(x0), .Y(ori_ori_n680_));
  NO3        o0631(.A(ori_ori_n57_), .B(x6), .C(x2), .Y(ori_ori_n681_));
  NA2        o0632(.A(ori_ori_n681_), .B(ori_ori_n205_), .Y(ori_ori_n682_));
  NO2        o0633(.A(ori_ori_n682_), .B(ori_ori_n680_), .Y(ori_ori_n683_));
  NO2        o0634(.A(ori_ori_n683_), .B(ori_ori_n676_), .Y(ori_ori_n684_));
  NA3        o0635(.A(ori_ori_n684_), .B(ori_ori_n673_), .C(ori_ori_n663_), .Y(ori_ori_n685_));
  AOI210     o0636(.A0(ori_ori_n658_), .A1(ori_ori_n57_), .B0(ori_ori_n685_), .Y(ori07));
  NA2        o0637(.A(ori_ori_n104_), .B(ori_ori_n59_), .Y(ori_ori_n687_));
  NOi21      o0638(.An(ori_ori_n674_), .B(ori_ori_n112_), .Y(ori_ori_n688_));
  NO3        o0639(.A(ori_ori_n57_), .B(x5), .C(x1), .Y(ori_ori_n689_));
  NA2        o0640(.A(ori_ori_n689_), .B(ori_ori_n336_), .Y(ori_ori_n690_));
  NO2        o0641(.A(ori_ori_n57_), .B(ori_ori_n71_), .Y(ori_ori_n691_));
  NO2        o0642(.A(ori_ori_n142_), .B(ori_ori_n105_), .Y(ori_ori_n692_));
  NAi21      o0643(.An(ori_ori_n143_), .B(ori_ori_n144_), .Y(ori_ori_n693_));
  NA3        o0644(.A(ori_ori_n693_), .B(ori_ori_n89_), .C(x3), .Y(ori_ori_n694_));
  NO3        o0645(.A(ori_ori_n55_), .B(x3), .C(x1), .Y(ori_ori_n695_));
  NO2        o0646(.A(ori_ori_n463_), .B(x2), .Y(ori_ori_n696_));
  AOI210     o0647(.A0(ori_ori_n696_), .A1(ori_ori_n465_), .B0(ori_ori_n695_), .Y(ori_ori_n697_));
  OAI210     o0648(.A0(ori_ori_n697_), .A1(ori_ori_n588_), .B0(ori_ori_n694_), .Y(ori_ori_n698_));
  NO2        o0649(.A(x8), .B(ori_ori_n53_), .Y(ori_ori_n699_));
  NA2        o0650(.A(ori_ori_n699_), .B(ori_ori_n59_), .Y(ori_ori_n700_));
  NO2        o0651(.A(x7), .B(x3), .Y(ori_ori_n701_));
  NA2        o0652(.A(ori_ori_n701_), .B(ori_ori_n97_), .Y(ori_ori_n702_));
  NO2        o0653(.A(ori_ori_n700_), .B(ori_ori_n702_), .Y(ori_ori_n703_));
  AOI210     o0654(.A0(ori_ori_n698_), .A1(ori_ori_n226_), .B0(ori_ori_n703_), .Y(ori_ori_n704_));
  NO2        o0655(.A(ori_ori_n704_), .B(x4), .Y(ori_ori_n705_));
  NO2        o0656(.A(ori_ori_n543_), .B(ori_ori_n106_), .Y(ori_ori_n706_));
  XO2        o0657(.A(x5), .B(x1), .Y(ori_ori_n707_));
  NO4        o0658(.A(ori_ori_n707_), .B(ori_ori_n152_), .C(ori_ori_n190_), .D(ori_ori_n55_), .Y(ori_ori_n708_));
  OAI210     o0659(.A0(ori_ori_n708_), .A1(ori_ori_n706_), .B0(ori_ori_n370_), .Y(ori_ori_n709_));
  NO3        o0660(.A(ori_ori_n50_), .B(x2), .C(x0), .Y(ori_ori_n710_));
  NO2        o0661(.A(ori_ori_n283_), .B(ori_ori_n104_), .Y(ori_ori_n711_));
  NA2        o0662(.A(x6), .B(x0), .Y(ori_ori_n712_));
  NO2        o0663(.A(ori_ori_n623_), .B(ori_ori_n712_), .Y(ori_ori_n713_));
  NO2        o0664(.A(ori_ori_n707_), .B(ori_ori_n634_), .Y(ori_ori_n714_));
  OAI210     o0665(.A0(ori_ori_n678_), .A1(ori_ori_n63_), .B0(ori_ori_n57_), .Y(ori_ori_n715_));
  OAI210     o0666(.A0(ori_ori_n715_), .A1(ori_ori_n714_), .B0(ori_ori_n690_), .Y(ori_ori_n716_));
  AOI220     o0667(.A0(ori_ori_n716_), .A1(ori_ori_n710_), .B0(ori_ori_n713_), .B1(ori_ori_n711_), .Y(ori_ori_n717_));
  AOI210     o0668(.A0(ori_ori_n717_), .A1(ori_ori_n709_), .B0(ori_ori_n56_), .Y(ori_ori_n718_));
  NOi21      o0669(.An(ori_ori_n212_), .B(ori_ori_n336_), .Y(ori_ori_n719_));
  NO2        o0670(.A(ori_ori_n719_), .B(ori_ori_n219_), .Y(ori_ori_n720_));
  NO2        o0671(.A(ori_ori_n283_), .B(x6), .Y(ori_ori_n721_));
  AN2        o0672(.A(ori_ori_n721_), .B(ori_ori_n300_), .Y(ori_ori_n722_));
  OAI210     o0673(.A0(ori_ori_n722_), .A1(ori_ori_n720_), .B0(ori_ori_n59_), .Y(ori_ori_n723_));
  NA2        o0674(.A(ori_ori_n90_), .B(ori_ori_n71_), .Y(ori_ori_n724_));
  NO2        o0675(.A(ori_ori_n724_), .B(ori_ori_n586_), .Y(ori_ori_n725_));
  NAi21      o0676(.An(x8), .B(x7), .Y(ori_ori_n726_));
  NA2        o0677(.A(ori_ori_n719_), .B(ori_ori_n726_), .Y(ori_ori_n727_));
  NA2        o0678(.A(ori_ori_n363_), .B(ori_ori_n106_), .Y(ori_ori_n728_));
  NO2        o0679(.A(ori_ori_n634_), .B(x1), .Y(ori_ori_n729_));
  NO3        o0680(.A(ori_ori_n729_), .B(ori_ori_n728_), .C(ori_ori_n518_), .Y(ori_ori_n730_));
  AOI210     o0681(.A0(ori_ori_n730_), .A1(ori_ori_n727_), .B0(ori_ori_n725_), .Y(ori_ori_n731_));
  AOI210     o0682(.A0(ori_ori_n731_), .A1(ori_ori_n723_), .B0(ori_ori_n133_), .Y(ori_ori_n732_));
  NO2        o0683(.A(x8), .B(x7), .Y(ori_ori_n733_));
  NO2        o0684(.A(ori_ori_n733_), .B(x3), .Y(ori_ori_n734_));
  NA3        o0685(.A(ori_ori_n734_), .B(ori_ori_n331_), .C(x1), .Y(ori_ori_n735_));
  NO2        o0686(.A(x8), .B(ori_ori_n106_), .Y(ori_ori_n736_));
  NA2        o0687(.A(ori_ori_n736_), .B(ori_ori_n230_), .Y(ori_ori_n737_));
  NO2        o0688(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n738_));
  NA2        o0689(.A(ori_ori_n738_), .B(ori_ori_n277_), .Y(ori_ori_n739_));
  AOI210     o0690(.A0(ori_ori_n737_), .A1(ori_ori_n735_), .B0(ori_ori_n739_), .Y(ori_ori_n740_));
  NO4        o0691(.A(ori_ori_n740_), .B(ori_ori_n732_), .C(ori_ori_n718_), .D(ori_ori_n705_), .Y(ori08));
  NA2        o0692(.A(ori_ori_n50_), .B(x1), .Y(ori_ori_n742_));
  XN2        o0693(.A(x5), .B(x4), .Y(ori_ori_n743_));
  INV        o0694(.A(ori_ori_n743_), .Y(ori_ori_n744_));
  NA2        o0695(.A(ori_ori_n744_), .B(ori_ori_n324_), .Y(ori_ori_n745_));
  NO2        o0696(.A(ori_ori_n220_), .B(ori_ori_n104_), .Y(ori_ori_n746_));
  AOI210     o0697(.A0(ori_ori_n746_), .A1(ori_ori_n251_), .B0(ori_ori_n176_), .Y(ori_ori_n747_));
  OAI220     o0698(.A0(ori_ori_n747_), .A1(x4), .B0(ori_ori_n745_), .B1(ori_ori_n742_), .Y(ori_ori_n748_));
  NA2        o0699(.A(ori_ori_n748_), .B(ori_ori_n246_), .Y(ori_ori_n749_));
  NO2        o0700(.A(ori_ori_n728_), .B(ori_ori_n562_), .Y(ori_ori_n750_));
  NA2        o0701(.A(ori_ori_n251_), .B(ori_ori_n138_), .Y(ori_ori_n751_));
  NA2        o0702(.A(ori_ori_n133_), .B(x7), .Y(ori_ori_n752_));
  OR3        o0703(.A(ori_ori_n675_), .B(ori_ori_n421_), .C(ori_ori_n654_), .Y(ori_ori_n753_));
  OAI220     o0704(.A0(ori_ori_n753_), .A1(ori_ori_n752_), .B0(ori_ori_n751_), .B1(ori_ori_n188_), .Y(ori_ori_n754_));
  AOI210     o0705(.A0(ori_ori_n750_), .A1(ori_ori_n265_), .B0(ori_ori_n754_), .Y(ori_ori_n755_));
  AOI210     o0706(.A0(ori_ori_n755_), .A1(ori_ori_n749_), .B0(ori_ori_n71_), .Y(ori_ori_n756_));
  NO2        o0707(.A(ori_ori_n733_), .B(ori_ori_n106_), .Y(ori_ori_n757_));
  INV        o0708(.A(ori_ori_n757_), .Y(ori_ori_n758_));
  NA2        o0709(.A(ori_ori_n366_), .B(ori_ori_n313_), .Y(ori_ori_n759_));
  NA2        o0710(.A(ori_ori_n392_), .B(ori_ori_n213_), .Y(ori_ori_n760_));
  NA2        o0711(.A(ori_ori_n651_), .B(ori_ori_n103_), .Y(ori_ori_n761_));
  OAI220     o0712(.A0(ori_ori_n761_), .A1(ori_ori_n760_), .B0(ori_ori_n759_), .B1(ori_ori_n758_), .Y(ori_ori_n762_));
  NA2        o0713(.A(ori_ori_n762_), .B(ori_ori_n261_), .Y(ori_ori_n763_));
  NA2        o0714(.A(ori_ori_n304_), .B(ori_ori_n53_), .Y(ori_ori_n764_));
  NO3        o0715(.A(ori_ori_n366_), .B(ori_ori_n129_), .C(ori_ori_n68_), .Y(ori_ori_n765_));
  NO2        o0716(.A(ori_ori_n639_), .B(ori_ori_n222_), .Y(ori_ori_n766_));
  NO2        o0717(.A(ori_ori_n422_), .B(ori_ori_n95_), .Y(ori_ori_n767_));
  AO220      o0718(.A0(ori_ori_n767_), .A1(ori_ori_n766_), .B0(ori_ori_n765_), .B1(ori_ori_n764_), .Y(ori_ori_n768_));
  NA2        o0719(.A(x7), .B(ori_ori_n59_), .Y(ori_ori_n769_));
  NO2        o0720(.A(ori_ori_n286_), .B(ori_ori_n769_), .Y(ori_ori_n770_));
  AOI210     o0721(.A0(ori_ori_n768_), .A1(x5), .B0(ori_ori_n770_), .Y(ori_ori_n771_));
  AOI210     o0722(.A0(ori_ori_n771_), .A1(ori_ori_n763_), .B0(ori_ori_n72_), .Y(ori_ori_n772_));
  NO2        o0723(.A(ori_ori_n70_), .B(x3), .Y(ori_ori_n773_));
  NA2        o0724(.A(ori_ori_n773_), .B(ori_ori_n136_), .Y(ori_ori_n774_));
  MUX2       o0725(.S(x3), .A(ori_ori_n152_), .B(ori_ori_n693_), .Y(ori_ori_n775_));
  NA2        o0726(.A(ori_ori_n775_), .B(ori_ori_n506_), .Y(ori_ori_n776_));
  NO3        o0727(.A(x6), .B(x4), .C(x0), .Y(ori_ori_n777_));
  INV        o0728(.A(ori_ori_n777_), .Y(ori_ori_n778_));
  AOI210     o0729(.A0(ori_ori_n776_), .A1(ori_ori_n774_), .B0(ori_ori_n778_), .Y(ori_ori_n779_));
  NO3        o0730(.A(x5), .B(x3), .C(ori_ori_n106_), .Y(ori_ori_n780_));
  AOI220     o0731(.A0(ori_ori_n744_), .A1(ori_ori_n282_), .B0(ori_ori_n780_), .B1(ori_ori_n59_), .Y(ori_ori_n781_));
  OR2        o0732(.A(x8), .B(x1), .Y(ori_ori_n782_));
  NO3        o0733(.A(ori_ori_n782_), .B(ori_ori_n781_), .C(ori_ori_n665_), .Y(ori_ori_n783_));
  NAi21      o0734(.An(x4), .B(x1), .Y(ori_ori_n784_));
  NO2        o0735(.A(ori_ori_n784_), .B(x0), .Y(ori_ori_n785_));
  NA2        o0736(.A(ori_ori_n557_), .B(ori_ori_n785_), .Y(ori_ori_n786_));
  NA3        o0737(.A(ori_ori_n55_), .B(x1), .C(x0), .Y(ori_ori_n787_));
  OAI210     o0738(.A0(ori_ori_n787_), .A1(ori_ori_n650_), .B0(ori_ori_n786_), .Y(ori_ori_n788_));
  OAI210     o0739(.A0(ori_ori_n788_), .A1(ori_ori_n783_), .B0(ori_ori_n291_), .Y(ori_ori_n789_));
  AO210      o0740(.A0(ori_ori_n263_), .A1(ori_ori_n239_), .B0(ori_ori_n664_), .Y(ori_ori_n790_));
  NA2        o0741(.A(ori_ori_n104_), .B(ori_ori_n56_), .Y(ori_ori_n791_));
  NO2        o0742(.A(ori_ori_n57_), .B(x2), .Y(ori_ori_n792_));
  NA2        o0743(.A(ori_ori_n790_), .B(ori_ori_n582_), .Y(ori_ori_n793_));
  NA2        o0744(.A(ori_ori_n793_), .B(ori_ori_n789_), .Y(ori_ori_n794_));
  NO4        o0745(.A(ori_ori_n794_), .B(ori_ori_n779_), .C(ori_ori_n772_), .D(ori_ori_n756_), .Y(ori09));
  NO3        o0746(.A(ori_ori_n707_), .B(ori_ori_n116_), .C(ori_ori_n92_), .Y(ori_ori_n796_));
  AOI220     o0747(.A0(ori_ori_n272_), .A1(ori_ori_n70_), .B0(ori_ori_n533_), .B1(ori_ori_n490_), .Y(ori_ori_n797_));
  OAI210     o0748(.A0(ori_ori_n796_), .A1(x2), .B0(ori_ori_n797_), .Y(ori_ori_n798_));
  AOI210     o0749(.A0(ori_ori_n798_), .A1(ori_ori_n679_), .B0(ori_ori_n400_), .Y(ori_ori_n799_));
  NO2        o0750(.A(ori_ori_n532_), .B(ori_ori_n238_), .Y(ori_ori_n800_));
  INV        o0751(.A(ori_ori_n310_), .Y(ori_ori_n801_));
  NO3        o0752(.A(ori_ori_n549_), .B(ori_ori_n98_), .C(ori_ori_n106_), .Y(ori_ori_n802_));
  AO220      o0753(.A0(ori_ori_n802_), .A1(ori_ori_n801_), .B0(ori_ori_n800_), .B1(ori_ori_n563_), .Y(ori_ori_n803_));
  OAI210     o0754(.A0(ori_ori_n803_), .A1(ori_ori_n799_), .B0(x4), .Y(ori_ori_n804_));
  NO2        o0755(.A(ori_ori_n351_), .B(ori_ori_n253_), .Y(ori_ori_n805_));
  NO2        o0756(.A(ori_ori_n175_), .B(ori_ori_n104_), .Y(ori_ori_n806_));
  NA2        o0757(.A(ori_ori_n805_), .B(ori_ori_n569_), .Y(ori_ori_n807_));
  NO2        o0758(.A(ori_ori_n707_), .B(ori_ori_n92_), .Y(ori_ori_n808_));
  NAi21      o0759(.An(x0), .B(x2), .Y(ori_ori_n809_));
  NO2        o0760(.A(ori_ori_n276_), .B(ori_ori_n809_), .Y(ori_ori_n810_));
  OAI210     o0761(.A0(ori_ori_n431_), .A1(ori_ori_n248_), .B0(ori_ori_n175_), .Y(ori_ori_n811_));
  AOI210     o0762(.A0(ori_ori_n154_), .A1(ori_ori_n726_), .B0(ori_ori_n323_), .Y(ori_ori_n812_));
  AOI220     o0763(.A0(ori_ori_n812_), .A1(ori_ori_n811_), .B0(ori_ori_n810_), .B1(ori_ori_n808_), .Y(ori_ori_n813_));
  OAI210     o0764(.A0(ori_ori_n807_), .A1(ori_ori_n55_), .B0(ori_ori_n813_), .Y(ori_ori_n814_));
  NA2        o0765(.A(ori_ori_n814_), .B(ori_ori_n56_), .Y(ori_ori_n815_));
  NO2        o0766(.A(ori_ori_n56_), .B(ori_ori_n59_), .Y(ori_ori_n816_));
  INV        o0767(.A(ori_ori_n121_), .Y(ori_ori_n817_));
  NA2        o0768(.A(ori_ori_n678_), .B(ori_ori_n55_), .Y(ori_ori_n818_));
  AOI210     o0769(.A0(x6), .A1(x1), .B0(x5), .Y(ori_ori_n819_));
  OAI210     o0770(.A0(ori_ori_n819_), .A1(ori_ori_n303_), .B0(x2), .Y(ori_ori_n820_));
  AOI210     o0771(.A0(ori_ori_n820_), .A1(ori_ori_n818_), .B0(ori_ori_n817_), .Y(ori_ori_n821_));
  NA2        o0772(.A(ori_ori_n505_), .B(ori_ori_n55_), .Y(ori_ori_n822_));
  NO2        o0773(.A(ori_ori_n211_), .B(ori_ori_n343_), .Y(ori_ori_n823_));
  NO2        o0774(.A(ori_ori_n283_), .B(ori_ori_n137_), .Y(ori_ori_n824_));
  INV        o0775(.A(ori_ori_n824_), .Y(ori_ori_n825_));
  OAI220     o0776(.A0(ori_ori_n825_), .A1(ori_ori_n55_), .B0(ori_ori_n822_), .B1(ori_ori_n412_), .Y(ori_ori_n826_));
  OAI210     o0777(.A0(ori_ori_n826_), .A1(ori_ori_n821_), .B0(ori_ori_n816_), .Y(ori_ori_n827_));
  NO2        o0778(.A(ori_ori_n359_), .B(ori_ori_n104_), .Y(ori_ori_n828_));
  NO2        o0779(.A(ori_ori_n304_), .B(ori_ori_n444_), .Y(ori_ori_n829_));
  AOI220     o0780(.A0(ori_ori_n829_), .A1(ori_ori_n828_), .B0(ori_ori_n191_), .B1(ori_ori_n209_), .Y(ori_ori_n830_));
  NA4        o0781(.A(ori_ori_n830_), .B(ori_ori_n827_), .C(ori_ori_n815_), .D(ori_ori_n804_), .Y(ori_ori_n831_));
  NA2        o0782(.A(ori_ori_n831_), .B(ori_ori_n50_), .Y(ori_ori_n832_));
  NO2        o0783(.A(ori_ori_n338_), .B(ori_ori_n148_), .Y(ori_ori_n833_));
  NO2        o0784(.A(ori_ori_n387_), .B(ori_ori_n736_), .Y(ori_ori_n834_));
  OAI210     o0785(.A0(ori_ori_n834_), .A1(ori_ori_n833_), .B0(x0), .Y(ori_ori_n835_));
  NO3        o0786(.A(x8), .B(x7), .C(x2), .Y(ori_ori_n836_));
  NO3        o0787(.A(ori_ori_n57_), .B(x5), .C(x2), .Y(ori_ori_n837_));
  OAI210     o0788(.A0(ori_ori_n837_), .A1(ori_ori_n836_), .B0(ori_ori_n465_), .Y(ori_ori_n838_));
  AOI210     o0789(.A0(ori_ori_n838_), .A1(ori_ori_n835_), .B0(x4), .Y(ori_ori_n839_));
  NO2        o0790(.A(ori_ori_n380_), .B(ori_ori_n136_), .Y(ori_ori_n840_));
  NO2        o0791(.A(ori_ori_n104_), .B(ori_ori_n56_), .Y(ori_ori_n841_));
  NA2        o0792(.A(ori_ori_n841_), .B(x8), .Y(ori_ori_n842_));
  OAI210     o0793(.A0(ori_ori_n840_), .A1(ori_ori_n839_), .B0(ori_ori_n561_), .Y(ori_ori_n843_));
  NO2        o0794(.A(ori_ori_n234_), .B(ori_ori_n115_), .Y(ori_ori_n844_));
  OAI210     o0795(.A0(x4), .A1(x2), .B0(x0), .Y(ori_ori_n845_));
  NA3        o0796(.A(ori_ori_n551_), .B(ori_ori_n562_), .C(ori_ori_n314_), .Y(ori_ori_n846_));
  OAI210     o0797(.A0(ori_ori_n845_), .A1(ori_ori_n260_), .B0(ori_ori_n53_), .Y(ori_ori_n847_));
  AOI210     o0798(.A0(ori_ori_n846_), .A1(ori_ori_n845_), .B0(ori_ori_n847_), .Y(ori_ori_n848_));
  OAI210     o0799(.A0(ori_ori_n848_), .A1(ori_ori_n844_), .B0(ori_ori_n299_), .Y(ori_ori_n849_));
  AOI220     o0800(.A0(ori_ori_n605_), .A1(ori_ori_n316_), .B0(ori_ori_n318_), .B1(ori_ori_n91_), .Y(ori_ori_n850_));
  NA2        o0801(.A(ori_ori_n91_), .B(x5), .Y(ori_ori_n851_));
  NO2        o0802(.A(ori_ori_n850_), .B(ori_ori_n292_), .Y(ori_ori_n852_));
  NA2        o0803(.A(ori_ori_n852_), .B(ori_ori_n68_), .Y(ori_ori_n853_));
  NA2        o0804(.A(ori_ori_n363_), .B(ori_ori_n693_), .Y(ori_ori_n854_));
  NA2        o0805(.A(ori_ori_n226_), .B(ori_ori_n152_), .Y(ori_ori_n855_));
  AO210      o0806(.A0(ori_ori_n855_), .A1(ori_ori_n854_), .B0(ori_ori_n126_), .Y(ori_ori_n856_));
  NO2        o0807(.A(ori_ori_n393_), .B(x2), .Y(ori_ori_n857_));
  NO2        o0808(.A(x7), .B(ori_ori_n53_), .Y(ori_ori_n858_));
  NA2        o0809(.A(ori_ori_n858_), .B(x5), .Y(ori_ori_n859_));
  NO2        o0810(.A(ori_ori_n859_), .B(ori_ori_n60_), .Y(ori_ori_n860_));
  AOI220     o0811(.A0(ori_ori_n860_), .A1(ori_ori_n857_), .B0(ori_ori_n606_), .B1(ori_ori_n221_), .Y(ori_ori_n861_));
  NA4        o0812(.A(ori_ori_n861_), .B(ori_ori_n856_), .C(ori_ori_n853_), .D(ori_ori_n849_), .Y(ori_ori_n862_));
  NO4        o0813(.A(ori_ori_n846_), .B(ori_ori_n576_), .C(ori_ori_n412_), .D(ori_ori_n50_), .Y(ori_ori_n863_));
  AOI220     o0814(.A0(ori_ori_n550_), .A1(ori_ori_n549_), .B0(ori_ori_n254_), .B1(x5), .Y(ori_ori_n864_));
  NO2        o0815(.A(ori_ori_n614_), .B(ori_ori_n175_), .Y(ori_ori_n865_));
  NA3        o0816(.A(ori_ori_n865_), .B(ori_ori_n607_), .C(x7), .Y(ori_ori_n866_));
  OAI210     o0817(.A0(ori_ori_n864_), .A1(ori_ori_n317_), .B0(ori_ori_n866_), .Y(ori_ori_n867_));
  OAI210     o0818(.A0(ori_ori_n867_), .A1(ori_ori_n863_), .B0(ori_ori_n82_), .Y(ori_ori_n868_));
  NA2        o0819(.A(ori_ori_n699_), .B(x2), .Y(ori_ori_n869_));
  NO2        o0820(.A(ori_ori_n869_), .B(ori_ori_n58_), .Y(ori_ori_n870_));
  NO2        o0821(.A(x5), .B(ori_ori_n53_), .Y(ori_ori_n871_));
  NAi21      o0822(.An(x1), .B(x4), .Y(ori_ori_n872_));
  NA2        o0823(.A(ori_ori_n872_), .B(ori_ori_n784_), .Y(ori_ori_n873_));
  NO3        o0824(.A(ori_ori_n873_), .B(ori_ori_n185_), .C(ori_ori_n871_), .Y(ori_ori_n874_));
  OAI210     o0825(.A0(ori_ori_n874_), .A1(ori_ori_n870_), .B0(ori_ori_n370_), .Y(ori_ori_n875_));
  NA2        o0826(.A(ori_ori_n875_), .B(ori_ori_n868_), .Y(ori_ori_n876_));
  AOI210     o0827(.A0(ori_ori_n862_), .A1(x6), .B0(ori_ori_n876_), .Y(ori_ori_n877_));
  NA3        o0828(.A(ori_ori_n877_), .B(ori_ori_n843_), .C(ori_ori_n832_), .Y(ori10));
  NO2        o0829(.A(x4), .B(x1), .Y(ori_ori_n879_));
  NO2        o0830(.A(ori_ori_n879_), .B(ori_ori_n138_), .Y(ori_ori_n880_));
  NA3        o0831(.A(x5), .B(x4), .C(x0), .Y(ori_ori_n881_));
  OAI220     o0832(.A0(ori_ori_n881_), .A1(ori_ori_n249_), .B0(ori_ori_n639_), .B1(ori_ori_n224_), .Y(ori_ori_n882_));
  NA2        o0833(.A(ori_ori_n882_), .B(ori_ori_n880_), .Y(ori_ori_n883_));
  NO3        o0834(.A(ori_ori_n324_), .B(ori_ori_n292_), .C(ori_ori_n90_), .Y(ori_ori_n884_));
  NA3        o0835(.A(ori_ori_n884_), .B(ori_ori_n341_), .C(ori_ori_n62_), .Y(ori_ori_n885_));
  AOI210     o0836(.A0(ori_ori_n885_), .A1(ori_ori_n883_), .B0(ori_ori_n276_), .Y(ori_ori_n886_));
  NOi21      o0837(.An(ori_ori_n233_), .B(ori_ori_n130_), .Y(ori_ori_n887_));
  AOI210     o0838(.A0(ori_ori_n451_), .A1(ori_ori_n563_), .B0(ori_ori_n300_), .Y(ori_ori_n888_));
  NO2        o0839(.A(ori_ori_n816_), .B(ori_ori_n312_), .Y(ori_ori_n889_));
  NOi31      o0840(.An(ori_ori_n889_), .B(ori_ori_n888_), .C(ori_ori_n887_), .Y(ori_ori_n890_));
  NA2        o0841(.A(x4), .B(ori_ori_n106_), .Y(ori_ori_n891_));
  NO2        o0842(.A(ori_ori_n295_), .B(ori_ori_n891_), .Y(ori_ori_n892_));
  NA2        o0843(.A(ori_ori_n95_), .B(x5), .Y(ori_ori_n893_));
  NO3        o0844(.A(ori_ori_n893_), .B(ori_ori_n107_), .C(ori_ori_n55_), .Y(ori_ori_n894_));
  NO3        o0845(.A(ori_ori_n894_), .B(ori_ori_n892_), .C(ori_ori_n890_), .Y(ori_ori_n895_));
  NA2        o0846(.A(ori_ori_n871_), .B(ori_ori_n50_), .Y(ori_ori_n896_));
  NA2        o0847(.A(ori_ori_n550_), .B(ori_ori_n245_), .Y(ori_ori_n897_));
  NO2        o0848(.A(ori_ori_n897_), .B(ori_ori_n896_), .Y(ori_ori_n898_));
  OAI220     o0849(.A0(ori_ori_n842_), .A1(ori_ori_n103_), .B0(ori_ori_n791_), .B1(ori_ori_n400_), .Y(ori_ori_n899_));
  AOI210     o0850(.A0(ori_ori_n899_), .A1(ori_ori_n251_), .B0(ori_ori_n898_), .Y(ori_ori_n900_));
  OAI210     o0851(.A0(ori_ori_n895_), .A1(ori_ori_n343_), .B0(ori_ori_n900_), .Y(ori_ori_n901_));
  OAI210     o0852(.A0(ori_ori_n901_), .A1(ori_ori_n886_), .B0(x7), .Y(ori_ori_n902_));
  NA2        o0853(.A(ori_ori_n55_), .B(ori_ori_n71_), .Y(ori_ori_n903_));
  AOI210     o0854(.A0(ori_ori_n400_), .A1(ori_ori_n323_), .B0(ori_ori_n891_), .Y(ori_ori_n904_));
  NO3        o0855(.A(ori_ori_n402_), .B(ori_ori_n809_), .C(x5), .Y(ori_ori_n905_));
  OAI210     o0856(.A0(ori_ori_n905_), .A1(ori_ori_n904_), .B0(ori_ori_n903_), .Y(ori_ori_n906_));
  NO2        o0857(.A(ori_ori_n324_), .B(ori_ori_n132_), .Y(ori_ori_n907_));
  NA2        o0858(.A(ori_ori_n907_), .B(ori_ori_n381_), .Y(ori_ori_n908_));
  AOI210     o0859(.A0(ori_ori_n908_), .A1(ori_ori_n906_), .B0(x3), .Y(ori_ori_n909_));
  NA2        o0860(.A(ori_ori_n634_), .B(ori_ori_n226_), .Y(ori_ori_n910_));
  NO2        o0861(.A(x5), .B(ori_ori_n106_), .Y(ori_ori_n911_));
  NA2        o0862(.A(ori_ori_n216_), .B(ori_ori_n851_), .Y(ori_ori_n912_));
  NA3        o0863(.A(ori_ori_n417_), .B(ori_ori_n124_), .C(ori_ori_n381_), .Y(ori_ori_n913_));
  OAI210     o0864(.A0(ori_ori_n402_), .A1(ori_ori_n195_), .B0(ori_ori_n913_), .Y(ori_ori_n914_));
  AOI210     o0865(.A0(ori_ori_n912_), .A1(ori_ori_n231_), .B0(ori_ori_n914_), .Y(ori_ori_n915_));
  OAI220     o0866(.A0(ori_ori_n915_), .A1(ori_ori_n59_), .B0(ori_ori_n910_), .B1(ori_ori_n644_), .Y(ori_ori_n916_));
  OAI210     o0867(.A0(ori_ori_n916_), .A1(ori_ori_n909_), .B0(ori_ori_n858_), .Y(ori_ori_n917_));
  NO2        o0868(.A(x4), .B(x3), .Y(ori_ori_n918_));
  NO3        o0869(.A(ori_ori_n918_), .B(ori_ori_n313_), .C(ori_ori_n87_), .Y(ori_ori_n919_));
  OAI210     o0870(.A0(ori_ori_n919_), .A1(ori_ori_n250_), .B0(ori_ori_n392_), .Y(ori_ori_n920_));
  AOI210     o0871(.A0(ori_ori_n354_), .A1(ori_ori_n123_), .B0(ori_ori_n227_), .Y(ori_ori_n921_));
  NA2        o0872(.A(ori_ori_n879_), .B(ori_ori_n55_), .Y(ori_ori_n922_));
  NO2        o0873(.A(ori_ori_n922_), .B(ori_ori_n893_), .Y(ori_ori_n923_));
  INV        o0874(.A(ori_ori_n475_), .Y(ori_ori_n924_));
  NO3        o0875(.A(x4), .B(ori_ori_n106_), .C(ori_ori_n59_), .Y(ori_ori_n925_));
  NO2        o0876(.A(ori_ori_n393_), .B(x1), .Y(ori_ori_n926_));
  NOi31      o0877(.An(ori_ori_n925_), .B(ori_ori_n926_), .C(ori_ori_n924_), .Y(ori_ori_n927_));
  NA2        o0878(.A(ori_ori_n55_), .B(x5), .Y(ori_ori_n928_));
  NO4        o0879(.A(ori_ori_n880_), .B(ori_ori_n464_), .C(ori_ori_n928_), .D(x2), .Y(ori_ori_n929_));
  NO4        o0880(.A(ori_ori_n929_), .B(ori_ori_n927_), .C(ori_ori_n923_), .D(ori_ori_n921_), .Y(ori_ori_n930_));
  AOI210     o0881(.A0(ori_ori_n930_), .A1(ori_ori_n920_), .B0(ori_ori_n190_), .Y(ori_ori_n931_));
  NO2        o0882(.A(ori_ori_n603_), .B(ori_ori_n450_), .Y(ori_ori_n932_));
  NO2        o0883(.A(x6), .B(x2), .Y(ori_ori_n933_));
  NO3        o0884(.A(ori_ori_n933_), .B(ori_ori_n634_), .C(ori_ori_n60_), .Y(ori_ori_n934_));
  NA2        o0885(.A(ori_ori_n934_), .B(ori_ori_n244_), .Y(ori_ori_n935_));
  NO2        o0886(.A(ori_ori_n791_), .B(ori_ori_n400_), .Y(ori_ori_n936_));
  NA3        o0887(.A(x4), .B(x3), .C(ori_ori_n106_), .Y(ori_ori_n937_));
  NO3        o0888(.A(ori_ori_n937_), .B(ori_ori_n637_), .C(ori_ori_n417_), .Y(ori_ori_n938_));
  AOI210     o0889(.A0(ori_ori_n936_), .A1(ori_ori_n424_), .B0(ori_ori_n938_), .Y(ori_ori_n939_));
  AOI210     o0890(.A0(ori_ori_n939_), .A1(ori_ori_n935_), .B0(ori_ori_n412_), .Y(ori_ori_n940_));
  NO2        o0891(.A(ori_ori_n55_), .B(ori_ori_n56_), .Y(ori_ori_n941_));
  NO2        o0892(.A(ori_ori_n744_), .B(ori_ori_n414_), .Y(ori_ori_n942_));
  NOi21      o0893(.An(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n943_));
  NO3        o0894(.A(ori_ori_n314_), .B(ori_ori_n295_), .C(ori_ori_n943_), .Y(ori_ori_n944_));
  AOI220     o0895(.A0(ori_ori_n944_), .A1(ori_ori_n230_), .B0(ori_ori_n942_), .B1(ori_ori_n112_), .Y(ori_ori_n945_));
  NO2        o0896(.A(ori_ori_n945_), .B(ori_ori_n941_), .Y(ori_ori_n946_));
  NA2        o0897(.A(ori_ori_n468_), .B(ori_ori_n235_), .Y(ori_ori_n947_));
  NO2        o0898(.A(ori_ori_n435_), .B(ori_ori_n532_), .Y(ori_ori_n948_));
  NA3        o0899(.A(ori_ori_n948_), .B(ori_ori_n947_), .C(ori_ori_n55_), .Y(ori_ori_n949_));
  NO2        o0900(.A(ori_ori_n168_), .B(ori_ori_n106_), .Y(ori_ori_n950_));
  INV        o0901(.A(ori_ori_n949_), .Y(ori_ori_n951_));
  NO4        o0902(.A(ori_ori_n951_), .B(ori_ori_n946_), .C(ori_ori_n940_), .D(ori_ori_n931_), .Y(ori_ori_n952_));
  NA3        o0903(.A(ori_ori_n952_), .B(ori_ori_n917_), .C(ori_ori_n902_), .Y(ori11));
  NA2        o0904(.A(ori_ori_n337_), .B(ori_ori_n90_), .Y(ori_ori_n954_));
  INV        o0905(.A(ori_ori_n810_), .Y(ori_ori_n955_));
  NO2        o0906(.A(ori_ori_n954_), .B(ori_ori_n332_), .Y(ori_ori_n956_));
  NO2        o0907(.A(ori_ori_n693_), .B(x5), .Y(ori_ori_n957_));
  NO2        o0908(.A(ori_ori_n155_), .B(ori_ori_n481_), .Y(ori_ori_n958_));
  AOI220     o0909(.A0(ori_ori_n958_), .A1(ori_ori_n957_), .B0(ori_ori_n956_), .B1(x5), .Y(ori_ori_n959_));
  OAI210     o0910(.A0(ori_ori_n887_), .A1(ori_ori_n198_), .B0(ori_ori_n196_), .Y(ori_ori_n960_));
  NO2        o0911(.A(ori_ori_n311_), .B(ori_ori_n382_), .Y(ori_ori_n961_));
  AOI220     o0912(.A0(ori_ori_n961_), .A1(ori_ori_n166_), .B0(ori_ori_n960_), .B1(ori_ori_n152_), .Y(ori_ori_n962_));
  NO2        o0913(.A(ori_ori_n962_), .B(ori_ori_n402_), .Y(ori_ori_n963_));
  NO2        o0914(.A(ori_ori_n55_), .B(ori_ori_n104_), .Y(ori_ori_n964_));
  NO2        o0915(.A(ori_ori_n71_), .B(x1), .Y(ori_ori_n965_));
  NA2        o0916(.A(ori_ori_n965_), .B(ori_ori_n78_), .Y(ori_ori_n966_));
  NO2        o0917(.A(ori_ori_n277_), .B(ori_ori_n53_), .Y(ori_ori_n967_));
  NO2        o0918(.A(ori_ori_n392_), .B(x3), .Y(ori_ori_n968_));
  NA3        o0919(.A(ori_ori_n968_), .B(ori_ori_n967_), .C(ori_ori_n809_), .Y(ori_ori_n969_));
  AOI210     o0920(.A0(ori_ori_n969_), .A1(ori_ori_n855_), .B0(ori_ori_n353_), .Y(ori_ori_n970_));
  NA2        o0921(.A(ori_ori_n106_), .B(x1), .Y(ori_ori_n971_));
  NO2        o0922(.A(ori_ori_n563_), .B(ori_ori_n200_), .Y(ori_ori_n972_));
  NA4        o0923(.A(ori_ori_n972_), .B(ori_ori_n801_), .C(ori_ori_n421_), .D(ori_ori_n971_), .Y(ori_ori_n973_));
  NA3        o0924(.A(x6), .B(x5), .C(ori_ori_n106_), .Y(ori_ori_n974_));
  NO2        o0925(.A(ori_ori_n974_), .B(ori_ori_n249_), .Y(ori_ori_n975_));
  NO2        o0926(.A(ori_ori_n402_), .B(x0), .Y(ori_ori_n976_));
  NOi31      o0927(.An(ori_ori_n976_), .B(ori_ori_n159_), .C(ori_ori_n51_), .Y(ori_ori_n977_));
  AOI210     o0928(.A0(ori_ori_n975_), .A1(ori_ori_n164_), .B0(ori_ori_n977_), .Y(ori_ori_n978_));
  NA2        o0929(.A(ori_ori_n978_), .B(ori_ori_n973_), .Y(ori_ori_n979_));
  NO3        o0930(.A(ori_ori_n979_), .B(ori_ori_n970_), .C(ori_ori_n963_), .Y(ori_ori_n980_));
  OAI210     o0931(.A0(ori_ori_n959_), .A1(ori_ori_n133_), .B0(ori_ori_n980_), .Y(ori_ori_n981_));
  NA2        o0932(.A(ori_ori_n782_), .B(ori_ori_n87_), .Y(ori_ori_n982_));
  NO3        o0933(.A(ori_ori_n418_), .B(ori_ori_n699_), .C(ori_ori_n119_), .Y(ori_ori_n983_));
  AOI210     o0934(.A0(ori_ori_n982_), .A1(ori_ori_n97_), .B0(ori_ori_n983_), .Y(ori_ori_n984_));
  NO2        o0935(.A(x8), .B(x1), .Y(ori_ori_n985_));
  NO3        o0936(.A(ori_ori_n985_), .B(ori_ori_n626_), .C(ori_ori_n404_), .Y(ori_ori_n986_));
  OAI210     o0937(.A0(ori_ori_n77_), .A1(ori_ori_n53_), .B0(ori_ori_n986_), .Y(ori_ori_n987_));
  OAI210     o0938(.A0(ori_ori_n984_), .A1(x3), .B0(ori_ori_n987_), .Y(ori_ori_n988_));
  NO2        o0939(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n989_));
  OAI210     o0940(.A0(ori_ori_n989_), .A1(x2), .B0(ori_ori_n213_), .Y(ori_ori_n990_));
  NO2        o0941(.A(ori_ori_n468_), .B(x4), .Y(ori_ori_n991_));
  NO3        o0942(.A(ori_ori_n55_), .B(x6), .C(x1), .Y(ori_ori_n992_));
  NOi21      o0943(.An(ori_ori_n992_), .B(ori_ori_n435_), .Y(ori_ori_n993_));
  AOI210     o0944(.A0(ori_ori_n991_), .A1(ori_ori_n522_), .B0(ori_ori_n993_), .Y(ori_ori_n994_));
  INV        o0945(.A(ori_ori_n994_), .Y(ori_ori_n995_));
  AOI210     o0946(.A0(ori_ori_n988_), .A1(x2), .B0(ori_ori_n995_), .Y(ori_ori_n996_));
  NO2        o0947(.A(ori_ori_n212_), .B(x2), .Y(ori_ori_n997_));
  NA2        o0948(.A(ori_ori_n997_), .B(ori_ori_n918_), .Y(ori_ori_n998_));
  NOi21      o0949(.An(ori_ori_n346_), .B(ori_ori_n514_), .Y(ori_ori_n999_));
  NO3        o0950(.A(ori_ori_n999_), .B(ori_ori_n550_), .C(ori_ori_n295_), .Y(ori_ori_n1000_));
  NA2        o0951(.A(x8), .B(ori_ori_n106_), .Y(ori_ori_n1001_));
  OAI220     o0952(.A0(ori_ori_n644_), .A1(ori_ori_n1001_), .B0(ori_ori_n295_), .B1(ori_ori_n341_), .Y(ori_ori_n1002_));
  OAI210     o0953(.A0(ori_ori_n1002_), .A1(ori_ori_n1000_), .B0(ori_ori_n71_), .Y(ori_ori_n1003_));
  NO2        o0954(.A(ori_ori_n104_), .B(x1), .Y(ori_ori_n1004_));
  NA2        o0955(.A(ori_ori_n1004_), .B(x7), .Y(ori_ori_n1005_));
  AOI210     o0956(.A0(ori_ori_n1003_), .A1(ori_ori_n998_), .B0(ori_ori_n1005_), .Y(ori_ori_n1006_));
  NA2        o0957(.A(ori_ori_n84_), .B(ori_ori_n71_), .Y(ori_ori_n1007_));
  INV        o0958(.A(ori_ori_n225_), .Y(ori_ori_n1008_));
  INV        o0959(.A(ori_ori_n1006_), .Y(ori_ori_n1009_));
  OAI210     o0960(.A0(ori_ori_n996_), .A1(ori_ori_n769_), .B0(ori_ori_n1009_), .Y(ori_ori_n1010_));
  AO210      o0961(.A0(ori_ori_n981_), .A1(ori_ori_n57_), .B0(ori_ori_n1010_), .Y(ori12));
  NA2        o0962(.A(ori_ori_n800_), .B(ori_ori_n224_), .Y(ori_ori_n1012_));
  NO2        o0963(.A(ori_ori_n567_), .B(x7), .Y(ori_ori_n1013_));
  NA2        o0964(.A(ori_ori_n636_), .B(ori_ori_n791_), .Y(ori_ori_n1014_));
  NO2        o0965(.A(ori_ori_n1012_), .B(ori_ori_n1014_), .Y(ori_ori_n1015_));
  NOi21      o0966(.An(ori_ori_n359_), .B(ori_ori_n501_), .Y(ori_ori_n1016_));
  NO2        o0967(.A(x7), .B(ori_ori_n50_), .Y(ori_ori_n1017_));
  NO2        o0968(.A(ori_ori_n551_), .B(ori_ori_n1017_), .Y(ori_ori_n1018_));
  NO3        o0969(.A(ori_ori_n784_), .B(ori_ori_n108_), .C(ori_ori_n95_), .Y(ori_ori_n1019_));
  AOI210     o0970(.A0(ori_ori_n1018_), .A1(ori_ori_n926_), .B0(ori_ori_n1019_), .Y(ori_ori_n1020_));
  NA2        o0971(.A(ori_ori_n964_), .B(ori_ori_n56_), .Y(ori_ori_n1021_));
  OAI220     o0972(.A0(ori_ori_n1021_), .A1(ori_ori_n523_), .B0(ori_ori_n1020_), .B1(ori_ori_n1016_), .Y(ori_ori_n1022_));
  OAI210     o0973(.A0(ori_ori_n1022_), .A1(ori_ori_n1015_), .B0(ori_ori_n527_), .Y(ori_ori_n1023_));
  NA2        o0974(.A(ori_ori_n87_), .B(x5), .Y(ori_ori_n1024_));
  OAI210     o0975(.A0(ori_ori_n1024_), .A1(ori_ori_n295_), .B0(ori_ori_n655_), .Y(ori_ori_n1025_));
  INV        o0976(.A(ori_ori_n1025_), .Y(ori_ori_n1026_));
  NA2        o0977(.A(ori_ori_n549_), .B(ori_ori_n53_), .Y(ori_ori_n1027_));
  NA2        o0978(.A(ori_ori_n260_), .B(ori_ori_n50_), .Y(ori_ori_n1028_));
  OAI220     o0979(.A0(ori_ori_n1028_), .A1(ori_ori_n283_), .B0(ori_ori_n1027_), .B1(ori_ori_n129_), .Y(ori_ori_n1029_));
  NO2        o0980(.A(ori_ori_n982_), .B(ori_ori_n463_), .Y(ori_ori_n1030_));
  NO3        o0981(.A(ori_ori_n218_), .B(ori_ori_n60_), .C(ori_ori_n57_), .Y(ori_ori_n1031_));
  AOI220     o0982(.A0(ori_ori_n1031_), .A1(ori_ori_n1030_), .B0(ori_ori_n1029_), .B1(ori_ori_n56_), .Y(ori_ori_n1032_));
  OAI210     o0983(.A0(ori_ori_n1026_), .A1(ori_ori_n64_), .B0(ori_ori_n1032_), .Y(ori_ori_n1033_));
  NO2        o0984(.A(ori_ori_n57_), .B(x0), .Y(ori_ori_n1034_));
  NO2        o0985(.A(ori_ori_n603_), .B(ori_ori_n292_), .Y(ori_ori_n1035_));
  NO2        o0986(.A(ori_ori_n680_), .B(x3), .Y(ori_ori_n1036_));
  NO2        o0987(.A(ori_ori_n601_), .B(x8), .Y(ori_ori_n1037_));
  NO2        o0988(.A(ori_ori_n626_), .B(x7), .Y(ori_ori_n1038_));
  NO3        o0989(.A(ori_ori_n1038_), .B(ori_ori_n552_), .C(x8), .Y(ori_ori_n1039_));
  NA4        o0990(.A(ori_ori_n605_), .B(ori_ori_n597_), .C(ori_ori_n188_), .D(x0), .Y(ori_ori_n1040_));
  NO2        o0991(.A(ori_ori_n1040_), .B(ori_ori_n1039_), .Y(ori_ori_n1041_));
  AOI210     o0992(.A0(ori_ori_n1033_), .A1(ori_ori_n933_), .B0(ori_ori_n1041_), .Y(ori_ori_n1042_));
  NO2        o0993(.A(ori_ori_n230_), .B(x8), .Y(ori_ori_n1043_));
  NO2        o0994(.A(ori_ori_n858_), .B(ori_ori_n96_), .Y(ori_ori_n1044_));
  NO2        o0995(.A(ori_ori_n154_), .B(ori_ori_n53_), .Y(ori_ori_n1045_));
  AOI210     o0996(.A0(ori_ori_n311_), .A1(x8), .B0(ori_ori_n1045_), .Y(ori_ori_n1046_));
  AOI210     o0997(.A0(ori_ori_n198_), .A1(ori_ori_n92_), .B0(ori_ori_n1046_), .Y(ori_ori_n1047_));
  OAI210     o0998(.A0(ori_ori_n1047_), .A1(ori_ori_n1044_), .B0(ori_ori_n614_), .Y(ori_ori_n1048_));
  NO2        o0999(.A(x7), .B(x0), .Y(ori_ori_n1049_));
  NO3        o1000(.A(ori_ori_n146_), .B(ori_ori_n1049_), .C(ori_ori_n135_), .Y(ori_ori_n1050_));
  XN2        o1001(.A(x8), .B(x7), .Y(ori_ori_n1051_));
  NO3        o1002(.A(ori_ori_n985_), .B(ori_ori_n233_), .C(ori_ori_n1051_), .Y(ori_ori_n1052_));
  OAI210     o1003(.A0(ori_ori_n1052_), .A1(ori_ori_n1050_), .B0(ori_ori_n665_), .Y(ori_ori_n1053_));
  NO2        o1004(.A(ori_ori_n242_), .B(ori_ori_n238_), .Y(ori_ori_n1054_));
  NO2        o1005(.A(ori_ori_n104_), .B(x4), .Y(ori_ori_n1055_));
  OAI210     o1006(.A0(ori_ori_n1054_), .A1(ori_ori_n250_), .B0(ori_ori_n1055_), .Y(ori_ori_n1056_));
  NA3        o1007(.A(ori_ori_n1056_), .B(ori_ori_n1053_), .C(ori_ori_n1048_), .Y(ori_ori_n1057_));
  NA2        o1008(.A(ori_ori_n1057_), .B(ori_ori_n505_), .Y(ori_ori_n1058_));
  NO2        o1009(.A(ori_ori_n55_), .B(x4), .Y(ori_ori_n1059_));
  NA2        o1010(.A(ori_ori_n1059_), .B(ori_ori_n151_), .Y(ori_ori_n1060_));
  NO2        o1011(.A(ori_ori_n607_), .B(ori_ori_n233_), .Y(ori_ori_n1061_));
  NA2        o1012(.A(ori_ori_n1061_), .B(ori_ori_n50_), .Y(ori_ori_n1062_));
  AOI210     o1013(.A0(ori_ori_n1062_), .A1(ori_ori_n1060_), .B0(ori_ori_n387_), .Y(ori_ori_n1063_));
  NA3        o1014(.A(ori_ori_n2466_), .B(ori_ori_n614_), .C(x1), .Y(ori_ori_n1064_));
  OAI210     o1015(.A0(x8), .A1(x0), .B0(x4), .Y(ori_ori_n1065_));
  NO2        o1016(.A(x7), .B(ori_ori_n56_), .Y(ori_ori_n1066_));
  NO2        o1017(.A(ori_ori_n68_), .B(ori_ori_n1066_), .Y(ori_ori_n1067_));
  NOi21      o1018(.An(ori_ori_n1065_), .B(ori_ori_n1067_), .Y(ori_ori_n1068_));
  NO2        o1019(.A(ori_ori_n605_), .B(ori_ori_n295_), .Y(ori_ori_n1069_));
  NO2        o1020(.A(ori_ori_n701_), .B(ori_ori_n201_), .Y(ori_ori_n1070_));
  OAI210     o1021(.A0(ori_ori_n1069_), .A1(ori_ori_n1068_), .B0(ori_ori_n1070_), .Y(ori_ori_n1071_));
  NO2        o1022(.A(ori_ori_n133_), .B(ori_ori_n132_), .Y(ori_ori_n1072_));
  NO2        o1023(.A(ori_ori_n551_), .B(ori_ori_n400_), .Y(ori_ori_n1073_));
  OAI210     o1024(.A0(ori_ori_n1073_), .A1(ori_ori_n1072_), .B0(ori_ori_n230_), .Y(ori_ori_n1074_));
  NO2        o1025(.A(ori_ori_n742_), .B(ori_ori_n378_), .Y(ori_ori_n1075_));
  NA2        o1026(.A(ori_ori_n299_), .B(ori_ori_n59_), .Y(ori_ori_n1076_));
  NO2        o1027(.A(ori_ori_n1021_), .B(ori_ori_n1076_), .Y(ori_ori_n1077_));
  AOI210     o1028(.A0(ori_ori_n1075_), .A1(ori_ori_n164_), .B0(ori_ori_n1077_), .Y(ori_ori_n1078_));
  NA4        o1029(.A(ori_ori_n1078_), .B(ori_ori_n1074_), .C(ori_ori_n1071_), .D(ori_ori_n1064_), .Y(ori_ori_n1079_));
  OAI210     o1030(.A0(ori_ori_n1079_), .A1(ori_ori_n1063_), .B0(ori_ori_n616_), .Y(ori_ori_n1080_));
  NA4        o1031(.A(ori_ori_n1080_), .B(ori_ori_n1058_), .C(ori_ori_n1042_), .D(ori_ori_n1023_), .Y(ori13));
  NO2        o1032(.A(ori_ori_n417_), .B(ori_ori_n318_), .Y(ori_ori_n1082_));
  NOi41      o1033(.An(ori_ori_n1082_), .B(ori_ori_n614_), .C(ori_ori_n264_), .D(ori_ori_n218_), .Y(ori_ori_n1083_));
  NO2        o1034(.A(ori_ori_n784_), .B(ori_ori_n168_), .Y(ori_ori_n1084_));
  NO2        o1035(.A(ori_ori_n145_), .B(ori_ori_n71_), .Y(ori_ori_n1085_));
  XN2        o1036(.A(x4), .B(x0), .Y(ori_ori_n1086_));
  NO3        o1037(.A(ori_ori_n1086_), .B(ori_ori_n107_), .C(ori_ori_n378_), .Y(ori_ori_n1087_));
  AO220      o1038(.A0(ori_ori_n1087_), .A1(ori_ori_n1085_), .B0(ori_ori_n1084_), .B1(ori_ori_n300_), .Y(ori_ori_n1088_));
  OAI210     o1039(.A0(ori_ori_n1088_), .A1(ori_ori_n1083_), .B0(x3), .Y(ori_ori_n1089_));
  NO2        o1040(.A(ori_ori_n784_), .B(x6), .Y(ori_ori_n1090_));
  NO2        o1041(.A(ori_ori_n1028_), .B(ori_ori_n351_), .Y(ori_ori_n1091_));
  NO3        o1042(.A(x8), .B(x5), .C(ori_ori_n106_), .Y(ori_ori_n1092_));
  NO2        o1043(.A(ori_ori_n551_), .B(ori_ori_n183_), .Y(ori_ori_n1093_));
  NA2        o1044(.A(ori_ori_n1093_), .B(ori_ori_n992_), .Y(ori_ori_n1094_));
  NA2        o1045(.A(ori_ori_n404_), .B(ori_ori_n53_), .Y(ori_ori_n1095_));
  NO2        o1046(.A(ori_ori_n1095_), .B(ori_ori_n851_), .Y(ori_ori_n1096_));
  INV        o1047(.A(ori_ori_n422_), .Y(ori_ori_n1097_));
  NA2        o1048(.A(ori_ori_n56_), .B(ori_ori_n106_), .Y(ori_ori_n1098_));
  NA2        o1049(.A(ori_ori_n1098_), .B(x1), .Y(ori_ori_n1099_));
  NO2        o1050(.A(ori_ori_n1099_), .B(ori_ori_n235_), .Y(ori_ori_n1100_));
  NO2        o1051(.A(ori_ori_n292_), .B(x6), .Y(ori_ori_n1101_));
  INV        o1052(.A(ori_ori_n869_), .Y(ori_ori_n1102_));
  AOI220     o1053(.A0(ori_ori_n1102_), .A1(ori_ori_n1101_), .B0(ori_ori_n1100_), .B1(ori_ori_n1097_), .Y(ori_ori_n1103_));
  NAi31      o1054(.An(ori_ori_n1096_), .B(ori_ori_n1103_), .C(ori_ori_n1094_), .Y(ori_ori_n1104_));
  AOI220     o1055(.A0(ori_ori_n1104_), .A1(ori_ori_n68_), .B0(ori_ori_n1091_), .B1(ori_ori_n1090_), .Y(ori_ori_n1105_));
  NA2        o1056(.A(ori_ori_n71_), .B(x3), .Y(ori_ori_n1106_));
  NA2        o1057(.A(ori_ori_n1106_), .B(ori_ori_n818_), .Y(ori_ori_n1107_));
  OAI220     o1058(.A0(ori_ori_n276_), .A1(ori_ori_n742_), .B0(ori_ori_n87_), .B1(ori_ori_n77_), .Y(ori_ori_n1108_));
  AOI210     o1059(.A0(ori_ori_n1024_), .A1(ori_ori_n561_), .B0(ori_ori_n891_), .Y(ori_ori_n1109_));
  OA210      o1060(.A0(ori_ori_n1108_), .A1(ori_ori_n1107_), .B0(ori_ori_n1109_), .Y(ori_ori_n1110_));
  NA2        o1061(.A(ori_ori_n563_), .B(ori_ori_n55_), .Y(ori_ori_n1111_));
  NA2        o1062(.A(ori_ori_n456_), .B(ori_ori_n444_), .Y(ori_ori_n1112_));
  NA2        o1063(.A(x6), .B(ori_ori_n50_), .Y(ori_ori_n1113_));
  NA2        o1064(.A(ori_ori_n1113_), .B(ori_ori_n490_), .Y(ori_ori_n1114_));
  NO2        o1065(.A(ori_ori_n148_), .B(ori_ori_n124_), .Y(ori_ori_n1115_));
  AOI210     o1066(.A0(ori_ori_n1114_), .A1(ori_ori_n388_), .B0(ori_ori_n1115_), .Y(ori_ori_n1116_));
  OAI220     o1067(.A0(ori_ori_n1116_), .A1(ori_ori_n791_), .B0(ori_ori_n1112_), .B1(ori_ori_n1111_), .Y(ori_ori_n1117_));
  OAI210     o1068(.A0(ori_ori_n1117_), .A1(ori_ori_n1110_), .B0(ori_ori_n1049_), .Y(ori_ori_n1118_));
  NAi21      o1069(.An(ori_ori_n84_), .B(ori_ori_n341_), .Y(ori_ori_n1119_));
  NO2        o1070(.A(ori_ori_n1119_), .B(ori_ori_n71_), .Y(ori_ori_n1120_));
  AOI210     o1071(.A0(ori_ori_n151_), .A1(x4), .B0(ori_ori_n160_), .Y(ori_ori_n1121_));
  NO2        o1072(.A(ori_ori_n1121_), .B(x0), .Y(ori_ori_n1122_));
  NO2        o1073(.A(ori_ori_n157_), .B(ori_ori_n267_), .Y(ori_ori_n1123_));
  OAI210     o1074(.A0(ori_ori_n1123_), .A1(ori_ori_n1122_), .B0(ori_ori_n1120_), .Y(ori_ori_n1124_));
  NA3        o1075(.A(ori_ori_n1055_), .B(ori_ori_n174_), .C(ori_ori_n71_), .Y(ori_ori_n1125_));
  NO2        o1076(.A(x4), .B(x0), .Y(ori_ori_n1126_));
  NA2        o1077(.A(ori_ori_n1125_), .B(ori_ori_n1124_), .Y(ori_ori_n1127_));
  NA2        o1078(.A(ori_ori_n226_), .B(ori_ori_n665_), .Y(ori_ori_n1128_));
  NA2        o1079(.A(ori_ori_n56_), .B(x0), .Y(ori_ori_n1129_));
  NO2        o1080(.A(ori_ori_n295_), .B(ori_ori_n341_), .Y(ori_ori_n1130_));
  NO2        o1081(.A(ori_ori_n626_), .B(x0), .Y(ori_ori_n1131_));
  OAI210     o1082(.A0(ori_ori_n1131_), .A1(ori_ori_n1130_), .B0(ori_ori_n303_), .Y(ori_ori_n1132_));
  NO2        o1083(.A(ori_ori_n712_), .B(x1), .Y(ori_ori_n1133_));
  AOI220     o1084(.A0(ori_ori_n1133_), .A1(ori_ori_n557_), .B0(ori_ori_n432_), .B1(ori_ori_n268_), .Y(ori_ori_n1134_));
  NA2        o1085(.A(ori_ori_n450_), .B(ori_ori_n50_), .Y(ori_ori_n1135_));
  AOI220     o1086(.A0(ori_ori_n1135_), .A1(ori_ori_n1084_), .B0(ori_ori_n892_), .B1(ori_ori_n97_), .Y(ori_ori_n1136_));
  NA3        o1087(.A(ori_ori_n1136_), .B(ori_ori_n1134_), .C(ori_ori_n1132_), .Y(ori_ori_n1137_));
  AOI220     o1088(.A0(ori_ori_n1137_), .A1(ori_ori_n125_), .B0(ori_ori_n1127_), .B1(ori_ori_n67_), .Y(ori_ori_n1138_));
  NA4        o1089(.A(ori_ori_n1138_), .B(ori_ori_n1118_), .C(ori_ori_n1105_), .D(ori_ori_n1089_), .Y(ori14));
  NO2        o1090(.A(ori_ori_n335_), .B(ori_ori_n71_), .Y(ori_ori_n1140_));
  NO3        o1091(.A(x7), .B(x6), .C(x0), .Y(ori_ori_n1141_));
  OAI210     o1092(.A0(ori_ori_n1141_), .A1(ori_ori_n1140_), .B0(x8), .Y(ori_ori_n1142_));
  NA2        o1093(.A(ori_ori_n1037_), .B(ori_ori_n85_), .Y(ori_ori_n1143_));
  AOI210     o1094(.A0(ori_ori_n1143_), .A1(ori_ori_n1142_), .B0(ori_ori_n144_), .Y(ori_ori_n1144_));
  AOI220     o1095(.A0(ori_ori_n336_), .A1(ori_ori_n769_), .B0(ori_ori_n404_), .B1(ori_ori_n378_), .Y(ori_ori_n1145_));
  NA2        o1096(.A(ori_ori_n251_), .B(ori_ori_n887_), .Y(ori_ori_n1146_));
  OAI220     o1097(.A0(ori_ori_n1146_), .A1(ori_ori_n1145_), .B0(ori_ori_n420_), .B1(ori_ori_n726_), .Y(ori_ori_n1147_));
  OA210      o1098(.A0(ori_ori_n1147_), .A1(ori_ori_n1144_), .B0(x4), .Y(ori_ori_n1148_));
  NO2        o1099(.A(ori_ori_n132_), .B(ori_ori_n555_), .Y(ori_ori_n1149_));
  NA2        o1100(.A(x6), .B(x2), .Y(ori_ori_n1150_));
  NO3        o1101(.A(ori_ori_n551_), .B(ori_ori_n337_), .C(ori_ori_n272_), .Y(ori_ori_n1151_));
  NA2        o1102(.A(ori_ori_n1151_), .B(ori_ori_n59_), .Y(ori_ori_n1152_));
  NA2        o1103(.A(x6), .B(ori_ori_n104_), .Y(ori_ori_n1153_));
  NO2        o1104(.A(ori_ori_n603_), .B(ori_ori_n1153_), .Y(ori_ori_n1154_));
  AOI210     o1105(.A0(ori_ori_n1037_), .A1(ori_ori_n925_), .B0(x1), .Y(ori_ori_n1155_));
  NO2        o1106(.A(ori_ori_n485_), .B(x5), .Y(ori_ori_n1156_));
  NA3        o1107(.A(ori_ori_n1156_), .B(ori_ori_n118_), .C(x0), .Y(ori_ori_n1157_));
  NA3        o1108(.A(ori_ori_n633_), .B(ori_ori_n841_), .C(ori_ori_n68_), .Y(ori_ori_n1158_));
  AN3        o1109(.A(ori_ori_n1158_), .B(ori_ori_n1157_), .C(ori_ori_n1155_), .Y(ori_ori_n1159_));
  NO2        o1110(.A(ori_ori_n637_), .B(ori_ori_n1001_), .Y(ori_ori_n1160_));
  NO2        o1111(.A(ori_ori_n77_), .B(ori_ori_n58_), .Y(ori_ori_n1161_));
  OAI210     o1112(.A0(ori_ori_n1160_), .A1(ori_ori_n401_), .B0(ori_ori_n1161_), .Y(ori_ori_n1162_));
  AO210      o1113(.A0(ori_ori_n1140_), .A1(ori_ori_n925_), .B0(ori_ori_n53_), .Y(ori_ori_n1163_));
  AOI210     o1114(.A0(ori_ori_n692_), .A1(ori_ori_n736_), .B0(ori_ori_n1163_), .Y(ori_ori_n1164_));
  AOI220     o1115(.A0(ori_ori_n1164_), .A1(ori_ori_n1162_), .B0(ori_ori_n1159_), .B1(ori_ori_n1152_), .Y(ori_ori_n1165_));
  NO2        o1116(.A(ori_ori_n1165_), .B(ori_ori_n1148_), .Y(ori_ori_n1166_));
  NO2        o1117(.A(ori_ori_n292_), .B(x2), .Y(ori_ori_n1167_));
  XN2        o1118(.A(x4), .B(x1), .Y(ori_ori_n1168_));
  NO2        o1119(.A(ori_ori_n1168_), .B(ori_ori_n276_), .Y(ori_ori_n1169_));
  NOi21      o1120(.An(ori_ori_n1169_), .B(ori_ori_n366_), .Y(ori_ori_n1170_));
  NO2        o1121(.A(ori_ori_n310_), .B(ori_ori_n60_), .Y(ori_ori_n1171_));
  OAI210     o1122(.A0(ori_ori_n1171_), .A1(ori_ori_n1170_), .B0(ori_ori_n1167_), .Y(ori_ori_n1172_));
  NA2        o1123(.A(ori_ori_n627_), .B(ori_ori_n56_), .Y(ori_ori_n1173_));
  OAI220     o1124(.A0(ori_ori_n1173_), .A1(ori_ori_n145_), .B0(ori_ori_n175_), .B1(ori_ori_n71_), .Y(ori_ori_n1174_));
  NO2        o1125(.A(ori_ori_n198_), .B(ori_ori_n233_), .Y(ori_ori_n1175_));
  NA2        o1126(.A(ori_ori_n226_), .B(ori_ori_n322_), .Y(ori_ori_n1176_));
  NA2        o1127(.A(ori_ori_n581_), .B(ori_ori_n943_), .Y(ori_ori_n1177_));
  NO2        o1128(.A(ori_ori_n1177_), .B(ori_ori_n1176_), .Y(ori_ori_n1178_));
  AOI210     o1129(.A0(ori_ori_n1175_), .A1(ori_ori_n1174_), .B0(ori_ori_n1178_), .Y(ori_ori_n1179_));
  AOI210     o1130(.A0(ori_ori_n1179_), .A1(ori_ori_n1172_), .B0(x7), .Y(ori_ori_n1180_));
  NO2        o1131(.A(ori_ori_n443_), .B(x6), .Y(ori_ori_n1181_));
  NO2        o1132(.A(ori_ori_n738_), .B(ori_ori_n1181_), .Y(ori_ori_n1182_));
  OAI220     o1133(.A0(ori_ori_n1182_), .A1(ori_ori_n55_), .B0(ori_ori_n443_), .B1(ori_ori_n100_), .Y(ori_ori_n1183_));
  NA2        o1134(.A(ori_ori_n1183_), .B(ori_ori_n324_), .Y(ori_ori_n1184_));
  NA3        o1135(.A(ori_ori_n558_), .B(ori_ori_n971_), .C(ori_ori_n70_), .Y(ori_ori_n1185_));
  NO3        o1136(.A(ori_ori_n966_), .B(ori_ori_n744_), .C(ori_ori_n433_), .Y(ori_ori_n1186_));
  NO2        o1137(.A(ori_ori_n1186_), .B(ori_ori_n948_), .Y(ori_ori_n1187_));
  AOI210     o1138(.A0(ori_ori_n1187_), .A1(ori_ori_n1184_), .B0(ori_ori_n278_), .Y(ori_ori_n1188_));
  NA2        o1139(.A(ori_ori_n816_), .B(ori_ori_n53_), .Y(ori_ori_n1189_));
  OAI210     o1140(.A0(ori_ori_n222_), .A1(ori_ori_n114_), .B0(x2), .Y(ori_ori_n1190_));
  NA2        o1141(.A(ori_ori_n333_), .B(ori_ori_n56_), .Y(ori_ori_n1191_));
  OA220      o1142(.A0(ori_ori_n1191_), .A1(ori_ori_n1190_), .B0(ori_ori_n1189_), .B1(ori_ori_n336_), .Y(ori_ori_n1192_));
  NA2        o1143(.A(ori_ori_n56_), .B(x2), .Y(ori_ori_n1193_));
  NO2        o1144(.A(ori_ori_n1193_), .B(ori_ori_n182_), .Y(ori_ori_n1194_));
  NA4        o1145(.A(ori_ori_n1194_), .B(ori_ori_n333_), .C(ori_ori_n233_), .D(ori_ori_n67_), .Y(ori_ori_n1195_));
  OAI210     o1146(.A0(ori_ori_n1192_), .A1(ori_ori_n288_), .B0(ori_ori_n1195_), .Y(ori_ori_n1196_));
  NO3        o1147(.A(ori_ori_n1196_), .B(ori_ori_n1188_), .C(ori_ori_n1180_), .Y(ori_ori_n1197_));
  OAI210     o1148(.A0(ori_ori_n1166_), .A1(x3), .B0(ori_ori_n1197_), .Y(ori15));
  NA2        o1149(.A(ori_ori_n533_), .B(ori_ori_n59_), .Y(ori_ori_n1199_));
  NAi41      o1150(.An(x2), .B(x7), .C(x6), .D(x0), .Y(ori_ori_n1200_));
  AOI210     o1151(.A0(ori_ori_n1200_), .A1(ori_ori_n1199_), .B0(ori_ori_n53_), .Y(ori_ori_n1201_));
  NA2        o1152(.A(ori_ori_n1201_), .B(ori_ori_n1055_), .Y(ori_ori_n1202_));
  NA2        o1153(.A(ori_ori_n108_), .B(ori_ori_n106_), .Y(ori_ori_n1203_));
  NA4        o1154(.A(ori_ori_n1203_), .B(ori_ori_n580_), .C(ori_ori_n282_), .D(x6), .Y(ori_ori_n1204_));
  AOI210     o1155(.A0(ori_ori_n664_), .A1(ori_ori_n76_), .B0(x3), .Y(ori_ori_n1205_));
  NA3        o1156(.A(ori_ori_n1205_), .B(ori_ori_n1204_), .C(ori_ori_n1202_), .Y(ori_ori_n1206_));
  AOI210     o1157(.A0(ori_ori_n976_), .A1(ori_ori_n537_), .B0(ori_ori_n50_), .Y(ori_ori_n1207_));
  NO2        o1158(.A(ori_ori_n267_), .B(ori_ori_n106_), .Y(ori_ori_n1208_));
  NO2        o1159(.A(ori_ori_n216_), .B(x5), .Y(ori_ori_n1209_));
  NA2        o1160(.A(ori_ori_n1209_), .B(ori_ori_n1208_), .Y(ori_ori_n1210_));
  NA3        o1161(.A(ori_ori_n1133_), .B(ori_ori_n570_), .C(ori_ori_n1066_), .Y(ori_ori_n1211_));
  NA4        o1162(.A(ori_ori_n1211_), .B(ori_ori_n1210_), .C(ori_ori_n1207_), .D(ori_ori_n1157_), .Y(ori_ori_n1212_));
  NA2        o1163(.A(ori_ori_n304_), .B(ori_ori_n312_), .Y(ori_ori_n1213_));
  AOI210     o1164(.A0(ori_ori_n1099_), .A1(ori_ori_n58_), .B0(ori_ori_n1213_), .Y(ori_ori_n1214_));
  NA4        o1165(.A(ori_ori_n1099_), .B(ori_ori_n636_), .C(ori_ori_n1034_), .D(ori_ori_n341_), .Y(ori_ori_n1215_));
  NA2        o1166(.A(ori_ori_n537_), .B(ori_ori_n421_), .Y(ori_ori_n1216_));
  NO2        o1167(.A(ori_ori_n680_), .B(ori_ori_n53_), .Y(ori_ori_n1217_));
  NO2        o1168(.A(ori_ori_n701_), .B(ori_ori_n272_), .Y(ori_ori_n1218_));
  NA2        o1169(.A(ori_ori_n1218_), .B(ori_ori_n1217_), .Y(ori_ori_n1219_));
  NA3        o1170(.A(ori_ori_n1219_), .B(ori_ori_n1216_), .C(ori_ori_n1215_), .Y(ori_ori_n1220_));
  OAI210     o1171(.A0(ori_ori_n1220_), .A1(ori_ori_n1214_), .B0(ori_ori_n77_), .Y(ori_ori_n1221_));
  NA2        o1172(.A(ori_ori_n334_), .B(ori_ori_n639_), .Y(ori_ori_n1222_));
  NA2        o1173(.A(ori_ori_n518_), .B(ori_ori_n56_), .Y(ori_ori_n1223_));
  NA3        o1174(.A(ori_ori_n1223_), .B(ori_ori_n312_), .C(ori_ori_n108_), .Y(ori_ori_n1224_));
  AOI210     o1175(.A0(ori_ori_n1224_), .A1(ori_ori_n1222_), .B0(ori_ori_n450_), .Y(ori_ori_n1225_));
  NO3        o1176(.A(ori_ori_n724_), .B(ori_ori_n568_), .C(ori_ori_n183_), .Y(ori_ori_n1226_));
  OAI210     o1177(.A0(ori_ori_n1226_), .A1(ori_ori_n1225_), .B0(ori_ori_n443_), .Y(ori_ori_n1227_));
  NO2        o1178(.A(ori_ori_n791_), .B(ori_ori_n50_), .Y(ori_ori_n1228_));
  NO2        o1179(.A(ori_ori_n224_), .B(ori_ori_n64_), .Y(ori_ori_n1229_));
  OA210      o1180(.A0(ori_ori_n1229_), .A1(ori_ori_n1228_), .B0(ori_ori_n366_), .Y(ori_ori_n1230_));
  NA2        o1181(.A(ori_ori_n57_), .B(x3), .Y(ori_ori_n1231_));
  AOI210     o1182(.A0(ori_ori_n893_), .A1(ori_ori_n1231_), .B0(ori_ori_n621_), .Y(ori_ori_n1232_));
  OAI210     o1183(.A0(ori_ori_n1232_), .A1(ori_ori_n1230_), .B0(ori_ori_n933_), .Y(ori_ori_n1233_));
  NA2        o1184(.A(ori_ori_n1194_), .B(ori_ori_n68_), .Y(ori_ori_n1234_));
  NO2        o1185(.A(ori_ori_n1150_), .B(x0), .Y(ori_ori_n1235_));
  AOI210     o1186(.A0(ori_ori_n1235_), .A1(ori_ori_n552_), .B0(x8), .Y(ori_ori_n1236_));
  NO2        o1187(.A(ori_ori_n387_), .B(ori_ori_n81_), .Y(ori_ori_n1237_));
  NO2        o1188(.A(ori_ori_n845_), .B(ori_ori_n71_), .Y(ori_ori_n1238_));
  NA2        o1189(.A(ori_ori_n1238_), .B(ori_ori_n1237_), .Y(ori_ori_n1239_));
  NO2        o1190(.A(ori_ori_n891_), .B(x6), .Y(ori_ori_n1240_));
  NA3        o1191(.A(ori_ori_n1240_), .B(ori_ori_n542_), .C(ori_ori_n370_), .Y(ori_ori_n1241_));
  AN4        o1192(.A(ori_ori_n1241_), .B(ori_ori_n1239_), .C(ori_ori_n1236_), .D(ori_ori_n1234_), .Y(ori_ori_n1242_));
  NA4        o1193(.A(ori_ori_n1242_), .B(ori_ori_n1233_), .C(ori_ori_n1227_), .D(ori_ori_n1221_), .Y(ori_ori_n1243_));
  NA2        o1194(.A(ori_ori_n152_), .B(ori_ori_n670_), .Y(ori_ori_n1244_));
  NO2        o1195(.A(ori_ori_n588_), .B(x2), .Y(ori_ori_n1245_));
  OAI210     o1196(.A0(ori_ori_n1245_), .A1(ori_ori_n85_), .B0(x1), .Y(ori_ori_n1246_));
  AOI210     o1197(.A0(ori_ori_n1246_), .A1(ori_ori_n1244_), .B0(ori_ori_n292_), .Y(ori_ori_n1247_));
  NA3        o1198(.A(ori_ori_n57_), .B(x1), .C(x0), .Y(ori_ori_n1248_));
  NA4        o1199(.A(x7), .B(x3), .C(ori_ori_n53_), .D(x0), .Y(ori_ori_n1249_));
  NAi21      o1200(.An(ori_ori_n112_), .B(ori_ori_n674_), .Y(ori_ori_n1250_));
  NA3        o1201(.A(ori_ori_n1250_), .B(ori_ori_n290_), .C(ori_ori_n570_), .Y(ori_ori_n1251_));
  OAI220     o1202(.A0(ori_ori_n295_), .A1(x7), .B0(ori_ori_n124_), .B1(ori_ori_n71_), .Y(ori_ori_n1252_));
  NA2        o1203(.A(ori_ori_n1252_), .B(ori_ori_n1004_), .Y(ori_ori_n1253_));
  NA2        o1204(.A(ori_ori_n82_), .B(ori_ori_n50_), .Y(ori_ori_n1254_));
  AO210      o1205(.A0(ori_ori_n1254_), .A1(ori_ori_n287_), .B0(ori_ori_n144_), .Y(ori_ori_n1255_));
  NA4        o1206(.A(ori_ori_n1255_), .B(ori_ori_n1253_), .C(ori_ori_n1251_), .D(ori_ori_n1249_), .Y(ori_ori_n1256_));
  OAI210     o1207(.A0(ori_ori_n1256_), .A1(ori_ori_n1247_), .B0(ori_ori_n56_), .Y(ori_ori_n1257_));
  AOI210     o1208(.A0(ori_ori_n629_), .A1(x4), .B0(ori_ori_n871_), .Y(ori_ori_n1258_));
  OAI220     o1209(.A0(ori_ori_n1258_), .A1(ori_ori_n273_), .B0(ori_ori_n937_), .B1(ori_ori_n859_), .Y(ori_ori_n1259_));
  NA2        o1210(.A(ori_ori_n752_), .B(ori_ori_n363_), .Y(ori_ori_n1260_));
  OAI210     o1211(.A0(ori_ori_n1237_), .A1(ori_ori_n1229_), .B0(ori_ori_n263_), .Y(ori_ori_n1261_));
  OAI210     o1212(.A0(ori_ori_n1260_), .A1(ori_ori_n764_), .B0(ori_ori_n1261_), .Y(ori_ori_n1262_));
  OAI210     o1213(.A0(ori_ori_n1262_), .A1(ori_ori_n1259_), .B0(x6), .Y(ori_ori_n1263_));
  NO2        o1214(.A(ori_ori_n57_), .B(ori_ori_n59_), .Y(ori_ori_n1264_));
  NO2        o1215(.A(x7), .B(x5), .Y(ori_ori_n1265_));
  AOI220     o1216(.A0(ori_ori_n773_), .A1(ori_ori_n1264_), .B0(ori_ori_n489_), .B1(ori_ori_n1265_), .Y(ori_ori_n1266_));
  NA2        o1217(.A(ori_ori_n689_), .B(ori_ori_n263_), .Y(ori_ori_n1267_));
  NA3        o1218(.A(ori_ori_n563_), .B(ori_ori_n265_), .C(ori_ori_n220_), .Y(ori_ori_n1268_));
  NA3        o1219(.A(ori_ori_n1268_), .B(ori_ori_n1267_), .C(ori_ori_n1266_), .Y(ori_ori_n1269_));
  NA2        o1220(.A(ori_ori_n1269_), .B(ori_ori_n381_), .Y(ori_ori_n1270_));
  AOI210     o1221(.A0(ori_ori_n339_), .A1(ori_ori_n311_), .B0(ori_ori_n55_), .Y(ori_ori_n1271_));
  NA4        o1222(.A(ori_ori_n1271_), .B(ori_ori_n1270_), .C(ori_ori_n1263_), .D(ori_ori_n1257_), .Y(ori_ori_n1272_));
  AO220      o1223(.A0(ori_ori_n1272_), .A1(ori_ori_n1243_), .B0(ori_ori_n1212_), .B1(ori_ori_n1206_), .Y(ori16));
  NO2        o1224(.A(x4), .B(ori_ori_n59_), .Y(ori_ori_n1274_));
  NA2        o1225(.A(ori_ori_n602_), .B(ori_ori_n486_), .Y(ori_ori_n1275_));
  NA3        o1226(.A(ori_ori_n212_), .B(ori_ori_n388_), .C(ori_ori_n871_), .Y(ori_ori_n1276_));
  NA2        o1227(.A(ori_ori_n127_), .B(ori_ori_n190_), .Y(ori_ori_n1277_));
  AOI210     o1228(.A0(ori_ori_n1276_), .A1(ori_ori_n1275_), .B0(ori_ori_n1277_), .Y(ori_ori_n1278_));
  NO3        o1229(.A(x8), .B(x6), .C(ori_ori_n50_), .Y(ori_ori_n1279_));
  NO2        o1230(.A(ori_ori_n668_), .B(ori_ori_n170_), .Y(ori_ori_n1280_));
  OAI210     o1231(.A0(ori_ori_n1279_), .A1(ori_ori_n218_), .B0(ori_ori_n1280_), .Y(ori_ori_n1281_));
  NO2        o1232(.A(ori_ori_n148_), .B(x5), .Y(ori_ori_n1282_));
  NA3        o1233(.A(ori_ori_n527_), .B(ori_ori_n488_), .C(ori_ori_n431_), .Y(ori_ori_n1283_));
  NA2        o1234(.A(ori_ori_n1283_), .B(ori_ori_n1281_), .Y(ori_ori_n1284_));
  OAI210     o1235(.A0(ori_ori_n1284_), .A1(ori_ori_n1278_), .B0(ori_ori_n1274_), .Y(ori_ori_n1285_));
  NO2        o1236(.A(ori_ori_n292_), .B(x7), .Y(ori_ori_n1286_));
  NA2        o1237(.A(ori_ori_n985_), .B(ori_ori_n183_), .Y(ori_ori_n1287_));
  NA2        o1238(.A(ori_ori_n55_), .B(ori_ori_n104_), .Y(ori_ori_n1288_));
  NA2        o1239(.A(ori_ori_n1288_), .B(ori_ori_n623_), .Y(ori_ori_n1289_));
  NA2        o1240(.A(ori_ori_n338_), .B(ori_ori_n989_), .Y(ori_ori_n1290_));
  OA220      o1241(.A0(ori_ori_n1290_), .A1(ori_ori_n1289_), .B0(ori_ori_n1287_), .B1(ori_ori_n577_), .Y(ori_ori_n1291_));
  NO2        o1242(.A(ori_ori_n1291_), .B(ori_ori_n592_), .Y(ori_ori_n1292_));
  INV        o1243(.A(ori_ori_n933_), .Y(ori_ori_n1293_));
  NO2        o1244(.A(ori_ori_n1293_), .B(ori_ori_n62_), .Y(ori_ori_n1294_));
  NA2        o1245(.A(ori_ori_n1154_), .B(ori_ori_n122_), .Y(ori_ori_n1295_));
  NA2        o1246(.A(ori_ori_n580_), .B(ori_ori_n330_), .Y(ori_ori_n1296_));
  NA2        o1247(.A(ori_ori_n418_), .B(ori_ori_n534_), .Y(ori_ori_n1297_));
  OAI220     o1248(.A0(ori_ori_n1297_), .A1(ori_ori_n1296_), .B0(ori_ori_n1295_), .B1(ori_ori_n283_), .Y(ori_ori_n1298_));
  NO2        o1249(.A(ori_ori_n1298_), .B(ori_ori_n1292_), .Y(ori_ori_n1299_));
  NA4        o1250(.A(ori_ori_n644_), .B(ori_ori_n170_), .C(ori_ori_n58_), .D(x6), .Y(ori_ori_n1300_));
  NO2        o1251(.A(ori_ori_n1300_), .B(ori_ori_n54_), .Y(ori_ori_n1301_));
  NO2        o1252(.A(ori_ori_n659_), .B(x3), .Y(ori_ori_n1302_));
  NO2        o1253(.A(ori_ori_n689_), .B(ori_ori_n462_), .Y(ori_ori_n1303_));
  NO3        o1254(.A(ori_ori_n1303_), .B(ori_ori_n235_), .C(ori_ori_n143_), .Y(ori_ori_n1304_));
  NO2        o1255(.A(ori_ori_n1304_), .B(ori_ori_n1301_), .Y(ori_ori_n1305_));
  NA2        o1256(.A(ori_ori_n364_), .B(ori_ori_n871_), .Y(ori_ori_n1306_));
  NA4        o1257(.A(ori_ori_n433_), .B(ori_ori_n335_), .C(ori_ori_n203_), .D(x6), .Y(ori_ori_n1307_));
  INV        o1258(.A(ori_ori_n1307_), .Y(ori_ori_n1308_));
  NA2        o1259(.A(ori_ori_n824_), .B(ori_ori_n1193_), .Y(ori_ori_n1309_));
  NA2        o1260(.A(ori_ori_n665_), .B(x7), .Y(ori_ori_n1310_));
  INV        o1261(.A(ori_ori_n1309_), .Y(ori_ori_n1311_));
  NA2        o1262(.A(ori_ori_n249_), .B(x2), .Y(ori_ori_n1312_));
  NO3        o1263(.A(ori_ori_n1312_), .B(ori_ori_n542_), .C(ori_ori_n72_), .Y(ori_ori_n1313_));
  BUFFER     o1264(.A(ori_ori_n702_), .Y(ori_ori_n1314_));
  AOI210     o1265(.A0(ori_ori_n527_), .A1(ori_ori_n50_), .B0(ori_ori_n537_), .Y(ori_ori_n1315_));
  OAI210     o1266(.A0(ori_ori_n841_), .A1(ori_ori_n858_), .B0(ori_ori_n343_), .Y(ori_ori_n1316_));
  OAI220     o1267(.A0(ori_ori_n1316_), .A1(ori_ori_n1315_), .B0(ori_ori_n1314_), .B1(ori_ori_n175_), .Y(ori_ori_n1317_));
  NO4        o1268(.A(ori_ori_n1317_), .B(ori_ori_n1313_), .C(ori_ori_n1311_), .D(ori_ori_n1308_), .Y(ori_ori_n1318_));
  OA220      o1269(.A0(ori_ori_n1318_), .A1(ori_ori_n400_), .B0(ori_ori_n1305_), .B1(ori_ori_n189_), .Y(ori_ori_n1319_));
  NO2        o1270(.A(ori_ori_n837_), .B(ori_ori_n55_), .Y(ori_ori_n1320_));
  NA2        o1271(.A(ori_ori_n375_), .B(ori_ori_n726_), .Y(ori_ori_n1321_));
  NO2        o1272(.A(ori_ori_n1321_), .B(ori_ori_n1320_), .Y(ori_ori_n1322_));
  NO3        o1273(.A(ori_ori_n872_), .B(ori_ori_n304_), .C(x8), .Y(ori_ori_n1323_));
  OAI210     o1274(.A0(ori_ori_n1323_), .A1(ori_ori_n1322_), .B0(x6), .Y(ori_ori_n1324_));
  NO2        o1275(.A(ori_ori_n999_), .B(ori_ori_n965_), .Y(ori_ori_n1325_));
  NA2        o1276(.A(ori_ori_n175_), .B(x7), .Y(ori_ori_n1326_));
  OAI220     o1277(.A0(ori_ori_n1326_), .A1(ori_ori_n1325_), .B0(ori_ori_n691_), .B1(ori_ori_n87_), .Y(ori_ori_n1327_));
  NA2        o1278(.A(ori_ori_n1327_), .B(ori_ori_n841_), .Y(ori_ori_n1328_));
  NA2        o1279(.A(ori_ori_n792_), .B(ori_ori_n71_), .Y(ori_ori_n1329_));
  INV        o1280(.A(ori_ori_n922_), .Y(ori_ori_n1330_));
  AOI210     o1281(.A0(ori_ori_n450_), .A1(ori_ori_n57_), .B0(ori_ori_n577_), .Y(ori_ori_n1331_));
  NA2        o1282(.A(ori_ori_n1331_), .B(ori_ori_n1330_), .Y(ori_ori_n1332_));
  NA3        o1283(.A(ori_ori_n1332_), .B(ori_ori_n1328_), .C(ori_ori_n1324_), .Y(ori_ori_n1333_));
  NA2        o1284(.A(ori_ori_n343_), .B(ori_ori_n341_), .Y(ori_ori_n1334_));
  AN2        o1285(.A(ori_ori_n1334_), .B(ori_ori_n125_), .Y(ori_ori_n1335_));
  NO3        o1286(.A(ori_ori_n402_), .B(ori_ori_n346_), .C(x7), .Y(ori_ori_n1336_));
  NO3        o1287(.A(ori_ori_n148_), .B(ori_ori_n75_), .C(x2), .Y(ori_ori_n1337_));
  NO3        o1288(.A(ori_ori_n1337_), .B(ori_ori_n1336_), .C(ori_ori_n1335_), .Y(ori_ori_n1338_));
  NO2        o1289(.A(ori_ori_n212_), .B(x1), .Y(ori_ori_n1339_));
  OAI210     o1290(.A0(ori_ori_n1339_), .A1(ori_ori_n407_), .B0(ori_ori_n462_), .Y(ori_ori_n1340_));
  NO2        o1291(.A(ori_ori_n57_), .B(ori_ori_n104_), .Y(ori_ori_n1341_));
  NA2        o1292(.A(ori_ori_n992_), .B(ori_ori_n1341_), .Y(ori_ori_n1342_));
  AOI210     o1293(.A0(ori_ori_n1342_), .A1(ori_ori_n1340_), .B0(ori_ori_n56_), .Y(ori_ori_n1343_));
  NA2        o1294(.A(ori_ori_n691_), .B(ori_ori_n699_), .Y(ori_ori_n1344_));
  NO2        o1295(.A(ori_ori_n1344_), .B(ori_ori_n1193_), .Y(ori_ori_n1345_));
  NO3        o1296(.A(ori_ori_n485_), .B(ori_ori_n159_), .C(ori_ori_n965_), .Y(ori_ori_n1346_));
  NA2        o1297(.A(ori_ori_n858_), .B(x4), .Y(ori_ori_n1347_));
  NO2        o1298(.A(ori_ori_n1347_), .B(ori_ori_n628_), .Y(ori_ori_n1348_));
  NO4        o1299(.A(ori_ori_n1348_), .B(ori_ori_n1346_), .C(ori_ori_n1345_), .D(ori_ori_n1343_), .Y(ori_ori_n1349_));
  OAI210     o1300(.A0(ori_ori_n1338_), .A1(x5), .B0(ori_ori_n1349_), .Y(ori_ori_n1350_));
  AOI220     o1301(.A0(ori_ori_n1350_), .A1(ori_ori_n95_), .B0(ori_ori_n1333_), .B1(ori_ori_n311_), .Y(ori_ori_n1351_));
  NA4        o1302(.A(ori_ori_n1351_), .B(ori_ori_n1319_), .C(ori_ori_n1299_), .D(ori_ori_n1285_), .Y(ori17));
  NO2        o1303(.A(ori_ori_n121_), .B(ori_ori_n1066_), .Y(ori_ori_n1353_));
  NA2        o1304(.A(ori_ori_n1353_), .B(ori_ori_n654_), .Y(ori_ori_n1354_));
  NA2        o1305(.A(ori_ori_n152_), .B(ori_ori_n78_), .Y(ori_ori_n1355_));
  NOi21      o1306(.An(ori_ori_n341_), .B(ori_ori_n84_), .Y(ori_ori_n1356_));
  OAI210     o1307(.A0(ori_ori_n570_), .A1(ori_ori_n55_), .B0(ori_ori_n1356_), .Y(ori_ori_n1357_));
  NA2        o1308(.A(ori_ori_n1119_), .B(ori_ori_n928_), .Y(ori_ori_n1358_));
  NA4        o1309(.A(ori_ori_n1358_), .B(ori_ori_n1357_), .C(ori_ori_n668_), .D(ori_ori_n57_), .Y(ori_ori_n1359_));
  OAI210     o1310(.A0(ori_ori_n644_), .A1(x8), .B0(ori_ori_n1193_), .Y(ori_ori_n1360_));
  NA3        o1311(.A(ori_ori_n1360_), .B(ori_ori_n1140_), .C(ori_ori_n357_), .Y(ori_ori_n1361_));
  NA3        o1312(.A(ori_ori_n352_), .B(ori_ori_n244_), .C(ori_ori_n533_), .Y(ori_ori_n1362_));
  NA4        o1313(.A(ori_ori_n682_), .B(ori_ori_n1362_), .C(ori_ori_n1361_), .D(ori_ori_n1359_), .Y(ori_ori_n1363_));
  AOI210     o1314(.A0(ori_ori_n1363_), .A1(x1), .B0(ori_ori_n59_), .Y(ori_ori_n1364_));
  NO2        o1315(.A(ori_ori_n896_), .B(ori_ori_n450_), .Y(ori_ori_n1365_));
  OAI210     o1316(.A0(ori_ori_n1365_), .A1(ori_ori_n975_), .B0(ori_ori_n555_), .Y(ori_ori_n1366_));
  NO3        o1317(.A(ori_ori_n577_), .B(ori_ori_n505_), .C(ori_ori_n476_), .Y(ori_ori_n1367_));
  OAI210     o1318(.A0(ori_ori_n1367_), .A1(ori_ori_n823_), .B0(ori_ori_n1302_), .Y(ori_ori_n1368_));
  AOI210     o1319(.A0(ori_ori_n1368_), .A1(ori_ori_n1366_), .B0(x8), .Y(ori_ori_n1369_));
  NO2        o1320(.A(ori_ori_n134_), .B(ori_ori_n133_), .Y(ori_ori_n1370_));
  NO3        o1321(.A(ori_ori_n819_), .B(ori_ori_n699_), .C(ori_ori_n638_), .Y(ori_ori_n1371_));
  AOI210     o1322(.A0(ori_ori_n1371_), .A1(ori_ori_n1370_), .B0(x0), .Y(ori_ori_n1372_));
  INV        o1323(.A(ori_ori_n1372_), .Y(ori_ori_n1373_));
  NO2        o1324(.A(ori_ori_n1373_), .B(ori_ori_n1369_), .Y(ori_ori_n1374_));
  OAI220     o1325(.A0(ori_ori_n1374_), .A1(ori_ori_n1364_), .B0(ori_ori_n1355_), .B1(ori_ori_n1354_), .Y(ori18));
  AOI210     o1326(.A0(x8), .A1(x0), .B0(x5), .Y(ori_ori_n1376_));
  NOi31      o1327(.An(ori_ori_n279_), .B(ori_ori_n1376_), .C(ori_ori_n964_), .Y(ori_ori_n1377_));
  NA2        o1328(.A(ori_ori_n549_), .B(ori_ori_n59_), .Y(ori_ori_n1378_));
  AOI210     o1329(.A0(ori_ori_n1287_), .A1(ori_ori_n319_), .B0(ori_ori_n1378_), .Y(ori_ori_n1379_));
  NO2        o1330(.A(ori_ori_n564_), .B(ori_ori_n700_), .Y(ori_ori_n1380_));
  NO4        o1331(.A(ori_ori_n231_), .B(ori_ori_n736_), .C(ori_ori_n142_), .D(ori_ori_n70_), .Y(ori_ori_n1381_));
  NO4        o1332(.A(ori_ori_n1381_), .B(ori_ori_n1380_), .C(ori_ori_n1379_), .D(ori_ori_n1377_), .Y(ori_ori_n1382_));
  NA3        o1333(.A(ori_ori_n471_), .B(ori_ori_n198_), .C(x0), .Y(ori_ori_n1383_));
  NAi21      o1334(.An(ori_ori_n347_), .B(ori_ori_n1383_), .Y(ori_ori_n1384_));
  OA220      o1335(.A0(ori_ori_n471_), .A1(ori_ori_n304_), .B0(ori_ori_n357_), .B1(x5), .Y(ori_ori_n1385_));
  NO2        o1336(.A(ori_ori_n1385_), .B(ori_ori_n267_), .Y(ori_ori_n1386_));
  AOI210     o1337(.A0(ori_ori_n1384_), .A1(ori_ori_n265_), .B0(ori_ori_n1386_), .Y(ori_ori_n1387_));
  AOI210     o1338(.A0(ori_ori_n1387_), .A1(ori_ori_n1382_), .B0(x6), .Y(ori_ori_n1388_));
  NA3        o1339(.A(ori_ori_n475_), .B(ori_ori_n378_), .C(x2), .Y(ori_ori_n1389_));
  NA2        o1340(.A(ori_ori_n964_), .B(ori_ori_n57_), .Y(ori_ori_n1390_));
  AOI210     o1341(.A0(ori_ori_n1390_), .A1(ori_ori_n1389_), .B0(ori_ori_n712_), .Y(ori_ori_n1391_));
  AOI210     o1342(.A0(ori_ori_n382_), .A1(ori_ori_n130_), .B0(ori_ori_n710_), .Y(ori_ori_n1392_));
  NA2        o1343(.A(ori_ori_n244_), .B(x6), .Y(ori_ori_n1393_));
  NA2        o1344(.A(ori_ori_n106_), .B(ori_ori_n1051_), .Y(ori_ori_n1394_));
  OAI220     o1345(.A0(ori_ori_n1394_), .A1(ori_ori_n1393_), .B0(ori_ori_n1392_), .B1(ori_ori_n674_), .Y(ori_ori_n1395_));
  OAI210     o1346(.A0(ori_ori_n1395_), .A1(ori_ori_n1391_), .B0(ori_ori_n53_), .Y(ori_ori_n1396_));
  NO2        o1347(.A(ori_ori_n627_), .B(ori_ori_n238_), .Y(ori_ori_n1397_));
  NO2        o1348(.A(ori_ori_n241_), .B(x3), .Y(ori_ori_n1398_));
  NO3        o1349(.A(ori_ori_n392_), .B(ori_ori_n549_), .C(ori_ori_n757_), .Y(ori_ori_n1399_));
  OAI210     o1350(.A0(ori_ori_n1399_), .A1(ori_ori_n1397_), .B0(ori_ori_n1398_), .Y(ori_ori_n1400_));
  AOI210     o1351(.A0(ori_ori_n1054_), .A1(ori_ori_n563_), .B0(x4), .Y(ori_ori_n1401_));
  OAI210     o1352(.A0(ori_ori_n505_), .A1(ori_ori_n549_), .B0(ori_ori_n59_), .Y(ori_ori_n1402_));
  OAI210     o1353(.A0(ori_ori_n570_), .A1(ori_ori_n588_), .B0(ori_ori_n1402_), .Y(ori_ori_n1403_));
  AO220      o1354(.A0(ori_ori_n1156_), .A1(ori_ori_n668_), .B0(ori_ori_n506_), .B1(ori_ori_n324_), .Y(ori_ori_n1404_));
  AOI220     o1355(.A0(ori_ori_n1404_), .A1(x1), .B0(ori_ori_n1403_), .B1(ori_ori_n149_), .Y(ori_ori_n1405_));
  NA4        o1356(.A(ori_ori_n1405_), .B(ori_ori_n1401_), .C(ori_ori_n1400_), .D(ori_ori_n1396_), .Y(ori_ori_n1406_));
  NO2        o1357(.A(ori_ori_n982_), .B(ori_ori_n124_), .Y(ori_ori_n1407_));
  OAI210     o1358(.A0(ori_ori_n1407_), .A1(ori_ori_n593_), .B0(ori_ori_n104_), .Y(ori_ori_n1408_));
  AOI210     o1359(.A0(ori_ori_n1408_), .A1(ori_ori_n511_), .B0(ori_ori_n712_), .Y(ori_ori_n1409_));
  NA3        o1360(.A(ori_ori_n1111_), .B(ori_ori_n175_), .C(ori_ori_n132_), .Y(ori_ori_n1410_));
  NA3        o1361(.A(ori_ori_n985_), .B(ori_ori_n701_), .C(ori_ori_n314_), .Y(ori_ori_n1411_));
  NA2        o1362(.A(ori_ori_n157_), .B(ori_ori_n699_), .Y(ori_ori_n1412_));
  OAI210     o1363(.A0(ori_ori_n1412_), .A1(ori_ori_n1203_), .B0(ori_ori_n1411_), .Y(ori_ori_n1413_));
  AOI210     o1364(.A0(ori_ori_n1410_), .A1(ori_ori_n163_), .B0(ori_ori_n1413_), .Y(ori_ori_n1414_));
  OAI210     o1365(.A0(ori_ori_n1414_), .A1(ori_ori_n494_), .B0(x4), .Y(ori_ori_n1415_));
  OAI220     o1366(.A0(ori_ori_n1415_), .A1(ori_ori_n1409_), .B0(ori_ori_n1406_), .B1(ori_ori_n1388_), .Y(ori_ori_n1416_));
  NO2        o1367(.A(ori_ori_n136_), .B(ori_ori_n119_), .Y(ori_ori_n1417_));
  NO2        o1368(.A(ori_ori_n175_), .B(ori_ori_n726_), .Y(ori_ori_n1418_));
  AOI210     o1369(.A0(ori_ori_n550_), .A1(ori_ori_n462_), .B0(ori_ori_n1418_), .Y(ori_ori_n1419_));
  NO2        o1370(.A(ori_ori_n1419_), .B(x6), .Y(ori_ori_n1420_));
  NO2        o1371(.A(ori_ori_n346_), .B(ori_ori_n230_), .Y(ori_ori_n1421_));
  NO2        o1372(.A(ori_ori_n125_), .B(ori_ori_n670_), .Y(ori_ori_n1422_));
  NO2        o1373(.A(ori_ori_n872_), .B(ori_ori_n533_), .Y(ori_ori_n1423_));
  AO220      o1374(.A0(ori_ori_n1423_), .A1(ori_ori_n1422_), .B0(ori_ori_n1421_), .B1(ori_ori_n121_), .Y(ori_ori_n1424_));
  NO3        o1375(.A(ori_ori_n1424_), .B(ori_ori_n1420_), .C(ori_ori_n1417_), .Y(ori_ori_n1425_));
  NA2        o1376(.A(ori_ori_n982_), .B(x3), .Y(ori_ori_n1426_));
  NA2        o1377(.A(ori_ori_n1240_), .B(ori_ori_n127_), .Y(ori_ori_n1427_));
  OAI220     o1378(.A0(ori_ori_n1427_), .A1(ori_ori_n1426_), .B0(ori_ori_n1425_), .B1(x3), .Y(ori_ori_n1428_));
  NO3        o1379(.A(ori_ori_n918_), .B(ori_ori_n627_), .C(ori_ori_n299_), .Y(ori_ori_n1429_));
  AO210      o1380(.A0(ori_ori_n947_), .A1(ori_ori_n272_), .B0(ori_ori_n1429_), .Y(ori_ori_n1430_));
  AOI220     o1381(.A0(ori_ori_n1430_), .A1(x8), .B0(ori_ori_n1240_), .B1(ori_ori_n393_), .Y(ori_ori_n1431_));
  NA2        o1382(.A(ori_ori_n678_), .B(ori_ori_n291_), .Y(ori_ori_n1432_));
  NO4        o1383(.A(ori_ori_n334_), .B(ori_ori_n187_), .C(ori_ori_n310_), .D(x2), .Y(ori_ori_n1433_));
  NA2        o1384(.A(ori_ori_n1288_), .B(ori_ori_n106_), .Y(ori_ori_n1434_));
  NO3        o1385(.A(ori_ori_n1113_), .B(ori_ori_n911_), .C(ori_ori_n1051_), .Y(ori_ori_n1435_));
  AOI210     o1386(.A0(ori_ori_n1435_), .A1(ori_ori_n1434_), .B0(ori_ori_n1433_), .Y(ori_ori_n1436_));
  OA220      o1387(.A0(ori_ori_n1436_), .A1(ori_ori_n872_), .B0(ori_ori_n1432_), .B1(ori_ori_n517_), .Y(ori_ori_n1437_));
  OAI210     o1388(.A0(ori_ori_n1431_), .A1(ori_ori_n367_), .B0(ori_ori_n1437_), .Y(ori_ori_n1438_));
  AOI210     o1389(.A0(ori_ori_n1428_), .A1(ori_ori_n130_), .B0(ori_ori_n1438_), .Y(ori_ori_n1439_));
  NA2        o1390(.A(ori_ori_n1439_), .B(ori_ori_n1416_), .Y(ori19));
  NO2        o1391(.A(ori_ori_n1329_), .B(ori_ori_n234_), .Y(ori_ori_n1441_));
  NA2        o1392(.A(ori_ori_n588_), .B(x3), .Y(ori_ori_n1442_));
  NO2        o1393(.A(ori_ori_n142_), .B(ori_ori_n105_), .Y(ori_ori_n1443_));
  NA2        o1394(.A(ori_ori_n1443_), .B(ori_ori_n220_), .Y(ori_ori_n1444_));
  NO2        o1395(.A(ori_ori_n1200_), .B(ori_ori_n157_), .Y(ori_ori_n1445_));
  INV        o1396(.A(ori_ori_n1445_), .Y(ori_ori_n1446_));
  AOI210     o1397(.A0(ori_ori_n1446_), .A1(ori_ori_n1444_), .B0(ori_ori_n56_), .Y(ori_ori_n1447_));
  NO2        o1398(.A(ori_ori_n782_), .B(ori_ori_n1126_), .Y(ori_ori_n1448_));
  OAI210     o1399(.A0(ori_ori_n1447_), .A1(ori_ori_n1441_), .B0(ori_ori_n1448_), .Y(ori_ori_n1449_));
  AOI210     o1400(.A0(ori_ori_n322_), .A1(x6), .B0(ori_ori_n118_), .Y(ori_ori_n1450_));
  NO3        o1401(.A(ori_ori_n1450_), .B(ori_ori_n687_), .C(ori_ori_n122_), .Y(ori_ori_n1451_));
  NA2        o1402(.A(ori_ori_n1106_), .B(ori_ori_n119_), .Y(ori_ori_n1452_));
  NO4        o1403(.A(ori_ori_n1452_), .B(ori_ori_n918_), .C(ori_ori_n809_), .D(ori_ori_n77_), .Y(ori_ori_n1453_));
  NO3        o1404(.A(ori_ori_n1453_), .B(ori_ori_n1451_), .C(ori_ori_n944_), .Y(ori_ori_n1454_));
  NO2        o1405(.A(ori_ori_n494_), .B(ori_ori_n567_), .Y(ori_ori_n1455_));
  NA2        o1406(.A(ori_ori_n1153_), .B(ori_ori_n50_), .Y(ori_ori_n1456_));
  NO3        o1407(.A(ori_ori_n469_), .B(ori_ori_n281_), .C(ori_ori_n64_), .Y(ori_ori_n1457_));
  AOI220     o1408(.A0(ori_ori_n1457_), .A1(ori_ori_n1456_), .B0(ori_ori_n1455_), .B1(ori_ori_n701_), .Y(ori_ori_n1458_));
  OAI210     o1409(.A0(ori_ori_n1454_), .A1(ori_ori_n57_), .B0(ori_ori_n1458_), .Y(ori_ori_n1459_));
  NA2        o1410(.A(ori_ori_n1459_), .B(ori_ori_n699_), .Y(ori_ori_n1460_));
  AOI210     o1411(.A0(ori_ori_n746_), .A1(ori_ori_n670_), .B0(ori_ori_n692_), .Y(ori_ori_n1461_));
  NO2        o1412(.A(ori_ori_n1461_), .B(x4), .Y(ori_ori_n1462_));
  NA3        o1413(.A(ori_ori_n668_), .B(ori_ori_n233_), .C(x7), .Y(ori_ori_n1463_));
  AOI220     o1414(.A0(ori_ori_n1286_), .A1(ori_ori_n712_), .B0(ori_ori_n638_), .B1(ori_ori_n1066_), .Y(ori_ori_n1464_));
  AOI210     o1415(.A0(ori_ori_n1464_), .A1(ori_ori_n1463_), .B0(ori_ori_n454_), .Y(ori_ori_n1465_));
  OAI210     o1416(.A0(ori_ori_n1465_), .A1(ori_ori_n1462_), .B0(ori_ori_n736_), .Y(ori_ori_n1466_));
  NO2        o1417(.A(ori_ori_n674_), .B(ori_ori_n295_), .Y(ori_ori_n1467_));
  NO2        o1418(.A(ori_ori_n142_), .B(ori_ori_n943_), .Y(ori_ori_n1468_));
  AOI220     o1419(.A0(ori_ori_n1468_), .A1(ori_ori_n1167_), .B0(ori_ori_n1467_), .B1(ori_ori_n432_), .Y(ori_ori_n1469_));
  AO210      o1420(.A0(ori_ori_n1469_), .A1(ori_ori_n1466_), .B0(x1), .Y(ori_ori_n1470_));
  NA2        o1421(.A(ori_ori_n577_), .B(ori_ori_n965_), .Y(ori_ori_n1471_));
  NA2        o1422(.A(ori_ori_n137_), .B(ori_ori_n107_), .Y(ori_ori_n1472_));
  NOi21      o1423(.An(x1), .B(x6), .Y(ori_ori_n1473_));
  NA2        o1424(.A(ori_ori_n1473_), .B(ori_ori_n84_), .Y(ori_ori_n1474_));
  NA3        o1425(.A(ori_ori_n1474_), .B(ori_ori_n1472_), .C(ori_ori_n1471_), .Y(ori_ori_n1475_));
  AOI220     o1426(.A0(ori_ori_n1475_), .A1(x3), .B0(ori_ori_n1114_), .B1(ori_ori_n342_), .Y(ori_ori_n1476_));
  NA2        o1427(.A(ori_ori_n1119_), .B(ori_ori_n721_), .Y(ori_ori_n1477_));
  AOI220     o1428(.A0(ori_ori_n1156_), .A1(ori_ori_n118_), .B0(ori_ori_n837_), .B1(ori_ori_n738_), .Y(ori_ori_n1478_));
  AOI210     o1429(.A0(ori_ori_n1478_), .A1(ori_ori_n1477_), .B0(ori_ori_n295_), .Y(ori_ori_n1479_));
  NA3        o1430(.A(ori_ori_n1106_), .B(ori_ori_n343_), .C(ori_ori_n106_), .Y(ori_ori_n1480_));
  NO2        o1431(.A(ori_ori_n1480_), .B(ori_ori_n881_), .Y(ori_ori_n1481_));
  NO3        o1432(.A(ori_ori_n565_), .B(ori_ori_n468_), .C(ori_ori_n1129_), .Y(ori_ori_n1482_));
  NO3        o1433(.A(ori_ori_n1482_), .B(ori_ori_n1481_), .C(ori_ori_n1479_), .Y(ori_ori_n1483_));
  OAI210     o1434(.A0(ori_ori_n1476_), .A1(ori_ori_n769_), .B0(ori_ori_n1483_), .Y(ori_ori_n1484_));
  NO2        o1435(.A(ori_ori_n505_), .B(ori_ori_n68_), .Y(ori_ori_n1485_));
  OAI220     o1436(.A0(ori_ori_n1485_), .A1(ori_ori_n1442_), .B0(ori_ori_n280_), .B1(ori_ori_n817_), .Y(ori_ori_n1486_));
  AOI220     o1437(.A0(ori_ori_n1486_), .A1(ori_ori_n56_), .B0(ori_ori_n1245_), .B1(ori_ori_n665_), .Y(ori_ori_n1487_));
  NO2        o1438(.A(ori_ori_n54_), .B(ori_ori_n71_), .Y(ori_ori_n1488_));
  AO220      o1439(.A0(ori_ori_n1488_), .A1(ori_ori_n918_), .B0(ori_ori_n738_), .B1(ori_ori_n871_), .Y(ori_ori_n1489_));
  INV        o1440(.A(ori_ori_n1473_), .Y(ori_ori_n1490_));
  NA2        o1441(.A(ori_ori_n450_), .B(ori_ori_n665_), .Y(ori_ori_n1491_));
  NO2        o1442(.A(ori_ori_n1491_), .B(ori_ori_n1490_), .Y(ori_ori_n1492_));
  AOI210     o1443(.A0(ori_ori_n1489_), .A1(x2), .B0(ori_ori_n1492_), .Y(ori_ori_n1493_));
  OAI220     o1444(.A0(ori_ori_n1493_), .A1(ori_ori_n142_), .B0(ori_ori_n1487_), .B1(ori_ori_n54_), .Y(ori_ori_n1494_));
  OAI210     o1445(.A0(ori_ori_n1494_), .A1(ori_ori_n1484_), .B0(x8), .Y(ori_ori_n1495_));
  NA4        o1446(.A(ori_ori_n1495_), .B(ori_ori_n1470_), .C(ori_ori_n1460_), .D(ori_ori_n1449_), .Y(ori20));
  NA2        o1447(.A(ori_ori_n432_), .B(ori_ori_n371_), .Y(ori_ori_n1497_));
  NO2        o1448(.A(ori_ori_n1497_), .B(ori_ori_n87_), .Y(ori_ori_n1498_));
  AOI210     o1449(.A0(ori_ori_n967_), .A1(ori_ori_n62_), .B0(ori_ori_n1455_), .Y(ori_ori_n1499_));
  AOI210     o1450(.A0(ori_ori_n905_), .A1(ori_ori_n318_), .B0(ori_ori_n1096_), .Y(ori_ori_n1500_));
  OAI210     o1451(.A0(ori_ori_n1499_), .A1(ori_ori_n623_), .B0(ori_ori_n1500_), .Y(ori_ori_n1501_));
  OAI210     o1452(.A0(ori_ori_n1501_), .A1(ori_ori_n1498_), .B0(ori_ori_n1017_), .Y(ori_ori_n1502_));
  NAi21      o1453(.An(ori_ori_n501_), .B(ori_ori_n359_), .Y(ori_ori_n1503_));
  NA3        o1454(.A(ori_ori_n1503_), .B(ori_ori_n903_), .C(ori_ori_n871_), .Y(ori_ori_n1504_));
  NA2        o1455(.A(ori_ori_n1016_), .B(ori_ori_n253_), .Y(ori_ori_n1505_));
  AOI210     o1456(.A0(ori_ori_n1505_), .A1(ori_ori_n1504_), .B0(ori_ori_n1193_), .Y(ori_ori_n1506_));
  NO2        o1457(.A(ori_ori_n678_), .B(ori_ori_n891_), .Y(ori_ori_n1507_));
  NOi31      o1458(.An(ori_ori_n1507_), .B(ori_ori_n1082_), .C(ori_ori_n481_), .Y(ori_ori_n1508_));
  OAI210     o1459(.A0(ori_ori_n1508_), .A1(ori_ori_n1506_), .B0(ori_ori_n299_), .Y(ori_ori_n1509_));
  NA2        o1460(.A(ori_ori_n291_), .B(ori_ori_n91_), .Y(ori_ori_n1510_));
  NA2        o1461(.A(ori_ori_n300_), .B(ori_ori_n104_), .Y(ori_ori_n1511_));
  INV        o1462(.A(ori_ori_n381_), .Y(ori_ori_n1512_));
  OAI220     o1463(.A0(ori_ori_n1512_), .A1(ori_ori_n1511_), .B0(ori_ori_n1510_), .B1(ori_ori_n248_), .Y(ori_ori_n1513_));
  NA2        o1464(.A(ori_ori_n1513_), .B(ori_ori_n203_), .Y(ori_ori_n1514_));
  NO2        o1465(.A(ori_ori_n607_), .B(ori_ori_n555_), .Y(ori_ori_n1515_));
  NA2        o1466(.A(ori_ori_n872_), .B(ori_ori_n50_), .Y(ori_ori_n1516_));
  NO3        o1467(.A(ori_ori_n1516_), .B(ori_ori_n333_), .C(ori_ori_n211_), .Y(ori_ori_n1517_));
  NA4        o1468(.A(ori_ori_n311_), .B(ori_ori_n218_), .C(ori_ori_n726_), .D(ori_ori_n64_), .Y(ori_ori_n1518_));
  OAI220     o1469(.A0(ori_ori_n1518_), .A1(ori_ori_n617_), .B0(ori_ori_n1347_), .B1(ori_ori_n955_), .Y(ori_ori_n1519_));
  AOI210     o1470(.A0(ori_ori_n1517_), .A1(ori_ori_n1515_), .B0(ori_ori_n1519_), .Y(ori_ori_n1520_));
  NA4        o1471(.A(ori_ori_n1520_), .B(ori_ori_n1514_), .C(ori_ori_n1509_), .D(ori_ori_n1502_), .Y(ori21));
  OAI210     o1472(.A0(ori_ori_n364_), .A1(ori_ori_n54_), .B0(x7), .Y(ori_ori_n1522_));
  OAI220     o1473(.A0(ori_ori_n1522_), .A1(ori_ori_n1185_), .B0(ori_ori_n968_), .B1(ori_ori_n92_), .Y(ori_ori_n1523_));
  NA2        o1474(.A(ori_ori_n1523_), .B(ori_ori_n78_), .Y(ori_ori_n1524_));
  NA2        o1475(.A(ori_ori_n265_), .B(ori_ori_n780_), .Y(ori_ori_n1525_));
  AOI220     o1476(.A0(ori_ori_n1525_), .A1(ori_ori_n283_), .B0(ori_ori_n517_), .B1(ori_ori_n416_), .Y(ori_ori_n1526_));
  NA2        o1477(.A(ori_ori_n858_), .B(ori_ori_n247_), .Y(ori_ori_n1527_));
  NA2        o1478(.A(ori_ori_n489_), .B(ori_ori_n417_), .Y(ori_ori_n1528_));
  NA4        o1479(.A(ori_ori_n1528_), .B(ori_ori_n1527_), .C(ori_ori_n1267_), .D(ori_ori_n56_), .Y(ori_ori_n1529_));
  NO2        o1480(.A(ori_ori_n701_), .B(ori_ori_n392_), .Y(ori_ori_n1530_));
  NO3        o1481(.A(ori_ori_n1530_), .B(ori_ori_n660_), .C(ori_ori_n227_), .Y(ori_ori_n1531_));
  NOi31      o1482(.An(ori_ori_n178_), .B(ori_ori_n577_), .C(ori_ori_n1004_), .Y(ori_ori_n1532_));
  NO4        o1483(.A(ori_ori_n1532_), .B(ori_ori_n1531_), .C(ori_ori_n1529_), .D(ori_ori_n1526_), .Y(ori_ori_n1533_));
  NO2        o1484(.A(ori_ori_n251_), .B(ori_ori_n52_), .Y(ori_ori_n1534_));
  OA210      o1485(.A0(ori_ori_n1534_), .A1(ori_ori_n806_), .B0(x3), .Y(ori_ori_n1535_));
  OAI210     o1486(.A0(ori_ori_n711_), .A1(ori_ori_n537_), .B0(ori_ori_n312_), .Y(ori_ori_n1536_));
  NO2        o1487(.A(ori_ori_n70_), .B(x2), .Y(ori_ori_n1537_));
  OAI210     o1488(.A0(ori_ori_n163_), .A1(x0), .B0(ori_ori_n1537_), .Y(ori_ori_n1538_));
  NA2        o1489(.A(ori_ori_n1538_), .B(ori_ori_n1536_), .Y(ori_ori_n1539_));
  OAI210     o1490(.A0(ori_ori_n1539_), .A1(ori_ori_n1535_), .B0(x8), .Y(ori_ori_n1540_));
  NO3        o1491(.A(ori_ori_n700_), .B(ori_ori_n568_), .C(ori_ori_n533_), .Y(ori_ori_n1541_));
  NA2        o1492(.A(ori_ori_n55_), .B(ori_ori_n50_), .Y(ori_ori_n1542_));
  MUX2       o1493(.S(ori_ori_n549_), .A(ori_ori_n1542_), .B(ori_ori_n103_), .Y(ori_ori_n1543_));
  AOI210     o1494(.A0(ori_ori_n1248_), .A1(ori_ori_n219_), .B0(ori_ori_n1543_), .Y(ori_ori_n1544_));
  OAI210     o1495(.A0(ori_ori_n586_), .A1(ori_ori_n532_), .B0(x4), .Y(ori_ori_n1545_));
  NO3        o1496(.A(ori_ori_n1545_), .B(ori_ori_n1544_), .C(ori_ori_n1541_), .Y(ori_ori_n1546_));
  AO220      o1497(.A0(ori_ori_n1546_), .A1(ori_ori_n1540_), .B0(ori_ori_n1533_), .B1(ori_ori_n1524_), .Y(ori_ori_n1547_));
  AO220      o1498(.A0(ori_ori_n578_), .A1(ori_ori_n295_), .B0(ori_ori_n538_), .B1(x8), .Y(ori_ori_n1548_));
  NO2        o1499(.A(ori_ori_n782_), .B(x0), .Y(ori_ori_n1549_));
  NO3        o1500(.A(ori_ori_n1549_), .B(ori_ori_n499_), .C(ori_ori_n88_), .Y(ori_ori_n1550_));
  NO2        o1501(.A(ori_ori_n148_), .B(x2), .Y(ori_ori_n1551_));
  NO3        o1502(.A(ori_ori_n340_), .B(ori_ori_n231_), .C(ori_ori_n170_), .Y(ori_ori_n1552_));
  AOI210     o1503(.A0(ori_ori_n1551_), .A1(ori_ori_n68_), .B0(ori_ori_n1552_), .Y(ori_ori_n1553_));
  OAI210     o1504(.A0(ori_ori_n1550_), .A1(ori_ori_n357_), .B0(ori_ori_n1553_), .Y(ori_ori_n1554_));
  AOI220     o1505(.A0(ori_ori_n1554_), .A1(x5), .B0(ori_ori_n1548_), .B1(ori_ori_n678_), .Y(ori_ori_n1555_));
  AOI210     o1506(.A0(ori_ori_n1555_), .A1(ori_ori_n1547_), .B0(ori_ori_n71_), .Y(ori_ori_n1556_));
  NO2        o1507(.A(ori_ori_n828_), .B(ori_ori_n156_), .Y(ori_ori_n1557_));
  NOi41      o1508(.An(ori_ori_n1312_), .B(ori_ori_n1376_), .C(ori_ori_n1065_), .D(ori_ori_n773_), .Y(ori_ori_n1558_));
  NA2        o1509(.A(ori_ori_n1558_), .B(ori_ori_n1557_), .Y(ori_ori_n1559_));
  NO2        o1510(.A(ori_ori_n78_), .B(x4), .Y(ori_ori_n1560_));
  OAI210     o1511(.A0(ori_ori_n263_), .A1(ori_ori_n146_), .B0(ori_ori_n1560_), .Y(ori_ori_n1561_));
  OAI210     o1512(.A0(ori_ori_n366_), .A1(ori_ori_n382_), .B0(ori_ori_n211_), .Y(ori_ori_n1562_));
  NO2        o1513(.A(ori_ori_n233_), .B(ori_ori_n50_), .Y(ori_ori_n1563_));
  NO2        o1514(.A(ori_ori_n1563_), .B(ori_ori_n57_), .Y(ori_ori_n1564_));
  NA2        o1515(.A(ori_ori_n1564_), .B(ori_ori_n1562_), .Y(ori_ori_n1565_));
  AOI210     o1516(.A0(ori_ori_n1561_), .A1(ori_ori_n1559_), .B0(ori_ori_n1565_), .Y(ori_ori_n1566_));
  NO2        o1517(.A(ori_ori_n1503_), .B(ori_ori_n1126_), .Y(ori_ori_n1567_));
  AOI220     o1518(.A0(ori_ori_n1567_), .A1(ori_ori_n1075_), .B0(ori_ori_n1217_), .B1(ori_ori_n964_), .Y(ori_ori_n1568_));
  NO2        o1519(.A(ori_ori_n1568_), .B(ori_ori_n106_), .Y(ori_ori_n1569_));
  NA2        o1520(.A(ori_ori_n272_), .B(ori_ori_n104_), .Y(ori_ori_n1570_));
  NA2        o1521(.A(ori_ori_n816_), .B(ori_ori_n55_), .Y(ori_ori_n1571_));
  NO2        o1522(.A(ori_ori_n612_), .B(ori_ori_n971_), .Y(ori_ori_n1572_));
  NO3        o1523(.A(ori_ori_n1572_), .B(ori_ori_n1569_), .C(ori_ori_n1566_), .Y(ori_ori_n1573_));
  NO2        o1524(.A(ori_ori_n1573_), .B(x6), .Y(ori_ori_n1574_));
  NO2        o1525(.A(ori_ori_n558_), .B(ori_ori_n1376_), .Y(ori_ori_n1575_));
  OAI210     o1526(.A0(ori_ori_n1575_), .A1(ori_ori_n630_), .B0(ori_ori_n56_), .Y(ori_ori_n1576_));
  NO2        o1527(.A(ori_ori_n680_), .B(ori_ori_n54_), .Y(ori_ori_n1577_));
  NO2        o1528(.A(ori_ori_n787_), .B(x5), .Y(ori_ori_n1578_));
  NO3        o1529(.A(ori_ori_n1578_), .B(ori_ori_n1577_), .C(ori_ori_n865_), .Y(ori_ori_n1579_));
  AOI210     o1530(.A0(ori_ori_n1579_), .A1(ori_ori_n1576_), .B0(ori_ori_n50_), .Y(ori_ori_n1580_));
  NA2        o1531(.A(ori_ori_n148_), .B(ori_ori_n104_), .Y(ori_ori_n1581_));
  OA210      o1532(.A0(ori_ori_n1581_), .A1(ori_ori_n395_), .B0(ori_ori_n422_), .Y(ori_ori_n1582_));
  NA3        o1533(.A(ori_ori_n55_), .B(x2), .C(x0), .Y(ori_ori_n1583_));
  AOI220     o1534(.A0(ori_ori_n1583_), .A1(ori_ori_n157_), .B0(ori_ori_n787_), .B1(ori_ori_n144_), .Y(ori_ori_n1584_));
  NO2        o1535(.A(ori_ori_n623_), .B(ori_ori_n233_), .Y(ori_ori_n1585_));
  NO3        o1536(.A(ori_ori_n223_), .B(ori_ori_n209_), .C(ori_ori_n328_), .Y(ori_ori_n1586_));
  NO3        o1537(.A(ori_ori_n1586_), .B(ori_ori_n1585_), .C(ori_ori_n1584_), .Y(ori_ori_n1587_));
  OAI220     o1538(.A0(ori_ori_n1587_), .A1(ori_ori_n56_), .B0(ori_ori_n1582_), .B1(ori_ori_n636_), .Y(ori_ori_n1588_));
  OAI210     o1539(.A0(ori_ori_n1588_), .A1(ori_ori_n1580_), .B0(ori_ori_n112_), .Y(ori_ori_n1589_));
  NO2        o1540(.A(ori_ori_n562_), .B(ori_ori_n278_), .Y(ori_ori_n1590_));
  AOI210     o1541(.A0(ori_ori_n556_), .A1(x5), .B0(ori_ori_n1590_), .Y(ori_ori_n1591_));
  NO2        o1542(.A(ori_ori_n1591_), .B(ori_ori_n106_), .Y(ori_ori_n1592_));
  NA2        o1543(.A(ori_ori_n644_), .B(ori_ori_n81_), .Y(ori_ori_n1593_));
  NA3        o1544(.A(ori_ori_n1593_), .B(ori_ori_n389_), .C(ori_ori_n57_), .Y(ori_ori_n1594_));
  OAI210     o1545(.A0(ori_ori_n1571_), .A1(ori_ori_n1570_), .B0(ori_ori_n1594_), .Y(ori_ori_n1595_));
  OAI210     o1546(.A0(ori_ori_n1595_), .A1(ori_ori_n1592_), .B0(x1), .Y(ori_ori_n1596_));
  NO4        o1547(.A(ori_ori_n375_), .B(ori_ori_n78_), .C(ori_ori_n138_), .D(x3), .Y(ori_ori_n1597_));
  NO2        o1548(.A(ori_ori_n300_), .B(ori_ori_n108_), .Y(ori_ori_n1598_));
  OAI210     o1549(.A0(ori_ori_n1597_), .A1(ori_ori_n1194_), .B0(ori_ori_n1598_), .Y(ori_ori_n1599_));
  NO2        o1550(.A(ori_ori_n60_), .B(ori_ori_n104_), .Y(ori_ori_n1600_));
  NO4        o1551(.A(ori_ori_n1570_), .B(ori_ori_n879_), .C(ori_ori_n607_), .D(ori_ori_n50_), .Y(ori_ori_n1601_));
  AOI210     o1552(.A0(ori_ori_n1600_), .A1(ori_ori_n1418_), .B0(ori_ori_n1601_), .Y(ori_ori_n1602_));
  NA4        o1553(.A(ori_ori_n1602_), .B(ori_ori_n1599_), .C(ori_ori_n1596_), .D(ori_ori_n1589_), .Y(ori_ori_n1603_));
  NO3        o1554(.A(ori_ori_n1603_), .B(ori_ori_n1574_), .C(ori_ori_n1556_), .Y(ori22));
  AOI210     o1555(.A0(ori_ori_n475_), .A1(ori_ori_n71_), .B0(ori_ori_n425_), .Y(ori_ori_n1605_));
  NO3        o1556(.A(ori_ori_n1101_), .B(ori_ori_n505_), .C(ori_ori_n638_), .Y(ori_ori_n1606_));
  AOI210     o1557(.A0(x5), .A1(x2), .B0(x8), .Y(ori_ori_n1607_));
  NA2        o1558(.A(ori_ori_n1607_), .B(ori_ori_n59_), .Y(ori_ori_n1608_));
  OAI220     o1559(.A0(ori_ori_n1608_), .A1(ori_ori_n1606_), .B0(ori_ori_n1605_), .B1(ori_ori_n357_), .Y(ori_ori_n1609_));
  NA2        o1560(.A(ori_ori_n532_), .B(ori_ori_n87_), .Y(ori_ori_n1610_));
  NA2        o1561(.A(ori_ori_n248_), .B(ori_ori_n77_), .Y(ori_ori_n1611_));
  OA220      o1562(.A0(ori_ori_n1611_), .A1(ori_ori_n1610_), .B0(ori_ori_n766_), .B1(ori_ori_n928_), .Y(ori_ori_n1612_));
  NO3        o1563(.A(ori_ori_n1150_), .B(ori_ori_n87_), .C(x0), .Y(ori_ori_n1613_));
  OAI210     o1564(.A0(ori_ori_n357_), .A1(ori_ori_n189_), .B0(x4), .Y(ori_ori_n1614_));
  NO2        o1565(.A(ori_ori_n1614_), .B(ori_ori_n1613_), .Y(ori_ori_n1615_));
  OAI210     o1566(.A0(ori_ori_n1612_), .A1(ori_ori_n183_), .B0(ori_ori_n1615_), .Y(ori_ori_n1616_));
  AOI210     o1567(.A0(ori_ori_n1609_), .A1(ori_ori_n53_), .B0(ori_ori_n1616_), .Y(ori_ori_n1617_));
  NA2        o1568(.A(ori_ori_n276_), .B(ori_ori_n281_), .Y(ori_ori_n1618_));
  NA3        o1569(.A(ori_ori_n1618_), .B(ori_ori_n203_), .C(ori_ori_n280_), .Y(ori_ori_n1619_));
  NA2        o1570(.A(ori_ori_n527_), .B(ori_ori_n222_), .Y(ori_ori_n1620_));
  NO3        o1571(.A(ori_ori_n450_), .B(ori_ori_n241_), .C(ori_ori_n196_), .Y(ori_ori_n1621_));
  NA2        o1572(.A(ori_ori_n1620_), .B(ori_ori_n1619_), .Y(ori_ori_n1622_));
  NO2        o1573(.A(ori_ori_n422_), .B(ori_ori_n235_), .Y(ori_ori_n1623_));
  OAI210     o1574(.A0(ori_ori_n999_), .A1(ori_ori_n172_), .B0(ori_ori_n56_), .Y(ori_ori_n1624_));
  NA3        o1575(.A(ori_ori_n55_), .B(ori_ori_n71_), .C(x0), .Y(ori_ori_n1625_));
  OAI220     o1576(.A0(ori_ori_n1625_), .A1(ori_ori_n971_), .B0(ori_ori_n333_), .B1(ori_ori_n195_), .Y(ori_ori_n1626_));
  NO2        o1577(.A(ori_ori_n1626_), .B(ori_ori_n1624_), .Y(ori_ori_n1627_));
  INV        o1578(.A(ori_ori_n1627_), .Y(ori_ori_n1628_));
  AOI210     o1579(.A0(ori_ori_n1622_), .A1(ori_ori_n104_), .B0(ori_ori_n1628_), .Y(ori_ori_n1629_));
  OAI210     o1580(.A0(ori_ori_n728_), .A1(ori_ori_n148_), .B0(ori_ori_n855_), .Y(ori_ori_n1630_));
  NA2        o1581(.A(ori_ori_n1630_), .B(ori_ori_n561_), .Y(ori_ori_n1631_));
  OA210      o1582(.A0(ori_ori_n1629_), .A1(ori_ori_n1617_), .B0(ori_ori_n1631_), .Y(ori_ori_n1632_));
  OAI210     o1583(.A0(ori_ori_n1084_), .A1(ori_ori_n643_), .B0(ori_ori_n634_), .Y(ori_ori_n1633_));
  NO2        o1584(.A(ori_ori_n323_), .B(x0), .Y(ori_ori_n1634_));
  NO2        o1585(.A(ori_ori_n1633_), .B(ori_ori_n357_), .Y(ori_ori_n1635_));
  NO3        o1586(.A(ori_ori_n157_), .B(ori_ori_n148_), .C(ori_ori_n62_), .Y(ori_ori_n1636_));
  OAI210     o1587(.A0(ori_ori_n1636_), .A1(ori_ori_n377_), .B0(ori_ori_n106_), .Y(ori_ori_n1637_));
  NA2        o1588(.A(ori_ori_n132_), .B(ori_ori_n712_), .Y(ori_ori_n1638_));
  NA2        o1589(.A(ori_ori_n375_), .B(x3), .Y(ori_ori_n1639_));
  NAi31      o1590(.An(ori_ori_n1639_), .B(ori_ori_n1638_), .C(ori_ori_n1434_), .Y(ori_ori_n1640_));
  NO3        o1591(.A(ori_ori_n782_), .B(ori_ori_n421_), .C(ori_ori_n106_), .Y(ori_ori_n1641_));
  NA2        o1592(.A(ori_ori_n1641_), .B(ori_ori_n1634_), .Y(ori_ori_n1642_));
  NA3        o1593(.A(ori_ori_n371_), .B(ori_ori_n91_), .C(ori_ori_n81_), .Y(ori_ori_n1643_));
  NO2        o1594(.A(ori_ori_n413_), .B(ori_ori_n447_), .Y(ori_ori_n1644_));
  NA2        o1595(.A(ori_ori_n1086_), .B(x3), .Y(ori_ori_n1645_));
  OAI210     o1596(.A0(ori_ori_n1645_), .A1(ori_ori_n1644_), .B0(ori_ori_n1643_), .Y(ori_ori_n1646_));
  NA3        o1597(.A(ori_ori_n56_), .B(ori_ori_n50_), .C(x0), .Y(ori_ori_n1647_));
  BUFFER     o1598(.A(ori_ori_n83_), .Y(ori_ori_n1648_));
  NA3        o1599(.A(x6), .B(x4), .C(ori_ori_n50_), .Y(ori_ori_n1649_));
  NA3        o1600(.A(ori_ori_n1649_), .B(ori_ori_n911_), .C(ori_ori_n242_), .Y(ori_ori_n1650_));
  OAI220     o1601(.A0(ori_ori_n1650_), .A1(ori_ori_n1648_), .B0(ori_ori_n974_), .B1(ori_ori_n1647_), .Y(ori_ori_n1651_));
  AOI220     o1602(.A0(ori_ori_n1651_), .A1(ori_ori_n985_), .B0(ori_ori_n1646_), .B1(ori_ori_n318_), .Y(ori_ori_n1652_));
  NA4        o1603(.A(ori_ori_n1652_), .B(ori_ori_n1642_), .C(ori_ori_n1640_), .D(ori_ori_n1637_), .Y(ori_ori_n1653_));
  AOI210     o1604(.A0(ori_ori_n1653_), .A1(x7), .B0(ori_ori_n1635_), .Y(ori_ori_n1654_));
  OAI210     o1605(.A0(ori_ori_n1632_), .A1(x7), .B0(ori_ori_n1654_), .Y(ori23));
  OR2        o1606(.A(ori_ori_n469_), .B(ori_ori_n203_), .Y(ori_ori_n1656_));
  AOI220     o1607(.A0(ori_ori_n1656_), .A1(ori_ori_n1507_), .B0(ori_ori_n563_), .B1(ori_ori_n268_), .Y(ori_ori_n1657_));
  NO3        o1608(.A(ori_ori_n766_), .B(ori_ori_n541_), .C(ori_ori_n440_), .Y(ori_ori_n1658_));
  NO3        o1609(.A(ori_ori_n873_), .B(ori_ori_n139_), .C(ori_ori_n113_), .Y(ori_ori_n1659_));
  AOI210     o1610(.A0(ori_ori_n1659_), .A1(ori_ori_n950_), .B0(ori_ori_n1658_), .Y(ori_ori_n1660_));
  OAI210     o1611(.A0(ori_ori_n1657_), .A1(ori_ori_n142_), .B0(ori_ori_n1660_), .Y(ori_ori_n1661_));
  NA2        o1612(.A(ori_ori_n1661_), .B(ori_ori_n55_), .Y(ori_ori_n1662_));
  NO2        o1613(.A(ori_ori_n879_), .B(ori_ori_n467_), .Y(ori_ori_n1663_));
  AO220      o1614(.A0(ori_ori_n1181_), .A1(ori_ori_n167_), .B0(ori_ori_n918_), .B1(ori_ori_n678_), .Y(ori_ori_n1664_));
  OAI210     o1615(.A0(ori_ori_n1664_), .A1(ori_ori_n1663_), .B0(ori_ori_n538_), .Y(ori_ori_n1665_));
  NA3        o1616(.A(ori_ori_n791_), .B(ori_ori_n382_), .C(ori_ori_n233_), .Y(ori_ori_n1666_));
  AOI210     o1617(.A0(ori_ori_n1666_), .A1(ori_ori_n452_), .B0(ori_ori_n343_), .Y(ori_ori_n1667_));
  NA2        o1618(.A(ori_ori_n1667_), .B(ori_ori_n272_), .Y(ori_ori_n1668_));
  NA3        o1619(.A(ori_ori_n57_), .B(x4), .C(x3), .Y(ori_ori_n1669_));
  NO3        o1620(.A(ori_ori_n1669_), .B(ori_ori_n675_), .C(ori_ori_n132_), .Y(ori_ori_n1670_));
  INV        o1621(.A(ori_ori_n1670_), .Y(ori_ori_n1671_));
  NA4        o1622(.A(ori_ori_n1671_), .B(ori_ori_n1668_), .C(ori_ori_n1665_), .D(ori_ori_n1662_), .Y(ori24));
  NO2        o1623(.A(ori_ori_n220_), .B(x1), .Y(ori_ori_n1673_));
  NA2        o1624(.A(ori_ori_n311_), .B(ori_ori_n444_), .Y(ori_ori_n1674_));
  BUFFER     o1625(.A(ori_ori_n1673_), .Y(ori_ori_n1675_));
  NO3        o1626(.A(ori_ori_n494_), .B(ori_ori_n626_), .C(ori_ori_n144_), .Y(ori_ori_n1676_));
  AOI210     o1627(.A0(ori_ori_n1675_), .A1(ori_ori_n91_), .B0(ori_ori_n1676_), .Y(ori_ori_n1677_));
  NA2        o1628(.A(ori_ori_n98_), .B(x8), .Y(ori_ori_n1678_));
  AN2        o1629(.A(ori_ori_n1169_), .B(ori_ori_n299_), .Y(ori_ori_n1679_));
  NA2        o1630(.A(ori_ori_n413_), .B(x8), .Y(ori_ori_n1680_));
  NA2        o1631(.A(ori_ori_n608_), .B(ori_ori_n121_), .Y(ori_ori_n1681_));
  OAI220     o1632(.A0(ori_ori_n1681_), .A1(ori_ori_n1321_), .B0(ori_ori_n1680_), .B1(ori_ori_n764_), .Y(ori_ori_n1682_));
  AOI220     o1633(.A0(ori_ori_n1682_), .A1(ori_ori_n1563_), .B0(ori_ori_n1679_), .B1(ori_ori_n950_), .Y(ori_ori_n1683_));
  OAI210     o1634(.A0(ori_ori_n1678_), .A1(ori_ori_n1677_), .B0(ori_ori_n1683_), .Y(ori25));
  NA2        o1635(.A(ori_ori_n300_), .B(ori_ori_n59_), .Y(ori_ori_n1685_));
  NO2        o1636(.A(ori_ori_n1279_), .B(ori_ori_n406_), .Y(ori_ori_n1686_));
  NO3        o1637(.A(ori_ori_n1686_), .B(ori_ori_n485_), .C(ori_ori_n95_), .Y(ori_ori_n1687_));
  NA2        o1638(.A(ori_ori_n462_), .B(ori_ori_n55_), .Y(ori_ori_n1688_));
  NO2        o1639(.A(ori_ori_n1688_), .B(ori_ori_n220_), .Y(ori_ori_n1689_));
  OAI210     o1640(.A0(ori_ori_n1689_), .A1(ori_ori_n1687_), .B0(ori_ori_n580_), .Y(ori_ori_n1690_));
  NA2        o1641(.A(ori_ori_n1623_), .B(ori_ori_n1045_), .Y(ori_ori_n1691_));
  NA2        o1642(.A(ori_ori_n1691_), .B(ori_ori_n1690_), .Y(ori_ori_n1692_));
  AN2        o1643(.A(ori_ori_n1692_), .B(ori_ori_n104_), .Y(ori26));
  NA2        o1644(.A(ori_ori_n699_), .B(ori_ori_n50_), .Y(ori_ori_n1694_));
  OAI220     o1645(.A0(ori_ori_n278_), .A1(ori_ori_n227_), .B0(ori_ori_n1694_), .B1(x7), .Y(ori_ori_n1695_));
  AOI220     o1646(.A0(ori_ori_n1695_), .A1(ori_ori_n91_), .B0(ori_ori_n1194_), .B1(ori_ori_n1051_), .Y(ori_ori_n1696_));
  NA2        o1647(.A(ori_ori_n571_), .B(ori_ori_n527_), .Y(ori_ori_n1697_));
  OAI210     o1648(.A0(ori_ori_n578_), .A1(ori_ori_n571_), .B0(ori_ori_n678_), .Y(ori_ori_n1698_));
  AOI210     o1649(.A0(ori_ori_n1697_), .A1(ori_ori_n1113_), .B0(ori_ori_n1698_), .Y(ori_ori_n1699_));
  NO2        o1650(.A(ori_ori_n1001_), .B(ori_ori_n75_), .Y(ori_ori_n1700_));
  NA2        o1651(.A(ori_ori_n736_), .B(ori_ori_n163_), .Y(ori_ori_n1701_));
  NA2        o1652(.A(ori_ori_n550_), .B(ori_ori_n462_), .Y(ori_ori_n1702_));
  NO2        o1653(.A(ori_ori_n128_), .B(ori_ori_n125_), .Y(ori_ori_n1703_));
  NA2        o1654(.A(ori_ori_n678_), .B(x3), .Y(ori_ori_n1704_));
  NO2        o1655(.A(ori_ori_n1702_), .B(ori_ori_n1704_), .Y(ori_ori_n1705_));
  NO2        o1656(.A(ori_ori_n928_), .B(x3), .Y(ori_ori_n1706_));
  AOI210     o1657(.A0(ori_ori_n404_), .A1(ori_ori_n104_), .B0(ori_ori_n1706_), .Y(ori_ori_n1707_));
  NA3        o1658(.A(ori_ori_n518_), .B(ori_ori_n51_), .C(ori_ori_n56_), .Y(ori_ori_n1708_));
  AOI210     o1659(.A0(ori_ori_n1515_), .A1(ori_ori_n975_), .B0(x0), .Y(ori_ori_n1709_));
  OAI210     o1660(.A0(ori_ori_n1708_), .A1(ori_ori_n1707_), .B0(ori_ori_n1709_), .Y(ori_ori_n1710_));
  NO3        o1661(.A(ori_ori_n1710_), .B(ori_ori_n1705_), .C(ori_ori_n1699_), .Y(ori_ori_n1711_));
  AOI210     o1662(.A0(x8), .A1(x6), .B0(x5), .Y(ori_ori_n1712_));
  AO220      o1663(.A0(ori_ori_n1712_), .A1(ori_ori_n135_), .B0(ori_ori_n541_), .B1(ori_ori_n132_), .Y(ori_ori_n1713_));
  NA2        o1664(.A(ori_ori_n1713_), .B(ori_ori_n405_), .Y(ori_ori_n1714_));
  NO2        o1665(.A(ori_ori_n688_), .B(ori_ori_n135_), .Y(ori_ori_n1715_));
  NA3        o1666(.A(ori_ori_n1715_), .B(ori_ori_n1537_), .C(ori_ori_n129_), .Y(ori_ori_n1716_));
  NO2        o1667(.A(ori_ori_n357_), .B(ori_ori_n1265_), .Y(ori_ori_n1717_));
  OAI210     o1668(.A0(ori_ori_n1717_), .A1(ori_ori_n1237_), .B0(ori_ori_n404_), .Y(ori_ori_n1718_));
  NA3        o1669(.A(ori_ori_n1718_), .B(ori_ori_n1716_), .C(ori_ori_n1714_), .Y(ori_ori_n1719_));
  INV        o1670(.A(ori_ori_n445_), .Y(ori_ori_n1720_));
  NO2        o1671(.A(ori_ori_n1720_), .B(ori_ori_n113_), .Y(ori_ori_n1721_));
  NA3        o1672(.A(ori_ori_n738_), .B(ori_ori_n928_), .C(x7), .Y(ori_ori_n1722_));
  AOI210     o1673(.A0(ori_ori_n314_), .A1(ori_ori_n198_), .B0(ori_ori_n1722_), .Y(ori_ori_n1723_));
  OAI220     o1674(.A0(ori_ori_n822_), .A1(ori_ori_n278_), .B0(ori_ori_n586_), .B1(ori_ori_n626_), .Y(ori_ori_n1724_));
  NO3        o1675(.A(ori_ori_n1724_), .B(ori_ori_n1723_), .C(ori_ori_n1721_), .Y(ori_ori_n1725_));
  OAI210     o1676(.A0(ori_ori_n1725_), .A1(ori_ori_n53_), .B0(x0), .Y(ori_ori_n1726_));
  AOI210     o1677(.A0(ori_ori_n1719_), .A1(x4), .B0(ori_ori_n1726_), .Y(ori_ori_n1727_));
  OA220      o1678(.A0(ori_ori_n1727_), .A1(ori_ori_n1711_), .B0(ori_ori_n1696_), .B1(ori_ori_n105_), .Y(ori27));
  NA2        o1679(.A(ori_ori_n1055_), .B(ori_ori_n404_), .Y(ori_ori_n1729_));
  NO2        o1680(.A(ori_ori_n1729_), .B(ori_ori_n273_), .Y(ori_ori_n1730_));
  NA2        o1681(.A(ori_ori_n837_), .B(ori_ori_n738_), .Y(ori_ori_n1731_));
  NA3        o1682(.A(ori_ori_n744_), .B(ori_ori_n331_), .C(ori_ori_n943_), .Y(ori_ori_n1732_));
  AOI210     o1683(.A0(ori_ori_n1732_), .A1(ori_ori_n1731_), .B0(ori_ori_n198_), .Y(ori_ori_n1733_));
  OAI210     o1684(.A0(ori_ori_n1733_), .A1(ori_ori_n1730_), .B0(ori_ori_n639_), .Y(ori_ori_n1734_));
  XO2        o1685(.A(x8), .B(x4), .Y(ori_ori_n1735_));
  NO2        o1686(.A(ori_ori_n1735_), .B(ori_ori_n157_), .Y(ori_ori_n1736_));
  OA210      o1687(.A0(ori_ori_n1736_), .A1(ori_ori_n1154_), .B0(ori_ori_n251_), .Y(ori_ori_n1737_));
  NA2        o1688(.A(ori_ori_n1737_), .B(ori_ori_n1034_), .Y(ori_ori_n1738_));
  AOI210     o1689(.A0(ori_ori_n578_), .A1(ori_ori_n56_), .B0(ori_ori_n1700_), .Y(ori_ori_n1739_));
  NO2        o1690(.A(ori_ori_n1739_), .B(ori_ori_n1153_), .Y(ori_ori_n1740_));
  NA2        o1691(.A(ori_ori_n1740_), .B(ori_ori_n489_), .Y(ori_ori_n1741_));
  NA3        o1692(.A(ori_ori_n1741_), .B(ori_ori_n1738_), .C(ori_ori_n1734_), .Y(ori28));
  NO3        o1693(.A(ori_ori_n1735_), .B(ori_ori_n1274_), .C(ori_ori_n137_), .Y(ori_ori_n1743_));
  OAI210     o1694(.A0(ori_ori_n1743_), .A1(ori_ori_n1171_), .B0(ori_ori_n533_), .Y(ori_ori_n1744_));
  NA3        o1695(.A(ori_ori_n1092_), .B(ori_ori_n816_), .C(x7), .Y(ori_ori_n1745_));
  NA3        o1696(.A(ori_ori_n447_), .B(ori_ori_n78_), .C(ori_ori_n555_), .Y(ori_ori_n1746_));
  NA3        o1697(.A(ori_ori_n1746_), .B(ori_ori_n1745_), .C(ori_ori_n1744_), .Y(ori_ori_n1747_));
  NA2        o1698(.A(ori_ori_n1150_), .B(ori_ori_n402_), .Y(ori_ori_n1748_));
  NA3        o1699(.A(ori_ori_n1748_), .B(ori_ori_n1289_), .C(ori_ori_n370_), .Y(ori_ori_n1749_));
  NO2        o1700(.A(ori_ori_n281_), .B(x4), .Y(ori_ori_n1750_));
  AOI220     o1701(.A0(ori_ori_n1750_), .A1(ori_ori_n1706_), .B0(ori_ori_n1035_), .B1(ori_ori_n616_), .Y(ori_ori_n1751_));
  NA2        o1702(.A(ori_ori_n1751_), .B(ori_ori_n1749_), .Y(ori_ori_n1752_));
  NO2        o1703(.A(ori_ori_n1150_), .B(ori_ori_n1129_), .Y(ori_ori_n1753_));
  NO4        o1704(.A(x6), .B(ori_ori_n56_), .C(x2), .D(x0), .Y(ori_ori_n1754_));
  OAI210     o1705(.A0(ori_ori_n1754_), .A1(ori_ori_n1753_), .B0(ori_ori_n964_), .Y(ori_ori_n1755_));
  NA2        o1706(.A(ori_ori_n1086_), .B(ori_ori_n104_), .Y(ori_ori_n1756_));
  NA2        o1707(.A(ori_ori_n997_), .B(ori_ori_n103_), .Y(ori_ori_n1757_));
  OAI210     o1708(.A0(ori_ori_n1757_), .A1(ori_ori_n1756_), .B0(ori_ori_n1755_), .Y(ori_ori_n1758_));
  OAI210     o1709(.A0(ori_ori_n1758_), .A1(ori_ori_n1752_), .B0(x7), .Y(ori_ori_n1759_));
  NO2        o1710(.A(ori_ori_n346_), .B(x7), .Y(ori_ori_n1760_));
  NO3        o1711(.A(ori_ori_n357_), .B(ori_ori_n246_), .C(ori_ori_n119_), .Y(ori_ori_n1761_));
  INV        o1712(.A(ori_ori_n81_), .Y(ori_ori_n1762_));
  OAI220     o1713(.A0(ori_ori_n1762_), .A1(ori_ori_n1761_), .B0(ori_ori_n1760_), .B1(ori_ori_n107_), .Y(ori_ori_n1763_));
  NA2        o1714(.A(ori_ori_n1649_), .B(ori_ori_n596_), .Y(ori_ori_n1764_));
  NO2        o1715(.A(ori_ori_n1688_), .B(ori_ori_n77_), .Y(ori_ori_n1765_));
  NA2        o1716(.A(ori_ori_n1765_), .B(ori_ori_n1764_), .Y(ori_ori_n1766_));
  AOI210     o1717(.A0(ori_ori_n1766_), .A1(ori_ori_n1763_), .B0(ori_ori_n59_), .Y(ori_ori_n1767_));
  NA2        o1718(.A(ori_ori_n369_), .B(ori_ori_n413_), .Y(ori_ori_n1768_));
  OAI210     o1719(.A0(ori_ori_n1768_), .A1(ori_ori_n134_), .B0(x1), .Y(ori_ori_n1769_));
  NO2        o1720(.A(ori_ori_n1769_), .B(ori_ori_n1767_), .Y(ori_ori_n1770_));
  AOI210     o1721(.A0(ori_ori_n1452_), .A1(ori_ori_n357_), .B0(ori_ori_n606_), .Y(ori_ori_n1771_));
  NO2        o1722(.A(ori_ori_n357_), .B(x5), .Y(ori_ori_n1772_));
  NO2        o1723(.A(ori_ori_n1772_), .B(ori_ori_n209_), .Y(ori_ori_n1773_));
  NO2        o1724(.A(ori_ori_n1773_), .B(ori_ori_n1771_), .Y(ori_ori_n1774_));
  NOi21      o1725(.An(ori_ori_n644_), .B(ori_ori_n918_), .Y(ori_ori_n1775_));
  NA2        o1726(.A(ori_ori_n1775_), .B(ori_ori_n997_), .Y(ori_ori_n1776_));
  INV        o1727(.A(ori_ori_n1776_), .Y(ori_ori_n1777_));
  OAI210     o1728(.A0(ori_ori_n1777_), .A1(ori_ori_n1774_), .B0(ori_ori_n1034_), .Y(ori_ori_n1778_));
  OAI210     o1729(.A0(ori_ori_n402_), .A1(ori_ori_n51_), .B0(ori_ori_n937_), .Y(ori_ori_n1779_));
  AOI220     o1730(.A0(ori_ori_n1779_), .A1(ori_ori_n417_), .B0(ori_ori_n402_), .B1(ori_ori_n347_), .Y(ori_ori_n1780_));
  NO2        o1731(.A(ori_ori_n1780_), .B(ori_ori_n142_), .Y(ori_ori_n1781_));
  NO2        o1732(.A(ori_ori_n276_), .B(x4), .Y(ori_ori_n1782_));
  NO2        o1733(.A(ori_ori_n644_), .B(ori_ori_n57_), .Y(ori_ori_n1783_));
  NA2        o1734(.A(ori_ori_n1783_), .B(ori_ori_n404_), .Y(ori_ori_n1784_));
  NA2        o1735(.A(ori_ori_n604_), .B(ori_ori_n670_), .Y(ori_ori_n1785_));
  AOI210     o1736(.A0(ori_ori_n1785_), .A1(ori_ori_n1784_), .B0(ori_ori_n233_), .Y(ori_ori_n1786_));
  NO3        o1737(.A(ori_ori_n1786_), .B(x1), .C(ori_ori_n1781_), .Y(ori_ori_n1787_));
  AOI220     o1738(.A0(ori_ori_n1787_), .A1(ori_ori_n1778_), .B0(ori_ori_n1770_), .B1(ori_ori_n1759_), .Y(ori_ori_n1788_));
  AOI210     o1739(.A0(ori_ori_n1747_), .A1(x3), .B0(ori_ori_n1788_), .Y(ori29));
  OAI210     o1740(.A0(ori_ori_n506_), .A1(ori_ori_n239_), .B0(ori_ori_n665_), .Y(ori_ori_n1790_));
  NA2        o1741(.A(ori_ori_n680_), .B(ori_ori_n964_), .Y(ori_ori_n1791_));
  AO210      o1742(.A0(ori_ori_n1067_), .A1(ori_ori_n1076_), .B0(ori_ori_n1791_), .Y(ori_ori_n1792_));
  NO2        o1743(.A(ori_ori_n168_), .B(ori_ori_n644_), .Y(ori_ori_n1793_));
  INV        o1744(.A(ori_ori_n1793_), .Y(ori_ori_n1794_));
  NA3        o1745(.A(ori_ori_n1794_), .B(ori_ori_n1792_), .C(ori_ori_n1790_), .Y(ori_ori_n1795_));
  NO2        o1746(.A(ori_ori_n1051_), .B(ori_ori_n50_), .Y(ori_ori_n1796_));
  NO3        o1747(.A(ori_ori_n1796_), .B(ori_ori_n1149_), .C(ori_ori_n506_), .Y(ori_ori_n1797_));
  NO2        o1748(.A(ori_ori_n400_), .B(ori_ori_n58_), .Y(ori_ori_n1798_));
  AOI220     o1749(.A0(ori_ori_n1798_), .A1(ori_ori_n1113_), .B0(ori_ori_n611_), .B1(ori_ori_n1264_), .Y(ori_ori_n1799_));
  OAI210     o1750(.A0(ori_ori_n1797_), .A1(ori_ori_n494_), .B0(ori_ori_n1799_), .Y(ori_ori_n1800_));
  AOI210     o1751(.A0(ori_ori_n1795_), .A1(x6), .B0(ori_ori_n1800_), .Y(ori_ori_n1801_));
  OAI210     o1752(.A0(x8), .A1(x4), .B0(x5), .Y(ori_ori_n1802_));
  NA2        o1753(.A(ori_ori_n1802_), .B(ori_ori_n108_), .Y(ori_ori_n1803_));
  NA2        o1754(.A(ori_ori_n276_), .B(ori_ori_n137_), .Y(ori_ori_n1804_));
  NA4        o1755(.A(ori_ori_n1804_), .B(ori_ori_n1803_), .C(ori_ori_n605_), .D(ori_ori_n64_), .Y(ori_ori_n1805_));
  AOI210     o1756(.A0(ori_ori_n1209_), .A1(ori_ori_n246_), .B0(ori_ori_n1590_), .Y(ori_ori_n1806_));
  AOI210     o1757(.A0(ori_ori_n1806_), .A1(ori_ori_n1805_), .B0(ori_ori_n809_), .Y(ori_ori_n1807_));
  NA4        o1758(.A(ori_ori_n606_), .B(ori_ori_n281_), .C(ori_ori_n168_), .D(ori_ori_n154_), .Y(ori_ori_n1808_));
  NA3        o1759(.A(ori_ori_n576_), .B(ori_ori_n269_), .C(ori_ori_n726_), .Y(ori_ori_n1809_));
  AOI210     o1760(.A0(ori_ori_n1809_), .A1(ori_ori_n1808_), .B0(ori_ori_n1113_), .Y(ori_ori_n1810_));
  OAI210     o1761(.A0(ori_ori_n816_), .A1(x8), .B0(x7), .Y(ori_ori_n1811_));
  NO2        o1762(.A(ori_ori_n1811_), .B(ori_ori_n123_), .Y(ori_ori_n1812_));
  OA210      o1763(.A0(ori_ori_n791_), .A1(ori_ori_n248_), .B0(ori_ori_n1802_), .Y(ori_ori_n1813_));
  OAI220     o1764(.A0(ori_ori_n1813_), .A1(ori_ori_n535_), .B0(ori_ori_n1378_), .B1(ori_ori_n353_), .Y(ori_ori_n1814_));
  NO4        o1765(.A(ori_ori_n1814_), .B(ori_ori_n1812_), .C(ori_ori_n1810_), .D(ori_ori_n1807_), .Y(ori_ori_n1815_));
  OAI210     o1766(.A0(ori_ori_n1801_), .A1(x2), .B0(ori_ori_n1815_), .Y(ori_ori_n1816_));
  NA3        o1767(.A(x6), .B(ori_ori_n50_), .C(x2), .Y(ori_ori_n1817_));
  NO2        o1768(.A(ori_ori_n1129_), .B(ori_ori_n322_), .Y(ori_ori_n1818_));
  NO2        o1769(.A(ori_ori_n402_), .B(x3), .Y(ori_ori_n1819_));
  AO220      o1770(.A0(ori_ori_n1819_), .A1(x5), .B0(ori_ori_n1754_), .B1(ori_ori_n81_), .Y(ori_ori_n1820_));
  AOI210     o1771(.A0(ori_ori_n1818_), .A1(ori_ori_n314_), .B0(ori_ori_n1820_), .Y(ori_ori_n1821_));
  NO3        o1772(.A(ori_ori_n637_), .B(ori_ori_n332_), .C(ori_ori_n133_), .Y(ori_ori_n1822_));
  AOI210     o1773(.A0(ori_ori_n664_), .A1(ori_ori_n561_), .B0(ori_ori_n1822_), .Y(ori_ori_n1823_));
  OAI210     o1774(.A0(ori_ori_n1821_), .A1(x7), .B0(ori_ori_n1823_), .Y(ori_ori_n1824_));
  AOI210     o1775(.A0(ori_ori_n1007_), .A1(ori_ori_n357_), .B0(ori_ori_n1288_), .Y(ori_ori_n1825_));
  AN2        o1776(.A(ori_ori_n575_), .B(ori_ori_n606_), .Y(ori_ori_n1826_));
  OAI210     o1777(.A0(ori_ori_n1826_), .A1(ori_ori_n1825_), .B0(ori_ori_n68_), .Y(ori_ori_n1827_));
  NO2        o1778(.A(ori_ori_n183_), .B(ori_ori_n85_), .Y(ori_ori_n1828_));
  OAI210     o1779(.A0(ori_ori_n1828_), .A1(ori_ori_n713_), .B0(ori_ori_n1013_), .Y(ori_ori_n1829_));
  NA3        o1780(.A(ori_ori_n1772_), .B(ori_ori_n212_), .C(ori_ori_n83_), .Y(ori_ori_n1830_));
  NA3        o1781(.A(ori_ori_n1830_), .B(ori_ori_n1829_), .C(ori_ori_n1827_), .Y(ori_ori_n1831_));
  AOI210     o1782(.A0(ori_ori_n1824_), .A1(x8), .B0(ori_ori_n1831_), .Y(ori_ori_n1832_));
  NO2        o1783(.A(ori_ori_n400_), .B(ori_ori_n224_), .Y(ori_ori_n1833_));
  OAI210     o1784(.A0(ori_ori_n1833_), .A1(ori_ori_n1035_), .B0(ori_ori_n616_), .Y(ori_ori_n1834_));
  NO3        o1785(.A(ori_ori_n941_), .B(ori_ori_n323_), .C(ori_ori_n138_), .Y(ori_ori_n1835_));
  NA3        o1786(.A(ori_ori_n1835_), .B(ori_ori_n1193_), .C(ori_ori_n50_), .Y(ori_ori_n1836_));
  NO2        o1787(.A(ori_ori_n129_), .B(ori_ori_n91_), .Y(ori_ori_n1837_));
  AOI220     o1788(.A0(ori_ori_n1837_), .A1(ori_ori_n536_), .B0(ori_ori_n1753_), .B1(ori_ori_n328_), .Y(ori_ori_n1838_));
  NOi31      o1789(.An(ori_ori_n1036_), .B(ori_ori_n1712_), .C(ori_ori_n570_), .Y(ori_ori_n1839_));
  NA2        o1790(.A(ori_ori_n159_), .B(x4), .Y(ori_ori_n1840_));
  NO3        o1791(.A(ori_ori_n1356_), .B(ori_ori_n220_), .C(ori_ori_n71_), .Y(ori_ori_n1841_));
  AOI210     o1792(.A0(ori_ori_n1841_), .A1(ori_ori_n1840_), .B0(ori_ori_n1839_), .Y(ori_ori_n1842_));
  NA4        o1793(.A(ori_ori_n1842_), .B(ori_ori_n1838_), .C(ori_ori_n1836_), .D(ori_ori_n1834_), .Y(ori_ori_n1843_));
  NO4        o1794(.A(ori_ori_n1129_), .B(ori_ori_n157_), .C(ori_ori_n55_), .D(ori_ori_n71_), .Y(ori_ori_n1844_));
  NO4        o1795(.A(ori_ori_n1106_), .B(ori_ori_n454_), .C(ori_ori_n1264_), .D(ori_ori_n104_), .Y(ori_ori_n1845_));
  OAI210     o1796(.A0(ori_ori_n1845_), .A1(ori_ori_n1844_), .B0(ori_ori_n106_), .Y(ori_ori_n1846_));
  AOI210     o1797(.A0(ori_ori_n280_), .A1(x4), .B0(ori_ori_n177_), .Y(ori_ori_n1847_));
  OAI210     o1798(.A0(ori_ori_n1847_), .A1(ori_ori_n1798_), .B0(ori_ori_n661_), .Y(ori_ori_n1848_));
  OR3        o1799(.A(ori_ori_n1611_), .B(ori_ori_n1310_), .C(ori_ori_n999_), .Y(ori_ori_n1849_));
  NA2        o1800(.A(ori_ori_n1754_), .B(ori_ori_n733_), .Y(ori_ori_n1850_));
  OR2        o1801(.A(ori_ori_n1850_), .B(ori_ori_n224_), .Y(ori_ori_n1851_));
  NA4        o1802(.A(ori_ori_n1851_), .B(ori_ori_n1849_), .C(ori_ori_n1848_), .D(ori_ori_n1846_), .Y(ori_ori_n1852_));
  AOI210     o1803(.A0(ori_ori_n1843_), .A1(ori_ori_n265_), .B0(ori_ori_n1852_), .Y(ori_ori_n1853_));
  OAI210     o1804(.A0(ori_ori_n1832_), .A1(x1), .B0(ori_ori_n1853_), .Y(ori_ori_n1854_));
  AO210      o1805(.A0(ori_ori_n1816_), .A1(x1), .B0(ori_ori_n1854_), .Y(ori30));
  NO3        o1806(.A(ori_ori_n1634_), .B(ori_ori_n524_), .C(ori_ori_n95_), .Y(ori_ori_n1856_));
  NO3        o1807(.A(ori_ori_n1049_), .B(ori_ori_n130_), .C(ori_ori_n343_), .Y(ori_ori_n1857_));
  AOI210     o1808(.A0(ori_ori_n661_), .A1(ori_ori_n230_), .B0(ori_ori_n1857_), .Y(ori_ori_n1858_));
  AOI210     o1809(.A0(ori_ori_n1858_), .A1(ori_ori_n1856_), .B0(ori_ori_n56_), .Y(ori_ori_n1859_));
  NA2        o1810(.A(ori_ori_n738_), .B(ori_ori_n312_), .Y(ori_ori_n1860_));
  NA2        o1811(.A(ori_ori_n1860_), .B(ori_ori_n1249_), .Y(ori_ori_n1861_));
  OAI210     o1812(.A0(ori_ori_n1861_), .A1(ori_ori_n1859_), .B0(ori_ori_n106_), .Y(ori_ori_n1862_));
  OAI210     o1813(.A0(ori_ori_n918_), .A1(ori_ori_n518_), .B0(ori_ori_n616_), .Y(ori_ori_n1863_));
  AOI220     o1814(.A0(ori_ori_n405_), .A1(ori_ori_n858_), .B0(ori_ori_n299_), .B1(ori_ori_n413_), .Y(ori_ori_n1864_));
  AOI210     o1815(.A0(ori_ori_n1864_), .A1(ori_ori_n1863_), .B0(ori_ori_n233_), .Y(ori_ori_n1865_));
  NO3        o1816(.A(ori_ori_n254_), .B(ori_ori_n120_), .C(x0), .Y(ori_ori_n1866_));
  AOI210     o1817(.A0(ori_ori_n456_), .A1(x6), .B0(ori_ori_n1866_), .Y(ori_ori_n1867_));
  AOI220     o1818(.A0(ori_ori_n1045_), .A1(ori_ori_n381_), .B0(ori_ori_n691_), .B1(ori_ori_n90_), .Y(ori_ori_n1868_));
  OAI220     o1819(.A0(ori_ori_n1868_), .A1(ori_ori_n224_), .B0(ori_ori_n1867_), .B1(ori_ori_n54_), .Y(ori_ori_n1869_));
  NA2        o1820(.A(ori_ori_n152_), .B(ori_ori_n71_), .Y(ori_ori_n1870_));
  AO210      o1821(.A0(ori_ori_n517_), .A1(ori_ori_n470_), .B0(x5), .Y(ori_ori_n1871_));
  AOI210     o1822(.A0(ori_ori_n1870_), .A1(ori_ori_n659_), .B0(ori_ori_n1871_), .Y(ori_ori_n1872_));
  AOI210     o1823(.A0(ori_ori_n1473_), .A1(ori_ori_n50_), .B0(ori_ori_n413_), .Y(ori_ori_n1873_));
  NA2        o1824(.A(ori_ori_n182_), .B(x2), .Y(ori_ori_n1874_));
  OR2        o1825(.A(ori_ori_n1874_), .B(ori_ori_n1873_), .Y(ori_ori_n1875_));
  OAI210     o1826(.A0(x7), .A1(x6), .B0(x1), .Y(ori_ori_n1876_));
  NA3        o1827(.A(ori_ori_n57_), .B(x4), .C(ori_ori_n59_), .Y(ori_ori_n1877_));
  AOI220     o1828(.A0(ori_ori_n1877_), .A1(ori_ori_n1254_), .B0(ori_ori_n1876_), .B1(ori_ori_n1669_), .Y(ori_ori_n1878_));
  NO3        o1829(.A(ori_ori_n1250_), .B(ori_ori_n314_), .C(ori_ori_n943_), .Y(ori_ori_n1879_));
  NO2        o1830(.A(ori_ori_n468_), .B(ori_ori_n784_), .Y(ori_ori_n1880_));
  NOi21      o1831(.An(ori_ori_n1880_), .B(ori_ori_n769_), .Y(ori_ori_n1881_));
  NO3        o1832(.A(ori_ori_n1193_), .B(ori_ori_n213_), .C(ori_ori_n588_), .Y(ori_ori_n1882_));
  NO4        o1833(.A(ori_ori_n1882_), .B(ori_ori_n1881_), .C(ori_ori_n1879_), .D(ori_ori_n1878_), .Y(ori_ori_n1883_));
  OAI210     o1834(.A0(ori_ori_n1875_), .A1(ori_ori_n687_), .B0(ori_ori_n1883_), .Y(ori_ori_n1884_));
  NO4        o1835(.A(ori_ori_n1884_), .B(ori_ori_n1872_), .C(ori_ori_n1869_), .D(ori_ori_n1865_), .Y(ori_ori_n1885_));
  AOI210     o1836(.A0(ori_ori_n1885_), .A1(ori_ori_n1862_), .B0(x8), .Y(ori_ori_n1886_));
  NO3        o1837(.A(ori_ori_n443_), .B(ori_ori_n710_), .C(ori_ori_n53_), .Y(ori_ori_n1887_));
  OAI220     o1838(.A0(ori_ori_n1647_), .A1(ori_ori_n314_), .B0(ori_ori_n435_), .B1(ori_ori_n532_), .Y(ori_ori_n1888_));
  OAI210     o1839(.A0(ori_ori_n1888_), .A1(ori_ori_n1887_), .B0(x6), .Y(ori_ori_n1889_));
  OAI210     o1840(.A0(ori_ori_n957_), .A1(ori_ori_n489_), .B0(ori_ori_n738_), .Y(ori_ori_n1890_));
  OAI210     o1841(.A0(ori_ori_n1600_), .A1(ori_ori_n302_), .B0(ori_ori_n122_), .Y(ori_ori_n1891_));
  AOI210     o1842(.A0(ori_ori_n340_), .A1(ori_ori_n211_), .B0(ori_ori_n72_), .Y(ori_ori_n1892_));
  INV        o1843(.A(ori_ori_n1892_), .Y(ori_ori_n1893_));
  NA4        o1844(.A(ori_ori_n1893_), .B(ori_ori_n1891_), .C(ori_ori_n1890_), .D(ori_ori_n1889_), .Y(ori_ori_n1894_));
  NA2        o1845(.A(ori_ori_n1004_), .B(ori_ori_n59_), .Y(ori_ori_n1895_));
  AOI210     o1846(.A0(ori_ori_n841_), .A1(ori_ori_n444_), .B0(ori_ori_n622_), .Y(ori_ori_n1896_));
  OAI220     o1847(.A0(ori_ori_n1896_), .A1(ori_ori_n280_), .B0(ori_ori_n1895_), .B1(ori_ori_n434_), .Y(ori_ori_n1897_));
  AOI210     o1848(.A0(ori_ori_n1894_), .A1(x8), .B0(ori_ori_n1897_), .Y(ori_ori_n1898_));
  NO2        o1849(.A(ori_ori_n1898_), .B(ori_ori_n57_), .Y(ori_ori_n1899_));
  INV        o1850(.A(ori_ori_n392_), .Y(ori_ori_n1900_));
  INV        o1851(.A(ori_ori_n602_), .Y(ori_ori_n1901_));
  AOI210     o1852(.A0(ori_ori_n1901_), .A1(ori_ori_n1900_), .B0(ori_ori_n402_), .Y(ori_ori_n1902_));
  NO3        o1853(.A(ori_ori_n580_), .B(ori_ori_n366_), .C(ori_ori_n1049_), .Y(ori_ori_n1903_));
  NO2        o1854(.A(ori_ori_n1903_), .B(ori_ori_n1153_), .Y(ori_ori_n1904_));
  NA2        o1855(.A(ori_ori_n277_), .B(x1), .Y(ori_ori_n1905_));
  NO2        o1856(.A(ori_ori_n283_), .B(x5), .Y(ori_ori_n1906_));
  NO2        o1857(.A(ori_ori_n1906_), .B(ori_ori_n777_), .Y(ori_ori_n1907_));
  OAI220     o1858(.A0(ori_ori_n1907_), .A1(ori_ori_n972_), .B0(ori_ori_n1905_), .B1(ori_ori_n190_), .Y(ori_ori_n1908_));
  NO3        o1859(.A(ori_ori_n1908_), .B(ori_ori_n1904_), .C(ori_ori_n1902_), .Y(ori_ori_n1909_));
  NA2        o1860(.A(ori_ori_n879_), .B(ori_ori_n82_), .Y(ori_ori_n1910_));
  OR2        o1861(.A(ori_ori_n1474_), .B(x3), .Y(ori_ori_n1911_));
  NO2        o1862(.A(ori_ori_n200_), .B(ori_ori_n56_), .Y(ori_ori_n1912_));
  NO2        o1863(.A(ori_ori_n323_), .B(ori_ori_n213_), .Y(ori_ori_n1913_));
  AOI220     o1864(.A0(ori_ori_n1913_), .A1(x2), .B0(ori_ori_n1912_), .B1(ori_ori_n1488_), .Y(ori_ori_n1914_));
  AOI210     o1865(.A0(ori_ori_n1914_), .A1(ori_ori_n1911_), .B0(ori_ori_n238_), .Y(ori_ori_n1915_));
  NO2        o1866(.A(ori_ori_n277_), .B(ori_ori_n119_), .Y(ori_ori_n1916_));
  NO3        o1867(.A(ori_ori_n743_), .B(ori_ori_n638_), .C(ori_ori_n154_), .Y(ori_ori_n1917_));
  OAI210     o1868(.A0(ori_ori_n1917_), .A1(ori_ori_n1916_), .B0(ori_ori_n143_), .Y(ori_ori_n1918_));
  NA2        o1869(.A(x4), .B(ori_ori_n59_), .Y(ori_ori_n1919_));
  AOI210     o1870(.A0(ori_ori_n1919_), .A1(ori_ori_n1199_), .B0(ori_ori_n490_), .Y(ori_ori_n1920_));
  AOI210     o1871(.A0(ori_ori_n1217_), .A1(x2), .B0(ori_ori_n1920_), .Y(ori_ori_n1921_));
  AOI210     o1872(.A0(ori_ori_n1921_), .A1(ori_ori_n1918_), .B0(ori_ori_n50_), .Y(ori_ori_n1922_));
  NA3        o1873(.A(ori_ori_n1353_), .B(ori_ori_n1043_), .C(ori_ori_n431_), .Y(ori_ori_n1923_));
  AOI210     o1874(.A0(ori_ori_n1923_), .A1(ori_ori_n1910_), .B0(ori_ori_n558_), .Y(ori_ori_n1924_));
  AOI210     o1875(.A0(ori_ori_n943_), .A1(x1), .B0(ori_ori_n1209_), .Y(ori_ori_n1925_));
  OAI220     o1876(.A0(ori_ori_n281_), .A1(x4), .B0(ori_ori_n51_), .B1(x6), .Y(ori_ori_n1926_));
  NO2        o1877(.A(ori_ori_n118_), .B(ori_ori_n108_), .Y(ori_ori_n1927_));
  AOI220     o1878(.A0(ori_ori_n1927_), .A1(ori_ori_n1926_), .B0(ori_ori_n1069_), .B1(ori_ori_n570_), .Y(ori_ori_n1928_));
  OAI210     o1879(.A0(ori_ori_n1925_), .A1(ori_ori_n438_), .B0(ori_ori_n1928_), .Y(ori_ori_n1929_));
  NO4        o1880(.A(ori_ori_n1929_), .B(ori_ori_n1924_), .C(ori_ori_n1922_), .D(ori_ori_n1915_), .Y(ori_ori_n1930_));
  OAI210     o1881(.A0(ori_ori_n1909_), .A1(ori_ori_n129_), .B0(ori_ori_n1930_), .Y(ori_ori_n1931_));
  NO3        o1882(.A(ori_ori_n1931_), .B(ori_ori_n1899_), .C(ori_ori_n1886_), .Y(ori31));
  INV        o1883(.A(ori_ori_n324_), .Y(ori_ori_n1933_));
  NO2        o1884(.A(ori_ori_n406_), .B(ori_ori_n616_), .Y(ori_ori_n1934_));
  AOI210     o1885(.A0(ori_ori_n1934_), .A1(ori_ori_n1933_), .B0(ori_ori_n58_), .Y(ori_ori_n1935_));
  NO2        o1886(.A(ori_ori_n712_), .B(ori_ori_n56_), .Y(ori_ori_n1936_));
  AOI220     o1887(.A0(ori_ori_n1936_), .A1(x2), .B0(ori_ori_n89_), .B1(x0), .Y(ori_ori_n1937_));
  NA3        o1888(.A(ori_ori_n1937_), .B(ori_ori_n1850_), .C(ori_ori_n1697_), .Y(ori_ori_n1938_));
  OAI210     o1889(.A0(ori_ori_n1938_), .A1(ori_ori_n1935_), .B0(ori_ori_n53_), .Y(ori_ori_n1939_));
  INV        o1890(.A(ori_ori_n616_), .Y(ori_ori_n1940_));
  NO2        o1891(.A(ori_ori_n1782_), .B(ori_ori_n810_), .Y(ori_ori_n1941_));
  OA220      o1892(.A0(ori_ori_n1941_), .A1(ori_ori_n431_), .B0(ori_ori_n1940_), .B1(ori_ori_n1347_), .Y(ori_ori_n1942_));
  AOI210     o1893(.A0(ori_ori_n1942_), .A1(ori_ori_n1939_), .B0(ori_ori_n104_), .Y(ori_ori_n1943_));
  NO2        o1894(.A(ori_ori_n450_), .B(ori_ori_n75_), .Y(ori_ori_n1944_));
  NA2        o1895(.A(ori_ori_n402_), .B(ori_ori_n57_), .Y(ori_ori_n1945_));
  AOI210     o1896(.A0(ori_ori_n280_), .A1(ori_ori_n86_), .B0(ori_ori_n1945_), .Y(ori_ori_n1946_));
  OAI210     o1897(.A0(ori_ori_n1946_), .A1(ori_ori_n1944_), .B0(ori_ori_n699_), .Y(ori_ori_n1947_));
  NO4        o1898(.A(ori_ori_n1065_), .B(ori_ori_n332_), .C(ori_ori_n1473_), .D(ori_ori_n67_), .Y(ori_ori_n1948_));
  AOI210     o1899(.A0(ori_ori_n1510_), .A1(ori_ori_n1244_), .B0(ori_ori_n400_), .Y(ori_ori_n1949_));
  NO2        o1900(.A(ori_ori_n1200_), .B(ori_ori_n872_), .Y(ori_ori_n1950_));
  NO3        o1901(.A(ori_ori_n1950_), .B(ori_ori_n1949_), .C(ori_ori_n1948_), .Y(ori_ori_n1951_));
  AOI210     o1902(.A0(ori_ori_n1951_), .A1(ori_ori_n1947_), .B0(x5), .Y(ori_ori_n1952_));
  AOI220     o1903(.A0(ori_ori_n404_), .A1(ori_ori_n570_), .B0(ori_ori_n518_), .B1(ori_ori_n63_), .Y(ori_ori_n1953_));
  AOI210     o1904(.A0(ori_ori_n1953_), .A1(ori_ori_n528_), .B0(ori_ori_n1129_), .Y(ori_ori_n1954_));
  AOI220     o1905(.A0(ori_ori_n880_), .A1(ori_ori_n670_), .B0(ori_ori_n1049_), .B1(ori_ori_n117_), .Y(ori_ori_n1955_));
  OAI220     o1906(.A0(ori_ori_n1955_), .A1(ori_ori_n346_), .B0(ori_ori_n434_), .B1(ori_ori_n700_), .Y(ori_ori_n1956_));
  NO4        o1907(.A(ori_ori_n1956_), .B(ori_ori_n1954_), .C(ori_ori_n1952_), .D(ori_ori_n1943_), .Y(ori_ori_n1957_));
  NA2        o1908(.A(ori_ori_n444_), .B(ori_ori_n59_), .Y(ori_ori_n1958_));
  AOI210     o1909(.A0(ori_ori_n494_), .A1(ori_ori_n1958_), .B0(ori_ori_n132_), .Y(ori_ori_n1959_));
  OAI210     o1910(.A0(ori_ori_n100_), .A1(ori_ori_n248_), .B0(ori_ori_n1895_), .Y(ori_ori_n1960_));
  OAI210     o1911(.A0(ori_ori_n1960_), .A1(ori_ori_n1959_), .B0(x7), .Y(ori_ori_n1961_));
  NA2        o1912(.A(ori_ori_n1001_), .B(ori_ori_n90_), .Y(ori_ori_n1962_));
  AOI210     o1913(.A0(ori_ori_n822_), .A1(ori_ori_n108_), .B0(ori_ori_n1962_), .Y(ori_ori_n1963_));
  NA2        o1914(.A(ori_ori_n1421_), .B(x6), .Y(ori_ori_n1964_));
  AOI210     o1915(.A0(ori_ori_n1964_), .A1(ori_ori_n264_), .B0(ori_ori_n104_), .Y(ori_ori_n1965_));
  NA2        o1916(.A(ori_ori_n1092_), .B(ori_ori_n291_), .Y(ori_ori_n1966_));
  AOI210     o1917(.A0(ori_ori_n1966_), .A1(ori_ori_n586_), .B0(ori_ori_n53_), .Y(ori_ori_n1967_));
  NO3        o1918(.A(ori_ori_n1967_), .B(ori_ori_n1965_), .C(ori_ori_n1963_), .Y(ori_ori_n1968_));
  AOI210     o1919(.A0(ori_ori_n1968_), .A1(ori_ori_n1961_), .B0(ori_ori_n626_), .Y(ori_ori_n1969_));
  NOi21      o1920(.An(ori_ori_n1625_), .B(ori_ori_n976_), .Y(ori_ori_n1970_));
  OAI220     o1921(.A0(ori_ori_n1970_), .A1(ori_ori_n1756_), .B0(ori_ori_n842_), .B1(ori_ori_n1958_), .Y(ori_ori_n1971_));
  NA2        o1922(.A(ori_ori_n1971_), .B(x3), .Y(ori_ori_n1972_));
  AOI220     o1923(.A0(ori_ori_n1274_), .A1(x8), .B0(ori_ori_n60_), .B1(x1), .Y(ori_ori_n1973_));
  NO3        o1924(.A(ori_ori_n1973_), .B(ori_ori_n1024_), .C(x6), .Y(ori_ori_n1974_));
  NA2        o1925(.A(ori_ori_n561_), .B(ori_ori_n366_), .Y(ori_ori_n1975_));
  NA2        o1926(.A(ori_ori_n114_), .B(ori_ori_n481_), .Y(ori_ori_n1976_));
  OAI220     o1927(.A0(ori_ori_n1976_), .A1(ori_ori_n1756_), .B0(ori_ori_n1975_), .B1(x4), .Y(ori_ori_n1977_));
  NO2        o1928(.A(ori_ori_n1977_), .B(ori_ori_n1974_), .Y(ori_ori_n1978_));
  AOI210     o1929(.A0(ori_ori_n1978_), .A1(ori_ori_n1972_), .B0(ori_ori_n170_), .Y(ori_ori_n1979_));
  NO4        o1930(.A(ori_ori_n562_), .B(ori_ori_n536_), .C(ori_ori_n639_), .D(ori_ori_n638_), .Y(ori_ori_n1980_));
  OAI210     o1931(.A0(ori_ori_n1980_), .A1(ori_ori_n992_), .B0(x3), .Y(ori_ori_n1981_));
  NO4        o1932(.A(ori_ori_n729_), .B(ori_ori_n1129_), .C(ori_ori_n699_), .D(x5), .Y(ori_ori_n1982_));
  NO3        o1933(.A(x6), .B(ori_ori_n56_), .C(x1), .Y(ori_ori_n1983_));
  NO2        o1934(.A(ori_ori_n1729_), .B(ori_ori_n340_), .Y(ori_ori_n1984_));
  NA4        o1935(.A(ori_ori_n580_), .B(ori_ori_n164_), .C(x6), .D(ori_ori_n104_), .Y(ori_ori_n1985_));
  NO2        o1936(.A(ori_ori_n778_), .B(ori_ori_n227_), .Y(ori_ori_n1986_));
  NOi41      o1937(.An(ori_ori_n1985_), .B(ori_ori_n1986_), .C(ori_ori_n1984_), .D(ori_ori_n1982_), .Y(ori_ori_n1987_));
  AOI210     o1938(.A0(ori_ori_n1987_), .A1(ori_ori_n1981_), .B0(ori_ori_n485_), .Y(ori_ori_n1988_));
  OAI210     o1939(.A0(ori_ori_n561_), .A1(ori_ori_n425_), .B0(ori_ori_n858_), .Y(ori_ori_n1989_));
  NO3        o1940(.A(ori_ori_n336_), .B(ori_ori_n77_), .C(ori_ori_n53_), .Y(ori_ori_n1990_));
  NO3        o1941(.A(ori_ori_n417_), .B(ori_ori_n318_), .C(ori_ori_n50_), .Y(ori_ori_n1991_));
  OAI210     o1942(.A0(ori_ori_n1991_), .A1(ori_ori_n1990_), .B0(ori_ori_n1066_), .Y(ori_ori_n1992_));
  AOI210     o1943(.A0(ori_ori_n1992_), .A1(ori_ori_n1989_), .B0(ori_ori_n351_), .Y(ori_ori_n1993_));
  NO2        o1944(.A(ori_ori_n198_), .B(ori_ori_n490_), .Y(ori_ori_n1994_));
  OAI210     o1945(.A0(ori_ori_n130_), .A1(x2), .B0(ori_ori_n1994_), .Y(ori_ori_n1995_));
  NO2        o1946(.A(ori_ori_n1995_), .B(ori_ori_n64_), .Y(ori_ori_n1996_));
  NA2        o1947(.A(ori_ori_n118_), .B(ori_ori_n57_), .Y(ori_ori_n1997_));
  AOI220     o1948(.A0(ori_ori_n1452_), .A1(ori_ori_n828_), .B0(ori_ori_n247_), .B1(x4), .Y(ori_ori_n1998_));
  AOI220     o1949(.A0(ori_ori_n1503_), .A1(ori_ori_n563_), .B0(ori_ori_n660_), .B1(ori_ori_n699_), .Y(ori_ori_n1999_));
  OAI220     o1950(.A0(ori_ori_n1999_), .A1(ori_ori_n1997_), .B0(ori_ori_n1998_), .B1(ori_ori_n175_), .Y(ori_ori_n2000_));
  OR3        o1951(.A(ori_ori_n2000_), .B(ori_ori_n1996_), .C(ori_ori_n1993_), .Y(ori_ori_n2001_));
  NO4        o1952(.A(ori_ori_n2001_), .B(ori_ori_n1988_), .C(ori_ori_n1979_), .D(ori_ori_n1969_), .Y(ori_ori_n2002_));
  OAI210     o1953(.A0(ori_ori_n1957_), .A1(x3), .B0(ori_ori_n2002_), .Y(ori32));
  OAI210     o1954(.A0(ori_ori_n514_), .A1(ori_ori_n53_), .B0(ori_ori_n371_), .Y(ori_ori_n2004_));
  NA2        o1955(.A(ori_ori_n465_), .B(x2), .Y(ori_ori_n2005_));
  AOI210     o1956(.A0(ori_ori_n2005_), .A1(ori_ori_n2004_), .B0(ori_ori_n57_), .Y(ori_ori_n2006_));
  OAI210     o1957(.A0(ori_ori_n2006_), .A1(ori_ori_n713_), .B0(ori_ori_n56_), .Y(ori_ori_n2007_));
  OAI210     o1958(.A0(ori_ori_n1571_), .A1(ori_ori_n1329_), .B0(ori_ori_n1355_), .Y(ori_ori_n2008_));
  AOI210     o1959(.A0(ori_ori_n1936_), .A1(ori_ori_n251_), .B0(ori_ori_n2008_), .Y(ori_ori_n2009_));
  AOI210     o1960(.A0(ori_ori_n2009_), .A1(ori_ori_n2007_), .B0(ori_ori_n50_), .Y(ori_ori_n2010_));
  NA3        o1961(.A(ori_ori_n1422_), .B(ori_ori_n727_), .C(ori_ori_n263_), .Y(ori_ori_n2011_));
  NA2        o1962(.A(ori_ori_n675_), .B(ori_ori_n498_), .Y(ori_ori_n2012_));
  OAI220     o1963(.A0(ori_ori_n971_), .A1(ori_ori_n212_), .B0(ori_ori_n623_), .B1(ori_ori_n190_), .Y(ori_ori_n2013_));
  NO3        o1964(.A(ori_ori_n337_), .B(ori_ori_n521_), .C(ori_ori_n733_), .Y(ori_ori_n2014_));
  NO2        o1965(.A(ori_ori_n1250_), .B(ori_ori_n532_), .Y(ori_ori_n2015_));
  NO4        o1966(.A(ori_ori_n2015_), .B(ori_ori_n2014_), .C(ori_ori_n2013_), .D(ori_ori_n2012_), .Y(ori_ori_n2016_));
  AOI210     o1967(.A0(ori_ori_n2016_), .A1(ori_ori_n2011_), .B0(ori_ori_n133_), .Y(ori_ori_n2017_));
  OAI220     o1968(.A0(ori_ori_n359_), .A1(x7), .B0(ori_ori_n276_), .B1(ori_ori_n269_), .Y(ori_ori_n2018_));
  NA2        o1969(.A(ori_ori_n2018_), .B(ori_ori_n879_), .Y(ori_ori_n2019_));
  NO2        o1970(.A(ori_ori_n501_), .B(ori_ori_n784_), .Y(ori_ori_n2020_));
  NA2        o1971(.A(ori_ori_n2020_), .B(ori_ori_n1715_), .Y(ori_ori_n2021_));
  AOI210     o1972(.A0(ori_ori_n2021_), .A1(ori_ori_n2019_), .B0(ori_ori_n106_), .Y(ori_ori_n2022_));
  NA2        o1973(.A(ori_ori_n1208_), .B(ori_ori_n1051_), .Y(ori_ori_n2023_));
  NA2        o1974(.A(ori_ori_n1245_), .B(ori_ori_n639_), .Y(ori_ori_n2024_));
  AOI210     o1975(.A0(ori_ori_n2024_), .A1(ori_ori_n2023_), .B0(ori_ori_n56_), .Y(ori_ori_n2025_));
  NA2        o1976(.A(ori_ori_n879_), .B(ori_ori_n57_), .Y(ori_ori_n2026_));
  NOi21      o1977(.An(ori_ori_n2026_), .B(ori_ori_n125_), .Y(ori_ori_n2027_));
  NA2        o1978(.A(ori_ori_n933_), .B(ori_ori_n227_), .Y(ori_ori_n2028_));
  NO3        o1979(.A(ori_ori_n2028_), .B(ori_ori_n2027_), .C(ori_ori_n59_), .Y(ori_ori_n2029_));
  OR4        o1980(.A(ori_ori_n2029_), .B(ori_ori_n2025_), .C(ori_ori_n2022_), .D(ori_ori_n2017_), .Y(ori_ori_n2030_));
  OAI210     o1981(.A0(ori_ori_n2030_), .A1(ori_ori_n2010_), .B0(ori_ori_n104_), .Y(ori_ori_n2031_));
  NO3        o1982(.A(ori_ori_n1129_), .B(ori_ori_n135_), .C(ori_ori_n121_), .Y(ori_ori_n2032_));
  NO2        o1983(.A(ori_ori_n341_), .B(ori_ori_n55_), .Y(ori_ori_n2033_));
  NA2        o1984(.A(ori_ori_n2033_), .B(ori_ori_n112_), .Y(ori_ori_n2034_));
  OAI210     o1985(.A0(ori_ori_n578_), .A1(ori_ori_n538_), .B0(ori_ori_n738_), .Y(ori_ori_n2035_));
  NA2        o1986(.A(ori_ori_n2035_), .B(ori_ori_n2034_), .Y(ori_ori_n2036_));
  OAI210     o1987(.A0(ori_ori_n2036_), .A1(ori_ori_n2032_), .B0(x3), .Y(ori_ori_n2037_));
  OAI210     o1988(.A0(ori_ori_n816_), .A1(ori_ori_n246_), .B0(ori_ori_n50_), .Y(ori_ori_n2038_));
  AOI210     o1989(.A0(ori_ori_n62_), .A1(ori_ori_n106_), .B0(ori_ori_n2038_), .Y(ori_ori_n2039_));
  OAI210     o1990(.A0(ori_ori_n2039_), .A1(ori_ori_n1700_), .B0(ori_ori_n638_), .Y(ori_ori_n2040_));
  NO3        o1991(.A(ori_ori_n278_), .B(ori_ori_n159_), .C(ori_ori_n119_), .Y(ori_ori_n2041_));
  NO3        o1992(.A(ori_ori_n727_), .B(ori_ori_n330_), .C(ori_ori_n133_), .Y(ori_ori_n2042_));
  OAI210     o1993(.A0(ori_ori_n2042_), .A1(ori_ori_n2041_), .B0(ori_ori_n59_), .Y(ori_ori_n2043_));
  NA2        o1994(.A(ori_ori_n1055_), .B(ori_ori_n71_), .Y(ori_ori_n2044_));
  NO2        o1995(.A(ori_ori_n1760_), .B(ori_ori_n538_), .Y(ori_ori_n2045_));
  AOI210     o1996(.A0(ori_ori_n2045_), .A1(ori_ori_n1701_), .B0(ori_ori_n2044_), .Y(ori_ori_n2046_));
  NO2        o1997(.A(ori_ori_n248_), .B(ori_ori_n57_), .Y(ori_ori_n2047_));
  NO2        o1998(.A(ori_ori_n2047_), .B(ori_ori_n925_), .Y(ori_ori_n2048_));
  NOi31      o1999(.An(ori_ori_n661_), .B(ori_ori_n2048_), .C(ori_ori_n254_), .Y(ori_ori_n2049_));
  NO3        o2000(.A(ori_ori_n2049_), .B(ori_ori_n2046_), .C(x1), .Y(ori_ori_n2050_));
  NA4        o2001(.A(ori_ori_n2050_), .B(ori_ori_n2043_), .C(ori_ori_n2040_), .D(ori_ori_n2037_), .Y(ori_ori_n2051_));
  AO210      o2002(.A0(ori_ori_n1007_), .A1(ori_ori_n354_), .B0(ori_ori_n928_), .Y(ori_ori_n2052_));
  NA3        o2003(.A(ori_ori_n1735_), .B(ori_ori_n505_), .C(ori_ori_n248_), .Y(ori_ori_n2053_));
  AOI210     o2004(.A0(ori_ori_n2053_), .A1(ori_ori_n2052_), .B0(ori_ori_n278_), .Y(ori_ori_n2054_));
  NA3        o2005(.A(ori_ori_n1161_), .B(ori_ori_n479_), .C(ori_ori_n212_), .Y(ori_ori_n2055_));
  NO3        o2006(.A(ori_ori_n1310_), .B(ori_ori_n928_), .C(x2), .Y(ori_ori_n2056_));
  NO2        o2007(.A(ori_ori_n1685_), .B(ori_ori_n64_), .Y(ori_ori_n2057_));
  NO3        o2008(.A(ori_ori_n2057_), .B(ori_ori_n2056_), .C(ori_ori_n53_), .Y(ori_ori_n2058_));
  NO3        o2009(.A(ori_ori_n421_), .B(ori_ori_n1001_), .C(ori_ori_n118_), .Y(ori_ori_n2059_));
  OAI220     o2010(.A0(ori_ori_n626_), .A1(ori_ori_n159_), .B0(ori_ori_n323_), .B1(ori_ori_n133_), .Y(ori_ori_n2060_));
  OAI210     o2011(.A0(ori_ori_n2060_), .A1(ori_ori_n2059_), .B0(ori_ori_n68_), .Y(ori_ori_n2061_));
  NO2        o2012(.A(ori_ori_n1802_), .B(ori_ori_n333_), .Y(ori_ori_n2062_));
  OAI210     o2013(.A0(ori_ori_n1703_), .A1(ori_ori_n556_), .B0(ori_ori_n2062_), .Y(ori_ori_n2063_));
  NA4        o2014(.A(ori_ori_n2063_), .B(ori_ori_n2061_), .C(ori_ori_n2058_), .D(ori_ori_n2055_), .Y(ori_ori_n2064_));
  OAI210     o2015(.A0(ori_ori_n2064_), .A1(ori_ori_n2054_), .B0(ori_ori_n2051_), .Y(ori_ori_n2065_));
  NO3        o2016(.A(ori_ori_n1119_), .B(ori_ori_n103_), .C(ori_ori_n71_), .Y(ori_ori_n2066_));
  NO2        o2017(.A(ori_ori_n514_), .B(ori_ori_n335_), .Y(ori_ori_n2067_));
  OAI210     o2018(.A0(ori_ori_n2066_), .A1(ori_ori_n1294_), .B0(ori_ori_n2067_), .Y(ori_ori_n2068_));
  NO3        o2019(.A(x8), .B(ori_ori_n71_), .C(x2), .Y(ori_ori_n2069_));
  OAI220     o2020(.A0(ori_ori_n2069_), .A1(ori_ori_n570_), .B0(ori_ori_n1302_), .B1(ori_ori_n89_), .Y(ori_ori_n2070_));
  AOI220     o2021(.A0(ori_ori_n506_), .A1(ori_ori_n738_), .B0(ori_ori_n616_), .B1(ori_ori_n231_), .Y(ori_ori_n2071_));
  AOI210     o2022(.A0(ori_ori_n2071_), .A1(ori_ori_n2070_), .B0(ori_ori_n241_), .Y(ori_ori_n2072_));
  NA2        o2023(.A(ori_ori_n933_), .B(ori_ori_n1049_), .Y(ori_ori_n2073_));
  AOI210     o2024(.A0(ori_ori_n612_), .A1(ori_ori_n626_), .B0(ori_ori_n2073_), .Y(ori_ori_n2074_));
  AOI210     o2025(.A0(ori_ori_n536_), .A1(ori_ori_n570_), .B0(ori_ori_n632_), .Y(ori_ori_n2075_));
  NO2        o2026(.A(ori_ori_n2075_), .B(ori_ori_n1669_), .Y(ori_ori_n2076_));
  INV        o2027(.A(ori_ori_n407_), .Y(ori_ori_n2077_));
  NOi31      o2028(.An(ori_ori_n1370_), .B(ori_ori_n2077_), .C(ori_ori_n536_), .Y(ori_ori_n2078_));
  NO4        o2029(.A(ori_ori_n2078_), .B(ori_ori_n2076_), .C(ori_ori_n2074_), .D(ori_ori_n2072_), .Y(ori_ori_n2079_));
  NA4        o2030(.A(ori_ori_n2079_), .B(ori_ori_n2068_), .C(ori_ori_n2065_), .D(ori_ori_n2031_), .Y(ori33));
  NA2        o2031(.A(x1), .B(ori_ori_n185_), .Y(ori_ori_n2081_));
  OAI210     o2032(.A0(ori_ori_n1906_), .A1(ori_ori_n163_), .B0(ori_ori_n300_), .Y(ori_ori_n2082_));
  OAI220     o2033(.A0(ori_ori_n989_), .A1(ori_ori_n733_), .B0(ori_ori_n1537_), .B1(ori_ori_n322_), .Y(ori_ori_n2083_));
  NA3        o2034(.A(ori_ori_n2083_), .B(ori_ori_n2082_), .C(ori_ori_n579_), .Y(ori_ori_n2084_));
  AOI210     o2035(.A0(ori_ori_n2081_), .A1(x5), .B0(ori_ori_n2084_), .Y(ori_ori_n2085_));
  NA2        o2036(.A(ori_ori_n211_), .B(ori_ori_n76_), .Y(ori_ori_n2086_));
  NO2        o2037(.A(ori_ori_n2086_), .B(ori_ori_n322_), .Y(ori_ori_n2087_));
  OAI210     o2038(.A0(ori_ori_n392_), .A1(ori_ori_n244_), .B0(ori_ori_n53_), .Y(ori_ori_n2088_));
  AOI210     o2039(.A0(ori_ori_n2088_), .A1(ori_ori_n394_), .B0(ori_ori_n64_), .Y(ori_ori_n2089_));
  NO3        o2040(.A(x6), .B(ori_ori_n2089_), .C(ori_ori_n2087_), .Y(ori_ori_n2090_));
  OAI210     o2041(.A0(ori_ori_n2085_), .A1(x4), .B0(ori_ori_n2090_), .Y(ori_ori_n2091_));
  INV        o2042(.A(ori_ori_n219_), .Y(ori_ori_n2092_));
  NA2        o2043(.A(ori_ori_n170_), .B(x4), .Y(ori_ori_n2093_));
  NA2        o2044(.A(ori_ori_n283_), .B(ori_ori_n260_), .Y(ori_ori_n2094_));
  NO2        o2045(.A(ori_ori_n879_), .B(ori_ori_n209_), .Y(ori_ori_n2095_));
  NA2        o2046(.A(ori_ori_n581_), .B(x7), .Y(ori_ori_n2096_));
  OAI220     o2047(.A0(ori_ori_n2096_), .A1(ori_ori_n2095_), .B0(ori_ori_n2094_), .B1(ori_ori_n2093_), .Y(ori_ori_n2097_));
  AOI210     o2048(.A0(ori_ori_n2092_), .A1(ori_ori_n941_), .B0(ori_ori_n2097_), .Y(ori_ori_n2098_));
  NA2        o2049(.A(ori_ori_n194_), .B(ori_ori_n871_), .Y(ori_ori_n2099_));
  AOI210     o2050(.A0(ori_ori_n2099_), .A1(ori_ori_n2026_), .B0(ori_ori_n196_), .Y(ori_ori_n2100_));
  OAI210     o2051(.A0(ori_ori_n784_), .A1(ori_ori_n51_), .B0(x6), .Y(ori_ori_n2101_));
  NA3        o2052(.A(ori_ori_n837_), .B(ori_ori_n665_), .C(ori_ori_n55_), .Y(ori_ori_n2102_));
  OAI210     o2053(.A0(ori_ori_n565_), .A1(ori_ori_n456_), .B0(ori_ori_n2102_), .Y(ori_ori_n2103_));
  NO3        o2054(.A(ori_ori_n2103_), .B(ori_ori_n2101_), .C(ori_ori_n2100_), .Y(ori_ori_n2104_));
  OAI210     o2055(.A0(ori_ori_n2098_), .A1(ori_ori_n50_), .B0(ori_ori_n2104_), .Y(ori_ori_n2105_));
  NA3        o2056(.A(ori_ori_n2105_), .B(ori_ori_n2091_), .C(ori_ori_n59_), .Y(ori_ori_n2106_));
  NO3        o2057(.A(ori_ori_n1434_), .B(ori_ori_n336_), .C(x4), .Y(ori_ori_n2107_));
  NA2        o2058(.A(ori_ori_n2107_), .B(ori_ori_n129_), .Y(ori_ori_n2108_));
  NA2        o2059(.A(ori_ori_n736_), .B(ori_ori_n104_), .Y(ori_ori_n2109_));
  NO2        o2060(.A(ori_ori_n644_), .B(ori_ori_n337_), .Y(ori_ori_n2110_));
  NA2        o2061(.A(ori_ori_n452_), .B(ori_ori_n53_), .Y(ori_ori_n2111_));
  AOI210     o2062(.A0(ori_ori_n2110_), .A1(ori_ori_n389_), .B0(ori_ori_n2111_), .Y(ori_ori_n2112_));
  OAI210     o2063(.A0(ori_ori_n2108_), .A1(ori_ori_n59_), .B0(ori_ori_n2112_), .Y(ori_ori_n2113_));
  AOI220     o2064(.A0(ori_ori_n626_), .A1(ori_ori_n216_), .B0(ori_ori_n346_), .B1(ori_ori_n212_), .Y(ori_ori_n2114_));
  NA2        o2065(.A(ori_ori_n666_), .B(ori_ori_n891_), .Y(ori_ori_n2115_));
  OAI210     o2066(.A0(ori_ori_n2115_), .A1(ori_ori_n2114_), .B0(ori_ori_n277_), .Y(ori_ori_n2116_));
  AOI210     o2067(.A0(ori_ori_n1936_), .A1(ori_ori_n197_), .B0(ori_ori_n53_), .Y(ori_ori_n2117_));
  NO2        o2068(.A(ori_ori_n133_), .B(ori_ori_n310_), .Y(ori_ori_n2118_));
  AOI220     o2069(.A0(ori_ori_n2118_), .A1(ori_ori_n911_), .B0(ori_ori_n611_), .B1(ori_ori_n322_), .Y(ori_ori_n2119_));
  NA2        o2070(.A(ori_ori_n402_), .B(ori_ori_n450_), .Y(ori_ori_n2120_));
  NO3        o2071(.A(ori_ori_n2120_), .B(ori_ori_n947_), .C(ori_ori_n168_), .Y(ori_ori_n2121_));
  AOI210     o2072(.A0(ori_ori_n1648_), .A1(ori_ori_n1092_), .B0(ori_ori_n2121_), .Y(ori_ori_n2122_));
  NA4        o2073(.A(ori_ori_n2122_), .B(ori_ori_n2119_), .C(ori_ori_n2117_), .D(ori_ori_n2116_), .Y(ori_ori_n2123_));
  NA3        o2074(.A(ori_ori_n2123_), .B(ori_ori_n2113_), .C(ori_ori_n57_), .Y(ori_ori_n2124_));
  BUFFER     o2075(.A(ori_ori_n1093_), .Y(ori_ori_n2125_));
  NA4        o2076(.A(ori_ori_n581_), .B(ori_ori_n1193_), .C(ori_ori_n425_), .D(ori_ori_n50_), .Y(ori_ori_n2126_));
  OAI210     o2077(.A0(ori_ori_n2118_), .A1(ori_ori_n1880_), .B0(x2), .Y(ori_ori_n2127_));
  NA4        o2078(.A(ori_ori_n260_), .B(ori_ori_n144_), .C(ori_ori_n249_), .D(ori_ori_n118_), .Y(ori_ori_n2128_));
  NA3        o2079(.A(ori_ori_n2128_), .B(ori_ori_n2127_), .C(ori_ori_n2126_), .Y(ori_ori_n2129_));
  AO220      o2080(.A0(ori_ori_n2129_), .A1(x0), .B0(ori_ori_n2125_), .B1(ori_ori_n131_), .Y(ori_ori_n2130_));
  NA3        o2081(.A(ori_ori_n699_), .B(ori_ori_n322_), .C(ori_ori_n60_), .Y(ori_ori_n2131_));
  NO2        o2082(.A(ori_ori_n2069_), .B(ori_ori_n370_), .Y(ori_ori_n2132_));
  NA2        o2083(.A(ori_ori_n580_), .B(ori_ori_n468_), .Y(ori_ori_n2133_));
  OAI220     o2084(.A0(ori_ori_n2133_), .A1(ori_ori_n2132_), .B0(ori_ori_n2131_), .B1(ori_ori_n71_), .Y(ori_ori_n2134_));
  OAI210     o2085(.A0(ori_ori_n1398_), .A1(ori_ori_n318_), .B0(ori_ori_n107_), .Y(ori_ori_n2135_));
  AOI210     o2086(.A0(ori_ori_n536_), .A1(ori_ori_n421_), .B0(ori_ori_n131_), .Y(ori_ori_n2136_));
  OAI210     o2087(.A0(ori_ori_n2136_), .A1(ori_ori_n346_), .B0(ori_ori_n2135_), .Y(ori_ori_n2137_));
  OAI210     o2088(.A0(ori_ori_n2137_), .A1(ori_ori_n2134_), .B0(ori_ori_n98_), .Y(ori_ori_n2138_));
  NA2        o2089(.A(ori_ori_n1111_), .B(ori_ori_n341_), .Y(ori_ori_n2139_));
  NA2        o2090(.A(ori_ori_n2139_), .B(ori_ori_n1673_), .Y(ori_ori_n2140_));
  NA2        o2091(.A(ori_ori_n1091_), .B(ori_ori_n647_), .Y(ori_ori_n2141_));
  NA2        o2092(.A(ori_ori_n1245_), .B(ori_ori_n1072_), .Y(ori_ori_n2142_));
  NA4        o2093(.A(ori_ori_n2142_), .B(ori_ori_n2141_), .C(ori_ori_n2140_), .D(ori_ori_n2138_), .Y(ori_ori_n2143_));
  AOI210     o2094(.A0(ori_ori_n2130_), .A1(x7), .B0(ori_ori_n2143_), .Y(ori_ori_n2144_));
  NA3        o2095(.A(ori_ori_n2144_), .B(ori_ori_n2124_), .C(ori_ori_n2106_), .Y(ori34));
  NA2        o2096(.A(ori_ori_n389_), .B(x4), .Y(ori_ori_n2146_));
  NO2        o2097(.A(ori_ori_n1782_), .B(ori_ori_n777_), .Y(ori_ori_n2147_));
  AOI210     o2098(.A0(ori_ori_n2147_), .A1(ori_ori_n2146_), .B0(ori_ori_n292_), .Y(ori_ori_n2148_));
  NA2        o2099(.A(ori_ori_n260_), .B(ori_ori_n119_), .Y(ori_ori_n2149_));
  NO2        o2100(.A(ori_ori_n889_), .B(ori_ori_n2149_), .Y(ori_ori_n2150_));
  AOI210     o2101(.A0(ori_ori_n1860_), .A1(ori_ori_n494_), .B0(ori_ori_n132_), .Y(ori_ori_n2151_));
  NO2        o2102(.A(ori_ori_n1680_), .B(ori_ori_n893_), .Y(ori_ori_n2152_));
  NO4        o2103(.A(ori_ori_n2152_), .B(ori_ori_n2151_), .C(ori_ori_n2150_), .D(ori_ori_n2148_), .Y(ori_ori_n2153_));
  NO2        o2104(.A(ori_ori_n2153_), .B(ori_ori_n431_), .Y(ori_ori_n2154_));
  NA2        o2105(.A(ori_ori_n668_), .B(x8), .Y(ori_ori_n2155_));
  AO210      o2106(.A0(ori_ori_n2155_), .A1(ori_ori_n437_), .B0(ori_ori_n601_), .Y(ori_ori_n2156_));
  NA2        o2107(.A(ori_ori_n611_), .B(ori_ori_n575_), .Y(ori_ori_n2157_));
  AOI210     o2108(.A0(ori_ori_n2157_), .A1(ori_ori_n2156_), .B0(ori_ori_n241_), .Y(ori_ori_n2158_));
  OAI210     o2109(.A0(ori_ori_n118_), .A1(ori_ori_n965_), .B0(ori_ori_n1341_), .Y(ori_ori_n2159_));
  OAI210     o2110(.A0(ori_ori_n1473_), .A1(ori_ori_n58_), .B0(ori_ori_n2159_), .Y(ori_ori_n2160_));
  NA3        o2111(.A(ori_ori_n2160_), .B(ori_ori_n311_), .C(x8), .Y(ori_ori_n2161_));
  NO3        o2112(.A(ori_ori_n910_), .B(ori_ori_n644_), .C(ori_ori_n412_), .Y(ori_ori_n2162_));
  AOI210     o2113(.A0(ori_ori_n1455_), .A1(ori_ori_n299_), .B0(ori_ori_n2162_), .Y(ori_ori_n2163_));
  NA2        o2114(.A(ori_ori_n605_), .B(ori_ori_n292_), .Y(ori_ori_n2164_));
  NA2        o2115(.A(ori_ori_n129_), .B(x0), .Y(ori_ori_n2165_));
  NAi31      o2116(.An(ori_ori_n2165_), .B(ori_ori_n2164_), .C(ori_ori_n721_), .Y(ori_ori_n2166_));
  NA3        o2117(.A(ori_ori_n1468_), .B(ori_ori_n1282_), .C(ori_ori_n50_), .Y(ori_ori_n2167_));
  NA4        o2118(.A(ori_ori_n2167_), .B(ori_ori_n2166_), .C(ori_ori_n2163_), .D(ori_ori_n2161_), .Y(ori_ori_n2168_));
  NA2        o2119(.A(ori_ori_n1016_), .B(ori_ori_n678_), .Y(ori_ori_n2169_));
  NA3        o2120(.A(ori_ori_n1051_), .B(ori_ori_n154_), .C(ori_ori_n1004_), .Y(ori_ori_n2170_));
  AOI210     o2121(.A0(ori_ori_n2170_), .A1(ori_ori_n2169_), .B0(ori_ori_n688_), .Y(ori_ori_n2171_));
  INV        o2122(.A(ori_ori_n2171_), .Y(ori_ori_n2172_));
  INV        o2123(.A(ori_ori_n506_), .Y(ori_ori_n2173_));
  OAI220     o2124(.A0(ori_ori_n2173_), .A1(ori_ori_n59_), .B0(ori_ori_n1027_), .B1(ori_ori_n55_), .Y(ori_ori_n2174_));
  NA3        o2125(.A(ori_ori_n2174_), .B(ori_ori_n668_), .C(ori_ori_n56_), .Y(ori_ori_n2175_));
  OAI210     o2126(.A0(ori_ori_n2172_), .A1(ori_ori_n133_), .B0(ori_ori_n2175_), .Y(ori_ori_n2176_));
  NO4        o2127(.A(ori_ori_n2176_), .B(ori_ori_n2168_), .C(ori_ori_n2158_), .D(ori_ori_n2154_), .Y(ori_ori_n2177_));
  NO2        o2128(.A(ori_ori_n284_), .B(ori_ori_n871_), .Y(ori_ori_n2178_));
  NO3        o2129(.A(ori_ori_n2178_), .B(ori_ori_n400_), .C(ori_ori_n299_), .Y(ori_ori_n2179_));
  NA2        o2130(.A(ori_ori_n707_), .B(ori_ori_n148_), .Y(ori_ori_n2180_));
  NO3        o2131(.A(ori_ori_n2047_), .B(ori_ori_n277_), .C(ori_ori_n1004_), .Y(ori_ori_n2181_));
  OAI220     o2132(.A0(ori_ori_n2181_), .A1(ori_ori_n1426_), .B0(ori_ori_n2180_), .B1(ori_ori_n1076_), .Y(ori_ori_n2182_));
  OAI210     o2133(.A0(ori_ori_n2182_), .A1(ori_ori_n2179_), .B0(x2), .Y(ori_ori_n2183_));
  OAI210     o2134(.A0(ori_ori_n787_), .A1(ori_ori_n335_), .B0(ori_ori_n2183_), .Y(ori_ori_n2184_));
  NA2        o2135(.A(ori_ori_n287_), .B(x4), .Y(ori_ori_n2185_));
  OAI220     o2136(.A0(ori_ori_n674_), .A1(ori_ori_n55_), .B0(ori_ori_n253_), .B1(ori_ori_n103_), .Y(ori_ori_n2186_));
  NO4        o2137(.A(ori_ori_n404_), .B(ori_ori_n77_), .C(x7), .D(x3), .Y(ori_ori_n2187_));
  NO2        o2138(.A(ori_ori_n1016_), .B(ori_ori_n261_), .Y(ori_ori_n2188_));
  NO4        o2139(.A(ori_ori_n2188_), .B(ori_ori_n2187_), .C(ori_ori_n2186_), .D(ori_ori_n2185_), .Y(ori_ori_n2189_));
  NA2        o2140(.A(ori_ori_n1141_), .B(ori_ori_n964_), .Y(ori_ori_n2190_));
  NA3        o2141(.A(ori_ori_n1279_), .B(ori_ori_n233_), .C(x7), .Y(ori_ori_n2191_));
  NA2        o2142(.A(ori_ori_n2191_), .B(ori_ori_n2190_), .Y(ori_ori_n2192_));
  OAI210     o2143(.A0(ori_ori_n2192_), .A1(ori_ori_n2189_), .B0(ori_ori_n152_), .Y(ori_ori_n2193_));
  NA3        o2144(.A(ori_ori_n782_), .B(ori_ori_n87_), .C(x0), .Y(ori_ori_n2194_));
  NA4        o2145(.A(ori_ori_n2194_), .B(ori_ori_n1055_), .C(ori_ori_n270_), .D(ori_ori_n534_), .Y(ori_ori_n2195_));
  NA2        o2146(.A(ori_ori_n1059_), .B(ori_ori_n616_), .Y(ori_ori_n2196_));
  OAI210     o2147(.A0(ori_ori_n2196_), .A1(ori_ori_n242_), .B0(ori_ori_n1985_), .Y(ori_ori_n2197_));
  AOI220     o2148(.A0(ori_ori_n2197_), .A1(x7), .B0(ori_ori_n932_), .B1(ori_ori_n602_), .Y(ori_ori_n2198_));
  NA2        o2149(.A(ori_ori_n90_), .B(x2), .Y(ori_ori_n2199_));
  AOI210     o2150(.A0(ori_ori_n245_), .A1(ori_ori_n53_), .B0(ori_ori_n593_), .Y(ori_ori_n2200_));
  OAI220     o2151(.A0(ori_ori_n2200_), .A1(ori_ori_n93_), .B0(ori_ori_n2199_), .B1(ori_ori_n1231_), .Y(ori_ori_n2201_));
  NA2        o2152(.A(ori_ori_n2201_), .B(ori_ori_n1209_), .Y(ori_ori_n2202_));
  NA4        o2153(.A(ori_ori_n2202_), .B(ori_ori_n2198_), .C(ori_ori_n2195_), .D(ori_ori_n2193_), .Y(ori_ori_n2203_));
  AOI210     o2154(.A0(ori_ori_n2184_), .A1(ori_ori_n738_), .B0(ori_ori_n2203_), .Y(ori_ori_n2204_));
  OAI210     o2155(.A0(ori_ori_n2177_), .A1(x2), .B0(ori_ori_n2204_), .Y(ori35));
  AOI220     o2156(.A0(ori_ori_n580_), .A1(ori_ori_n55_), .B0(ori_ori_n699_), .B1(ori_ori_n1126_), .Y(ori_ori_n2206_));
  NO2        o2157(.A(ori_ori_n2206_), .B(ori_ori_n71_), .Y(ori_ori_n2207_));
  NO2        o2158(.A(ori_ori_n464_), .B(ori_ori_n310_), .Y(ori_ori_n2208_));
  OAI210     o2159(.A0(ori_ori_n2208_), .A1(ori_ori_n2207_), .B0(x2), .Y(ori_ori_n2209_));
  INV        o2160(.A(ori_ori_n247_), .Y(ori_ori_n2210_));
  OAI220     o2161(.A0(ori_ori_n2210_), .A1(ori_ori_n607_), .B0(ori_ori_n183_), .B1(x4), .Y(ori_ori_n2211_));
  NA2        o2162(.A(ori_ori_n2211_), .B(ori_ori_n131_), .Y(ori_ori_n2212_));
  NO2        o2163(.A(ori_ori_n1583_), .B(ori_ori_n626_), .Y(ori_ori_n2213_));
  OAI210     o2164(.A0(ori_ori_n2131_), .A1(x6), .B0(ori_ori_n677_), .Y(ori_ori_n2214_));
  NO2        o2165(.A(ori_ori_n2214_), .B(ori_ori_n2213_), .Y(ori_ori_n2215_));
  NA3        o2166(.A(ori_ori_n2215_), .B(ori_ori_n2212_), .C(ori_ori_n2209_), .Y(ori_ori_n2216_));
  NAi21      o2167(.An(ori_ori_n1551_), .B(ori_ori_n1190_), .Y(ori_ori_n2217_));
  NA2        o2168(.A(ori_ori_n196_), .B(ori_ori_n521_), .Y(ori_ori_n2218_));
  NO2        o2169(.A(ori_ori_n389_), .B(ori_ori_n382_), .Y(ori_ori_n2219_));
  AOI220     o2170(.A0(ori_ori_n2219_), .A1(ori_ori_n2218_), .B0(ori_ori_n2217_), .B1(ori_ori_n56_), .Y(ori_ori_n2220_));
  NA2        o2171(.A(ori_ori_n691_), .B(ori_ori_n636_), .Y(ori_ori_n2221_));
  NO3        o2172(.A(ori_ori_n621_), .B(ori_ori_n55_), .C(x6), .Y(ori_ori_n2222_));
  OAI210     o2173(.A0(ori_ori_n2222_), .A1(ori_ori_n647_), .B0(ori_ori_n200_), .Y(ori_ori_n2223_));
  NA2        o2174(.A(ori_ori_n1217_), .B(ori_ori_n63_), .Y(ori_ori_n2224_));
  NA2        o2175(.A(x6), .B(ori_ori_n426_), .Y(ori_ori_n2225_));
  NA3        o2176(.A(ori_ori_n2225_), .B(ori_ori_n2224_), .C(ori_ori_n2223_), .Y(ori_ori_n2226_));
  NA2        o2177(.A(ori_ori_n2226_), .B(ori_ori_n50_), .Y(ori_ori_n2227_));
  OAI210     o2178(.A0(ori_ori_n2221_), .A1(ori_ori_n2220_), .B0(ori_ori_n2227_), .Y(ori_ori_n2228_));
  AOI210     o2179(.A0(ori_ori_n2216_), .A1(ori_ori_n57_), .B0(ori_ori_n2228_), .Y(ori_ori_n2229_));
  NO3        o2180(.A(ori_ori_n985_), .B(ori_ori_n514_), .C(ori_ori_n119_), .Y(ori_ori_n2230_));
  OAI210     o2181(.A0(ori_ori_n145_), .A1(ori_ori_n67_), .B0(ori_ori_n2230_), .Y(ori_ori_n2231_));
  NO2        o2182(.A(ori_ori_n2231_), .B(ori_ori_n50_), .Y(ori_ori_n2232_));
  NA3        o2183(.A(ori_ori_n421_), .B(ori_ori_n792_), .C(ori_ori_n100_), .Y(ori_ori_n2233_));
  NA2        o2184(.A(ori_ori_n879_), .B(ori_ori_n681_), .Y(ori_ori_n2234_));
  OAI210     o2185(.A0(ori_ori_n231_), .A1(ori_ori_n533_), .B0(ori_ori_n1983_), .Y(ori_ori_n2235_));
  NA3        o2186(.A(ori_ori_n2235_), .B(ori_ori_n2234_), .C(ori_ori_n2233_), .Y(ori_ori_n2236_));
  OAI210     o2187(.A0(ori_ori_n2236_), .A1(ori_ori_n2232_), .B0(ori_ori_n59_), .Y(ori_ori_n2237_));
  AOI210     o2188(.A0(ori_ori_n782_), .A1(ori_ori_n485_), .B0(ori_ori_n1735_), .Y(ori_ori_n2238_));
  AOI210     o2189(.A0(ori_ori_n514_), .A1(ori_ori_n555_), .B0(ori_ori_n2238_), .Y(ori_ori_n2239_));
  XN2        o2190(.A(x4), .B(x3), .Y(ori_ori_n2240_));
  NO3        o2191(.A(ori_ori_n2240_), .B(ori_ori_n606_), .C(ori_ori_n283_), .Y(ori_ori_n2241_));
  NO2        o2192(.A(ori_ori_n2241_), .B(ori_ori_n1337_), .Y(ori_ori_n2242_));
  OAI210     o2193(.A0(ori_ori_n2239_), .A1(x3), .B0(ori_ori_n2242_), .Y(ori_ori_n2243_));
  NO3        o2194(.A(ori_ori_n674_), .B(ori_ori_n784_), .C(ori_ori_n248_), .Y(ori_ori_n2244_));
  OAI210     o2195(.A0(ori_ori_n2244_), .A1(ori_ori_n1337_), .B0(ori_ori_n50_), .Y(ori_ori_n2245_));
  NA3        o2196(.A(ori_ori_n991_), .B(ori_ori_n736_), .C(ori_ori_n230_), .Y(ori_ori_n2246_));
  NA2        o2197(.A(ori_ori_n2246_), .B(ori_ori_n2245_), .Y(ori_ori_n2247_));
  AOI210     o2198(.A0(ori_ori_n2243_), .A1(ori_ori_n536_), .B0(ori_ori_n2247_), .Y(ori_ori_n2248_));
  AOI210     o2199(.A0(ori_ori_n1310_), .A1(ori_ori_n585_), .B0(ori_ori_n623_), .Y(ori_ori_n2249_));
  INV        o2200(.A(ori_ori_n792_), .Y(ori_ori_n2250_));
  OAI210     o2201(.A0(ori_ori_n1783_), .A1(ori_ori_n555_), .B0(ori_ori_n2069_), .Y(ori_ori_n2251_));
  OAI210     o2202(.A0(ori_ori_n2155_), .A1(ori_ori_n2250_), .B0(ori_ori_n2251_), .Y(ori_ori_n2252_));
  OAI210     o2203(.A0(ori_ori_n2252_), .A1(ori_ori_n2249_), .B0(ori_ori_n90_), .Y(ori_ori_n2253_));
  NO2        o2204(.A(ori_ori_n775_), .B(ori_ori_n603_), .Y(ori_ori_n2254_));
  NO2        o2205(.A(ori_ori_n261_), .B(x6), .Y(ori_ori_n2255_));
  OAI210     o2206(.A0(ori_ori_n2254_), .A1(ori_ori_n1641_), .B0(ori_ori_n2255_), .Y(ori_ori_n2256_));
  NA4        o2207(.A(ori_ori_n2256_), .B(ori_ori_n2253_), .C(ori_ori_n2248_), .D(ori_ori_n2237_), .Y(ori_ori_n2257_));
  NO2        o2208(.A(ori_ori_n383_), .B(x1), .Y(ori_ori_n2258_));
  OAI210     o2209(.A0(ori_ori_n421_), .A1(ori_ori_n155_), .B0(ori_ori_n719_), .Y(ori_ori_n2259_));
  AOI210     o2210(.A0(ori_ori_n2259_), .A1(ori_ori_n937_), .B0(ori_ori_n53_), .Y(ori_ori_n2260_));
  NO2        o2211(.A(ori_ori_n2260_), .B(ori_ori_n2258_), .Y(ori_ori_n2261_));
  NA3        o2212(.A(ori_ori_n1312_), .B(ori_ori_n1169_), .C(ori_ori_n742_), .Y(ori_ori_n2262_));
  AOI220     o2213(.A0(ori_ori_n1775_), .A1(ori_ori_n131_), .B0(ori_ori_n375_), .B1(ori_ori_n122_), .Y(ori_ori_n2263_));
  AOI210     o2214(.A0(ori_ori_n2263_), .A1(ori_ori_n2262_), .B0(ori_ori_n1378_), .Y(ori_ori_n2264_));
  NO2        o2215(.A(ori_ori_n580_), .B(x3), .Y(ori_ori_n2265_));
  NO3        o2216(.A(ori_ori_n634_), .B(ori_ori_n1473_), .C(x2), .Y(ori_ori_n2266_));
  AOI220     o2217(.A0(ori_ori_n2266_), .A1(ori_ori_n2265_), .B0(ori_ori_n1748_), .B1(ori_ori_n695_), .Y(ori_ori_n2267_));
  NO2        o2218(.A(ori_ori_n621_), .B(ori_ori_n481_), .Y(ori_ori_n2268_));
  OAI220     o2219(.A0(ori_ori_n1200_), .A1(x8), .B0(ori_ori_n336_), .B1(ori_ori_n321_), .Y(ori_ori_n2269_));
  AOI220     o2220(.A0(ori_ori_n2269_), .A1(ori_ori_n375_), .B0(ori_ori_n2268_), .B1(ori_ori_n836_), .Y(ori_ori_n2270_));
  OAI210     o2221(.A0(ori_ori_n2267_), .A1(ori_ori_n1067_), .B0(ori_ori_n2270_), .Y(ori_ori_n2271_));
  NO2        o2222(.A(ori_ori_n2271_), .B(ori_ori_n2264_), .Y(ori_ori_n2272_));
  OAI210     o2223(.A0(ori_ori_n2261_), .A1(ori_ori_n287_), .B0(ori_ori_n2272_), .Y(ori_ori_n2273_));
  AOI210     o2224(.A0(ori_ori_n2257_), .A1(x5), .B0(ori_ori_n2273_), .Y(ori_ori_n2274_));
  OAI210     o2225(.A0(ori_ori_n2229_), .A1(x5), .B0(ori_ori_n2274_), .Y(ori36));
  NO2        o2226(.A(ori_ori_n784_), .B(ori_ori_n276_), .Y(ori_ori_n2276_));
  NO3        o2227(.A(ori_ori_n118_), .B(ori_ori_n965_), .C(ori_ori_n55_), .Y(ori_ori_n2277_));
  NO3        o2228(.A(ori_ori_n2277_), .B(ori_ori_n1802_), .C(ori_ori_n985_), .Y(ori_ori_n2278_));
  OAI210     o2229(.A0(ori_ori_n2278_), .A1(ori_ori_n2276_), .B0(ori_ori_n106_), .Y(ori_ori_n2279_));
  INV        o2230(.A(ori_ori_n922_), .Y(ori_ori_n2280_));
  OAI210     o2231(.A0(ori_ori_n2033_), .A1(ori_ori_n2280_), .B0(ori_ori_n253_), .Y(ori_ori_n2281_));
  NA2        o2232(.A(ori_ori_n402_), .B(ori_ori_n209_), .Y(ori_ori_n2282_));
  NA3        o2233(.A(ori_ori_n2282_), .B(ori_ori_n2281_), .C(ori_ori_n2279_), .Y(ori_ori_n2283_));
  INV        o2234(.A(x8), .Y(ori_ori_n2284_));
  NO3        o2235(.A(ori_ori_n2284_), .B(ori_ori_n907_), .C(ori_ori_n490_), .Y(ori_ori_n2285_));
  AOI220     o2236(.A0(ori_ori_n277_), .A1(x1), .B0(ori_ori_n130_), .B1(x6), .Y(ori_ori_n2286_));
  AOI210     o2237(.A0(ori_ori_n1004_), .A1(x6), .B0(ori_ori_n379_), .Y(ori_ori_n2287_));
  OAI220     o2238(.A0(ori_ori_n2287_), .A1(ori_ori_n329_), .B0(ori_ori_n2286_), .B1(ori_ori_n422_), .Y(ori_ori_n2288_));
  OAI210     o2239(.A0(ori_ori_n2288_), .A1(ori_ori_n2285_), .B0(ori_ori_n421_), .Y(ori_ori_n2289_));
  NA2        o2240(.A(ori_ori_n611_), .B(ori_ori_n444_), .Y(ori_ori_n2290_));
  AOI210     o2241(.A0(ori_ori_n2290_), .A1(ori_ori_n590_), .B0(ori_ori_n242_), .Y(ori_ori_n2291_));
  NO3        o2242(.A(ori_ori_n1712_), .B(ori_ori_n1472_), .C(ori_ori_n249_), .Y(ori_ori_n2292_));
  NO3        o2243(.A(ori_ori_n2292_), .B(ori_ori_n2291_), .C(ori_ori_n377_), .Y(ori_ori_n2293_));
  OAI210     o2244(.A0(ori_ori_n581_), .A1(ori_ori_n728_), .B0(ori_ori_n897_), .Y(ori_ori_n2294_));
  OAI210     o2245(.A0(ori_ori_n1516_), .A1(ori_ori_n1511_), .B0(ori_ori_n897_), .Y(ori_ori_n2295_));
  AOI220     o2246(.A0(ori_ori_n2295_), .A1(ori_ori_n116_), .B0(ori_ori_n2294_), .B1(ori_ori_n575_), .Y(ori_ori_n2296_));
  NA3        o2247(.A(ori_ori_n2296_), .B(ori_ori_n2293_), .C(ori_ori_n2289_), .Y(ori_ori_n2297_));
  AOI210     o2248(.A0(ori_ori_n2283_), .A1(ori_ori_n311_), .B0(ori_ori_n2297_), .Y(ori_ori_n2298_));
  OAI210     o2249(.A0(ori_ori_n541_), .A1(ori_ori_n469_), .B0(ori_ori_n155_), .Y(ori_ori_n2299_));
  OAI210     o2250(.A0(ori_ori_n1817_), .A1(ori_ori_n70_), .B0(ori_ori_n2299_), .Y(ori_ori_n2300_));
  OAI210     o2251(.A0(ori_ori_n447_), .A1(ori_ori_n218_), .B0(ori_ori_n231_), .Y(ori_ori_n2301_));
  INV        o2252(.A(ori_ori_n160_), .Y(ori_ori_n2302_));
  NA2        o2253(.A(ori_ori_n1113_), .B(ori_ori_n55_), .Y(ori_ori_n2303_));
  OAI210     o2254(.A0(ori_ori_n2303_), .A1(ori_ori_n2302_), .B0(ori_ori_n2301_), .Y(ori_ori_n2304_));
  OAI210     o2255(.A0(ori_ori_n2304_), .A1(ori_ori_n2300_), .B0(ori_ori_n816_), .Y(ori_ori_n2305_));
  AOI210     o2256(.A0(ori_ori_n103_), .A1(ori_ori_n106_), .B0(ori_ori_n312_), .Y(ori_ori_n2306_));
  NA2        o2257(.A(ori_ori_n611_), .B(ori_ori_n1473_), .Y(ori_ori_n2307_));
  OAI220     o2258(.A0(ori_ori_n2307_), .A1(ori_ori_n2306_), .B0(ori_ori_n677_), .B1(ori_ori_n1153_), .Y(ori_ori_n2308_));
  NO2        o2259(.A(ori_ori_n1282_), .B(ori_ori_n527_), .Y(ori_ori_n2309_));
  NO3        o2260(.A(ori_ori_n2309_), .B(ori_ori_n1647_), .C(ori_ori_n634_), .Y(ori_ori_n2310_));
  NO2        o2261(.A(ori_ori_n2310_), .B(ori_ori_n2308_), .Y(ori_ori_n2311_));
  AOI210     o2262(.A0(ori_ori_n2311_), .A1(ori_ori_n2305_), .B0(x7), .Y(ori_ori_n2312_));
  AOI210     o2263(.A0(ori_ori_n536_), .A1(ori_ori_n570_), .B0(ori_ori_n1092_), .Y(ori_ori_n2313_));
  NA3        o2264(.A(ori_ori_n2313_), .B(ori_ori_n910_), .C(ori_ori_n809_), .Y(ori_ori_n2314_));
  NA2        o2265(.A(ori_ori_n2314_), .B(ori_ori_n456_), .Y(ori_ori_n2315_));
  AOI220     o2266(.A0(ori_ori_n1607_), .A1(ori_ori_n234_), .B0(ori_ori_n964_), .B1(ori_ori_n122_), .Y(ori_ori_n2316_));
  NO2        o2267(.A(ori_ori_n2316_), .B(ori_ori_n402_), .Y(ori_ori_n2317_));
  NO2        o2268(.A(ori_ori_n364_), .B(ori_ori_n209_), .Y(ori_ori_n2318_));
  NO3        o2269(.A(ori_ori_n2318_), .B(ori_ori_n1173_), .C(ori_ori_n59_), .Y(ori_ori_n2319_));
  NO2        o2270(.A(ori_ori_n1128_), .B(x6), .Y(ori_ori_n2320_));
  NA3        o2271(.A(ori_ori_n1542_), .B(ori_ori_n253_), .C(ori_ori_n245_), .Y(ori_ori_n2321_));
  NA2        o2272(.A(ori_ori_n2321_), .B(ori_ori_n1497_), .Y(ori_ori_n2322_));
  NO4        o2273(.A(ori_ori_n2322_), .B(ori_ori_n2320_), .C(ori_ori_n2319_), .D(ori_ori_n2317_), .Y(ori_ori_n2323_));
  AOI210     o2274(.A0(ori_ori_n2323_), .A1(ori_ori_n2315_), .B0(ori_ori_n412_), .Y(ori_ori_n2324_));
  NO3        o2275(.A(ori_ori_n2240_), .B(ori_ori_n822_), .C(ori_ori_n455_), .Y(ori_ori_n2325_));
  AOI210     o2276(.A0(ori_ori_n1171_), .A1(ori_ori_n244_), .B0(ori_ori_n2325_), .Y(ori_ori_n2326_));
  OAI210     o2277(.A0(ori_ori_n791_), .A1(ori_ori_n248_), .B0(ori_ori_n354_), .Y(ori_ori_n2327_));
  NA2        o2278(.A(ori_ori_n1113_), .B(ori_ori_n159_), .Y(ori_ori_n2328_));
  NO2        o2279(.A(ori_ori_n561_), .B(ori_ori_n106_), .Y(ori_ori_n2329_));
  AO210      o2280(.A0(ori_ori_n2329_), .A1(ori_ori_n2328_), .B0(ori_ori_n1623_), .Y(ori_ori_n2330_));
  NO2        o2281(.A(ori_ori_n417_), .B(ori_ori_n376_), .Y(ori_ori_n2331_));
  AOI220     o2282(.A0(ori_ori_n2331_), .A1(ori_ori_n2330_), .B0(ori_ori_n2327_), .B1(ori_ori_n268_), .Y(ori_ori_n2332_));
  OAI210     o2283(.A0(ori_ori_n2326_), .A1(x1), .B0(ori_ori_n2332_), .Y(ori_ori_n2333_));
  NO3        o2284(.A(ori_ori_n2333_), .B(ori_ori_n2324_), .C(ori_ori_n2312_), .Y(ori_ori_n2334_));
  OAI210     o2285(.A0(ori_ori_n2298_), .A1(ori_ori_n57_), .B0(ori_ori_n2334_), .Y(ori37));
  NA2        o2286(.A(ori_ori_n982_), .B(x3), .Y(ori_ori_n2336_));
  NA3        o2287(.A(ori_ori_n707_), .B(ori_ori_n148_), .C(ori_ori_n50_), .Y(ori_ori_n2337_));
  AOI210     o2288(.A0(ori_ori_n2337_), .A1(ori_ori_n2336_), .B0(ori_ori_n627_), .Y(ori_ori_n2338_));
  NO3        o2289(.A(ori_ori_n982_), .B(ori_ori_n338_), .C(ori_ori_n463_), .Y(ori_ori_n2339_));
  OAI210     o2290(.A0(ori_ori_n2339_), .A1(ori_ori_n2338_), .B0(ori_ori_n56_), .Y(ori_ori_n2340_));
  AOI220     o2291(.A0(ori_ori_n550_), .A1(ori_ori_n678_), .B0(ori_ori_n421_), .B1(ori_ori_n964_), .Y(ori_ori_n2341_));
  NO2        o2292(.A(ori_ori_n606_), .B(ori_ori_n167_), .Y(ori_ori_n2342_));
  OAI220     o2293(.A0(ori_ori_n2342_), .A1(ori_ori_n760_), .B0(ori_ori_n2341_), .B1(ori_ori_n106_), .Y(ori_ori_n2343_));
  NA2        o2294(.A(ori_ori_n2343_), .B(ori_ori_n71_), .Y(ori_ori_n2344_));
  NA2        o2295(.A(ori_ori_n176_), .B(ori_ori_n413_), .Y(ori_ori_n2345_));
  NA3        o2296(.A(ori_ori_n2345_), .B(ori_ori_n2344_), .C(ori_ori_n2340_), .Y(ori_ori_n2346_));
  NA2        o2297(.A(ori_ori_n382_), .B(ori_ori_n130_), .Y(ori_ori_n2347_));
  NO2        o2298(.A(ori_ori_n1571_), .B(ori_ori_n105_), .Y(ori_ori_n2348_));
  AOI210     o2299(.A0(ori_ori_n1804_), .A1(ori_ori_n785_), .B0(ori_ori_n2348_), .Y(ori_ori_n2349_));
  OAI220     o2300(.A0(ori_ori_n2349_), .A1(ori_ori_n51_), .B0(ori_ori_n1474_), .B1(ori_ori_n2347_), .Y(ori_ori_n2350_));
  AOI210     o2301(.A0(ori_ori_n2346_), .A1(ori_ori_n68_), .B0(ori_ori_n2350_), .Y(ori_ori_n2351_));
  OAI210     o2302(.A0(ori_ori_n245_), .A1(ori_ori_n1008_), .B0(ori_ori_n438_), .Y(ori_ori_n2352_));
  NA3        o2303(.A(ori_ori_n2352_), .B(ori_ori_n242_), .C(ori_ori_n965_), .Y(ori_ori_n2353_));
  OAI210     o2304(.A0(ori_ori_n212_), .A1(ori_ori_n200_), .B0(ori_ori_n1583_), .Y(ori_ori_n2354_));
  NA2        o2305(.A(ori_ori_n316_), .B(ori_ori_n247_), .Y(ori_ori_n2355_));
  NA3        o2306(.A(ori_ori_n360_), .B(ori_ori_n742_), .C(ori_ori_n106_), .Y(ori_ori_n2356_));
  NO2        o2307(.A(ori_ori_n482_), .B(ori_ori_n56_), .Y(ori_ori_n2357_));
  NA3        o2308(.A(ori_ori_n2357_), .B(ori_ori_n2356_), .C(ori_ori_n2355_), .Y(ori_ori_n2358_));
  AOI210     o2309(.A0(ori_ori_n2354_), .A1(ori_ori_n463_), .B0(ori_ori_n2358_), .Y(ori_ori_n2359_));
  NO2        o2310(.A(ori_ori_n1085_), .B(ori_ori_n248_), .Y(ori_ori_n2360_));
  OAI210     o2311(.A0(ori_ori_n268_), .A1(ori_ori_n240_), .B0(ori_ori_n2360_), .Y(ori_ori_n2361_));
  OAI210     o2312(.A0(ori_ori_n608_), .A1(ori_ori_n131_), .B0(x3), .Y(ori_ori_n2362_));
  AOI210     o2313(.A0(ori_ori_n608_), .A1(ori_ori_n333_), .B0(ori_ori_n2362_), .Y(ori_ori_n2363_));
  AOI210     o2314(.A0(ori_ori_n1473_), .A1(ori_ori_n50_), .B0(ori_ori_n316_), .Y(ori_ori_n2364_));
  OAI210     o2315(.A0(ori_ori_n2364_), .A1(ori_ori_n359_), .B0(ori_ori_n56_), .Y(ori_ori_n2365_));
  NO2        o2316(.A(ori_ori_n2365_), .B(ori_ori_n2363_), .Y(ori_ori_n2366_));
  AOI220     o2317(.A0(ori_ori_n2366_), .A1(ori_ori_n2361_), .B0(ori_ori_n2359_), .B1(ori_ori_n2353_), .Y(ori_ori_n2367_));
  OAI210     o2318(.A0(ori_ori_n2367_), .A1(ori_ori_n1621_), .B0(ori_ori_n98_), .Y(ori_ori_n2368_));
  NA2        o2319(.A(ori_ori_n634_), .B(ori_ori_n1098_), .Y(ori_ori_n2369_));
  INV        o2320(.A(ori_ori_n107_), .Y(ori_ori_n2370_));
  AOI210     o2321(.A0(ori_ori_n2370_), .A1(ori_ori_n2369_), .B0(ori_ori_n392_), .Y(ori_ori_n2371_));
  NO2        o2322(.A(ori_ori_n2044_), .B(ori_ori_n55_), .Y(ori_ori_n2372_));
  OAI210     o2323(.A0(ori_ori_n2372_), .A1(ori_ori_n2371_), .B0(ori_ori_n1673_), .Y(ori_ori_n2373_));
  AOI210     o2324(.A0(ori_ori_n323_), .A1(ori_ori_n132_), .B0(ori_ori_n133_), .Y(ori_ori_n2374_));
  NA2        o2325(.A(ori_ori_n2374_), .B(ori_ori_n316_), .Y(ori_ori_n2375_));
  AOI210     o2326(.A0(ori_ori_n562_), .A1(ori_ori_n392_), .B0(ori_ori_n1181_), .Y(ori_ori_n2376_));
  NO3        o2327(.A(ori_ori_n2376_), .B(ori_ori_n242_), .C(ori_ori_n63_), .Y(ori_ori_n2377_));
  NO2        o2328(.A(ori_ori_n1919_), .B(ori_ori_n346_), .Y(ori_ori_n2378_));
  OAI210     o2329(.A0(ori_ori_n2378_), .A1(ori_ori_n2377_), .B0(ori_ori_n53_), .Y(ori_ori_n2379_));
  NO4        o2330(.A(ori_ori_n2165_), .B(ori_ori_n851_), .C(ori_ori_n393_), .D(ori_ori_n203_), .Y(ori_ori_n2380_));
  NO4        o2331(.A(ori_ori_n668_), .B(ori_ori_n551_), .C(ori_ori_n400_), .D(ori_ori_n971_), .Y(ori_ori_n2381_));
  NO3        o2332(.A(ori_ori_n2381_), .B(ori_ori_n2380_), .C(ori_ori_n977_), .Y(ori_ori_n2382_));
  NA4        o2333(.A(ori_ori_n2382_), .B(ori_ori_n2379_), .C(ori_ori_n2375_), .D(ori_ori_n2373_), .Y(ori_ori_n2383_));
  NO3        o2334(.A(ori_ori_n227_), .B(ori_ori_n322_), .C(ori_ori_n84_), .Y(ori_ori_n2384_));
  NO2        o2335(.A(ori_ori_n251_), .B(ori_ori_n699_), .Y(ori_ori_n2385_));
  NO3        o2336(.A(ori_ori_n2385_), .B(ori_ori_n1113_), .C(ori_ori_n1129_), .Y(ori_ori_n2386_));
  OAI220     o2337(.A0(ori_ori_n2386_), .A1(ori_ori_n2384_), .B0(ori_ori_n421_), .B1(ori_ori_n85_), .Y(ori_ori_n2387_));
  OR2        o2338(.A(ori_ori_n857_), .B(ori_ori_n680_), .Y(ori_ori_n2388_));
  NA2        o2339(.A(ori_ori_n1126_), .B(ori_ori_n55_), .Y(ori_ori_n2389_));
  NOi21      o2340(.An(ori_ori_n2389_), .B(ori_ori_n347_), .Y(ori_ori_n2390_));
  AOI210     o2341(.A0(ori_ori_n2390_), .A1(ori_ori_n2388_), .B0(x1), .Y(ori_ori_n2391_));
  NA2        o2342(.A(ori_ori_n241_), .B(ori_ori_n84_), .Y(ori_ori_n2392_));
  AOI210     o2343(.A0(ori_ori_n1426_), .A1(ori_ori_n359_), .B0(ori_ori_n2392_), .Y(ori_ori_n2393_));
  NA2        o2344(.A(ori_ori_n1016_), .B(ori_ori_n62_), .Y(ori_ori_n2394_));
  NA2        o2345(.A(ori_ori_n1059_), .B(ori_ori_n160_), .Y(ori_ori_n2395_));
  OAI210     o2346(.A0(ori_ori_n2394_), .A1(ori_ori_n286_), .B0(ori_ori_n2395_), .Y(ori_ori_n2396_));
  NO3        o2347(.A(ori_ori_n2396_), .B(ori_ori_n2393_), .C(ori_ori_n2391_), .Y(ori_ori_n2397_));
  OAI210     o2348(.A0(ori_ori_n2397_), .A1(x6), .B0(ori_ori_n2387_), .Y(ori_ori_n2398_));
  AOI220     o2349(.A0(ori_ori_n2398_), .A1(ori_ori_n1341_), .B0(ori_ori_n2383_), .B1(ori_ori_n57_), .Y(ori_ori_n2399_));
  NA3        o2350(.A(ori_ori_n2399_), .B(ori_ori_n2368_), .C(ori_ori_n2351_), .Y(ori38));
  NO2        o2351(.A(ori_ori_n172_), .B(ori_ori_n891_), .Y(ori_ori_n2401_));
  NO2        o2352(.A(ori_ori_n526_), .B(ori_ori_n1001_), .Y(ori_ori_n2402_));
  AOI210     o2353(.A0(ori_ori_n2389_), .A1(ori_ori_n1694_), .B0(ori_ori_n211_), .Y(ori_ori_n2403_));
  NO3        o2354(.A(ori_ori_n2403_), .B(ori_ori_n2402_), .C(ori_ori_n2401_), .Y(ori_ori_n2404_));
  NO2        o2355(.A(ori_ori_n2404_), .B(x6), .Y(ori_ori_n2405_));
  NA4        o2356(.A(ori_ori_n340_), .B(ori_ori_n233_), .C(ori_ori_n175_), .D(x8), .Y(ori_ori_n2406_));
  NA2        o2357(.A(ori_ori_n358_), .B(ori_ori_n104_), .Y(ori_ori_n2407_));
  AOI210     o2358(.A0(ori_ori_n2407_), .A1(ori_ori_n2406_), .B0(ori_ori_n133_), .Y(ori_ori_n2408_));
  AOI210     o2359(.A0(ori_ori_n393_), .A1(ori_ori_n363_), .B0(ori_ori_n1593_), .Y(ori_ori_n2409_));
  NO2        o2360(.A(ori_ori_n736_), .B(ori_ori_n90_), .Y(ori_ori_n2410_));
  OAI210     o2361(.A0(ori_ori_n941_), .A1(ori_ori_n138_), .B0(ori_ori_n328_), .Y(ori_ori_n2411_));
  OAI220     o2362(.A0(ori_ori_n2411_), .A1(ori_ori_n2410_), .B0(ori_ori_n2409_), .B1(ori_ori_n175_), .Y(ori_ori_n2412_));
  OAI210     o2363(.A0(ori_ori_n2412_), .A1(ori_ori_n2408_), .B0(x6), .Y(ori_ori_n2413_));
  NO2        o2364(.A(ori_ori_n225_), .B(ori_ori_n699_), .Y(ori_ori_n2414_));
  NO3        o2365(.A(ori_ori_n2414_), .B(ori_ori_n1551_), .C(ori_ori_n233_), .Y(ori_ori_n2415_));
  NO3        o2366(.A(x3), .B(ori_ori_n53_), .C(x0), .Y(ori_ori_n2416_));
  INV        o2367(.A(ori_ori_n2416_), .Y(ori_ori_n2417_));
  NA3        o2368(.A(ori_ori_n392_), .B(ori_ori_n382_), .C(ori_ori_n267_), .Y(ori_ori_n2418_));
  NA2        o2369(.A(ori_ori_n2418_), .B(ori_ori_n2417_), .Y(ori_ori_n2419_));
  OAI210     o2370(.A0(ori_ori_n2419_), .A1(ori_ori_n2415_), .B0(ori_ori_n738_), .Y(ori_ori_n2420_));
  AN3        o2371(.A(ori_ori_n743_), .B(ori_ori_n707_), .C(x0), .Y(ori_ori_n2421_));
  NA2        o2372(.A(ori_ori_n2421_), .B(ori_ori_n300_), .Y(ori_ori_n2422_));
  OAI220     o2373(.A0(ori_ori_n551_), .A1(ori_ori_n249_), .B0(ori_ori_n742_), .B1(ori_ori_n91_), .Y(ori_ori_n2423_));
  OAI210     o2374(.A0(ori_ori_n626_), .A1(x0), .B0(ori_ori_n51_), .Y(ori_ori_n2424_));
  AOI210     o2375(.A0(ori_ori_n532_), .A1(x4), .B0(ori_ori_n210_), .Y(ori_ori_n2425_));
  AOI220     o2376(.A0(ori_ori_n2425_), .A1(ori_ori_n2424_), .B0(ori_ori_n2423_), .B1(ori_ori_n360_), .Y(ori_ori_n2426_));
  NA4        o2377(.A(ori_ori_n2426_), .B(ori_ori_n2422_), .C(ori_ori_n2420_), .D(ori_ori_n2413_), .Y(ori_ori_n2427_));
  OAI210     o2378(.A0(ori_ori_n2427_), .A1(ori_ori_n2405_), .B0(x7), .Y(ori_ori_n2428_));
  AOI210     o2379(.A0(ori_ori_n337_), .A1(x1), .B0(ori_ori_n1133_), .Y(ori_ori_n2429_));
  NO2        o2380(.A(ori_ori_n2429_), .B(ori_ori_n51_), .Y(ori_ori_n2430_));
  AOI210     o2381(.A0(ori_ori_n90_), .A1(ori_ori_n71_), .B0(ori_ori_n2069_), .Y(ori_ori_n2431_));
  NA2        o2382(.A(ori_ori_n346_), .B(x3), .Y(ori_ori_n2432_));
  NO2        o2383(.A(ori_ori_n1613_), .B(ori_ori_n482_), .Y(ori_ori_n2433_));
  OAI210     o2384(.A0(ori_ori_n2432_), .A1(ori_ori_n2431_), .B0(ori_ori_n2433_), .Y(ori_ori_n2434_));
  OAI210     o2385(.A0(ori_ori_n2434_), .A1(ori_ori_n2430_), .B0(x4), .Y(ori_ori_n2435_));
  AOI210     o2386(.A0(ori_ori_n971_), .A1(ori_ori_n220_), .B0(ori_ori_n353_), .Y(ori_ori_n2436_));
  AO210      o2387(.A0(ori_ori_n1194_), .A1(x6), .B0(ori_ori_n2436_), .Y(ori_ori_n2437_));
  NA2        o2388(.A(ori_ori_n1782_), .B(ori_ori_n295_), .Y(ori_ori_n2438_));
  NO2        o2389(.A(ori_ori_n2438_), .B(ori_ori_n990_), .Y(ori_ori_n2439_));
  NO2        o2390(.A(ori_ori_n2439_), .B(ori_ori_n2437_), .Y(ori_ori_n2440_));
  AOI210     o2391(.A0(ori_ori_n2440_), .A1(ori_ori_n2435_), .B0(ori_ori_n104_), .Y(ori_ori_n2441_));
  NA3        o2392(.A(ori_ori_n1775_), .B(ori_ori_n551_), .C(ori_ori_n152_), .Y(ori_ori_n2442_));
  AOI210     o2393(.A0(ori_ori_n2442_), .A1(ori_ori_n1306_), .B0(ori_ori_n212_), .Y(ori_ori_n2443_));
  NO2        o2394(.A(ori_ori_n183_), .B(ori_ori_n115_), .Y(ori_ori_n2444_));
  OAI210     o2395(.A0(ori_ori_n2444_), .A1(ori_ori_n2443_), .B0(x0), .Y(ori_ori_n2445_));
  NA3        o2396(.A(ori_ori_n363_), .B(ori_ori_n742_), .C(ori_ori_n249_), .Y(ori_ori_n2446_));
  AOI210     o2397(.A0(ori_ori_n2446_), .A1(ori_ori_n655_), .B0(ori_ori_n2028_), .Y(ori_ori_n2447_));
  NA2        o2398(.A(ori_ori_n1036_), .B(ori_ori_n871_), .Y(ori_ori_n2448_));
  NA2        o2399(.A(ori_ori_n164_), .B(x3), .Y(ori_ori_n2449_));
  AOI210     o2400(.A0(ori_ori_n2449_), .A1(ori_ori_n2448_), .B0(ori_ori_n450_), .Y(ori_ori_n2450_));
  NO4        o2401(.A(ori_ori_n1293_), .B(ori_ori_n471_), .C(ori_ori_n1129_), .D(ori_ori_n699_), .Y(ori_ori_n2451_));
  NO2        o2402(.A(ori_ori_n1639_), .B(ori_ori_n2109_), .Y(ori_ori_n2452_));
  NO4        o2403(.A(ori_ori_n2452_), .B(ori_ori_n2451_), .C(ori_ori_n2450_), .D(ori_ori_n2447_), .Y(ori_ori_n2453_));
  NA2        o2404(.A(ori_ori_n2453_), .B(ori_ori_n2445_), .Y(ori_ori_n2454_));
  OAI210     o2405(.A0(ori_ori_n2454_), .A1(ori_ori_n2441_), .B0(ori_ori_n57_), .Y(ori_ori_n2455_));
  NO2        o2406(.A(ori_ori_n1674_), .B(ori_ori_n623_), .Y(ori_ori_n2456_));
  OAI210     o2407(.A0(ori_ori_n1620_), .A1(ori_ori_n196_), .B0(ori_ori_n446_), .Y(ori_ori_n2457_));
  OAI210     o2408(.A0(ori_ori_n2457_), .A1(ori_ori_n2456_), .B0(ori_ori_n576_), .Y(ori_ori_n2458_));
  NO2        o2409(.A(ori_ori_n1625_), .B(ori_ori_n249_), .Y(ori_ori_n2459_));
  NA2        o2410(.A(ori_ori_n1706_), .B(ori_ori_n324_), .Y(ori_ori_n2460_));
  OAI220     o2411(.A0(ori_ori_n2460_), .A1(ori_ori_n581_), .B0(ori_ori_n633_), .B1(ori_ori_n140_), .Y(ori_ori_n2461_));
  AOI210     o2412(.A0(ori_ori_n2459_), .A1(ori_ori_n911_), .B0(ori_ori_n2461_), .Y(ori_ori_n2462_));
  NA4        o2413(.A(ori_ori_n2462_), .B(ori_ori_n2458_), .C(ori_ori_n2455_), .D(ori_ori_n2428_), .Y(ori39));
  INV        o2414(.A(ori_ori_n248_), .Y(ori_ori_n2466_));
  INV        m0000(.A(x3), .Y(mai_mai_n50_));
  NA2        m0001(.A(mai_mai_n50_), .B(x2), .Y(mai_mai_n51_));
  NA2        m0002(.A(x7), .B(x0), .Y(mai_mai_n52_));
  INV        m0003(.A(x1), .Y(mai_mai_n53_));
  NA2        m0004(.A(x5), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  INV        m0005(.A(x8), .Y(mai_mai_n55_));
  INV        m0006(.A(x4), .Y(mai_mai_n56_));
  INV        m0007(.A(x7), .Y(mai_mai_n57_));
  NA2        m0008(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0009(.A(x0), .Y(mai_mai_n59_));
  NA2        m0010(.A(x4), .B(mai_mai_n59_), .Y(mai_mai_n60_));
  NA2        m0011(.A(mai_mai_n56_), .B(mai_mai_n59_), .Y(mai_mai_n61_));
  NO2        m0012(.A(mai_mai_n55_), .B(x6), .Y(mai_mai_n62_));
  NA2        m0013(.A(mai_mai_n57_), .B(x4), .Y(mai_mai_n63_));
  NO2        m0014(.A(x8), .B(mai_mai_n57_), .Y(mai_mai_n64_));
  NO2        m0015(.A(x7), .B(mai_mai_n59_), .Y(mai_mai_n65_));
  NAi21      m0016(.An(x5), .B(x1), .Y(mai_mai_n66_));
  INV        m0017(.A(x6), .Y(mai_mai_n67_));
  NA2        m0018(.A(mai_mai_n67_), .B(x4), .Y(mai_mai_n68_));
  NA2        m0019(.A(x7), .B(x4), .Y(mai_mai_n69_));
  NO2        m0020(.A(mai_mai_n69_), .B(x1), .Y(mai_mai_n70_));
  NO2        m0021(.A(mai_mai_n67_), .B(x5), .Y(mai_mai_n71_));
  NO2        m0022(.A(x8), .B(mai_mai_n59_), .Y(mai_mai_n72_));
  NA2        m0023(.A(x5), .B(x3), .Y(mai_mai_n73_));
  NO2        m0024(.A(x6), .B(x0), .Y(mai_mai_n74_));
  NO2        m0025(.A(mai_mai_n74_), .B(x4), .Y(mai_mai_n75_));
  NO2        m0026(.A(x4), .B(x2), .Y(mai_mai_n76_));
  NO2        m0027(.A(mai_mai_n67_), .B(mai_mai_n59_), .Y(mai_mai_n77_));
  NO2        m0028(.A(mai_mai_n77_), .B(mai_mai_n76_), .Y(mai_mai_n78_));
  NA2        m0029(.A(x8), .B(x1), .Y(mai_mai_n79_));
  NO2        m0030(.A(mai_mai_n79_), .B(x7), .Y(mai_mai_n80_));
  INV        m0031(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  OR3        m0032(.A(mai_mai_n81_), .B(mai_mai_n78_), .C(mai_mai_n75_), .Y(mai_mai_n82_));
  NO3        m0033(.A(x8), .B(mai_mai_n57_), .C(x6), .Y(mai_mai_n83_));
  NO2        m0034(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n84_));
  NO2        m0035(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n85_));
  NA3        m0036(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n83_), .Y(mai_mai_n86_));
  AOI210     m0037(.A0(mai_mai_n86_), .A1(mai_mai_n82_), .B0(mai_mai_n73_), .Y(mai_mai_n87_));
  XO2        m0038(.A(x7), .B(x1), .Y(mai_mai_n88_));
  INV        m0039(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  NO2        m0040(.A(mai_mai_n50_), .B(x0), .Y(mai_mai_n90_));
  NA2        m0041(.A(mai_mai_n90_), .B(mai_mai_n55_), .Y(mai_mai_n91_));
  NO2        m0042(.A(x6), .B(x5), .Y(mai_mai_n92_));
  NO2        m0043(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n93_));
  NA2        m0044(.A(x6), .B(x1), .Y(mai_mai_n94_));
  NA2        m0045(.A(x3), .B(x0), .Y(mai_mai_n95_));
  INV        m0046(.A(x5), .Y(mai_mai_n96_));
  NA2        m0047(.A(mai_mai_n67_), .B(mai_mai_n96_), .Y(mai_mai_n97_));
  INV        m0048(.A(x2), .Y(mai_mai_n98_));
  NO2        m0049(.A(mai_mai_n56_), .B(mai_mai_n98_), .Y(mai_mai_n99_));
  NA2        m0050(.A(mai_mai_n57_), .B(mai_mai_n96_), .Y(mai_mai_n100_));
  NA3        m0051(.A(mai_mai_n100_), .B(mai_mai_n99_), .C(mai_mai_n97_), .Y(mai_mai_n101_));
  NO3        m0052(.A(mai_mai_n101_), .B(mai_mai_n95_), .C(mai_mai_n53_), .Y(mai_mai_n102_));
  NO2        m0053(.A(mai_mai_n102_), .B(mai_mai_n87_), .Y(mai00));
  NO2        m0054(.A(x7), .B(x6), .Y(mai_mai_n104_));
  INV        m0055(.A(mai_mai_n104_), .Y(mai_mai_n105_));
  NO2        m0056(.A(mai_mai_n55_), .B(mai_mai_n53_), .Y(mai_mai_n106_));
  NA2        m0057(.A(mai_mai_n106_), .B(mai_mai_n56_), .Y(mai_mai_n107_));
  NO2        m0058(.A(mai_mai_n107_), .B(mai_mai_n105_), .Y(mai_mai_n108_));
  XN2        m0059(.A(x6), .B(x1), .Y(mai_mai_n109_));
  INV        m0060(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NO2        m0061(.A(x6), .B(x4), .Y(mai_mai_n111_));
  NA2        m0062(.A(x6), .B(x4), .Y(mai_mai_n112_));
  NAi21      m0063(.An(mai_mai_n111_), .B(mai_mai_n112_), .Y(mai_mai_n113_));
  XN2        m0064(.A(x7), .B(x6), .Y(mai_mai_n114_));
  NO4        m0065(.A(mai_mai_n114_), .B(mai_mai_n113_), .C(mai_mai_n110_), .D(x8), .Y(mai_mai_n115_));
  NO2        m0066(.A(x3), .B(mai_mai_n98_), .Y(mai_mai_n116_));
  NA2        m0067(.A(mai_mai_n116_), .B(mai_mai_n96_), .Y(mai_mai_n117_));
  NO2        m0068(.A(mai_mai_n117_), .B(mai_mai_n59_), .Y(mai_mai_n118_));
  OAI210     m0069(.A0(mai_mai_n115_), .A1(mai_mai_n108_), .B0(mai_mai_n118_), .Y(mai_mai_n119_));
  NA2        m0070(.A(x3), .B(mai_mai_n98_), .Y(mai_mai_n120_));
  NO2        m0071(.A(mai_mai_n55_), .B(mai_mai_n57_), .Y(mai_mai_n121_));
  NA2        m0072(.A(mai_mai_n121_), .B(mai_mai_n56_), .Y(mai_mai_n122_));
  NA2        m0073(.A(mai_mai_n55_), .B(mai_mai_n57_), .Y(mai_mai_n123_));
  NA2        m0074(.A(mai_mai_n123_), .B(x2), .Y(mai_mai_n124_));
  NA2        m0075(.A(x8), .B(x3), .Y(mai_mai_n125_));
  NA2        m0076(.A(mai_mai_n125_), .B(mai_mai_n69_), .Y(mai_mai_n126_));
  OAI220     m0077(.A0(mai_mai_n126_), .A1(mai_mai_n124_), .B0(mai_mai_n122_), .B1(mai_mai_n120_), .Y(mai_mai_n127_));
  NO2        m0078(.A(x5), .B(x0), .Y(mai_mai_n128_));
  NO2        m0079(.A(x6), .B(x1), .Y(mai_mai_n129_));
  NA3        m0080(.A(mai_mai_n129_), .B(mai_mai_n128_), .C(mai_mai_n127_), .Y(mai_mai_n130_));
  NA2        m0081(.A(x8), .B(mai_mai_n96_), .Y(mai_mai_n131_));
  NA2        m0082(.A(x4), .B(mai_mai_n50_), .Y(mai_mai_n132_));
  NO3        m0083(.A(mai_mai_n132_), .B(mai_mai_n131_), .C(mai_mai_n94_), .Y(mai_mai_n133_));
  NAi21      m0084(.An(x7), .B(x2), .Y(mai_mai_n134_));
  NO2        m0085(.A(mai_mai_n134_), .B(x0), .Y(mai_mai_n135_));
  XO2        m0086(.A(x8), .B(x7), .Y(mai_mai_n136_));
  NA2        m0087(.A(mai_mai_n136_), .B(mai_mai_n98_), .Y(mai_mai_n137_));
  NA2        m0088(.A(x6), .B(x5), .Y(mai_mai_n138_));
  NO2        m0089(.A(mai_mai_n56_), .B(x0), .Y(mai_mai_n139_));
  NO2        m0090(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n140_));
  NA2        m0091(.A(mai_mai_n140_), .B(mai_mai_n139_), .Y(mai_mai_n141_));
  NA2        m0092(.A(mai_mai_n135_), .B(mai_mai_n133_), .Y(mai_mai_n142_));
  NA3        m0093(.A(mai_mai_n142_), .B(mai_mai_n130_), .C(mai_mai_n119_), .Y(mai01));
  NA2        m0094(.A(mai_mai_n57_), .B(mai_mai_n59_), .Y(mai_mai_n144_));
  NO2        m0095(.A(x2), .B(x1), .Y(mai_mai_n145_));
  NA2        m0096(.A(x2), .B(x1), .Y(mai_mai_n146_));
  NOi21      m0097(.An(mai_mai_n146_), .B(mai_mai_n145_), .Y(mai_mai_n147_));
  NA2        m0098(.A(mai_mai_n96_), .B(mai_mai_n53_), .Y(mai_mai_n148_));
  NAi21      m0099(.An(x8), .B(x1), .Y(mai_mai_n149_));
  NO2        m0100(.A(mai_mai_n149_), .B(x3), .Y(mai_mai_n150_));
  NA2        m0101(.A(mai_mai_n150_), .B(mai_mai_n147_), .Y(mai_mai_n151_));
  NO2        m0102(.A(x5), .B(mai_mai_n50_), .Y(mai_mai_n152_));
  NO2        m0103(.A(mai_mai_n98_), .B(x1), .Y(mai_mai_n153_));
  NA2        m0104(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  AOI210     m0105(.A0(mai_mai_n154_), .A1(mai_mai_n151_), .B0(mai_mai_n144_), .Y(mai_mai_n155_));
  NAi21      m0106(.An(x7), .B(x0), .Y(mai_mai_n156_));
  NO2        m0107(.A(mai_mai_n55_), .B(x2), .Y(mai_mai_n157_));
  NO2        m0108(.A(mai_mai_n73_), .B(x1), .Y(mai_mai_n158_));
  NA2        m0109(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NA2        m0110(.A(x5), .B(mai_mai_n50_), .Y(mai_mai_n160_));
  NO2        m0111(.A(mai_mai_n160_), .B(mai_mai_n149_), .Y(mai_mai_n161_));
  NA2        m0112(.A(x8), .B(x5), .Y(mai_mai_n162_));
  NO2        m0113(.A(mai_mai_n162_), .B(mai_mai_n51_), .Y(mai_mai_n163_));
  NO3        m0114(.A(x3), .B(mai_mai_n98_), .C(mai_mai_n53_), .Y(mai_mai_n164_));
  NO3        m0115(.A(mai_mai_n164_), .B(mai_mai_n163_), .C(mai_mai_n161_), .Y(mai_mai_n165_));
  AOI210     m0116(.A0(mai_mai_n165_), .A1(mai_mai_n159_), .B0(mai_mai_n156_), .Y(mai_mai_n166_));
  NO2        m0117(.A(mai_mai_n57_), .B(x3), .Y(mai_mai_n167_));
  NO2        m0118(.A(mai_mai_n55_), .B(x0), .Y(mai_mai_n168_));
  NA3        m0119(.A(mai_mai_n96_), .B(mai_mai_n98_), .C(x1), .Y(mai_mai_n169_));
  NO2        m0120(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  NO2        m0121(.A(mai_mai_n79_), .B(mai_mai_n50_), .Y(mai_mai_n171_));
  NA2        m0122(.A(mai_mai_n96_), .B(x0), .Y(mai_mai_n172_));
  NO2        m0123(.A(mai_mai_n172_), .B(x2), .Y(mai_mai_n173_));
  AOI220     m0124(.A0(mai_mai_n173_), .A1(mai_mai_n171_), .B0(mai_mai_n170_), .B1(mai_mai_n167_), .Y(mai_mai_n174_));
  NA2        m0125(.A(x7), .B(mai_mai_n98_), .Y(mai_mai_n175_));
  NA2        m0126(.A(mai_mai_n152_), .B(x8), .Y(mai_mai_n176_));
  NA4        m0127(.A(x5), .B(x3), .C(x1), .D(x0), .Y(mai_mai_n177_));
  AO210      m0128(.A0(mai_mai_n177_), .A1(mai_mai_n176_), .B0(mai_mai_n175_), .Y(mai_mai_n178_));
  NO2        m0129(.A(mai_mai_n146_), .B(mai_mai_n50_), .Y(mai_mai_n179_));
  NAi21      m0130(.An(x1), .B(x2), .Y(mai_mai_n180_));
  NO2        m0131(.A(mai_mai_n160_), .B(mai_mai_n180_), .Y(mai_mai_n181_));
  NA2        m0132(.A(x8), .B(x7), .Y(mai_mai_n182_));
  NO2        m0133(.A(mai_mai_n182_), .B(x0), .Y(mai_mai_n183_));
  OAI210     m0134(.A0(mai_mai_n181_), .A1(mai_mai_n179_), .B0(mai_mai_n183_), .Y(mai_mai_n184_));
  NA3        m0135(.A(mai_mai_n184_), .B(mai_mai_n178_), .C(mai_mai_n174_), .Y(mai_mai_n185_));
  NO3        m0136(.A(mai_mai_n185_), .B(mai_mai_n166_), .C(mai_mai_n155_), .Y(mai_mai_n186_));
  NA2        m0137(.A(x3), .B(x1), .Y(mai_mai_n187_));
  NA2        m0138(.A(mai_mai_n50_), .B(mai_mai_n98_), .Y(mai_mai_n188_));
  NO2        m0139(.A(mai_mai_n188_), .B(mai_mai_n66_), .Y(mai_mai_n189_));
  OAI210     m0140(.A0(mai_mai_n189_), .A1(mai_mai_n181_), .B0(mai_mai_n64_), .Y(mai_mai_n190_));
  NA2        m0141(.A(mai_mai_n121_), .B(mai_mai_n98_), .Y(mai_mai_n191_));
  OAI210     m0142(.A0(mai_mai_n191_), .A1(mai_mai_n187_), .B0(mai_mai_n190_), .Y(mai_mai_n192_));
  XO2        m0143(.A(x5), .B(x3), .Y(mai_mai_n193_));
  NA2        m0144(.A(mai_mai_n193_), .B(x8), .Y(mai_mai_n194_));
  NA2        m0145(.A(x8), .B(mai_mai_n59_), .Y(mai_mai_n195_));
  NA2        m0146(.A(mai_mai_n195_), .B(mai_mai_n125_), .Y(mai_mai_n196_));
  NA2        m0147(.A(x7), .B(mai_mai_n67_), .Y(mai_mai_n197_));
  NO2        m0148(.A(mai_mai_n180_), .B(mai_mai_n197_), .Y(mai_mai_n198_));
  OA210      m0149(.A0(mai_mai_n196_), .A1(mai_mai_n193_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  AOI220     m0150(.A0(mai_mai_n199_), .A1(mai_mai_n194_), .B0(mai_mai_n192_), .B1(x0), .Y(mai_mai_n200_));
  OAI210     m0151(.A0(mai_mai_n186_), .A1(mai_mai_n67_), .B0(mai_mai_n200_), .Y(mai_mai_n201_));
  NO2        m0152(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n202_));
  NA4        m0153(.A(mai_mai_n55_), .B(x5), .C(x3), .D(x2), .Y(mai_mai_n203_));
  NA2        m0154(.A(x8), .B(mai_mai_n50_), .Y(mai_mai_n204_));
  NA2        m0155(.A(mai_mai_n204_), .B(x2), .Y(mai_mai_n205_));
  NA2        m0156(.A(mai_mai_n55_), .B(x3), .Y(mai_mai_n206_));
  NA3        m0157(.A(mai_mai_n205_), .B(mai_mai_n193_), .C(mai_mai_n74_), .Y(mai_mai_n207_));
  AOI210     m0158(.A0(mai_mai_n207_), .A1(mai_mai_n203_), .B0(mai_mai_n53_), .Y(mai_mai_n208_));
  NO2        m0159(.A(mai_mai_n98_), .B(mai_mai_n59_), .Y(mai_mai_n209_));
  NA2        m0160(.A(x5), .B(x1), .Y(mai_mai_n210_));
  NO2        m0161(.A(mai_mai_n210_), .B(x6), .Y(mai_mai_n211_));
  NO2        m0162(.A(x3), .B(x1), .Y(mai_mai_n212_));
  NO2        m0163(.A(mai_mai_n73_), .B(mai_mai_n55_), .Y(mai_mai_n213_));
  NO2        m0164(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n214_));
  NA2        m0165(.A(mai_mai_n214_), .B(mai_mai_n67_), .Y(mai_mai_n215_));
  NAi21      m0166(.An(x2), .B(x5), .Y(mai_mai_n216_));
  NA2        m0167(.A(x8), .B(x6), .Y(mai_mai_n217_));
  OAI210     m0168(.A0(mai_mai_n217_), .A1(mai_mai_n216_), .B0(mai_mai_n215_), .Y(mai_mai_n218_));
  NA2        m0169(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n219_));
  NO2        m0170(.A(mai_mai_n219_), .B(mai_mai_n59_), .Y(mai_mai_n220_));
  AO220      m0171(.A0(mai_mai_n220_), .A1(mai_mai_n218_), .B0(mai_mai_n211_), .B1(mai_mai_n209_), .Y(mai_mai_n221_));
  OAI210     m0172(.A0(mai_mai_n221_), .A1(mai_mai_n208_), .B0(mai_mai_n202_), .Y(mai_mai_n222_));
  NA2        m0173(.A(mai_mai_n67_), .B(mai_mai_n56_), .Y(mai_mai_n223_));
  NO2        m0174(.A(mai_mai_n223_), .B(x7), .Y(mai_mai_n224_));
  NO2        m0175(.A(mai_mai_n96_), .B(mai_mai_n53_), .Y(mai_mai_n225_));
  NA2        m0176(.A(mai_mai_n225_), .B(mai_mai_n98_), .Y(mai_mai_n226_));
  AOI210     m0177(.A0(mai_mai_n226_), .A1(mai_mai_n154_), .B0(mai_mai_n59_), .Y(mai_mai_n227_));
  NA2        m0178(.A(x3), .B(mai_mai_n59_), .Y(mai_mai_n228_));
  NO2        m0179(.A(mai_mai_n169_), .B(mai_mai_n228_), .Y(mai_mai_n229_));
  OA210      m0180(.A0(mai_mai_n229_), .A1(mai_mai_n227_), .B0(x8), .Y(mai_mai_n230_));
  NO2        m0181(.A(x1), .B(x0), .Y(mai_mai_n231_));
  NA2        m0182(.A(mai_mai_n231_), .B(mai_mai_n98_), .Y(mai_mai_n232_));
  NA2        m0183(.A(mai_mai_n96_), .B(mai_mai_n50_), .Y(mai_mai_n233_));
  XN2        m0184(.A(x3), .B(x2), .Y(mai_mai_n234_));
  NA2        m0185(.A(mai_mai_n234_), .B(mai_mai_n147_), .Y(mai_mai_n235_));
  NO2        m0186(.A(mai_mai_n96_), .B(x0), .Y(mai_mai_n236_));
  NA2        m0187(.A(x8), .B(mai_mai_n53_), .Y(mai_mai_n237_));
  NA2        m0188(.A(mai_mai_n237_), .B(mai_mai_n236_), .Y(mai_mai_n238_));
  OAI220     m0189(.A0(mai_mai_n238_), .A1(mai_mai_n235_), .B0(mai_mai_n233_), .B1(mai_mai_n232_), .Y(mai_mai_n239_));
  OAI210     m0190(.A0(mai_mai_n239_), .A1(mai_mai_n230_), .B0(mai_mai_n224_), .Y(mai_mai_n240_));
  NO2        m0191(.A(x7), .B(x1), .Y(mai_mai_n241_));
  NOi21      m0192(.An(x8), .B(x3), .Y(mai_mai_n242_));
  NA2        m0193(.A(mai_mai_n242_), .B(mai_mai_n59_), .Y(mai_mai_n243_));
  NA2        m0194(.A(x5), .B(x0), .Y(mai_mai_n244_));
  NAi21      m0195(.An(mai_mai_n128_), .B(mai_mai_n244_), .Y(mai_mai_n245_));
  NA2        m0196(.A(mai_mai_n67_), .B(mai_mai_n50_), .Y(mai_mai_n246_));
  OAI210     m0197(.A0(mai_mai_n246_), .A1(mai_mai_n245_), .B0(mai_mai_n243_), .Y(mai_mai_n247_));
  NA3        m0198(.A(mai_mai_n247_), .B(mai_mai_n131_), .C(mai_mai_n241_), .Y(mai_mai_n248_));
  NA2        m0199(.A(x8), .B(mai_mai_n57_), .Y(mai_mai_n249_));
  NO2        m0200(.A(mai_mai_n249_), .B(x5), .Y(mai_mai_n250_));
  NO2        m0201(.A(mai_mai_n140_), .B(mai_mai_n67_), .Y(mai_mai_n251_));
  NA2        m0202(.A(x1), .B(x0), .Y(mai_mai_n252_));
  NA2        m0203(.A(mai_mai_n50_), .B(mai_mai_n59_), .Y(mai_mai_n253_));
  NA4        m0204(.A(mai_mai_n253_), .B(mai_mai_n252_), .C(mai_mai_n251_), .D(mai_mai_n250_), .Y(mai_mai_n254_));
  NA3        m0205(.A(mai_mai_n254_), .B(mai_mai_n248_), .C(mai_mai_n177_), .Y(mai_mai_n255_));
  NO2        m0206(.A(mai_mai_n96_), .B(x3), .Y(mai_mai_n256_));
  NO2        m0207(.A(mai_mai_n98_), .B(x0), .Y(mai_mai_n257_));
  NA2        m0208(.A(mai_mai_n257_), .B(mai_mai_n256_), .Y(mai_mai_n258_));
  NO2        m0209(.A(mai_mai_n55_), .B(x7), .Y(mai_mai_n259_));
  NA2        m0210(.A(mai_mai_n259_), .B(mai_mai_n129_), .Y(mai_mai_n260_));
  NO3        m0211(.A(x8), .B(mai_mai_n50_), .C(x0), .Y(mai_mai_n261_));
  NAi21      m0212(.An(x8), .B(x0), .Y(mai_mai_n262_));
  NAi21      m0213(.An(x1), .B(x3), .Y(mai_mai_n263_));
  NO2        m0214(.A(mai_mai_n263_), .B(mai_mai_n262_), .Y(mai_mai_n264_));
  NO2        m0215(.A(x2), .B(mai_mai_n53_), .Y(mai_mai_n265_));
  AOI210     m0216(.A0(mai_mai_n265_), .A1(mai_mai_n261_), .B0(mai_mai_n264_), .Y(mai_mai_n266_));
  NOi21      m0217(.An(x5), .B(x6), .Y(mai_mai_n267_));
  NO2        m0218(.A(mai_mai_n57_), .B(x4), .Y(mai_mai_n268_));
  NA2        m0219(.A(mai_mai_n268_), .B(mai_mai_n267_), .Y(mai_mai_n269_));
  OAI220     m0220(.A0(mai_mai_n269_), .A1(mai_mai_n266_), .B0(mai_mai_n260_), .B1(mai_mai_n258_), .Y(mai_mai_n270_));
  AOI210     m0221(.A0(mai_mai_n255_), .A1(mai_mai_n99_), .B0(mai_mai_n270_), .Y(mai_mai_n271_));
  NA3        m0222(.A(mai_mai_n271_), .B(mai_mai_n240_), .C(mai_mai_n222_), .Y(mai_mai_n272_));
  AOI210     m0223(.A0(mai_mai_n201_), .A1(mai_mai_n56_), .B0(mai_mai_n272_), .Y(mai02));
  NO2        m0224(.A(x8), .B(mai_mai_n96_), .Y(mai_mai_n274_));
  XN2        m0225(.A(x7), .B(x3), .Y(mai_mai_n275_));
  INV        m0226(.A(mai_mai_n275_), .Y(mai_mai_n276_));
  NO2        m0227(.A(x2), .B(x0), .Y(mai_mai_n277_));
  NA2        m0228(.A(mai_mai_n277_), .B(mai_mai_n67_), .Y(mai_mai_n278_));
  NO2        m0229(.A(mai_mai_n57_), .B(x1), .Y(mai_mai_n279_));
  NO3        m0230(.A(mai_mai_n279_), .B(mai_mai_n278_), .C(mai_mai_n276_), .Y(mai_mai_n280_));
  NA2        m0231(.A(mai_mai_n53_), .B(x0), .Y(mai_mai_n281_));
  NO2        m0232(.A(mai_mai_n263_), .B(x6), .Y(mai_mai_n282_));
  XO2        m0233(.A(x7), .B(x0), .Y(mai_mai_n283_));
  NO2        m0234(.A(mai_mai_n283_), .B(mai_mai_n277_), .Y(mai_mai_n284_));
  NA2        m0235(.A(mai_mai_n284_), .B(mai_mai_n282_), .Y(mai_mai_n285_));
  AN2        m0236(.A(x7), .B(x2), .Y(mai_mai_n286_));
  NA2        m0237(.A(mai_mai_n286_), .B(mai_mai_n50_), .Y(mai_mai_n287_));
  OAI210     m0238(.A0(mai_mai_n287_), .A1(mai_mai_n281_), .B0(mai_mai_n285_), .Y(mai_mai_n288_));
  OAI210     m0239(.A0(mai_mai_n288_), .A1(mai_mai_n280_), .B0(mai_mai_n274_), .Y(mai_mai_n289_));
  NAi21      m0240(.An(x8), .B(x6), .Y(mai_mai_n290_));
  NO2        m0241(.A(mai_mai_n96_), .B(mai_mai_n59_), .Y(mai_mai_n291_));
  NA2        m0242(.A(x7), .B(x3), .Y(mai_mai_n292_));
  NO2        m0243(.A(mai_mai_n292_), .B(x2), .Y(mai_mai_n293_));
  NA2        m0244(.A(x2), .B(x0), .Y(mai_mai_n294_));
  NA2        m0245(.A(mai_mai_n98_), .B(mai_mai_n59_), .Y(mai_mai_n295_));
  NA2        m0246(.A(mai_mai_n295_), .B(mai_mai_n294_), .Y(mai_mai_n296_));
  NAi21      m0247(.An(x7), .B(x1), .Y(mai_mai_n297_));
  NO2        m0248(.A(mai_mai_n297_), .B(x3), .Y(mai_mai_n298_));
  AOI220     m0249(.A0(mai_mai_n298_), .A1(mai_mai_n296_), .B0(mai_mai_n293_), .B1(mai_mai_n291_), .Y(mai_mai_n299_));
  NA2        m0250(.A(mai_mai_n265_), .B(mai_mai_n50_), .Y(mai_mai_n300_));
  NA3        m0251(.A(x7), .B(mai_mai_n96_), .C(x0), .Y(mai_mai_n301_));
  NA2        m0252(.A(mai_mai_n257_), .B(mai_mai_n53_), .Y(mai_mai_n302_));
  NA2        m0253(.A(mai_mai_n152_), .B(mai_mai_n57_), .Y(mai_mai_n303_));
  OA220      m0254(.A0(mai_mai_n303_), .A1(mai_mai_n302_), .B0(mai_mai_n301_), .B1(mai_mai_n300_), .Y(mai_mai_n304_));
  AOI210     m0255(.A0(mai_mai_n304_), .A1(mai_mai_n299_), .B0(mai_mai_n290_), .Y(mai_mai_n305_));
  INV        m0256(.A(mai_mai_n283_), .Y(mai_mai_n306_));
  NO2        m0257(.A(x7), .B(mai_mai_n67_), .Y(mai_mai_n307_));
  NA2        m0258(.A(mai_mai_n96_), .B(x3), .Y(mai_mai_n308_));
  NO2        m0259(.A(mai_mai_n308_), .B(mai_mai_n307_), .Y(mai_mai_n309_));
  NA2        m0260(.A(mai_mai_n309_), .B(mai_mai_n306_), .Y(mai_mai_n310_));
  NA2        m0261(.A(mai_mai_n50_), .B(x0), .Y(mai_mai_n311_));
  NO2        m0262(.A(mai_mai_n311_), .B(x7), .Y(mai_mai_n312_));
  NA2        m0263(.A(mai_mai_n312_), .B(mai_mai_n267_), .Y(mai_mai_n313_));
  NA2        m0264(.A(mai_mai_n157_), .B(x1), .Y(mai_mai_n314_));
  AOI210     m0265(.A0(mai_mai_n313_), .A1(mai_mai_n310_), .B0(mai_mai_n314_), .Y(mai_mai_n315_));
  NO2        m0266(.A(mai_mai_n57_), .B(mai_mai_n50_), .Y(mai_mai_n316_));
  NO2        m0267(.A(mai_mai_n55_), .B(mai_mai_n98_), .Y(mai_mai_n317_));
  NA3        m0268(.A(mai_mai_n317_), .B(mai_mai_n316_), .C(mai_mai_n59_), .Y(mai_mai_n318_));
  NO2        m0269(.A(mai_mai_n148_), .B(x6), .Y(mai_mai_n319_));
  NO2        m0270(.A(mai_mai_n94_), .B(mai_mai_n96_), .Y(mai_mai_n320_));
  NA2        m0271(.A(mai_mai_n57_), .B(mai_mai_n98_), .Y(mai_mai_n321_));
  NO2        m0272(.A(mai_mai_n321_), .B(mai_mai_n253_), .Y(mai_mai_n322_));
  OAI210     m0273(.A0(mai_mai_n320_), .A1(mai_mai_n319_), .B0(mai_mai_n322_), .Y(mai_mai_n323_));
  OAI210     m0274(.A0(mai_mai_n318_), .A1(mai_mai_n94_), .B0(mai_mai_n323_), .Y(mai_mai_n324_));
  NO3        m0275(.A(mai_mai_n324_), .B(mai_mai_n315_), .C(mai_mai_n305_), .Y(mai_mai_n325_));
  AOI210     m0276(.A0(mai_mai_n325_), .A1(mai_mai_n289_), .B0(x4), .Y(mai_mai_n326_));
  NA2        m0277(.A(x8), .B(mai_mai_n67_), .Y(mai_mai_n327_));
  NO2        m0278(.A(x3), .B(mai_mai_n59_), .Y(mai_mai_n328_));
  NA3        m0279(.A(mai_mai_n328_), .B(mai_mai_n96_), .C(mai_mai_n53_), .Y(mai_mai_n329_));
  NO2        m0280(.A(x3), .B(x0), .Y(mai_mai_n330_));
  NAi21      m0281(.An(mai_mai_n330_), .B(mai_mai_n95_), .Y(mai_mai_n331_));
  NA2        m0282(.A(x5), .B(x2), .Y(mai_mai_n332_));
  NO2        m0283(.A(mai_mai_n332_), .B(mai_mai_n212_), .Y(mai_mai_n333_));
  AOI210     m0284(.A0(mai_mai_n333_), .A1(mai_mai_n331_), .B0(mai_mai_n229_), .Y(mai_mai_n334_));
  AO210      m0285(.A0(mai_mai_n334_), .A1(mai_mai_n329_), .B0(mai_mai_n327_), .Y(mai_mai_n335_));
  NO2        m0286(.A(mai_mai_n98_), .B(mai_mai_n53_), .Y(mai_mai_n336_));
  NA2        m0287(.A(mai_mai_n336_), .B(x3), .Y(mai_mai_n337_));
  NO2        m0288(.A(mai_mai_n55_), .B(x1), .Y(mai_mai_n338_));
  NA2        m0289(.A(mai_mai_n338_), .B(mai_mai_n98_), .Y(mai_mai_n339_));
  NO2        m0290(.A(mai_mai_n339_), .B(mai_mai_n160_), .Y(mai_mai_n340_));
  NAi32      m0291(.An(x3), .Bn(x0), .C(x2), .Y(mai_mai_n341_));
  NO2        m0292(.A(mai_mai_n50_), .B(x2), .Y(mai_mai_n342_));
  NAi21      m0293(.An(x6), .B(x5), .Y(mai_mai_n343_));
  NO2        m0294(.A(x2), .B(mai_mai_n59_), .Y(mai_mai_n344_));
  NO4        m0295(.A(mai_mai_n344_), .B(mai_mai_n343_), .C(mai_mai_n149_), .D(mai_mai_n342_), .Y(mai_mai_n345_));
  AOI220     m0296(.A0(mai_mai_n345_), .A1(mai_mai_n341_), .B0(mai_mai_n340_), .B1(mai_mai_n77_), .Y(mai_mai_n346_));
  AOI210     m0297(.A0(mai_mai_n346_), .A1(mai_mai_n335_), .B0(mai_mai_n69_), .Y(mai_mai_n347_));
  NA2        m0298(.A(mai_mai_n338_), .B(mai_mai_n56_), .Y(mai_mai_n348_));
  NO2        m0299(.A(mai_mai_n96_), .B(mai_mai_n50_), .Y(mai_mai_n349_));
  NO2        m0300(.A(mai_mai_n277_), .B(mai_mai_n209_), .Y(mai_mai_n350_));
  XO2        m0301(.A(x7), .B(x2), .Y(mai_mai_n351_));
  INV        m0302(.A(mai_mai_n351_), .Y(mai_mai_n352_));
  XO2        m0303(.A(x6), .B(x2), .Y(mai_mai_n353_));
  NA4        m0304(.A(mai_mai_n353_), .B(mai_mai_n352_), .C(mai_mai_n350_), .D(mai_mai_n349_), .Y(mai_mai_n354_));
  NAi21      m0305(.An(x0), .B(x6), .Y(mai_mai_n355_));
  AOI210     m0306(.A0(mai_mai_n355_), .A1(mai_mai_n134_), .B0(mai_mai_n257_), .Y(mai_mai_n356_));
  XN2        m0307(.A(x7), .B(x5), .Y(mai_mai_n357_));
  NA2        m0308(.A(mai_mai_n357_), .B(mai_mai_n67_), .Y(mai_mai_n358_));
  NA2        m0309(.A(x7), .B(x5), .Y(mai_mai_n359_));
  AOI210     m0310(.A0(mai_mai_n359_), .A1(x6), .B0(mai_mai_n341_), .Y(mai_mai_n360_));
  AOI220     m0311(.A0(mai_mai_n360_), .A1(mai_mai_n358_), .B0(mai_mai_n356_), .B1(mai_mai_n309_), .Y(mai_mai_n361_));
  AOI210     m0312(.A0(mai_mai_n361_), .A1(mai_mai_n354_), .B0(mai_mai_n348_), .Y(mai_mai_n362_));
  NO2        m0313(.A(x8), .B(x6), .Y(mai_mai_n363_));
  NAi21      m0314(.An(mai_mai_n363_), .B(mai_mai_n217_), .Y(mai_mai_n364_));
  AOI210     m0315(.A0(mai_mai_n364_), .A1(mai_mai_n84_), .B0(x3), .Y(mai_mai_n365_));
  NA2        m0316(.A(mai_mai_n96_), .B(x2), .Y(mai_mai_n366_));
  NO2        m0317(.A(mai_mai_n366_), .B(mai_mai_n63_), .Y(mai_mai_n367_));
  NA2        m0318(.A(x1), .B(mai_mai_n59_), .Y(mai_mai_n368_));
  NO2        m0319(.A(mai_mai_n368_), .B(mai_mai_n217_), .Y(mai_mai_n369_));
  OAI210     m0320(.A0(mai_mai_n369_), .A1(mai_mai_n50_), .B0(mai_mai_n367_), .Y(mai_mai_n370_));
  NA2        m0321(.A(x4), .B(x2), .Y(mai_mai_n371_));
  NO2        m0322(.A(mai_mai_n371_), .B(mai_mai_n96_), .Y(mai_mai_n372_));
  NAi21      m0323(.An(x1), .B(x6), .Y(mai_mai_n373_));
  NA2        m0324(.A(mai_mai_n330_), .B(mai_mai_n259_), .Y(mai_mai_n374_));
  OAI220     m0325(.A0(mai_mai_n374_), .A1(mai_mai_n373_), .B0(mai_mai_n95_), .B1(mai_mai_n53_), .Y(mai_mai_n375_));
  NA2        m0326(.A(x8), .B(x2), .Y(mai_mai_n376_));
  NO2        m0327(.A(mai_mai_n376_), .B(mai_mai_n50_), .Y(mai_mai_n377_));
  INV        m0328(.A(mai_mai_n211_), .Y(mai_mai_n378_));
  NO2        m0329(.A(mai_mai_n378_), .B(mai_mai_n52_), .Y(mai_mai_n379_));
  AOI220     m0330(.A0(mai_mai_n379_), .A1(mai_mai_n377_), .B0(mai_mai_n375_), .B1(mai_mai_n372_), .Y(mai_mai_n380_));
  OAI210     m0331(.A0(mai_mai_n370_), .A1(mai_mai_n365_), .B0(mai_mai_n380_), .Y(mai_mai_n381_));
  NO4        m0332(.A(mai_mai_n381_), .B(mai_mai_n362_), .C(mai_mai_n347_), .D(mai_mai_n326_), .Y(mai03));
  NAi21      m0333(.An(x2), .B(x0), .Y(mai_mai_n383_));
  NO3        m0334(.A(x8), .B(x6), .C(x4), .Y(mai_mai_n384_));
  INV        m0335(.A(mai_mai_n384_), .Y(mai_mai_n385_));
  NO2        m0336(.A(mai_mai_n385_), .B(mai_mai_n383_), .Y(mai_mai_n386_));
  NA2        m0337(.A(mai_mai_n99_), .B(mai_mai_n59_), .Y(mai_mai_n387_));
  NO2        m0338(.A(mai_mai_n387_), .B(mai_mai_n55_), .Y(mai_mai_n388_));
  OAI210     m0339(.A0(mai_mai_n388_), .A1(mai_mai_n386_), .B0(mai_mai_n152_), .Y(mai_mai_n389_));
  NA2        m0340(.A(x3), .B(x2), .Y(mai_mai_n390_));
  NO2        m0341(.A(mai_mai_n149_), .B(x0), .Y(mai_mai_n391_));
  NA2        m0342(.A(x8), .B(x0), .Y(mai_mai_n392_));
  NO2        m0343(.A(mai_mai_n392_), .B(x6), .Y(mai_mai_n393_));
  AOI210     m0344(.A0(mai_mai_n393_), .A1(x5), .B0(mai_mai_n391_), .Y(mai_mai_n394_));
  NO2        m0345(.A(mai_mai_n394_), .B(mai_mai_n390_), .Y(mai_mai_n395_));
  NO2        m0346(.A(x5), .B(mai_mai_n59_), .Y(mai_mai_n396_));
  NO2        m0347(.A(x3), .B(x2), .Y(mai_mai_n397_));
  NA2        m0348(.A(mai_mai_n397_), .B(mai_mai_n396_), .Y(mai_mai_n398_));
  NO2        m0349(.A(mai_mai_n53_), .B(x0), .Y(mai_mai_n399_));
  NA2        m0350(.A(mai_mai_n399_), .B(x5), .Y(mai_mai_n400_));
  NO2        m0351(.A(mai_mai_n400_), .B(mai_mai_n290_), .Y(mai_mai_n401_));
  NA2        m0352(.A(mai_mai_n243_), .B(mai_mai_n162_), .Y(mai_mai_n402_));
  NO2        m0353(.A(mai_mai_n50_), .B(mai_mai_n59_), .Y(mai_mai_n403_));
  NO2        m0354(.A(mai_mai_n67_), .B(x0), .Y(mai_mai_n404_));
  NO4        m0355(.A(mai_mai_n404_), .B(mai_mai_n403_), .C(x2), .D(mai_mai_n53_), .Y(mai_mai_n405_));
  AO210      m0356(.A0(mai_mai_n405_), .A1(mai_mai_n402_), .B0(mai_mai_n401_), .Y(mai_mai_n406_));
  OAI210     m0357(.A0(mai_mai_n406_), .A1(mai_mai_n395_), .B0(x4), .Y(mai_mai_n407_));
  NO2        m0358(.A(x4), .B(mai_mai_n53_), .Y(mai_mai_n408_));
  NA2        m0359(.A(mai_mai_n408_), .B(mai_mai_n59_), .Y(mai_mai_n409_));
  NO3        m0360(.A(mai_mai_n409_), .B(mai_mai_n217_), .C(x5), .Y(mai_mai_n410_));
  NA2        m0361(.A(x7), .B(mai_mai_n96_), .Y(mai_mai_n411_));
  NO3        m0362(.A(x5), .B(mai_mai_n53_), .C(x0), .Y(mai_mai_n412_));
  INV        m0363(.A(mai_mai_n412_), .Y(mai_mai_n413_));
  NO2        m0364(.A(x6), .B(mai_mai_n56_), .Y(mai_mai_n414_));
  NO2        m0365(.A(x8), .B(mai_mai_n50_), .Y(mai_mai_n415_));
  NA2        m0366(.A(mai_mai_n415_), .B(mai_mai_n414_), .Y(mai_mai_n416_));
  OAI210     m0367(.A0(mai_mai_n416_), .A1(mai_mai_n413_), .B0(mai_mai_n411_), .Y(mai_mai_n417_));
  AOI210     m0368(.A0(mai_mai_n410_), .A1(x2), .B0(mai_mai_n417_), .Y(mai_mai_n418_));
  AOI220     m0369(.A0(mai_mai_n418_), .A1(mai_mai_n407_), .B0(mai_mai_n389_), .B1(x7), .Y(mai_mai_n419_));
  NA2        m0370(.A(x7), .B(mai_mai_n53_), .Y(mai_mai_n420_));
  NO2        m0371(.A(mai_mai_n242_), .B(mai_mai_n98_), .Y(mai_mai_n421_));
  NO2        m0372(.A(mai_mai_n55_), .B(mai_mai_n59_), .Y(mai_mai_n422_));
  NO3        m0373(.A(mai_mai_n422_), .B(mai_mai_n421_), .C(mai_mai_n138_), .Y(mai_mai_n423_));
  AOI210     m0374(.A0(mai_mai_n196_), .A1(mai_mai_n92_), .B0(mai_mai_n423_), .Y(mai_mai_n424_));
  NO2        m0375(.A(x5), .B(x2), .Y(mai_mai_n425_));
  NO2        m0376(.A(x8), .B(x3), .Y(mai_mai_n426_));
  NA2        m0377(.A(mai_mai_n426_), .B(mai_mai_n425_), .Y(mai_mai_n427_));
  NO2        m0378(.A(mai_mai_n427_), .B(x6), .Y(mai_mai_n428_));
  NA2        m0379(.A(mai_mai_n195_), .B(x2), .Y(mai_mai_n429_));
  NO3        m0380(.A(mai_mai_n426_), .B(mai_mai_n331_), .C(mai_mai_n343_), .Y(mai_mai_n430_));
  AOI210     m0381(.A0(mai_mai_n430_), .A1(mai_mai_n429_), .B0(mai_mai_n428_), .Y(mai_mai_n431_));
  OAI210     m0382(.A0(mai_mai_n424_), .A1(mai_mai_n277_), .B0(mai_mai_n431_), .Y(mai_mai_n432_));
  NA2        m0383(.A(mai_mai_n432_), .B(x4), .Y(mai_mai_n433_));
  NA2        m0384(.A(mai_mai_n55_), .B(mai_mai_n59_), .Y(mai_mai_n434_));
  NO2        m0385(.A(mai_mai_n434_), .B(x5), .Y(mai_mai_n435_));
  NAi21      m0386(.An(x4), .B(x6), .Y(mai_mai_n436_));
  NO2        m0387(.A(mai_mai_n55_), .B(mai_mai_n67_), .Y(mai_mai_n437_));
  NO2        m0388(.A(mai_mai_n50_), .B(mai_mai_n98_), .Y(mai_mai_n438_));
  NO2        m0389(.A(mai_mai_n217_), .B(x0), .Y(mai_mai_n439_));
  NO2        m0390(.A(mai_mai_n343_), .B(x8), .Y(mai_mai_n440_));
  OAI210     m0391(.A0(mai_mai_n440_), .A1(mai_mai_n439_), .B0(mai_mai_n438_), .Y(mai_mai_n441_));
  OAI210     m0392(.A0(mai_mai_n398_), .A1(mai_mai_n437_), .B0(mai_mai_n441_), .Y(mai_mai_n442_));
  NA2        m0393(.A(mai_mai_n442_), .B(mai_mai_n56_), .Y(mai_mai_n443_));
  AOI210     m0394(.A0(mai_mai_n443_), .A1(mai_mai_n433_), .B0(mai_mai_n420_), .Y(mai_mai_n444_));
  NA2        m0395(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n445_));
  NO2        m0396(.A(mai_mai_n67_), .B(mai_mai_n56_), .Y(mai_mai_n446_));
  NA2        m0397(.A(mai_mai_n342_), .B(mai_mai_n59_), .Y(mai_mai_n447_));
  OAI220     m0398(.A0(mai_mai_n447_), .A1(mai_mai_n55_), .B0(mai_mai_n188_), .B1(mai_mai_n262_), .Y(mai_mai_n448_));
  NA2        m0399(.A(mai_mai_n448_), .B(mai_mai_n446_), .Y(mai_mai_n449_));
  NO3        m0400(.A(x6), .B(x4), .C(mai_mai_n50_), .Y(mai_mai_n450_));
  NA2        m0401(.A(mai_mai_n422_), .B(x5), .Y(mai_mai_n451_));
  NO2        m0402(.A(x8), .B(x5), .Y(mai_mai_n452_));
  NAi21      m0403(.An(mai_mai_n452_), .B(mai_mai_n162_), .Y(mai_mai_n453_));
  INV        m0404(.A(mai_mai_n451_), .Y(mai_mai_n454_));
  NA2        m0405(.A(mai_mai_n350_), .B(mai_mai_n71_), .Y(mai_mai_n455_));
  NOi21      m0406(.An(x3), .B(x4), .Y(mai_mai_n456_));
  NA2        m0407(.A(mai_mai_n55_), .B(mai_mai_n98_), .Y(mai_mai_n457_));
  NA2        m0408(.A(mai_mai_n457_), .B(mai_mai_n456_), .Y(mai_mai_n458_));
  NO2        m0409(.A(mai_mai_n51_), .B(x6), .Y(mai_mai_n459_));
  NO2        m0410(.A(mai_mai_n138_), .B(mai_mai_n55_), .Y(mai_mai_n460_));
  NO3        m0411(.A(mai_mai_n56_), .B(x2), .C(x0), .Y(mai_mai_n461_));
  AOI220     m0412(.A0(mai_mai_n461_), .A1(mai_mai_n460_), .B0(mai_mai_n459_), .B1(mai_mai_n435_), .Y(mai_mai_n462_));
  OAI210     m0413(.A0(mai_mai_n458_), .A1(mai_mai_n455_), .B0(mai_mai_n462_), .Y(mai_mai_n463_));
  AOI210     m0414(.A0(mai_mai_n454_), .A1(mai_mai_n450_), .B0(mai_mai_n463_), .Y(mai_mai_n464_));
  AOI210     m0415(.A0(mai_mai_n464_), .A1(mai_mai_n449_), .B0(mai_mai_n445_), .Y(mai_mai_n465_));
  NA2        m0416(.A(x7), .B(x1), .Y(mai_mai_n466_));
  NO3        m0417(.A(x5), .B(x4), .C(x2), .Y(mai_mai_n467_));
  AN2        m0418(.A(mai_mai_n467_), .B(mai_mai_n363_), .Y(mai_mai_n468_));
  NO3        m0419(.A(mai_mai_n468_), .B(mai_mai_n460_), .C(mai_mai_n372_), .Y(mai_mai_n469_));
  OAI210     m0420(.A0(mai_mai_n363_), .A1(mai_mai_n76_), .B0(mai_mai_n330_), .Y(mai_mai_n470_));
  NO2        m0421(.A(mai_mai_n470_), .B(mai_mai_n469_), .Y(mai_mai_n471_));
  NO2        m0422(.A(x4), .B(mai_mai_n98_), .Y(mai_mai_n472_));
  NA2        m0423(.A(mai_mai_n472_), .B(x6), .Y(mai_mai_n473_));
  NA3        m0424(.A(mai_mai_n96_), .B(x4), .C(mai_mai_n98_), .Y(mai_mai_n474_));
  NO2        m0425(.A(mai_mai_n473_), .B(mai_mai_n91_), .Y(mai_mai_n475_));
  NA2        m0426(.A(mai_mai_n456_), .B(mai_mai_n67_), .Y(mai_mai_n476_));
  NA2        m0427(.A(mai_mai_n157_), .B(mai_mai_n59_), .Y(mai_mai_n477_));
  NO2        m0428(.A(mai_mai_n477_), .B(mai_mai_n476_), .Y(mai_mai_n478_));
  NA2        m0429(.A(mai_mai_n438_), .B(x4), .Y(mai_mai_n479_));
  NO3        m0430(.A(mai_mai_n479_), .B(mai_mai_n363_), .C(mai_mai_n404_), .Y(mai_mai_n480_));
  NO4        m0431(.A(mai_mai_n480_), .B(mai_mai_n478_), .C(mai_mai_n475_), .D(mai_mai_n471_), .Y(mai_mai_n481_));
  NA2        m0432(.A(x5), .B(x4), .Y(mai_mai_n482_));
  NO2        m0433(.A(mai_mai_n67_), .B(mai_mai_n53_), .Y(mai_mai_n483_));
  NO3        m0434(.A(x8), .B(x3), .C(x2), .Y(mai_mai_n484_));
  NO3        m0435(.A(x6), .B(x5), .C(x2), .Y(mai_mai_n485_));
  NA3        m0436(.A(mai_mai_n485_), .B(mai_mai_n279_), .C(mai_mai_n72_), .Y(mai_mai_n486_));
  INV        m0437(.A(mai_mai_n486_), .Y(mai_mai_n487_));
  NA2        m0438(.A(mai_mai_n67_), .B(x2), .Y(mai_mai_n488_));
  NO3        m0439(.A(x4), .B(x3), .C(mai_mai_n59_), .Y(mai_mai_n489_));
  NA2        m0440(.A(mai_mai_n489_), .B(mai_mai_n214_), .Y(mai_mai_n490_));
  NO3        m0441(.A(mai_mai_n490_), .B(mai_mai_n488_), .C(mai_mai_n88_), .Y(mai_mai_n491_));
  XO2        m0442(.A(x4), .B(x0), .Y(mai_mai_n492_));
  NA2        m0443(.A(mai_mai_n253_), .B(x5), .Y(mai_mai_n493_));
  NO2        m0444(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n494_));
  NO2        m0445(.A(mai_mai_n494_), .B(mai_mai_n62_), .Y(mai_mai_n495_));
  NO4        m0446(.A(mai_mai_n495_), .B(mai_mai_n493_), .C(mai_mai_n492_), .D(mai_mai_n146_), .Y(mai_mai_n496_));
  NO3        m0447(.A(mai_mai_n496_), .B(mai_mai_n491_), .C(mai_mai_n487_), .Y(mai_mai_n497_));
  OAI210     m0448(.A0(mai_mai_n481_), .A1(mai_mai_n466_), .B0(mai_mai_n497_), .Y(mai_mai_n498_));
  NO4        m0449(.A(mai_mai_n498_), .B(mai_mai_n465_), .C(mai_mai_n444_), .D(mai_mai_n419_), .Y(mai04));
  NO2        m0450(.A(x7), .B(x2), .Y(mai_mai_n500_));
  NO2        m0451(.A(x3), .B(mai_mai_n53_), .Y(mai_mai_n501_));
  NO2        m0452(.A(mai_mai_n501_), .B(mai_mai_n140_), .Y(mai_mai_n502_));
  XN2        m0453(.A(x8), .B(x1), .Y(mai_mai_n503_));
  NO2        m0454(.A(mai_mai_n503_), .B(mai_mai_n138_), .Y(mai_mai_n504_));
  NA2        m0455(.A(mai_mai_n504_), .B(mai_mai_n502_), .Y(mai_mai_n505_));
  NA2        m0456(.A(x6), .B(x3), .Y(mai_mai_n506_));
  NO2        m0457(.A(mai_mai_n506_), .B(x5), .Y(mai_mai_n507_));
  NA2        m0458(.A(mai_mai_n67_), .B(x1), .Y(mai_mai_n508_));
  NO2        m0459(.A(mai_mai_n452_), .B(mai_mai_n242_), .Y(mai_mai_n509_));
  NO2        m0460(.A(mai_mai_n509_), .B(mai_mai_n508_), .Y(mai_mai_n510_));
  AOI210     m0461(.A0(mai_mai_n507_), .A1(mai_mai_n338_), .B0(mai_mai_n510_), .Y(mai_mai_n511_));
  AOI210     m0462(.A0(mai_mai_n511_), .A1(mai_mai_n505_), .B0(x0), .Y(mai_mai_n512_));
  NOi21      m0463(.An(mai_mai_n162_), .B(mai_mai_n452_), .Y(mai_mai_n513_));
  NA2        m0464(.A(mai_mai_n97_), .B(x1), .Y(mai_mai_n514_));
  NO3        m0465(.A(mai_mai_n514_), .B(mai_mai_n513_), .C(mai_mai_n311_), .Y(mai_mai_n515_));
  OAI210     m0466(.A0(mai_mai_n515_), .A1(mai_mai_n512_), .B0(mai_mai_n500_), .Y(mai_mai_n516_));
  NA2        m0467(.A(mai_mai_n125_), .B(mai_mai_n228_), .Y(mai_mai_n517_));
  OR4        m0468(.A(mai_mai_n517_), .B(mai_mai_n364_), .C(mai_mai_n74_), .D(mai_mai_n54_), .Y(mai_mai_n518_));
  OR2        m0469(.A(x6), .B(x0), .Y(mai_mai_n519_));
  NO3        m0470(.A(mai_mai_n519_), .B(x3), .C(x1), .Y(mai_mai_n520_));
  AOI220     m0471(.A0(mai_mai_n520_), .A1(mai_mai_n96_), .B0(mai_mai_n267_), .B1(mai_mai_n261_), .Y(mai_mai_n521_));
  AOI210     m0472(.A0(mai_mai_n521_), .A1(mai_mai_n518_), .B0(mai_mai_n175_), .Y(mai_mai_n522_));
  NA2        m0473(.A(x7), .B(x2), .Y(mai_mai_n523_));
  INV        m0474(.A(mai_mai_n125_), .Y(mai_mai_n524_));
  OAI210     m0475(.A0(mai_mai_n161_), .A1(mai_mai_n524_), .B0(mai_mai_n74_), .Y(mai_mai_n525_));
  NO2        m0476(.A(mai_mai_n308_), .B(mai_mai_n55_), .Y(mai_mai_n526_));
  NO3        m0477(.A(x3), .B(x1), .C(x0), .Y(mai_mai_n527_));
  OR2        m0478(.A(x6), .B(x1), .Y(mai_mai_n528_));
  NA2        m0479(.A(mai_mai_n528_), .B(x0), .Y(mai_mai_n529_));
  AOI220     m0480(.A0(mai_mai_n529_), .A1(mai_mai_n526_), .B0(mai_mai_n527_), .B1(mai_mai_n460_), .Y(mai_mai_n530_));
  AOI210     m0481(.A0(mai_mai_n530_), .A1(mai_mai_n525_), .B0(mai_mai_n523_), .Y(mai_mai_n531_));
  NA2        m0482(.A(mai_mai_n67_), .B(x0), .Y(mai_mai_n532_));
  NOi31      m0483(.An(mai_mai_n333_), .B(mai_mai_n532_), .C(mai_mai_n249_), .Y(mai_mai_n533_));
  NO4        m0484(.A(mai_mai_n533_), .B(mai_mai_n531_), .C(mai_mai_n522_), .D(mai_mai_n56_), .Y(mai_mai_n534_));
  NA2        m0485(.A(mai_mai_n534_), .B(mai_mai_n516_), .Y(mai_mai_n535_));
  NA3        m0486(.A(x8), .B(x7), .C(x0), .Y(mai_mai_n536_));
  INV        m0487(.A(mai_mai_n536_), .Y(mai_mai_n537_));
  AOI210     m0488(.A0(mai_mai_n259_), .A1(mai_mai_n90_), .B0(mai_mai_n537_), .Y(mai_mai_n538_));
  NO2        m0489(.A(mai_mai_n538_), .B(mai_mai_n146_), .Y(mai_mai_n539_));
  NA2        m0490(.A(mai_mai_n422_), .B(mai_mai_n57_), .Y(mai_mai_n540_));
  NO2        m0491(.A(x8), .B(x0), .Y(mai_mai_n541_));
  NA2        m0492(.A(mai_mai_n541_), .B(mai_mai_n352_), .Y(mai_mai_n542_));
  AOI210     m0493(.A0(mai_mai_n542_), .A1(mai_mai_n540_), .B0(mai_mai_n263_), .Y(mai_mai_n543_));
  OAI210     m0494(.A0(mai_mai_n543_), .A1(mai_mai_n539_), .B0(mai_mai_n267_), .Y(mai_mai_n544_));
  NO2        m0495(.A(mai_mai_n67_), .B(mai_mai_n98_), .Y(mai_mai_n545_));
  NO2        m0496(.A(mai_mai_n359_), .B(x8), .Y(mai_mai_n546_));
  NO2        m0497(.A(mai_mai_n546_), .B(mai_mai_n250_), .Y(mai_mai_n547_));
  NO2        m0498(.A(mai_mai_n547_), .B(mai_mai_n368_), .Y(mai_mai_n548_));
  NO2        m0499(.A(mai_mai_n276_), .B(x8), .Y(mai_mai_n549_));
  OAI210     m0500(.A0(mai_mai_n452_), .A1(mai_mai_n316_), .B0(mai_mai_n231_), .Y(mai_mai_n550_));
  NA2        m0501(.A(mai_mai_n338_), .B(mai_mai_n167_), .Y(mai_mai_n551_));
  OAI220     m0502(.A0(mai_mai_n551_), .A1(mai_mai_n59_), .B0(mai_mai_n550_), .B1(mai_mai_n549_), .Y(mai_mai_n552_));
  OAI210     m0503(.A0(mai_mai_n552_), .A1(mai_mai_n548_), .B0(mai_mai_n545_), .Y(mai_mai_n553_));
  NO2        m0504(.A(x8), .B(x2), .Y(mai_mai_n554_));
  NO2        m0505(.A(mai_mai_n212_), .B(mai_mai_n57_), .Y(mai_mai_n555_));
  NA3        m0506(.A(mai_mai_n555_), .B(mai_mai_n554_), .C(mai_mai_n331_), .Y(mai_mai_n556_));
  NO2        m0507(.A(mai_mai_n232_), .B(mai_mai_n125_), .Y(mai_mai_n557_));
  AOI210     m0508(.A0(mai_mai_n312_), .A1(mai_mai_n153_), .B0(mai_mai_n557_), .Y(mai_mai_n558_));
  AOI210     m0509(.A0(mai_mai_n558_), .A1(mai_mai_n556_), .B0(mai_mai_n97_), .Y(mai_mai_n559_));
  NA2        m0510(.A(mai_mai_n328_), .B(x2), .Y(mai_mai_n560_));
  NO2        m0511(.A(mai_mai_n57_), .B(mai_mai_n53_), .Y(mai_mai_n561_));
  NA2        m0512(.A(mai_mai_n561_), .B(mai_mai_n62_), .Y(mai_mai_n562_));
  AOI210     m0513(.A0(mai_mai_n560_), .A1(mai_mai_n447_), .B0(mai_mai_n562_), .Y(mai_mai_n563_));
  NA2        m0514(.A(mai_mai_n98_), .B(mai_mai_n53_), .Y(mai_mai_n564_));
  NA2        m0515(.A(x7), .B(mai_mai_n50_), .Y(mai_mai_n565_));
  NO2        m0516(.A(mai_mai_n172_), .B(mai_mai_n565_), .Y(mai_mai_n566_));
  NA2        m0517(.A(mai_mai_n396_), .B(mai_mai_n140_), .Y(mai_mai_n567_));
  NO2        m0518(.A(mai_mai_n67_), .B(x2), .Y(mai_mai_n568_));
  NA2        m0519(.A(mai_mai_n568_), .B(mai_mai_n259_), .Y(mai_mai_n569_));
  NO3        m0520(.A(x4), .B(mai_mai_n563_), .C(mai_mai_n559_), .Y(mai_mai_n570_));
  NA3        m0521(.A(mai_mai_n570_), .B(mai_mai_n553_), .C(mai_mai_n544_), .Y(mai_mai_n571_));
  NA2        m0522(.A(mai_mai_n53_), .B(mai_mai_n59_), .Y(mai_mai_n572_));
  NOi21      m0523(.An(x2), .B(x7), .Y(mai_mai_n573_));
  NO2        m0524(.A(x6), .B(x3), .Y(mai_mai_n574_));
  NA2        m0525(.A(mai_mai_n574_), .B(mai_mai_n573_), .Y(mai_mai_n575_));
  NO2        m0526(.A(x6), .B(mai_mai_n59_), .Y(mai_mai_n576_));
  NO3        m0527(.A(mai_mai_n57_), .B(x2), .C(x1), .Y(mai_mai_n577_));
  NO3        m0528(.A(mai_mai_n57_), .B(x2), .C(x0), .Y(mai_mai_n578_));
  NA2        m0529(.A(mai_mai_n577_), .B(mai_mai_n576_), .Y(mai_mai_n579_));
  OAI210     m0530(.A0(mai_mai_n575_), .A1(mai_mai_n572_), .B0(mai_mai_n579_), .Y(mai_mai_n580_));
  NO2        m0531(.A(mai_mai_n92_), .B(mai_mai_n53_), .Y(mai_mai_n581_));
  NA2        m0532(.A(mai_mai_n210_), .B(mai_mai_n57_), .Y(mai_mai_n582_));
  OAI210     m0533(.A0(mai_mai_n581_), .A1(mai_mai_n440_), .B0(mai_mai_n582_), .Y(mai_mai_n583_));
  NO3        m0534(.A(mai_mai_n583_), .B(mai_mai_n479_), .C(mai_mai_n59_), .Y(mai_mai_n584_));
  AO210      m0535(.A0(mai_mai_n580_), .A1(mai_mai_n452_), .B0(mai_mai_n584_), .Y(mai_mai_n585_));
  AOI210     m0536(.A0(mai_mai_n571_), .A1(mai_mai_n535_), .B0(mai_mai_n585_), .Y(mai05));
  NO2        m0537(.A(x7), .B(mai_mai_n96_), .Y(mai_mai_n587_));
  NO2        m0538(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n588_));
  NA2        m0539(.A(x5), .B(mai_mai_n56_), .Y(mai_mai_n589_));
  NO2        m0540(.A(mai_mai_n589_), .B(mai_mai_n565_), .Y(mai_mai_n590_));
  NO2        m0541(.A(x7), .B(x4), .Y(mai_mai_n591_));
  NO2        m0542(.A(mai_mai_n63_), .B(mai_mai_n55_), .Y(mai_mai_n592_));
  NO2        m0543(.A(mai_mai_n188_), .B(x5), .Y(mai_mai_n593_));
  NA2        m0544(.A(mai_mai_n96_), .B(mai_mai_n98_), .Y(mai_mai_n594_));
  NO2        m0545(.A(mai_mai_n594_), .B(mai_mai_n206_), .Y(mai_mai_n595_));
  AN2        m0546(.A(mai_mai_n595_), .B(mai_mai_n591_), .Y(mai_mai_n596_));
  NA2        m0547(.A(mai_mai_n596_), .B(mai_mai_n483_), .Y(mai_mai_n597_));
  NO2        m0548(.A(x6), .B(mai_mai_n50_), .Y(mai_mai_n598_));
  NA2        m0549(.A(mai_mai_n55_), .B(x4), .Y(mai_mai_n599_));
  NO2        m0550(.A(mai_mai_n96_), .B(mai_mai_n98_), .Y(mai_mai_n600_));
  NA2        m0551(.A(mai_mai_n600_), .B(x7), .Y(mai_mai_n601_));
  NA2        m0552(.A(mai_mai_n425_), .B(mai_mai_n241_), .Y(mai_mai_n602_));
  AOI210     m0553(.A0(mai_mai_n602_), .A1(mai_mai_n601_), .B0(mai_mai_n599_), .Y(mai_mai_n603_));
  NA2        m0554(.A(mai_mai_n96_), .B(x4), .Y(mai_mai_n604_));
  XO2        m0555(.A(x7), .B(x5), .Y(mai_mai_n605_));
  NO2        m0556(.A(mai_mai_n605_), .B(mai_mai_n53_), .Y(mai_mai_n606_));
  NA3        m0557(.A(mai_mai_n606_), .B(mai_mai_n604_), .C(mai_mai_n317_), .Y(mai_mai_n607_));
  NO2        m0558(.A(mai_mai_n96_), .B(x2), .Y(mai_mai_n608_));
  NO2        m0559(.A(mai_mai_n69_), .B(mai_mai_n55_), .Y(mai_mai_n609_));
  NA2        m0560(.A(mai_mai_n609_), .B(mai_mai_n608_), .Y(mai_mai_n610_));
  NA2        m0561(.A(mai_mai_n610_), .B(mai_mai_n607_), .Y(mai_mai_n611_));
  OAI210     m0562(.A0(mai_mai_n611_), .A1(mai_mai_n603_), .B0(mai_mai_n598_), .Y(mai_mai_n612_));
  NO2        m0563(.A(mai_mai_n67_), .B(mai_mai_n50_), .Y(mai_mai_n613_));
  NO2        m0564(.A(mai_mai_n182_), .B(x4), .Y(mai_mai_n614_));
  NO2        m0565(.A(x5), .B(mai_mai_n56_), .Y(mai_mai_n615_));
  XO2        m0566(.A(x5), .B(x2), .Y(mai_mai_n616_));
  NO3        m0567(.A(x8), .B(x7), .C(mai_mai_n98_), .Y(mai_mai_n617_));
  AO220      m0568(.A0(mai_mai_n617_), .A1(mai_mai_n615_), .B0(mai_mai_n616_), .B1(mai_mai_n614_), .Y(mai_mai_n618_));
  NA3        m0569(.A(mai_mai_n618_), .B(mai_mai_n613_), .C(mai_mai_n53_), .Y(mai_mai_n619_));
  NA2        m0570(.A(mai_mai_n256_), .B(mai_mai_n573_), .Y(mai_mai_n620_));
  NOi21      m0571(.An(x4), .B(x1), .Y(mai_mai_n621_));
  NA2        m0572(.A(mai_mai_n621_), .B(mai_mai_n62_), .Y(mai_mai_n622_));
  NA2        m0573(.A(x4), .B(x1), .Y(mai_mai_n623_));
  NO2        m0574(.A(mai_mai_n623_), .B(mai_mai_n50_), .Y(mai_mai_n624_));
  AOI210     m0575(.A0(mai_mai_n624_), .A1(mai_mai_n600_), .B0(mai_mai_n59_), .Y(mai_mai_n625_));
  OA210      m0576(.A0(mai_mai_n622_), .A1(mai_mai_n620_), .B0(mai_mai_n625_), .Y(mai_mai_n626_));
  NA4        m0577(.A(mai_mai_n626_), .B(mai_mai_n619_), .C(mai_mai_n612_), .D(mai_mai_n597_), .Y(mai_mai_n627_));
  NA2        m0578(.A(mai_mai_n613_), .B(mai_mai_n56_), .Y(mai_mai_n628_));
  NA2        m0579(.A(mai_mai_n554_), .B(mai_mai_n587_), .Y(mai_mai_n629_));
  NO2        m0580(.A(mai_mai_n629_), .B(mai_mai_n628_), .Y(mai_mai_n630_));
  NA2        m0581(.A(mai_mai_n259_), .B(mai_mai_n111_), .Y(mai_mai_n631_));
  OAI210     m0582(.A0(mai_mai_n631_), .A1(mai_mai_n154_), .B0(mai_mai_n59_), .Y(mai_mai_n632_));
  NA2        m0583(.A(mai_mai_n57_), .B(x6), .Y(mai_mai_n633_));
  AOI210     m0584(.A0(mai_mai_n633_), .A1(x3), .B0(mai_mai_n83_), .Y(mai_mai_n634_));
  NA2        m0585(.A(mai_mai_n615_), .B(mai_mai_n145_), .Y(mai_mai_n635_));
  NO3        m0586(.A(mai_mai_n635_), .B(mai_mai_n634_), .C(mai_mai_n415_), .Y(mai_mai_n636_));
  NA2        m0587(.A(mai_mai_n268_), .B(mai_mai_n67_), .Y(mai_mai_n637_));
  NO2        m0588(.A(mai_mai_n376_), .B(x3), .Y(mai_mai_n638_));
  NO2        m0589(.A(mai_mai_n415_), .B(mai_mai_n614_), .Y(mai_mai_n639_));
  NO2        m0590(.A(mai_mai_n456_), .B(mai_mai_n96_), .Y(mai_mai_n640_));
  NO2        m0591(.A(mai_mai_n564_), .B(x6), .Y(mai_mai_n641_));
  NA2        m0592(.A(mai_mai_n641_), .B(mai_mai_n640_), .Y(mai_mai_n642_));
  NO2        m0593(.A(mai_mai_n642_), .B(mai_mai_n639_), .Y(mai_mai_n643_));
  NO4        m0594(.A(mai_mai_n643_), .B(mai_mai_n636_), .C(mai_mai_n632_), .D(mai_mai_n630_), .Y(mai_mai_n644_));
  NA2        m0595(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n645_));
  NO2        m0596(.A(mai_mai_n645_), .B(x1), .Y(mai_mai_n646_));
  NA2        m0597(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n647_));
  NA2        m0598(.A(x8), .B(x4), .Y(mai_mai_n648_));
  NO2        m0599(.A(x8), .B(x4), .Y(mai_mai_n649_));
  NAi21      m0600(.An(mai_mai_n649_), .B(mai_mai_n648_), .Y(mai_mai_n650_));
  NAi21      m0601(.An(mai_mai_n554_), .B(mai_mai_n376_), .Y(mai_mai_n651_));
  NO3        m0602(.A(x8), .B(mai_mai_n96_), .C(x4), .Y(mai_mai_n652_));
  INV        m0603(.A(mai_mai_n652_), .Y(mai_mai_n653_));
  NO2        m0604(.A(mai_mai_n653_), .B(mai_mai_n98_), .Y(mai_mai_n654_));
  NO2        m0605(.A(x5), .B(x4), .Y(mai_mai_n655_));
  NA3        m0606(.A(mai_mai_n655_), .B(mai_mai_n62_), .C(mai_mai_n98_), .Y(mai_mai_n656_));
  NO2        m0607(.A(x6), .B(mai_mai_n98_), .Y(mai_mai_n657_));
  INV        m0608(.A(mai_mai_n656_), .Y(mai_mai_n658_));
  OAI210     m0609(.A0(mai_mai_n658_), .A1(mai_mai_n654_), .B0(mai_mai_n298_), .Y(mai_mai_n659_));
  NA2        m0610(.A(mai_mai_n659_), .B(mai_mai_n644_), .Y(mai_mai_n660_));
  OR2        m0611(.A(x4), .B(x1), .Y(mai_mai_n661_));
  NO2        m0612(.A(mai_mai_n661_), .B(x3), .Y(mai_mai_n662_));
  NA2        m0613(.A(mai_mai_n55_), .B(x2), .Y(mai_mai_n663_));
  NO3        m0614(.A(mai_mai_n357_), .B(mai_mai_n663_), .C(x6), .Y(mai_mai_n664_));
  AOI220     m0615(.A0(mai_mai_n664_), .A1(mai_mai_n662_), .B0(mai_mai_n660_), .B1(mai_mai_n627_), .Y(mai06));
  NA2        m0616(.A(mai_mai_n56_), .B(x3), .Y(mai_mai_n666_));
  NA2        m0617(.A(x6), .B(mai_mai_n98_), .Y(mai_mai_n667_));
  NA2        m0618(.A(mai_mai_n667_), .B(mai_mai_n55_), .Y(mai_mai_n668_));
  NA2        m0619(.A(x5), .B(mai_mai_n59_), .Y(mai_mai_n669_));
  NO2        m0620(.A(mai_mai_n669_), .B(mai_mai_n106_), .Y(mai_mai_n670_));
  NA3        m0621(.A(mai_mai_n670_), .B(mai_mai_n668_), .C(mai_mai_n488_), .Y(mai_mai_n671_));
  NO2        m0622(.A(mai_mai_n376_), .B(x0), .Y(mai_mai_n672_));
  NA2        m0623(.A(mai_mai_n327_), .B(x2), .Y(mai_mai_n673_));
  NOi21      m0624(.An(x6), .B(x8), .Y(mai_mai_n674_));
  NO2        m0625(.A(mai_mai_n674_), .B(x2), .Y(mai_mai_n675_));
  NO3        m0626(.A(mai_mai_n675_), .B(mai_mai_n66_), .C(mai_mai_n59_), .Y(mai_mai_n676_));
  AOI220     m0627(.A0(mai_mai_n676_), .A1(mai_mai_n673_), .B0(mai_mai_n672_), .B1(mai_mai_n319_), .Y(mai_mai_n677_));
  AOI210     m0628(.A0(mai_mai_n677_), .A1(mai_mai_n671_), .B0(mai_mai_n666_), .Y(mai_mai_n678_));
  NA2        m0629(.A(mai_mai_n56_), .B(mai_mai_n50_), .Y(mai_mai_n679_));
  NA2        m0630(.A(mai_mai_n355_), .B(mai_mai_n343_), .Y(mai_mai_n680_));
  NO2        m0631(.A(mai_mai_n67_), .B(mai_mai_n96_), .Y(mai_mai_n681_));
  NO2        m0632(.A(mai_mai_n53_), .B(mai_mai_n59_), .Y(mai_mai_n682_));
  NO2        m0633(.A(mai_mai_n663_), .B(mai_mai_n681_), .Y(mai_mai_n683_));
  AOI220     m0634(.A0(mai_mai_n683_), .A1(mai_mai_n680_), .B0(mai_mai_n412_), .B1(mai_mai_n62_), .Y(mai_mai_n684_));
  NO2        m0635(.A(mai_mai_n684_), .B(mai_mai_n679_), .Y(mai_mai_n685_));
  NO2        m0636(.A(mai_mai_n54_), .B(x0), .Y(mai_mai_n686_));
  NA2        m0637(.A(x4), .B(x3), .Y(mai_mai_n687_));
  NO2        m0638(.A(mai_mai_n94_), .B(mai_mai_n56_), .Y(mai_mai_n688_));
  NO2        m0639(.A(x5), .B(x3), .Y(mai_mai_n689_));
  NA2        m0640(.A(mai_mai_n588_), .B(mai_mai_n545_), .Y(mai_mai_n690_));
  OR2        m0641(.A(mai_mai_n690_), .B(mai_mai_n567_), .Y(mai_mai_n691_));
  INV        m0642(.A(mai_mai_n691_), .Y(mai_mai_n692_));
  OR3        m0643(.A(mai_mai_n692_), .B(mai_mai_n685_), .C(mai_mai_n678_), .Y(mai_mai_n693_));
  NA2        m0644(.A(x7), .B(mai_mai_n56_), .Y(mai_mai_n694_));
  NO2        m0645(.A(mai_mai_n600_), .B(mai_mai_n59_), .Y(mai_mai_n695_));
  NA2        m0646(.A(mai_mai_n695_), .B(mai_mai_n613_), .Y(mai_mai_n696_));
  NO2        m0647(.A(mai_mai_n160_), .B(x6), .Y(mai_mai_n697_));
  NA2        m0648(.A(mai_mai_n697_), .B(mai_mai_n277_), .Y(mai_mai_n698_));
  AOI210     m0649(.A0(mai_mai_n698_), .A1(mai_mai_n696_), .B0(mai_mai_n694_), .Y(mai_mai_n699_));
  AN2        m0650(.A(mai_mai_n461_), .B(mai_mai_n309_), .Y(mai_mai_n700_));
  OAI210     m0651(.A0(mai_mai_n700_), .A1(mai_mai_n699_), .B0(mai_mai_n338_), .Y(mai_mai_n701_));
  NO2        m0652(.A(mai_mai_n294_), .B(mai_mai_n96_), .Y(mai_mai_n702_));
  NO2        m0653(.A(mai_mai_n56_), .B(x3), .Y(mai_mai_n703_));
  NA2        m0654(.A(mai_mai_n703_), .B(mai_mai_n67_), .Y(mai_mai_n704_));
  NO2        m0655(.A(mai_mai_n704_), .B(mai_mai_n237_), .Y(mai_mai_n705_));
  NO2        m0656(.A(mai_mai_n67_), .B(x3), .Y(mai_mai_n706_));
  NO2        m0657(.A(mai_mai_n57_), .B(x6), .Y(mai_mai_n707_));
  NA2        m0658(.A(mai_mai_n171_), .B(mai_mai_n707_), .Y(mai_mai_n708_));
  NA3        m0659(.A(mai_mai_n588_), .B(mai_mai_n316_), .C(mai_mai_n67_), .Y(mai_mai_n709_));
  NA2        m0660(.A(mai_mai_n709_), .B(mai_mai_n708_), .Y(mai_mai_n710_));
  OR3        m0661(.A(mai_mai_n710_), .B(mai_mai_n705_), .C(mai_mai_n624_), .Y(mai_mai_n711_));
  NA2        m0662(.A(mai_mai_n711_), .B(mai_mai_n702_), .Y(mai_mai_n712_));
  NA2        m0663(.A(mai_mai_n686_), .B(mai_mai_n613_), .Y(mai_mai_n713_));
  NA4        m0664(.A(mai_mai_n252_), .B(mai_mai_n574_), .C(mai_mai_n210_), .D(mai_mai_n244_), .Y(mai_mai_n714_));
  NA2        m0665(.A(mai_mai_n472_), .B(mai_mai_n64_), .Y(mai_mai_n715_));
  AOI210     m0666(.A0(mai_mai_n714_), .A1(mai_mai_n713_), .B0(mai_mai_n715_), .Y(mai_mai_n716_));
  NA2        m0667(.A(x7), .B(x6), .Y(mai_mai_n717_));
  NA3        m0668(.A(x2), .B(x1), .C(x0), .Y(mai_mai_n718_));
  NA2        m0669(.A(mai_mai_n484_), .B(mai_mai_n139_), .Y(mai_mai_n719_));
  NO2        m0670(.A(x5), .B(x1), .Y(mai_mai_n720_));
  NA2        m0671(.A(mai_mai_n720_), .B(mai_mai_n707_), .Y(mai_mai_n721_));
  NA2        m0672(.A(x4), .B(x0), .Y(mai_mai_n722_));
  NO3        m0673(.A(mai_mai_n57_), .B(x6), .C(x2), .Y(mai_mai_n723_));
  NA2        m0674(.A(mai_mai_n723_), .B(mai_mai_n213_), .Y(mai_mai_n724_));
  OAI220     m0675(.A0(mai_mai_n724_), .A1(mai_mai_n722_), .B0(mai_mai_n721_), .B1(mai_mai_n719_), .Y(mai_mai_n725_));
  NO2        m0676(.A(mai_mai_n725_), .B(mai_mai_n716_), .Y(mai_mai_n726_));
  NA3        m0677(.A(mai_mai_n726_), .B(mai_mai_n712_), .C(mai_mai_n701_), .Y(mai_mai_n727_));
  AOI210     m0678(.A0(mai_mai_n693_), .A1(mai_mai_n57_), .B0(mai_mai_n727_), .Y(mai07));
  NA2        m0679(.A(mai_mai_n96_), .B(mai_mai_n59_), .Y(mai_mai_n729_));
  NOi21      m0680(.An(mai_mai_n717_), .B(mai_mai_n104_), .Y(mai_mai_n730_));
  NO4        m0681(.A(mai_mai_n730_), .B(mai_mai_n613_), .C(mai_mai_n237_), .D(mai_mai_n729_), .Y(mai_mai_n731_));
  NO3        m0682(.A(mai_mai_n57_), .B(x5), .C(x1), .Y(mai_mai_n732_));
  NA2        m0683(.A(mai_mai_n732_), .B(mai_mai_n363_), .Y(mai_mai_n733_));
  NO2        m0684(.A(mai_mai_n57_), .B(mai_mai_n67_), .Y(mai_mai_n734_));
  NO2        m0685(.A(mai_mai_n144_), .B(mai_mai_n97_), .Y(mai_mai_n735_));
  AOI210     m0686(.A0(mai_mai_n734_), .A1(mai_mai_n84_), .B0(mai_mai_n735_), .Y(mai_mai_n736_));
  OAI220     m0687(.A0(mai_mai_n736_), .A1(mai_mai_n125_), .B0(mai_mai_n733_), .B1(mai_mai_n311_), .Y(mai_mai_n737_));
  OAI210     m0688(.A0(mai_mai_n737_), .A1(mai_mai_n731_), .B0(x2), .Y(mai_mai_n738_));
  NAi21      m0689(.An(mai_mai_n145_), .B(mai_mai_n146_), .Y(mai_mai_n739_));
  NA3        m0690(.A(mai_mai_n739_), .B(mai_mai_n83_), .C(x3), .Y(mai_mai_n740_));
  NO3        m0691(.A(mai_mai_n55_), .B(x3), .C(x1), .Y(mai_mai_n741_));
  NO2        m0692(.A(mai_mai_n501_), .B(x2), .Y(mai_mai_n742_));
  NA2        m0693(.A(mai_mai_n742_), .B(mai_mai_n503_), .Y(mai_mai_n743_));
  OAI210     m0694(.A0(mai_mai_n743_), .A1(mai_mai_n633_), .B0(mai_mai_n740_), .Y(mai_mai_n744_));
  NO2        m0695(.A(x8), .B(mai_mai_n53_), .Y(mai_mai_n745_));
  NA2        m0696(.A(mai_mai_n745_), .B(mai_mai_n59_), .Y(mai_mai_n746_));
  NA2        m0697(.A(mai_mai_n344_), .B(mai_mai_n338_), .Y(mai_mai_n747_));
  NO2        m0698(.A(x7), .B(x3), .Y(mai_mai_n748_));
  NA2        m0699(.A(mai_mai_n748_), .B(mai_mai_n92_), .Y(mai_mai_n749_));
  AOI210     m0700(.A0(mai_mai_n747_), .A1(mai_mai_n746_), .B0(mai_mai_n749_), .Y(mai_mai_n750_));
  AOI210     m0701(.A0(mai_mai_n744_), .A1(mai_mai_n236_), .B0(mai_mai_n750_), .Y(mai_mai_n751_));
  AOI210     m0702(.A0(mai_mai_n751_), .A1(mai_mai_n738_), .B0(x4), .Y(mai_mai_n752_));
  NA3        m0703(.A(mai_mai_n720_), .B(mai_mai_n307_), .C(mai_mai_n55_), .Y(mai_mai_n753_));
  AOI210     m0704(.A0(mai_mai_n753_), .A1(mai_mai_n583_), .B0(mai_mai_n98_), .Y(mai_mai_n754_));
  XO2        m0705(.A(x5), .B(x1), .Y(mai_mai_n755_));
  NA2        m0706(.A(mai_mai_n754_), .B(mai_mai_n403_), .Y(mai_mai_n756_));
  NO3        m0707(.A(mai_mai_n50_), .B(x2), .C(x0), .Y(mai_mai_n757_));
  NA2        m0708(.A(x6), .B(x0), .Y(mai_mai_n758_));
  NO2        m0709(.A(mai_mai_n663_), .B(mai_mai_n758_), .Y(mai_mai_n759_));
  NO2        m0710(.A(mai_mai_n756_), .B(mai_mai_n56_), .Y(mai_mai_n760_));
  NOi21      m0711(.An(mai_mai_n217_), .B(mai_mai_n363_), .Y(mai_mai_n761_));
  NO3        m0712(.A(mai_mai_n761_), .B(mai_mai_n226_), .C(mai_mai_n64_), .Y(mai_mai_n762_));
  NO2        m0713(.A(mai_mai_n180_), .B(mai_mai_n67_), .Y(mai_mai_n763_));
  NO2        m0714(.A(mai_mai_n297_), .B(x6), .Y(mai_mai_n764_));
  AO220      m0715(.A0(mai_mai_n764_), .A1(mai_mai_n317_), .B0(mai_mai_n763_), .B1(mai_mai_n546_), .Y(mai_mai_n765_));
  OAI210     m0716(.A0(mai_mai_n765_), .A1(mai_mai_n762_), .B0(mai_mai_n59_), .Y(mai_mai_n766_));
  NA2        m0717(.A(mai_mai_n84_), .B(mai_mai_n67_), .Y(mai_mai_n767_));
  NAi21      m0718(.An(x8), .B(x7), .Y(mai_mai_n768_));
  NA2        m0719(.A(mai_mai_n761_), .B(mai_mai_n768_), .Y(mai_mai_n769_));
  NA2        m0720(.A(mai_mai_n396_), .B(mai_mai_n98_), .Y(mai_mai_n770_));
  NO2        m0721(.A(mai_mai_n674_), .B(x1), .Y(mai_mai_n771_));
  NO2        m0722(.A(mai_mai_n766_), .B(mai_mai_n132_), .Y(mai_mai_n772_));
  NO2        m0723(.A(x8), .B(x7), .Y(mai_mai_n773_));
  NO2        m0724(.A(mai_mai_n773_), .B(x3), .Y(mai_mai_n774_));
  NA3        m0725(.A(mai_mai_n774_), .B(mai_mai_n352_), .C(x1), .Y(mai_mai_n775_));
  NO2        m0726(.A(x8), .B(mai_mai_n98_), .Y(mai_mai_n776_));
  AOI220     m0727(.A0(mai_mai_n316_), .A1(mai_mai_n338_), .B0(mai_mai_n776_), .B1(mai_mai_n241_), .Y(mai_mai_n777_));
  NO2        m0728(.A(mai_mai_n67_), .B(x4), .Y(mai_mai_n778_));
  NA2        m0729(.A(mai_mai_n778_), .B(mai_mai_n291_), .Y(mai_mai_n779_));
  AOI210     m0730(.A0(mai_mai_n777_), .A1(mai_mai_n775_), .B0(mai_mai_n779_), .Y(mai_mai_n780_));
  NO4        m0731(.A(mai_mai_n780_), .B(mai_mai_n772_), .C(mai_mai_n760_), .D(mai_mai_n752_), .Y(mai08));
  NA2        m0732(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n782_));
  XN2        m0733(.A(x5), .B(x4), .Y(mai_mai_n783_));
  INV        m0734(.A(mai_mai_n783_), .Y(mai_mai_n784_));
  AOI220     m0735(.A0(mai_mai_n784_), .A1(mai_mai_n344_), .B0(mai_mai_n128_), .B1(mai_mai_n56_), .Y(mai_mai_n785_));
  NO2        m0736(.A(mai_mai_n228_), .B(mai_mai_n96_), .Y(mai_mai_n786_));
  AOI210     m0737(.A0(mai_mai_n786_), .A1(mai_mai_n265_), .B0(mai_mai_n181_), .Y(mai_mai_n787_));
  OAI220     m0738(.A0(mai_mai_n787_), .A1(x4), .B0(mai_mai_n785_), .B1(mai_mai_n782_), .Y(mai_mai_n788_));
  NA2        m0739(.A(mai_mai_n788_), .B(mai_mai_n259_), .Y(mai_mai_n789_));
  NO2        m0740(.A(mai_mai_n258_), .B(mai_mai_n599_), .Y(mai_mai_n790_));
  NA2        m0741(.A(mai_mai_n594_), .B(mai_mai_n160_), .Y(mai_mai_n791_));
  OAI220     m0742(.A0(mai_mai_n791_), .A1(mai_mai_n647_), .B0(mai_mai_n474_), .B1(mai_mai_n50_), .Y(mai_mai_n792_));
  AO210      m0743(.A0(mai_mai_n792_), .A1(mai_mai_n331_), .B0(mai_mai_n790_), .Y(mai_mai_n793_));
  NA2        m0744(.A(mai_mai_n265_), .B(mai_mai_n139_), .Y(mai_mai_n794_));
  NA2        m0745(.A(mai_mai_n132_), .B(x7), .Y(mai_mai_n795_));
  NO2        m0746(.A(mai_mai_n794_), .B(mai_mai_n194_), .Y(mai_mai_n796_));
  AOI210     m0747(.A0(mai_mai_n793_), .A1(mai_mai_n279_), .B0(mai_mai_n796_), .Y(mai_mai_n797_));
  AOI210     m0748(.A0(mai_mai_n797_), .A1(mai_mai_n789_), .B0(mai_mai_n67_), .Y(mai_mai_n798_));
  NO2        m0749(.A(mai_mai_n773_), .B(mai_mai_n98_), .Y(mai_mai_n799_));
  NA2        m0750(.A(mai_mai_n799_), .B(mai_mai_n182_), .Y(mai_mai_n800_));
  OAI210     m0751(.A0(mai_mai_n399_), .A1(mai_mai_n291_), .B0(mai_mai_n331_), .Y(mai_mai_n801_));
  NA2        m0752(.A(mai_mai_n425_), .B(mai_mai_n219_), .Y(mai_mai_n802_));
  NO2        m0753(.A(mai_mai_n801_), .B(mai_mai_n800_), .Y(mai_mai_n803_));
  NA2        m0754(.A(mai_mai_n803_), .B(mai_mai_n275_), .Y(mai_mai_n804_));
  NA2        m0755(.A(mai_mai_n321_), .B(mai_mai_n53_), .Y(mai_mai_n805_));
  NO2        m0756(.A(mai_mai_n682_), .B(mai_mai_n231_), .Y(mai_mai_n806_));
  NO3        m0757(.A(mai_mai_n555_), .B(mai_mai_n457_), .C(mai_mai_n90_), .Y(mai_mai_n807_));
  AN2        m0758(.A(mai_mai_n807_), .B(mai_mai_n806_), .Y(mai_mai_n808_));
  NA2        m0759(.A(x7), .B(mai_mai_n59_), .Y(mai_mai_n809_));
  NO3        m0760(.A(mai_mai_n300_), .B(mai_mai_n809_), .C(mai_mai_n274_), .Y(mai_mai_n810_));
  AOI210     m0761(.A0(mai_mai_n808_), .A1(x5), .B0(mai_mai_n810_), .Y(mai_mai_n811_));
  AOI210     m0762(.A0(mai_mai_n811_), .A1(mai_mai_n804_), .B0(mai_mai_n68_), .Y(mai_mai_n812_));
  NO2        m0763(.A(mai_mai_n66_), .B(x3), .Y(mai_mai_n813_));
  OAI210     m0764(.A0(mai_mai_n813_), .A1(mai_mai_n250_), .B0(mai_mai_n137_), .Y(mai_mai_n814_));
  MUX2       m0765(.S(x3), .A(mai_mai_n153_), .B(mai_mai_n739_), .Y(mai_mai_n815_));
  NA2        m0766(.A(mai_mai_n815_), .B(mai_mai_n546_), .Y(mai_mai_n816_));
  NO3        m0767(.A(x6), .B(x4), .C(x0), .Y(mai_mai_n817_));
  INV        m0768(.A(mai_mai_n817_), .Y(mai_mai_n818_));
  AOI210     m0769(.A0(mai_mai_n816_), .A1(mai_mai_n814_), .B0(mai_mai_n818_), .Y(mai_mai_n819_));
  NO3        m0770(.A(x5), .B(x3), .C(mai_mai_n98_), .Y(mai_mai_n820_));
  NA2        m0771(.A(mai_mai_n784_), .B(mai_mai_n296_), .Y(mai_mai_n821_));
  OR2        m0772(.A(x8), .B(x1), .Y(mai_mai_n822_));
  NO3        m0773(.A(mai_mai_n822_), .B(mai_mai_n821_), .C(mai_mai_n703_), .Y(mai_mai_n823_));
  NAi21      m0774(.An(x4), .B(x1), .Y(mai_mai_n824_));
  NA3        m0775(.A(mai_mai_n55_), .B(x1), .C(x0), .Y(mai_mai_n825_));
  NA2        m0776(.A(mai_mai_n823_), .B(mai_mai_n307_), .Y(mai_mai_n826_));
  BUFFER     m0777(.A(mai_mai_n702_), .Y(mai_mai_n827_));
  NA2        m0778(.A(mai_mai_n96_), .B(mai_mai_n56_), .Y(mai_mai_n828_));
  NO2        m0779(.A(mai_mai_n828_), .B(mai_mai_n246_), .Y(mai_mai_n829_));
  NO2        m0780(.A(mai_mai_n57_), .B(x2), .Y(mai_mai_n830_));
  NO4        m0781(.A(mai_mai_n317_), .B(mai_mai_n830_), .C(mai_mai_n773_), .D(mai_mai_n281_), .Y(mai_mai_n831_));
  AOI220     m0782(.A0(mai_mai_n831_), .A1(mai_mai_n829_), .B0(mai_mai_n827_), .B1(mai_mai_n624_), .Y(mai_mai_n832_));
  NA2        m0783(.A(mai_mai_n832_), .B(mai_mai_n826_), .Y(mai_mai_n833_));
  NO4        m0784(.A(mai_mai_n833_), .B(mai_mai_n819_), .C(mai_mai_n812_), .D(mai_mai_n798_), .Y(mai09));
  NO3        m0785(.A(mai_mai_n755_), .B(mai_mai_n109_), .C(mai_mai_n88_), .Y(mai_mai_n835_));
  AOI220     m0786(.A0(mai_mai_n286_), .A1(mai_mai_n66_), .B0(mai_mai_n573_), .B1(mai_mai_n528_), .Y(mai_mai_n836_));
  OAI210     m0787(.A0(mai_mai_n835_), .A1(x2), .B0(mai_mai_n836_), .Y(mai_mai_n837_));
  AOI210     m0788(.A0(mai_mai_n837_), .A1(mai_mai_n721_), .B0(mai_mai_n434_), .Y(mai_mai_n838_));
  NO2        m0789(.A(mai_mai_n572_), .B(mai_mai_n249_), .Y(mai_mai_n839_));
  NO2        m0790(.A(mai_mai_n720_), .B(mai_mai_n327_), .Y(mai_mai_n840_));
  NO3        m0791(.A(mai_mai_n587_), .B(mai_mai_n93_), .C(mai_mai_n98_), .Y(mai_mai_n841_));
  AO220      m0792(.A0(mai_mai_n841_), .A1(mai_mai_n840_), .B0(mai_mai_n839_), .B1(mai_mai_n600_), .Y(mai_mai_n842_));
  OAI210     m0793(.A0(mai_mai_n842_), .A1(mai_mai_n838_), .B0(x4), .Y(mai_mai_n843_));
  OAI220     m0794(.A0(mai_mai_n355_), .A1(mai_mai_n134_), .B0(mai_mai_n383_), .B1(mai_mai_n267_), .Y(mai_mai_n844_));
  NO2        m0795(.A(mai_mai_n180_), .B(mai_mai_n96_), .Y(mai_mai_n845_));
  AOI220     m0796(.A0(mai_mai_n845_), .A1(mai_mai_n114_), .B0(mai_mai_n844_), .B1(mai_mai_n606_), .Y(mai_mai_n846_));
  NAi21      m0797(.An(x0), .B(x2), .Y(mai_mai_n847_));
  NO2        m0798(.A(mai_mai_n290_), .B(mai_mai_n847_), .Y(mai_mai_n848_));
  OAI210     m0799(.A0(mai_mai_n466_), .A1(mai_mai_n262_), .B0(mai_mai_n180_), .Y(mai_mai_n849_));
  AOI210     m0800(.A0(mai_mai_n156_), .A1(mai_mai_n768_), .B0(mai_mai_n343_), .Y(mai_mai_n850_));
  NA2        m0801(.A(mai_mai_n850_), .B(mai_mai_n849_), .Y(mai_mai_n851_));
  OAI210     m0802(.A0(mai_mai_n846_), .A1(mai_mai_n55_), .B0(mai_mai_n851_), .Y(mai_mai_n852_));
  NA2        m0803(.A(mai_mai_n852_), .B(mai_mai_n56_), .Y(mai_mai_n853_));
  NO2        m0804(.A(mai_mai_n56_), .B(mai_mai_n59_), .Y(mai_mai_n854_));
  INV        m0805(.A(mai_mai_n114_), .Y(mai_mai_n855_));
  NA2        m0806(.A(mai_mai_n720_), .B(mai_mai_n55_), .Y(mai_mai_n856_));
  AOI210     m0807(.A0(x6), .A1(x1), .B0(x5), .Y(mai_mai_n857_));
  OAI210     m0808(.A0(mai_mai_n857_), .A1(mai_mai_n320_), .B0(x2), .Y(mai_mai_n858_));
  AOI210     m0809(.A0(mai_mai_n858_), .A1(mai_mai_n856_), .B0(mai_mai_n855_), .Y(mai_mai_n859_));
  NA2        m0810(.A(mai_mai_n545_), .B(mai_mai_n55_), .Y(mai_mai_n860_));
  NO4        m0811(.A(mai_mai_n57_), .B(x6), .C(x5), .D(x1), .Y(mai_mai_n861_));
  NO2        m0812(.A(mai_mai_n216_), .B(mai_mai_n373_), .Y(mai_mai_n862_));
  NO2        m0813(.A(mai_mai_n297_), .B(mai_mai_n138_), .Y(mai_mai_n863_));
  NO3        m0814(.A(mai_mai_n863_), .B(mai_mai_n862_), .C(mai_mai_n861_), .Y(mai_mai_n864_));
  OAI220     m0815(.A0(mai_mai_n864_), .A1(mai_mai_n55_), .B0(mai_mai_n860_), .B1(mai_mai_n445_), .Y(mai_mai_n865_));
  OAI210     m0816(.A0(mai_mai_n865_), .A1(mai_mai_n859_), .B0(mai_mai_n854_), .Y(mai_mai_n866_));
  NO2        m0817(.A(mai_mai_n392_), .B(mai_mai_n96_), .Y(mai_mai_n867_));
  NO2        m0818(.A(mai_mai_n321_), .B(mai_mai_n483_), .Y(mai_mai_n868_));
  AOI220     m0819(.A0(mai_mai_n868_), .A1(mai_mai_n867_), .B0(mai_mai_n198_), .B1(mai_mai_n214_), .Y(mai_mai_n869_));
  NA4        m0820(.A(mai_mai_n869_), .B(mai_mai_n866_), .C(mai_mai_n853_), .D(mai_mai_n843_), .Y(mai_mai_n870_));
  NA2        m0821(.A(mai_mai_n870_), .B(mai_mai_n50_), .Y(mai_mai_n871_));
  NO2        m0822(.A(mai_mai_n366_), .B(mai_mai_n149_), .Y(mai_mai_n872_));
  NA2        m0823(.A(mai_mai_n225_), .B(mai_mai_n573_), .Y(mai_mai_n873_));
  OAI210     m0824(.A0(mai_mai_n420_), .A1(mai_mai_n776_), .B0(mai_mai_n873_), .Y(mai_mai_n874_));
  OAI210     m0825(.A0(mai_mai_n874_), .A1(mai_mai_n872_), .B0(x0), .Y(mai_mai_n875_));
  NO3        m0826(.A(x8), .B(x7), .C(x2), .Y(mai_mai_n876_));
  NO3        m0827(.A(mai_mai_n57_), .B(x5), .C(x2), .Y(mai_mai_n877_));
  OAI210     m0828(.A0(mai_mai_n877_), .A1(mai_mai_n876_), .B0(mai_mai_n503_), .Y(mai_mai_n878_));
  AOI210     m0829(.A0(mai_mai_n878_), .A1(mai_mai_n875_), .B0(x4), .Y(mai_mai_n879_));
  NO2        m0830(.A(mai_mai_n413_), .B(mai_mai_n137_), .Y(mai_mai_n880_));
  NO2        m0831(.A(mai_mai_n52_), .B(x2), .Y(mai_mai_n881_));
  NO2        m0832(.A(mai_mai_n96_), .B(mai_mai_n56_), .Y(mai_mai_n882_));
  NA2        m0833(.A(mai_mai_n882_), .B(x8), .Y(mai_mai_n883_));
  NA2        m0834(.A(mai_mai_n883_), .B(mai_mai_n856_), .Y(mai_mai_n884_));
  AO210      m0835(.A0(mai_mai_n884_), .A1(mai_mai_n881_), .B0(mai_mai_n880_), .Y(mai_mai_n885_));
  OAI210     m0836(.A0(mai_mai_n885_), .A1(mai_mai_n879_), .B0(mai_mai_n598_), .Y(mai_mai_n886_));
  NO2        m0837(.A(mai_mai_n245_), .B(mai_mai_n107_), .Y(mai_mai_n887_));
  OAI210     m0838(.A0(x4), .A1(x2), .B0(x0), .Y(mai_mai_n888_));
  NA3        m0839(.A(mai_mai_n589_), .B(mai_mai_n599_), .C(mai_mai_n332_), .Y(mai_mai_n889_));
  OAI210     m0840(.A0(mai_mai_n888_), .A1(mai_mai_n274_), .B0(mai_mai_n53_), .Y(mai_mai_n890_));
  AOI210     m0841(.A0(mai_mai_n889_), .A1(mai_mai_n888_), .B0(mai_mai_n890_), .Y(mai_mai_n891_));
  OAI210     m0842(.A0(mai_mai_n891_), .A1(mai_mai_n887_), .B0(mai_mai_n316_), .Y(mai_mai_n892_));
  AOI220     m0843(.A0(mai_mai_n648_), .A1(mai_mai_n336_), .B0(mai_mai_n338_), .B1(mai_mai_n85_), .Y(mai_mai_n893_));
  NA2        m0844(.A(mai_mai_n85_), .B(x5), .Y(mai_mai_n894_));
  OAI220     m0845(.A0(mai_mai_n894_), .A1(mai_mai_n822_), .B0(mai_mai_n893_), .B1(mai_mai_n308_), .Y(mai_mai_n895_));
  NA2        m0846(.A(mai_mai_n895_), .B(mai_mai_n65_), .Y(mai_mai_n896_));
  NA2        m0847(.A(mai_mai_n396_), .B(mai_mai_n739_), .Y(mai_mai_n897_));
  NA2        m0848(.A(mai_mai_n236_), .B(mai_mai_n153_), .Y(mai_mai_n898_));
  AO210      m0849(.A0(mai_mai_n898_), .A1(mai_mai_n897_), .B0(mai_mai_n122_), .Y(mai_mai_n899_));
  NO2        m0850(.A(mai_mai_n426_), .B(x2), .Y(mai_mai_n900_));
  NO2        m0851(.A(x7), .B(mai_mai_n53_), .Y(mai_mai_n901_));
  NA2        m0852(.A(mai_mai_n649_), .B(mai_mai_n229_), .Y(mai_mai_n902_));
  NA4        m0853(.A(mai_mai_n902_), .B(mai_mai_n899_), .C(mai_mai_n896_), .D(mai_mai_n892_), .Y(mai_mai_n903_));
  NO4        m0854(.A(mai_mai_n889_), .B(mai_mai_n615_), .C(mai_mai_n445_), .D(mai_mai_n50_), .Y(mai_mai_n904_));
  AOI220     m0855(.A0(mai_mai_n588_), .A1(mai_mai_n587_), .B0(mai_mai_n268_), .B1(x5), .Y(mai_mai_n905_));
  NO2        m0856(.A(mai_mai_n655_), .B(mai_mai_n180_), .Y(mai_mai_n906_));
  NA3        m0857(.A(mai_mai_n906_), .B(mai_mai_n650_), .C(x7), .Y(mai_mai_n907_));
  OAI210     m0858(.A0(mai_mai_n905_), .A1(mai_mai_n337_), .B0(mai_mai_n907_), .Y(mai_mai_n908_));
  OAI210     m0859(.A0(mai_mai_n908_), .A1(mai_mai_n904_), .B0(mai_mai_n74_), .Y(mai_mai_n909_));
  NA2        m0860(.A(mai_mai_n745_), .B(x2), .Y(mai_mai_n910_));
  NO2        m0861(.A(mai_mai_n910_), .B(mai_mai_n58_), .Y(mai_mai_n911_));
  NO2        m0862(.A(x5), .B(mai_mai_n53_), .Y(mai_mai_n912_));
  NAi21      m0863(.An(x1), .B(x4), .Y(mai_mai_n913_));
  NA2        m0864(.A(mai_mai_n913_), .B(mai_mai_n824_), .Y(mai_mai_n914_));
  NO3        m0865(.A(mai_mai_n914_), .B(mai_mai_n191_), .C(mai_mai_n912_), .Y(mai_mai_n915_));
  OAI210     m0866(.A0(mai_mai_n915_), .A1(mai_mai_n911_), .B0(mai_mai_n403_), .Y(mai_mai_n916_));
  NA3        m0867(.A(mai_mai_n386_), .B(mai_mai_n720_), .C(mai_mai_n57_), .Y(mai_mai_n917_));
  NA3        m0868(.A(mai_mai_n917_), .B(mai_mai_n916_), .C(mai_mai_n909_), .Y(mai_mai_n918_));
  AOI210     m0869(.A0(mai_mai_n903_), .A1(x6), .B0(mai_mai_n918_), .Y(mai_mai_n919_));
  NA3        m0870(.A(mai_mai_n919_), .B(mai_mai_n886_), .C(mai_mai_n871_), .Y(mai10));
  NO2        m0871(.A(x4), .B(x1), .Y(mai_mai_n921_));
  NO2        m0872(.A(mai_mai_n921_), .B(mai_mai_n139_), .Y(mai_mai_n922_));
  NA3        m0873(.A(x5), .B(x4), .C(x0), .Y(mai_mai_n923_));
  NO2        m0874(.A(mai_mai_n923_), .B(mai_mai_n263_), .Y(mai_mai_n924_));
  NO2        m0875(.A(mai_mai_n2517_), .B(mai_mai_n290_), .Y(mai_mai_n925_));
  NOi21      m0876(.An(mai_mai_n244_), .B(mai_mai_n128_), .Y(mai_mai_n926_));
  AOI210     m0877(.A0(mai_mai_n489_), .A1(mai_mai_n600_), .B0(mai_mai_n317_), .Y(mai_mai_n927_));
  NO2        m0878(.A(mai_mai_n854_), .B(mai_mai_n330_), .Y(mai_mai_n928_));
  NOi31      m0879(.An(mai_mai_n928_), .B(mai_mai_n927_), .C(mai_mai_n926_), .Y(mai_mai_n929_));
  NA2        m0880(.A(x4), .B(mai_mai_n98_), .Y(mai_mai_n930_));
  NO2        m0881(.A(mai_mai_n311_), .B(mai_mai_n930_), .Y(mai_mai_n931_));
  NA2        m0882(.A(mai_mai_n90_), .B(x5), .Y(mai_mai_n932_));
  NO3        m0883(.A(mai_mai_n932_), .B(mai_mai_n99_), .C(mai_mai_n55_), .Y(mai_mai_n933_));
  NO3        m0884(.A(mai_mai_n933_), .B(mai_mai_n931_), .C(mai_mai_n929_), .Y(mai_mai_n934_));
  NA2        m0885(.A(mai_mai_n588_), .B(mai_mai_n257_), .Y(mai_mai_n935_));
  OAI220     m0886(.A0(mai_mai_n883_), .A1(mai_mai_n95_), .B0(mai_mai_n828_), .B1(mai_mai_n434_), .Y(mai_mai_n936_));
  NA2        m0887(.A(mai_mai_n936_), .B(mai_mai_n265_), .Y(mai_mai_n937_));
  OAI210     m0888(.A0(mai_mai_n934_), .A1(mai_mai_n373_), .B0(mai_mai_n937_), .Y(mai_mai_n938_));
  OAI210     m0889(.A0(mai_mai_n938_), .A1(mai_mai_n925_), .B0(x7), .Y(mai_mai_n939_));
  NA2        m0890(.A(mai_mai_n55_), .B(mai_mai_n67_), .Y(mai_mai_n940_));
  AOI210     m0891(.A0(mai_mai_n434_), .A1(mai_mai_n343_), .B0(mai_mai_n930_), .Y(mai_mai_n941_));
  NO3        m0892(.A(mai_mai_n436_), .B(mai_mai_n847_), .C(x5), .Y(mai_mai_n942_));
  OAI210     m0893(.A0(mai_mai_n942_), .A1(mai_mai_n941_), .B0(mai_mai_n940_), .Y(mai_mai_n943_));
  NO2        m0894(.A(mai_mai_n344_), .B(mai_mai_n131_), .Y(mai_mai_n944_));
  NA2        m0895(.A(mai_mai_n944_), .B(mai_mai_n414_), .Y(mai_mai_n945_));
  AOI210     m0896(.A0(mai_mai_n945_), .A1(mai_mai_n943_), .B0(x3), .Y(mai_mai_n946_));
  NO2        m0897(.A(x5), .B(mai_mai_n98_), .Y(mai_mai_n947_));
  OAI210     m0898(.A0(mai_mai_n947_), .A1(mai_mai_n223_), .B0(mai_mai_n894_), .Y(mai_mai_n948_));
  NO2        m0899(.A(mai_mai_n436_), .B(mai_mai_n203_), .Y(mai_mai_n949_));
  AOI210     m0900(.A0(mai_mai_n948_), .A1(mai_mai_n242_), .B0(mai_mai_n949_), .Y(mai_mai_n950_));
  NO2        m0901(.A(mai_mai_n950_), .B(mai_mai_n59_), .Y(mai_mai_n951_));
  OAI210     m0902(.A0(mai_mai_n951_), .A1(mai_mai_n946_), .B0(mai_mai_n901_), .Y(mai_mai_n952_));
  NO2        m0903(.A(x4), .B(x3), .Y(mai_mai_n953_));
  NO3        m0904(.A(mai_mai_n953_), .B(mai_mai_n331_), .C(mai_mai_n79_), .Y(mai_mai_n954_));
  OAI210     m0905(.A0(mai_mai_n954_), .A1(mai_mai_n264_), .B0(mai_mai_n425_), .Y(mai_mai_n955_));
  AOI210     m0906(.A0(mai_mai_n387_), .A1(mai_mai_n117_), .B0(mai_mai_n237_), .Y(mai_mai_n956_));
  NA2        m0907(.A(mai_mai_n921_), .B(mai_mai_n55_), .Y(mai_mai_n957_));
  NO2        m0908(.A(mai_mai_n957_), .B(mai_mai_n932_), .Y(mai_mai_n958_));
  NO2        m0909(.A(mai_mai_n513_), .B(mai_mai_n349_), .Y(mai_mai_n959_));
  NO3        m0910(.A(x4), .B(mai_mai_n98_), .C(mai_mai_n59_), .Y(mai_mai_n960_));
  NO2        m0911(.A(mai_mai_n426_), .B(x1), .Y(mai_mai_n961_));
  NOi31      m0912(.An(mai_mai_n960_), .B(mai_mai_n961_), .C(mai_mai_n959_), .Y(mai_mai_n962_));
  NA2        m0913(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n963_));
  NO4        m0914(.A(mai_mai_n922_), .B(mai_mai_n502_), .C(mai_mai_n963_), .D(x2), .Y(mai_mai_n964_));
  NO4        m0915(.A(mai_mai_n964_), .B(mai_mai_n962_), .C(mai_mai_n958_), .D(mai_mai_n956_), .Y(mai_mai_n965_));
  AOI210     m0916(.A0(mai_mai_n965_), .A1(mai_mai_n955_), .B0(mai_mai_n197_), .Y(mai_mai_n966_));
  NO2        m0917(.A(mai_mai_n647_), .B(mai_mai_n488_), .Y(mai_mai_n967_));
  NO2        m0918(.A(x6), .B(x2), .Y(mai_mai_n968_));
  NO3        m0919(.A(mai_mai_n968_), .B(mai_mai_n674_), .C(mai_mai_n60_), .Y(mai_mai_n969_));
  OAI210     m0920(.A0(mai_mai_n969_), .A1(mai_mai_n967_), .B0(mai_mai_n256_), .Y(mai_mai_n970_));
  NO2        m0921(.A(mai_mai_n828_), .B(mai_mai_n434_), .Y(mai_mai_n971_));
  NA3        m0922(.A(x4), .B(x3), .C(mai_mai_n98_), .Y(mai_mai_n972_));
  NO3        m0923(.A(mai_mai_n972_), .B(mai_mai_n680_), .C(mai_mai_n452_), .Y(mai_mai_n973_));
  AOI210     m0924(.A0(mai_mai_n971_), .A1(mai_mai_n459_), .B0(mai_mai_n973_), .Y(mai_mai_n974_));
  AOI210     m0925(.A0(mai_mai_n974_), .A1(mai_mai_n970_), .B0(mai_mai_n445_), .Y(mai_mai_n975_));
  NO2        m0926(.A(mai_mai_n55_), .B(mai_mai_n56_), .Y(mai_mai_n976_));
  OAI220     m0927(.A0(mai_mai_n784_), .A1(mai_mai_n447_), .B0(mai_mai_n722_), .B1(mai_mai_n117_), .Y(mai_mai_n977_));
  NOi21      m0928(.An(mai_mai_n112_), .B(mai_mai_n111_), .Y(mai_mai_n978_));
  NO3        m0929(.A(mai_mai_n332_), .B(mai_mai_n311_), .C(mai_mai_n978_), .Y(mai_mai_n979_));
  AOI220     m0930(.A0(mai_mai_n979_), .A1(mai_mai_n241_), .B0(mai_mai_n977_), .B1(mai_mai_n104_), .Y(mai_mai_n980_));
  NO2        m0931(.A(mai_mai_n980_), .B(mai_mai_n976_), .Y(mai_mai_n981_));
  NA2        m0932(.A(mai_mai_n506_), .B(mai_mai_n246_), .Y(mai_mai_n982_));
  NO2        m0933(.A(mai_mai_n474_), .B(mai_mai_n572_), .Y(mai_mai_n983_));
  NA3        m0934(.A(mai_mai_n983_), .B(mai_mai_n982_), .C(mai_mai_n55_), .Y(mai_mai_n984_));
  NO2        m0935(.A(mai_mai_n172_), .B(mai_mai_n98_), .Y(mai_mai_n985_));
  NA3        m0936(.A(mai_mai_n985_), .B(mai_mai_n171_), .C(mai_mai_n111_), .Y(mai_mai_n986_));
  NA2        m0937(.A(mai_mai_n986_), .B(mai_mai_n984_), .Y(mai_mai_n987_));
  NO4        m0938(.A(mai_mai_n987_), .B(mai_mai_n981_), .C(mai_mai_n975_), .D(mai_mai_n966_), .Y(mai_mai_n988_));
  NA3        m0939(.A(mai_mai_n988_), .B(mai_mai_n952_), .C(mai_mai_n939_), .Y(mai11));
  INV        m0940(.A(mai_mai_n848_), .Y(mai_mai_n990_));
  NO2        m0941(.A(mai_mai_n739_), .B(x5), .Y(mai_mai_n991_));
  NO2        m0942(.A(mai_mai_n157_), .B(mai_mai_n519_), .Y(mai_mai_n992_));
  AOI220     m0943(.A0(mai_mai_n992_), .A1(mai_mai_n991_), .B0(mai_mai_n848_), .B1(x5), .Y(mai_mai_n993_));
  OAI220     m0944(.A0(mai_mai_n926_), .A1(mai_mai_n206_), .B0(mai_mai_n204_), .B1(mai_mai_n172_), .Y(mai_mai_n994_));
  NO2        m0945(.A(mai_mai_n328_), .B(mai_mai_n415_), .Y(mai_mai_n995_));
  AOI220     m0946(.A0(mai_mai_n995_), .A1(mai_mai_n170_), .B0(mai_mai_n994_), .B1(mai_mai_n153_), .Y(mai_mai_n996_));
  NO2        m0947(.A(mai_mai_n996_), .B(mai_mai_n436_), .Y(mai_mai_n997_));
  NO2        m0948(.A(mai_mai_n237_), .B(x2), .Y(mai_mai_n998_));
  OAI210     m0949(.A0(mai_mai_n872_), .A1(mai_mai_n998_), .B0(mai_mai_n404_), .Y(mai_mai_n999_));
  NO2        m0950(.A(mai_mai_n55_), .B(mai_mai_n96_), .Y(mai_mai_n1000_));
  NA2        m0951(.A(mai_mai_n265_), .B(mai_mai_n1000_), .Y(mai_mai_n1001_));
  NO2        m0952(.A(mai_mai_n67_), .B(x1), .Y(mai_mai_n1002_));
  NA2        m0953(.A(mai_mai_n1002_), .B(mai_mai_n72_), .Y(mai_mai_n1003_));
  OA220      m0954(.A0(mai_mai_n1003_), .A1(mai_mai_n594_), .B0(mai_mai_n1001_), .B1(mai_mai_n519_), .Y(mai_mai_n1004_));
  AOI210     m0955(.A0(mai_mai_n1004_), .A1(mai_mai_n999_), .B0(mai_mai_n687_), .Y(mai_mai_n1005_));
  NO2        m0956(.A(mai_mai_n291_), .B(mai_mai_n53_), .Y(mai_mai_n1006_));
  NO2        m0957(.A(mai_mai_n425_), .B(x3), .Y(mai_mai_n1007_));
  NA3        m0958(.A(mai_mai_n1007_), .B(mai_mai_n1006_), .C(mai_mai_n847_), .Y(mai_mai_n1008_));
  AOI210     m0959(.A0(mai_mai_n1008_), .A1(mai_mai_n898_), .B0(mai_mai_n385_), .Y(mai_mai_n1009_));
  NA2        m0960(.A(mai_mai_n98_), .B(x1), .Y(mai_mai_n1010_));
  NO2        m0961(.A(mai_mai_n600_), .B(mai_mai_n209_), .Y(mai_mai_n1011_));
  NA4        m0962(.A(mai_mai_n1011_), .B(mai_mai_n840_), .C(mai_mai_n456_), .D(mai_mai_n1010_), .Y(mai_mai_n1012_));
  INV        m0963(.A(mai_mai_n1012_), .Y(mai_mai_n1013_));
  NO4        m0964(.A(mai_mai_n1013_), .B(mai_mai_n1009_), .C(mai_mai_n1005_), .D(mai_mai_n997_), .Y(mai_mai_n1014_));
  OAI210     m0965(.A0(mai_mai_n993_), .A1(mai_mai_n132_), .B0(mai_mai_n1014_), .Y(mai_mai_n1015_));
  NA2        m0966(.A(mai_mai_n822_), .B(mai_mai_n79_), .Y(mai_mai_n1016_));
  NO3        m0967(.A(mai_mai_n453_), .B(mai_mai_n745_), .C(mai_mai_n112_), .Y(mai_mai_n1017_));
  AOI210     m0968(.A0(mai_mai_n1016_), .A1(mai_mai_n92_), .B0(mai_mai_n1017_), .Y(mai_mai_n1018_));
  NO2        m0969(.A(x8), .B(x1), .Y(mai_mai_n1019_));
  NO3        m0970(.A(mai_mai_n1019_), .B(mai_mai_n666_), .C(mai_mai_n437_), .Y(mai_mai_n1020_));
  OAI210     m0971(.A0(mai_mai_n71_), .A1(mai_mai_n53_), .B0(mai_mai_n1020_), .Y(mai_mai_n1021_));
  OAI210     m0972(.A0(mai_mai_n1018_), .A1(x3), .B0(mai_mai_n1021_), .Y(mai_mai_n1022_));
  NO2        m0973(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n1023_));
  OAI210     m0974(.A0(mai_mai_n1023_), .A1(x2), .B0(mai_mai_n219_), .Y(mai_mai_n1024_));
  NO2        m0975(.A(mai_mai_n589_), .B(mai_mai_n217_), .Y(mai_mai_n1025_));
  NA2        m0976(.A(mai_mai_n1025_), .B(mai_mai_n1024_), .Y(mai_mai_n1026_));
  NO3        m0977(.A(mai_mai_n55_), .B(x6), .C(x1), .Y(mai_mai_n1027_));
  INV        m0978(.A(mai_mai_n1026_), .Y(mai_mai_n1028_));
  AOI210     m0979(.A0(mai_mai_n1022_), .A1(x2), .B0(mai_mai_n1028_), .Y(mai_mai_n1029_));
  NO2        m0980(.A(mai_mai_n217_), .B(x2), .Y(mai_mai_n1030_));
  NA2        m0981(.A(mai_mai_n1030_), .B(mai_mai_n953_), .Y(mai_mai_n1031_));
  NOi21      m0982(.An(mai_mai_n376_), .B(mai_mai_n554_), .Y(mai_mai_n1032_));
  NO3        m0983(.A(mai_mai_n1032_), .B(mai_mai_n588_), .C(mai_mai_n311_), .Y(mai_mai_n1033_));
  NA2        m0984(.A(x8), .B(mai_mai_n98_), .Y(mai_mai_n1034_));
  OAI220     m0985(.A0(mai_mai_n687_), .A1(mai_mai_n1034_), .B0(mai_mai_n311_), .B1(mai_mai_n371_), .Y(mai_mai_n1035_));
  OAI210     m0986(.A0(mai_mai_n1035_), .A1(mai_mai_n1033_), .B0(mai_mai_n67_), .Y(mai_mai_n1036_));
  NO2        m0987(.A(mai_mai_n96_), .B(x1), .Y(mai_mai_n1037_));
  NA2        m0988(.A(mai_mai_n1037_), .B(x7), .Y(mai_mai_n1038_));
  AOI210     m0989(.A0(mai_mai_n1036_), .A1(mai_mai_n1031_), .B0(mai_mai_n1038_), .Y(mai_mai_n1039_));
  NA2        m0990(.A(mai_mai_n76_), .B(mai_mai_n67_), .Y(mai_mai_n1040_));
  INV        m0991(.A(mai_mai_n234_), .Y(mai_mai_n1041_));
  NA2        m0992(.A(mai_mai_n1041_), .B(mai_mai_n139_), .Y(mai_mai_n1042_));
  OAI220     m0993(.A0(mai_mai_n1042_), .A1(mai_mai_n353_), .B0(mai_mai_n1040_), .B1(mai_mai_n311_), .Y(mai_mai_n1043_));
  NO2        m0994(.A(mai_mai_n148_), .B(mai_mai_n55_), .Y(mai_mai_n1044_));
  AOI210     m0995(.A0(mai_mai_n1044_), .A1(mai_mai_n1043_), .B0(mai_mai_n1039_), .Y(mai_mai_n1045_));
  OAI210     m0996(.A0(mai_mai_n1029_), .A1(mai_mai_n809_), .B0(mai_mai_n1045_), .Y(mai_mai_n1046_));
  AO210      m0997(.A0(mai_mai_n1015_), .A1(mai_mai_n57_), .B0(mai_mai_n1046_), .Y(mai12));
  NA2        m0998(.A(mai_mai_n839_), .B(mai_mai_n233_), .Y(mai_mai_n1048_));
  NO2        m0999(.A(mai_mai_n604_), .B(x7), .Y(mai_mai_n1049_));
  NA2        m1000(.A(mai_mai_n1049_), .B(mai_mai_n264_), .Y(mai_mai_n1050_));
  AOI210     m1001(.A0(mai_mai_n1050_), .A1(mai_mai_n1048_), .B0(mai_mai_n56_), .Y(mai_mai_n1051_));
  NOi21      m1002(.An(mai_mai_n392_), .B(mai_mai_n541_), .Y(mai_mai_n1052_));
  NO2        m1003(.A(x7), .B(mai_mai_n50_), .Y(mai_mai_n1053_));
  NO2        m1004(.A(mai_mai_n589_), .B(mai_mai_n1053_), .Y(mai_mai_n1054_));
  NO3        m1005(.A(mai_mai_n824_), .B(mai_mai_n100_), .C(mai_mai_n90_), .Y(mai_mai_n1055_));
  AOI210     m1006(.A0(mai_mai_n1054_), .A1(mai_mai_n961_), .B0(mai_mai_n1055_), .Y(mai_mai_n1056_));
  NA2        m1007(.A(mai_mai_n1000_), .B(mai_mai_n56_), .Y(mai_mai_n1057_));
  OAI220     m1008(.A0(mai_mai_n1057_), .A1(mai_mai_n565_), .B0(mai_mai_n1056_), .B1(mai_mai_n1052_), .Y(mai_mai_n1058_));
  OAI210     m1009(.A0(mai_mai_n1058_), .A1(mai_mai_n1051_), .B0(mai_mai_n568_), .Y(mai_mai_n1059_));
  NA2        m1010(.A(mai_mai_n79_), .B(x5), .Y(mai_mai_n1060_));
  NO2        m1011(.A(mai_mai_n1060_), .B(mai_mai_n311_), .Y(mai_mai_n1061_));
  AOI210     m1012(.A0(mai_mai_n786_), .A1(mai_mai_n106_), .B0(mai_mai_n1061_), .Y(mai_mai_n1062_));
  NA2        m1013(.A(mai_mai_n274_), .B(mai_mai_n50_), .Y(mai_mai_n1063_));
  NO2        m1014(.A(mai_mai_n1063_), .B(mai_mai_n297_), .Y(mai_mai_n1064_));
  NA2        m1015(.A(mai_mai_n1064_), .B(mai_mai_n56_), .Y(mai_mai_n1065_));
  OAI210     m1016(.A0(mai_mai_n1062_), .A1(mai_mai_n63_), .B0(mai_mai_n1065_), .Y(mai_mai_n1066_));
  NO2        m1017(.A(mai_mai_n57_), .B(x0), .Y(mai_mai_n1067_));
  NO2        m1018(.A(mai_mai_n647_), .B(mai_mai_n308_), .Y(mai_mai_n1068_));
  NO2        m1019(.A(mai_mai_n722_), .B(x3), .Y(mai_mai_n1069_));
  NO2        m1020(.A(mai_mai_n645_), .B(x8), .Y(mai_mai_n1070_));
  AOI220     m1021(.A0(mai_mai_n1070_), .A1(mai_mai_n1069_), .B0(mai_mai_n1068_), .B1(mai_mai_n1067_), .Y(mai_mai_n1071_));
  AOI210     m1022(.A0(mai_mai_n666_), .A1(mai_mai_n233_), .B0(x7), .Y(mai_mai_n1072_));
  NO3        m1023(.A(mai_mai_n1072_), .B(mai_mai_n590_), .C(x8), .Y(mai_mai_n1073_));
  NA4        m1024(.A(mai_mai_n648_), .B(mai_mai_n641_), .C(mai_mai_n194_), .D(x0), .Y(mai_mai_n1074_));
  OAI220     m1025(.A0(mai_mai_n1074_), .A1(mai_mai_n1073_), .B0(mai_mai_n1071_), .B1(mai_mai_n564_), .Y(mai_mai_n1075_));
  AOI210     m1026(.A0(mai_mai_n1066_), .A1(mai_mai_n968_), .B0(mai_mai_n1075_), .Y(mai_mai_n1076_));
  NO2        m1027(.A(mai_mai_n233_), .B(mai_mai_n55_), .Y(mai_mai_n1077_));
  NO2        m1028(.A(mai_mai_n241_), .B(x8), .Y(mai_mai_n1078_));
  NOi32      m1029(.An(mai_mai_n1078_), .Bn(mai_mai_n193_), .C(mai_mai_n555_), .Y(mai_mai_n1079_));
  NO2        m1030(.A(mai_mai_n80_), .B(mai_mai_n60_), .Y(mai_mai_n1080_));
  OAI210     m1031(.A0(mai_mai_n1079_), .A1(mai_mai_n1077_), .B0(mai_mai_n1080_), .Y(mai_mai_n1081_));
  NO2        m1032(.A(mai_mai_n901_), .B(mai_mai_n91_), .Y(mai_mai_n1082_));
  NO2        m1033(.A(mai_mai_n156_), .B(mai_mai_n53_), .Y(mai_mai_n1083_));
  AOI210     m1034(.A0(mai_mai_n328_), .A1(x8), .B0(mai_mai_n1083_), .Y(mai_mai_n1084_));
  AOI210     m1035(.A0(mai_mai_n206_), .A1(mai_mai_n88_), .B0(mai_mai_n1084_), .Y(mai_mai_n1085_));
  OAI210     m1036(.A0(mai_mai_n1085_), .A1(mai_mai_n1082_), .B0(mai_mai_n655_), .Y(mai_mai_n1086_));
  NO2        m1037(.A(x7), .B(x0), .Y(mai_mai_n1087_));
  NO2        m1038(.A(mai_mai_n148_), .B(mai_mai_n136_), .Y(mai_mai_n1088_));
  XN2        m1039(.A(x8), .B(x7), .Y(mai_mai_n1089_));
  NO3        m1040(.A(mai_mai_n1019_), .B(mai_mai_n244_), .C(mai_mai_n1089_), .Y(mai_mai_n1090_));
  OAI210     m1041(.A0(mai_mai_n1090_), .A1(mai_mai_n1088_), .B0(mai_mai_n703_), .Y(mai_mai_n1091_));
  NO2        m1042(.A(mai_mai_n253_), .B(mai_mai_n249_), .Y(mai_mai_n1092_));
  NO2        m1043(.A(mai_mai_n96_), .B(x4), .Y(mai_mai_n1093_));
  NA2        m1044(.A(mai_mai_n264_), .B(mai_mai_n1093_), .Y(mai_mai_n1094_));
  NA4        m1045(.A(mai_mai_n1094_), .B(mai_mai_n1091_), .C(mai_mai_n1086_), .D(mai_mai_n1081_), .Y(mai_mai_n1095_));
  NA2        m1046(.A(mai_mai_n1095_), .B(mai_mai_n545_), .Y(mai_mai_n1096_));
  NO2        m1047(.A(mai_mai_n55_), .B(x4), .Y(mai_mai_n1097_));
  NA2        m1048(.A(mai_mai_n1097_), .B(mai_mai_n152_), .Y(mai_mai_n1098_));
  NO2        m1049(.A(mai_mai_n650_), .B(mai_mai_n244_), .Y(mai_mai_n1099_));
  OAI210     m1050(.A0(mai_mai_n1099_), .A1(mai_mai_n971_), .B0(mai_mai_n50_), .Y(mai_mai_n1100_));
  AOI210     m1051(.A0(mai_mai_n1100_), .A1(mai_mai_n1098_), .B0(mai_mai_n420_), .Y(mai_mai_n1101_));
  OAI220     m1052(.A0(mai_mai_n276_), .A1(mai_mai_n262_), .B0(mai_mai_n249_), .B1(mai_mai_n228_), .Y(mai_mai_n1102_));
  NA3        m1053(.A(mai_mai_n1102_), .B(mai_mai_n655_), .C(x1), .Y(mai_mai_n1103_));
  OAI210     m1054(.A0(x8), .A1(x0), .B0(x4), .Y(mai_mai_n1104_));
  NO2        m1055(.A(x7), .B(mai_mai_n56_), .Y(mai_mai_n1105_));
  NO2        m1056(.A(mai_mai_n65_), .B(mai_mai_n1105_), .Y(mai_mai_n1106_));
  NOi21      m1057(.An(mai_mai_n1104_), .B(mai_mai_n1106_), .Y(mai_mai_n1107_));
  NO2        m1058(.A(mai_mai_n648_), .B(mai_mai_n311_), .Y(mai_mai_n1108_));
  NO2        m1059(.A(mai_mai_n748_), .B(mai_mai_n210_), .Y(mai_mai_n1109_));
  NA2        m1060(.A(mai_mai_n1107_), .B(mai_mai_n1109_), .Y(mai_mai_n1110_));
  NO2        m1061(.A(mai_mai_n132_), .B(mai_mai_n131_), .Y(mai_mai_n1111_));
  NO2        m1062(.A(mai_mai_n589_), .B(mai_mai_n434_), .Y(mai_mai_n1112_));
  OAI210     m1063(.A0(mai_mai_n1112_), .A1(mai_mai_n1111_), .B0(mai_mai_n241_), .Y(mai_mai_n1113_));
  NO2        m1064(.A(mai_mai_n782_), .B(mai_mai_n411_), .Y(mai_mai_n1114_));
  NA2        m1065(.A(mai_mai_n316_), .B(mai_mai_n59_), .Y(mai_mai_n1115_));
  NO2        m1066(.A(mai_mai_n1057_), .B(mai_mai_n1115_), .Y(mai_mai_n1116_));
  AOI210     m1067(.A0(mai_mai_n1114_), .A1(mai_mai_n168_), .B0(mai_mai_n1116_), .Y(mai_mai_n1117_));
  NA4        m1068(.A(mai_mai_n1117_), .B(mai_mai_n1113_), .C(mai_mai_n1110_), .D(mai_mai_n1103_), .Y(mai_mai_n1118_));
  OAI210     m1069(.A0(mai_mai_n1118_), .A1(mai_mai_n1101_), .B0(mai_mai_n657_), .Y(mai_mai_n1119_));
  NA4        m1070(.A(mai_mai_n1119_), .B(mai_mai_n1096_), .C(mai_mai_n1076_), .D(mai_mai_n1059_), .Y(mai13));
  NO2        m1071(.A(mai_mai_n824_), .B(mai_mai_n172_), .Y(mai_mai_n1121_));
  NO2        m1072(.A(mai_mai_n147_), .B(mai_mai_n67_), .Y(mai_mai_n1122_));
  XN2        m1073(.A(x4), .B(x0), .Y(mai_mai_n1123_));
  NO3        m1074(.A(mai_mai_n1123_), .B(mai_mai_n99_), .C(mai_mai_n411_), .Y(mai_mai_n1124_));
  AO220      m1075(.A0(mai_mai_n1124_), .A1(mai_mai_n1122_), .B0(mai_mai_n1121_), .B1(mai_mai_n317_), .Y(mai_mai_n1125_));
  NA2        m1076(.A(mai_mai_n1125_), .B(x3), .Y(mai_mai_n1126_));
  NO2        m1077(.A(mai_mai_n824_), .B(x6), .Y(mai_mai_n1127_));
  NO2        m1078(.A(mai_mai_n1063_), .B(mai_mai_n383_), .Y(mai_mai_n1128_));
  NO3        m1079(.A(x8), .B(x5), .C(mai_mai_n98_), .Y(mai_mai_n1129_));
  NA2        m1080(.A(mai_mai_n1129_), .B(mai_mai_n624_), .Y(mai_mai_n1130_));
  NO2        m1081(.A(mai_mai_n589_), .B(mai_mai_n188_), .Y(mai_mai_n1131_));
  NA2        m1082(.A(mai_mai_n437_), .B(mai_mai_n53_), .Y(mai_mai_n1132_));
  NO2        m1083(.A(mai_mai_n1132_), .B(mai_mai_n894_), .Y(mai_mai_n1133_));
  NA2        m1084(.A(mai_mai_n1057_), .B(mai_mai_n457_), .Y(mai_mai_n1134_));
  NA2        m1085(.A(mai_mai_n56_), .B(mai_mai_n98_), .Y(mai_mai_n1135_));
  NA2        m1086(.A(mai_mai_n1135_), .B(x1), .Y(mai_mai_n1136_));
  NO2        m1087(.A(mai_mai_n1136_), .B(mai_mai_n246_), .Y(mai_mai_n1137_));
  NO2        m1088(.A(mai_mai_n308_), .B(x6), .Y(mai_mai_n1138_));
  OAI210     m1089(.A0(mai_mai_n237_), .A1(mai_mai_n930_), .B0(mai_mai_n910_), .Y(mai_mai_n1139_));
  AOI220     m1090(.A0(mai_mai_n1139_), .A1(mai_mai_n1138_), .B0(mai_mai_n1137_), .B1(mai_mai_n1134_), .Y(mai_mai_n1140_));
  NAi31      m1091(.An(mai_mai_n1133_), .B(mai_mai_n1140_), .C(mai_mai_n1130_), .Y(mai_mai_n1141_));
  AOI220     m1092(.A0(mai_mai_n1141_), .A1(mai_mai_n65_), .B0(mai_mai_n1128_), .B1(mai_mai_n1127_), .Y(mai_mai_n1142_));
  NA2        m1093(.A(mai_mai_n67_), .B(x3), .Y(mai_mai_n1143_));
  NA2        m1094(.A(mai_mai_n1143_), .B(mai_mai_n856_), .Y(mai_mai_n1144_));
  OAI220     m1095(.A0(mai_mai_n290_), .A1(mai_mai_n782_), .B0(mai_mai_n79_), .B1(mai_mai_n71_), .Y(mai_mai_n1145_));
  AOI210     m1096(.A0(mai_mai_n1060_), .A1(mai_mai_n598_), .B0(mai_mai_n930_), .Y(mai_mai_n1146_));
  OA210      m1097(.A0(mai_mai_n1145_), .A1(mai_mai_n1144_), .B0(mai_mai_n1146_), .Y(mai_mai_n1147_));
  NA2        m1098(.A(mai_mai_n600_), .B(mai_mai_n55_), .Y(mai_mai_n1148_));
  NA2        m1099(.A(x6), .B(mai_mai_n50_), .Y(mai_mai_n1149_));
  NA2        m1100(.A(mai_mai_n1149_), .B(mai_mai_n528_), .Y(mai_mai_n1150_));
  NO2        m1101(.A(mai_mai_n149_), .B(mai_mai_n120_), .Y(mai_mai_n1151_));
  AOI210     m1102(.A0(mai_mai_n1150_), .A1(mai_mai_n421_), .B0(mai_mai_n1151_), .Y(mai_mai_n1152_));
  NO2        m1103(.A(mai_mai_n1152_), .B(mai_mai_n828_), .Y(mai_mai_n1153_));
  OAI210     m1104(.A0(mai_mai_n1153_), .A1(mai_mai_n1147_), .B0(mai_mai_n1087_), .Y(mai_mai_n1154_));
  NAi21      m1105(.An(mai_mai_n76_), .B(mai_mai_n371_), .Y(mai_mai_n1155_));
  NO2        m1106(.A(mai_mai_n1155_), .B(mai_mai_n67_), .Y(mai_mai_n1156_));
  NO2        m1107(.A(mai_mai_n160_), .B(mai_mai_n281_), .Y(mai_mai_n1157_));
  NA2        m1108(.A(mai_mai_n1157_), .B(mai_mai_n1156_), .Y(mai_mai_n1158_));
  NA3        m1109(.A(mai_mai_n1093_), .B(mai_mai_n179_), .C(mai_mai_n67_), .Y(mai_mai_n1159_));
  NO2        m1110(.A(x4), .B(x0), .Y(mai_mai_n1160_));
  NO3        m1111(.A(mai_mai_n947_), .B(mai_mai_n234_), .C(mai_mai_n528_), .Y(mai_mai_n1161_));
  OAI210     m1112(.A0(mai_mai_n1161_), .A1(mai_mai_n189_), .B0(mai_mai_n1160_), .Y(mai_mai_n1162_));
  NA3        m1113(.A(mai_mai_n1162_), .B(mai_mai_n1159_), .C(mai_mai_n1158_), .Y(mai_mai_n1163_));
  NA2        m1114(.A(mai_mai_n236_), .B(mai_mai_n703_), .Y(mai_mai_n1164_));
  NO2        m1115(.A(mai_mai_n1164_), .B(mai_mai_n508_), .Y(mai_mai_n1165_));
  NA2        m1116(.A(mai_mai_n56_), .B(x0), .Y(mai_mai_n1166_));
  NO3        m1117(.A(mai_mai_n1166_), .B(mai_mai_n483_), .C(mai_mai_n73_), .Y(mai_mai_n1167_));
  OAI210     m1118(.A0(mai_mai_n1167_), .A1(mai_mai_n1165_), .B0(x2), .Y(mai_mai_n1168_));
  NO2        m1119(.A(mai_mai_n311_), .B(mai_mai_n371_), .Y(mai_mai_n1169_));
  NO2        m1120(.A(mai_mai_n666_), .B(x0), .Y(mai_mai_n1170_));
  OAI210     m1121(.A0(mai_mai_n1170_), .A1(mai_mai_n1169_), .B0(mai_mai_n320_), .Y(mai_mai_n1171_));
  NO2        m1122(.A(mai_mai_n758_), .B(x1), .Y(mai_mai_n1172_));
  AOI220     m1123(.A0(mai_mai_n1172_), .A1(mai_mai_n593_), .B0(mai_mai_n467_), .B1(mai_mai_n282_), .Y(mai_mai_n1173_));
  NA2        m1124(.A(mai_mai_n488_), .B(mai_mai_n50_), .Y(mai_mai_n1174_));
  AOI220     m1125(.A0(mai_mai_n1174_), .A1(mai_mai_n1121_), .B0(mai_mai_n931_), .B1(mai_mai_n92_), .Y(mai_mai_n1175_));
  NA4        m1126(.A(mai_mai_n1175_), .B(mai_mai_n1173_), .C(mai_mai_n1171_), .D(mai_mai_n1168_), .Y(mai_mai_n1176_));
  AOI220     m1127(.A0(mai_mai_n1176_), .A1(mai_mai_n121_), .B0(mai_mai_n1163_), .B1(mai_mai_n64_), .Y(mai_mai_n1177_));
  NA4        m1128(.A(mai_mai_n1177_), .B(mai_mai_n1154_), .C(mai_mai_n1142_), .D(mai_mai_n1126_), .Y(mai14));
  NO2        m1129(.A(mai_mai_n359_), .B(mai_mai_n67_), .Y(mai_mai_n1179_));
  NO3        m1130(.A(x7), .B(x6), .C(x0), .Y(mai_mai_n1180_));
  OAI210     m1131(.A0(mai_mai_n1180_), .A1(mai_mai_n1179_), .B0(x8), .Y(mai_mai_n1181_));
  NO2        m1132(.A(mai_mai_n1181_), .B(mai_mai_n146_), .Y(mai_mai_n1182_));
  AOI220     m1133(.A0(mai_mai_n363_), .A1(mai_mai_n809_), .B0(mai_mai_n437_), .B1(mai_mai_n411_), .Y(mai_mai_n1183_));
  NA2        m1134(.A(mai_mai_n265_), .B(mai_mai_n926_), .Y(mai_mai_n1184_));
  OAI220     m1135(.A0(mai_mai_n1184_), .A1(mai_mai_n1183_), .B0(mai_mai_n455_), .B1(mai_mai_n768_), .Y(mai_mai_n1185_));
  OA210      m1136(.A0(mai_mai_n1185_), .A1(mai_mai_n1182_), .B0(x4), .Y(mai_mai_n1186_));
  NO2        m1137(.A(mai_mai_n131_), .B(mai_mai_n591_), .Y(mai_mai_n1187_));
  NA2        m1138(.A(x6), .B(x2), .Y(mai_mai_n1188_));
  NO2        m1139(.A(mai_mai_n609_), .B(mai_mai_n1188_), .Y(mai_mai_n1189_));
  OA210      m1140(.A0(mai_mai_n1187_), .A1(mai_mai_n202_), .B0(mai_mai_n1189_), .Y(mai_mai_n1190_));
  NO4        m1141(.A(mai_mai_n589_), .B(mai_mai_n364_), .C(mai_mai_n286_), .D(mai_mai_n104_), .Y(mai_mai_n1191_));
  OAI210     m1142(.A0(mai_mai_n1191_), .A1(mai_mai_n1190_), .B0(mai_mai_n59_), .Y(mai_mai_n1192_));
  NA2        m1143(.A(x6), .B(mai_mai_n96_), .Y(mai_mai_n1193_));
  NO2        m1144(.A(mai_mai_n647_), .B(mai_mai_n1193_), .Y(mai_mai_n1194_));
  NA2        m1145(.A(mai_mai_n1194_), .B(mai_mai_n881_), .Y(mai_mai_n1195_));
  AOI210     m1146(.A0(mai_mai_n1070_), .A1(mai_mai_n960_), .B0(x1), .Y(mai_mai_n1196_));
  NO2        m1147(.A(mai_mai_n523_), .B(x5), .Y(mai_mai_n1197_));
  NA3        m1148(.A(mai_mai_n1197_), .B(mai_mai_n111_), .C(x0), .Y(mai_mai_n1198_));
  NA4        m1149(.A(mai_mai_n673_), .B(mai_mai_n882_), .C(mai_mai_n290_), .D(mai_mai_n65_), .Y(mai_mai_n1199_));
  AN4        m1150(.A(mai_mai_n1199_), .B(mai_mai_n1198_), .C(mai_mai_n1196_), .D(mai_mai_n1195_), .Y(mai_mai_n1200_));
  NO2        m1151(.A(mai_mai_n680_), .B(mai_mai_n1034_), .Y(mai_mai_n1201_));
  NO2        m1152(.A(mai_mai_n71_), .B(mai_mai_n58_), .Y(mai_mai_n1202_));
  OAI210     m1153(.A0(mai_mai_n1201_), .A1(mai_mai_n435_), .B0(mai_mai_n1202_), .Y(mai_mai_n1203_));
  AOI220     m1154(.A0(x1), .A1(mai_mai_n1203_), .B0(mai_mai_n1200_), .B1(mai_mai_n1192_), .Y(mai_mai_n1204_));
  NO2        m1155(.A(mai_mai_n656_), .B(mai_mai_n156_), .Y(mai_mai_n1205_));
  NO3        m1156(.A(mai_mai_n1205_), .B(mai_mai_n1204_), .C(mai_mai_n1186_), .Y(mai_mai_n1206_));
  NO2        m1157(.A(mai_mai_n308_), .B(x2), .Y(mai_mai_n1207_));
  XN2        m1158(.A(x4), .B(x1), .Y(mai_mai_n1208_));
  NO2        m1159(.A(mai_mai_n1208_), .B(mai_mai_n290_), .Y(mai_mai_n1209_));
  NO2        m1160(.A(mai_mai_n327_), .B(mai_mai_n60_), .Y(mai_mai_n1210_));
  NA2        m1161(.A(mai_mai_n1210_), .B(mai_mai_n1207_), .Y(mai_mai_n1211_));
  NA2        m1162(.A(mai_mai_n667_), .B(mai_mai_n56_), .Y(mai_mai_n1212_));
  OAI220     m1163(.A0(mai_mai_n1212_), .A1(mai_mai_n147_), .B0(mai_mai_n180_), .B1(mai_mai_n67_), .Y(mai_mai_n1213_));
  NO2        m1164(.A(mai_mai_n206_), .B(mai_mai_n244_), .Y(mai_mai_n1214_));
  AOI220     m1165(.A0(mai_mai_n128_), .A1(mai_mai_n56_), .B0(mai_mai_n85_), .B1(x5), .Y(mai_mai_n1215_));
  NA2        m1166(.A(mai_mai_n1027_), .B(mai_mai_n295_), .Y(mai_mai_n1216_));
  NA2        m1167(.A(mai_mai_n236_), .B(mai_mai_n342_), .Y(mai_mai_n1217_));
  OAI220     m1168(.A0(mai_mai_n2513_), .A1(mai_mai_n1217_), .B0(mai_mai_n1216_), .B1(mai_mai_n1215_), .Y(mai_mai_n1218_));
  AOI210     m1169(.A0(mai_mai_n1214_), .A1(mai_mai_n1213_), .B0(mai_mai_n1218_), .Y(mai_mai_n1219_));
  AOI210     m1170(.A0(mai_mai_n1219_), .A1(mai_mai_n1211_), .B0(x7), .Y(mai_mai_n1220_));
  NO2        m1171(.A(mai_mai_n482_), .B(x6), .Y(mai_mai_n1221_));
  AOI210     m1172(.A0(mai_mai_n778_), .A1(mai_mai_n912_), .B0(mai_mai_n1221_), .Y(mai_mai_n1222_));
  OAI220     m1173(.A0(mai_mai_n1222_), .A1(mai_mai_n55_), .B0(mai_mai_n482_), .B1(mai_mai_n94_), .Y(mai_mai_n1223_));
  NA2        m1174(.A(mai_mai_n1223_), .B(mai_mai_n344_), .Y(mai_mai_n1224_));
  NA3        m1175(.A(mai_mai_n594_), .B(mai_mai_n1010_), .C(mai_mai_n66_), .Y(mai_mai_n1225_));
  NO4        m1176(.A(mai_mai_n1225_), .B(mai_mai_n1166_), .C(mai_mai_n109_), .D(mai_mai_n55_), .Y(mai_mai_n1226_));
  NO2        m1177(.A(mai_mai_n1003_), .B(mai_mai_n784_), .Y(mai_mai_n1227_));
  NO3        m1178(.A(mai_mai_n722_), .B(mai_mai_n488_), .C(mai_mai_n54_), .Y(mai_mai_n1228_));
  NO3        m1179(.A(mai_mai_n1228_), .B(mai_mai_n1227_), .C(mai_mai_n1226_), .Y(mai_mai_n1229_));
  AOI210     m1180(.A0(mai_mai_n1229_), .A1(mai_mai_n1224_), .B0(mai_mai_n292_), .Y(mai_mai_n1230_));
  NA2        m1181(.A(mai_mai_n854_), .B(mai_mai_n53_), .Y(mai_mai_n1231_));
  OAI210     m1182(.A0(mai_mai_n231_), .A1(mai_mai_n106_), .B0(x2), .Y(mai_mai_n1232_));
  NA2        m1183(.A(mai_mai_n355_), .B(mai_mai_n56_), .Y(mai_mai_n1233_));
  OA220      m1184(.A0(mai_mai_n1233_), .A1(mai_mai_n1232_), .B0(mai_mai_n1231_), .B1(mai_mai_n363_), .Y(mai_mai_n1234_));
  NA3        m1185(.A(mai_mai_n983_), .B(mai_mai_n707_), .C(mai_mai_n55_), .Y(mai_mai_n1235_));
  NA2        m1186(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n1236_));
  NO2        m1187(.A(mai_mai_n1236_), .B(mai_mai_n187_), .Y(mai_mai_n1237_));
  NA4        m1188(.A(mai_mai_n1237_), .B(mai_mai_n355_), .C(mai_mai_n244_), .D(mai_mai_n64_), .Y(mai_mai_n1238_));
  NA3        m1189(.A(mai_mai_n1172_), .B(mai_mai_n600_), .C(mai_mai_n614_), .Y(mai_mai_n1239_));
  AN3        m1190(.A(mai_mai_n1239_), .B(mai_mai_n1238_), .C(mai_mai_n1235_), .Y(mai_mai_n1240_));
  OAI210     m1191(.A0(mai_mai_n1234_), .A1(mai_mai_n303_), .B0(mai_mai_n1240_), .Y(mai_mai_n1241_));
  NO3        m1192(.A(mai_mai_n1241_), .B(mai_mai_n1230_), .C(mai_mai_n1220_), .Y(mai_mai_n1242_));
  OAI210     m1193(.A0(mai_mai_n1206_), .A1(x3), .B0(mai_mai_n1242_), .Y(mai15));
  NA2        m1194(.A(mai_mai_n573_), .B(mai_mai_n59_), .Y(mai_mai_n1244_));
  NAi41      m1195(.An(x2), .B(x7), .C(x6), .D(x0), .Y(mai_mai_n1245_));
  AOI210     m1196(.A0(mai_mai_n1245_), .A1(mai_mai_n1244_), .B0(mai_mai_n53_), .Y(mai_mai_n1246_));
  NA3        m1197(.A(mai_mai_n57_), .B(x6), .C(mai_mai_n98_), .Y(mai_mai_n1247_));
  NO2        m1198(.A(mai_mai_n1247_), .B(mai_mai_n281_), .Y(mai_mai_n1248_));
  OAI210     m1199(.A0(mai_mai_n1248_), .A1(mai_mai_n1246_), .B0(mai_mai_n1093_), .Y(mai_mai_n1249_));
  NA2        m1200(.A(mai_mai_n100_), .B(mai_mai_n98_), .Y(mai_mai_n1250_));
  NA4        m1201(.A(mai_mai_n1250_), .B(mai_mai_n621_), .C(mai_mai_n296_), .D(x6), .Y(mai_mai_n1251_));
  AOI210     m1202(.A0(mai_mai_n702_), .A1(mai_mai_n70_), .B0(x3), .Y(mai_mai_n1252_));
  NA3        m1203(.A(mai_mai_n1252_), .B(mai_mai_n1251_), .C(mai_mai_n1249_), .Y(mai_mai_n1253_));
  NO2        m1204(.A(mai_mai_n281_), .B(mai_mai_n98_), .Y(mai_mai_n1254_));
  NO2        m1205(.A(mai_mai_n223_), .B(x5), .Y(mai_mai_n1255_));
  NA2        m1206(.A(mai_mai_n1255_), .B(mai_mai_n1254_), .Y(mai_mai_n1256_));
  NA3        m1207(.A(mai_mai_n1172_), .B(mai_mai_n608_), .C(mai_mai_n1105_), .Y(mai_mai_n1257_));
  NA4        m1208(.A(mai_mai_n1257_), .B(mai_mai_n1256_), .C(x3), .D(mai_mai_n1198_), .Y(mai_mai_n1258_));
  NA2        m1209(.A(mai_mai_n577_), .B(mai_mai_n456_), .Y(mai_mai_n1259_));
  NO2        m1210(.A(mai_mai_n722_), .B(mai_mai_n53_), .Y(mai_mai_n1260_));
  NO2        m1211(.A(mai_mai_n748_), .B(mai_mai_n286_), .Y(mai_mai_n1261_));
  NA2        m1212(.A(mai_mai_n1261_), .B(mai_mai_n1260_), .Y(mai_mai_n1262_));
  NA2        m1213(.A(mai_mai_n1262_), .B(mai_mai_n1259_), .Y(mai_mai_n1263_));
  NA2        m1214(.A(mai_mai_n1263_), .B(mai_mai_n71_), .Y(mai_mai_n1264_));
  NA2        m1215(.A(mai_mai_n357_), .B(mai_mai_n682_), .Y(mai_mai_n1265_));
  NA3        m1216(.A(mai_mai_n53_), .B(mai_mai_n330_), .C(mai_mai_n100_), .Y(mai_mai_n1266_));
  AOI210     m1217(.A0(mai_mai_n1266_), .A1(mai_mai_n1265_), .B0(mai_mai_n488_), .Y(mai_mai_n1267_));
  NO3        m1218(.A(mai_mai_n767_), .B(mai_mai_n605_), .C(mai_mai_n188_), .Y(mai_mai_n1268_));
  OAI210     m1219(.A0(mai_mai_n1268_), .A1(mai_mai_n1267_), .B0(mai_mai_n482_), .Y(mai_mai_n1269_));
  NO2        m1220(.A(mai_mai_n233_), .B(mai_mai_n63_), .Y(mai_mai_n1270_));
  NA2        m1221(.A(mai_mai_n57_), .B(x3), .Y(mai_mai_n1271_));
  AOI210     m1222(.A0(mai_mai_n932_), .A1(mai_mai_n1271_), .B0(mai_mai_n661_), .Y(mai_mai_n1272_));
  NA2        m1223(.A(mai_mai_n1272_), .B(mai_mai_n968_), .Y(mai_mai_n1273_));
  NA2        m1224(.A(mai_mai_n1237_), .B(mai_mai_n65_), .Y(mai_mai_n1274_));
  NO2        m1225(.A(mai_mai_n420_), .B(mai_mai_n73_), .Y(mai_mai_n1275_));
  NO2        m1226(.A(mai_mai_n888_), .B(mai_mai_n67_), .Y(mai_mai_n1276_));
  NA2        m1227(.A(mai_mai_n1276_), .B(mai_mai_n1275_), .Y(mai_mai_n1277_));
  NO2        m1228(.A(mai_mai_n930_), .B(x6), .Y(mai_mai_n1278_));
  NA4        m1229(.A(mai_mai_n1278_), .B(mai_mai_n582_), .C(mai_mai_n148_), .D(mai_mai_n403_), .Y(mai_mai_n1279_));
  AN4        m1230(.A(mai_mai_n1279_), .B(mai_mai_n1277_), .C(mai_mai_n2512_), .D(mai_mai_n1274_), .Y(mai_mai_n1280_));
  NA4        m1231(.A(mai_mai_n1280_), .B(mai_mai_n1273_), .C(mai_mai_n1269_), .D(mai_mai_n1264_), .Y(mai_mai_n1281_));
  NA2        m1232(.A(mai_mai_n153_), .B(mai_mai_n707_), .Y(mai_mai_n1282_));
  NO2        m1233(.A(mai_mai_n633_), .B(x2), .Y(mai_mai_n1283_));
  OAI210     m1234(.A0(mai_mai_n65_), .A1(mai_mai_n53_), .B0(mai_mai_n134_), .Y(mai_mai_n1284_));
  OAI210     m1235(.A0(mai_mai_n1283_), .A1(mai_mai_n77_), .B0(mai_mai_n1284_), .Y(mai_mai_n1285_));
  AOI210     m1236(.A0(mai_mai_n1285_), .A1(mai_mai_n1282_), .B0(mai_mai_n308_), .Y(mai_mai_n1286_));
  NO3        m1237(.A(mai_mai_n1247_), .B(mai_mai_n252_), .C(mai_mai_n233_), .Y(mai_mai_n1287_));
  NA3        m1238(.A(mai_mai_n57_), .B(x1), .C(x0), .Y(mai_mai_n1288_));
  NA3        m1239(.A(mai_mai_n67_), .B(x5), .C(x2), .Y(mai_mai_n1289_));
  NA4        m1240(.A(x7), .B(x3), .C(mai_mai_n53_), .D(x0), .Y(mai_mai_n1290_));
  OAI220     m1241(.A0(mai_mai_n1290_), .A1(x6), .B0(mai_mai_n1289_), .B1(mai_mai_n1288_), .Y(mai_mai_n1291_));
  NO2        m1242(.A(mai_mai_n1291_), .B(mai_mai_n1287_), .Y(mai_mai_n1292_));
  NAi21      m1243(.An(mai_mai_n104_), .B(mai_mai_n717_), .Y(mai_mai_n1293_));
  NA4        m1244(.A(mai_mai_n1293_), .B(mai_mai_n306_), .C(mai_mai_n276_), .D(mai_mai_n608_), .Y(mai_mai_n1294_));
  NA2        m1245(.A(mai_mai_n74_), .B(mai_mai_n50_), .Y(mai_mai_n1295_));
  AO210      m1246(.A0(mai_mai_n1295_), .A1(mai_mai_n301_), .B0(mai_mai_n146_), .Y(mai_mai_n1296_));
  NA3        m1247(.A(mai_mai_n1296_), .B(mai_mai_n1294_), .C(mai_mai_n1292_), .Y(mai_mai_n1297_));
  OAI210     m1248(.A0(mai_mai_n1297_), .A1(mai_mai_n1286_), .B0(mai_mai_n56_), .Y(mai_mai_n1298_));
  AOI210     m1249(.A0(mai_mai_n669_), .A1(x4), .B0(mai_mai_n912_), .Y(mai_mai_n1299_));
  NO2        m1250(.A(mai_mai_n1299_), .B(mai_mai_n287_), .Y(mai_mai_n1300_));
  NA2        m1251(.A(mai_mai_n795_), .B(mai_mai_n396_), .Y(mai_mai_n1301_));
  OAI210     m1252(.A0(mai_mai_n1275_), .A1(mai_mai_n1270_), .B0(mai_mai_n277_), .Y(mai_mai_n1302_));
  OAI210     m1253(.A0(mai_mai_n1301_), .A1(mai_mai_n805_), .B0(mai_mai_n1302_), .Y(mai_mai_n1303_));
  OAI210     m1254(.A0(mai_mai_n1303_), .A1(mai_mai_n1300_), .B0(x6), .Y(mai_mai_n1304_));
  NO2        m1255(.A(mai_mai_n57_), .B(mai_mai_n59_), .Y(mai_mai_n1305_));
  NO2        m1256(.A(x7), .B(x5), .Y(mai_mai_n1306_));
  AOI220     m1257(.A0(mai_mai_n813_), .A1(mai_mai_n1305_), .B0(mai_mai_n527_), .B1(mai_mai_n1306_), .Y(mai_mai_n1307_));
  NA2        m1258(.A(mai_mai_n732_), .B(mai_mai_n277_), .Y(mai_mai_n1308_));
  INV        m1259(.A(mai_mai_n1307_), .Y(mai_mai_n1309_));
  NA2        m1260(.A(mai_mai_n1309_), .B(mai_mai_n414_), .Y(mai_mai_n1310_));
  AOI210     m1261(.A0(mai_mai_n367_), .A1(mai_mai_n328_), .B0(mai_mai_n55_), .Y(mai_mai_n1311_));
  NA4        m1262(.A(mai_mai_n1311_), .B(mai_mai_n1310_), .C(mai_mai_n1304_), .D(mai_mai_n1298_), .Y(mai_mai_n1312_));
  AO220      m1263(.A0(mai_mai_n1312_), .A1(mai_mai_n1281_), .B0(mai_mai_n1258_), .B1(mai_mai_n1253_), .Y(mai16));
  NO2        m1264(.A(x4), .B(mai_mai_n59_), .Y(mai_mai_n1314_));
  NA2        m1265(.A(mai_mai_n646_), .B(mai_mai_n524_), .Y(mai_mai_n1315_));
  NA3        m1266(.A(mai_mai_n217_), .B(mai_mai_n421_), .C(mai_mai_n912_), .Y(mai_mai_n1316_));
  NA2        m1267(.A(mai_mai_n123_), .B(mai_mai_n197_), .Y(mai_mai_n1317_));
  AOI210     m1268(.A0(mai_mai_n1316_), .A1(mai_mai_n1315_), .B0(mai_mai_n1317_), .Y(mai_mai_n1318_));
  NO3        m1269(.A(x8), .B(x6), .C(mai_mai_n50_), .Y(mai_mai_n1319_));
  NO2        m1270(.A(mai_mai_n706_), .B(mai_mai_n175_), .Y(mai_mai_n1320_));
  OAI210     m1271(.A0(mai_mai_n1319_), .A1(mai_mai_n225_), .B0(mai_mai_n1320_), .Y(mai_mai_n1321_));
  NO2        m1272(.A(mai_mai_n149_), .B(x5), .Y(mai_mai_n1322_));
  NA2        m1273(.A(mai_mai_n1322_), .B(mai_mai_n1283_), .Y(mai_mai_n1323_));
  NA3        m1274(.A(mai_mai_n568_), .B(mai_mai_n526_), .C(mai_mai_n466_), .Y(mai_mai_n1324_));
  NA3        m1275(.A(mai_mai_n1324_), .B(mai_mai_n1323_), .C(mai_mai_n1321_), .Y(mai_mai_n1325_));
  OAI210     m1276(.A0(mai_mai_n1325_), .A1(mai_mai_n1318_), .B0(mai_mai_n1314_), .Y(mai_mai_n1326_));
  OAI210     m1277(.A0(mai_mai_n1207_), .A1(mai_mai_n881_), .B0(mai_mai_n411_), .Y(mai_mai_n1327_));
  NO2        m1278(.A(mai_mai_n308_), .B(x7), .Y(mai_mai_n1328_));
  NA2        m1279(.A(mai_mai_n1328_), .B(x0), .Y(mai_mai_n1329_));
  AOI210     m1280(.A0(mai_mai_n1329_), .A1(mai_mai_n1327_), .B0(mai_mai_n622_), .Y(mai_mai_n1330_));
  NA2        m1281(.A(mai_mai_n1019_), .B(mai_mai_n188_), .Y(mai_mai_n1331_));
  NA2        m1282(.A(mai_mai_n55_), .B(mai_mai_n96_), .Y(mai_mai_n1332_));
  NA2        m1283(.A(mai_mai_n1332_), .B(mai_mai_n663_), .Y(mai_mai_n1333_));
  NA2        m1284(.A(mai_mai_n366_), .B(mai_mai_n1023_), .Y(mai_mai_n1334_));
  OA220      m1285(.A0(mai_mai_n1334_), .A1(mai_mai_n1333_), .B0(mai_mai_n1331_), .B1(mai_mai_n616_), .Y(mai_mai_n1335_));
  OAI210     m1286(.A0(mai_mai_n1335_), .A1(mai_mai_n637_), .B0(mai_mai_n486_), .Y(mai_mai_n1336_));
  INV        m1287(.A(mai_mai_n968_), .Y(mai_mai_n1337_));
  NO2        m1288(.A(mai_mai_n1337_), .B(mai_mai_n61_), .Y(mai_mai_n1338_));
  AOI220     m1289(.A0(mai_mai_n1338_), .A1(mai_mai_n256_), .B0(mai_mai_n1194_), .B1(mai_mai_n116_), .Y(mai_mai_n1339_));
  AOI220     m1290(.A0(mai_mai_n621_), .A1(mai_mai_n351_), .B0(mai_mai_n608_), .B1(mai_mai_n80_), .Y(mai_mai_n1340_));
  NA3        m1291(.A(mai_mai_n453_), .B(mai_mai_n574_), .C(mai_mai_n182_), .Y(mai_mai_n1341_));
  OAI220     m1292(.A0(mai_mai_n1341_), .A1(mai_mai_n1340_), .B0(mai_mai_n1339_), .B1(mai_mai_n297_), .Y(mai_mai_n1342_));
  NO3        m1293(.A(mai_mai_n1342_), .B(mai_mai_n1336_), .C(mai_mai_n1330_), .Y(mai_mai_n1343_));
  NO3        m1294(.A(x6), .B(x4), .C(x3), .Y(mai_mai_n1344_));
  NA2        m1295(.A(mai_mai_n1344_), .B(mai_mai_n523_), .Y(mai_mai_n1345_));
  NA4        m1296(.A(mai_mai_n687_), .B(mai_mai_n175_), .C(mai_mai_n58_), .D(x6), .Y(mai_mai_n1346_));
  AOI210     m1297(.A0(mai_mai_n1346_), .A1(mai_mai_n1345_), .B0(mai_mai_n54_), .Y(mai_mai_n1347_));
  NO2        m1298(.A(mai_mai_n694_), .B(x3), .Y(mai_mai_n1348_));
  AOI210     m1299(.A0(mai_mai_n645_), .A1(mai_mai_n138_), .B0(mai_mai_n1010_), .Y(mai_mai_n1349_));
  OA210      m1300(.A0(mai_mai_n1348_), .A1(mai_mai_n414_), .B0(mai_mai_n1349_), .Y(mai_mai_n1350_));
  NO3        m1301(.A(mai_mai_n488_), .B(mai_mai_n210_), .C(mai_mai_n69_), .Y(mai_mai_n1351_));
  NO2        m1302(.A(mai_mai_n732_), .B(mai_mai_n500_), .Y(mai_mai_n1352_));
  NO3        m1303(.A(mai_mai_n1352_), .B(mai_mai_n246_), .C(mai_mai_n145_), .Y(mai_mai_n1353_));
  NO4        m1304(.A(mai_mai_n1353_), .B(mai_mai_n1351_), .C(mai_mai_n1350_), .D(mai_mai_n1347_), .Y(mai_mai_n1354_));
  NA2        m1305(.A(mai_mai_n397_), .B(mai_mai_n912_), .Y(mai_mai_n1355_));
  NA4        m1306(.A(mai_mai_n472_), .B(mai_mai_n359_), .C(mai_mai_n212_), .D(x6), .Y(mai_mai_n1356_));
  OAI210     m1307(.A0(mai_mai_n694_), .A1(mai_mai_n1355_), .B0(mai_mai_n1356_), .Y(mai_mai_n1357_));
  NA2        m1308(.A(mai_mai_n863_), .B(mai_mai_n1236_), .Y(mai_mai_n1358_));
  NA2        m1309(.A(mai_mai_n703_), .B(x7), .Y(mai_mai_n1359_));
  OAI210     m1310(.A0(mai_mai_n1359_), .A1(mai_mai_n378_), .B0(mai_mai_n1358_), .Y(mai_mai_n1360_));
  NA2        m1311(.A(mai_mai_n263_), .B(x2), .Y(mai_mai_n1361_));
  OA210      m1312(.A0(mai_mai_n1193_), .A1(mai_mai_n58_), .B0(mai_mai_n749_), .Y(mai_mai_n1362_));
  NO2        m1313(.A(mai_mai_n1362_), .B(mai_mai_n180_), .Y(mai_mai_n1363_));
  NO3        m1314(.A(mai_mai_n1363_), .B(mai_mai_n1360_), .C(mai_mai_n1357_), .Y(mai_mai_n1364_));
  OA220      m1315(.A0(mai_mai_n1364_), .A1(mai_mai_n434_), .B0(mai_mai_n1354_), .B1(mai_mai_n195_), .Y(mai_mai_n1365_));
  NO2        m1316(.A(mai_mai_n877_), .B(mai_mai_n55_), .Y(mai_mai_n1366_));
  NA2        m1317(.A(mai_mai_n408_), .B(mai_mai_n768_), .Y(mai_mai_n1367_));
  NO2        m1318(.A(mai_mai_n1367_), .B(mai_mai_n1366_), .Y(mai_mai_n1368_));
  NO3        m1319(.A(mai_mai_n913_), .B(mai_mai_n321_), .C(x8), .Y(mai_mai_n1369_));
  OAI210     m1320(.A0(mai_mai_n1369_), .A1(mai_mai_n1368_), .B0(x6), .Y(mai_mai_n1370_));
  NO2        m1321(.A(mai_mai_n1032_), .B(mai_mai_n1002_), .Y(mai_mai_n1371_));
  NA2        m1322(.A(mai_mai_n180_), .B(x7), .Y(mai_mai_n1372_));
  OAI220     m1323(.A0(mai_mai_n1372_), .A1(mai_mai_n1371_), .B0(mai_mai_n734_), .B1(mai_mai_n79_), .Y(mai_mai_n1373_));
  NA2        m1324(.A(mai_mai_n1373_), .B(mai_mai_n882_), .Y(mai_mai_n1374_));
  NA2        m1325(.A(mai_mai_n830_), .B(mai_mai_n67_), .Y(mai_mai_n1375_));
  OAI210     m1326(.A0(mai_mai_n1375_), .A1(mai_mai_n148_), .B0(mai_mai_n957_), .Y(mai_mai_n1376_));
  AOI210     m1327(.A0(mai_mai_n488_), .A1(mai_mai_n57_), .B0(mai_mai_n616_), .Y(mai_mai_n1377_));
  NA3        m1328(.A(mai_mai_n214_), .B(mai_mai_n70_), .C(mai_mai_n67_), .Y(mai_mai_n1378_));
  OAI210     m1329(.A0(mai_mai_n873_), .A1(mai_mai_n217_), .B0(mai_mai_n1378_), .Y(mai_mai_n1379_));
  AOI210     m1330(.A0(mai_mai_n1377_), .A1(mai_mai_n1376_), .B0(mai_mai_n1379_), .Y(mai_mai_n1380_));
  NA3        m1331(.A(mai_mai_n1380_), .B(mai_mai_n1374_), .C(mai_mai_n1370_), .Y(mai_mai_n1381_));
  NO2        m1332(.A(mai_mai_n623_), .B(x6), .Y(mai_mai_n1382_));
  OAI210     m1333(.A0(mai_mai_n373_), .A1(mai_mai_n76_), .B0(mai_mai_n371_), .Y(mai_mai_n1383_));
  OA210      m1334(.A0(mai_mai_n1383_), .A1(mai_mai_n1382_), .B0(mai_mai_n121_), .Y(mai_mai_n1384_));
  NO3        m1335(.A(mai_mai_n436_), .B(mai_mai_n376_), .C(x7), .Y(mai_mai_n1385_));
  NO3        m1336(.A(mai_mai_n149_), .B(mai_mai_n69_), .C(x2), .Y(mai_mai_n1386_));
  NO2        m1337(.A(mai_mai_n1385_), .B(mai_mai_n1384_), .Y(mai_mai_n1387_));
  NO2        m1338(.A(mai_mai_n57_), .B(mai_mai_n96_), .Y(mai_mai_n1388_));
  AOI220     m1339(.A0(mai_mai_n734_), .A1(mai_mai_n745_), .B0(mai_mai_n503_), .B1(mai_mai_n267_), .Y(mai_mai_n1389_));
  NO2        m1340(.A(mai_mai_n1389_), .B(mai_mai_n1236_), .Y(mai_mai_n1390_));
  NO3        m1341(.A(mai_mai_n523_), .B(mai_mai_n162_), .C(mai_mai_n1002_), .Y(mai_mai_n1391_));
  NA2        m1342(.A(mai_mai_n901_), .B(x4), .Y(mai_mai_n1392_));
  OAI220     m1343(.A0(mai_mai_n1392_), .A1(mai_mai_n668_), .B0(mai_mai_n631_), .B1(mai_mai_n594_), .Y(mai_mai_n1393_));
  NO3        m1344(.A(mai_mai_n1393_), .B(mai_mai_n1391_), .C(mai_mai_n1390_), .Y(mai_mai_n1394_));
  OAI210     m1345(.A0(mai_mai_n1387_), .A1(x5), .B0(mai_mai_n1394_), .Y(mai_mai_n1395_));
  AOI220     m1346(.A0(mai_mai_n1395_), .A1(mai_mai_n90_), .B0(mai_mai_n1381_), .B1(mai_mai_n328_), .Y(mai_mai_n1396_));
  NA4        m1347(.A(mai_mai_n1396_), .B(mai_mai_n1365_), .C(mai_mai_n1343_), .D(mai_mai_n1326_), .Y(mai17));
  NO4        m1348(.A(mai_mai_n587_), .B(mai_mai_n681_), .C(mai_mai_n93_), .D(mai_mai_n92_), .Y(mai_mai_n1398_));
  NO2        m1349(.A(mai_mai_n114_), .B(mai_mai_n1105_), .Y(mai_mai_n1399_));
  AOI220     m1350(.A0(mai_mai_n1399_), .A1(mai_mai_n689_), .B0(mai_mai_n1398_), .B1(mai_mai_n494_), .Y(mai_mai_n1400_));
  NA2        m1351(.A(mai_mai_n153_), .B(mai_mai_n72_), .Y(mai_mai_n1401_));
  INV        m1352(.A(mai_mai_n76_), .Y(mai_mai_n1402_));
  OAI210     m1353(.A0(mai_mai_n608_), .A1(mai_mai_n55_), .B0(mai_mai_n1402_), .Y(mai_mai_n1403_));
  NA2        m1354(.A(mai_mai_n1155_), .B(mai_mai_n963_), .Y(mai_mai_n1404_));
  NA4        m1355(.A(mai_mai_n1404_), .B(mai_mai_n1403_), .C(mai_mai_n706_), .D(mai_mai_n57_), .Y(mai_mai_n1405_));
  OA210      m1356(.A0(mai_mai_n1247_), .A1(mai_mai_n1098_), .B0(mai_mai_n724_), .Y(mai_mai_n1406_));
  NA2        m1357(.A(mai_mai_n1406_), .B(mai_mai_n1405_), .Y(mai_mai_n1407_));
  NA3        m1358(.A(mai_mai_n152_), .B(mai_mai_n614_), .C(mai_mai_n1002_), .Y(mai_mai_n1408_));
  AOI210     m1359(.A0(mai_mai_n1025_), .A1(mai_mai_n293_), .B0(mai_mai_n59_), .Y(mai_mai_n1409_));
  NA2        m1360(.A(mai_mai_n1409_), .B(mai_mai_n1408_), .Y(mai_mai_n1410_));
  AOI210     m1361(.A0(mai_mai_n1407_), .A1(x1), .B0(mai_mai_n1410_), .Y(mai_mai_n1411_));
  NO2        m1362(.A(mai_mai_n616_), .B(mai_mai_n514_), .Y(mai_mai_n1412_));
  OAI210     m1363(.A0(mai_mai_n1412_), .A1(mai_mai_n862_), .B0(mai_mai_n1348_), .Y(mai_mai_n1413_));
  NO2        m1364(.A(mai_mai_n1413_), .B(x8), .Y(mai_mai_n1414_));
  NA3        m1365(.A(mai_mai_n616_), .B(mai_mai_n259_), .C(mai_mai_n111_), .Y(mai_mai_n1415_));
  NO2        m1366(.A(mai_mai_n134_), .B(mai_mai_n132_), .Y(mai_mai_n1416_));
  NO3        m1367(.A(mai_mai_n857_), .B(mai_mai_n745_), .C(mai_mai_n681_), .Y(mai_mai_n1417_));
  AOI210     m1368(.A0(mai_mai_n1417_), .A1(mai_mai_n1416_), .B0(x0), .Y(mai_mai_n1418_));
  OAI210     m1369(.A0(mai_mai_n1415_), .A1(mai_mai_n235_), .B0(mai_mai_n1418_), .Y(mai_mai_n1419_));
  NO2        m1370(.A(mai_mai_n1419_), .B(mai_mai_n1414_), .Y(mai_mai_n1420_));
  OAI220     m1371(.A0(mai_mai_n1420_), .A1(mai_mai_n1411_), .B0(mai_mai_n1401_), .B1(mai_mai_n1400_), .Y(mai18));
  AOI210     m1372(.A0(x8), .A1(x0), .B0(x5), .Y(mai_mai_n1422_));
  NOi31      m1373(.An(mai_mai_n293_), .B(mai_mai_n1422_), .C(mai_mai_n1000_), .Y(mai_mai_n1423_));
  NA2        m1374(.A(mai_mai_n587_), .B(mai_mai_n59_), .Y(mai_mai_n1424_));
  AOI210     m1375(.A0(mai_mai_n1331_), .A1(mai_mai_n339_), .B0(mai_mai_n1424_), .Y(mai_mai_n1425_));
  NO2        m1376(.A(mai_mai_n601_), .B(mai_mai_n746_), .Y(mai_mai_n1426_));
  NO4        m1377(.A(mai_mai_n242_), .B(mai_mai_n776_), .C(mai_mai_n144_), .D(mai_mai_n66_), .Y(mai_mai_n1427_));
  NO4        m1378(.A(mai_mai_n1427_), .B(mai_mai_n1426_), .C(mai_mai_n1425_), .D(mai_mai_n1423_), .Y(mai_mai_n1428_));
  NA3        m1379(.A(mai_mai_n509_), .B(mai_mai_n206_), .C(x0), .Y(mai_mai_n1429_));
  NAi21      m1380(.An(mai_mai_n377_), .B(mai_mai_n1429_), .Y(mai_mai_n1430_));
  NO2        m1381(.A(mai_mai_n847_), .B(x5), .Y(mai_mai_n1431_));
  AOI210     m1382(.A0(mai_mai_n1083_), .A1(x5), .B0(mai_mai_n1431_), .Y(mai_mai_n1432_));
  OA220      m1383(.A0(mai_mai_n509_), .A1(mai_mai_n321_), .B0(mai_mai_n390_), .B1(x5), .Y(mai_mai_n1433_));
  OAI220     m1384(.A0(mai_mai_n1433_), .A1(mai_mai_n281_), .B0(mai_mai_n1432_), .B1(mai_mai_n204_), .Y(mai_mai_n1434_));
  AOI210     m1385(.A0(mai_mai_n1430_), .A1(mai_mai_n279_), .B0(mai_mai_n1434_), .Y(mai_mai_n1435_));
  AOI210     m1386(.A0(mai_mai_n1435_), .A1(mai_mai_n1428_), .B0(x6), .Y(mai_mai_n1436_));
  NA3        m1387(.A(mai_mai_n513_), .B(mai_mai_n411_), .C(x2), .Y(mai_mai_n1437_));
  NA3        m1388(.A(mai_mai_n1000_), .B(mai_mai_n51_), .C(mai_mai_n57_), .Y(mai_mai_n1438_));
  AOI210     m1389(.A0(mai_mai_n1438_), .A1(mai_mai_n1437_), .B0(mai_mai_n758_), .Y(mai_mai_n1439_));
  NA2        m1390(.A(mai_mai_n256_), .B(x6), .Y(mai_mai_n1440_));
  OAI210     m1391(.A0(mai_mai_n168_), .A1(mai_mai_n98_), .B0(mai_mai_n1089_), .Y(mai_mai_n1441_));
  NO2        m1392(.A(mai_mai_n1441_), .B(mai_mai_n1440_), .Y(mai_mai_n1442_));
  OAI210     m1393(.A0(mai_mai_n1442_), .A1(mai_mai_n1439_), .B0(mai_mai_n53_), .Y(mai_mai_n1443_));
  NO2        m1394(.A(mai_mai_n667_), .B(mai_mai_n249_), .Y(mai_mai_n1444_));
  NO2        m1395(.A(mai_mai_n252_), .B(x3), .Y(mai_mai_n1445_));
  NO3        m1396(.A(mai_mai_n425_), .B(mai_mai_n587_), .C(mai_mai_n799_), .Y(mai_mai_n1446_));
  OAI210     m1397(.A0(mai_mai_n1446_), .A1(mai_mai_n1444_), .B0(mai_mai_n1445_), .Y(mai_mai_n1447_));
  AOI210     m1398(.A0(mai_mai_n1092_), .A1(mai_mai_n600_), .B0(x4), .Y(mai_mai_n1448_));
  NA2        m1399(.A(mai_mai_n587_), .B(mai_mai_n59_), .Y(mai_mai_n1449_));
  OAI210     m1400(.A0(mai_mai_n608_), .A1(mai_mai_n633_), .B0(mai_mai_n1449_), .Y(mai_mai_n1450_));
  AO220      m1401(.A0(mai_mai_n1197_), .A1(mai_mai_n706_), .B0(mai_mai_n546_), .B1(mai_mai_n344_), .Y(mai_mai_n1451_));
  AOI220     m1402(.A0(mai_mai_n1451_), .A1(x1), .B0(mai_mai_n1450_), .B1(mai_mai_n150_), .Y(mai_mai_n1452_));
  NA4        m1403(.A(mai_mai_n1452_), .B(mai_mai_n1448_), .C(mai_mai_n1447_), .D(mai_mai_n1443_), .Y(mai_mai_n1453_));
  NO3        m1404(.A(mai_mai_n1016_), .B(mai_mai_n121_), .C(mai_mai_n120_), .Y(mai_mai_n1454_));
  OAI210     m1405(.A0(mai_mai_n1454_), .A1(mai_mai_n638_), .B0(mai_mai_n96_), .Y(mai_mai_n1455_));
  AOI210     m1406(.A0(mai_mai_n1455_), .A1(mai_mai_n551_), .B0(mai_mai_n758_), .Y(mai_mai_n1456_));
  NA3        m1407(.A(mai_mai_n1148_), .B(mai_mai_n180_), .C(mai_mai_n131_), .Y(mai_mai_n1457_));
  NA3        m1408(.A(mai_mai_n1019_), .B(mai_mai_n748_), .C(mai_mai_n332_), .Y(mai_mai_n1458_));
  NA2        m1409(.A(mai_mai_n160_), .B(mai_mai_n745_), .Y(mai_mai_n1459_));
  OAI210     m1410(.A0(mai_mai_n1459_), .A1(mai_mai_n1250_), .B0(mai_mai_n1458_), .Y(mai_mai_n1460_));
  AOI210     m1411(.A0(mai_mai_n1457_), .A1(mai_mai_n167_), .B0(mai_mai_n1460_), .Y(mai_mai_n1461_));
  OAI210     m1412(.A0(mai_mai_n1461_), .A1(mai_mai_n532_), .B0(x4), .Y(mai_mai_n1462_));
  OAI220     m1413(.A0(mai_mai_n1462_), .A1(mai_mai_n1456_), .B0(mai_mai_n1453_), .B1(mai_mai_n1436_), .Y(mai_mai_n1463_));
  NO2        m1414(.A(mai_mai_n137_), .B(mai_mai_n112_), .Y(mai_mai_n1464_));
  NO2        m1415(.A(mai_mai_n180_), .B(mai_mai_n768_), .Y(mai_mai_n1465_));
  NO2        m1416(.A(mai_mai_n376_), .B(mai_mai_n241_), .Y(mai_mai_n1466_));
  NO2        m1417(.A(mai_mai_n913_), .B(mai_mai_n573_), .Y(mai_mai_n1467_));
  AO220      m1418(.A0(mai_mai_n1467_), .A1(mai_mai_n57_), .B0(mai_mai_n1466_), .B1(mai_mai_n114_), .Y(mai_mai_n1468_));
  NO3        m1419(.A(mai_mai_n1468_), .B(mai_mai_n1465_), .C(mai_mai_n1464_), .Y(mai_mai_n1469_));
  NA2        m1420(.A(mai_mai_n1016_), .B(x3), .Y(mai_mai_n1470_));
  NO2        m1421(.A(mai_mai_n1469_), .B(x3), .Y(mai_mai_n1471_));
  NO3        m1422(.A(mai_mai_n953_), .B(mai_mai_n667_), .C(mai_mai_n316_), .Y(mai_mai_n1472_));
  AO210      m1423(.A0(mai_mai_n982_), .A1(mai_mai_n286_), .B0(mai_mai_n1472_), .Y(mai_mai_n1473_));
  AOI220     m1424(.A0(mai_mai_n1473_), .A1(x8), .B0(mai_mai_n1278_), .B1(mai_mai_n426_), .Y(mai_mai_n1474_));
  NA2        m1425(.A(mai_mai_n720_), .B(mai_mai_n307_), .Y(mai_mai_n1475_));
  NA2        m1426(.A(mai_mai_n1332_), .B(mai_mai_n98_), .Y(mai_mai_n1476_));
  NO3        m1427(.A(mai_mai_n1149_), .B(mai_mai_n947_), .C(mai_mai_n1089_), .Y(mai_mai_n1477_));
  NA2        m1428(.A(mai_mai_n1477_), .B(mai_mai_n1476_), .Y(mai_mai_n1478_));
  OA220      m1429(.A0(mai_mai_n1478_), .A1(mai_mai_n913_), .B0(mai_mai_n1475_), .B1(mai_mai_n560_), .Y(mai_mai_n1479_));
  OAI210     m1430(.A0(mai_mai_n1474_), .A1(mai_mai_n400_), .B0(mai_mai_n1479_), .Y(mai_mai_n1480_));
  AOI210     m1431(.A0(mai_mai_n1471_), .A1(mai_mai_n128_), .B0(mai_mai_n1480_), .Y(mai_mai_n1481_));
  NA2        m1432(.A(mai_mai_n1481_), .B(mai_mai_n1463_), .Y(mai19));
  NO2        m1433(.A(mai_mai_n1375_), .B(mai_mai_n245_), .Y(mai_mai_n1483_));
  NA2        m1434(.A(mai_mai_n633_), .B(x3), .Y(mai_mai_n1484_));
  OAI210     m1435(.A0(mai_mai_n144_), .A1(mai_mai_n97_), .B0(mai_mai_n73_), .Y(mai_mai_n1485_));
  NA3        m1436(.A(mai_mai_n1485_), .B(mai_mai_n1484_), .C(mai_mai_n228_), .Y(mai_mai_n1486_));
  NO2        m1437(.A(mai_mai_n1245_), .B(mai_mai_n160_), .Y(mai_mai_n1487_));
  AOI210     m1438(.A0(mai_mai_n1398_), .A1(mai_mai_n342_), .B0(mai_mai_n1487_), .Y(mai_mai_n1488_));
  AOI210     m1439(.A0(mai_mai_n1488_), .A1(mai_mai_n1486_), .B0(mai_mai_n56_), .Y(mai_mai_n1489_));
  NO2        m1440(.A(mai_mai_n822_), .B(mai_mai_n1160_), .Y(mai_mai_n1490_));
  OAI210     m1441(.A0(mai_mai_n1489_), .A1(mai_mai_n1483_), .B0(mai_mai_n1490_), .Y(mai_mai_n1491_));
  NOi21      m1442(.An(mai_mai_n595_), .B(mai_mai_n637_), .Y(mai_mai_n1492_));
  NO3        m1443(.A(mai_mai_n2514_), .B(mai_mai_n729_), .C(mai_mai_n116_), .Y(mai_mai_n1493_));
  NA2        m1444(.A(mai_mai_n1143_), .B(mai_mai_n112_), .Y(mai_mai_n1494_));
  NO4        m1445(.A(mai_mai_n1494_), .B(mai_mai_n953_), .C(mai_mai_n847_), .D(mai_mai_n71_), .Y(mai_mai_n1495_));
  NO3        m1446(.A(mai_mai_n1495_), .B(mai_mai_n1493_), .C(mai_mai_n979_), .Y(mai_mai_n1496_));
  NO2        m1447(.A(mai_mai_n532_), .B(mai_mai_n604_), .Y(mai_mai_n1497_));
  NO3        m1448(.A(mai_mai_n507_), .B(mai_mai_n295_), .C(mai_mai_n63_), .Y(mai_mai_n1498_));
  NA2        m1449(.A(mai_mai_n1498_), .B(x3), .Y(mai_mai_n1499_));
  OAI210     m1450(.A0(mai_mai_n1496_), .A1(mai_mai_n57_), .B0(mai_mai_n1499_), .Y(mai_mai_n1500_));
  AOI210     m1451(.A0(mai_mai_n1500_), .A1(mai_mai_n745_), .B0(mai_mai_n1492_), .Y(mai_mai_n1501_));
  AOI210     m1452(.A0(mai_mai_n786_), .A1(mai_mai_n707_), .B0(mai_mai_n735_), .Y(mai_mai_n1502_));
  NO2        m1453(.A(mai_mai_n1502_), .B(x4), .Y(mai_mai_n1503_));
  NA2        m1454(.A(mai_mai_n1328_), .B(mai_mai_n758_), .Y(mai_mai_n1504_));
  NO2        m1455(.A(mai_mai_n1504_), .B(mai_mai_n492_), .Y(mai_mai_n1505_));
  OAI210     m1456(.A0(mai_mai_n1505_), .A1(mai_mai_n1503_), .B0(mai_mai_n776_), .Y(mai_mai_n1506_));
  OR2        m1457(.A(mai_mai_n1506_), .B(x1), .Y(mai_mai_n1507_));
  NA2        m1458(.A(mai_mai_n1002_), .B(mai_mai_n1135_), .Y(mai_mai_n1508_));
  NA2        m1459(.A(mai_mai_n138_), .B(mai_mai_n99_), .Y(mai_mai_n1509_));
  NOi21      m1460(.An(x1), .B(x6), .Y(mai_mai_n1510_));
  NA2        m1461(.A(mai_mai_n1510_), .B(mai_mai_n76_), .Y(mai_mai_n1511_));
  NA3        m1462(.A(mai_mai_n1511_), .B(mai_mai_n1509_), .C(mai_mai_n1508_), .Y(mai_mai_n1512_));
  AOI220     m1463(.A0(mai_mai_n1512_), .A1(x3), .B0(mai_mai_n1150_), .B1(mai_mai_n372_), .Y(mai_mai_n1513_));
  AOI220     m1464(.A0(mai_mai_n1197_), .A1(mai_mai_n111_), .B0(mai_mai_n877_), .B1(mai_mai_n778_), .Y(mai_mai_n1514_));
  NO2        m1465(.A(mai_mai_n1514_), .B(mai_mai_n311_), .Y(mai_mai_n1515_));
  NA2        m1466(.A(mai_mai_n901_), .B(mai_mai_n50_), .Y(mai_mai_n1516_));
  NA3        m1467(.A(mai_mai_n1143_), .B(mai_mai_n373_), .C(mai_mai_n98_), .Y(mai_mai_n1517_));
  AOI210     m1468(.A0(mai_mai_n1517_), .A1(mai_mai_n1516_), .B0(mai_mai_n923_), .Y(mai_mai_n1518_));
  NO2        m1469(.A(mai_mai_n1518_), .B(mai_mai_n1515_), .Y(mai_mai_n1519_));
  OAI210     m1470(.A0(mai_mai_n1513_), .A1(mai_mai_n809_), .B0(mai_mai_n1519_), .Y(mai_mai_n1520_));
  INV        m1471(.A(mai_mai_n65_), .Y(mai_mai_n1521_));
  OAI220     m1472(.A0(mai_mai_n1521_), .A1(mai_mai_n1484_), .B0(mai_mai_n294_), .B1(mai_mai_n855_), .Y(mai_mai_n1522_));
  AOI220     m1473(.A0(mai_mai_n1522_), .A1(mai_mai_n56_), .B0(mai_mai_n1283_), .B1(mai_mai_n703_), .Y(mai_mai_n1523_));
  NO2        m1474(.A(mai_mai_n54_), .B(mai_mai_n67_), .Y(mai_mai_n1524_));
  AN2        m1475(.A(mai_mai_n778_), .B(mai_mai_n912_), .Y(mai_mai_n1525_));
  NA2        m1476(.A(mai_mai_n1127_), .B(mai_mai_n349_), .Y(mai_mai_n1526_));
  NO2        m1477(.A(mai_mai_n947_), .B(mai_mai_n1510_), .Y(mai_mai_n1527_));
  NA2        m1478(.A(mai_mai_n488_), .B(mai_mai_n703_), .Y(mai_mai_n1528_));
  OAI210     m1479(.A0(mai_mai_n1528_), .A1(mai_mai_n1527_), .B0(mai_mai_n1526_), .Y(mai_mai_n1529_));
  AOI210     m1480(.A0(mai_mai_n1525_), .A1(x2), .B0(mai_mai_n1529_), .Y(mai_mai_n1530_));
  OAI220     m1481(.A0(mai_mai_n1530_), .A1(mai_mai_n144_), .B0(mai_mai_n1523_), .B1(mai_mai_n54_), .Y(mai_mai_n1531_));
  OAI210     m1482(.A0(mai_mai_n1531_), .A1(mai_mai_n1520_), .B0(x8), .Y(mai_mai_n1532_));
  NA4        m1483(.A(mai_mai_n1532_), .B(mai_mai_n1507_), .C(mai_mai_n1501_), .D(mai_mai_n1491_), .Y(mai20));
  NA4        m1484(.A(mai_mai_n383_), .B(mai_mai_n267_), .C(mai_mai_n371_), .D(mai_mai_n61_), .Y(mai_mai_n1534_));
  NA2        m1485(.A(mai_mai_n467_), .B(mai_mai_n404_), .Y(mai_mai_n1535_));
  AOI210     m1486(.A0(mai_mai_n1535_), .A1(mai_mai_n1534_), .B0(mai_mai_n79_), .Y(mai_mai_n1536_));
  AOI210     m1487(.A0(mai_mai_n1006_), .A1(mai_mai_n61_), .B0(mai_mai_n1497_), .Y(mai_mai_n1537_));
  AOI210     m1488(.A0(mai_mai_n942_), .A1(mai_mai_n338_), .B0(mai_mai_n1133_), .Y(mai_mai_n1538_));
  OAI210     m1489(.A0(mai_mai_n1537_), .A1(mai_mai_n663_), .B0(mai_mai_n1538_), .Y(mai_mai_n1539_));
  OAI210     m1490(.A0(mai_mai_n1539_), .A1(mai_mai_n1536_), .B0(mai_mai_n1053_), .Y(mai_mai_n1540_));
  NAi21      m1491(.An(mai_mai_n541_), .B(mai_mai_n392_), .Y(mai_mai_n1541_));
  NA3        m1492(.A(mai_mai_n1541_), .B(mai_mai_n940_), .C(mai_mai_n912_), .Y(mai_mai_n1542_));
  NA3        m1493(.A(mai_mai_n1052_), .B(mai_mai_n267_), .C(mai_mai_n572_), .Y(mai_mai_n1543_));
  AOI210     m1494(.A0(mai_mai_n1543_), .A1(mai_mai_n1542_), .B0(mai_mai_n1236_), .Y(mai_mai_n1544_));
  NO2        m1495(.A(mai_mai_n720_), .B(mai_mai_n930_), .Y(mai_mai_n1545_));
  NA2        m1496(.A(mai_mai_n1544_), .B(mai_mai_n316_), .Y(mai_mai_n1546_));
  NO4        m1497(.A(mai_mai_n536_), .B(mai_mai_n223_), .C(x5), .D(x2), .Y(mai_mai_n1547_));
  NA2        m1498(.A(mai_mai_n307_), .B(mai_mai_n85_), .Y(mai_mai_n1548_));
  NA2        m1499(.A(mai_mai_n317_), .B(mai_mai_n96_), .Y(mai_mai_n1549_));
  NA2        m1500(.A(mai_mai_n414_), .B(mai_mai_n52_), .Y(mai_mai_n1550_));
  OAI220     m1501(.A0(mai_mai_n1550_), .A1(mai_mai_n1549_), .B0(mai_mai_n1548_), .B1(mai_mai_n262_), .Y(mai_mai_n1551_));
  OAI210     m1502(.A0(mai_mai_n1551_), .A1(mai_mai_n1547_), .B0(mai_mai_n212_), .Y(mai_mai_n1552_));
  NO2        m1503(.A(mai_mai_n650_), .B(mai_mai_n591_), .Y(mai_mai_n1553_));
  NA2        m1504(.A(mai_mai_n913_), .B(mai_mai_n50_), .Y(mai_mai_n1554_));
  NO3        m1505(.A(mai_mai_n1554_), .B(mai_mai_n355_), .C(mai_mai_n216_), .Y(mai_mai_n1555_));
  NO2        m1506(.A(mai_mai_n1392_), .B(mai_mai_n990_), .Y(mai_mai_n1556_));
  AOI210     m1507(.A0(mai_mai_n1555_), .A1(mai_mai_n1553_), .B0(mai_mai_n1556_), .Y(mai_mai_n1557_));
  NA4        m1508(.A(mai_mai_n1557_), .B(mai_mai_n1552_), .C(mai_mai_n1546_), .D(mai_mai_n1540_), .Y(mai21));
  NO2        m1509(.A(mai_mai_n1007_), .B(mai_mai_n88_), .Y(mai_mai_n1559_));
  NA2        m1510(.A(mai_mai_n1559_), .B(mai_mai_n72_), .Y(mai_mai_n1560_));
  NA2        m1511(.A(mai_mai_n279_), .B(mai_mai_n820_), .Y(mai_mai_n1561_));
  AOI220     m1512(.A0(mai_mai_n1561_), .A1(mai_mai_n297_), .B0(mai_mai_n560_), .B1(mai_mai_n451_), .Y(mai_mai_n1562_));
  NA2        m1513(.A(mai_mai_n901_), .B(mai_mai_n261_), .Y(mai_mai_n1563_));
  NA2        m1514(.A(mai_mai_n527_), .B(mai_mai_n452_), .Y(mai_mai_n1564_));
  NA3        m1515(.A(mai_mai_n1563_), .B(mai_mai_n1308_), .C(mai_mai_n56_), .Y(mai_mai_n1565_));
  NO2        m1516(.A(mai_mai_n748_), .B(mai_mai_n425_), .Y(mai_mai_n1566_));
  NO3        m1517(.A(mai_mai_n1566_), .B(mai_mai_n695_), .C(mai_mai_n237_), .Y(mai_mai_n1567_));
  NOi31      m1518(.An(mai_mai_n183_), .B(mai_mai_n616_), .C(mai_mai_n1037_), .Y(mai_mai_n1568_));
  NO4        m1519(.A(mai_mai_n1568_), .B(mai_mai_n1567_), .C(mai_mai_n1565_), .D(mai_mai_n1562_), .Y(mai_mai_n1569_));
  AN2        m1520(.A(mai_mai_n845_), .B(x3), .Y(mai_mai_n1570_));
  NO2        m1521(.A(mai_mai_n66_), .B(x2), .Y(mai_mai_n1571_));
  OAI210     m1522(.A0(mai_mai_n167_), .A1(x0), .B0(mai_mai_n1571_), .Y(mai_mai_n1572_));
  NA2        m1523(.A(mai_mai_n135_), .B(mai_mai_n96_), .Y(mai_mai_n1573_));
  NA2        m1524(.A(mai_mai_n1573_), .B(mai_mai_n1572_), .Y(mai_mai_n1574_));
  OAI210     m1525(.A0(mai_mai_n1574_), .A1(mai_mai_n1570_), .B0(x8), .Y(mai_mai_n1575_));
  NO3        m1526(.A(mai_mai_n746_), .B(mai_mai_n605_), .C(mai_mai_n573_), .Y(mai_mai_n1576_));
  NA2        m1527(.A(mai_mai_n55_), .B(mai_mai_n50_), .Y(mai_mai_n1577_));
  MUX2       m1528(.S(mai_mai_n587_), .A(mai_mai_n1577_), .B(mai_mai_n95_), .Y(mai_mai_n1578_));
  AOI210     m1529(.A0(mai_mai_n1288_), .A1(mai_mai_n226_), .B0(mai_mai_n1578_), .Y(mai_mai_n1579_));
  OAI210     m1530(.A0(mai_mai_n629_), .A1(mai_mai_n572_), .B0(x4), .Y(mai_mai_n1580_));
  NO3        m1531(.A(mai_mai_n1580_), .B(mai_mai_n1579_), .C(mai_mai_n1576_), .Y(mai_mai_n1581_));
  AO220      m1532(.A0(mai_mai_n1581_), .A1(mai_mai_n1575_), .B0(mai_mai_n1569_), .B1(mai_mai_n1560_), .Y(mai_mai_n1582_));
  AN2        m1533(.A(mai_mai_n617_), .B(mai_mai_n311_), .Y(mai_mai_n1583_));
  NO2        m1534(.A(mai_mai_n822_), .B(x0), .Y(mai_mai_n1584_));
  NO3        m1535(.A(mai_mai_n1584_), .B(mai_mai_n537_), .C(mai_mai_n80_), .Y(mai_mai_n1585_));
  NO2        m1536(.A(mai_mai_n149_), .B(x2), .Y(mai_mai_n1586_));
  NO3        m1537(.A(mai_mai_n368_), .B(mai_mai_n242_), .C(mai_mai_n175_), .Y(mai_mai_n1587_));
  AOI210     m1538(.A0(mai_mai_n1586_), .A1(mai_mai_n65_), .B0(mai_mai_n1587_), .Y(mai_mai_n1588_));
  OAI210     m1539(.A0(mai_mai_n1585_), .A1(mai_mai_n390_), .B0(mai_mai_n1588_), .Y(mai_mai_n1589_));
  AOI220     m1540(.A0(mai_mai_n1589_), .A1(x5), .B0(mai_mai_n1583_), .B1(mai_mai_n720_), .Y(mai_mai_n1590_));
  AOI210     m1541(.A0(mai_mai_n1590_), .A1(mai_mai_n1582_), .B0(mai_mai_n67_), .Y(mai_mai_n1591_));
  NO2        m1542(.A(mai_mai_n867_), .B(mai_mai_n158_), .Y(mai_mai_n1592_));
  NOi41      m1543(.An(mai_mai_n1361_), .B(mai_mai_n1422_), .C(mai_mai_n1104_), .D(mai_mai_n813_), .Y(mai_mai_n1593_));
  NA2        m1544(.A(mai_mai_n1593_), .B(mai_mai_n1592_), .Y(mai_mai_n1594_));
  NO2        m1545(.A(mai_mai_n72_), .B(x4), .Y(mai_mai_n1595_));
  OAI210     m1546(.A0(mai_mai_n277_), .A1(mai_mai_n148_), .B0(mai_mai_n1595_), .Y(mai_mai_n1596_));
  OAI210     m1547(.A0(mai_mai_n399_), .A1(mai_mai_n415_), .B0(mai_mai_n216_), .Y(mai_mai_n1597_));
  NO2        m1548(.A(mai_mai_n244_), .B(mai_mai_n50_), .Y(mai_mai_n1598_));
  NO2        m1549(.A(mai_mai_n1598_), .B(mai_mai_n57_), .Y(mai_mai_n1599_));
  NA2        m1550(.A(mai_mai_n1599_), .B(mai_mai_n1597_), .Y(mai_mai_n1600_));
  AOI210     m1551(.A0(mai_mai_n1596_), .A1(mai_mai_n1594_), .B0(mai_mai_n1600_), .Y(mai_mai_n1601_));
  NA2        m1552(.A(mai_mai_n732_), .B(mai_mai_n541_), .Y(mai_mai_n1602_));
  AO210      m1553(.A0(mai_mai_n1602_), .A1(mai_mai_n923_), .B0(mai_mai_n50_), .Y(mai_mai_n1603_));
  NO2        m1554(.A(mai_mai_n1541_), .B(mai_mai_n1160_), .Y(mai_mai_n1604_));
  NA2        m1555(.A(mai_mai_n1604_), .B(mai_mai_n1114_), .Y(mai_mai_n1605_));
  AOI210     m1556(.A0(mai_mai_n1605_), .A1(mai_mai_n1603_), .B0(mai_mai_n98_), .Y(mai_mai_n1606_));
  NA2        m1557(.A(mai_mai_n286_), .B(mai_mai_n96_), .Y(mai_mai_n1607_));
  NA2        m1558(.A(mai_mai_n854_), .B(mai_mai_n55_), .Y(mai_mai_n1608_));
  NO2        m1559(.A(mai_mai_n1608_), .B(mai_mai_n1607_), .Y(mai_mai_n1609_));
  NO2        m1560(.A(mai_mai_n653_), .B(mai_mai_n1010_), .Y(mai_mai_n1610_));
  NO4        m1561(.A(mai_mai_n1610_), .B(mai_mai_n1609_), .C(mai_mai_n1606_), .D(mai_mai_n1601_), .Y(mai_mai_n1611_));
  NO2        m1562(.A(mai_mai_n1611_), .B(x6), .Y(mai_mai_n1612_));
  AOI210     m1563(.A0(mai_mai_n594_), .A1(mai_mai_n1010_), .B0(mai_mai_n1422_), .Y(mai_mai_n1613_));
  OAI210     m1564(.A0(mai_mai_n1613_), .A1(mai_mai_n670_), .B0(mai_mai_n56_), .Y(mai_mai_n1614_));
  NO2        m1565(.A(mai_mai_n722_), .B(mai_mai_n54_), .Y(mai_mai_n1615_));
  NO4        m1566(.A(mai_mai_n921_), .B(mai_mai_n265_), .C(mai_mai_n745_), .D(mai_mai_n729_), .Y(mai_mai_n1616_));
  NO2        m1567(.A(mai_mai_n825_), .B(x5), .Y(mai_mai_n1617_));
  NO4        m1568(.A(mai_mai_n1617_), .B(mai_mai_n1616_), .C(mai_mai_n1615_), .D(mai_mai_n906_), .Y(mai_mai_n1618_));
  AOI210     m1569(.A0(mai_mai_n1618_), .A1(mai_mai_n1614_), .B0(mai_mai_n50_), .Y(mai_mai_n1619_));
  NA2        m1570(.A(mai_mai_n149_), .B(mai_mai_n96_), .Y(mai_mai_n1620_));
  OA220      m1571(.A0(mai_mai_n1620_), .A1(mai_mai_n429_), .B0(mai_mai_n457_), .B1(mai_mai_n720_), .Y(mai_mai_n1621_));
  NA3        m1572(.A(mai_mai_n55_), .B(x2), .C(x0), .Y(mai_mai_n1622_));
  AOI220     m1573(.A0(mai_mai_n1622_), .A1(mai_mai_n160_), .B0(mai_mai_n825_), .B1(mai_mai_n146_), .Y(mai_mai_n1623_));
  NO2        m1574(.A(mai_mai_n663_), .B(mai_mai_n244_), .Y(mai_mai_n1624_));
  NO3        m1575(.A(mai_mai_n232_), .B(mai_mai_n214_), .C(mai_mai_n349_), .Y(mai_mai_n1625_));
  NO3        m1576(.A(mai_mai_n1625_), .B(mai_mai_n1624_), .C(mai_mai_n1623_), .Y(mai_mai_n1626_));
  OAI220     m1577(.A0(mai_mai_n1626_), .A1(mai_mai_n56_), .B0(mai_mai_n1621_), .B1(mai_mai_n679_), .Y(mai_mai_n1627_));
  OAI210     m1578(.A0(mai_mai_n1627_), .A1(mai_mai_n1619_), .B0(mai_mai_n104_), .Y(mai_mai_n1628_));
  NO2        m1579(.A(mai_mai_n599_), .B(mai_mai_n292_), .Y(mai_mai_n1629_));
  AOI210     m1580(.A0(mai_mai_n592_), .A1(x5), .B0(mai_mai_n1629_), .Y(mai_mai_n1630_));
  NO2        m1581(.A(mai_mai_n1630_), .B(mai_mai_n98_), .Y(mai_mai_n1631_));
  NA2        m1582(.A(mai_mai_n687_), .B(mai_mai_n73_), .Y(mai_mai_n1632_));
  NA3        m1583(.A(mai_mai_n1632_), .B(mai_mai_n422_), .C(mai_mai_n57_), .Y(mai_mai_n1633_));
  OAI210     m1584(.A0(mai_mai_n1608_), .A1(mai_mai_n1607_), .B0(mai_mai_n1633_), .Y(mai_mai_n1634_));
  OAI210     m1585(.A0(mai_mai_n1634_), .A1(mai_mai_n1631_), .B0(x1), .Y(mai_mai_n1635_));
  NO4        m1586(.A(mai_mai_n408_), .B(mai_mai_n72_), .C(mai_mai_n139_), .D(x3), .Y(mai_mai_n1636_));
  NO2        m1587(.A(mai_mai_n317_), .B(mai_mai_n100_), .Y(mai_mai_n1637_));
  OAI210     m1588(.A0(mai_mai_n1636_), .A1(mai_mai_n1237_), .B0(mai_mai_n1637_), .Y(mai_mai_n1638_));
  NO2        m1589(.A(mai_mai_n60_), .B(mai_mai_n96_), .Y(mai_mai_n1639_));
  NO4        m1590(.A(mai_mai_n1607_), .B(mai_mai_n921_), .C(mai_mai_n650_), .D(mai_mai_n50_), .Y(mai_mai_n1640_));
  AOI210     m1591(.A0(mai_mai_n1639_), .A1(mai_mai_n1465_), .B0(mai_mai_n1640_), .Y(mai_mai_n1641_));
  NA4        m1592(.A(mai_mai_n1641_), .B(mai_mai_n1638_), .C(mai_mai_n1635_), .D(mai_mai_n1628_), .Y(mai_mai_n1642_));
  NO3        m1593(.A(mai_mai_n1642_), .B(mai_mai_n1612_), .C(mai_mai_n1591_), .Y(mai22));
  AOI210     m1594(.A0(mai_mai_n513_), .A1(mai_mai_n67_), .B0(mai_mai_n460_), .Y(mai_mai_n1644_));
  AOI210     m1595(.A0(x5), .A1(x2), .B0(x8), .Y(mai_mai_n1645_));
  NA2        m1596(.A(mai_mai_n1645_), .B(mai_mai_n59_), .Y(mai_mai_n1646_));
  OAI220     m1597(.A0(mai_mai_n1646_), .A1(mai_mai_n308_), .B0(mai_mai_n1644_), .B1(mai_mai_n390_), .Y(mai_mai_n1647_));
  NA2        m1598(.A(mai_mai_n262_), .B(mai_mai_n71_), .Y(mai_mai_n1648_));
  OA220      m1599(.A0(mai_mai_n1648_), .A1(mai_mai_n59_), .B0(mai_mai_n806_), .B1(mai_mai_n963_), .Y(mai_mai_n1649_));
  NO4        m1600(.A(mai_mai_n376_), .B(mai_mai_n210_), .C(mai_mai_n67_), .D(x3), .Y(mai_mai_n1650_));
  NO3        m1601(.A(mai_mai_n1188_), .B(mai_mai_n79_), .C(x0), .Y(mai_mai_n1651_));
  OAI210     m1602(.A0(mai_mai_n390_), .A1(mai_mai_n195_), .B0(x4), .Y(mai_mai_n1652_));
  NO3        m1603(.A(mai_mai_n1652_), .B(mai_mai_n1651_), .C(mai_mai_n1650_), .Y(mai_mai_n1653_));
  OAI210     m1604(.A0(mai_mai_n1649_), .A1(mai_mai_n188_), .B0(mai_mai_n1653_), .Y(mai_mai_n1654_));
  AOI210     m1605(.A0(mai_mai_n1647_), .A1(mai_mai_n53_), .B0(mai_mai_n1654_), .Y(mai_mai_n1655_));
  NA2        m1606(.A(mai_mai_n290_), .B(mai_mai_n295_), .Y(mai_mai_n1656_));
  NA3        m1607(.A(mai_mai_n1656_), .B(mai_mai_n212_), .C(mai_mai_n294_), .Y(mai_mai_n1657_));
  NA2        m1608(.A(mai_mai_n568_), .B(mai_mai_n231_), .Y(mai_mai_n1658_));
  NO3        m1609(.A(mai_mai_n488_), .B(mai_mai_n252_), .C(mai_mai_n204_), .Y(mai_mai_n1659_));
  NAi31      m1610(.An(mai_mai_n1659_), .B(mai_mai_n1658_), .C(mai_mai_n1657_), .Y(mai_mai_n1660_));
  NO2        m1611(.A(mai_mai_n457_), .B(mai_mai_n246_), .Y(mai_mai_n1661_));
  NO2        m1612(.A(mai_mai_n1188_), .B(x3), .Y(mai_mai_n1662_));
  AOI210     m1613(.A0(mai_mai_n1662_), .A1(mai_mai_n338_), .B0(mai_mai_n1661_), .Y(mai_mai_n1663_));
  OAI210     m1614(.A0(mai_mai_n1032_), .A1(mai_mai_n177_), .B0(mai_mai_n56_), .Y(mai_mai_n1664_));
  NA3        m1615(.A(mai_mai_n55_), .B(mai_mai_n67_), .C(x0), .Y(mai_mai_n1665_));
  OAI220     m1616(.A0(mai_mai_n1665_), .A1(mai_mai_n1010_), .B0(mai_mai_n355_), .B1(mai_mai_n203_), .Y(mai_mai_n1666_));
  NO2        m1617(.A(mai_mai_n1666_), .B(mai_mai_n1664_), .Y(mai_mai_n1667_));
  OAI210     m1618(.A0(mai_mai_n1663_), .A1(mai_mai_n244_), .B0(mai_mai_n1667_), .Y(mai_mai_n1668_));
  AOI210     m1619(.A0(mai_mai_n1660_), .A1(mai_mai_n96_), .B0(mai_mai_n1668_), .Y(mai_mai_n1669_));
  AOI210     m1620(.A0(mai_mai_n910_), .A1(mai_mai_n747_), .B0(mai_mai_n828_), .Y(mai_mai_n1670_));
  OAI210     m1621(.A0(mai_mai_n770_), .A1(mai_mai_n149_), .B0(mai_mai_n898_), .Y(mai_mai_n1671_));
  OAI210     m1622(.A0(mai_mai_n1671_), .A1(mai_mai_n1670_), .B0(mai_mai_n598_), .Y(mai_mai_n1672_));
  OA210      m1623(.A0(mai_mai_n1669_), .A1(mai_mai_n1655_), .B0(mai_mai_n1672_), .Y(mai_mai_n1673_));
  OAI210     m1624(.A0(mai_mai_n1121_), .A1(mai_mai_n686_), .B0(mai_mai_n674_), .Y(mai_mai_n1674_));
  NO2        m1625(.A(mai_mai_n343_), .B(x0), .Y(mai_mai_n1675_));
  NA3        m1626(.A(mai_mai_n1675_), .B(mai_mai_n338_), .C(mai_mai_n56_), .Y(mai_mai_n1676_));
  AOI210     m1627(.A0(mai_mai_n1676_), .A1(mai_mai_n1674_), .B0(mai_mai_n390_), .Y(mai_mai_n1677_));
  NO3        m1628(.A(mai_mai_n160_), .B(mai_mai_n149_), .C(mai_mai_n61_), .Y(mai_mai_n1678_));
  OAI210     m1629(.A0(mai_mai_n1678_), .A1(mai_mai_n410_), .B0(mai_mai_n98_), .Y(mai_mai_n1679_));
  NA2        m1630(.A(mai_mai_n131_), .B(mai_mai_n758_), .Y(mai_mai_n1680_));
  NA2        m1631(.A(mai_mai_n408_), .B(x3), .Y(mai_mai_n1681_));
  NAi31      m1632(.An(mai_mai_n1681_), .B(mai_mai_n1680_), .C(mai_mai_n1476_), .Y(mai_mai_n1682_));
  NO3        m1633(.A(mai_mai_n822_), .B(mai_mai_n456_), .C(mai_mai_n98_), .Y(mai_mai_n1683_));
  NO2        m1634(.A(mai_mai_n1034_), .B(mai_mai_n132_), .Y(mai_mai_n1684_));
  NO3        m1635(.A(mai_mai_n857_), .B(mai_mai_n404_), .C(mai_mai_n291_), .Y(mai_mai_n1685_));
  AOI220     m1636(.A0(mai_mai_n1685_), .A1(mai_mai_n1684_), .B0(mai_mai_n1683_), .B1(mai_mai_n1675_), .Y(mai_mai_n1686_));
  NA3        m1637(.A(mai_mai_n56_), .B(mai_mai_n50_), .C(x0), .Y(mai_mai_n1687_));
  NOi21      m1638(.An(mai_mai_n75_), .B(mai_mai_n706_), .Y(mai_mai_n1688_));
  NA2        m1639(.A(mai_mai_n947_), .B(mai_mai_n253_), .Y(mai_mai_n1689_));
  NO2        m1640(.A(mai_mai_n1689_), .B(mai_mai_n1688_), .Y(mai_mai_n1690_));
  NA2        m1641(.A(mai_mai_n1690_), .B(mai_mai_n1019_), .Y(mai_mai_n1691_));
  NA4        m1642(.A(mai_mai_n1691_), .B(mai_mai_n1686_), .C(mai_mai_n1682_), .D(mai_mai_n1679_), .Y(mai_mai_n1692_));
  AOI210     m1643(.A0(mai_mai_n1692_), .A1(x7), .B0(mai_mai_n1677_), .Y(mai_mai_n1693_));
  OAI210     m1644(.A0(mai_mai_n1673_), .A1(x7), .B0(mai_mai_n1693_), .Y(mai23));
  OR2        m1645(.A(mai_mai_n507_), .B(mai_mai_n212_), .Y(mai_mai_n1695_));
  AOI220     m1646(.A0(mai_mai_n1695_), .A1(mai_mai_n1545_), .B0(mai_mai_n600_), .B1(mai_mai_n282_), .Y(mai_mai_n1696_));
  NO3        m1647(.A(mai_mai_n806_), .B(mai_mai_n581_), .C(mai_mai_n479_), .Y(mai_mai_n1697_));
  INV        m1648(.A(mai_mai_n1697_), .Y(mai_mai_n1698_));
  OAI210     m1649(.A0(mai_mai_n1696_), .A1(mai_mai_n144_), .B0(mai_mai_n1698_), .Y(mai_mai_n1699_));
  NA2        m1650(.A(mai_mai_n1699_), .B(mai_mai_n55_), .Y(mai_mai_n1700_));
  NO2        m1651(.A(mai_mai_n921_), .B(mai_mai_n505_), .Y(mai_mai_n1701_));
  AO220      m1652(.A0(mai_mai_n1221_), .A1(mai_mai_n171_), .B0(mai_mai_n953_), .B1(mai_mai_n720_), .Y(mai_mai_n1702_));
  OAI210     m1653(.A0(mai_mai_n1702_), .A1(mai_mai_n1701_), .B0(mai_mai_n578_), .Y(mai_mai_n1703_));
  NA2        m1654(.A(mai_mai_n168_), .B(mai_mai_n158_), .Y(mai_mai_n1704_));
  NA2        m1655(.A(mai_mai_n396_), .B(mai_mai_n150_), .Y(mai_mai_n1705_));
  AOI210     m1656(.A0(mai_mai_n1705_), .A1(mai_mai_n1704_), .B0(mai_mai_n223_), .Y(mai_mai_n1706_));
  NA2        m1657(.A(mai_mai_n415_), .B(mai_mai_n244_), .Y(mai_mai_n1707_));
  AOI210     m1658(.A0(mai_mai_n1707_), .A1(mai_mai_n490_), .B0(mai_mai_n373_), .Y(mai_mai_n1708_));
  OAI210     m1659(.A0(mai_mai_n1708_), .A1(mai_mai_n1706_), .B0(mai_mai_n286_), .Y(mai_mai_n1709_));
  NA3        m1660(.A(mai_mai_n57_), .B(x4), .C(x3), .Y(mai_mai_n1710_));
  NO3        m1661(.A(mai_mai_n1710_), .B(mai_mai_n718_), .C(mai_mai_n131_), .Y(mai_mai_n1711_));
  AOI210     m1662(.A0(mai_mai_n881_), .A1(mai_mai_n133_), .B0(mai_mai_n1711_), .Y(mai_mai_n1712_));
  NA4        m1663(.A(mai_mai_n1712_), .B(mai_mai_n1709_), .C(mai_mai_n1703_), .D(mai_mai_n1700_), .Y(mai24));
  NO2        m1664(.A(mai_mai_n228_), .B(x1), .Y(mai_mai_n1714_));
  NA2        m1665(.A(mai_mai_n328_), .B(mai_mai_n483_), .Y(mai_mai_n1715_));
  INV        m1666(.A(mai_mai_n1715_), .Y(mai_mai_n1716_));
  NA2        m1667(.A(mai_mai_n1716_), .B(mai_mai_n85_), .Y(mai_mai_n1717_));
  NA2        m1668(.A(mai_mai_n93_), .B(x8), .Y(mai_mai_n1718_));
  NO3        m1669(.A(mai_mai_n1016_), .B(mai_mai_n1271_), .C(mai_mai_n1002_), .Y(mai_mai_n1719_));
  NA2        m1670(.A(mai_mai_n940_), .B(mai_mai_n56_), .Y(mai_mai_n1720_));
  AO220      m1671(.A0(mai_mai_n1720_), .A1(mai_mai_n1719_), .B0(mai_mai_n1209_), .B1(mai_mai_n316_), .Y(mai_mai_n1721_));
  NA2        m1672(.A(mai_mai_n446_), .B(x8), .Y(mai_mai_n1722_));
  NA2        m1673(.A(mai_mai_n651_), .B(mai_mai_n114_), .Y(mai_mai_n1723_));
  NO2        m1674(.A(mai_mai_n1723_), .B(mai_mai_n1367_), .Y(mai_mai_n1724_));
  AOI220     m1675(.A0(mai_mai_n1724_), .A1(mai_mai_n1598_), .B0(mai_mai_n1721_), .B1(mai_mai_n985_), .Y(mai_mai_n1725_));
  OAI210     m1676(.A0(mai_mai_n1718_), .A1(mai_mai_n1717_), .B0(mai_mai_n1725_), .Y(mai25));
  NA2        m1677(.A(mai_mai_n317_), .B(mai_mai_n59_), .Y(mai_mai_n1727_));
  NO2        m1678(.A(mai_mai_n1727_), .B(mai_mai_n308_), .Y(mai_mai_n1728_));
  OAI210     m1679(.A0(mai_mai_n1728_), .A1(mai_mai_n1128_), .B0(mai_mai_n104_), .Y(mai_mai_n1729_));
  INV        m1680(.A(mai_mai_n1217_), .Y(mai_mai_n1730_));
  AOI220     m1681(.A0(x6), .A1(mai_mai_n1730_), .B0(mai_mai_n2516_), .B1(mai_mai_n1129_), .Y(mai_mai_n1731_));
  AOI210     m1682(.A0(mai_mai_n1731_), .A1(mai_mai_n1729_), .B0(mai_mai_n661_), .Y(mai_mai_n1732_));
  NO3        m1683(.A(mai_mai_n995_), .B(mai_mai_n134_), .C(mai_mai_n72_), .Y(mai_mai_n1733_));
  OAI210     m1684(.A0(mai_mai_n188_), .A1(mai_mai_n262_), .B0(mai_mai_n318_), .Y(mai_mai_n1734_));
  OAI210     m1685(.A0(mai_mai_n1734_), .A1(mai_mai_n1733_), .B0(mai_mai_n1127_), .Y(mai_mai_n1735_));
  NA2        m1686(.A(mai_mai_n500_), .B(mai_mai_n55_), .Y(mai_mai_n1736_));
  OAI220     m1687(.A0(mai_mai_n1736_), .A1(mai_mai_n228_), .B0(mai_mai_n575_), .B1(mai_mai_n262_), .Y(mai_mai_n1737_));
  NA2        m1688(.A(mai_mai_n1737_), .B(mai_mai_n621_), .Y(mai_mai_n1738_));
  NA2        m1689(.A(mai_mai_n1416_), .B(mai_mai_n369_), .Y(mai_mai_n1739_));
  NA3        m1690(.A(mai_mai_n1739_), .B(mai_mai_n1738_), .C(mai_mai_n1735_), .Y(mai_mai_n1740_));
  AO210      m1691(.A0(mai_mai_n1740_), .A1(mai_mai_n96_), .B0(mai_mai_n1732_), .Y(mai26));
  NA2        m1692(.A(mai_mai_n745_), .B(mai_mai_n50_), .Y(mai_mai_n1742_));
  NA2        m1693(.A(mai_mai_n1237_), .B(mai_mai_n1089_), .Y(mai_mai_n1743_));
  NA2        m1694(.A(mai_mai_n609_), .B(mai_mai_n568_), .Y(mai_mai_n1744_));
  NA2        m1695(.A(mai_mai_n976_), .B(mai_mai_n573_), .Y(mai_mai_n1745_));
  NO2        m1696(.A(mai_mai_n1745_), .B(mai_mai_n1193_), .Y(mai_mai_n1746_));
  AOI210     m1697(.A0(mai_mai_n1684_), .A1(mai_mai_n1388_), .B0(mai_mai_n1746_), .Y(mai_mai_n1747_));
  NO2        m1698(.A(mai_mai_n1034_), .B(mai_mai_n69_), .Y(mai_mai_n1748_));
  NA2        m1699(.A(mai_mai_n776_), .B(mai_mai_n167_), .Y(mai_mai_n1749_));
  NO2        m1700(.A(mai_mai_n1749_), .B(mai_mai_n528_), .Y(mai_mai_n1750_));
  AOI210     m1701(.A0(mai_mai_n1748_), .A1(mai_mai_n574_), .B0(mai_mai_n1750_), .Y(mai_mai_n1751_));
  OAI220     m1702(.A0(mai_mai_n1751_), .A1(mai_mai_n96_), .B0(mai_mai_n1747_), .B1(mai_mai_n53_), .Y(mai_mai_n1752_));
  NA2        m1703(.A(mai_mai_n588_), .B(mai_mai_n500_), .Y(mai_mai_n1753_));
  NO2        m1704(.A(mai_mai_n124_), .B(mai_mai_n121_), .Y(mai_mai_n1754_));
  NA2        m1705(.A(mai_mai_n1754_), .B(mai_mai_n111_), .Y(mai_mai_n1755_));
  NA2        m1706(.A(mai_mai_n720_), .B(x3), .Y(mai_mai_n1756_));
  AOI210     m1707(.A0(mai_mai_n1755_), .A1(mai_mai_n1753_), .B0(mai_mai_n1756_), .Y(mai_mai_n1757_));
  NO2        m1708(.A(mai_mai_n963_), .B(x3), .Y(mai_mai_n1758_));
  AOI210     m1709(.A0(mai_mai_n437_), .A1(mai_mai_n96_), .B0(mai_mai_n1758_), .Y(mai_mai_n1759_));
  NA3        m1710(.A(mai_mai_n561_), .B(mai_mai_n51_), .C(mai_mai_n56_), .Y(mai_mai_n1760_));
  INV        m1711(.A(x0), .Y(mai_mai_n1761_));
  OAI210     m1712(.A0(mai_mai_n1760_), .A1(mai_mai_n1759_), .B0(mai_mai_n1761_), .Y(mai_mai_n1762_));
  NO3        m1713(.A(mai_mai_n1762_), .B(mai_mai_n1757_), .C(mai_mai_n1752_), .Y(mai_mai_n1763_));
  AOI210     m1714(.A0(x8), .A1(x6), .B0(x5), .Y(mai_mai_n1764_));
  AO220      m1715(.A0(mai_mai_n1764_), .A1(mai_mai_n136_), .B0(mai_mai_n581_), .B1(mai_mai_n131_), .Y(mai_mai_n1765_));
  NA2        m1716(.A(mai_mai_n1765_), .B(mai_mai_n438_), .Y(mai_mai_n1766_));
  NO2        m1717(.A(mai_mai_n730_), .B(mai_mai_n136_), .Y(mai_mai_n1767_));
  NA3        m1718(.A(mai_mai_n1767_), .B(mai_mai_n1571_), .C(mai_mai_n125_), .Y(mai_mai_n1768_));
  NA3        m1719(.A(mai_mai_n363_), .B(mai_mai_n820_), .C(mai_mai_n241_), .Y(mai_mai_n1769_));
  NA3        m1720(.A(mai_mai_n1769_), .B(mai_mai_n1768_), .C(mai_mai_n1766_), .Y(mai_mai_n1770_));
  AOI210     m1721(.A0(mai_mai_n213_), .A1(x2), .B0(mai_mai_n484_), .Y(mai_mai_n1771_));
  NO2        m1722(.A(mai_mai_n1771_), .B(mai_mai_n105_), .Y(mai_mai_n1772_));
  NA3        m1723(.A(mai_mai_n778_), .B(mai_mai_n963_), .C(x7), .Y(mai_mai_n1773_));
  AOI210     m1724(.A0(mai_mai_n332_), .A1(mai_mai_n206_), .B0(mai_mai_n1773_), .Y(mai_mai_n1774_));
  OAI220     m1725(.A0(mai_mai_n860_), .A1(mai_mai_n292_), .B0(mai_mai_n629_), .B1(mai_mai_n666_), .Y(mai_mai_n1775_));
  NO3        m1726(.A(mai_mai_n1775_), .B(mai_mai_n1774_), .C(mai_mai_n1772_), .Y(mai_mai_n1776_));
  NA3        m1727(.A(mai_mai_n651_), .B(mai_mai_n182_), .C(mai_mai_n912_), .Y(mai_mai_n1777_));
  NA2        m1728(.A(mai_mai_n1777_), .B(mai_mai_n629_), .Y(mai_mai_n1778_));
  NA2        m1729(.A(mai_mai_n131_), .B(mai_mai_n123_), .Y(mai_mai_n1779_));
  OAI210     m1730(.A0(mai_mai_n1779_), .A1(mai_mai_n1356_), .B0(x0), .Y(mai_mai_n1780_));
  AOI210     m1731(.A0(mai_mai_n1778_), .A1(mai_mai_n1344_), .B0(mai_mai_n1780_), .Y(mai_mai_n1781_));
  OAI210     m1732(.A0(mai_mai_n1776_), .A1(mai_mai_n53_), .B0(mai_mai_n1781_), .Y(mai_mai_n1782_));
  AOI210     m1733(.A0(mai_mai_n1770_), .A1(x4), .B0(mai_mai_n1782_), .Y(mai_mai_n1783_));
  OA220      m1734(.A0(mai_mai_n1783_), .A1(mai_mai_n1763_), .B0(mai_mai_n1743_), .B1(mai_mai_n97_), .Y(mai27));
  NA2        m1735(.A(mai_mai_n877_), .B(mai_mai_n778_), .Y(mai_mai_n1785_));
  NA3        m1736(.A(mai_mai_n784_), .B(mai_mai_n352_), .C(mai_mai_n978_), .Y(mai_mai_n1786_));
  AOI210     m1737(.A0(mai_mai_n1786_), .A1(mai_mai_n1785_), .B0(mai_mai_n206_), .Y(mai_mai_n1787_));
  NA2        m1738(.A(mai_mai_n1787_), .B(mai_mai_n682_), .Y(mai_mai_n1788_));
  XO2        m1739(.A(x8), .B(x4), .Y(mai_mai_n1789_));
  NO3        m1740(.A(mai_mai_n1789_), .B(mai_mai_n437_), .C(mai_mai_n160_), .Y(mai_mai_n1790_));
  OA210      m1741(.A0(mai_mai_n1790_), .A1(mai_mai_n1194_), .B0(mai_mai_n265_), .Y(mai_mai_n1791_));
  NO2        m1742(.A(mai_mai_n385_), .B(mai_mai_n154_), .Y(mai_mai_n1792_));
  OAI210     m1743(.A0(mai_mai_n1792_), .A1(mai_mai_n1791_), .B0(mai_mai_n1067_), .Y(mai_mai_n1793_));
  NO2        m1744(.A(mai_mai_n1148_), .B(mai_mai_n197_), .Y(mai_mai_n1794_));
  NO2        m1745(.A(mai_mai_n679_), .B(mai_mai_n134_), .Y(mai_mai_n1795_));
  NO2        m1746(.A(mai_mai_n1132_), .B(mai_mai_n244_), .Y(mai_mai_n1796_));
  AOI220     m1747(.A0(mai_mai_n1796_), .A1(mai_mai_n1795_), .B0(mai_mai_n1794_), .B1(mai_mai_n527_), .Y(mai_mai_n1797_));
  NA3        m1748(.A(mai_mai_n1797_), .B(mai_mai_n1793_), .C(mai_mai_n1788_), .Y(mai28));
  NO3        m1749(.A(mai_mai_n1789_), .B(mai_mai_n1314_), .C(mai_mai_n138_), .Y(mai_mai_n1799_));
  OAI210     m1750(.A0(mai_mai_n1799_), .A1(mai_mai_n1210_), .B0(mai_mai_n573_), .Y(mai_mai_n1800_));
  NA3        m1751(.A(mai_mai_n1129_), .B(mai_mai_n854_), .C(x7), .Y(mai_mai_n1801_));
  NA2        m1752(.A(mai_mai_n1801_), .B(mai_mai_n1800_), .Y(mai_mai_n1802_));
  NA2        m1753(.A(mai_mai_n1188_), .B(mai_mai_n436_), .Y(mai_mai_n1803_));
  NA3        m1754(.A(mai_mai_n1803_), .B(mai_mai_n1333_), .C(mai_mai_n403_), .Y(mai_mai_n1804_));
  NO2        m1755(.A(mai_mai_n295_), .B(x4), .Y(mai_mai_n1805_));
  NA2        m1756(.A(mai_mai_n1805_), .B(mai_mai_n1758_), .Y(mai_mai_n1806_));
  NA2        m1757(.A(mai_mai_n1806_), .B(mai_mai_n1804_), .Y(mai_mai_n1807_));
  NO2        m1758(.A(mai_mai_n1188_), .B(mai_mai_n1166_), .Y(mai_mai_n1808_));
  NO4        m1759(.A(x6), .B(mai_mai_n56_), .C(x2), .D(x0), .Y(mai_mai_n1809_));
  OAI210     m1760(.A0(mai_mai_n1809_), .A1(mai_mai_n1808_), .B0(mai_mai_n1000_), .Y(mai_mai_n1810_));
  NA2        m1761(.A(mai_mai_n1123_), .B(mai_mai_n96_), .Y(mai_mai_n1811_));
  NA2        m1762(.A(mai_mai_n1030_), .B(mai_mai_n95_), .Y(mai_mai_n1812_));
  OAI210     m1763(.A0(mai_mai_n1812_), .A1(mai_mai_n1811_), .B0(mai_mai_n1810_), .Y(mai_mai_n1813_));
  OAI210     m1764(.A0(mai_mai_n1813_), .A1(mai_mai_n1807_), .B0(x7), .Y(mai_mai_n1814_));
  NO2        m1765(.A(mai_mai_n376_), .B(x7), .Y(mai_mai_n1815_));
  NO3        m1766(.A(mai_mai_n390_), .B(mai_mai_n259_), .C(mai_mai_n112_), .Y(mai_mai_n1816_));
  OAI210     m1767(.A0(mai_mai_n828_), .A1(mai_mai_n246_), .B0(mai_mai_n73_), .Y(mai_mai_n1817_));
  OAI220     m1768(.A0(mai_mai_n1817_), .A1(mai_mai_n1816_), .B0(mai_mai_n1815_), .B1(mai_mai_n99_), .Y(mai_mai_n1818_));
  INV        m1769(.A(mai_mai_n640_), .Y(mai_mai_n1819_));
  NO2        m1770(.A(mai_mai_n1736_), .B(mai_mai_n71_), .Y(mai_mai_n1820_));
  AOI220     m1771(.A0(mai_mai_n1820_), .A1(mai_mai_n1819_), .B0(mai_mai_n468_), .B1(mai_mai_n50_), .Y(mai_mai_n1821_));
  AOI210     m1772(.A0(mai_mai_n1821_), .A1(mai_mai_n1818_), .B0(mai_mai_n59_), .Y(mai_mai_n1822_));
  AOI220     m1773(.A0(mai_mai_n1319_), .A1(mai_mai_n655_), .B0(mai_mai_n402_), .B1(mai_mai_n446_), .Y(mai_mai_n1823_));
  OAI210     m1774(.A0(mai_mai_n1823_), .A1(mai_mai_n134_), .B0(x1), .Y(mai_mai_n1824_));
  NO2        m1775(.A(mai_mai_n1824_), .B(mai_mai_n1822_), .Y(mai_mai_n1825_));
  NO2        m1776(.A(mai_mai_n390_), .B(x5), .Y(mai_mai_n1826_));
  NOi21      m1777(.An(mai_mai_n687_), .B(mai_mai_n953_), .Y(mai_mai_n1827_));
  NO2        m1778(.A(mai_mai_n1289_), .B(mai_mai_n1577_), .Y(mai_mai_n1828_));
  NA2        m1779(.A(mai_mai_n1828_), .B(mai_mai_n1067_), .Y(mai_mai_n1829_));
  INV        m1780(.A(mai_mai_n972_), .Y(mai_mai_n1830_));
  AOI220     m1781(.A0(mai_mai_n1830_), .A1(mai_mai_n452_), .B0(mai_mai_n436_), .B1(mai_mai_n377_), .Y(mai_mai_n1831_));
  NO2        m1782(.A(mai_mai_n1831_), .B(mai_mai_n144_), .Y(mai_mai_n1832_));
  NA2        m1783(.A(mai_mai_n152_), .B(mai_mai_n67_), .Y(mai_mai_n1833_));
  OAI210     m1784(.A0(mai_mai_n1745_), .A1(mai_mai_n1833_), .B0(mai_mai_n53_), .Y(mai_mai_n1834_));
  OAI220     m1785(.A0(mai_mai_n667_), .A1(mai_mai_n249_), .B0(mai_mai_n663_), .B1(x6), .Y(mai_mai_n1835_));
  NO2        m1786(.A(mai_mai_n290_), .B(x4), .Y(mai_mai_n1836_));
  AOI220     m1787(.A0(mai_mai_n1836_), .A1(mai_mai_n352_), .B0(mai_mai_n1835_), .B1(x4), .Y(mai_mai_n1837_));
  NO3        m1788(.A(mai_mai_n1837_), .B(mai_mai_n311_), .C(x5), .Y(mai_mai_n1838_));
  NO2        m1789(.A(mai_mai_n687_), .B(mai_mai_n57_), .Y(mai_mai_n1839_));
  NA2        m1790(.A(mai_mai_n1795_), .B(mai_mai_n437_), .Y(mai_mai_n1840_));
  NA2        m1791(.A(mai_mai_n484_), .B(mai_mai_n224_), .Y(mai_mai_n1841_));
  AOI210     m1792(.A0(mai_mai_n1841_), .A1(mai_mai_n1840_), .B0(mai_mai_n244_), .Y(mai_mai_n1842_));
  NO4        m1793(.A(mai_mai_n1842_), .B(mai_mai_n1838_), .C(mai_mai_n1834_), .D(mai_mai_n1832_), .Y(mai_mai_n1843_));
  AOI220     m1794(.A0(mai_mai_n1843_), .A1(mai_mai_n1829_), .B0(mai_mai_n1825_), .B1(mai_mai_n1814_), .Y(mai_mai_n1844_));
  AOI210     m1795(.A0(mai_mai_n1802_), .A1(x3), .B0(mai_mai_n1844_), .Y(mai29));
  OAI210     m1796(.A0(mai_mai_n546_), .A1(mai_mai_n250_), .B0(mai_mai_n703_), .Y(mai_mai_n1846_));
  NA2        m1797(.A(mai_mai_n722_), .B(mai_mai_n1000_), .Y(mai_mai_n1847_));
  AO210      m1798(.A0(mai_mai_n1106_), .A1(mai_mai_n1115_), .B0(mai_mai_n1847_), .Y(mai_mai_n1848_));
  AOI210     m1799(.A0(mai_mai_n172_), .A1(mai_mai_n156_), .B0(mai_mai_n687_), .Y(mai_mai_n1849_));
  AOI210     m1800(.A0(mai_mai_n1348_), .A1(mai_mai_n72_), .B0(mai_mai_n1849_), .Y(mai_mai_n1850_));
  NA3        m1801(.A(mai_mai_n1850_), .B(mai_mai_n1848_), .C(mai_mai_n1846_), .Y(mai_mai_n1851_));
  NO3        m1802(.A(mai_mai_n649_), .B(mai_mai_n1089_), .C(mai_mai_n50_), .Y(mai_mai_n1852_));
  NO3        m1803(.A(mai_mai_n1852_), .B(mai_mai_n1187_), .C(mai_mai_n546_), .Y(mai_mai_n1853_));
  NO2        m1804(.A(mai_mai_n434_), .B(mai_mai_n58_), .Y(mai_mai_n1854_));
  AOI220     m1805(.A0(mai_mai_n1854_), .A1(mai_mai_n1149_), .B0(mai_mai_n652_), .B1(mai_mai_n1305_), .Y(mai_mai_n1855_));
  OAI210     m1806(.A0(mai_mai_n1853_), .A1(mai_mai_n532_), .B0(mai_mai_n1855_), .Y(mai_mai_n1856_));
  AOI210     m1807(.A0(mai_mai_n1851_), .A1(x6), .B0(mai_mai_n1856_), .Y(mai_mai_n1857_));
  OAI210     m1808(.A0(x8), .A1(x4), .B0(x5), .Y(mai_mai_n1858_));
  NA2        m1809(.A(mai_mai_n290_), .B(mai_mai_n138_), .Y(mai_mai_n1859_));
  NA4        m1810(.A(mai_mai_n1859_), .B(mai_mai_n2519_), .C(mai_mai_n648_), .D(mai_mai_n63_), .Y(mai_mai_n1860_));
  AOI210     m1811(.A0(mai_mai_n1255_), .A1(mai_mai_n259_), .B0(mai_mai_n1629_), .Y(mai_mai_n1861_));
  AOI210     m1812(.A0(mai_mai_n1861_), .A1(mai_mai_n1860_), .B0(mai_mai_n847_), .Y(mai_mai_n1862_));
  NA2        m1813(.A(mai_mai_n615_), .B(mai_mai_n283_), .Y(mai_mai_n1863_));
  NO2        m1814(.A(mai_mai_n1863_), .B(mai_mai_n1149_), .Y(mai_mai_n1864_));
  OAI210     m1815(.A0(mai_mai_n854_), .A1(x8), .B0(x7), .Y(mai_mai_n1865_));
  NO2        m1816(.A(mai_mai_n1865_), .B(mai_mai_n117_), .Y(mai_mai_n1866_));
  AN2        m1817(.A(mai_mai_n262_), .B(mai_mai_n1858_), .Y(mai_mai_n1867_));
  OAI220     m1818(.A0(mai_mai_n1867_), .A1(mai_mai_n575_), .B0(mai_mai_n1424_), .B1(mai_mai_n385_), .Y(mai_mai_n1868_));
  NO4        m1819(.A(mai_mai_n1868_), .B(mai_mai_n1866_), .C(mai_mai_n1864_), .D(mai_mai_n1862_), .Y(mai_mai_n1869_));
  OAI210     m1820(.A0(mai_mai_n1857_), .A1(x2), .B0(mai_mai_n1869_), .Y(mai_mai_n1870_));
  NA3        m1821(.A(x6), .B(mai_mai_n50_), .C(x2), .Y(mai_mai_n1871_));
  OAI210     m1822(.A0(mai_mai_n1166_), .A1(mai_mai_n342_), .B0(mai_mai_n1871_), .Y(mai_mai_n1872_));
  AOI210     m1823(.A0(mai_mai_n1872_), .A1(mai_mai_n332_), .B0(mai_mai_n1809_), .Y(mai_mai_n1873_));
  NO3        m1824(.A(mai_mai_n680_), .B(mai_mai_n353_), .C(mai_mai_n132_), .Y(mai_mai_n1874_));
  AOI210     m1825(.A0(mai_mai_n702_), .A1(mai_mai_n598_), .B0(mai_mai_n1874_), .Y(mai_mai_n1875_));
  OAI210     m1826(.A0(mai_mai_n1873_), .A1(x7), .B0(mai_mai_n1875_), .Y(mai_mai_n1876_));
  AOI210     m1827(.A0(mai_mai_n1040_), .A1(mai_mai_n390_), .B0(mai_mai_n1332_), .Y(mai_mai_n1877_));
  NO2        m1828(.A(mai_mai_n138_), .B(x2), .Y(mai_mai_n1878_));
  OA210      m1829(.A0(mai_mai_n1878_), .A1(mai_mai_n613_), .B0(mai_mai_n649_), .Y(mai_mai_n1879_));
  OAI210     m1830(.A0(mai_mai_n1879_), .A1(mai_mai_n1877_), .B0(mai_mai_n65_), .Y(mai_mai_n1880_));
  NO2        m1831(.A(mai_mai_n188_), .B(mai_mai_n77_), .Y(mai_mai_n1881_));
  OAI210     m1832(.A0(mai_mai_n1881_), .A1(mai_mai_n759_), .B0(mai_mai_n1049_), .Y(mai_mai_n1882_));
  NA3        m1833(.A(mai_mai_n1826_), .B(mai_mai_n217_), .C(mai_mai_n75_), .Y(mai_mai_n1883_));
  NA3        m1834(.A(mai_mai_n1883_), .B(mai_mai_n1882_), .C(mai_mai_n1880_), .Y(mai_mai_n1884_));
  AOI210     m1835(.A0(mai_mai_n1876_), .A1(x8), .B0(mai_mai_n1884_), .Y(mai_mai_n1885_));
  OAI210     m1836(.A0(mai_mai_n434_), .A1(mai_mai_n233_), .B0(mai_mai_n923_), .Y(mai_mai_n1886_));
  OAI210     m1837(.A0(mai_mai_n1886_), .A1(mai_mai_n1068_), .B0(mai_mai_n657_), .Y(mai_mai_n1887_));
  NO3        m1838(.A(mai_mai_n976_), .B(mai_mai_n343_), .C(mai_mai_n139_), .Y(mai_mai_n1888_));
  NA3        m1839(.A(mai_mai_n1888_), .B(mai_mai_n1236_), .C(mai_mai_n50_), .Y(mai_mai_n1889_));
  NO2        m1840(.A(mai_mai_n125_), .B(mai_mai_n85_), .Y(mai_mai_n1890_));
  AOI220     m1841(.A0(mai_mai_n1890_), .A1(mai_mai_n576_), .B0(mai_mai_n1808_), .B1(mai_mai_n349_), .Y(mai_mai_n1891_));
  NOi31      m1842(.An(mai_mai_n1069_), .B(mai_mai_n1764_), .C(mai_mai_n608_), .Y(mai_mai_n1892_));
  INV        m1843(.A(mai_mai_n1892_), .Y(mai_mai_n1893_));
  NA4        m1844(.A(mai_mai_n1893_), .B(mai_mai_n1891_), .C(mai_mai_n1889_), .D(mai_mai_n1887_), .Y(mai_mai_n1894_));
  NO4        m1845(.A(mai_mai_n1166_), .B(mai_mai_n160_), .C(mai_mai_n55_), .D(mai_mai_n67_), .Y(mai_mai_n1895_));
  NO4        m1846(.A(mai_mai_n1143_), .B(mai_mai_n492_), .C(mai_mai_n1305_), .D(mai_mai_n96_), .Y(mai_mai_n1896_));
  OAI210     m1847(.A0(mai_mai_n1896_), .A1(mai_mai_n1895_), .B0(mai_mai_n98_), .Y(mai_mai_n1897_));
  NO2        m1848(.A(x4), .B(mai_mai_n182_), .Y(mai_mai_n1898_));
  OAI210     m1849(.A0(mai_mai_n1898_), .A1(mai_mai_n1854_), .B0(mai_mai_n697_), .Y(mai_mai_n1899_));
  NA2        m1850(.A(mai_mai_n1809_), .B(mai_mai_n773_), .Y(mai_mai_n1900_));
  OR2        m1851(.A(mai_mai_n569_), .B(mai_mai_n1687_), .Y(mai_mai_n1901_));
  NA3        m1852(.A(mai_mai_n1901_), .B(mai_mai_n1899_), .C(mai_mai_n1897_), .Y(mai_mai_n1902_));
  AOI210     m1853(.A0(mai_mai_n1894_), .A1(mai_mai_n279_), .B0(mai_mai_n1902_), .Y(mai_mai_n1903_));
  OAI210     m1854(.A0(mai_mai_n1885_), .A1(x1), .B0(mai_mai_n1903_), .Y(mai_mai_n1904_));
  AO210      m1855(.A0(mai_mai_n1870_), .A1(x1), .B0(mai_mai_n1904_), .Y(mai30));
  NO3        m1856(.A(mai_mai_n1675_), .B(mai_mai_n566_), .C(mai_mai_n90_), .Y(mai_mai_n1906_));
  NO3        m1857(.A(mai_mai_n1087_), .B(mai_mai_n128_), .C(mai_mai_n373_), .Y(mai_mai_n1907_));
  INV        m1858(.A(mai_mai_n1907_), .Y(mai_mai_n1908_));
  AOI210     m1859(.A0(mai_mai_n1908_), .A1(mai_mai_n1906_), .B0(mai_mai_n56_), .Y(mai_mai_n1909_));
  NA2        m1860(.A(mai_mai_n778_), .B(mai_mai_n330_), .Y(mai_mai_n1910_));
  NA2        m1861(.A(mai_mai_n1910_), .B(mai_mai_n1290_), .Y(mai_mai_n1911_));
  OAI210     m1862(.A0(mai_mai_n1911_), .A1(mai_mai_n1909_), .B0(mai_mai_n98_), .Y(mai_mai_n1912_));
  OAI210     m1863(.A0(mai_mai_n953_), .A1(mai_mai_n561_), .B0(mai_mai_n657_), .Y(mai_mai_n1913_));
  AOI220     m1864(.A0(mai_mai_n438_), .A1(mai_mai_n901_), .B0(mai_mai_n316_), .B1(mai_mai_n446_), .Y(mai_mai_n1914_));
  AOI210     m1865(.A0(mai_mai_n1914_), .A1(mai_mai_n1913_), .B0(mai_mai_n244_), .Y(mai_mai_n1915_));
  NO2        m1866(.A(mai_mai_n113_), .B(x0), .Y(mai_mai_n1916_));
  AOI210     m1867(.A0(mai_mai_n494_), .A1(x6), .B0(mai_mai_n1916_), .Y(mai_mai_n1917_));
  NO2        m1868(.A(mai_mai_n1917_), .B(mai_mai_n54_), .Y(mai_mai_n1918_));
  AO210      m1869(.A0(mai_mai_n560_), .A1(mai_mai_n508_), .B0(x5), .Y(mai_mai_n1919_));
  NO2        m1870(.A(mai_mai_n694_), .B(mai_mai_n1919_), .Y(mai_mai_n1920_));
  AOI210     m1871(.A0(mai_mai_n1510_), .A1(mai_mai_n50_), .B0(mai_mai_n446_), .Y(mai_mai_n1921_));
  NA2        m1872(.A(mai_mai_n187_), .B(x2), .Y(mai_mai_n1922_));
  OA220      m1873(.A0(mai_mai_n1922_), .A1(mai_mai_n1921_), .B0(mai_mai_n263_), .B1(x6), .Y(mai_mai_n1923_));
  OAI210     m1874(.A0(x7), .A1(x6), .B0(x1), .Y(mai_mai_n1924_));
  NA3        m1875(.A(mai_mai_n57_), .B(x4), .C(mai_mai_n59_), .Y(mai_mai_n1925_));
  AOI220     m1876(.A0(mai_mai_n1925_), .A1(mai_mai_n1295_), .B0(mai_mai_n1924_), .B1(mai_mai_n1710_), .Y(mai_mai_n1926_));
  NO3        m1877(.A(mai_mai_n1293_), .B(mai_mai_n332_), .C(mai_mai_n978_), .Y(mai_mai_n1927_));
  NO2        m1878(.A(mai_mai_n506_), .B(mai_mai_n824_), .Y(mai_mai_n1928_));
  NOi21      m1879(.An(mai_mai_n1928_), .B(mai_mai_n809_), .Y(mai_mai_n1929_));
  NO3        m1880(.A(mai_mai_n1236_), .B(mai_mai_n219_), .C(mai_mai_n633_), .Y(mai_mai_n1930_));
  NO4        m1881(.A(mai_mai_n1930_), .B(mai_mai_n1929_), .C(mai_mai_n1927_), .D(mai_mai_n1926_), .Y(mai_mai_n1931_));
  OAI210     m1882(.A0(mai_mai_n1923_), .A1(mai_mai_n729_), .B0(mai_mai_n1931_), .Y(mai_mai_n1932_));
  NO4        m1883(.A(mai_mai_n1932_), .B(mai_mai_n1920_), .C(mai_mai_n1918_), .D(mai_mai_n1915_), .Y(mai_mai_n1933_));
  AOI210     m1884(.A0(mai_mai_n1933_), .A1(mai_mai_n1912_), .B0(x8), .Y(mai_mai_n1934_));
  NO3        m1885(.A(mai_mai_n482_), .B(mai_mai_n757_), .C(mai_mai_n53_), .Y(mai_mai_n1935_));
  NA2        m1886(.A(mai_mai_n1935_), .B(x6), .Y(mai_mai_n1936_));
  OAI210     m1887(.A0(mai_mai_n991_), .A1(mai_mai_n527_), .B0(mai_mai_n778_), .Y(mai_mai_n1937_));
  OAI210     m1888(.A0(mai_mai_n1639_), .A1(mai_mai_n319_), .B0(mai_mai_n116_), .Y(mai_mai_n1938_));
  AOI210     m1889(.A0(mai_mai_n368_), .A1(mai_mai_n216_), .B0(mai_mai_n68_), .Y(mai_mai_n1939_));
  AOI210     m1890(.A0(mai_mai_n953_), .A1(mai_mai_n720_), .B0(mai_mai_n1939_), .Y(mai_mai_n1940_));
  NA4        m1891(.A(mai_mai_n1940_), .B(mai_mai_n1938_), .C(mai_mai_n1937_), .D(mai_mai_n1936_), .Y(mai_mai_n1941_));
  NA2        m1892(.A(mai_mai_n1037_), .B(mai_mai_n59_), .Y(mai_mai_n1942_));
  AOI210     m1893(.A0(mai_mai_n882_), .A1(mai_mai_n483_), .B0(mai_mai_n662_), .Y(mai_mai_n1943_));
  OAI220     m1894(.A0(mai_mai_n1943_), .A1(mai_mai_n294_), .B0(mai_mai_n1942_), .B1(mai_mai_n473_), .Y(mai_mai_n1944_));
  AOI210     m1895(.A0(mai_mai_n1941_), .A1(x8), .B0(mai_mai_n1944_), .Y(mai_mai_n1945_));
  NO2        m1896(.A(mai_mai_n1945_), .B(mai_mai_n57_), .Y(mai_mai_n1946_));
  NA2        m1897(.A(mai_mai_n425_), .B(mai_mai_n809_), .Y(mai_mai_n1947_));
  NO2        m1898(.A(mai_mai_n881_), .B(mai_mai_n646_), .Y(mai_mai_n1948_));
  AOI210     m1899(.A0(mai_mai_n1948_), .A1(mai_mai_n1947_), .B0(mai_mai_n436_), .Y(mai_mai_n1949_));
  NO3        m1900(.A(mai_mai_n621_), .B(mai_mai_n399_), .C(mai_mai_n1087_), .Y(mai_mai_n1950_));
  NO3        m1901(.A(mai_mai_n1950_), .B(mai_mai_n1193_), .C(mai_mai_n1305_), .Y(mai_mai_n1951_));
  AOI210     m1902(.A0(mai_mai_n291_), .A1(x1), .B0(mai_mai_n139_), .Y(mai_mai_n1952_));
  NO2        m1903(.A(mai_mai_n297_), .B(x5), .Y(mai_mai_n1953_));
  NO2        m1904(.A(mai_mai_n1953_), .B(mai_mai_n817_), .Y(mai_mai_n1954_));
  OAI220     m1905(.A0(mai_mai_n1954_), .A1(mai_mai_n1011_), .B0(mai_mai_n1952_), .B1(mai_mai_n197_), .Y(mai_mai_n1955_));
  NO3        m1906(.A(mai_mai_n1955_), .B(mai_mai_n1951_), .C(mai_mai_n1949_), .Y(mai_mai_n1956_));
  NA2        m1907(.A(mai_mai_n921_), .B(mai_mai_n74_), .Y(mai_mai_n1957_));
  AO210      m1908(.A0(mai_mai_n1957_), .A1(mai_mai_n1511_), .B0(x3), .Y(mai_mai_n1958_));
  OAI220     m1909(.A0(mai_mai_n368_), .A1(mai_mai_n1193_), .B0(mai_mai_n343_), .B1(mai_mai_n219_), .Y(mai_mai_n1959_));
  AOI220     m1910(.A0(mai_mai_n1959_), .A1(x2), .B0(mai_mai_n59_), .B1(mai_mai_n1524_), .Y(mai_mai_n1960_));
  AOI210     m1911(.A0(mai_mai_n1960_), .A1(mai_mai_n1958_), .B0(mai_mai_n249_), .Y(mai_mai_n1961_));
  NO3        m1912(.A(mai_mai_n783_), .B(mai_mai_n681_), .C(mai_mai_n156_), .Y(mai_mai_n1962_));
  OAI210     m1913(.A0(mai_mai_n1962_), .A1(mai_mai_n2510_), .B0(mai_mai_n145_), .Y(mai_mai_n1963_));
  NA3        m1914(.A(x5), .B(x4), .C(mai_mai_n59_), .Y(mai_mai_n1964_));
  NO2        m1915(.A(mai_mai_n1244_), .B(mai_mai_n528_), .Y(mai_mai_n1965_));
  AOI210     m1916(.A0(mai_mai_n1260_), .A1(x2), .B0(mai_mai_n1965_), .Y(mai_mai_n1966_));
  AOI210     m1917(.A0(mai_mai_n1966_), .A1(mai_mai_n1963_), .B0(mai_mai_n50_), .Y(mai_mai_n1967_));
  NA3        m1918(.A(mai_mai_n1399_), .B(mai_mai_n1078_), .C(mai_mai_n466_), .Y(mai_mai_n1968_));
  AOI210     m1919(.A0(mai_mai_n1968_), .A1(mai_mai_n1957_), .B0(mai_mai_n594_), .Y(mai_mai_n1969_));
  AOI210     m1920(.A0(mai_mai_n978_), .A1(x1), .B0(mai_mai_n1255_), .Y(mai_mai_n1970_));
  OAI220     m1921(.A0(mai_mai_n295_), .A1(x4), .B0(mai_mai_n51_), .B1(x6), .Y(mai_mai_n1971_));
  NO2        m1922(.A(mai_mai_n111_), .B(mai_mai_n100_), .Y(mai_mai_n1972_));
  AOI220     m1923(.A0(mai_mai_n1972_), .A1(mai_mai_n1971_), .B0(mai_mai_n1108_), .B1(mai_mai_n608_), .Y(mai_mai_n1973_));
  OAI210     m1924(.A0(mai_mai_n1970_), .A1(mai_mai_n477_), .B0(mai_mai_n1973_), .Y(mai_mai_n1974_));
  NO4        m1925(.A(mai_mai_n1974_), .B(mai_mai_n1969_), .C(mai_mai_n1967_), .D(mai_mai_n1961_), .Y(mai_mai_n1975_));
  OAI210     m1926(.A0(mai_mai_n1956_), .A1(mai_mai_n125_), .B0(mai_mai_n1975_), .Y(mai_mai_n1976_));
  NO3        m1927(.A(mai_mai_n1976_), .B(mai_mai_n1946_), .C(mai_mai_n1934_), .Y(mai31));
  NA2        m1928(.A(mai_mai_n940_), .B(mai_mai_n344_), .Y(mai_mai_n1978_));
  NO2        m1929(.A(mai_mai_n439_), .B(mai_mai_n657_), .Y(mai_mai_n1979_));
  AOI210     m1930(.A0(mai_mai_n1979_), .A1(mai_mai_n1978_), .B0(mai_mai_n58_), .Y(mai_mai_n1980_));
  NO2        m1931(.A(mai_mai_n758_), .B(mai_mai_n56_), .Y(mai_mai_n1981_));
  AOI220     m1932(.A0(mai_mai_n1981_), .A1(x2), .B0(mai_mai_n83_), .B1(x0), .Y(mai_mai_n1982_));
  NA3        m1933(.A(mai_mai_n1982_), .B(mai_mai_n1900_), .C(mai_mai_n1744_), .Y(mai_mai_n1983_));
  OAI210     m1934(.A0(mai_mai_n1983_), .A1(mai_mai_n1980_), .B0(mai_mai_n53_), .Y(mai_mai_n1984_));
  NO2        m1935(.A(mai_mai_n422_), .B(mai_mai_n657_), .Y(mai_mai_n1985_));
  NO3        m1936(.A(mai_mai_n1836_), .B(mai_mai_n1809_), .C(mai_mai_n848_), .Y(mai_mai_n1986_));
  OA220      m1937(.A0(mai_mai_n1986_), .A1(mai_mai_n466_), .B0(mai_mai_n1985_), .B1(mai_mai_n1392_), .Y(mai_mai_n1987_));
  AOI210     m1938(.A0(mai_mai_n1987_), .A1(mai_mai_n1984_), .B0(mai_mai_n96_), .Y(mai_mai_n1988_));
  NO4        m1939(.A(mai_mai_n1104_), .B(mai_mai_n353_), .C(mai_mai_n1510_), .D(mai_mai_n64_), .Y(mai_mai_n1989_));
  AOI210     m1940(.A0(mai_mai_n1548_), .A1(mai_mai_n1282_), .B0(mai_mai_n434_), .Y(mai_mai_n1990_));
  OAI220     m1941(.A0(mai_mai_n1245_), .A1(mai_mai_n913_), .B0(mai_mai_n747_), .B1(mai_mai_n105_), .Y(mai_mai_n1991_));
  NO3        m1942(.A(mai_mai_n1991_), .B(mai_mai_n1990_), .C(mai_mai_n1989_), .Y(mai_mai_n1992_));
  NO2        m1943(.A(mai_mai_n1992_), .B(x5), .Y(mai_mai_n1993_));
  AOI220     m1944(.A0(mai_mai_n437_), .A1(mai_mai_n608_), .B0(mai_mai_n561_), .B1(mai_mai_n62_), .Y(mai_mai_n1994_));
  AOI210     m1945(.A0(mai_mai_n1994_), .A1(mai_mai_n569_), .B0(mai_mai_n1166_), .Y(mai_mai_n1995_));
  AOI220     m1946(.A0(mai_mai_n922_), .A1(mai_mai_n707_), .B0(mai_mai_n1087_), .B1(mai_mai_n110_), .Y(mai_mai_n1996_));
  NO2        m1947(.A(mai_mai_n1996_), .B(mai_mai_n376_), .Y(mai_mai_n1997_));
  NO4        m1948(.A(mai_mai_n1997_), .B(mai_mai_n1995_), .C(mai_mai_n1993_), .D(mai_mai_n1988_), .Y(mai_mai_n1998_));
  NA2        m1949(.A(mai_mai_n483_), .B(mai_mai_n59_), .Y(mai_mai_n1999_));
  AOI210     m1950(.A0(mai_mai_n532_), .A1(mai_mai_n1999_), .B0(mai_mai_n131_), .Y(mai_mai_n2000_));
  OAI210     m1951(.A0(mai_mai_n94_), .A1(mai_mai_n262_), .B0(mai_mai_n1942_), .Y(mai_mai_n2001_));
  OAI210     m1952(.A0(mai_mai_n2001_), .A1(mai_mai_n2000_), .B0(x7), .Y(mai_mai_n2002_));
  NO3        m1953(.A(mai_mai_n368_), .B(mai_mai_n55_), .C(x7), .Y(mai_mai_n2003_));
  OA210      m1954(.A0(mai_mai_n2003_), .A1(mai_mai_n1254_), .B0(mai_mai_n92_), .Y(mai_mai_n2004_));
  NA2        m1955(.A(mai_mai_n1034_), .B(mai_mai_n84_), .Y(mai_mai_n2005_));
  AOI210     m1956(.A0(mai_mai_n860_), .A1(mai_mai_n100_), .B0(mai_mai_n2005_), .Y(mai_mai_n2006_));
  NA2        m1957(.A(mai_mai_n1466_), .B(x6), .Y(mai_mai_n2007_));
  AOI210     m1958(.A0(mai_mai_n2007_), .A1(mai_mai_n278_), .B0(mai_mai_n96_), .Y(mai_mai_n2008_));
  NA2        m1959(.A(mai_mai_n1129_), .B(mai_mai_n307_), .Y(mai_mai_n2009_));
  AOI210     m1960(.A0(mai_mai_n2009_), .A1(mai_mai_n629_), .B0(mai_mai_n53_), .Y(mai_mai_n2010_));
  NO4        m1961(.A(mai_mai_n2010_), .B(mai_mai_n2008_), .C(mai_mai_n2006_), .D(mai_mai_n2004_), .Y(mai_mai_n2011_));
  AOI210     m1962(.A0(mai_mai_n2011_), .A1(mai_mai_n2002_), .B0(mai_mai_n666_), .Y(mai_mai_n2012_));
  OAI220     m1963(.A0(mai_mai_n1665_), .A1(mai_mai_n1811_), .B0(mai_mai_n883_), .B1(mai_mai_n1999_), .Y(mai_mai_n2013_));
  NA2        m1964(.A(mai_mai_n2013_), .B(x3), .Y(mai_mai_n2014_));
  AOI220     m1965(.A0(mai_mai_n1314_), .A1(x8), .B0(mai_mai_n60_), .B1(x1), .Y(mai_mai_n2015_));
  NO3        m1966(.A(mai_mai_n2015_), .B(mai_mai_n1060_), .C(x6), .Y(mai_mai_n2016_));
  AOI220     m1967(.A0(mai_mai_n598_), .A1(mai_mai_n399_), .B0(mai_mai_n483_), .B1(mai_mai_n72_), .Y(mai_mai_n2017_));
  NA2        m1968(.A(mai_mai_n106_), .B(mai_mai_n519_), .Y(mai_mai_n2018_));
  OAI220     m1969(.A0(mai_mai_n2018_), .A1(mai_mai_n1811_), .B0(mai_mai_n2017_), .B1(x4), .Y(mai_mai_n2019_));
  NO2        m1970(.A(mai_mai_n2019_), .B(mai_mai_n2016_), .Y(mai_mai_n2020_));
  AOI210     m1971(.A0(mai_mai_n2020_), .A1(mai_mai_n2014_), .B0(mai_mai_n175_), .Y(mai_mai_n2021_));
  NO3        m1972(.A(mai_mai_n599_), .B(mai_mai_n576_), .C(mai_mai_n681_), .Y(mai_mai_n2022_));
  OAI210     m1973(.A0(mai_mai_n2022_), .A1(mai_mai_n1027_), .B0(x3), .Y(mai_mai_n2023_));
  NO4        m1974(.A(mai_mai_n771_), .B(mai_mai_n1166_), .C(mai_mai_n745_), .D(x5), .Y(mai_mai_n2024_));
  NO3        m1975(.A(x6), .B(mai_mai_n56_), .C(x1), .Y(mai_mai_n2025_));
  NA2        m1976(.A(mai_mai_n2025_), .B(mai_mai_n274_), .Y(mai_mai_n2026_));
  INV        m1977(.A(mai_mai_n2026_), .Y(mai_mai_n2027_));
  NO2        m1978(.A(mai_mai_n818_), .B(mai_mai_n237_), .Y(mai_mai_n2028_));
  NO3        m1979(.A(mai_mai_n2028_), .B(mai_mai_n2027_), .C(mai_mai_n2024_), .Y(mai_mai_n2029_));
  AOI210     m1980(.A0(mai_mai_n2029_), .A1(mai_mai_n2023_), .B0(mai_mai_n523_), .Y(mai_mai_n2030_));
  OAI210     m1981(.A0(mai_mai_n598_), .A1(mai_mai_n460_), .B0(mai_mai_n901_), .Y(mai_mai_n2031_));
  NO3        m1982(.A(mai_mai_n452_), .B(mai_mai_n338_), .C(mai_mai_n50_), .Y(mai_mai_n2032_));
  NA2        m1983(.A(mai_mai_n2032_), .B(mai_mai_n1105_), .Y(mai_mai_n2033_));
  AOI210     m1984(.A0(mai_mai_n2033_), .A1(mai_mai_n2031_), .B0(mai_mai_n383_), .Y(mai_mai_n2034_));
  NO2        m1985(.A(mai_mai_n206_), .B(mai_mai_n528_), .Y(mai_mai_n2035_));
  OAI210     m1986(.A0(mai_mai_n128_), .A1(x2), .B0(mai_mai_n2035_), .Y(mai_mai_n2036_));
  NA3        m1987(.A(mai_mai_n399_), .B(mai_mai_n317_), .C(mai_mai_n71_), .Y(mai_mai_n2037_));
  OA210      m1988(.A0(mai_mai_n232_), .A1(mai_mai_n215_), .B0(mai_mai_n2037_), .Y(mai_mai_n2038_));
  AOI210     m1989(.A0(mai_mai_n2038_), .A1(mai_mai_n2036_), .B0(mai_mai_n63_), .Y(mai_mai_n2039_));
  NA2        m1990(.A(mai_mai_n111_), .B(mai_mai_n57_), .Y(mai_mai_n2040_));
  AOI220     m1991(.A0(mai_mai_n1494_), .A1(mai_mai_n867_), .B0(mai_mai_n261_), .B1(x4), .Y(mai_mai_n2041_));
  AOI220     m1992(.A0(mai_mai_n1541_), .A1(mai_mai_n600_), .B0(mai_mai_n695_), .B1(mai_mai_n745_), .Y(mai_mai_n2042_));
  OAI220     m1993(.A0(mai_mai_n2042_), .A1(mai_mai_n2040_), .B0(mai_mai_n2041_), .B1(mai_mai_n180_), .Y(mai_mai_n2043_));
  OR3        m1994(.A(mai_mai_n2043_), .B(mai_mai_n2039_), .C(mai_mai_n2034_), .Y(mai_mai_n2044_));
  NO4        m1995(.A(mai_mai_n2044_), .B(mai_mai_n2030_), .C(mai_mai_n2021_), .D(mai_mai_n2012_), .Y(mai_mai_n2045_));
  OAI210     m1996(.A0(mai_mai_n1998_), .A1(x3), .B0(mai_mai_n2045_), .Y(mai32));
  NA2        m1997(.A(mai_mai_n759_), .B(mai_mai_n56_), .Y(mai_mai_n2047_));
  OAI210     m1998(.A0(mai_mai_n1608_), .A1(mai_mai_n1375_), .B0(mai_mai_n1401_), .Y(mai_mai_n2048_));
  AOI210     m1999(.A0(mai_mai_n1981_), .A1(mai_mai_n265_), .B0(mai_mai_n2048_), .Y(mai_mai_n2049_));
  AOI210     m2000(.A0(mai_mai_n2049_), .A1(mai_mai_n2047_), .B0(mai_mai_n50_), .Y(mai_mai_n2050_));
  NA3        m2001(.A(mai_mai_n57_), .B(mai_mai_n769_), .C(mai_mai_n277_), .Y(mai_mai_n2051_));
  NA2        m2002(.A(mai_mai_n718_), .B(mai_mai_n536_), .Y(mai_mai_n2052_));
  NO3        m2003(.A(mai_mai_n364_), .B(mai_mai_n564_), .C(mai_mai_n773_), .Y(mai_mai_n2053_));
  NO3        m2004(.A(mai_mai_n1293_), .B(mai_mai_n572_), .C(mai_mai_n259_), .Y(mai_mai_n2054_));
  NO3        m2005(.A(mai_mai_n2054_), .B(mai_mai_n2053_), .C(mai_mai_n2052_), .Y(mai_mai_n2055_));
  AOI210     m2006(.A0(mai_mai_n2055_), .A1(mai_mai_n2051_), .B0(mai_mai_n132_), .Y(mai_mai_n2056_));
  OAI220     m2007(.A0(mai_mai_n392_), .A1(x7), .B0(mai_mai_n290_), .B1(mai_mai_n283_), .Y(mai_mai_n2057_));
  NA2        m2008(.A(mai_mai_n2057_), .B(mai_mai_n921_), .Y(mai_mai_n2058_));
  INV        m2009(.A(mai_mai_n824_), .Y(mai_mai_n2059_));
  AOI220     m2010(.A0(mai_mai_n2059_), .A1(mai_mai_n1767_), .B0(mai_mai_n520_), .B1(mai_mai_n121_), .Y(mai_mai_n2060_));
  AOI210     m2011(.A0(mai_mai_n2060_), .A1(mai_mai_n2058_), .B0(mai_mai_n98_), .Y(mai_mai_n2061_));
  NA3        m2012(.A(mai_mai_n1254_), .B(mai_mai_n1089_), .C(mai_mai_n105_), .Y(mai_mai_n2062_));
  NA2        m2013(.A(mai_mai_n1180_), .B(mai_mai_n998_), .Y(mai_mai_n2063_));
  AOI210     m2014(.A0(mai_mai_n2063_), .A1(mai_mai_n2062_), .B0(mai_mai_n56_), .Y(mai_mai_n2064_));
  NA2        m2015(.A(mai_mai_n921_), .B(mai_mai_n57_), .Y(mai_mai_n2065_));
  NOi21      m2016(.An(mai_mai_n2065_), .B(mai_mai_n121_), .Y(mai_mai_n2066_));
  NA2        m2017(.A(mai_mai_n968_), .B(mai_mai_n237_), .Y(mai_mai_n2067_));
  NO3        m2018(.A(mai_mai_n2067_), .B(mai_mai_n2066_), .C(mai_mai_n59_), .Y(mai_mai_n2068_));
  OR4        m2019(.A(mai_mai_n2068_), .B(mai_mai_n2064_), .C(mai_mai_n2061_), .D(mai_mai_n2056_), .Y(mai_mai_n2069_));
  OAI210     m2020(.A0(mai_mai_n2069_), .A1(mai_mai_n2050_), .B0(mai_mai_n96_), .Y(mai_mai_n2070_));
  NO3        m2021(.A(mai_mai_n1166_), .B(mai_mai_n136_), .C(mai_mai_n114_), .Y(mai_mai_n2071_));
  NO2        m2022(.A(mai_mai_n371_), .B(mai_mai_n55_), .Y(mai_mai_n2072_));
  NA2        m2023(.A(mai_mai_n2072_), .B(mai_mai_n104_), .Y(mai_mai_n2073_));
  INV        m2024(.A(mai_mai_n2073_), .Y(mai_mai_n2074_));
  OAI210     m2025(.A0(mai_mai_n2074_), .A1(mai_mai_n2071_), .B0(x3), .Y(mai_mai_n2075_));
  OAI210     m2026(.A0(mai_mai_n854_), .A1(mai_mai_n259_), .B0(mai_mai_n50_), .Y(mai_mai_n2076_));
  NO2        m2027(.A(mai_mai_n98_), .B(mai_mai_n2076_), .Y(mai_mai_n2077_));
  OAI210     m2028(.A0(mai_mai_n2077_), .A1(mai_mai_n1748_), .B0(mai_mai_n681_), .Y(mai_mai_n2078_));
  NO3        m2029(.A(mai_mai_n769_), .B(mai_mai_n351_), .C(mai_mai_n132_), .Y(mai_mai_n2079_));
  NA2        m2030(.A(mai_mai_n2079_), .B(mai_mai_n59_), .Y(mai_mai_n2080_));
  NA2        m2031(.A(mai_mai_n1093_), .B(mai_mai_n67_), .Y(mai_mai_n2081_));
  NO2        m2032(.A(mai_mai_n1815_), .B(mai_mai_n578_), .Y(mai_mai_n2082_));
  AOI210     m2033(.A0(mai_mai_n2082_), .A1(mai_mai_n1749_), .B0(mai_mai_n2081_), .Y(mai_mai_n2083_));
  NO2        m2034(.A(mai_mai_n262_), .B(mai_mai_n57_), .Y(mai_mai_n2084_));
  NO2        m2035(.A(mai_mai_n2084_), .B(mai_mai_n960_), .Y(mai_mai_n2085_));
  NOi31      m2036(.An(mai_mai_n697_), .B(mai_mai_n2085_), .C(mai_mai_n268_), .Y(mai_mai_n2086_));
  NO3        m2037(.A(mai_mai_n1247_), .B(mai_mai_n206_), .C(mai_mai_n244_), .Y(mai_mai_n2087_));
  NO4        m2038(.A(mai_mai_n2087_), .B(mai_mai_n2086_), .C(mai_mai_n2083_), .D(x1), .Y(mai_mai_n2088_));
  NA4        m2039(.A(mai_mai_n2088_), .B(mai_mai_n2080_), .C(mai_mai_n2078_), .D(mai_mai_n2075_), .Y(mai_mai_n2089_));
  AO210      m2040(.A0(mai_mai_n1040_), .A1(mai_mai_n387_), .B0(mai_mai_n963_), .Y(mai_mai_n2090_));
  NA3        m2041(.A(mai_mai_n1789_), .B(mai_mai_n545_), .C(mai_mai_n262_), .Y(mai_mai_n2091_));
  AOI210     m2042(.A0(mai_mai_n2091_), .A1(mai_mai_n2090_), .B0(mai_mai_n292_), .Y(mai_mai_n2092_));
  NA4        m2043(.A(mai_mai_n1202_), .B(mai_mai_n517_), .C(mai_mai_n376_), .D(mai_mai_n217_), .Y(mai_mai_n2093_));
  NO3        m2044(.A(mai_mai_n1359_), .B(mai_mai_n963_), .C(x2), .Y(mai_mai_n2094_));
  NO2        m2045(.A(mai_mai_n1188_), .B(mai_mai_n374_), .Y(mai_mai_n2095_));
  NO2        m2046(.A(mai_mai_n1727_), .B(mai_mai_n63_), .Y(mai_mai_n2096_));
  NO4        m2047(.A(mai_mai_n2096_), .B(mai_mai_n2095_), .C(mai_mai_n2094_), .D(mai_mai_n53_), .Y(mai_mai_n2097_));
  NO3        m2048(.A(mai_mai_n456_), .B(mai_mai_n1034_), .C(mai_mai_n111_), .Y(mai_mai_n2098_));
  OAI220     m2049(.A0(mai_mai_n666_), .A1(mai_mai_n162_), .B0(mai_mai_n343_), .B1(mai_mai_n132_), .Y(mai_mai_n2099_));
  OAI210     m2050(.A0(mai_mai_n2099_), .A1(mai_mai_n2098_), .B0(mai_mai_n65_), .Y(mai_mai_n2100_));
  NO2        m2051(.A(mai_mai_n1858_), .B(mai_mai_n355_), .Y(mai_mai_n2101_));
  NA2        m2052(.A(mai_mai_n1754_), .B(mai_mai_n2101_), .Y(mai_mai_n2102_));
  NA4        m2053(.A(mai_mai_n2102_), .B(mai_mai_n2100_), .C(mai_mai_n2097_), .D(mai_mai_n2093_), .Y(mai_mai_n2103_));
  OAI210     m2054(.A0(mai_mai_n2103_), .A1(mai_mai_n2092_), .B0(mai_mai_n2089_), .Y(mai_mai_n2104_));
  NO3        m2055(.A(mai_mai_n1155_), .B(mai_mai_n95_), .C(mai_mai_n67_), .Y(mai_mai_n2105_));
  NO2        m2056(.A(mai_mai_n554_), .B(mai_mai_n359_), .Y(mai_mai_n2106_));
  OAI210     m2057(.A0(mai_mai_n2105_), .A1(mai_mai_n1338_), .B0(mai_mai_n2106_), .Y(mai_mai_n2107_));
  NO3        m2058(.A(x8), .B(mai_mai_n67_), .C(x2), .Y(mai_mai_n2108_));
  OAI220     m2059(.A0(mai_mai_n2108_), .A1(mai_mai_n608_), .B0(mai_mai_n1348_), .B1(mai_mai_n83_), .Y(mai_mai_n2109_));
  AOI220     m2060(.A0(mai_mai_n546_), .A1(mai_mai_n778_), .B0(mai_mai_n657_), .B1(mai_mai_n242_), .Y(mai_mai_n2110_));
  AOI210     m2061(.A0(mai_mai_n2110_), .A1(mai_mai_n2109_), .B0(mai_mai_n252_), .Y(mai_mai_n2111_));
  NA2        m2062(.A(mai_mai_n968_), .B(mai_mai_n1087_), .Y(mai_mai_n2112_));
  NO2        m2063(.A(mai_mai_n653_), .B(mai_mai_n2112_), .Y(mai_mai_n2113_));
  AOI210     m2064(.A0(mai_mai_n576_), .A1(mai_mai_n608_), .B0(mai_mai_n672_), .Y(mai_mai_n2114_));
  NO2        m2065(.A(mai_mai_n2114_), .B(mai_mai_n1710_), .Y(mai_mai_n2115_));
  NO2        m2066(.A(mai_mai_n440_), .B(mai_mai_n422_), .Y(mai_mai_n2116_));
  NOi31      m2067(.An(mai_mai_n1416_), .B(mai_mai_n2116_), .C(mai_mai_n576_), .Y(mai_mai_n2117_));
  NO4        m2068(.A(mai_mai_n2117_), .B(mai_mai_n2115_), .C(mai_mai_n2113_), .D(mai_mai_n2111_), .Y(mai_mai_n2118_));
  NA4        m2069(.A(mai_mai_n2118_), .B(mai_mai_n2107_), .C(mai_mai_n2104_), .D(mai_mai_n2070_), .Y(mai33));
  OAI210     m2070(.A0(mai_mai_n774_), .A1(x1), .B0(mai_mai_n191_), .Y(mai_mai_n2120_));
  OAI210     m2071(.A0(mai_mai_n1953_), .A1(mai_mai_n167_), .B0(mai_mai_n317_), .Y(mai_mai_n2121_));
  NA2        m2072(.A(mai_mai_n1023_), .B(mai_mai_n342_), .Y(mai_mai_n2122_));
  NA3        m2073(.A(mai_mai_n2122_), .B(mai_mai_n2121_), .C(mai_mai_n620_), .Y(mai_mai_n2123_));
  AOI210     m2074(.A0(mai_mai_n2120_), .A1(x5), .B0(mai_mai_n2123_), .Y(mai_mai_n2124_));
  NA2        m2075(.A(mai_mai_n216_), .B(mai_mai_n70_), .Y(mai_mai_n2125_));
  NA4        m2076(.A(mai_mai_n1645_), .B(mai_mai_n555_), .C(mai_mai_n233_), .D(x4), .Y(mai_mai_n2126_));
  AOI210     m2077(.A0(mai_mai_n2126_), .A1(mai_mai_n2125_), .B0(mai_mai_n342_), .Y(mai_mai_n2127_));
  OAI210     m2078(.A0(mai_mai_n425_), .A1(mai_mai_n256_), .B0(mai_mai_n53_), .Y(mai_mai_n2128_));
  NO2        m2079(.A(mai_mai_n2128_), .B(mai_mai_n63_), .Y(mai_mai_n2129_));
  NA2        m2080(.A(mai_mai_n1561_), .B(mai_mai_n67_), .Y(mai_mai_n2130_));
  NO3        m2081(.A(mai_mai_n2130_), .B(mai_mai_n2129_), .C(mai_mai_n2127_), .Y(mai_mai_n2131_));
  OAI210     m2082(.A0(mai_mai_n2124_), .A1(x4), .B0(mai_mai_n2131_), .Y(mai_mai_n2132_));
  OAI210     m2083(.A0(mai_mai_n134_), .A1(x5), .B0(mai_mai_n226_), .Y(mai_mai_n2133_));
  NO2        m2084(.A(mai_mai_n921_), .B(mai_mai_n214_), .Y(mai_mai_n2134_));
  NA2        m2085(.A(mai_mai_n623_), .B(x7), .Y(mai_mai_n2135_));
  NO2        m2086(.A(mai_mai_n2135_), .B(mai_mai_n2134_), .Y(mai_mai_n2136_));
  AOI210     m2087(.A0(mai_mai_n2133_), .A1(mai_mai_n976_), .B0(mai_mai_n2136_), .Y(mai_mai_n2137_));
  NO2        m2088(.A(mai_mai_n2065_), .B(mai_mai_n204_), .Y(mai_mai_n2138_));
  NO2        m2089(.A(mai_mai_n1549_), .B(mai_mai_n913_), .Y(mai_mai_n2139_));
  OAI210     m2090(.A0(mai_mai_n824_), .A1(mai_mai_n51_), .B0(x6), .Y(mai_mai_n2140_));
  NO2        m2091(.A(mai_mai_n602_), .B(mai_mai_n494_), .Y(mai_mai_n2141_));
  NO4        m2092(.A(mai_mai_n2141_), .B(mai_mai_n2140_), .C(mai_mai_n2139_), .D(mai_mai_n2138_), .Y(mai_mai_n2142_));
  OAI210     m2093(.A0(mai_mai_n2137_), .A1(mai_mai_n50_), .B0(mai_mai_n2142_), .Y(mai_mai_n2143_));
  NA3        m2094(.A(mai_mai_n2143_), .B(mai_mai_n2132_), .C(mai_mai_n59_), .Y(mai_mai_n2144_));
  NA2        m2095(.A(mai_mai_n524_), .B(mai_mai_n97_), .Y(mai_mai_n2145_));
  NO3        m2096(.A(mai_mai_n1476_), .B(mai_mai_n363_), .C(x4), .Y(mai_mai_n2146_));
  AOI210     m2097(.A0(mai_mai_n2146_), .A1(mai_mai_n2145_), .B0(mai_mai_n428_), .Y(mai_mai_n2147_));
  NA2        m2098(.A(mai_mai_n776_), .B(mai_mai_n96_), .Y(mai_mai_n2148_));
  INV        m2099(.A(mai_mai_n2148_), .Y(mai_mai_n2149_));
  NO2        m2100(.A(mai_mai_n687_), .B(mai_mai_n364_), .Y(mai_mai_n2150_));
  NA2        m2101(.A(mai_mai_n490_), .B(mai_mai_n53_), .Y(mai_mai_n2151_));
  AOI210     m2102(.A0(mai_mai_n2150_), .A1(mai_mai_n2149_), .B0(mai_mai_n2151_), .Y(mai_mai_n2152_));
  OAI210     m2103(.A0(mai_mai_n2147_), .A1(mai_mai_n59_), .B0(mai_mai_n2152_), .Y(mai_mai_n2153_));
  AOI220     m2104(.A0(mai_mai_n666_), .A1(mai_mai_n223_), .B0(mai_mai_n376_), .B1(mai_mai_n217_), .Y(mai_mai_n2154_));
  NA2        m2105(.A(mai_mai_n704_), .B(mai_mai_n930_), .Y(mai_mai_n2155_));
  OAI210     m2106(.A0(mai_mai_n2155_), .A1(mai_mai_n2154_), .B0(mai_mai_n291_), .Y(mai_mai_n2156_));
  AOI210     m2107(.A0(mai_mai_n1981_), .A1(mai_mai_n205_), .B0(mai_mai_n53_), .Y(mai_mai_n2157_));
  NO2        m2108(.A(mai_mai_n132_), .B(mai_mai_n327_), .Y(mai_mai_n2158_));
  AOI220     m2109(.A0(mai_mai_n2158_), .A1(mai_mai_n947_), .B0(mai_mai_n652_), .B1(mai_mai_n342_), .Y(mai_mai_n2159_));
  NA2        m2110(.A(mai_mai_n436_), .B(mai_mai_n488_), .Y(mai_mai_n2160_));
  NO3        m2111(.A(mai_mai_n2160_), .B(mai_mai_n982_), .C(mai_mai_n172_), .Y(mai_mai_n2161_));
  AOI210     m2112(.A0(mai_mai_n1688_), .A1(mai_mai_n1129_), .B0(mai_mai_n2161_), .Y(mai_mai_n2162_));
  NA4        m2113(.A(mai_mai_n2162_), .B(mai_mai_n2159_), .C(mai_mai_n2157_), .D(mai_mai_n2156_), .Y(mai_mai_n2163_));
  NA3        m2114(.A(mai_mai_n2163_), .B(mai_mai_n2153_), .C(mai_mai_n57_), .Y(mai_mai_n2164_));
  NAi21      m2115(.An(mai_mai_n1131_), .B(mai_mai_n479_), .Y(mai_mai_n2165_));
  NA4        m2116(.A(mai_mai_n623_), .B(mai_mai_n1236_), .C(mai_mai_n460_), .D(mai_mai_n50_), .Y(mai_mai_n2166_));
  OAI210     m2117(.A0(mai_mai_n2158_), .A1(mai_mai_n1928_), .B0(x2), .Y(mai_mai_n2167_));
  NA4        m2118(.A(mai_mai_n274_), .B(mai_mai_n146_), .C(mai_mai_n263_), .D(mai_mai_n111_), .Y(mai_mai_n2168_));
  NA3        m2119(.A(mai_mai_n2168_), .B(mai_mai_n2167_), .C(mai_mai_n2166_), .Y(mai_mai_n2169_));
  AO220      m2120(.A0(mai_mai_n2169_), .A1(x0), .B0(mai_mai_n2165_), .B1(mai_mai_n129_), .Y(mai_mai_n2170_));
  NA3        m2121(.A(mai_mai_n745_), .B(mai_mai_n342_), .C(mai_mai_n60_), .Y(mai_mai_n2171_));
  NA2        m2122(.A(mai_mai_n621_), .B(mai_mai_n506_), .Y(mai_mai_n2172_));
  OAI220     m2123(.A0(mai_mai_n2172_), .A1(mai_mai_n50_), .B0(mai_mai_n2171_), .B1(mai_mai_n67_), .Y(mai_mai_n2173_));
  OAI210     m2124(.A0(mai_mai_n1445_), .A1(mai_mai_n338_), .B0(mai_mai_n99_), .Y(mai_mai_n2174_));
  OAI210     m2125(.A0(mai_mai_n2511_), .A1(mai_mai_n376_), .B0(mai_mai_n2174_), .Y(mai_mai_n2175_));
  OAI210     m2126(.A0(mai_mai_n2175_), .A1(mai_mai_n2173_), .B0(mai_mai_n93_), .Y(mai_mai_n2176_));
  NA2        m2127(.A(mai_mai_n122_), .B(mai_mai_n371_), .Y(mai_mai_n2177_));
  NA2        m2128(.A(mai_mai_n2177_), .B(mai_mai_n1714_), .Y(mai_mai_n2178_));
  NA2        m2129(.A(mai_mai_n1128_), .B(mai_mai_n688_), .Y(mai_mai_n2179_));
  AOI220     m2130(.A0(mai_mai_n2072_), .A1(mai_mai_n282_), .B0(mai_mai_n1283_), .B1(mai_mai_n1111_), .Y(mai_mai_n2180_));
  NA4        m2131(.A(mai_mai_n2180_), .B(mai_mai_n2179_), .C(mai_mai_n2178_), .D(mai_mai_n2176_), .Y(mai_mai_n2181_));
  AOI210     m2132(.A0(mai_mai_n2170_), .A1(x7), .B0(mai_mai_n2181_), .Y(mai_mai_n2182_));
  NA3        m2133(.A(mai_mai_n2182_), .B(mai_mai_n2164_), .C(mai_mai_n2144_), .Y(mai34));
  NA2        m2134(.A(mai_mai_n422_), .B(x4), .Y(mai_mai_n2184_));
  AOI210     m2135(.A0(mai_mai_n2515_), .A1(mai_mai_n2184_), .B0(mai_mai_n308_), .Y(mai_mai_n2185_));
  NA2        m2136(.A(mai_mai_n274_), .B(mai_mai_n112_), .Y(mai_mai_n2186_));
  NO2        m2137(.A(mai_mai_n928_), .B(mai_mai_n2186_), .Y(mai_mai_n2187_));
  AOI210     m2138(.A0(mai_mai_n1910_), .A1(mai_mai_n532_), .B0(mai_mai_n131_), .Y(mai_mai_n2188_));
  NA2        m2139(.A(mai_mai_n1836_), .B(x0), .Y(mai_mai_n2189_));
  OAI210     m2140(.A0(mai_mai_n1722_), .A1(mai_mai_n932_), .B0(mai_mai_n2189_), .Y(mai_mai_n2190_));
  NO4        m2141(.A(mai_mai_n2190_), .B(mai_mai_n2188_), .C(mai_mai_n2187_), .D(mai_mai_n2185_), .Y(mai_mai_n2191_));
  NO2        m2142(.A(mai_mai_n2191_), .B(mai_mai_n466_), .Y(mai_mai_n2192_));
  NA2        m2143(.A(mai_mai_n706_), .B(x8), .Y(mai_mai_n2193_));
  AO210      m2144(.A0(mai_mai_n2193_), .A1(mai_mai_n476_), .B0(mai_mai_n645_), .Y(mai_mai_n2194_));
  NA2        m2145(.A(mai_mai_n652_), .B(mai_mai_n613_), .Y(mai_mai_n2195_));
  AOI210     m2146(.A0(mai_mai_n2195_), .A1(mai_mai_n2194_), .B0(mai_mai_n252_), .Y(mai_mai_n2196_));
  OAI210     m2147(.A0(mai_mai_n111_), .A1(mai_mai_n1002_), .B0(mai_mai_n1388_), .Y(mai_mai_n2197_));
  OAI210     m2148(.A0(mai_mai_n1510_), .A1(mai_mai_n58_), .B0(mai_mai_n2197_), .Y(mai_mai_n2198_));
  NA3        m2149(.A(mai_mai_n2198_), .B(mai_mai_n328_), .C(x8), .Y(mai_mai_n2199_));
  NA2        m2150(.A(mai_mai_n1497_), .B(mai_mai_n316_), .Y(mai_mai_n2200_));
  NA2        m2151(.A(mai_mai_n648_), .B(mai_mai_n308_), .Y(mai_mai_n2201_));
  NA2        m2152(.A(mai_mai_n125_), .B(x0), .Y(mai_mai_n2202_));
  NAi31      m2153(.An(mai_mai_n2202_), .B(mai_mai_n2201_), .C(mai_mai_n764_), .Y(mai_mai_n2203_));
  NA3        m2154(.A(mai_mai_n2203_), .B(mai_mai_n2200_), .C(mai_mai_n2199_), .Y(mai_mai_n2204_));
  NA2        m2155(.A(mai_mai_n1052_), .B(mai_mai_n720_), .Y(mai_mai_n2205_));
  NA3        m2156(.A(mai_mai_n1089_), .B(mai_mai_n156_), .C(mai_mai_n1037_), .Y(mai_mai_n2206_));
  AOI210     m2157(.A0(mai_mai_n2206_), .A1(mai_mai_n2205_), .B0(mai_mai_n730_), .Y(mai_mai_n2207_));
  AOI210     m2158(.A0(mai_mai_n1675_), .A1(mai_mai_n121_), .B0(mai_mai_n2207_), .Y(mai_mai_n2208_));
  INV        m2159(.A(mai_mai_n241_), .Y(mai_mai_n2209_));
  NO2        m2160(.A(mai_mai_n2209_), .B(mai_mai_n59_), .Y(mai_mai_n2210_));
  NA3        m2161(.A(mai_mai_n2210_), .B(mai_mai_n706_), .C(mai_mai_n56_), .Y(mai_mai_n2211_));
  OAI210     m2162(.A0(mai_mai_n2208_), .A1(mai_mai_n132_), .B0(mai_mai_n2211_), .Y(mai_mai_n2212_));
  NO4        m2163(.A(mai_mai_n2212_), .B(mai_mai_n2204_), .C(mai_mai_n2196_), .D(mai_mai_n2192_), .Y(mai_mai_n2213_));
  NA2        m2164(.A(mai_mai_n755_), .B(mai_mai_n149_), .Y(mai_mai_n2214_));
  NO2        m2165(.A(mai_mai_n291_), .B(mai_mai_n1037_), .Y(mai_mai_n2215_));
  OAI220     m2166(.A0(mai_mai_n2215_), .A1(mai_mai_n1470_), .B0(mai_mai_n2214_), .B1(mai_mai_n1115_), .Y(mai_mai_n2216_));
  NA2        m2167(.A(mai_mai_n2216_), .B(x2), .Y(mai_mai_n2217_));
  OAI210     m2168(.A0(mai_mai_n825_), .A1(mai_mai_n359_), .B0(mai_mai_n2217_), .Y(mai_mai_n2218_));
  OAI220     m2169(.A0(mai_mai_n717_), .A1(mai_mai_n55_), .B0(mai_mai_n267_), .B1(mai_mai_n95_), .Y(mai_mai_n2219_));
  NO4        m2170(.A(mai_mai_n437_), .B(mai_mai_n71_), .C(x7), .D(x3), .Y(mai_mai_n2220_));
  NO2        m2171(.A(mai_mai_n1052_), .B(mai_mai_n275_), .Y(mai_mai_n2221_));
  NO4        m2172(.A(mai_mai_n2221_), .B(mai_mai_n2220_), .C(mai_mai_n2219_), .D(mai_mai_n2518_), .Y(mai_mai_n2222_));
  NA2        m2173(.A(mai_mai_n1180_), .B(mai_mai_n1000_), .Y(mai_mai_n2223_));
  NA4        m2174(.A(mai_mai_n706_), .B(mai_mai_n168_), .C(mai_mai_n57_), .D(mai_mai_n96_), .Y(mai_mai_n2224_));
  NA3        m2175(.A(mai_mai_n1319_), .B(mai_mai_n244_), .C(x7), .Y(mai_mai_n2225_));
  NA3        m2176(.A(mai_mai_n2225_), .B(mai_mai_n2224_), .C(mai_mai_n2223_), .Y(mai_mai_n2226_));
  OAI210     m2177(.A0(mai_mai_n2226_), .A1(mai_mai_n2222_), .B0(mai_mai_n153_), .Y(mai_mai_n2227_));
  NA3        m2178(.A(mai_mai_n822_), .B(mai_mai_n79_), .C(x0), .Y(mai_mai_n2228_));
  NA4        m2179(.A(mai_mai_n2228_), .B(mai_mai_n1093_), .C(mai_mai_n284_), .D(mai_mai_n574_), .Y(mai_mai_n2229_));
  NA2        m2180(.A(mai_mai_n1097_), .B(mai_mai_n657_), .Y(mai_mai_n2230_));
  NO2        m2181(.A(mai_mai_n2230_), .B(mai_mai_n253_), .Y(mai_mai_n2231_));
  AOI220     m2182(.A0(mai_mai_n2231_), .A1(x7), .B0(mai_mai_n967_), .B1(mai_mai_n646_), .Y(mai_mai_n2232_));
  OAI210     m2183(.A0(mai_mai_n1921_), .A1(mai_mai_n249_), .B0(mai_mai_n709_), .Y(mai_mai_n2233_));
  AOI220     m2184(.A0(mai_mai_n399_), .A1(x8), .B0(mai_mai_n84_), .B1(x2), .Y(mai_mai_n2234_));
  AOI210     m2185(.A0(mai_mai_n257_), .A1(mai_mai_n53_), .B0(mai_mai_n638_), .Y(mai_mai_n2235_));
  OAI220     m2186(.A0(mai_mai_n2235_), .A1(mai_mai_n89_), .B0(mai_mai_n2234_), .B1(mai_mai_n1271_), .Y(mai_mai_n2236_));
  AOI220     m2187(.A0(mai_mai_n2236_), .A1(mai_mai_n1255_), .B0(mai_mai_n2233_), .B1(mai_mai_n1431_), .Y(mai_mai_n2237_));
  NA4        m2188(.A(mai_mai_n2237_), .B(mai_mai_n2232_), .C(mai_mai_n2229_), .D(mai_mai_n2227_), .Y(mai_mai_n2238_));
  AOI210     m2189(.A0(mai_mai_n2218_), .A1(mai_mai_n778_), .B0(mai_mai_n2238_), .Y(mai_mai_n2239_));
  OAI210     m2190(.A0(mai_mai_n2213_), .A1(x2), .B0(mai_mai_n2239_), .Y(mai35));
  NA2        m2191(.A(mai_mai_n494_), .B(mai_mai_n168_), .Y(mai_mai_n2241_));
  AOI220     m2192(.A0(mai_mai_n621_), .A1(mai_mai_n55_), .B0(mai_mai_n745_), .B1(mai_mai_n1160_), .Y(mai_mai_n2242_));
  AOI210     m2193(.A0(mai_mai_n2242_), .A1(mai_mai_n2241_), .B0(mai_mai_n67_), .Y(mai_mai_n2243_));
  NO3        m2194(.A(mai_mai_n502_), .B(mai_mai_n456_), .C(mai_mai_n327_), .Y(mai_mai_n2244_));
  OAI210     m2195(.A0(mai_mai_n2244_), .A1(mai_mai_n2243_), .B0(x2), .Y(mai_mai_n2245_));
  AOI210     m2196(.A0(mai_mai_n206_), .A1(x0), .B0(mai_mai_n261_), .Y(mai_mai_n2246_));
  OAI220     m2197(.A0(mai_mai_n2246_), .A1(mai_mai_n650_), .B0(mai_mai_n188_), .B1(x4), .Y(mai_mai_n2247_));
  NA2        m2198(.A(mai_mai_n2247_), .B(mai_mai_n129_), .Y(mai_mai_n2248_));
  NA3        m2199(.A(mai_mai_n399_), .B(x8), .C(mai_mai_n67_), .Y(mai_mai_n2249_));
  AOI210     m2200(.A0(mai_mai_n2249_), .A1(mai_mai_n1622_), .B0(mai_mai_n666_), .Y(mai_mai_n2250_));
  OAI210     m2201(.A0(mai_mai_n2171_), .A1(x6), .B0(mai_mai_n719_), .Y(mai_mai_n2251_));
  NO2        m2202(.A(mai_mai_n2251_), .B(mai_mai_n2250_), .Y(mai_mai_n2252_));
  NA3        m2203(.A(mai_mai_n2252_), .B(mai_mai_n2248_), .C(mai_mai_n2245_), .Y(mai_mai_n2253_));
  INV        m2204(.A(mai_mai_n1232_), .Y(mai_mai_n2254_));
  NA2        m2205(.A(mai_mai_n2254_), .B(mai_mai_n56_), .Y(mai_mai_n2255_));
  NA2        m2206(.A(mai_mai_n734_), .B(mai_mai_n679_), .Y(mai_mai_n2256_));
  NA2        m2207(.A(mai_mai_n688_), .B(mai_mai_n209_), .Y(mai_mai_n2257_));
  NA2        m2208(.A(mai_mai_n1260_), .B(mai_mai_n62_), .Y(mai_mai_n2258_));
  OAI210     m2209(.A0(mai_mai_n1019_), .A1(x6), .B0(mai_mai_n461_), .Y(mai_mai_n2259_));
  NA3        m2210(.A(mai_mai_n2259_), .B(mai_mai_n2258_), .C(mai_mai_n2257_), .Y(mai_mai_n2260_));
  NA3        m2211(.A(mai_mai_n1208_), .B(mai_mai_n722_), .C(x3), .Y(mai_mai_n2261_));
  NO3        m2212(.A(mai_mai_n2261_), .B(mai_mai_n663_), .C(mai_mai_n197_), .Y(mai_mai_n2262_));
  AOI210     m2213(.A0(mai_mai_n2260_), .A1(mai_mai_n50_), .B0(mai_mai_n2262_), .Y(mai_mai_n2263_));
  OAI210     m2214(.A0(mai_mai_n2256_), .A1(mai_mai_n2255_), .B0(mai_mai_n2263_), .Y(mai_mai_n2264_));
  AOI210     m2215(.A0(mai_mai_n2253_), .A1(mai_mai_n57_), .B0(mai_mai_n2264_), .Y(mai_mai_n2265_));
  NA2        m2216(.A(mai_mai_n921_), .B(mai_mai_n62_), .Y(mai_mai_n2266_));
  NO3        m2217(.A(mai_mai_n1019_), .B(mai_mai_n554_), .C(mai_mai_n112_), .Y(mai_mai_n2267_));
  OAI210     m2218(.A0(mai_mai_n147_), .A1(mai_mai_n64_), .B0(mai_mai_n2267_), .Y(mai_mai_n2268_));
  AOI210     m2219(.A0(mai_mai_n2268_), .A1(mai_mai_n2266_), .B0(mai_mai_n50_), .Y(mai_mai_n2269_));
  NA4        m2220(.A(mai_mai_n456_), .B(mai_mai_n217_), .C(mai_mai_n830_), .D(mai_mai_n94_), .Y(mai_mai_n2270_));
  OAI210     m2221(.A0(mai_mai_n921_), .A1(mai_mai_n242_), .B0(mai_mai_n723_), .Y(mai_mai_n2271_));
  NA2        m2222(.A(mai_mai_n573_), .B(mai_mai_n2025_), .Y(mai_mai_n2272_));
  NA3        m2223(.A(mai_mai_n2272_), .B(mai_mai_n2271_), .C(mai_mai_n2270_), .Y(mai_mai_n2273_));
  OAI210     m2224(.A0(mai_mai_n2273_), .A1(mai_mai_n2269_), .B0(mai_mai_n59_), .Y(mai_mai_n2274_));
  AOI210     m2225(.A0(mai_mai_n822_), .A1(mai_mai_n523_), .B0(mai_mai_n1789_), .Y(mai_mai_n2275_));
  AOI210     m2226(.A0(mai_mai_n554_), .A1(mai_mai_n591_), .B0(mai_mai_n2275_), .Y(mai_mai_n2276_));
  NO4        m2227(.A(mai_mai_n913_), .B(mai_mai_n554_), .C(mai_mai_n351_), .D(mai_mai_n397_), .Y(mai_mai_n2277_));
  XN2        m2228(.A(x4), .B(x3), .Y(mai_mai_n2278_));
  NO3        m2229(.A(mai_mai_n2278_), .B(mai_mai_n649_), .C(mai_mai_n297_), .Y(mai_mai_n2279_));
  NO3        m2230(.A(mai_mai_n2279_), .B(mai_mai_n2277_), .C(mai_mai_n1386_), .Y(mai_mai_n2280_));
  OAI210     m2231(.A0(mai_mai_n2276_), .A1(x3), .B0(mai_mai_n2280_), .Y(mai_mai_n2281_));
  NA2        m2232(.A(mai_mai_n1386_), .B(mai_mai_n50_), .Y(mai_mai_n2282_));
  INV        m2233(.A(mai_mai_n2282_), .Y(mai_mai_n2283_));
  AOI210     m2234(.A0(mai_mai_n2281_), .A1(mai_mai_n576_), .B0(mai_mai_n2283_), .Y(mai_mai_n2284_));
  AOI210     m2235(.A0(mai_mai_n1359_), .A1(mai_mai_n628_), .B0(mai_mai_n663_), .Y(mai_mai_n2285_));
  NO2        m2236(.A(mai_mai_n830_), .B(mai_mai_n56_), .Y(mai_mai_n2286_));
  OAI210     m2237(.A0(mai_mai_n1839_), .A1(mai_mai_n591_), .B0(mai_mai_n2108_), .Y(mai_mai_n2287_));
  OAI210     m2238(.A0(mai_mai_n2193_), .A1(mai_mai_n2286_), .B0(mai_mai_n2287_), .Y(mai_mai_n2288_));
  OAI210     m2239(.A0(mai_mai_n2288_), .A1(mai_mai_n2285_), .B0(mai_mai_n84_), .Y(mai_mai_n2289_));
  NO2        m2240(.A(mai_mai_n815_), .B(mai_mai_n647_), .Y(mai_mai_n2290_));
  NO2        m2241(.A(mai_mai_n275_), .B(x6), .Y(mai_mai_n2291_));
  OAI210     m2242(.A0(mai_mai_n2290_), .A1(mai_mai_n1683_), .B0(mai_mai_n2291_), .Y(mai_mai_n2292_));
  NA4        m2243(.A(mai_mai_n2292_), .B(mai_mai_n2289_), .C(mai_mai_n2284_), .D(mai_mai_n2274_), .Y(mai_mai_n2293_));
  NA4        m2244(.A(mai_mai_n599_), .B(mai_mai_n666_), .C(mai_mai_n421_), .D(x6), .Y(mai_mai_n2294_));
  AOI210     m2245(.A0(mai_mai_n2294_), .A1(mai_mai_n416_), .B0(x1), .Y(mai_mai_n2295_));
  NO2        m2246(.A(mai_mai_n704_), .B(mai_mai_n663_), .Y(mai_mai_n2296_));
  OAI210     m2247(.A0(mai_mai_n456_), .A1(mai_mai_n157_), .B0(mai_mai_n761_), .Y(mai_mai_n2297_));
  AOI210     m2248(.A0(mai_mai_n2297_), .A1(mai_mai_n972_), .B0(mai_mai_n53_), .Y(mai_mai_n2298_));
  NO3        m2249(.A(mai_mai_n2298_), .B(mai_mai_n2296_), .C(mai_mai_n2295_), .Y(mai_mai_n2299_));
  NA3        m2250(.A(mai_mai_n1361_), .B(mai_mai_n1209_), .C(mai_mai_n782_), .Y(mai_mai_n2300_));
  AOI220     m2251(.A0(mai_mai_n1827_), .A1(mai_mai_n129_), .B0(mai_mai_n408_), .B1(mai_mai_n116_), .Y(mai_mai_n2301_));
  AOI210     m2252(.A0(mai_mai_n2301_), .A1(mai_mai_n2300_), .B0(mai_mai_n1424_), .Y(mai_mai_n2302_));
  NO2        m2253(.A(mai_mai_n621_), .B(x3), .Y(mai_mai_n2303_));
  NO3        m2254(.A(mai_mai_n674_), .B(mai_mai_n1510_), .C(x2), .Y(mai_mai_n2304_));
  AOI220     m2255(.A0(mai_mai_n2304_), .A1(mai_mai_n2303_), .B0(mai_mai_n1803_), .B1(mai_mai_n741_), .Y(mai_mai_n2305_));
  NA3        m2256(.A(x6), .B(x4), .C(x0), .Y(mai_mai_n2306_));
  OAI220     m2257(.A0(mai_mai_n2306_), .A1(mai_mai_n187_), .B0(mai_mai_n661_), .B1(mai_mai_n519_), .Y(mai_mai_n2307_));
  OAI220     m2258(.A0(mai_mai_n1245_), .A1(x8), .B0(mai_mai_n363_), .B1(mai_mai_n341_), .Y(mai_mai_n2308_));
  AOI220     m2259(.A0(mai_mai_n2308_), .A1(mai_mai_n408_), .B0(mai_mai_n2307_), .B1(mai_mai_n876_), .Y(mai_mai_n2309_));
  OAI210     m2260(.A0(mai_mai_n2305_), .A1(mai_mai_n1106_), .B0(mai_mai_n2309_), .Y(mai_mai_n2310_));
  NO2        m2261(.A(mai_mai_n2310_), .B(mai_mai_n2302_), .Y(mai_mai_n2311_));
  OAI210     m2262(.A0(mai_mai_n2299_), .A1(mai_mai_n301_), .B0(mai_mai_n2311_), .Y(mai_mai_n2312_));
  AOI210     m2263(.A0(mai_mai_n2293_), .A1(x5), .B0(mai_mai_n2312_), .Y(mai_mai_n2313_));
  OAI210     m2264(.A0(mai_mai_n2265_), .A1(x5), .B0(mai_mai_n2313_), .Y(mai36));
  NO2        m2265(.A(mai_mai_n824_), .B(mai_mai_n290_), .Y(mai_mai_n2315_));
  NO3        m2266(.A(mai_mai_n111_), .B(mai_mai_n1002_), .C(mai_mai_n55_), .Y(mai_mai_n2316_));
  NO3        m2267(.A(mai_mai_n2316_), .B(mai_mai_n1858_), .C(mai_mai_n1019_), .Y(mai_mai_n2317_));
  OAI210     m2268(.A0(mai_mai_n2317_), .A1(mai_mai_n2315_), .B0(mai_mai_n98_), .Y(mai_mai_n2318_));
  OR4        m2269(.A(mai_mai_n914_), .B(mai_mai_n771_), .C(mai_mai_n366_), .D(mai_mai_n483_), .Y(mai_mai_n2319_));
  INV        m2270(.A(mai_mai_n957_), .Y(mai_mai_n2320_));
  OAI210     m2271(.A0(mai_mai_n2072_), .A1(mai_mai_n2320_), .B0(mai_mai_n267_), .Y(mai_mai_n2321_));
  NA3        m2272(.A(mai_mai_n436_), .B(mai_mai_n214_), .C(mai_mai_n110_), .Y(mai_mai_n2322_));
  NA4        m2273(.A(mai_mai_n2322_), .B(mai_mai_n2321_), .C(mai_mai_n2319_), .D(mai_mai_n2318_), .Y(mai_mai_n2323_));
  NO2        m2274(.A(mai_mai_n947_), .B(x8), .Y(mai_mai_n2324_));
  NO3        m2275(.A(mai_mai_n2324_), .B(mai_mai_n944_), .C(mai_mai_n528_), .Y(mai_mai_n2325_));
  AOI220     m2276(.A0(mai_mai_n291_), .A1(x1), .B0(mai_mai_n128_), .B1(x6), .Y(mai_mai_n2326_));
  AOI210     m2277(.A0(mai_mai_n1037_), .A1(x6), .B0(mai_mai_n412_), .Y(mai_mai_n2327_));
  OAI220     m2278(.A0(mai_mai_n2327_), .A1(mai_mai_n350_), .B0(mai_mai_n2326_), .B1(mai_mai_n457_), .Y(mai_mai_n2328_));
  OAI210     m2279(.A0(mai_mai_n2328_), .A1(mai_mai_n2325_), .B0(mai_mai_n456_), .Y(mai_mai_n2329_));
  NA2        m2280(.A(mai_mai_n652_), .B(mai_mai_n483_), .Y(mai_mai_n2330_));
  AOI210     m2281(.A0(mai_mai_n2330_), .A1(mai_mai_n635_), .B0(mai_mai_n253_), .Y(mai_mai_n2331_));
  NO3        m2282(.A(mai_mai_n1764_), .B(mai_mai_n1509_), .C(mai_mai_n263_), .Y(mai_mai_n2332_));
  NO2        m2283(.A(mai_mai_n2266_), .B(mai_mai_n216_), .Y(mai_mai_n2333_));
  NO4        m2284(.A(mai_mai_n2333_), .B(mai_mai_n2332_), .C(mai_mai_n2331_), .D(mai_mai_n410_), .Y(mai_mai_n2334_));
  OAI210     m2285(.A0(mai_mai_n623_), .A1(mai_mai_n770_), .B0(mai_mai_n935_), .Y(mai_mai_n2335_));
  OAI220     m2286(.A0(mai_mai_n1554_), .A1(mai_mai_n1549_), .B0(mai_mai_n935_), .B1(mai_mai_n1037_), .Y(mai_mai_n2336_));
  AOI220     m2287(.A0(mai_mai_n2336_), .A1(mai_mai_n109_), .B0(mai_mai_n2335_), .B1(mai_mai_n613_), .Y(mai_mai_n2337_));
  NA3        m2288(.A(mai_mai_n2337_), .B(mai_mai_n2334_), .C(mai_mai_n2329_), .Y(mai_mai_n2338_));
  AOI210     m2289(.A0(mai_mai_n2323_), .A1(mai_mai_n328_), .B0(mai_mai_n2338_), .Y(mai_mai_n2339_));
  OAI210     m2290(.A0(mai_mai_n581_), .A1(mai_mai_n507_), .B0(mai_mai_n157_), .Y(mai_mai_n2340_));
  OAI210     m2291(.A0(mai_mai_n1871_), .A1(mai_mai_n66_), .B0(mai_mai_n2340_), .Y(mai_mai_n2341_));
  NA2        m2292(.A(mai_mai_n225_), .B(mai_mai_n242_), .Y(mai_mai_n2342_));
  NO2        m2293(.A(mai_mai_n1878_), .B(mai_mai_n164_), .Y(mai_mai_n2343_));
  NA2        m2294(.A(mai_mai_n1149_), .B(mai_mai_n55_), .Y(mai_mai_n2344_));
  OAI210     m2295(.A0(mai_mai_n2344_), .A1(mai_mai_n2343_), .B0(mai_mai_n2342_), .Y(mai_mai_n2345_));
  OAI210     m2296(.A0(mai_mai_n2345_), .A1(mai_mai_n2341_), .B0(mai_mai_n854_), .Y(mai_mai_n2346_));
  AOI210     m2297(.A0(mai_mai_n95_), .A1(mai_mai_n98_), .B0(mai_mai_n330_), .Y(mai_mai_n2347_));
  NA2        m2298(.A(mai_mai_n652_), .B(mai_mai_n1510_), .Y(mai_mai_n2348_));
  OAI220     m2299(.A0(mai_mai_n2348_), .A1(mai_mai_n2347_), .B0(mai_mai_n719_), .B1(mai_mai_n1193_), .Y(mai_mai_n2349_));
  NO2        m2300(.A(mai_mai_n1322_), .B(mai_mai_n568_), .Y(mai_mai_n2350_));
  NO3        m2301(.A(mai_mai_n2350_), .B(mai_mai_n1687_), .C(mai_mai_n674_), .Y(mai_mai_n2351_));
  NOi31      m2302(.An(mai_mai_n1890_), .B(mai_mai_n2160_), .C(mai_mai_n729_), .Y(mai_mai_n2352_));
  NO3        m2303(.A(mai_mai_n2352_), .B(mai_mai_n2351_), .C(mai_mai_n2349_), .Y(mai_mai_n2353_));
  AOI210     m2304(.A0(mai_mai_n2353_), .A1(mai_mai_n2346_), .B0(x7), .Y(mai_mai_n2354_));
  NA2        m2305(.A(mai_mai_n128_), .B(mai_mai_n62_), .Y(mai_mai_n2355_));
  AOI210     m2306(.A0(mai_mai_n576_), .A1(mai_mai_n608_), .B0(mai_mai_n1129_), .Y(mai_mai_n2356_));
  NA3        m2307(.A(mai_mai_n2356_), .B(mai_mai_n2355_), .C(mai_mai_n847_), .Y(mai_mai_n2357_));
  NA2        m2308(.A(mai_mai_n2357_), .B(mai_mai_n494_), .Y(mai_mai_n2358_));
  AOI220     m2309(.A0(mai_mai_n1645_), .A1(mai_mai_n245_), .B0(mai_mai_n1000_), .B1(mai_mai_n116_), .Y(mai_mai_n2359_));
  NO2        m2310(.A(mai_mai_n2359_), .B(mai_mai_n436_), .Y(mai_mai_n2360_));
  NO2        m2311(.A(mai_mai_n397_), .B(mai_mai_n214_), .Y(mai_mai_n2361_));
  NO3        m2312(.A(mai_mai_n2361_), .B(mai_mai_n1212_), .C(mai_mai_n59_), .Y(mai_mai_n2362_));
  AOI210     m2313(.A0(mai_mai_n1164_), .A1(mai_mai_n398_), .B0(x6), .Y(mai_mai_n2363_));
  NA3        m2314(.A(mai_mai_n1577_), .B(mai_mai_n267_), .C(mai_mai_n257_), .Y(mai_mai_n2364_));
  NA2        m2315(.A(mai_mai_n2364_), .B(mai_mai_n1535_), .Y(mai_mai_n2365_));
  NO4        m2316(.A(mai_mai_n2365_), .B(mai_mai_n2363_), .C(mai_mai_n2362_), .D(mai_mai_n2360_), .Y(mai_mai_n2366_));
  AOI210     m2317(.A0(mai_mai_n2366_), .A1(mai_mai_n2358_), .B0(mai_mai_n445_), .Y(mai_mai_n2367_));
  NO3        m2318(.A(mai_mai_n2278_), .B(mai_mai_n860_), .C(mai_mai_n493_), .Y(mai_mai_n2368_));
  AOI210     m2319(.A0(mai_mai_n1210_), .A1(mai_mai_n256_), .B0(mai_mai_n2368_), .Y(mai_mai_n2369_));
  OAI210     m2320(.A0(mai_mai_n828_), .A1(mai_mai_n262_), .B0(mai_mai_n387_), .Y(mai_mai_n2370_));
  NA2        m2321(.A(mai_mai_n1149_), .B(mai_mai_n162_), .Y(mai_mai_n2371_));
  NO2        m2322(.A(mai_mai_n598_), .B(mai_mai_n98_), .Y(mai_mai_n2372_));
  AO210      m2323(.A0(mai_mai_n2372_), .A1(mai_mai_n2371_), .B0(mai_mai_n1661_), .Y(mai_mai_n2373_));
  NO2        m2324(.A(mai_mai_n452_), .B(mai_mai_n409_), .Y(mai_mai_n2374_));
  AOI220     m2325(.A0(mai_mai_n2374_), .A1(mai_mai_n2373_), .B0(mai_mai_n2370_), .B1(mai_mai_n282_), .Y(mai_mai_n2375_));
  OAI210     m2326(.A0(mai_mai_n2369_), .A1(x1), .B0(mai_mai_n2375_), .Y(mai_mai_n2376_));
  NO3        m2327(.A(mai_mai_n2376_), .B(mai_mai_n2367_), .C(mai_mai_n2354_), .Y(mai_mai_n2377_));
  OAI210     m2328(.A0(mai_mai_n2339_), .A1(mai_mai_n57_), .B0(mai_mai_n2377_), .Y(mai37));
  NA3        m2329(.A(mai_mai_n1016_), .B(mai_mai_n131_), .C(x3), .Y(mai_mai_n2379_));
  NA3        m2330(.A(mai_mai_n755_), .B(mai_mai_n149_), .C(mai_mai_n50_), .Y(mai_mai_n2380_));
  AOI210     m2331(.A0(mai_mai_n2380_), .A1(mai_mai_n2379_), .B0(mai_mai_n667_), .Y(mai_mai_n2381_));
  NO3        m2332(.A(mai_mai_n1016_), .B(mai_mai_n366_), .C(mai_mai_n501_), .Y(mai_mai_n2382_));
  OAI210     m2333(.A0(mai_mai_n2382_), .A1(mai_mai_n2381_), .B0(mai_mai_n56_), .Y(mai_mai_n2383_));
  NA2        m2334(.A(mai_mai_n588_), .B(mai_mai_n720_), .Y(mai_mai_n2384_));
  AOI210     m2335(.A0(mai_mai_n2384_), .A1(mai_mai_n1001_), .B0(x3), .Y(mai_mai_n2385_));
  AOI220     m2336(.A0(mai_mai_n588_), .A1(mai_mai_n720_), .B0(mai_mai_n456_), .B1(mai_mai_n1000_), .Y(mai_mai_n2386_));
  NO2        m2337(.A(mai_mai_n649_), .B(mai_mai_n171_), .Y(mai_mai_n2387_));
  OAI220     m2338(.A0(mai_mai_n2387_), .A1(mai_mai_n802_), .B0(mai_mai_n2386_), .B1(mai_mai_n98_), .Y(mai_mai_n2388_));
  OAI210     m2339(.A0(mai_mai_n2388_), .A1(mai_mai_n2385_), .B0(mai_mai_n67_), .Y(mai_mai_n2389_));
  NA2        m2340(.A(mai_mai_n1131_), .B(mai_mai_n1019_), .Y(mai_mai_n2390_));
  NA2        m2341(.A(mai_mai_n1151_), .B(mai_mai_n446_), .Y(mai_mai_n2391_));
  NA4        m2342(.A(mai_mai_n2391_), .B(mai_mai_n2390_), .C(mai_mai_n2389_), .D(mai_mai_n2383_), .Y(mai_mai_n2392_));
  NA2        m2343(.A(mai_mai_n2392_), .B(mai_mai_n65_), .Y(mai_mai_n2393_));
  NO2        m2344(.A(mai_mai_n257_), .B(mai_mai_n1041_), .Y(mai_mai_n2394_));
  NA2        m2345(.A(mai_mai_n2394_), .B(mai_mai_n1002_), .Y(mai_mai_n2395_));
  OAI210     m2346(.A0(mai_mai_n217_), .A1(mai_mai_n209_), .B0(mai_mai_n1622_), .Y(mai_mai_n2396_));
  NA2        m2347(.A(mai_mai_n336_), .B(mai_mai_n261_), .Y(mai_mai_n2397_));
  NA3        m2348(.A(mai_mai_n393_), .B(mai_mai_n782_), .C(mai_mai_n98_), .Y(mai_mai_n2398_));
  NO2        m2349(.A(mai_mai_n520_), .B(mai_mai_n56_), .Y(mai_mai_n2399_));
  NA3        m2350(.A(mai_mai_n2399_), .B(mai_mai_n2398_), .C(mai_mai_n2397_), .Y(mai_mai_n2400_));
  AOI210     m2351(.A0(mai_mai_n2396_), .A1(mai_mai_n501_), .B0(mai_mai_n2400_), .Y(mai_mai_n2401_));
  NO2        m2352(.A(mai_mai_n1122_), .B(mai_mai_n262_), .Y(mai_mai_n2402_));
  OAI210     m2353(.A0(mai_mai_n282_), .A1(mai_mai_n251_), .B0(mai_mai_n2402_), .Y(mai_mai_n2403_));
  OAI210     m2354(.A0(mai_mai_n651_), .A1(mai_mai_n129_), .B0(x3), .Y(mai_mai_n2404_));
  AOI210     m2355(.A0(mai_mai_n651_), .A1(mai_mai_n355_), .B0(mai_mai_n2404_), .Y(mai_mai_n2405_));
  AOI210     m2356(.A0(mai_mai_n1510_), .A1(mai_mai_n50_), .B0(mai_mai_n336_), .Y(mai_mai_n2406_));
  OAI210     m2357(.A0(mai_mai_n2406_), .A1(mai_mai_n392_), .B0(mai_mai_n56_), .Y(mai_mai_n2407_));
  NO2        m2358(.A(mai_mai_n2407_), .B(mai_mai_n2405_), .Y(mai_mai_n2408_));
  AOI220     m2359(.A0(mai_mai_n2408_), .A1(mai_mai_n2403_), .B0(mai_mai_n2401_), .B1(mai_mai_n2395_), .Y(mai_mai_n2409_));
  OAI210     m2360(.A0(mai_mai_n2409_), .A1(mai_mai_n1659_), .B0(mai_mai_n93_), .Y(mai_mai_n2410_));
  NA2        m2361(.A(mai_mai_n674_), .B(mai_mai_n1135_), .Y(mai_mai_n2411_));
  NOi21      m2362(.An(mai_mai_n1289_), .B(mai_mai_n99_), .Y(mai_mai_n2412_));
  NA2        m2363(.A(mai_mai_n2412_), .B(mai_mai_n2411_), .Y(mai_mai_n2413_));
  NA2        m2364(.A(mai_mai_n2413_), .B(mai_mai_n1714_), .Y(mai_mai_n2414_));
  NA2        m2365(.A(mai_mai_n168_), .B(mai_mai_n96_), .Y(mai_mai_n2415_));
  NA2        m2366(.A(mai_mai_n666_), .B(x6), .Y(mai_mai_n2416_));
  AOI210     m2367(.A0(mai_mai_n2416_), .A1(mai_mai_n476_), .B0(mai_mai_n2415_), .Y(mai_mai_n2417_));
  AOI210     m2368(.A0(mai_mai_n343_), .A1(mai_mai_n131_), .B0(mai_mai_n132_), .Y(mai_mai_n2418_));
  OAI210     m2369(.A0(mai_mai_n2418_), .A1(mai_mai_n2417_), .B0(mai_mai_n336_), .Y(mai_mai_n2419_));
  AOI210     m2370(.A0(mai_mai_n599_), .A1(mai_mai_n425_), .B0(mai_mai_n1221_), .Y(mai_mai_n2420_));
  NO3        m2371(.A(mai_mai_n2420_), .B(mai_mai_n253_), .C(mai_mai_n62_), .Y(mai_mai_n2421_));
  OAI220     m2372(.A0(mai_mai_n2193_), .A1(mai_mai_n474_), .B0(mai_mai_n1964_), .B1(mai_mai_n376_), .Y(mai_mai_n2422_));
  OAI210     m2373(.A0(mai_mai_n2422_), .A1(mai_mai_n2421_), .B0(mai_mai_n53_), .Y(mai_mai_n2423_));
  NO4        m2374(.A(mai_mai_n2202_), .B(mai_mai_n894_), .C(mai_mai_n426_), .D(mai_mai_n212_), .Y(mai_mai_n2424_));
  NO4        m2375(.A(mai_mai_n706_), .B(mai_mai_n589_), .C(mai_mai_n434_), .D(mai_mai_n1010_), .Y(mai_mai_n2425_));
  NO2        m2376(.A(mai_mai_n2425_), .B(mai_mai_n2424_), .Y(mai_mai_n2426_));
  NA4        m2377(.A(mai_mai_n2426_), .B(mai_mai_n2423_), .C(mai_mai_n2419_), .D(mai_mai_n2414_), .Y(mai_mai_n2427_));
  NO3        m2378(.A(mai_mai_n237_), .B(mai_mai_n342_), .C(mai_mai_n76_), .Y(mai_mai_n2428_));
  NO3        m2379(.A(mai_mai_n53_), .B(mai_mai_n1149_), .C(mai_mai_n1166_), .Y(mai_mai_n2429_));
  OAI220     m2380(.A0(mai_mai_n2429_), .A1(mai_mai_n2428_), .B0(mai_mai_n456_), .B1(mai_mai_n77_), .Y(mai_mai_n2430_));
  OR2        m2381(.A(mai_mai_n900_), .B(mai_mai_n722_), .Y(mai_mai_n2431_));
  NA2        m2382(.A(mai_mai_n1160_), .B(mai_mai_n55_), .Y(mai_mai_n2432_));
  NOi21      m2383(.An(mai_mai_n2432_), .B(mai_mai_n377_), .Y(mai_mai_n2433_));
  AOI210     m2384(.A0(mai_mai_n2433_), .A1(mai_mai_n2431_), .B0(x1), .Y(mai_mai_n2434_));
  NA2        m2385(.A(mai_mai_n252_), .B(mai_mai_n76_), .Y(mai_mai_n2435_));
  AOI210     m2386(.A0(mai_mai_n1470_), .A1(mai_mai_n392_), .B0(mai_mai_n2435_), .Y(mai_mai_n2436_));
  NA2        m2387(.A(mai_mai_n1052_), .B(mai_mai_n61_), .Y(mai_mai_n2437_));
  NA2        m2388(.A(mai_mai_n1097_), .B(mai_mai_n164_), .Y(mai_mai_n2438_));
  OAI210     m2389(.A0(mai_mai_n2437_), .A1(mai_mai_n300_), .B0(mai_mai_n2438_), .Y(mai_mai_n2439_));
  NO3        m2390(.A(mai_mai_n2439_), .B(mai_mai_n2436_), .C(mai_mai_n2434_), .Y(mai_mai_n2440_));
  OAI210     m2391(.A0(mai_mai_n2440_), .A1(x6), .B0(mai_mai_n2430_), .Y(mai_mai_n2441_));
  AOI220     m2392(.A0(mai_mai_n2441_), .A1(mai_mai_n1388_), .B0(mai_mai_n2427_), .B1(mai_mai_n57_), .Y(mai_mai_n2442_));
  NA3        m2393(.A(mai_mai_n2442_), .B(mai_mai_n2410_), .C(mai_mai_n2393_), .Y(mai38));
  AOI210     m2394(.A0(mai_mai_n1564_), .A1(mai_mai_n177_), .B0(mai_mai_n930_), .Y(mai_mai_n2444_));
  AOI210     m2395(.A0(mai_mai_n1164_), .A1(mai_mai_n567_), .B0(mai_mai_n1034_), .Y(mai_mai_n2445_));
  AOI210     m2396(.A0(mai_mai_n2432_), .A1(mai_mai_n1742_), .B0(mai_mai_n216_), .Y(mai_mai_n2446_));
  NO3        m2397(.A(mai_mai_n1231_), .B(mai_mai_n308_), .C(x8), .Y(mai_mai_n2447_));
  NO4        m2398(.A(mai_mai_n2447_), .B(mai_mai_n2446_), .C(mai_mai_n2445_), .D(mai_mai_n2444_), .Y(mai_mai_n2448_));
  NO2        m2399(.A(mai_mai_n2448_), .B(x6), .Y(mai_mai_n2449_));
  NA4        m2400(.A(mai_mai_n368_), .B(mai_mai_n244_), .C(mai_mai_n180_), .D(x8), .Y(mai_mai_n2450_));
  NO2        m2401(.A(mai_mai_n2450_), .B(mai_mai_n132_), .Y(mai_mai_n2451_));
  AOI210     m2402(.A0(mai_mai_n426_), .A1(mai_mai_n396_), .B0(mai_mai_n1632_), .Y(mai_mai_n2452_));
  NO2        m2403(.A(mai_mai_n2452_), .B(mai_mai_n180_), .Y(mai_mai_n2453_));
  OAI210     m2404(.A0(mai_mai_n2453_), .A1(mai_mai_n2451_), .B0(x6), .Y(mai_mai_n2454_));
  INV        m2405(.A(mai_mai_n234_), .Y(mai_mai_n2455_));
  NO3        m2406(.A(mai_mai_n2455_), .B(mai_mai_n1586_), .C(mai_mai_n244_), .Y(mai_mai_n2456_));
  NO3        m2407(.A(x3), .B(mai_mai_n53_), .C(x0), .Y(mai_mai_n2457_));
  OAI210     m2408(.A0(mai_mai_n513_), .A1(x2), .B0(mai_mai_n2457_), .Y(mai_mai_n2458_));
  NA3        m2409(.A(mai_mai_n425_), .B(mai_mai_n415_), .C(mai_mai_n281_), .Y(mai_mai_n2459_));
  NA3        m2410(.A(mai_mai_n2459_), .B(mai_mai_n2458_), .C(mai_mai_n1704_), .Y(mai_mai_n2460_));
  OAI210     m2411(.A0(mai_mai_n2460_), .A1(mai_mai_n2456_), .B0(mai_mai_n778_), .Y(mai_mai_n2461_));
  NO2        m2412(.A(mai_mai_n589_), .B(mai_mai_n263_), .Y(mai_mai_n2462_));
  AN3        m2413(.A(mai_mai_n783_), .B(mai_mai_n755_), .C(x0), .Y(mai_mai_n2463_));
  OAI210     m2414(.A0(mai_mai_n2463_), .A1(mai_mai_n2462_), .B0(mai_mai_n317_), .Y(mai_mai_n2464_));
  NO2        m2415(.A(mai_mai_n782_), .B(mai_mai_n85_), .Y(mai_mai_n2465_));
  OAI210     m2416(.A0(mai_mai_n666_), .A1(x0), .B0(mai_mai_n51_), .Y(mai_mai_n2466_));
  AOI210     m2417(.A0(mai_mai_n572_), .A1(x4), .B0(mai_mai_n215_), .Y(mai_mai_n2467_));
  AOI220     m2418(.A0(mai_mai_n2467_), .A1(mai_mai_n2466_), .B0(mai_mai_n2465_), .B1(mai_mai_n393_), .Y(mai_mai_n2468_));
  NA4        m2419(.A(mai_mai_n2468_), .B(mai_mai_n2464_), .C(mai_mai_n2461_), .D(mai_mai_n2454_), .Y(mai_mai_n2469_));
  OAI210     m2420(.A0(mai_mai_n2469_), .A1(mai_mai_n2449_), .B0(x7), .Y(mai_mai_n2470_));
  NA2        m2421(.A(mai_mai_n364_), .B(x1), .Y(mai_mai_n2471_));
  NO2        m2422(.A(mai_mai_n2471_), .B(mai_mai_n51_), .Y(mai_mai_n2472_));
  AOI210     m2423(.A0(mai_mai_n84_), .A1(mai_mai_n67_), .B0(mai_mai_n2108_), .Y(mai_mai_n2473_));
  NA2        m2424(.A(mai_mai_n376_), .B(x3), .Y(mai_mai_n2474_));
  NO2        m2425(.A(mai_mai_n1651_), .B(mai_mai_n520_), .Y(mai_mai_n2475_));
  OAI210     m2426(.A0(mai_mai_n2474_), .A1(mai_mai_n2473_), .B0(mai_mai_n2475_), .Y(mai_mai_n2476_));
  OAI210     m2427(.A0(mai_mai_n2476_), .A1(mai_mai_n2472_), .B0(x4), .Y(mai_mai_n2477_));
  NO2        m2428(.A(mai_mai_n1662_), .B(mai_mai_n450_), .Y(mai_mai_n2478_));
  NO3        m2429(.A(mai_mai_n2478_), .B(mai_mai_n392_), .C(mai_mai_n109_), .Y(mai_mai_n2479_));
  AOI210     m2430(.A0(mai_mai_n1010_), .A1(mai_mai_n228_), .B0(mai_mai_n385_), .Y(mai_mai_n2480_));
  AO210      m2431(.A0(mai_mai_n1237_), .A1(x6), .B0(mai_mai_n2480_), .Y(mai_mai_n2481_));
  NO2        m2432(.A(mai_mai_n1344_), .B(mai_mai_n129_), .Y(mai_mai_n2482_));
  NA2        m2433(.A(mai_mai_n1836_), .B(mai_mai_n311_), .Y(mai_mai_n2483_));
  OAI220     m2434(.A0(mai_mai_n2483_), .A1(mai_mai_n1024_), .B0(mai_mai_n2482_), .B1(mai_mai_n1727_), .Y(mai_mai_n2484_));
  NO3        m2435(.A(mai_mai_n2484_), .B(mai_mai_n2481_), .C(mai_mai_n2479_), .Y(mai_mai_n2485_));
  AOI210     m2436(.A0(mai_mai_n2485_), .A1(mai_mai_n2477_), .B0(mai_mai_n96_), .Y(mai_mai_n2486_));
  NA3        m2437(.A(mai_mai_n1827_), .B(mai_mai_n589_), .C(mai_mai_n153_), .Y(mai_mai_n2487_));
  AOI210     m2438(.A0(mai_mai_n2487_), .A1(mai_mai_n1355_), .B0(mai_mai_n217_), .Y(mai_mai_n2488_));
  AOI210     m2439(.A0(mai_mai_n494_), .A1(mai_mai_n483_), .B0(mai_mai_n662_), .Y(mai_mai_n2489_));
  OAI220     m2440(.A0(mai_mai_n2489_), .A1(mai_mai_n457_), .B0(mai_mai_n188_), .B1(mai_mai_n107_), .Y(mai_mai_n2490_));
  OAI210     m2441(.A0(mai_mai_n2490_), .A1(mai_mai_n2488_), .B0(x0), .Y(mai_mai_n2491_));
  NA3        m2442(.A(mai_mai_n396_), .B(mai_mai_n782_), .C(mai_mai_n263_), .Y(mai_mai_n2492_));
  NO2        m2443(.A(mai_mai_n2492_), .B(mai_mai_n2067_), .Y(mai_mai_n2493_));
  NA4        m2444(.A(mai_mai_n661_), .B(mai_mai_n589_), .C(mai_mai_n168_), .D(x3), .Y(mai_mai_n2494_));
  NO2        m2445(.A(mai_mai_n2494_), .B(mai_mai_n488_), .Y(mai_mai_n2495_));
  OAI220     m2446(.A0(mai_mai_n1681_), .A1(mai_mai_n2148_), .B0(mai_mai_n215_), .B1(mai_mai_n141_), .Y(mai_mai_n2496_));
  NO3        m2447(.A(mai_mai_n2496_), .B(mai_mai_n2495_), .C(mai_mai_n2493_), .Y(mai_mai_n2497_));
  NA2        m2448(.A(mai_mai_n2497_), .B(mai_mai_n2491_), .Y(mai_mai_n2498_));
  OAI210     m2449(.A0(mai_mai_n2498_), .A1(mai_mai_n2486_), .B0(mai_mai_n57_), .Y(mai_mai_n2499_));
  AOI210     m2450(.A0(mai_mai_n1715_), .A1(mai_mai_n263_), .B0(mai_mai_n663_), .Y(mai_mai_n2500_));
  NO2        m2451(.A(mai_mai_n1658_), .B(mai_mai_n204_), .Y(mai_mai_n2501_));
  OAI210     m2452(.A0(mai_mai_n2501_), .A1(mai_mai_n2500_), .B0(mai_mai_n615_), .Y(mai_mai_n2502_));
  OAI220     m2453(.A0(mai_mai_n1665_), .A1(mai_mai_n263_), .B0(mai_mai_n243_), .B1(mai_mai_n94_), .Y(mai_mai_n2503_));
  NA2        m2454(.A(mai_mai_n1758_), .B(mai_mai_n344_), .Y(mai_mai_n2504_));
  OAI220     m2455(.A0(mai_mai_n2504_), .A1(mai_mai_n623_), .B0(mai_mai_n673_), .B1(mai_mai_n141_), .Y(mai_mai_n2505_));
  AOI210     m2456(.A0(mai_mai_n2503_), .A1(mai_mai_n947_), .B0(mai_mai_n2505_), .Y(mai_mai_n2506_));
  NA4        m2457(.A(mai_mai_n2506_), .B(mai_mai_n2502_), .C(mai_mai_n2499_), .D(mai_mai_n2470_), .Y(mai39));
  INV        m2458(.A(mai_mai_n112_), .Y(mai_mai_n2510_));
  INV        m2459(.A(mai_mai_n129_), .Y(mai_mai_n2511_));
  INV        m2460(.A(x8), .Y(mai_mai_n2512_));
  INV        m2461(.A(x6), .Y(mai_mai_n2513_));
  INV        m2462(.A(mai_mai_n111_), .Y(mai_mai_n2514_));
  INV        m2463(.A(mai_mai_n817_), .Y(mai_mai_n2515_));
  INV        m2464(.A(mai_mai_n717_), .Y(mai_mai_n2516_));
  INV        m2465(.A(mai_mai_n924_), .Y(mai_mai_n2517_));
  INV        m2466(.A(x4), .Y(mai_mai_n2518_));
  INV        m2467(.A(mai_mai_n1858_), .Y(mai_mai_n2519_));
  INV        u0000(.A(x3), .Y(men_men_n50_));
  NA2        u0001(.A(men_men_n50_), .B(x2), .Y(men_men_n51_));
  NA2        u0002(.A(x7), .B(x0), .Y(men_men_n52_));
  INV        u0003(.A(x1), .Y(men_men_n53_));
  NA2        u0004(.A(x5), .B(men_men_n53_), .Y(men_men_n54_));
  INV        u0005(.A(x8), .Y(men_men_n55_));
  INV        u0006(.A(x4), .Y(men_men_n56_));
  INV        u0007(.A(x7), .Y(men_men_n57_));
  NA2        u0008(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0009(.A(x0), .Y(men_men_n59_));
  NA2        u0010(.A(x4), .B(men_men_n59_), .Y(men_men_n60_));
  NA4        u0011(.A(men_men_n60_), .B(men_men_n58_), .C(men_men_n55_), .D(x6), .Y(men_men_n61_));
  NA2        u0012(.A(men_men_n56_), .B(men_men_n59_), .Y(men_men_n62_));
  NO2        u0013(.A(men_men_n55_), .B(x6), .Y(men_men_n63_));
  NA2        u0014(.A(men_men_n57_), .B(x4), .Y(men_men_n64_));
  NA3        u0015(.A(men_men_n64_), .B(men_men_n63_), .C(men_men_n62_), .Y(men_men_n65_));
  AOI210     u0016(.A0(men_men_n65_), .A1(men_men_n61_), .B0(men_men_n54_), .Y(men_men_n66_));
  NO2        u0017(.A(x8), .B(men_men_n57_), .Y(men_men_n67_));
  NO2        u0018(.A(x7), .B(men_men_n59_), .Y(men_men_n68_));
  NO2        u0019(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi21      u0020(.An(x5), .B(x1), .Y(men_men_n70_));
  INV        u0021(.A(x6), .Y(men_men_n71_));
  NA2        u0022(.A(men_men_n71_), .B(x4), .Y(men_men_n72_));
  NO3        u0023(.A(men_men_n72_), .B(men_men_n70_), .C(men_men_n69_), .Y(men_men_n73_));
  OAI210     u0024(.A0(men_men_n73_), .A1(men_men_n66_), .B0(men_men_n52_), .Y(men_men_n74_));
  NA2        u0025(.A(x7), .B(x4), .Y(men_men_n75_));
  NO2        u0026(.A(men_men_n75_), .B(x1), .Y(men_men_n76_));
  NO2        u0027(.A(men_men_n71_), .B(x5), .Y(men_men_n77_));
  NO2        u0028(.A(x8), .B(men_men_n59_), .Y(men_men_n78_));
  NA3        u0029(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n76_), .Y(men_men_n79_));
  AOI210     u0030(.A0(men_men_n79_), .A1(men_men_n74_), .B0(men_men_n51_), .Y(men_men_n80_));
  NA2        u0031(.A(x5), .B(x3), .Y(men_men_n81_));
  NO2        u0032(.A(x6), .B(x0), .Y(men_men_n82_));
  NO2        u0033(.A(men_men_n82_), .B(x4), .Y(men_men_n83_));
  NO2        u0034(.A(x4), .B(x2), .Y(men_men_n84_));
  NO2        u0035(.A(men_men_n71_), .B(men_men_n59_), .Y(men_men_n85_));
  NO2        u0036(.A(men_men_n85_), .B(men_men_n84_), .Y(men_men_n86_));
  NA2        u0037(.A(x8), .B(x1), .Y(men_men_n87_));
  NO2        u0038(.A(men_men_n87_), .B(x7), .Y(men_men_n88_));
  OR3        u0039(.A(men_men_n87_), .B(men_men_n86_), .C(men_men_n83_), .Y(men_men_n89_));
  NO3        u0040(.A(x8), .B(men_men_n57_), .C(x6), .Y(men_men_n90_));
  NO2        u0041(.A(x1), .B(men_men_n59_), .Y(men_men_n91_));
  NO2        u0042(.A(men_men_n56_), .B(x2), .Y(men_men_n92_));
  NA3        u0043(.A(men_men_n92_), .B(men_men_n91_), .C(men_men_n90_), .Y(men_men_n93_));
  AOI210     u0044(.A0(men_men_n93_), .A1(men_men_n89_), .B0(men_men_n81_), .Y(men_men_n94_));
  XO2        u0045(.A(x7), .B(x1), .Y(men_men_n95_));
  INV        u0046(.A(men_men_n95_), .Y(men_men_n96_));
  NO2        u0047(.A(men_men_n96_), .B(x6), .Y(men_men_n97_));
  NO2        u0048(.A(men_men_n50_), .B(x0), .Y(men_men_n98_));
  NA2        u0049(.A(men_men_n98_), .B(men_men_n55_), .Y(men_men_n99_));
  NO2        u0050(.A(x6), .B(x5), .Y(men_men_n100_));
  NO2        u0051(.A(men_men_n57_), .B(x5), .Y(men_men_n101_));
  NO2        u0052(.A(men_men_n101_), .B(men_men_n100_), .Y(men_men_n102_));
  NA2        u0053(.A(x6), .B(x1), .Y(men_men_n103_));
  NA2        u0054(.A(men_men_n103_), .B(men_men_n84_), .Y(men_men_n104_));
  NO4        u0055(.A(men_men_n104_), .B(men_men_n102_), .C(men_men_n99_), .D(men_men_n97_), .Y(men_men_n105_));
  NA2        u0056(.A(x3), .B(x0), .Y(men_men_n106_));
  INV        u0057(.A(x5), .Y(men_men_n107_));
  NA2        u0058(.A(men_men_n71_), .B(men_men_n107_), .Y(men_men_n108_));
  INV        u0059(.A(x2), .Y(men_men_n109_));
  NO2        u0060(.A(men_men_n56_), .B(men_men_n109_), .Y(men_men_n110_));
  NA2        u0061(.A(men_men_n57_), .B(men_men_n107_), .Y(men_men_n111_));
  NA3        u0062(.A(men_men_n111_), .B(men_men_n110_), .C(men_men_n108_), .Y(men_men_n112_));
  NO3        u0063(.A(men_men_n112_), .B(men_men_n106_), .C(men_men_n53_), .Y(men_men_n113_));
  NO4        u0064(.A(men_men_n113_), .B(men_men_n105_), .C(men_men_n94_), .D(men_men_n80_), .Y(men00));
  NO2        u0065(.A(x7), .B(x6), .Y(men_men_n115_));
  INV        u0066(.A(men_men_n115_), .Y(men_men_n116_));
  NO2        u0067(.A(men_men_n55_), .B(men_men_n53_), .Y(men_men_n117_));
  NA2        u0068(.A(men_men_n117_), .B(men_men_n56_), .Y(men_men_n118_));
  NO2        u0069(.A(men_men_n118_), .B(men_men_n116_), .Y(men_men_n119_));
  XN2        u0070(.A(x6), .B(x1), .Y(men_men_n120_));
  INV        u0071(.A(men_men_n120_), .Y(men_men_n121_));
  NO2        u0072(.A(x6), .B(x4), .Y(men_men_n122_));
  NA2        u0073(.A(x6), .B(x4), .Y(men_men_n123_));
  NAi21      u0074(.An(men_men_n122_), .B(men_men_n123_), .Y(men_men_n124_));
  XN2        u0075(.A(x7), .B(x6), .Y(men_men_n125_));
  NO4        u0076(.A(men_men_n125_), .B(men_men_n124_), .C(men_men_n121_), .D(x8), .Y(men_men_n126_));
  NO2        u0077(.A(x3), .B(men_men_n109_), .Y(men_men_n127_));
  NA2        u0078(.A(men_men_n127_), .B(men_men_n107_), .Y(men_men_n128_));
  NO2        u0079(.A(men_men_n128_), .B(men_men_n59_), .Y(men_men_n129_));
  OAI210     u0080(.A0(men_men_n126_), .A1(men_men_n119_), .B0(men_men_n129_), .Y(men_men_n130_));
  NA2        u0081(.A(x3), .B(men_men_n109_), .Y(men_men_n131_));
  NO2        u0082(.A(men_men_n55_), .B(men_men_n57_), .Y(men_men_n132_));
  NA2        u0083(.A(men_men_n132_), .B(men_men_n56_), .Y(men_men_n133_));
  NA2        u0084(.A(men_men_n55_), .B(men_men_n57_), .Y(men_men_n134_));
  NA2        u0085(.A(men_men_n134_), .B(x2), .Y(men_men_n135_));
  NA2        u0086(.A(x8), .B(x3), .Y(men_men_n136_));
  NA2        u0087(.A(men_men_n136_), .B(men_men_n75_), .Y(men_men_n137_));
  OAI220     u0088(.A0(men_men_n137_), .A1(men_men_n135_), .B0(men_men_n133_), .B1(men_men_n131_), .Y(men_men_n138_));
  NO2        u0089(.A(x5), .B(x0), .Y(men_men_n139_));
  NO2        u0090(.A(x6), .B(x1), .Y(men_men_n140_));
  NA3        u0091(.A(men_men_n140_), .B(men_men_n139_), .C(men_men_n138_), .Y(men_men_n141_));
  NA2        u0092(.A(x8), .B(men_men_n107_), .Y(men_men_n142_));
  NA2        u0093(.A(x4), .B(men_men_n50_), .Y(men_men_n143_));
  NO3        u0094(.A(men_men_n143_), .B(men_men_n142_), .C(men_men_n103_), .Y(men_men_n144_));
  NAi21      u0095(.An(x7), .B(x2), .Y(men_men_n145_));
  NO2        u0096(.A(men_men_n145_), .B(x0), .Y(men_men_n146_));
  XO2        u0097(.A(x8), .B(x7), .Y(men_men_n147_));
  NA2        u0098(.A(men_men_n147_), .B(men_men_n109_), .Y(men_men_n148_));
  NA2        u0099(.A(x6), .B(x5), .Y(men_men_n149_));
  NO2        u0100(.A(men_men_n56_), .B(x0), .Y(men_men_n150_));
  NO2        u0101(.A(men_men_n50_), .B(x1), .Y(men_men_n151_));
  NA2        u0102(.A(men_men_n151_), .B(men_men_n150_), .Y(men_men_n152_));
  NO3        u0103(.A(men_men_n152_), .B(men_men_n149_), .C(men_men_n148_), .Y(men_men_n153_));
  AOI210     u0104(.A0(men_men_n146_), .A1(men_men_n144_), .B0(men_men_n153_), .Y(men_men_n154_));
  NA3        u0105(.A(men_men_n154_), .B(men_men_n141_), .C(men_men_n130_), .Y(men01));
  NA2        u0106(.A(men_men_n57_), .B(men_men_n59_), .Y(men_men_n156_));
  NO2        u0107(.A(x2), .B(x1), .Y(men_men_n157_));
  NA2        u0108(.A(x2), .B(x1), .Y(men_men_n158_));
  NOi21      u0109(.An(men_men_n158_), .B(men_men_n157_), .Y(men_men_n159_));
  NA2        u0110(.A(men_men_n107_), .B(men_men_n53_), .Y(men_men_n160_));
  NO2        u0111(.A(men_men_n160_), .B(x8), .Y(men_men_n161_));
  NAi21      u0112(.An(x8), .B(x1), .Y(men_men_n162_));
  NO2        u0113(.A(men_men_n162_), .B(x3), .Y(men_men_n163_));
  OAI210     u0114(.A0(men_men_n163_), .A1(men_men_n161_), .B0(men_men_n159_), .Y(men_men_n164_));
  NO2        u0115(.A(x5), .B(men_men_n50_), .Y(men_men_n165_));
  NO2        u0116(.A(men_men_n109_), .B(x1), .Y(men_men_n166_));
  NA2        u0117(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  AOI210     u0118(.A0(men_men_n167_), .A1(men_men_n164_), .B0(men_men_n156_), .Y(men_men_n168_));
  NAi21      u0119(.An(x7), .B(x0), .Y(men_men_n169_));
  NO2        u0120(.A(men_men_n55_), .B(x2), .Y(men_men_n170_));
  NO2        u0121(.A(men_men_n81_), .B(x1), .Y(men_men_n171_));
  NA2        u0122(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  NA2        u0123(.A(x5), .B(men_men_n50_), .Y(men_men_n173_));
  NO2        u0124(.A(men_men_n173_), .B(men_men_n162_), .Y(men_men_n174_));
  NA2        u0125(.A(x8), .B(x5), .Y(men_men_n175_));
  NO2        u0126(.A(men_men_n175_), .B(men_men_n51_), .Y(men_men_n176_));
  NO3        u0127(.A(x3), .B(men_men_n109_), .C(men_men_n53_), .Y(men_men_n177_));
  NO3        u0128(.A(men_men_n177_), .B(men_men_n176_), .C(men_men_n174_), .Y(men_men_n178_));
  AOI210     u0129(.A0(men_men_n178_), .A1(men_men_n172_), .B0(men_men_n169_), .Y(men_men_n179_));
  NO2        u0130(.A(men_men_n57_), .B(x3), .Y(men_men_n180_));
  NO2        u0131(.A(men_men_n55_), .B(x0), .Y(men_men_n181_));
  NA3        u0132(.A(men_men_n107_), .B(men_men_n109_), .C(x1), .Y(men_men_n182_));
  NO2        u0133(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  NO2        u0134(.A(men_men_n87_), .B(men_men_n50_), .Y(men_men_n184_));
  NA2        u0135(.A(men_men_n107_), .B(x0), .Y(men_men_n185_));
  NO2        u0136(.A(men_men_n185_), .B(x2), .Y(men_men_n186_));
  AOI220     u0137(.A0(men_men_n186_), .A1(men_men_n184_), .B0(men_men_n183_), .B1(men_men_n180_), .Y(men_men_n187_));
  NA2        u0138(.A(x7), .B(men_men_n109_), .Y(men_men_n188_));
  NA2        u0139(.A(men_men_n165_), .B(x8), .Y(men_men_n189_));
  NA4        u0140(.A(x5), .B(x3), .C(x1), .D(x0), .Y(men_men_n190_));
  OR2        u0141(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n191_));
  NO2        u0142(.A(men_men_n158_), .B(men_men_n50_), .Y(men_men_n192_));
  NAi21      u0143(.An(x1), .B(x2), .Y(men_men_n193_));
  NO2        u0144(.A(men_men_n173_), .B(men_men_n193_), .Y(men_men_n194_));
  NA2        u0145(.A(x8), .B(x7), .Y(men_men_n195_));
  NO2        u0146(.A(men_men_n195_), .B(x0), .Y(men_men_n196_));
  OAI210     u0147(.A0(men_men_n194_), .A1(men_men_n192_), .B0(men_men_n196_), .Y(men_men_n197_));
  NA3        u0148(.A(men_men_n197_), .B(men_men_n191_), .C(men_men_n187_), .Y(men_men_n198_));
  NO3        u0149(.A(men_men_n198_), .B(men_men_n179_), .C(men_men_n168_), .Y(men_men_n199_));
  NA2        u0150(.A(x3), .B(x1), .Y(men_men_n200_));
  NA2        u0151(.A(men_men_n50_), .B(men_men_n109_), .Y(men_men_n201_));
  NO2        u0152(.A(men_men_n201_), .B(men_men_n70_), .Y(men_men_n202_));
  OAI210     u0153(.A0(men_men_n202_), .A1(men_men_n194_), .B0(men_men_n67_), .Y(men_men_n203_));
  NA2        u0154(.A(men_men_n132_), .B(men_men_n109_), .Y(men_men_n204_));
  OAI210     u0155(.A0(men_men_n204_), .A1(men_men_n200_), .B0(men_men_n203_), .Y(men_men_n205_));
  XO2        u0156(.A(x5), .B(x3), .Y(men_men_n206_));
  NA2        u0157(.A(men_men_n206_), .B(x8), .Y(men_men_n207_));
  NA2        u0158(.A(x8), .B(men_men_n59_), .Y(men_men_n208_));
  NA2        u0159(.A(men_men_n208_), .B(men_men_n136_), .Y(men_men_n209_));
  NA2        u0160(.A(x7), .B(men_men_n71_), .Y(men_men_n210_));
  NO2        u0161(.A(men_men_n193_), .B(men_men_n210_), .Y(men_men_n211_));
  OA210      u0162(.A0(men_men_n209_), .A1(men_men_n206_), .B0(men_men_n211_), .Y(men_men_n212_));
  AOI220     u0163(.A0(men_men_n212_), .A1(men_men_n207_), .B0(men_men_n205_), .B1(x0), .Y(men_men_n213_));
  OAI210     u0164(.A0(men_men_n199_), .A1(men_men_n71_), .B0(men_men_n213_), .Y(men_men_n214_));
  NO2        u0165(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n215_));
  NA2        u0166(.A(x8), .B(men_men_n50_), .Y(men_men_n216_));
  NA2        u0167(.A(men_men_n216_), .B(x2), .Y(men_men_n217_));
  NA2        u0168(.A(men_men_n55_), .B(x3), .Y(men_men_n218_));
  NA4        u0169(.A(men_men_n218_), .B(men_men_n217_), .C(men_men_n206_), .D(men_men_n82_), .Y(men_men_n219_));
  NO2        u0170(.A(men_men_n219_), .B(men_men_n53_), .Y(men_men_n220_));
  NO2        u0171(.A(men_men_n109_), .B(men_men_n59_), .Y(men_men_n221_));
  NA2        u0172(.A(x5), .B(x1), .Y(men_men_n222_));
  NO2        u0173(.A(men_men_n222_), .B(x6), .Y(men_men_n223_));
  NO2        u0174(.A(x3), .B(x1), .Y(men_men_n224_));
  AOI210     u0175(.A0(men_men_n224_), .A1(men_men_n77_), .B0(men_men_n223_), .Y(men_men_n225_));
  NO2        u0176(.A(men_men_n81_), .B(men_men_n55_), .Y(men_men_n226_));
  NO2        u0177(.A(men_men_n103_), .B(men_men_n50_), .Y(men_men_n227_));
  NO2        u0178(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n228_));
  OAI210     u0179(.A0(men_men_n225_), .A1(x8), .B0(men_men_n228_), .Y(men_men_n229_));
  NO2        u0180(.A(men_men_n55_), .B(x5), .Y(men_men_n230_));
  NA2        u0181(.A(men_men_n230_), .B(men_men_n71_), .Y(men_men_n231_));
  NAi21      u0182(.An(x2), .B(x5), .Y(men_men_n232_));
  NA2        u0183(.A(x8), .B(x6), .Y(men_men_n233_));
  OAI210     u0184(.A0(men_men_n233_), .A1(men_men_n232_), .B0(men_men_n231_), .Y(men_men_n234_));
  NA2        u0185(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n235_));
  NO2        u0186(.A(men_men_n235_), .B(men_men_n59_), .Y(men_men_n236_));
  AO220      u0187(.A0(men_men_n236_), .A1(men_men_n234_), .B0(men_men_n229_), .B1(men_men_n221_), .Y(men_men_n237_));
  OAI210     u0188(.A0(men_men_n237_), .A1(men_men_n220_), .B0(men_men_n215_), .Y(men_men_n238_));
  NA2        u0189(.A(men_men_n71_), .B(men_men_n56_), .Y(men_men_n239_));
  NO2        u0190(.A(men_men_n239_), .B(x7), .Y(men_men_n240_));
  NO2        u0191(.A(men_men_n107_), .B(men_men_n53_), .Y(men_men_n241_));
  NA2        u0192(.A(men_men_n241_), .B(men_men_n109_), .Y(men_men_n242_));
  AOI210     u0193(.A0(men_men_n242_), .A1(men_men_n167_), .B0(men_men_n59_), .Y(men_men_n243_));
  NA2        u0194(.A(x3), .B(men_men_n59_), .Y(men_men_n244_));
  NO2        u0195(.A(men_men_n182_), .B(men_men_n244_), .Y(men_men_n245_));
  OA210      u0196(.A0(men_men_n245_), .A1(men_men_n243_), .B0(x8), .Y(men_men_n246_));
  NO2        u0197(.A(x1), .B(x0), .Y(men_men_n247_));
  NA2        u0198(.A(men_men_n247_), .B(men_men_n109_), .Y(men_men_n248_));
  NA2        u0199(.A(men_men_n107_), .B(men_men_n50_), .Y(men_men_n249_));
  XN2        u0200(.A(x3), .B(x2), .Y(men_men_n250_));
  NA2        u0201(.A(men_men_n250_), .B(men_men_n159_), .Y(men_men_n251_));
  NO2        u0202(.A(men_men_n107_), .B(x0), .Y(men_men_n252_));
  NA2        u0203(.A(x8), .B(men_men_n53_), .Y(men_men_n253_));
  NA2        u0204(.A(men_men_n253_), .B(men_men_n252_), .Y(men_men_n254_));
  OAI220     u0205(.A0(men_men_n254_), .A1(men_men_n251_), .B0(men_men_n249_), .B1(men_men_n248_), .Y(men_men_n255_));
  OAI210     u0206(.A0(men_men_n255_), .A1(men_men_n246_), .B0(men_men_n240_), .Y(men_men_n256_));
  NO2        u0207(.A(x7), .B(x1), .Y(men_men_n257_));
  NOi21      u0208(.An(x8), .B(x3), .Y(men_men_n258_));
  NA2        u0209(.A(men_men_n258_), .B(men_men_n59_), .Y(men_men_n259_));
  NA2        u0210(.A(x5), .B(x0), .Y(men_men_n260_));
  NAi21      u0211(.An(men_men_n139_), .B(men_men_n260_), .Y(men_men_n261_));
  NA2        u0212(.A(men_men_n71_), .B(men_men_n50_), .Y(men_men_n262_));
  OAI210     u0213(.A0(men_men_n262_), .A1(men_men_n261_), .B0(men_men_n259_), .Y(men_men_n263_));
  NA3        u0214(.A(men_men_n263_), .B(men_men_n142_), .C(men_men_n257_), .Y(men_men_n264_));
  NA2        u0215(.A(x8), .B(men_men_n57_), .Y(men_men_n265_));
  NO2        u0216(.A(men_men_n265_), .B(x5), .Y(men_men_n266_));
  NO2        u0217(.A(men_men_n151_), .B(men_men_n71_), .Y(men_men_n267_));
  NA2        u0218(.A(x1), .B(x0), .Y(men_men_n268_));
  NA2        u0219(.A(men_men_n50_), .B(men_men_n59_), .Y(men_men_n269_));
  NA4        u0220(.A(men_men_n269_), .B(men_men_n268_), .C(men_men_n267_), .D(men_men_n266_), .Y(men_men_n270_));
  NA3        u0221(.A(men_men_n270_), .B(men_men_n264_), .C(men_men_n190_), .Y(men_men_n271_));
  NO2        u0222(.A(men_men_n107_), .B(x3), .Y(men_men_n272_));
  NO2        u0223(.A(men_men_n109_), .B(x0), .Y(men_men_n273_));
  NA2        u0224(.A(men_men_n273_), .B(men_men_n272_), .Y(men_men_n274_));
  NO2        u0225(.A(men_men_n55_), .B(x7), .Y(men_men_n275_));
  NA2        u0226(.A(men_men_n275_), .B(men_men_n140_), .Y(men_men_n276_));
  NO3        u0227(.A(x8), .B(men_men_n50_), .C(x0), .Y(men_men_n277_));
  NAi21      u0228(.An(x8), .B(x0), .Y(men_men_n278_));
  NAi21      u0229(.An(x1), .B(x3), .Y(men_men_n279_));
  NO2        u0230(.A(men_men_n279_), .B(men_men_n278_), .Y(men_men_n280_));
  NO2        u0231(.A(x2), .B(men_men_n53_), .Y(men_men_n281_));
  NOi21      u0232(.An(x5), .B(x6), .Y(men_men_n282_));
  NO2        u0233(.A(men_men_n57_), .B(x4), .Y(men_men_n283_));
  NO2        u0234(.A(men_men_n276_), .B(men_men_n274_), .Y(men_men_n284_));
  AOI210     u0235(.A0(men_men_n271_), .A1(men_men_n110_), .B0(men_men_n284_), .Y(men_men_n285_));
  NA3        u0236(.A(men_men_n285_), .B(men_men_n256_), .C(men_men_n238_), .Y(men_men_n286_));
  AOI210     u0237(.A0(men_men_n214_), .A1(men_men_n56_), .B0(men_men_n286_), .Y(men02));
  NO2        u0238(.A(x8), .B(men_men_n107_), .Y(men_men_n288_));
  XN2        u0239(.A(x7), .B(x3), .Y(men_men_n289_));
  INV        u0240(.A(men_men_n289_), .Y(men_men_n290_));
  NO2        u0241(.A(x2), .B(x0), .Y(men_men_n291_));
  NA2        u0242(.A(men_men_n291_), .B(men_men_n71_), .Y(men_men_n292_));
  NO2        u0243(.A(men_men_n57_), .B(x1), .Y(men_men_n293_));
  NA2        u0244(.A(men_men_n53_), .B(x0), .Y(men_men_n294_));
  NO2        u0245(.A(men_men_n279_), .B(x6), .Y(men_men_n295_));
  XO2        u0246(.A(x7), .B(x0), .Y(men_men_n296_));
  NO2        u0247(.A(men_men_n296_), .B(men_men_n291_), .Y(men_men_n297_));
  AN2        u0248(.A(x7), .B(x2), .Y(men_men_n298_));
  NA2        u0249(.A(men_men_n298_), .B(men_men_n50_), .Y(men_men_n299_));
  NAi21      u0250(.An(x8), .B(x6), .Y(men_men_n300_));
  NO2        u0251(.A(men_men_n107_), .B(men_men_n59_), .Y(men_men_n301_));
  NA2        u0252(.A(x7), .B(x3), .Y(men_men_n302_));
  NO2        u0253(.A(men_men_n302_), .B(x2), .Y(men_men_n303_));
  NA2        u0254(.A(x2), .B(x0), .Y(men_men_n304_));
  NA2        u0255(.A(men_men_n109_), .B(men_men_n59_), .Y(men_men_n305_));
  NA2        u0256(.A(men_men_n305_), .B(men_men_n304_), .Y(men_men_n306_));
  NAi21      u0257(.An(x7), .B(x1), .Y(men_men_n307_));
  NO2        u0258(.A(men_men_n307_), .B(x3), .Y(men_men_n308_));
  AOI220     u0259(.A0(men_men_n308_), .A1(men_men_n306_), .B0(men_men_n303_), .B1(men_men_n301_), .Y(men_men_n309_));
  NA2        u0260(.A(men_men_n281_), .B(men_men_n50_), .Y(men_men_n310_));
  NA3        u0261(.A(x7), .B(men_men_n107_), .C(x0), .Y(men_men_n311_));
  NA2        u0262(.A(men_men_n273_), .B(men_men_n53_), .Y(men_men_n312_));
  NA2        u0263(.A(men_men_n165_), .B(men_men_n57_), .Y(men_men_n313_));
  OA220      u0264(.A0(men_men_n313_), .A1(men_men_n312_), .B0(men_men_n311_), .B1(men_men_n310_), .Y(men_men_n314_));
  AOI210     u0265(.A0(men_men_n314_), .A1(men_men_n309_), .B0(men_men_n300_), .Y(men_men_n315_));
  INV        u0266(.A(men_men_n296_), .Y(men_men_n316_));
  NO2        u0267(.A(x7), .B(men_men_n71_), .Y(men_men_n317_));
  NA2        u0268(.A(men_men_n107_), .B(x3), .Y(men_men_n318_));
  NO2        u0269(.A(men_men_n318_), .B(men_men_n317_), .Y(men_men_n319_));
  NA2        u0270(.A(men_men_n319_), .B(men_men_n316_), .Y(men_men_n320_));
  NA2        u0271(.A(men_men_n50_), .B(x0), .Y(men_men_n321_));
  NO2        u0272(.A(men_men_n321_), .B(x7), .Y(men_men_n322_));
  NA2        u0273(.A(men_men_n322_), .B(men_men_n282_), .Y(men_men_n323_));
  NA2        u0274(.A(men_men_n170_), .B(x1), .Y(men_men_n324_));
  AOI210     u0275(.A0(men_men_n323_), .A1(men_men_n320_), .B0(men_men_n324_), .Y(men_men_n325_));
  NO2        u0276(.A(men_men_n57_), .B(men_men_n50_), .Y(men_men_n326_));
  NO2        u0277(.A(men_men_n55_), .B(men_men_n109_), .Y(men_men_n327_));
  NA3        u0278(.A(men_men_n327_), .B(men_men_n326_), .C(men_men_n59_), .Y(men_men_n328_));
  NO2        u0279(.A(men_men_n160_), .B(x6), .Y(men_men_n329_));
  NO2        u0280(.A(men_men_n103_), .B(men_men_n107_), .Y(men_men_n330_));
  NA2        u0281(.A(men_men_n57_), .B(men_men_n109_), .Y(men_men_n331_));
  NO2        u0282(.A(men_men_n331_), .B(men_men_n269_), .Y(men_men_n332_));
  OAI210     u0283(.A0(men_men_n330_), .A1(men_men_n329_), .B0(men_men_n332_), .Y(men_men_n333_));
  OAI210     u0284(.A0(men_men_n328_), .A1(men_men_n103_), .B0(men_men_n333_), .Y(men_men_n334_));
  NO3        u0285(.A(men_men_n334_), .B(men_men_n325_), .C(men_men_n315_), .Y(men_men_n335_));
  NO2        u0286(.A(men_men_n335_), .B(x4), .Y(men_men_n336_));
  NA2        u0287(.A(x8), .B(men_men_n71_), .Y(men_men_n337_));
  NO2        u0288(.A(x3), .B(men_men_n59_), .Y(men_men_n338_));
  NA3        u0289(.A(men_men_n338_), .B(men_men_n107_), .C(men_men_n53_), .Y(men_men_n339_));
  NO2        u0290(.A(x3), .B(x0), .Y(men_men_n340_));
  NAi21      u0291(.An(men_men_n340_), .B(men_men_n106_), .Y(men_men_n341_));
  NA2        u0292(.A(x5), .B(x2), .Y(men_men_n342_));
  NO2        u0293(.A(men_men_n342_), .B(men_men_n224_), .Y(men_men_n343_));
  AOI210     u0294(.A0(men_men_n343_), .A1(men_men_n341_), .B0(men_men_n245_), .Y(men_men_n344_));
  AO210      u0295(.A0(men_men_n344_), .A1(men_men_n339_), .B0(men_men_n337_), .Y(men_men_n345_));
  NO2        u0296(.A(men_men_n109_), .B(men_men_n53_), .Y(men_men_n346_));
  NA2        u0297(.A(men_men_n346_), .B(x3), .Y(men_men_n347_));
  NO2        u0298(.A(men_men_n55_), .B(x1), .Y(men_men_n348_));
  NA2        u0299(.A(men_men_n348_), .B(men_men_n109_), .Y(men_men_n349_));
  OAI210     u0300(.A0(men_men_n349_), .A1(men_men_n173_), .B0(men_men_n347_), .Y(men_men_n350_));
  NAi32      u0301(.An(x3), .Bn(x0), .C(x2), .Y(men_men_n351_));
  NO2        u0302(.A(men_men_n50_), .B(x2), .Y(men_men_n352_));
  NAi21      u0303(.An(x6), .B(x5), .Y(men_men_n353_));
  NO2        u0304(.A(x2), .B(men_men_n59_), .Y(men_men_n354_));
  NA2        u0305(.A(men_men_n350_), .B(men_men_n85_), .Y(men_men_n355_));
  AOI210     u0306(.A0(men_men_n355_), .A1(men_men_n345_), .B0(men_men_n75_), .Y(men_men_n356_));
  NA2        u0307(.A(men_men_n348_), .B(men_men_n56_), .Y(men_men_n357_));
  NO2        u0308(.A(men_men_n107_), .B(men_men_n50_), .Y(men_men_n358_));
  NO2        u0309(.A(men_men_n291_), .B(men_men_n221_), .Y(men_men_n359_));
  XO2        u0310(.A(x7), .B(x2), .Y(men_men_n360_));
  INV        u0311(.A(men_men_n360_), .Y(men_men_n361_));
  XO2        u0312(.A(x6), .B(x2), .Y(men_men_n362_));
  NA3        u0313(.A(men_men_n361_), .B(men_men_n359_), .C(men_men_n358_), .Y(men_men_n363_));
  NAi21      u0314(.An(x0), .B(x6), .Y(men_men_n364_));
  AOI210     u0315(.A0(men_men_n364_), .A1(men_men_n145_), .B0(men_men_n273_), .Y(men_men_n365_));
  XN2        u0316(.A(x7), .B(x5), .Y(men_men_n366_));
  NA2        u0317(.A(men_men_n366_), .B(men_men_n71_), .Y(men_men_n367_));
  NA2        u0318(.A(x7), .B(x5), .Y(men_men_n368_));
  AOI210     u0319(.A0(men_men_n368_), .A1(x6), .B0(men_men_n351_), .Y(men_men_n369_));
  AOI220     u0320(.A0(men_men_n369_), .A1(men_men_n367_), .B0(men_men_n365_), .B1(men_men_n319_), .Y(men_men_n370_));
  AOI210     u0321(.A0(men_men_n370_), .A1(men_men_n363_), .B0(men_men_n357_), .Y(men_men_n371_));
  NO2        u0322(.A(x8), .B(x6), .Y(men_men_n372_));
  NAi21      u0323(.An(men_men_n372_), .B(men_men_n233_), .Y(men_men_n373_));
  AOI210     u0324(.A0(men_men_n373_), .A1(men_men_n91_), .B0(x3), .Y(men_men_n374_));
  NA2        u0325(.A(men_men_n107_), .B(x2), .Y(men_men_n375_));
  NO2        u0326(.A(men_men_n375_), .B(men_men_n64_), .Y(men_men_n376_));
  NA2        u0327(.A(x1), .B(men_men_n59_), .Y(men_men_n377_));
  NO2        u0328(.A(men_men_n377_), .B(men_men_n233_), .Y(men_men_n378_));
  OAI210     u0329(.A0(men_men_n378_), .A1(men_men_n50_), .B0(men_men_n376_), .Y(men_men_n379_));
  NA2        u0330(.A(x4), .B(x2), .Y(men_men_n380_));
  NO2        u0331(.A(men_men_n380_), .B(men_men_n107_), .Y(men_men_n381_));
  NAi21      u0332(.An(x1), .B(x6), .Y(men_men_n382_));
  NA2        u0333(.A(men_men_n340_), .B(men_men_n275_), .Y(men_men_n383_));
  OAI220     u0334(.A0(men_men_n383_), .A1(men_men_n382_), .B0(men_men_n106_), .B1(men_men_n53_), .Y(men_men_n384_));
  NA2        u0335(.A(x8), .B(x2), .Y(men_men_n385_));
  NO2        u0336(.A(men_men_n385_), .B(men_men_n50_), .Y(men_men_n386_));
  INV        u0337(.A(men_men_n223_), .Y(men_men_n387_));
  NO2        u0338(.A(men_men_n387_), .B(men_men_n52_), .Y(men_men_n388_));
  AOI220     u0339(.A0(men_men_n388_), .A1(men_men_n386_), .B0(men_men_n384_), .B1(men_men_n381_), .Y(men_men_n389_));
  OAI210     u0340(.A0(men_men_n379_), .A1(men_men_n374_), .B0(men_men_n389_), .Y(men_men_n390_));
  NO4        u0341(.A(men_men_n390_), .B(men_men_n371_), .C(men_men_n356_), .D(men_men_n336_), .Y(men03));
  NAi21      u0342(.An(x2), .B(x0), .Y(men_men_n392_));
  NO3        u0343(.A(x8), .B(x6), .C(x4), .Y(men_men_n393_));
  INV        u0344(.A(men_men_n393_), .Y(men_men_n394_));
  NO2        u0345(.A(men_men_n394_), .B(men_men_n392_), .Y(men_men_n395_));
  NA2        u0346(.A(men_men_n395_), .B(men_men_n165_), .Y(men_men_n396_));
  NA2        u0347(.A(x3), .B(x2), .Y(men_men_n397_));
  NO2        u0348(.A(men_men_n162_), .B(x0), .Y(men_men_n398_));
  NA2        u0349(.A(x8), .B(x0), .Y(men_men_n399_));
  NO2        u0350(.A(men_men_n399_), .B(x6), .Y(men_men_n400_));
  AOI210     u0351(.A0(men_men_n400_), .A1(x5), .B0(men_men_n398_), .Y(men_men_n401_));
  NO2        u0352(.A(men_men_n401_), .B(men_men_n397_), .Y(men_men_n402_));
  NO2        u0353(.A(x5), .B(men_men_n59_), .Y(men_men_n403_));
  NO2        u0354(.A(x3), .B(x2), .Y(men_men_n404_));
  NA2        u0355(.A(men_men_n404_), .B(men_men_n403_), .Y(men_men_n405_));
  NO2        u0356(.A(men_men_n53_), .B(x0), .Y(men_men_n406_));
  NA2        u0357(.A(men_men_n406_), .B(x5), .Y(men_men_n407_));
  AOI210     u0358(.A0(men_men_n407_), .A1(men_men_n405_), .B0(men_men_n300_), .Y(men_men_n408_));
  NA2        u0359(.A(men_men_n259_), .B(men_men_n175_), .Y(men_men_n409_));
  NO2        u0360(.A(men_men_n50_), .B(men_men_n59_), .Y(men_men_n410_));
  NO2        u0361(.A(men_men_n71_), .B(x0), .Y(men_men_n411_));
  NO4        u0362(.A(men_men_n411_), .B(men_men_n410_), .C(x2), .D(men_men_n53_), .Y(men_men_n412_));
  AO210      u0363(.A0(men_men_n412_), .A1(men_men_n409_), .B0(men_men_n408_), .Y(men_men_n413_));
  OAI210     u0364(.A0(men_men_n413_), .A1(men_men_n402_), .B0(x4), .Y(men_men_n414_));
  NO2        u0365(.A(x4), .B(men_men_n53_), .Y(men_men_n415_));
  NA2        u0366(.A(men_men_n415_), .B(men_men_n59_), .Y(men_men_n416_));
  NO3        u0367(.A(men_men_n416_), .B(men_men_n233_), .C(x5), .Y(men_men_n417_));
  NA2        u0368(.A(x7), .B(men_men_n107_), .Y(men_men_n418_));
  NO3        u0369(.A(x5), .B(men_men_n53_), .C(x0), .Y(men_men_n419_));
  INV        u0370(.A(men_men_n419_), .Y(men_men_n420_));
  NO2        u0371(.A(x6), .B(men_men_n56_), .Y(men_men_n421_));
  NO2        u0372(.A(x8), .B(men_men_n50_), .Y(men_men_n422_));
  NA2        u0373(.A(men_men_n422_), .B(men_men_n421_), .Y(men_men_n423_));
  AOI210     u0374(.A0(men_men_n417_), .A1(x2), .B0(x7), .Y(men_men_n424_));
  AOI220     u0375(.A0(men_men_n424_), .A1(men_men_n414_), .B0(men_men_n396_), .B1(x7), .Y(men_men_n425_));
  NA2        u0376(.A(x7), .B(men_men_n53_), .Y(men_men_n426_));
  NO2        u0377(.A(men_men_n258_), .B(men_men_n109_), .Y(men_men_n427_));
  NO2        u0378(.A(men_men_n55_), .B(men_men_n59_), .Y(men_men_n428_));
  NO3        u0379(.A(men_men_n428_), .B(men_men_n427_), .C(men_men_n149_), .Y(men_men_n429_));
  AOI210     u0380(.A0(men_men_n209_), .A1(men_men_n100_), .B0(men_men_n429_), .Y(men_men_n430_));
  NO2        u0381(.A(x5), .B(x2), .Y(men_men_n431_));
  NO2        u0382(.A(x8), .B(x3), .Y(men_men_n432_));
  NA2        u0383(.A(men_men_n432_), .B(men_men_n431_), .Y(men_men_n433_));
  NO2        u0384(.A(men_men_n433_), .B(x6), .Y(men_men_n434_));
  NA2        u0385(.A(men_men_n208_), .B(x2), .Y(men_men_n435_));
  INV        u0386(.A(men_men_n434_), .Y(men_men_n436_));
  OAI210     u0387(.A0(men_men_n430_), .A1(men_men_n291_), .B0(men_men_n436_), .Y(men_men_n437_));
  NA2        u0388(.A(men_men_n437_), .B(x4), .Y(men_men_n438_));
  NA2        u0389(.A(men_men_n55_), .B(men_men_n59_), .Y(men_men_n439_));
  NO2        u0390(.A(men_men_n439_), .B(x5), .Y(men_men_n440_));
  NAi21      u0391(.An(x4), .B(x6), .Y(men_men_n441_));
  NO2        u0392(.A(men_men_n441_), .B(men_men_n51_), .Y(men_men_n442_));
  NO2        u0393(.A(men_men_n55_), .B(men_men_n71_), .Y(men_men_n443_));
  NO2        u0394(.A(men_men_n50_), .B(men_men_n109_), .Y(men_men_n444_));
  NO2        u0395(.A(men_men_n233_), .B(x0), .Y(men_men_n445_));
  NO2        u0396(.A(men_men_n353_), .B(x8), .Y(men_men_n446_));
  NO2        u0397(.A(men_men_n405_), .B(men_men_n443_), .Y(men_men_n447_));
  AOI220     u0398(.A0(men_men_n447_), .A1(men_men_n56_), .B0(men_men_n442_), .B1(men_men_n440_), .Y(men_men_n448_));
  AOI210     u0399(.A0(men_men_n448_), .A1(men_men_n438_), .B0(men_men_n426_), .Y(men_men_n449_));
  NA2        u0400(.A(men_men_n57_), .B(men_men_n53_), .Y(men_men_n450_));
  NO2        u0401(.A(men_men_n71_), .B(men_men_n56_), .Y(men_men_n451_));
  NA2        u0402(.A(men_men_n352_), .B(men_men_n59_), .Y(men_men_n452_));
  OAI220     u0403(.A0(men_men_n452_), .A1(men_men_n55_), .B0(men_men_n201_), .B1(men_men_n278_), .Y(men_men_n453_));
  NA2        u0404(.A(men_men_n453_), .B(men_men_n451_), .Y(men_men_n454_));
  NO3        u0405(.A(x6), .B(x4), .C(men_men_n50_), .Y(men_men_n455_));
  NA2        u0406(.A(men_men_n428_), .B(x5), .Y(men_men_n456_));
  NO2        u0407(.A(x8), .B(x5), .Y(men_men_n457_));
  NAi21      u0408(.An(men_men_n457_), .B(men_men_n175_), .Y(men_men_n458_));
  NO2        u0409(.A(men_men_n458_), .B(men_men_n305_), .Y(men_men_n459_));
  NA2        u0410(.A(men_men_n359_), .B(men_men_n77_), .Y(men_men_n460_));
  NOi21      u0411(.An(x3), .B(x4), .Y(men_men_n461_));
  NA2        u0412(.A(men_men_n55_), .B(men_men_n109_), .Y(men_men_n462_));
  NA2        u0413(.A(men_men_n462_), .B(men_men_n461_), .Y(men_men_n463_));
  NO2        u0414(.A(men_men_n149_), .B(men_men_n55_), .Y(men_men_n464_));
  NO3        u0415(.A(men_men_n56_), .B(x2), .C(x0), .Y(men_men_n465_));
  NO2        u0416(.A(men_men_n463_), .B(men_men_n460_), .Y(men_men_n466_));
  AOI210     u0417(.A0(men_men_n459_), .A1(men_men_n455_), .B0(men_men_n466_), .Y(men_men_n467_));
  AOI210     u0418(.A0(men_men_n467_), .A1(men_men_n454_), .B0(men_men_n450_), .Y(men_men_n468_));
  NA2        u0419(.A(x7), .B(x1), .Y(men_men_n469_));
  NO3        u0420(.A(x5), .B(x4), .C(x2), .Y(men_men_n470_));
  AN2        u0421(.A(men_men_n470_), .B(men_men_n372_), .Y(men_men_n471_));
  NO3        u0422(.A(men_men_n471_), .B(men_men_n464_), .C(men_men_n381_), .Y(men_men_n472_));
  OAI210     u0423(.A0(men_men_n372_), .A1(men_men_n84_), .B0(men_men_n340_), .Y(men_men_n473_));
  NO2        u0424(.A(men_men_n473_), .B(men_men_n472_), .Y(men_men_n474_));
  NO2        u0425(.A(x4), .B(men_men_n109_), .Y(men_men_n475_));
  NA2        u0426(.A(men_men_n475_), .B(x6), .Y(men_men_n476_));
  NA3        u0427(.A(men_men_n107_), .B(x4), .C(men_men_n109_), .Y(men_men_n477_));
  AOI210     u0428(.A0(men_men_n477_), .A1(men_men_n476_), .B0(men_men_n99_), .Y(men_men_n478_));
  NA2        u0429(.A(men_men_n461_), .B(men_men_n71_), .Y(men_men_n479_));
  NA2        u0430(.A(men_men_n170_), .B(men_men_n59_), .Y(men_men_n480_));
  NA2        u0431(.A(men_men_n444_), .B(x4), .Y(men_men_n481_));
  NO3        u0432(.A(men_men_n481_), .B(men_men_n372_), .C(men_men_n411_), .Y(men_men_n482_));
  NO3        u0433(.A(men_men_n482_), .B(men_men_n478_), .C(men_men_n474_), .Y(men_men_n483_));
  NA2        u0434(.A(x5), .B(x4), .Y(men_men_n484_));
  NO2        u0435(.A(men_men_n71_), .B(men_men_n53_), .Y(men_men_n485_));
  NO3        u0436(.A(x8), .B(x3), .C(x2), .Y(men_men_n486_));
  NA3        u0437(.A(men_men_n486_), .B(men_men_n485_), .C(men_men_n59_), .Y(men_men_n487_));
  NO3        u0438(.A(x6), .B(x5), .C(x2), .Y(men_men_n488_));
  NA3        u0439(.A(men_men_n488_), .B(men_men_n293_), .C(men_men_n78_), .Y(men_men_n489_));
  OAI210     u0440(.A0(men_men_n487_), .A1(men_men_n484_), .B0(men_men_n489_), .Y(men_men_n490_));
  NA2        u0441(.A(men_men_n71_), .B(x2), .Y(men_men_n491_));
  XO2        u0442(.A(x4), .B(x0), .Y(men_men_n492_));
  NA2        u0443(.A(men_men_n269_), .B(x5), .Y(men_men_n493_));
  NO2        u0444(.A(men_men_n56_), .B(men_men_n50_), .Y(men_men_n494_));
  NO2        u0445(.A(men_men_n494_), .B(men_men_n63_), .Y(men_men_n495_));
  NO4        u0446(.A(men_men_n495_), .B(men_men_n493_), .C(men_men_n492_), .D(men_men_n158_), .Y(men_men_n496_));
  NO2        u0447(.A(men_men_n496_), .B(men_men_n490_), .Y(men_men_n497_));
  OAI210     u0448(.A0(men_men_n483_), .A1(men_men_n469_), .B0(men_men_n497_), .Y(men_men_n498_));
  NO4        u0449(.A(men_men_n498_), .B(men_men_n468_), .C(men_men_n449_), .D(men_men_n425_), .Y(men04));
  NO2        u0450(.A(x7), .B(x2), .Y(men_men_n500_));
  NO2        u0451(.A(x3), .B(men_men_n53_), .Y(men_men_n501_));
  NO2        u0452(.A(men_men_n501_), .B(men_men_n151_), .Y(men_men_n502_));
  XN2        u0453(.A(x8), .B(x1), .Y(men_men_n503_));
  NO2        u0454(.A(men_men_n503_), .B(men_men_n149_), .Y(men_men_n504_));
  NA2        u0455(.A(men_men_n504_), .B(men_men_n502_), .Y(men_men_n505_));
  NA2        u0456(.A(x6), .B(x3), .Y(men_men_n506_));
  NO2        u0457(.A(men_men_n506_), .B(x5), .Y(men_men_n507_));
  NA2        u0458(.A(men_men_n71_), .B(x1), .Y(men_men_n508_));
  NO2        u0459(.A(men_men_n457_), .B(men_men_n258_), .Y(men_men_n509_));
  NO3        u0460(.A(men_men_n509_), .B(men_men_n432_), .C(men_men_n508_), .Y(men_men_n510_));
  AOI210     u0461(.A0(men_men_n507_), .A1(men_men_n348_), .B0(men_men_n510_), .Y(men_men_n511_));
  AOI210     u0462(.A0(men_men_n511_), .A1(men_men_n505_), .B0(x0), .Y(men_men_n512_));
  NOi21      u0463(.An(men_men_n175_), .B(men_men_n457_), .Y(men_men_n513_));
  NA2        u0464(.A(men_men_n108_), .B(x1), .Y(men_men_n514_));
  NO3        u0465(.A(men_men_n514_), .B(men_men_n513_), .C(men_men_n321_), .Y(men_men_n515_));
  OAI210     u0466(.A0(men_men_n515_), .A1(men_men_n512_), .B0(men_men_n500_), .Y(men_men_n516_));
  NA2        u0467(.A(men_men_n136_), .B(men_men_n244_), .Y(men_men_n517_));
  OR4        u0468(.A(men_men_n517_), .B(men_men_n373_), .C(men_men_n82_), .D(men_men_n54_), .Y(men_men_n518_));
  OR2        u0469(.A(x6), .B(x0), .Y(men_men_n519_));
  NO3        u0470(.A(men_men_n519_), .B(x3), .C(x1), .Y(men_men_n520_));
  AOI220     u0471(.A0(men_men_n520_), .A1(men_men_n107_), .B0(men_men_n282_), .B1(men_men_n277_), .Y(men_men_n521_));
  AOI210     u0472(.A0(men_men_n521_), .A1(men_men_n518_), .B0(men_men_n188_), .Y(men_men_n522_));
  NA2        u0473(.A(x7), .B(x2), .Y(men_men_n523_));
  INV        u0474(.A(men_men_n136_), .Y(men_men_n524_));
  OAI210     u0475(.A0(men_men_n174_), .A1(men_men_n524_), .B0(men_men_n82_), .Y(men_men_n525_));
  NO2        u0476(.A(men_men_n318_), .B(men_men_n55_), .Y(men_men_n526_));
  NO3        u0477(.A(x3), .B(x1), .C(x0), .Y(men_men_n527_));
  OR2        u0478(.A(x6), .B(x1), .Y(men_men_n528_));
  NA2        u0479(.A(men_men_n527_), .B(men_men_n464_), .Y(men_men_n529_));
  AOI210     u0480(.A0(men_men_n529_), .A1(men_men_n525_), .B0(men_men_n523_), .Y(men_men_n530_));
  NA2        u0481(.A(men_men_n71_), .B(x0), .Y(men_men_n531_));
  NOi31      u0482(.An(men_men_n343_), .B(men_men_n531_), .C(men_men_n265_), .Y(men_men_n532_));
  NO4        u0483(.A(men_men_n532_), .B(men_men_n530_), .C(men_men_n522_), .D(men_men_n56_), .Y(men_men_n533_));
  NA2        u0484(.A(men_men_n533_), .B(men_men_n516_), .Y(men_men_n534_));
  NA3        u0485(.A(x8), .B(x7), .C(x0), .Y(men_men_n535_));
  INV        u0486(.A(men_men_n535_), .Y(men_men_n536_));
  AOI210     u0487(.A0(men_men_n275_), .A1(men_men_n98_), .B0(men_men_n536_), .Y(men_men_n537_));
  NO2        u0488(.A(men_men_n537_), .B(men_men_n158_), .Y(men_men_n538_));
  NO2        u0489(.A(x8), .B(x0), .Y(men_men_n539_));
  NA2        u0490(.A(men_men_n538_), .B(men_men_n282_), .Y(men_men_n540_));
  NO2        u0491(.A(men_men_n71_), .B(men_men_n109_), .Y(men_men_n541_));
  NO2        u0492(.A(men_men_n368_), .B(x8), .Y(men_men_n542_));
  NO2        u0493(.A(men_men_n542_), .B(men_men_n266_), .Y(men_men_n543_));
  NO3        u0494(.A(men_men_n543_), .B(men_men_n377_), .C(men_men_n272_), .Y(men_men_n544_));
  OAI210     u0495(.A0(men_men_n457_), .A1(men_men_n326_), .B0(men_men_n247_), .Y(men_men_n545_));
  NO2        u0496(.A(men_men_n545_), .B(men_men_n289_), .Y(men_men_n546_));
  OAI210     u0497(.A0(men_men_n546_), .A1(men_men_n544_), .B0(men_men_n541_), .Y(men_men_n547_));
  NO2        u0498(.A(x8), .B(x2), .Y(men_men_n548_));
  NO2        u0499(.A(men_men_n224_), .B(men_men_n57_), .Y(men_men_n549_));
  NA3        u0500(.A(men_men_n549_), .B(men_men_n548_), .C(men_men_n341_), .Y(men_men_n550_));
  NO2        u0501(.A(men_men_n248_), .B(men_men_n136_), .Y(men_men_n551_));
  AOI210     u0502(.A0(men_men_n322_), .A1(men_men_n166_), .B0(men_men_n551_), .Y(men_men_n552_));
  AOI210     u0503(.A0(men_men_n552_), .A1(men_men_n550_), .B0(men_men_n108_), .Y(men_men_n553_));
  NA2        u0504(.A(men_men_n338_), .B(x2), .Y(men_men_n554_));
  NO2        u0505(.A(men_men_n57_), .B(men_men_n53_), .Y(men_men_n555_));
  NA2        u0506(.A(men_men_n109_), .B(men_men_n53_), .Y(men_men_n556_));
  NO2        u0507(.A(men_men_n556_), .B(x8), .Y(men_men_n557_));
  NA2        u0508(.A(x7), .B(men_men_n50_), .Y(men_men_n558_));
  NO2        u0509(.A(men_men_n185_), .B(men_men_n558_), .Y(men_men_n559_));
  AN2        u0510(.A(men_men_n559_), .B(men_men_n557_), .Y(men_men_n560_));
  NA2        u0511(.A(men_men_n403_), .B(men_men_n151_), .Y(men_men_n561_));
  NO2        u0512(.A(men_men_n71_), .B(x2), .Y(men_men_n562_));
  NA2        u0513(.A(men_men_n562_), .B(men_men_n275_), .Y(men_men_n563_));
  OAI210     u0514(.A0(men_men_n563_), .A1(men_men_n561_), .B0(men_men_n56_), .Y(men_men_n564_));
  NO3        u0515(.A(men_men_n564_), .B(men_men_n560_), .C(men_men_n553_), .Y(men_men_n565_));
  NA3        u0516(.A(men_men_n565_), .B(men_men_n547_), .C(men_men_n540_), .Y(men_men_n566_));
  NA2        u0517(.A(men_men_n53_), .B(men_men_n59_), .Y(men_men_n567_));
  NOi21      u0518(.An(x2), .B(x7), .Y(men_men_n568_));
  NO2        u0519(.A(x6), .B(x3), .Y(men_men_n569_));
  NA2        u0520(.A(men_men_n569_), .B(men_men_n568_), .Y(men_men_n570_));
  NO2        u0521(.A(x6), .B(men_men_n59_), .Y(men_men_n571_));
  NO3        u0522(.A(men_men_n57_), .B(x2), .C(x1), .Y(men_men_n572_));
  NO3        u0523(.A(men_men_n57_), .B(x2), .C(x0), .Y(men_men_n573_));
  AOI220     u0524(.A0(men_men_n573_), .A1(men_men_n227_), .B0(men_men_n572_), .B1(men_men_n571_), .Y(men_men_n574_));
  INV        u0525(.A(men_men_n574_), .Y(men_men_n575_));
  NO2        u0526(.A(men_men_n100_), .B(men_men_n53_), .Y(men_men_n576_));
  NA2        u0527(.A(men_men_n222_), .B(men_men_n57_), .Y(men_men_n577_));
  OAI210     u0528(.A0(men_men_n576_), .A1(men_men_n446_), .B0(men_men_n577_), .Y(men_men_n578_));
  NO3        u0529(.A(men_men_n578_), .B(men_men_n481_), .C(men_men_n59_), .Y(men_men_n579_));
  AO210      u0530(.A0(men_men_n575_), .A1(men_men_n457_), .B0(men_men_n579_), .Y(men_men_n580_));
  AOI210     u0531(.A0(men_men_n566_), .A1(men_men_n534_), .B0(men_men_n580_), .Y(men05));
  AOI210     u0532(.A0(men_men_n165_), .A1(men_men_n55_), .B0(men_men_n494_), .Y(men_men_n582_));
  OR2        u0533(.A(men_men_n582_), .B(men_men_n57_), .Y(men_men_n583_));
  NO2        u0534(.A(x7), .B(men_men_n107_), .Y(men_men_n584_));
  NO2        u0535(.A(x8), .B(men_men_n56_), .Y(men_men_n585_));
  NA2        u0536(.A(x5), .B(men_men_n56_), .Y(men_men_n586_));
  NO2        u0537(.A(men_men_n586_), .B(men_men_n558_), .Y(men_men_n587_));
  AOI210     u0538(.A0(men_men_n585_), .A1(men_men_n584_), .B0(men_men_n587_), .Y(men_men_n588_));
  AOI210     u0539(.A0(men_men_n588_), .A1(men_men_n583_), .B0(men_men_n109_), .Y(men_men_n589_));
  NO2        u0540(.A(x7), .B(x4), .Y(men_men_n590_));
  NO2        u0541(.A(men_men_n64_), .B(men_men_n55_), .Y(men_men_n591_));
  NO2        u0542(.A(men_men_n201_), .B(x5), .Y(men_men_n592_));
  NA2        u0543(.A(men_men_n107_), .B(men_men_n109_), .Y(men_men_n593_));
  NO2        u0544(.A(men_men_n593_), .B(men_men_n218_), .Y(men_men_n594_));
  AO220      u0545(.A0(men_men_n594_), .A1(men_men_n590_), .B0(men_men_n592_), .B1(men_men_n591_), .Y(men_men_n595_));
  OAI210     u0546(.A0(men_men_n595_), .A1(men_men_n589_), .B0(men_men_n485_), .Y(men_men_n596_));
  NO2        u0547(.A(x6), .B(men_men_n50_), .Y(men_men_n597_));
  NA2        u0548(.A(men_men_n55_), .B(x4), .Y(men_men_n598_));
  NO2        u0549(.A(men_men_n107_), .B(men_men_n109_), .Y(men_men_n599_));
  NA2        u0550(.A(men_men_n599_), .B(x7), .Y(men_men_n600_));
  NA2        u0551(.A(men_men_n431_), .B(men_men_n257_), .Y(men_men_n601_));
  AOI210     u0552(.A0(men_men_n601_), .A1(men_men_n600_), .B0(men_men_n598_), .Y(men_men_n602_));
  NA2        u0553(.A(men_men_n107_), .B(x4), .Y(men_men_n603_));
  XO2        u0554(.A(x7), .B(x5), .Y(men_men_n604_));
  NO2        u0555(.A(men_men_n604_), .B(men_men_n53_), .Y(men_men_n605_));
  NA3        u0556(.A(men_men_n605_), .B(men_men_n603_), .C(men_men_n327_), .Y(men_men_n606_));
  NO2        u0557(.A(men_men_n107_), .B(x2), .Y(men_men_n607_));
  NO2        u0558(.A(men_men_n75_), .B(men_men_n55_), .Y(men_men_n608_));
  NA2        u0559(.A(men_men_n608_), .B(men_men_n607_), .Y(men_men_n609_));
  NA2        u0560(.A(men_men_n609_), .B(men_men_n606_), .Y(men_men_n610_));
  OAI210     u0561(.A0(men_men_n610_), .A1(men_men_n602_), .B0(men_men_n597_), .Y(men_men_n611_));
  NO2        u0562(.A(men_men_n71_), .B(men_men_n50_), .Y(men_men_n612_));
  NO2        u0563(.A(men_men_n195_), .B(x4), .Y(men_men_n613_));
  NO2        u0564(.A(x5), .B(men_men_n56_), .Y(men_men_n614_));
  XO2        u0565(.A(x5), .B(x2), .Y(men_men_n615_));
  NO3        u0566(.A(x8), .B(x7), .C(men_men_n109_), .Y(men_men_n616_));
  AO220      u0567(.A0(men_men_n616_), .A1(men_men_n614_), .B0(men_men_n615_), .B1(men_men_n613_), .Y(men_men_n617_));
  NA3        u0568(.A(men_men_n617_), .B(men_men_n612_), .C(men_men_n53_), .Y(men_men_n618_));
  NA2        u0569(.A(men_men_n272_), .B(men_men_n568_), .Y(men_men_n619_));
  NOi21      u0570(.An(x4), .B(x1), .Y(men_men_n620_));
  NA2        u0571(.A(men_men_n620_), .B(men_men_n63_), .Y(men_men_n621_));
  NA2        u0572(.A(x4), .B(x1), .Y(men_men_n622_));
  NO2        u0573(.A(men_men_n622_), .B(men_men_n50_), .Y(men_men_n623_));
  AOI210     u0574(.A0(men_men_n623_), .A1(men_men_n599_), .B0(men_men_n59_), .Y(men_men_n624_));
  OA210      u0575(.A0(men_men_n621_), .A1(men_men_n619_), .B0(men_men_n624_), .Y(men_men_n625_));
  NA4        u0576(.A(men_men_n625_), .B(men_men_n618_), .C(men_men_n611_), .D(men_men_n596_), .Y(men_men_n626_));
  NA2        u0577(.A(men_men_n612_), .B(men_men_n56_), .Y(men_men_n627_));
  NA2        u0578(.A(men_men_n548_), .B(men_men_n584_), .Y(men_men_n628_));
  NO2        u0579(.A(men_men_n628_), .B(men_men_n627_), .Y(men_men_n629_));
  NA2        u0580(.A(men_men_n275_), .B(men_men_n122_), .Y(men_men_n630_));
  OAI210     u0581(.A0(men_men_n630_), .A1(men_men_n167_), .B0(men_men_n59_), .Y(men_men_n631_));
  NA2        u0582(.A(men_men_n57_), .B(x6), .Y(men_men_n632_));
  AOI210     u0583(.A0(men_men_n632_), .A1(x3), .B0(men_men_n90_), .Y(men_men_n633_));
  NA2        u0584(.A(men_men_n614_), .B(men_men_n157_), .Y(men_men_n634_));
  NO3        u0585(.A(men_men_n634_), .B(men_men_n633_), .C(men_men_n422_), .Y(men_men_n635_));
  NA2        u0586(.A(men_men_n283_), .B(men_men_n71_), .Y(men_men_n636_));
  NO2        u0587(.A(men_men_n385_), .B(x3), .Y(men_men_n637_));
  NA2        u0588(.A(men_men_n637_), .B(men_men_n241_), .Y(men_men_n638_));
  NO2        u0589(.A(men_men_n422_), .B(men_men_n613_), .Y(men_men_n639_));
  NO2        u0590(.A(men_men_n461_), .B(men_men_n107_), .Y(men_men_n640_));
  NO2        u0591(.A(men_men_n556_), .B(x6), .Y(men_men_n641_));
  NA2        u0592(.A(men_men_n641_), .B(men_men_n640_), .Y(men_men_n642_));
  OAI220     u0593(.A0(men_men_n642_), .A1(men_men_n639_), .B0(men_men_n638_), .B1(men_men_n636_), .Y(men_men_n643_));
  NO4        u0594(.A(men_men_n643_), .B(men_men_n635_), .C(men_men_n631_), .D(men_men_n629_), .Y(men_men_n644_));
  NA2        u0595(.A(men_men_n57_), .B(x5), .Y(men_men_n645_));
  NO2        u0596(.A(men_men_n645_), .B(x1), .Y(men_men_n646_));
  NA2        u0597(.A(x8), .B(men_men_n56_), .Y(men_men_n647_));
  NO2        u0598(.A(men_men_n647_), .B(men_men_n131_), .Y(men_men_n648_));
  NA2        u0599(.A(x8), .B(x4), .Y(men_men_n649_));
  NO2        u0600(.A(x8), .B(x4), .Y(men_men_n650_));
  NAi21      u0601(.An(men_men_n650_), .B(men_men_n649_), .Y(men_men_n651_));
  NAi21      u0602(.An(men_men_n548_), .B(men_men_n385_), .Y(men_men_n652_));
  NO4        u0603(.A(men_men_n652_), .B(men_men_n651_), .C(men_men_n422_), .D(men_men_n71_), .Y(men_men_n653_));
  OAI210     u0604(.A0(men_men_n653_), .A1(men_men_n648_), .B0(men_men_n646_), .Y(men_men_n654_));
  NO3        u0605(.A(x8), .B(men_men_n107_), .C(x4), .Y(men_men_n655_));
  INV        u0606(.A(men_men_n655_), .Y(men_men_n656_));
  NO2        u0607(.A(men_men_n656_), .B(men_men_n109_), .Y(men_men_n657_));
  NO2        u0608(.A(x5), .B(x4), .Y(men_men_n658_));
  NA3        u0609(.A(men_men_n658_), .B(men_men_n63_), .C(men_men_n109_), .Y(men_men_n659_));
  NO2        u0610(.A(x6), .B(men_men_n109_), .Y(men_men_n660_));
  NA2        u0611(.A(men_men_n647_), .B(men_men_n660_), .Y(men_men_n661_));
  OAI210     u0612(.A0(men_men_n661_), .A1(men_men_n513_), .B0(men_men_n659_), .Y(men_men_n662_));
  OAI210     u0613(.A0(men_men_n662_), .A1(men_men_n657_), .B0(men_men_n308_), .Y(men_men_n663_));
  NA3        u0614(.A(men_men_n663_), .B(men_men_n654_), .C(men_men_n644_), .Y(men_men_n664_));
  OR2        u0615(.A(x4), .B(x1), .Y(men_men_n665_));
  NO2        u0616(.A(men_men_n665_), .B(x3), .Y(men_men_n666_));
  NA2        u0617(.A(men_men_n55_), .B(x2), .Y(men_men_n667_));
  NO3        u0618(.A(men_men_n366_), .B(men_men_n667_), .C(x6), .Y(men_men_n668_));
  AOI220     u0619(.A0(men_men_n668_), .A1(men_men_n666_), .B0(men_men_n664_), .B1(men_men_n626_), .Y(men06));
  NA2        u0620(.A(men_men_n56_), .B(x3), .Y(men_men_n670_));
  NA2        u0621(.A(x6), .B(men_men_n109_), .Y(men_men_n671_));
  NA2        u0622(.A(men_men_n671_), .B(men_men_n55_), .Y(men_men_n672_));
  NA2        u0623(.A(x5), .B(men_men_n59_), .Y(men_men_n673_));
  NO2        u0624(.A(men_men_n673_), .B(men_men_n117_), .Y(men_men_n674_));
  NA3        u0625(.A(men_men_n674_), .B(men_men_n672_), .C(men_men_n491_), .Y(men_men_n675_));
  NO2        u0626(.A(men_men_n385_), .B(x0), .Y(men_men_n676_));
  NA2        u0627(.A(men_men_n337_), .B(x2), .Y(men_men_n677_));
  NOi21      u0628(.An(x6), .B(x8), .Y(men_men_n678_));
  NO2        u0629(.A(men_men_n678_), .B(x2), .Y(men_men_n679_));
  NO3        u0630(.A(men_men_n679_), .B(men_men_n70_), .C(men_men_n59_), .Y(men_men_n680_));
  AOI220     u0631(.A0(men_men_n680_), .A1(men_men_n677_), .B0(men_men_n676_), .B1(men_men_n329_), .Y(men_men_n681_));
  AOI210     u0632(.A0(men_men_n681_), .A1(men_men_n675_), .B0(men_men_n670_), .Y(men_men_n682_));
  NA2        u0633(.A(men_men_n56_), .B(men_men_n50_), .Y(men_men_n683_));
  NA2        u0634(.A(men_men_n364_), .B(men_men_n353_), .Y(men_men_n684_));
  NO2        u0635(.A(men_men_n71_), .B(men_men_n107_), .Y(men_men_n685_));
  NO2        u0636(.A(men_men_n53_), .B(men_men_n59_), .Y(men_men_n686_));
  NO4        u0637(.A(men_men_n686_), .B(men_men_n667_), .C(men_men_n685_), .D(men_men_n485_), .Y(men_men_n687_));
  AOI220     u0638(.A0(men_men_n687_), .A1(men_men_n684_), .B0(men_men_n419_), .B1(men_men_n63_), .Y(men_men_n688_));
  NO2        u0639(.A(men_men_n688_), .B(men_men_n683_), .Y(men_men_n689_));
  NO2        u0640(.A(men_men_n54_), .B(x0), .Y(men_men_n690_));
  NA2        u0641(.A(x4), .B(x3), .Y(men_men_n691_));
  NA2        u0642(.A(x3), .B(men_men_n690_), .Y(men_men_n692_));
  NO2        u0643(.A(men_men_n103_), .B(men_men_n56_), .Y(men_men_n693_));
  NA3        u0644(.A(men_men_n693_), .B(men_men_n258_), .C(men_men_n403_), .Y(men_men_n694_));
  AOI210     u0645(.A0(men_men_n694_), .A1(men_men_n692_), .B0(x2), .Y(men_men_n695_));
  INV        u0646(.A(men_men_n381_), .Y(men_men_n696_));
  NO2        u0647(.A(men_men_n406_), .B(x8), .Y(men_men_n697_));
  NO2        u0648(.A(men_men_n259_), .B(men_men_n508_), .Y(men_men_n698_));
  AOI210     u0649(.A0(men_men_n697_), .A1(men_men_n267_), .B0(men_men_n698_), .Y(men_men_n699_));
  NO2        u0650(.A(x5), .B(x3), .Y(men_men_n700_));
  NA3        u0651(.A(men_men_n539_), .B(men_men_n700_), .C(x1), .Y(men_men_n701_));
  NA2        u0652(.A(men_men_n585_), .B(men_men_n541_), .Y(men_men_n702_));
  OA220      u0653(.A0(men_men_n702_), .A1(men_men_n561_), .B0(men_men_n701_), .B1(men_men_n491_), .Y(men_men_n703_));
  OAI210     u0654(.A0(men_men_n699_), .A1(men_men_n696_), .B0(men_men_n703_), .Y(men_men_n704_));
  OR4        u0655(.A(men_men_n704_), .B(men_men_n695_), .C(men_men_n689_), .D(men_men_n682_), .Y(men_men_n705_));
  NA2        u0656(.A(x7), .B(men_men_n56_), .Y(men_men_n706_));
  NO2        u0657(.A(men_men_n599_), .B(men_men_n59_), .Y(men_men_n707_));
  NA2        u0658(.A(men_men_n707_), .B(men_men_n612_), .Y(men_men_n708_));
  NO2        u0659(.A(men_men_n173_), .B(x6), .Y(men_men_n709_));
  NA2        u0660(.A(men_men_n709_), .B(men_men_n291_), .Y(men_men_n710_));
  AOI210     u0661(.A0(men_men_n710_), .A1(men_men_n708_), .B0(men_men_n706_), .Y(men_men_n711_));
  AN2        u0662(.A(men_men_n465_), .B(men_men_n319_), .Y(men_men_n712_));
  OAI210     u0663(.A0(men_men_n712_), .A1(men_men_n711_), .B0(men_men_n348_), .Y(men_men_n713_));
  NO2        u0664(.A(men_men_n304_), .B(men_men_n107_), .Y(men_men_n714_));
  NO2        u0665(.A(men_men_n56_), .B(x3), .Y(men_men_n715_));
  NA2        u0666(.A(men_men_n715_), .B(men_men_n71_), .Y(men_men_n716_));
  NO2        u0667(.A(men_men_n716_), .B(men_men_n253_), .Y(men_men_n717_));
  NO2        u0668(.A(men_men_n71_), .B(x3), .Y(men_men_n718_));
  NA3        u0669(.A(men_men_n718_), .B(men_men_n555_), .C(men_men_n56_), .Y(men_men_n719_));
  NO2        u0670(.A(men_men_n57_), .B(x6), .Y(men_men_n720_));
  NA2        u0671(.A(men_men_n184_), .B(men_men_n720_), .Y(men_men_n721_));
  NA3        u0672(.A(men_men_n585_), .B(men_men_n326_), .C(men_men_n71_), .Y(men_men_n722_));
  NA3        u0673(.A(men_men_n722_), .B(men_men_n721_), .C(men_men_n719_), .Y(men_men_n723_));
  OR3        u0674(.A(men_men_n723_), .B(men_men_n717_), .C(men_men_n623_), .Y(men_men_n724_));
  NA2        u0675(.A(men_men_n724_), .B(men_men_n714_), .Y(men_men_n725_));
  NA2        u0676(.A(men_men_n690_), .B(men_men_n612_), .Y(men_men_n726_));
  NA4        u0677(.A(men_men_n268_), .B(men_men_n569_), .C(men_men_n222_), .D(men_men_n260_), .Y(men_men_n727_));
  NA2        u0678(.A(men_men_n475_), .B(men_men_n67_), .Y(men_men_n728_));
  AOI210     u0679(.A0(men_men_n727_), .A1(men_men_n726_), .B0(men_men_n728_), .Y(men_men_n729_));
  NA2        u0680(.A(x7), .B(x6), .Y(men_men_n730_));
  NA3        u0681(.A(x2), .B(x1), .C(x0), .Y(men_men_n731_));
  NO3        u0682(.A(men_men_n731_), .B(men_men_n730_), .C(men_men_n582_), .Y(men_men_n732_));
  NA2        u0683(.A(men_men_n486_), .B(men_men_n150_), .Y(men_men_n733_));
  NO2        u0684(.A(x5), .B(x1), .Y(men_men_n734_));
  NA2        u0685(.A(men_men_n734_), .B(men_men_n720_), .Y(men_men_n735_));
  NA2        u0686(.A(x4), .B(x0), .Y(men_men_n736_));
  NO3        u0687(.A(men_men_n57_), .B(x6), .C(x2), .Y(men_men_n737_));
  NA2        u0688(.A(men_men_n737_), .B(men_men_n226_), .Y(men_men_n738_));
  OAI220     u0689(.A0(men_men_n738_), .A1(men_men_n736_), .B0(men_men_n735_), .B1(men_men_n733_), .Y(men_men_n739_));
  NO3        u0690(.A(men_men_n739_), .B(men_men_n732_), .C(men_men_n729_), .Y(men_men_n740_));
  NA3        u0691(.A(men_men_n740_), .B(men_men_n725_), .C(men_men_n713_), .Y(men_men_n741_));
  AOI210     u0692(.A0(men_men_n705_), .A1(men_men_n57_), .B0(men_men_n741_), .Y(men07));
  NA2        u0693(.A(men_men_n107_), .B(men_men_n59_), .Y(men_men_n743_));
  NOi21      u0694(.An(men_men_n730_), .B(men_men_n115_), .Y(men_men_n744_));
  NO4        u0695(.A(men_men_n744_), .B(men_men_n612_), .C(men_men_n253_), .D(men_men_n743_), .Y(men_men_n745_));
  NO3        u0696(.A(men_men_n57_), .B(x5), .C(x1), .Y(men_men_n746_));
  NA2        u0697(.A(men_men_n746_), .B(men_men_n372_), .Y(men_men_n747_));
  NO2        u0698(.A(men_men_n57_), .B(men_men_n71_), .Y(men_men_n748_));
  NO2        u0699(.A(men_men_n156_), .B(men_men_n108_), .Y(men_men_n749_));
  AOI210     u0700(.A0(men_men_n748_), .A1(men_men_n91_), .B0(men_men_n749_), .Y(men_men_n750_));
  OAI220     u0701(.A0(men_men_n750_), .A1(men_men_n136_), .B0(men_men_n747_), .B1(men_men_n321_), .Y(men_men_n751_));
  OAI210     u0702(.A0(men_men_n751_), .A1(men_men_n745_), .B0(x2), .Y(men_men_n752_));
  NAi21      u0703(.An(men_men_n157_), .B(men_men_n158_), .Y(men_men_n753_));
  NO3        u0704(.A(men_men_n55_), .B(x3), .C(x1), .Y(men_men_n754_));
  NO2        u0705(.A(men_men_n501_), .B(x2), .Y(men_men_n755_));
  AOI210     u0706(.A0(men_men_n755_), .A1(men_men_n503_), .B0(men_men_n754_), .Y(men_men_n756_));
  NO2        u0707(.A(men_men_n756_), .B(men_men_n632_), .Y(men_men_n757_));
  NO2        u0708(.A(x8), .B(men_men_n53_), .Y(men_men_n758_));
  NA2        u0709(.A(men_men_n758_), .B(men_men_n59_), .Y(men_men_n759_));
  NA2        u0710(.A(men_men_n354_), .B(men_men_n348_), .Y(men_men_n760_));
  NO2        u0711(.A(x7), .B(x3), .Y(men_men_n761_));
  NA2        u0712(.A(men_men_n761_), .B(men_men_n100_), .Y(men_men_n762_));
  AOI210     u0713(.A0(men_men_n760_), .A1(men_men_n759_), .B0(men_men_n762_), .Y(men_men_n763_));
  AOI210     u0714(.A0(men_men_n757_), .A1(men_men_n252_), .B0(men_men_n763_), .Y(men_men_n764_));
  AOI210     u0715(.A0(men_men_n764_), .A1(men_men_n752_), .B0(x4), .Y(men_men_n765_));
  NA3        u0716(.A(men_men_n734_), .B(men_men_n317_), .C(men_men_n55_), .Y(men_men_n766_));
  AOI210     u0717(.A0(men_men_n766_), .A1(men_men_n578_), .B0(men_men_n109_), .Y(men_men_n767_));
  XO2        u0718(.A(x5), .B(x1), .Y(men_men_n768_));
  NO3        u0719(.A(men_men_n768_), .B(men_men_n210_), .C(men_men_n55_), .Y(men_men_n769_));
  OAI210     u0720(.A0(men_men_n769_), .A1(men_men_n767_), .B0(men_men_n410_), .Y(men_men_n770_));
  NO3        u0721(.A(men_men_n50_), .B(x2), .C(x0), .Y(men_men_n771_));
  NO2        u0722(.A(men_men_n307_), .B(men_men_n107_), .Y(men_men_n772_));
  NA2        u0723(.A(x6), .B(x0), .Y(men_men_n773_));
  NO2        u0724(.A(men_men_n667_), .B(men_men_n773_), .Y(men_men_n774_));
  NO2        u0725(.A(men_men_n768_), .B(men_men_n678_), .Y(men_men_n775_));
  OAI210     u0726(.A0(men_men_n734_), .A1(men_men_n63_), .B0(men_men_n57_), .Y(men_men_n776_));
  OAI210     u0727(.A0(men_men_n776_), .A1(men_men_n775_), .B0(men_men_n747_), .Y(men_men_n777_));
  AOI220     u0728(.A0(men_men_n777_), .A1(men_men_n771_), .B0(men_men_n774_), .B1(men_men_n772_), .Y(men_men_n778_));
  AOI210     u0729(.A0(men_men_n778_), .A1(men_men_n770_), .B0(men_men_n56_), .Y(men_men_n779_));
  NOi21      u0730(.An(men_men_n233_), .B(men_men_n372_), .Y(men_men_n780_));
  NO3        u0731(.A(men_men_n780_), .B(men_men_n242_), .C(men_men_n67_), .Y(men_men_n781_));
  NO2        u0732(.A(men_men_n193_), .B(men_men_n71_), .Y(men_men_n782_));
  NO2        u0733(.A(men_men_n307_), .B(x6), .Y(men_men_n783_));
  AO220      u0734(.A0(men_men_n783_), .A1(men_men_n327_), .B0(men_men_n782_), .B1(men_men_n542_), .Y(men_men_n784_));
  OAI210     u0735(.A0(men_men_n784_), .A1(men_men_n781_), .B0(men_men_n59_), .Y(men_men_n785_));
  NA2        u0736(.A(men_men_n91_), .B(men_men_n71_), .Y(men_men_n786_));
  NO2        u0737(.A(men_men_n786_), .B(men_men_n628_), .Y(men_men_n787_));
  NAi21      u0738(.An(x8), .B(x7), .Y(men_men_n788_));
  NA2        u0739(.A(men_men_n780_), .B(men_men_n788_), .Y(men_men_n789_));
  NA2        u0740(.A(men_men_n403_), .B(men_men_n109_), .Y(men_men_n790_));
  NO2        u0741(.A(men_men_n678_), .B(x1), .Y(men_men_n791_));
  NO3        u0742(.A(men_men_n791_), .B(men_men_n790_), .C(men_men_n555_), .Y(men_men_n792_));
  AOI210     u0743(.A0(men_men_n792_), .A1(men_men_n789_), .B0(men_men_n787_), .Y(men_men_n793_));
  AOI210     u0744(.A0(men_men_n793_), .A1(men_men_n785_), .B0(men_men_n143_), .Y(men_men_n794_));
  NO2        u0745(.A(x8), .B(x7), .Y(men_men_n795_));
  NO2        u0746(.A(x8), .B(men_men_n109_), .Y(men_men_n796_));
  AOI220     u0747(.A0(men_men_n326_), .A1(men_men_n348_), .B0(men_men_n796_), .B1(men_men_n257_), .Y(men_men_n797_));
  NO2        u0748(.A(men_men_n71_), .B(x4), .Y(men_men_n798_));
  NA2        u0749(.A(men_men_n798_), .B(men_men_n301_), .Y(men_men_n799_));
  NO2        u0750(.A(men_men_n797_), .B(men_men_n799_), .Y(men_men_n800_));
  NO4        u0751(.A(men_men_n800_), .B(men_men_n794_), .C(men_men_n779_), .D(men_men_n765_), .Y(men08));
  NA2        u0752(.A(men_men_n50_), .B(x1), .Y(men_men_n802_));
  XN2        u0753(.A(x5), .B(x4), .Y(men_men_n803_));
  INV        u0754(.A(men_men_n803_), .Y(men_men_n804_));
  AOI220     u0755(.A0(men_men_n804_), .A1(men_men_n354_), .B0(men_men_n139_), .B1(men_men_n56_), .Y(men_men_n805_));
  NO2        u0756(.A(men_men_n244_), .B(men_men_n107_), .Y(men_men_n806_));
  AOI210     u0757(.A0(men_men_n806_), .A1(men_men_n281_), .B0(men_men_n194_), .Y(men_men_n807_));
  OAI220     u0758(.A0(men_men_n807_), .A1(x4), .B0(men_men_n805_), .B1(men_men_n802_), .Y(men_men_n808_));
  NA2        u0759(.A(men_men_n808_), .B(men_men_n275_), .Y(men_men_n809_));
  AOI210     u0760(.A0(men_men_n274_), .A1(men_men_n790_), .B0(men_men_n598_), .Y(men_men_n810_));
  NA2        u0761(.A(men_men_n593_), .B(men_men_n173_), .Y(men_men_n811_));
  OAI220     u0762(.A0(men_men_n811_), .A1(men_men_n647_), .B0(men_men_n477_), .B1(men_men_n50_), .Y(men_men_n812_));
  AO210      u0763(.A0(men_men_n812_), .A1(men_men_n341_), .B0(men_men_n810_), .Y(men_men_n813_));
  NA2        u0764(.A(men_men_n281_), .B(men_men_n150_), .Y(men_men_n814_));
  NA2        u0765(.A(men_men_n143_), .B(x7), .Y(men_men_n815_));
  OR2        u0766(.A(men_men_n731_), .B(men_men_n461_), .Y(men_men_n816_));
  OAI220     u0767(.A0(men_men_n816_), .A1(men_men_n815_), .B0(men_men_n814_), .B1(men_men_n207_), .Y(men_men_n817_));
  AOI210     u0768(.A0(men_men_n813_), .A1(men_men_n293_), .B0(men_men_n817_), .Y(men_men_n818_));
  AOI210     u0769(.A0(men_men_n818_), .A1(men_men_n809_), .B0(men_men_n71_), .Y(men_men_n819_));
  NO2        u0770(.A(men_men_n795_), .B(men_men_n109_), .Y(men_men_n820_));
  NA2        u0771(.A(men_men_n820_), .B(men_men_n195_), .Y(men_men_n821_));
  OAI210     u0772(.A0(men_men_n406_), .A1(men_men_n301_), .B0(men_men_n341_), .Y(men_men_n822_));
  NA2        u0773(.A(men_men_n431_), .B(men_men_n235_), .Y(men_men_n823_));
  NA2        u0774(.A(men_men_n697_), .B(men_men_n106_), .Y(men_men_n824_));
  OAI220     u0775(.A0(men_men_n824_), .A1(men_men_n823_), .B0(men_men_n822_), .B1(men_men_n821_), .Y(men_men_n825_));
  NA2        u0776(.A(men_men_n825_), .B(men_men_n289_), .Y(men_men_n826_));
  NA2        u0777(.A(men_men_n331_), .B(men_men_n53_), .Y(men_men_n827_));
  NO3        u0778(.A(men_men_n406_), .B(men_men_n136_), .C(men_men_n68_), .Y(men_men_n828_));
  NO2        u0779(.A(men_men_n686_), .B(men_men_n247_), .Y(men_men_n829_));
  NO3        u0780(.A(men_men_n549_), .B(men_men_n462_), .C(men_men_n98_), .Y(men_men_n830_));
  AO220      u0781(.A0(men_men_n830_), .A1(men_men_n829_), .B0(men_men_n828_), .B1(men_men_n827_), .Y(men_men_n831_));
  NA2        u0782(.A(x7), .B(men_men_n59_), .Y(men_men_n832_));
  NO3        u0783(.A(men_men_n310_), .B(men_men_n832_), .C(men_men_n288_), .Y(men_men_n833_));
  AOI210     u0784(.A0(men_men_n831_), .A1(x5), .B0(men_men_n833_), .Y(men_men_n834_));
  AOI210     u0785(.A0(men_men_n834_), .A1(men_men_n826_), .B0(men_men_n72_), .Y(men_men_n835_));
  NO2        u0786(.A(men_men_n70_), .B(x3), .Y(men_men_n836_));
  OAI210     u0787(.A0(men_men_n836_), .A1(men_men_n266_), .B0(men_men_n148_), .Y(men_men_n837_));
  NO3        u0788(.A(x6), .B(x4), .C(x0), .Y(men_men_n838_));
  INV        u0789(.A(men_men_n838_), .Y(men_men_n839_));
  NO2        u0790(.A(men_men_n837_), .B(men_men_n839_), .Y(men_men_n840_));
  NO3        u0791(.A(x5), .B(x3), .C(men_men_n109_), .Y(men_men_n841_));
  AOI220     u0792(.A0(men_men_n804_), .A1(men_men_n306_), .B0(men_men_n841_), .B1(men_men_n59_), .Y(men_men_n842_));
  OR2        u0793(.A(x8), .B(x1), .Y(men_men_n843_));
  NO3        u0794(.A(men_men_n843_), .B(men_men_n842_), .C(men_men_n715_), .Y(men_men_n844_));
  NAi21      u0795(.An(x4), .B(x1), .Y(men_men_n845_));
  NO2        u0796(.A(men_men_n845_), .B(x0), .Y(men_men_n846_));
  NA2        u0797(.A(men_men_n592_), .B(men_men_n846_), .Y(men_men_n847_));
  NA3        u0798(.A(men_men_n55_), .B(x1), .C(x0), .Y(men_men_n848_));
  OAI210     u0799(.A0(men_men_n848_), .A1(men_men_n696_), .B0(men_men_n847_), .Y(men_men_n849_));
  OAI210     u0800(.A0(men_men_n849_), .A1(men_men_n844_), .B0(men_men_n317_), .Y(men_men_n850_));
  AO210      u0801(.A0(men_men_n291_), .A1(men_men_n266_), .B0(men_men_n714_), .Y(men_men_n851_));
  NA2        u0802(.A(men_men_n107_), .B(men_men_n56_), .Y(men_men_n852_));
  NO2        u0803(.A(men_men_n852_), .B(men_men_n262_), .Y(men_men_n853_));
  NO2        u0804(.A(men_men_n57_), .B(x2), .Y(men_men_n854_));
  NO4        u0805(.A(men_men_n327_), .B(men_men_n854_), .C(men_men_n795_), .D(men_men_n294_), .Y(men_men_n855_));
  AOI220     u0806(.A0(men_men_n855_), .A1(men_men_n853_), .B0(men_men_n851_), .B1(men_men_n623_), .Y(men_men_n856_));
  NA2        u0807(.A(men_men_n856_), .B(men_men_n850_), .Y(men_men_n857_));
  NO4        u0808(.A(men_men_n857_), .B(men_men_n840_), .C(men_men_n835_), .D(men_men_n819_), .Y(men09));
  AOI220     u0809(.A0(men_men_n298_), .A1(men_men_n70_), .B0(men_men_n568_), .B1(men_men_n528_), .Y(men_men_n859_));
  NA2        u0810(.A(x2), .B(men_men_n859_), .Y(men_men_n860_));
  AOI210     u0811(.A0(men_men_n860_), .A1(men_men_n735_), .B0(men_men_n439_), .Y(men_men_n861_));
  NO2        u0812(.A(men_men_n567_), .B(men_men_n265_), .Y(men_men_n862_));
  NO2        u0813(.A(men_men_n734_), .B(men_men_n337_), .Y(men_men_n863_));
  NO3        u0814(.A(men_men_n584_), .B(men_men_n101_), .C(men_men_n109_), .Y(men_men_n864_));
  AO220      u0815(.A0(men_men_n864_), .A1(men_men_n863_), .B0(men_men_n862_), .B1(men_men_n599_), .Y(men_men_n865_));
  OAI210     u0816(.A0(men_men_n865_), .A1(men_men_n861_), .B0(x4), .Y(men_men_n866_));
  OAI220     u0817(.A0(men_men_n364_), .A1(men_men_n145_), .B0(men_men_n392_), .B1(men_men_n282_), .Y(men_men_n867_));
  NO2        u0818(.A(men_men_n193_), .B(men_men_n107_), .Y(men_men_n868_));
  AOI220     u0819(.A0(men_men_n868_), .A1(men_men_n125_), .B0(men_men_n867_), .B1(men_men_n605_), .Y(men_men_n869_));
  NO2        u0820(.A(men_men_n768_), .B(men_men_n95_), .Y(men_men_n870_));
  NAi21      u0821(.An(x0), .B(x2), .Y(men_men_n871_));
  NO2        u0822(.A(men_men_n300_), .B(men_men_n871_), .Y(men_men_n872_));
  NA2        u0823(.A(men_men_n872_), .B(men_men_n870_), .Y(men_men_n873_));
  OAI210     u0824(.A0(men_men_n869_), .A1(men_men_n55_), .B0(men_men_n873_), .Y(men_men_n874_));
  NA2        u0825(.A(men_men_n874_), .B(men_men_n56_), .Y(men_men_n875_));
  NO2        u0826(.A(men_men_n56_), .B(men_men_n59_), .Y(men_men_n876_));
  INV        u0827(.A(men_men_n125_), .Y(men_men_n877_));
  NA2        u0828(.A(men_men_n734_), .B(men_men_n55_), .Y(men_men_n878_));
  AOI210     u0829(.A0(x6), .A1(x1), .B0(x5), .Y(men_men_n879_));
  NA2        u0830(.A(men_men_n879_), .B(x2), .Y(men_men_n880_));
  AOI210     u0831(.A0(men_men_n880_), .A1(men_men_n878_), .B0(men_men_n877_), .Y(men_men_n881_));
  NA2        u0832(.A(men_men_n541_), .B(men_men_n55_), .Y(men_men_n882_));
  NO4        u0833(.A(men_men_n57_), .B(x6), .C(x5), .D(x1), .Y(men_men_n883_));
  NO2        u0834(.A(men_men_n232_), .B(men_men_n382_), .Y(men_men_n884_));
  NO2        u0835(.A(men_men_n307_), .B(men_men_n149_), .Y(men_men_n885_));
  NO3        u0836(.A(men_men_n885_), .B(men_men_n884_), .C(men_men_n883_), .Y(men_men_n886_));
  OAI220     u0837(.A0(men_men_n886_), .A1(men_men_n55_), .B0(men_men_n882_), .B1(men_men_n450_), .Y(men_men_n887_));
  OAI210     u0838(.A0(men_men_n887_), .A1(men_men_n881_), .B0(men_men_n876_), .Y(men_men_n888_));
  NO2        u0839(.A(men_men_n399_), .B(men_men_n107_), .Y(men_men_n889_));
  NO2        u0840(.A(men_men_n331_), .B(men_men_n485_), .Y(men_men_n890_));
  AOI220     u0841(.A0(men_men_n890_), .A1(men_men_n889_), .B0(men_men_n211_), .B1(men_men_n230_), .Y(men_men_n891_));
  NA4        u0842(.A(men_men_n891_), .B(men_men_n888_), .C(men_men_n875_), .D(men_men_n866_), .Y(men_men_n892_));
  NA2        u0843(.A(men_men_n892_), .B(men_men_n50_), .Y(men_men_n893_));
  NO2        u0844(.A(men_men_n375_), .B(men_men_n162_), .Y(men_men_n894_));
  NA2        u0845(.A(men_men_n241_), .B(men_men_n568_), .Y(men_men_n895_));
  OAI210     u0846(.A0(men_men_n426_), .A1(men_men_n796_), .B0(men_men_n895_), .Y(men_men_n896_));
  OAI210     u0847(.A0(men_men_n896_), .A1(men_men_n894_), .B0(x0), .Y(men_men_n897_));
  NO3        u0848(.A(x8), .B(x7), .C(x2), .Y(men_men_n898_));
  NO3        u0849(.A(men_men_n57_), .B(x5), .C(x2), .Y(men_men_n899_));
  OAI210     u0850(.A0(men_men_n899_), .A1(men_men_n898_), .B0(men_men_n503_), .Y(men_men_n900_));
  AOI210     u0851(.A0(men_men_n900_), .A1(men_men_n897_), .B0(x4), .Y(men_men_n901_));
  NO2        u0852(.A(men_men_n420_), .B(men_men_n148_), .Y(men_men_n902_));
  NO2        u0853(.A(men_men_n52_), .B(x2), .Y(men_men_n903_));
  NO2        u0854(.A(men_men_n107_), .B(men_men_n56_), .Y(men_men_n904_));
  NA2        u0855(.A(men_men_n904_), .B(x8), .Y(men_men_n905_));
  NA2        u0856(.A(men_men_n905_), .B(men_men_n878_), .Y(men_men_n906_));
  AO210      u0857(.A0(men_men_n906_), .A1(men_men_n903_), .B0(men_men_n902_), .Y(men_men_n907_));
  OAI210     u0858(.A0(men_men_n907_), .A1(men_men_n901_), .B0(men_men_n597_), .Y(men_men_n908_));
  NO2        u0859(.A(men_men_n261_), .B(men_men_n118_), .Y(men_men_n909_));
  OAI210     u0860(.A0(x4), .A1(x2), .B0(x0), .Y(men_men_n910_));
  NA3        u0861(.A(men_men_n586_), .B(men_men_n598_), .C(men_men_n342_), .Y(men_men_n911_));
  OAI210     u0862(.A0(men_men_n910_), .A1(men_men_n288_), .B0(men_men_n53_), .Y(men_men_n912_));
  AOI210     u0863(.A0(men_men_n911_), .A1(men_men_n910_), .B0(men_men_n912_), .Y(men_men_n913_));
  OAI210     u0864(.A0(men_men_n913_), .A1(men_men_n909_), .B0(men_men_n326_), .Y(men_men_n914_));
  AOI220     u0865(.A0(men_men_n649_), .A1(men_men_n346_), .B0(men_men_n348_), .B1(men_men_n92_), .Y(men_men_n915_));
  NA2        u0866(.A(men_men_n92_), .B(x5), .Y(men_men_n916_));
  OAI220     u0867(.A0(men_men_n916_), .A1(men_men_n843_), .B0(men_men_n915_), .B1(men_men_n318_), .Y(men_men_n917_));
  NA2        u0868(.A(men_men_n917_), .B(men_men_n68_), .Y(men_men_n918_));
  NO2        u0869(.A(men_men_n432_), .B(x2), .Y(men_men_n919_));
  NO2        u0870(.A(x7), .B(men_men_n53_), .Y(men_men_n920_));
  NA2        u0871(.A(men_men_n920_), .B(x5), .Y(men_men_n921_));
  NO2        u0872(.A(men_men_n921_), .B(men_men_n60_), .Y(men_men_n922_));
  AOI220     u0873(.A0(men_men_n922_), .A1(men_men_n919_), .B0(men_men_n650_), .B1(men_men_n245_), .Y(men_men_n923_));
  NA3        u0874(.A(men_men_n923_), .B(men_men_n918_), .C(men_men_n914_), .Y(men_men_n924_));
  NO4        u0875(.A(men_men_n911_), .B(men_men_n614_), .C(men_men_n450_), .D(men_men_n50_), .Y(men_men_n925_));
  NO2        u0876(.A(men_men_n658_), .B(men_men_n193_), .Y(men_men_n926_));
  NA2        u0877(.A(men_men_n925_), .B(men_men_n82_), .Y(men_men_n927_));
  NA2        u0878(.A(men_men_n758_), .B(x2), .Y(men_men_n928_));
  NO2        u0879(.A(x5), .B(men_men_n53_), .Y(men_men_n929_));
  NAi21      u0880(.An(x1), .B(x4), .Y(men_men_n930_));
  NA2        u0881(.A(men_men_n930_), .B(men_men_n845_), .Y(men_men_n931_));
  NA3        u0882(.A(men_men_n395_), .B(men_men_n734_), .C(men_men_n57_), .Y(men_men_n932_));
  NA2        u0883(.A(men_men_n932_), .B(men_men_n927_), .Y(men_men_n933_));
  AOI210     u0884(.A0(men_men_n924_), .A1(x6), .B0(men_men_n933_), .Y(men_men_n934_));
  NA3        u0885(.A(men_men_n934_), .B(men_men_n908_), .C(men_men_n893_), .Y(men10));
  NO2        u0886(.A(x4), .B(x1), .Y(men_men_n936_));
  NO2        u0887(.A(men_men_n936_), .B(men_men_n150_), .Y(men_men_n937_));
  NA3        u0888(.A(x5), .B(x4), .C(x0), .Y(men_men_n938_));
  OAI220     u0889(.A0(men_men_n938_), .A1(men_men_n279_), .B0(men_men_n686_), .B1(men_men_n249_), .Y(men_men_n939_));
  NA2        u0890(.A(men_men_n939_), .B(men_men_n937_), .Y(men_men_n940_));
  NO3        u0891(.A(men_men_n354_), .B(men_men_n318_), .C(men_men_n91_), .Y(men_men_n941_));
  NA3        u0892(.A(men_men_n941_), .B(men_men_n380_), .C(men_men_n62_), .Y(men_men_n942_));
  AOI210     u0893(.A0(men_men_n942_), .A1(men_men_n940_), .B0(men_men_n300_), .Y(men_men_n943_));
  NOi21      u0894(.An(men_men_n260_), .B(men_men_n139_), .Y(men_men_n944_));
  NA2        u0895(.A(x4), .B(men_men_n109_), .Y(men_men_n945_));
  NO2        u0896(.A(men_men_n321_), .B(men_men_n945_), .Y(men_men_n946_));
  NA2        u0897(.A(men_men_n929_), .B(men_men_n50_), .Y(men_men_n947_));
  NA2        u0898(.A(men_men_n585_), .B(men_men_n273_), .Y(men_men_n948_));
  NO2        u0899(.A(men_men_n948_), .B(men_men_n947_), .Y(men_men_n949_));
  OAI220     u0900(.A0(men_men_n905_), .A1(men_men_n106_), .B0(men_men_n852_), .B1(men_men_n439_), .Y(men_men_n950_));
  AOI210     u0901(.A0(men_men_n950_), .A1(men_men_n281_), .B0(men_men_n949_), .Y(men_men_n951_));
  INV        u0902(.A(men_men_n951_), .Y(men_men_n952_));
  OAI210     u0903(.A0(men_men_n952_), .A1(men_men_n943_), .B0(x7), .Y(men_men_n953_));
  NA2        u0904(.A(men_men_n55_), .B(men_men_n71_), .Y(men_men_n954_));
  AOI210     u0905(.A0(men_men_n439_), .A1(men_men_n353_), .B0(men_men_n945_), .Y(men_men_n955_));
  NO3        u0906(.A(men_men_n441_), .B(men_men_n871_), .C(x5), .Y(men_men_n956_));
  OAI210     u0907(.A0(men_men_n956_), .A1(men_men_n955_), .B0(men_men_n954_), .Y(men_men_n957_));
  NO2        u0908(.A(men_men_n354_), .B(men_men_n142_), .Y(men_men_n958_));
  NA2        u0909(.A(men_men_n958_), .B(men_men_n421_), .Y(men_men_n959_));
  AOI210     u0910(.A0(men_men_n959_), .A1(men_men_n957_), .B0(x3), .Y(men_men_n960_));
  NA2        u0911(.A(men_men_n678_), .B(men_men_n252_), .Y(men_men_n961_));
  NO2        u0912(.A(x5), .B(men_men_n109_), .Y(men_men_n962_));
  OAI210     u0913(.A0(men_men_n962_), .A1(men_men_n239_), .B0(men_men_n916_), .Y(men_men_n963_));
  NA3        u0914(.A(men_men_n457_), .B(men_men_n131_), .C(men_men_n421_), .Y(men_men_n964_));
  INV        u0915(.A(men_men_n964_), .Y(men_men_n965_));
  AOI210     u0916(.A0(men_men_n963_), .A1(men_men_n258_), .B0(men_men_n965_), .Y(men_men_n966_));
  OAI220     u0917(.A0(men_men_n966_), .A1(men_men_n59_), .B0(men_men_n961_), .B1(men_men_n691_), .Y(men_men_n967_));
  OAI210     u0918(.A0(men_men_n967_), .A1(men_men_n960_), .B0(men_men_n920_), .Y(men_men_n968_));
  NO2        u0919(.A(x4), .B(x3), .Y(men_men_n969_));
  NO2        u0920(.A(men_men_n341_), .B(men_men_n87_), .Y(men_men_n970_));
  OAI210     u0921(.A0(men_men_n970_), .A1(men_men_n280_), .B0(men_men_n431_), .Y(men_men_n971_));
  NO2        u0922(.A(men_men_n128_), .B(men_men_n253_), .Y(men_men_n972_));
  INV        u0923(.A(men_men_n358_), .Y(men_men_n973_));
  NO3        u0924(.A(x4), .B(men_men_n109_), .C(men_men_n59_), .Y(men_men_n974_));
  NOi31      u0925(.An(men_men_n974_), .B(men_men_n2551_), .C(men_men_n973_), .Y(men_men_n975_));
  NA2        u0926(.A(men_men_n55_), .B(x5), .Y(men_men_n976_));
  NO2        u0927(.A(men_men_n975_), .B(men_men_n972_), .Y(men_men_n977_));
  AOI210     u0928(.A0(men_men_n977_), .A1(men_men_n971_), .B0(men_men_n210_), .Y(men_men_n978_));
  NO2        u0929(.A(men_men_n647_), .B(men_men_n491_), .Y(men_men_n979_));
  NO2        u0930(.A(x6), .B(x2), .Y(men_men_n980_));
  NO3        u0931(.A(men_men_n980_), .B(men_men_n678_), .C(men_men_n60_), .Y(men_men_n981_));
  OAI210     u0932(.A0(men_men_n981_), .A1(men_men_n979_), .B0(men_men_n272_), .Y(men_men_n982_));
  NO2        u0933(.A(men_men_n852_), .B(men_men_n439_), .Y(men_men_n983_));
  NA3        u0934(.A(x4), .B(x3), .C(men_men_n109_), .Y(men_men_n984_));
  NO3        u0935(.A(men_men_n984_), .B(men_men_n684_), .C(men_men_n457_), .Y(men_men_n985_));
  INV        u0936(.A(men_men_n985_), .Y(men_men_n986_));
  AOI210     u0937(.A0(men_men_n986_), .A1(men_men_n982_), .B0(men_men_n450_), .Y(men_men_n987_));
  NO2        u0938(.A(men_men_n55_), .B(men_men_n56_), .Y(men_men_n988_));
  OAI220     u0939(.A0(men_men_n804_), .A1(men_men_n452_), .B0(men_men_n736_), .B1(men_men_n128_), .Y(men_men_n989_));
  NOi21      u0940(.An(men_men_n123_), .B(men_men_n122_), .Y(men_men_n990_));
  NA2        u0941(.A(men_men_n989_), .B(men_men_n115_), .Y(men_men_n991_));
  NO2        u0942(.A(men_men_n991_), .B(men_men_n988_), .Y(men_men_n992_));
  NA2        u0943(.A(men_men_n506_), .B(men_men_n262_), .Y(men_men_n993_));
  NO2        u0944(.A(men_men_n477_), .B(men_men_n567_), .Y(men_men_n994_));
  NA3        u0945(.A(men_men_n994_), .B(men_men_n993_), .C(men_men_n55_), .Y(men_men_n995_));
  NO2        u0946(.A(men_men_n185_), .B(men_men_n109_), .Y(men_men_n996_));
  NA3        u0947(.A(men_men_n996_), .B(men_men_n184_), .C(men_men_n122_), .Y(men_men_n997_));
  NA2        u0948(.A(men_men_n997_), .B(men_men_n995_), .Y(men_men_n998_));
  NO4        u0949(.A(men_men_n998_), .B(men_men_n992_), .C(men_men_n987_), .D(men_men_n978_), .Y(men_men_n999_));
  NA3        u0950(.A(men_men_n999_), .B(men_men_n968_), .C(men_men_n953_), .Y(men11));
  NA2        u0951(.A(men_men_n373_), .B(men_men_n91_), .Y(men_men_n1001_));
  INV        u0952(.A(men_men_n872_), .Y(men_men_n1002_));
  OAI220     u0953(.A0(men_men_n1002_), .A1(men_men_n53_), .B0(men_men_n1001_), .B1(men_men_n362_), .Y(men_men_n1003_));
  NO2        u0954(.A(men_men_n753_), .B(x5), .Y(men_men_n1004_));
  NO2        u0955(.A(men_men_n170_), .B(men_men_n519_), .Y(men_men_n1005_));
  AOI220     u0956(.A0(men_men_n1005_), .A1(men_men_n1004_), .B0(men_men_n1003_), .B1(x5), .Y(men_men_n1006_));
  NO2        u0957(.A(men_men_n944_), .B(men_men_n218_), .Y(men_men_n1007_));
  NO2        u0958(.A(men_men_n338_), .B(men_men_n422_), .Y(men_men_n1008_));
  AOI220     u0959(.A0(men_men_n1008_), .A1(men_men_n183_), .B0(men_men_n1007_), .B1(men_men_n166_), .Y(men_men_n1009_));
  NO2        u0960(.A(men_men_n1009_), .B(men_men_n441_), .Y(men_men_n1010_));
  NO2        u0961(.A(men_men_n253_), .B(x2), .Y(men_men_n1011_));
  OAI210     u0962(.A0(men_men_n894_), .A1(men_men_n1011_), .B0(men_men_n411_), .Y(men_men_n1012_));
  NO2        u0963(.A(men_men_n55_), .B(men_men_n107_), .Y(men_men_n1013_));
  NA2        u0964(.A(men_men_n281_), .B(men_men_n1013_), .Y(men_men_n1014_));
  NO2        u0965(.A(men_men_n71_), .B(x1), .Y(men_men_n1015_));
  NA2        u0966(.A(men_men_n1015_), .B(men_men_n78_), .Y(men_men_n1016_));
  OA220      u0967(.A0(men_men_n1016_), .A1(men_men_n593_), .B0(men_men_n1014_), .B1(men_men_n519_), .Y(men_men_n1017_));
  AOI210     u0968(.A0(men_men_n1017_), .A1(men_men_n1012_), .B0(men_men_n691_), .Y(men_men_n1018_));
  NO2        u0969(.A(men_men_n301_), .B(men_men_n53_), .Y(men_men_n1019_));
  NO2        u0970(.A(men_men_n431_), .B(x3), .Y(men_men_n1020_));
  NA2        u0971(.A(men_men_n109_), .B(x1), .Y(men_men_n1021_));
  NO2        u0972(.A(men_men_n599_), .B(men_men_n221_), .Y(men_men_n1022_));
  NA4        u0973(.A(men_men_n1022_), .B(men_men_n863_), .C(men_men_n461_), .D(men_men_n1021_), .Y(men_men_n1023_));
  NA3        u0974(.A(x6), .B(x5), .C(men_men_n109_), .Y(men_men_n1024_));
  NO2        u0975(.A(men_men_n1024_), .B(men_men_n279_), .Y(men_men_n1025_));
  NO2        u0976(.A(men_men_n441_), .B(x0), .Y(men_men_n1026_));
  NOi31      u0977(.An(men_men_n1026_), .B(men_men_n175_), .C(men_men_n51_), .Y(men_men_n1027_));
  AOI210     u0978(.A0(men_men_n1025_), .A1(men_men_n181_), .B0(men_men_n1027_), .Y(men_men_n1028_));
  NA2        u0979(.A(men_men_n1028_), .B(men_men_n1023_), .Y(men_men_n1029_));
  NO3        u0980(.A(men_men_n1029_), .B(men_men_n1018_), .C(men_men_n1010_), .Y(men_men_n1030_));
  OAI210     u0981(.A0(men_men_n1006_), .A1(men_men_n143_), .B0(men_men_n1030_), .Y(men_men_n1031_));
  NA2        u0982(.A(men_men_n843_), .B(men_men_n87_), .Y(men_men_n1032_));
  NO3        u0983(.A(men_men_n458_), .B(men_men_n758_), .C(men_men_n123_), .Y(men_men_n1033_));
  AOI210     u0984(.A0(men_men_n1032_), .A1(men_men_n100_), .B0(men_men_n1033_), .Y(men_men_n1034_));
  NO2        u0985(.A(x8), .B(x1), .Y(men_men_n1035_));
  NO3        u0986(.A(men_men_n1035_), .B(men_men_n670_), .C(men_men_n443_), .Y(men_men_n1036_));
  OAI210     u0987(.A0(men_men_n77_), .A1(men_men_n53_), .B0(men_men_n1036_), .Y(men_men_n1037_));
  OAI210     u0988(.A0(men_men_n1034_), .A1(x3), .B0(men_men_n1037_), .Y(men_men_n1038_));
  NO2        u0989(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n1039_));
  OAI210     u0990(.A0(men_men_n1039_), .A1(x2), .B0(men_men_n235_), .Y(men_men_n1040_));
  NO2        u0991(.A(men_men_n586_), .B(men_men_n233_), .Y(men_men_n1041_));
  NA2        u0992(.A(men_men_n1041_), .B(men_men_n1040_), .Y(men_men_n1042_));
  NO2        u0993(.A(men_men_n506_), .B(x4), .Y(men_men_n1043_));
  NO3        u0994(.A(men_men_n55_), .B(x6), .C(x1), .Y(men_men_n1044_));
  NOi21      u0995(.An(men_men_n1044_), .B(men_men_n477_), .Y(men_men_n1045_));
  AOI210     u0996(.A0(men_men_n1043_), .A1(men_men_n557_), .B0(men_men_n1045_), .Y(men_men_n1046_));
  NA2        u0997(.A(men_men_n1046_), .B(men_men_n1042_), .Y(men_men_n1047_));
  AOI210     u0998(.A0(men_men_n1038_), .A1(x2), .B0(men_men_n1047_), .Y(men_men_n1048_));
  NO2        u0999(.A(men_men_n233_), .B(x2), .Y(men_men_n1049_));
  NOi21      u1000(.An(men_men_n385_), .B(men_men_n548_), .Y(men_men_n1050_));
  NA2        u1001(.A(x8), .B(men_men_n109_), .Y(men_men_n1051_));
  NO2        u1002(.A(men_men_n107_), .B(x1), .Y(men_men_n1052_));
  NA2        u1003(.A(men_men_n84_), .B(men_men_n71_), .Y(men_men_n1053_));
  INV        u1004(.A(men_men_n250_), .Y(men_men_n1054_));
  NA2        u1005(.A(men_men_n1054_), .B(men_men_n150_), .Y(men_men_n1055_));
  OAI220     u1006(.A0(men_men_n1055_), .A1(men_men_n362_), .B0(men_men_n1053_), .B1(men_men_n321_), .Y(men_men_n1056_));
  NO2        u1007(.A(men_men_n160_), .B(men_men_n55_), .Y(men_men_n1057_));
  NA2        u1008(.A(men_men_n1057_), .B(men_men_n1056_), .Y(men_men_n1058_));
  OAI210     u1009(.A0(men_men_n1048_), .A1(men_men_n832_), .B0(men_men_n1058_), .Y(men_men_n1059_));
  AO210      u1010(.A0(men_men_n1031_), .A1(men_men_n57_), .B0(men_men_n1059_), .Y(men12));
  NA2        u1011(.A(men_men_n862_), .B(men_men_n249_), .Y(men_men_n1061_));
  NO2        u1012(.A(men_men_n603_), .B(x7), .Y(men_men_n1062_));
  NA2        u1013(.A(men_men_n1062_), .B(men_men_n280_), .Y(men_men_n1063_));
  NA2        u1014(.A(men_men_n683_), .B(men_men_n852_), .Y(men_men_n1064_));
  AOI210     u1015(.A0(men_men_n1063_), .A1(men_men_n1061_), .B0(men_men_n1064_), .Y(men_men_n1065_));
  NOi21      u1016(.An(men_men_n399_), .B(men_men_n539_), .Y(men_men_n1066_));
  NO2        u1017(.A(x7), .B(men_men_n50_), .Y(men_men_n1067_));
  NO3        u1018(.A(men_men_n845_), .B(men_men_n111_), .C(men_men_n98_), .Y(men_men_n1068_));
  INV        u1019(.A(men_men_n1068_), .Y(men_men_n1069_));
  NA2        u1020(.A(men_men_n1013_), .B(men_men_n56_), .Y(men_men_n1070_));
  OAI220     u1021(.A0(men_men_n1070_), .A1(men_men_n558_), .B0(men_men_n1069_), .B1(men_men_n1066_), .Y(men_men_n1071_));
  OAI210     u1022(.A0(men_men_n1071_), .A1(men_men_n1065_), .B0(men_men_n562_), .Y(men_men_n1072_));
  NA2        u1023(.A(men_men_n87_), .B(x5), .Y(men_men_n1073_));
  OAI210     u1024(.A0(men_men_n1073_), .A1(men_men_n321_), .B0(men_men_n701_), .Y(men_men_n1074_));
  AOI210     u1025(.A0(men_men_n806_), .A1(men_men_n117_), .B0(men_men_n1074_), .Y(men_men_n1075_));
  NA2        u1026(.A(men_men_n584_), .B(men_men_n53_), .Y(men_men_n1076_));
  NA2        u1027(.A(men_men_n288_), .B(men_men_n50_), .Y(men_men_n1077_));
  NO2        u1028(.A(men_men_n1076_), .B(men_men_n136_), .Y(men_men_n1078_));
  NO2        u1029(.A(men_men_n1032_), .B(men_men_n501_), .Y(men_men_n1079_));
  NO4        u1030(.A(men_men_n241_), .B(men_men_n272_), .C(men_men_n60_), .D(men_men_n57_), .Y(men_men_n1080_));
  AOI220     u1031(.A0(men_men_n1080_), .A1(men_men_n1079_), .B0(men_men_n1078_), .B1(men_men_n56_), .Y(men_men_n1081_));
  OAI210     u1032(.A0(men_men_n1075_), .A1(men_men_n64_), .B0(men_men_n1081_), .Y(men_men_n1082_));
  NO2        u1033(.A(men_men_n57_), .B(x0), .Y(men_men_n1083_));
  NO2        u1034(.A(men_men_n647_), .B(men_men_n318_), .Y(men_men_n1084_));
  NO2        u1035(.A(men_men_n736_), .B(x3), .Y(men_men_n1085_));
  NO2        u1036(.A(men_men_n645_), .B(x8), .Y(men_men_n1086_));
  AOI220     u1037(.A0(men_men_n1086_), .A1(men_men_n1085_), .B0(men_men_n1084_), .B1(men_men_n1083_), .Y(men_men_n1087_));
  AOI210     u1038(.A0(men_men_n670_), .A1(men_men_n249_), .B0(x7), .Y(men_men_n1088_));
  NO2        u1039(.A(men_men_n1088_), .B(x8), .Y(men_men_n1089_));
  NA4        u1040(.A(men_men_n649_), .B(men_men_n641_), .C(men_men_n207_), .D(x0), .Y(men_men_n1090_));
  OAI220     u1041(.A0(men_men_n1090_), .A1(men_men_n1089_), .B0(men_men_n1087_), .B1(men_men_n556_), .Y(men_men_n1091_));
  AOI210     u1042(.A0(men_men_n1082_), .A1(men_men_n980_), .B0(men_men_n1091_), .Y(men_men_n1092_));
  NO2        u1043(.A(men_men_n249_), .B(men_men_n55_), .Y(men_men_n1093_));
  NO2        u1044(.A(men_men_n257_), .B(x8), .Y(men_men_n1094_));
  NOi32      u1045(.An(men_men_n1094_), .Bn(men_men_n206_), .C(men_men_n549_), .Y(men_men_n1095_));
  NO2        u1046(.A(men_men_n88_), .B(men_men_n60_), .Y(men_men_n1096_));
  OAI210     u1047(.A0(men_men_n1095_), .A1(men_men_n1093_), .B0(men_men_n1096_), .Y(men_men_n1097_));
  NO2        u1048(.A(men_men_n920_), .B(men_men_n99_), .Y(men_men_n1098_));
  NO2        u1049(.A(men_men_n169_), .B(men_men_n53_), .Y(men_men_n1099_));
  NA2        u1050(.A(men_men_n1098_), .B(men_men_n658_), .Y(men_men_n1100_));
  NO2        u1051(.A(x7), .B(x0), .Y(men_men_n1101_));
  NO3        u1052(.A(men_men_n160_), .B(men_men_n1101_), .C(men_men_n147_), .Y(men_men_n1102_));
  XN2        u1053(.A(x8), .B(x7), .Y(men_men_n1103_));
  NO3        u1054(.A(men_men_n1035_), .B(men_men_n260_), .C(men_men_n1103_), .Y(men_men_n1104_));
  OAI210     u1055(.A0(men_men_n1104_), .A1(men_men_n1102_), .B0(men_men_n715_), .Y(men_men_n1105_));
  NO2        u1056(.A(men_men_n269_), .B(men_men_n265_), .Y(men_men_n1106_));
  NO2        u1057(.A(men_men_n107_), .B(x4), .Y(men_men_n1107_));
  OAI210     u1058(.A0(men_men_n1106_), .A1(men_men_n280_), .B0(men_men_n1107_), .Y(men_men_n1108_));
  NA4        u1059(.A(men_men_n1108_), .B(men_men_n1105_), .C(men_men_n1100_), .D(men_men_n1097_), .Y(men_men_n1109_));
  NA2        u1060(.A(men_men_n1109_), .B(men_men_n541_), .Y(men_men_n1110_));
  NO2        u1061(.A(men_men_n55_), .B(x4), .Y(men_men_n1111_));
  NA2        u1062(.A(men_men_n1111_), .B(men_men_n165_), .Y(men_men_n1112_));
  NA2        u1063(.A(men_men_n983_), .B(men_men_n50_), .Y(men_men_n1113_));
  AOI210     u1064(.A0(men_men_n1113_), .A1(men_men_n1112_), .B0(men_men_n426_), .Y(men_men_n1114_));
  OAI220     u1065(.A0(men_men_n290_), .A1(men_men_n278_), .B0(men_men_n265_), .B1(men_men_n244_), .Y(men_men_n1115_));
  NA3        u1066(.A(men_men_n1115_), .B(men_men_n658_), .C(x1), .Y(men_men_n1116_));
  OAI210     u1067(.A0(x8), .A1(x0), .B0(x4), .Y(men_men_n1117_));
  NO2        u1068(.A(x7), .B(men_men_n56_), .Y(men_men_n1118_));
  NO2        u1069(.A(men_men_n68_), .B(men_men_n1118_), .Y(men_men_n1119_));
  NOi21      u1070(.An(men_men_n1117_), .B(men_men_n1119_), .Y(men_men_n1120_));
  NO2        u1071(.A(men_men_n649_), .B(men_men_n321_), .Y(men_men_n1121_));
  NO2        u1072(.A(men_men_n761_), .B(men_men_n222_), .Y(men_men_n1122_));
  OAI210     u1073(.A0(men_men_n1121_), .A1(men_men_n1120_), .B0(men_men_n1122_), .Y(men_men_n1123_));
  NO2        u1074(.A(men_men_n143_), .B(men_men_n142_), .Y(men_men_n1124_));
  NA2        u1075(.A(men_men_n1124_), .B(men_men_n257_), .Y(men_men_n1125_));
  NO2        u1076(.A(men_men_n802_), .B(men_men_n418_), .Y(men_men_n1126_));
  NA2        u1077(.A(men_men_n326_), .B(men_men_n59_), .Y(men_men_n1127_));
  NO2        u1078(.A(men_men_n1070_), .B(men_men_n1127_), .Y(men_men_n1128_));
  AOI210     u1079(.A0(men_men_n1126_), .A1(men_men_n181_), .B0(men_men_n1128_), .Y(men_men_n1129_));
  NA4        u1080(.A(men_men_n1129_), .B(men_men_n1125_), .C(men_men_n1123_), .D(men_men_n1116_), .Y(men_men_n1130_));
  OAI210     u1081(.A0(men_men_n1130_), .A1(men_men_n1114_), .B0(men_men_n660_), .Y(men_men_n1131_));
  NA4        u1082(.A(men_men_n1131_), .B(men_men_n1110_), .C(men_men_n1092_), .D(men_men_n1072_), .Y(men13));
  NO2        u1083(.A(men_men_n457_), .B(men_men_n348_), .Y(men_men_n1133_));
  NOi41      u1084(.An(men_men_n1133_), .B(men_men_n658_), .C(men_men_n292_), .D(men_men_n241_), .Y(men_men_n1134_));
  NO2        u1085(.A(men_men_n845_), .B(men_men_n185_), .Y(men_men_n1135_));
  NO2        u1086(.A(men_men_n159_), .B(men_men_n71_), .Y(men_men_n1136_));
  XN2        u1087(.A(x4), .B(x0), .Y(men_men_n1137_));
  NO3        u1088(.A(men_men_n1137_), .B(men_men_n110_), .C(men_men_n418_), .Y(men_men_n1138_));
  AO220      u1089(.A0(men_men_n1138_), .A1(men_men_n1136_), .B0(men_men_n1135_), .B1(men_men_n327_), .Y(men_men_n1139_));
  OAI210     u1090(.A0(men_men_n1139_), .A1(men_men_n1134_), .B0(x3), .Y(men_men_n1140_));
  NO2        u1091(.A(men_men_n845_), .B(x6), .Y(men_men_n1141_));
  INV        u1092(.A(men_men_n1077_), .Y(men_men_n1142_));
  NO3        u1093(.A(x8), .B(x5), .C(men_men_n109_), .Y(men_men_n1143_));
  NA2        u1094(.A(men_men_n1143_), .B(men_men_n623_), .Y(men_men_n1144_));
  NO2        u1095(.A(men_men_n586_), .B(men_men_n201_), .Y(men_men_n1145_));
  NA2        u1096(.A(men_men_n1145_), .B(men_men_n1044_), .Y(men_men_n1146_));
  NA2        u1097(.A(men_men_n443_), .B(men_men_n53_), .Y(men_men_n1147_));
  NO2        u1098(.A(men_men_n1147_), .B(men_men_n916_), .Y(men_men_n1148_));
  NA2        u1099(.A(men_men_n1070_), .B(men_men_n462_), .Y(men_men_n1149_));
  NA2        u1100(.A(men_men_n56_), .B(men_men_n109_), .Y(men_men_n1150_));
  NA2        u1101(.A(men_men_n1150_), .B(x1), .Y(men_men_n1151_));
  NO2        u1102(.A(men_men_n1151_), .B(men_men_n262_), .Y(men_men_n1152_));
  NO2        u1103(.A(men_men_n318_), .B(x6), .Y(men_men_n1153_));
  OAI210     u1104(.A0(men_men_n253_), .A1(men_men_n945_), .B0(men_men_n928_), .Y(men_men_n1154_));
  AOI220     u1105(.A0(men_men_n1154_), .A1(men_men_n1153_), .B0(men_men_n1152_), .B1(men_men_n1149_), .Y(men_men_n1155_));
  NAi41      u1106(.An(men_men_n1148_), .B(men_men_n1155_), .C(men_men_n1146_), .D(men_men_n1144_), .Y(men_men_n1156_));
  NA2        u1107(.A(men_men_n1156_), .B(men_men_n68_), .Y(men_men_n1157_));
  NA2        u1108(.A(men_men_n71_), .B(x3), .Y(men_men_n1158_));
  NA2        u1109(.A(men_men_n1158_), .B(men_men_n878_), .Y(men_men_n1159_));
  OAI220     u1110(.A0(men_men_n300_), .A1(men_men_n802_), .B0(men_men_n87_), .B1(men_men_n77_), .Y(men_men_n1160_));
  AOI210     u1111(.A0(men_men_n1073_), .A1(men_men_n597_), .B0(men_men_n945_), .Y(men_men_n1161_));
  OA210      u1112(.A0(men_men_n1160_), .A1(men_men_n1159_), .B0(men_men_n1161_), .Y(men_men_n1162_));
  NA2        u1113(.A(men_men_n599_), .B(men_men_n55_), .Y(men_men_n1163_));
  NA2        u1114(.A(men_men_n494_), .B(men_men_n485_), .Y(men_men_n1164_));
  NA2        u1115(.A(x6), .B(men_men_n50_), .Y(men_men_n1165_));
  NA2        u1116(.A(men_men_n1165_), .B(men_men_n528_), .Y(men_men_n1166_));
  NO2        u1117(.A(men_men_n162_), .B(men_men_n131_), .Y(men_men_n1167_));
  AOI210     u1118(.A0(men_men_n1166_), .A1(men_men_n427_), .B0(men_men_n1167_), .Y(men_men_n1168_));
  OAI220     u1119(.A0(men_men_n1168_), .A1(men_men_n852_), .B0(men_men_n1164_), .B1(men_men_n1163_), .Y(men_men_n1169_));
  OAI210     u1120(.A0(men_men_n1169_), .A1(men_men_n1162_), .B0(men_men_n1101_), .Y(men_men_n1170_));
  NAi21      u1121(.An(men_men_n84_), .B(men_men_n380_), .Y(men_men_n1171_));
  NO2        u1122(.A(men_men_n1171_), .B(men_men_n71_), .Y(men_men_n1172_));
  AOI210     u1123(.A0(men_men_n165_), .A1(x4), .B0(men_men_n177_), .Y(men_men_n1173_));
  NO2        u1124(.A(men_men_n1173_), .B(x0), .Y(men_men_n1174_));
  NA2        u1125(.A(men_men_n1174_), .B(men_men_n1172_), .Y(men_men_n1175_));
  NO2        u1126(.A(x4), .B(x0), .Y(men_men_n1176_));
  NO3        u1127(.A(men_men_n962_), .B(men_men_n250_), .C(men_men_n528_), .Y(men_men_n1177_));
  OAI210     u1128(.A0(men_men_n1177_), .A1(men_men_n202_), .B0(men_men_n1176_), .Y(men_men_n1178_));
  NA2        u1129(.A(men_men_n1178_), .B(men_men_n1175_), .Y(men_men_n1179_));
  NA2        u1130(.A(men_men_n252_), .B(men_men_n715_), .Y(men_men_n1180_));
  NO2        u1131(.A(men_men_n1180_), .B(men_men_n508_), .Y(men_men_n1181_));
  NA2        u1132(.A(men_men_n56_), .B(x0), .Y(men_men_n1182_));
  NO3        u1133(.A(men_men_n1182_), .B(men_men_n485_), .C(men_men_n81_), .Y(men_men_n1183_));
  OAI210     u1134(.A0(men_men_n1183_), .A1(men_men_n1181_), .B0(x2), .Y(men_men_n1184_));
  NO2        u1135(.A(men_men_n670_), .B(x0), .Y(men_men_n1185_));
  NA2        u1136(.A(men_men_n1185_), .B(men_men_n330_), .Y(men_men_n1186_));
  NO2        u1137(.A(men_men_n773_), .B(x1), .Y(men_men_n1187_));
  AOI220     u1138(.A0(men_men_n1187_), .A1(men_men_n592_), .B0(men_men_n470_), .B1(men_men_n295_), .Y(men_men_n1188_));
  AOI220     u1139(.A0(x3), .A1(men_men_n1135_), .B0(men_men_n946_), .B1(men_men_n100_), .Y(men_men_n1189_));
  NA4        u1140(.A(men_men_n1189_), .B(men_men_n1188_), .C(men_men_n1186_), .D(men_men_n1184_), .Y(men_men_n1190_));
  AOI220     u1141(.A0(men_men_n1190_), .A1(men_men_n132_), .B0(men_men_n1179_), .B1(men_men_n67_), .Y(men_men_n1191_));
  NA4        u1142(.A(men_men_n1191_), .B(men_men_n1170_), .C(men_men_n1157_), .D(men_men_n1140_), .Y(men14));
  NO2        u1143(.A(men_men_n368_), .B(men_men_n71_), .Y(men_men_n1193_));
  NO3        u1144(.A(x7), .B(x6), .C(x0), .Y(men_men_n1194_));
  OAI210     u1145(.A0(men_men_n1194_), .A1(men_men_n1193_), .B0(x8), .Y(men_men_n1195_));
  NA2        u1146(.A(men_men_n1086_), .B(men_men_n85_), .Y(men_men_n1196_));
  AOI210     u1147(.A0(men_men_n1196_), .A1(men_men_n1195_), .B0(men_men_n158_), .Y(men_men_n1197_));
  AOI220     u1148(.A0(men_men_n372_), .A1(men_men_n832_), .B0(men_men_n443_), .B1(men_men_n418_), .Y(men_men_n1198_));
  NA2        u1149(.A(men_men_n281_), .B(men_men_n944_), .Y(men_men_n1199_));
  OAI220     u1150(.A0(men_men_n1199_), .A1(men_men_n1198_), .B0(men_men_n460_), .B1(men_men_n788_), .Y(men_men_n1200_));
  OA210      u1151(.A0(men_men_n1200_), .A1(men_men_n1197_), .B0(x4), .Y(men_men_n1201_));
  NO2        u1152(.A(men_men_n142_), .B(men_men_n590_), .Y(men_men_n1202_));
  NA2        u1153(.A(x6), .B(x2), .Y(men_men_n1203_));
  NO2        u1154(.A(men_men_n608_), .B(men_men_n1203_), .Y(men_men_n1204_));
  OA210      u1155(.A0(men_men_n1202_), .A1(men_men_n215_), .B0(men_men_n1204_), .Y(men_men_n1205_));
  NO4        u1156(.A(men_men_n586_), .B(men_men_n373_), .C(men_men_n298_), .D(men_men_n115_), .Y(men_men_n1206_));
  OAI210     u1157(.A0(men_men_n1206_), .A1(men_men_n1205_), .B0(men_men_n59_), .Y(men_men_n1207_));
  NA2        u1158(.A(x6), .B(men_men_n107_), .Y(men_men_n1208_));
  NO2        u1159(.A(men_men_n647_), .B(men_men_n1208_), .Y(men_men_n1209_));
  NA2        u1160(.A(men_men_n1209_), .B(men_men_n903_), .Y(men_men_n1210_));
  AOI210     u1161(.A0(men_men_n1086_), .A1(men_men_n974_), .B0(x1), .Y(men_men_n1211_));
  NO2        u1162(.A(men_men_n523_), .B(x5), .Y(men_men_n1212_));
  NA3        u1163(.A(men_men_n1212_), .B(men_men_n122_), .C(x0), .Y(men_men_n1213_));
  NA4        u1164(.A(men_men_n677_), .B(men_men_n904_), .C(men_men_n300_), .D(men_men_n68_), .Y(men_men_n1214_));
  AN4        u1165(.A(men_men_n1214_), .B(men_men_n1213_), .C(men_men_n1211_), .D(men_men_n1210_), .Y(men_men_n1215_));
  NO2        u1166(.A(men_men_n684_), .B(men_men_n1051_), .Y(men_men_n1216_));
  NO2        u1167(.A(men_men_n77_), .B(men_men_n58_), .Y(men_men_n1217_));
  OAI210     u1168(.A0(men_men_n1216_), .A1(men_men_n440_), .B0(men_men_n1217_), .Y(men_men_n1218_));
  AO210      u1169(.A0(men_men_n1193_), .A1(men_men_n974_), .B0(men_men_n53_), .Y(men_men_n1219_));
  AOI210     u1170(.A0(men_men_n749_), .A1(men_men_n796_), .B0(men_men_n1219_), .Y(men_men_n1220_));
  AOI220     u1171(.A0(men_men_n1220_), .A1(men_men_n1218_), .B0(men_men_n1215_), .B1(men_men_n1207_), .Y(men_men_n1221_));
  NO2        u1172(.A(men_men_n659_), .B(men_men_n169_), .Y(men_men_n1222_));
  NO3        u1173(.A(men_men_n1222_), .B(men_men_n1221_), .C(men_men_n1201_), .Y(men_men_n1223_));
  NO2        u1174(.A(men_men_n318_), .B(x2), .Y(men_men_n1224_));
  XN2        u1175(.A(x4), .B(x1), .Y(men_men_n1225_));
  NO2        u1176(.A(men_men_n1225_), .B(men_men_n300_), .Y(men_men_n1226_));
  NO2        u1177(.A(men_men_n337_), .B(men_men_n60_), .Y(men_men_n1227_));
  OAI210     u1178(.A0(men_men_n1227_), .A1(men_men_n1226_), .B0(men_men_n1224_), .Y(men_men_n1228_));
  NA2        u1179(.A(men_men_n671_), .B(men_men_n56_), .Y(men_men_n1229_));
  OAI220     u1180(.A0(men_men_n1229_), .A1(men_men_n159_), .B0(men_men_n193_), .B1(men_men_n71_), .Y(men_men_n1230_));
  NO2        u1181(.A(men_men_n218_), .B(men_men_n260_), .Y(men_men_n1231_));
  AOI220     u1182(.A0(men_men_n139_), .A1(men_men_n56_), .B0(men_men_n92_), .B1(x5), .Y(men_men_n1232_));
  NA2        u1183(.A(men_men_n1044_), .B(men_men_n305_), .Y(men_men_n1233_));
  NA2        u1184(.A(men_men_n252_), .B(men_men_n352_), .Y(men_men_n1234_));
  NA2        u1185(.A(men_men_n622_), .B(men_men_n990_), .Y(men_men_n1235_));
  OAI220     u1186(.A0(men_men_n1235_), .A1(men_men_n1234_), .B0(men_men_n1233_), .B1(men_men_n1232_), .Y(men_men_n1236_));
  AOI210     u1187(.A0(men_men_n1231_), .A1(men_men_n1230_), .B0(men_men_n1236_), .Y(men_men_n1237_));
  AOI210     u1188(.A0(men_men_n1237_), .A1(men_men_n1228_), .B0(x7), .Y(men_men_n1238_));
  NO2        u1189(.A(men_men_n484_), .B(x6), .Y(men_men_n1239_));
  AOI210     u1190(.A0(men_men_n798_), .A1(men_men_n929_), .B0(men_men_n1239_), .Y(men_men_n1240_));
  OAI220     u1191(.A0(men_men_n1240_), .A1(men_men_n55_), .B0(men_men_n484_), .B1(men_men_n103_), .Y(men_men_n1241_));
  NA2        u1192(.A(men_men_n1241_), .B(men_men_n354_), .Y(men_men_n1242_));
  NA3        u1193(.A(men_men_n593_), .B(men_men_n1021_), .C(men_men_n70_), .Y(men_men_n1243_));
  NO4        u1194(.A(men_men_n1243_), .B(men_men_n1182_), .C(men_men_n120_), .D(men_men_n55_), .Y(men_men_n1244_));
  NO3        u1195(.A(men_men_n1016_), .B(men_men_n804_), .C(men_men_n475_), .Y(men_men_n1245_));
  NO3        u1196(.A(men_men_n736_), .B(men_men_n491_), .C(men_men_n54_), .Y(men_men_n1246_));
  NO4        u1197(.A(men_men_n1246_), .B(men_men_n1245_), .C(men_men_n1244_), .D(men_men_n994_), .Y(men_men_n1247_));
  AOI210     u1198(.A0(men_men_n1247_), .A1(men_men_n1242_), .B0(men_men_n302_), .Y(men_men_n1248_));
  NA2        u1199(.A(men_men_n876_), .B(men_men_n53_), .Y(men_men_n1249_));
  OAI210     u1200(.A0(men_men_n247_), .A1(men_men_n117_), .B0(x2), .Y(men_men_n1250_));
  NA2        u1201(.A(men_men_n364_), .B(men_men_n56_), .Y(men_men_n1251_));
  OA220      u1202(.A0(men_men_n1251_), .A1(men_men_n1250_), .B0(men_men_n1249_), .B1(men_men_n372_), .Y(men_men_n1252_));
  NA3        u1203(.A(men_men_n994_), .B(men_men_n720_), .C(men_men_n55_), .Y(men_men_n1253_));
  NA2        u1204(.A(men_men_n56_), .B(x2), .Y(men_men_n1254_));
  NO2        u1205(.A(men_men_n1254_), .B(men_men_n200_), .Y(men_men_n1255_));
  NA4        u1206(.A(men_men_n1255_), .B(men_men_n364_), .C(men_men_n260_), .D(men_men_n67_), .Y(men_men_n1256_));
  NA3        u1207(.A(men_men_n1187_), .B(men_men_n599_), .C(men_men_n613_), .Y(men_men_n1257_));
  AN3        u1208(.A(men_men_n1257_), .B(men_men_n1256_), .C(men_men_n1253_), .Y(men_men_n1258_));
  OAI210     u1209(.A0(men_men_n1252_), .A1(men_men_n313_), .B0(men_men_n1258_), .Y(men_men_n1259_));
  NO3        u1210(.A(men_men_n1259_), .B(men_men_n1248_), .C(men_men_n1238_), .Y(men_men_n1260_));
  OAI210     u1211(.A0(men_men_n1223_), .A1(x3), .B0(men_men_n1260_), .Y(men15));
  NA2        u1212(.A(men_men_n568_), .B(men_men_n59_), .Y(men_men_n1262_));
  NO2        u1213(.A(men_men_n1262_), .B(men_men_n53_), .Y(men_men_n1263_));
  NA3        u1214(.A(men_men_n57_), .B(x6), .C(men_men_n109_), .Y(men_men_n1264_));
  NO2        u1215(.A(men_men_n1264_), .B(men_men_n294_), .Y(men_men_n1265_));
  OAI210     u1216(.A0(men_men_n1265_), .A1(men_men_n1263_), .B0(men_men_n1107_), .Y(men_men_n1266_));
  NA2        u1217(.A(men_men_n111_), .B(men_men_n109_), .Y(men_men_n1267_));
  NA4        u1218(.A(men_men_n1267_), .B(men_men_n620_), .C(men_men_n306_), .D(x6), .Y(men_men_n1268_));
  INV        u1219(.A(x3), .Y(men_men_n1269_));
  NA3        u1220(.A(men_men_n1269_), .B(men_men_n1268_), .C(men_men_n1266_), .Y(men_men_n1270_));
  AOI210     u1221(.A0(men_men_n1026_), .A1(men_men_n572_), .B0(men_men_n50_), .Y(men_men_n1271_));
  NO2        u1222(.A(men_men_n294_), .B(men_men_n109_), .Y(men_men_n1272_));
  NO2        u1223(.A(men_men_n239_), .B(x5), .Y(men_men_n1273_));
  NA2        u1224(.A(men_men_n1273_), .B(men_men_n1272_), .Y(men_men_n1274_));
  NA3        u1225(.A(men_men_n1187_), .B(men_men_n607_), .C(men_men_n1118_), .Y(men_men_n1275_));
  NA4        u1226(.A(men_men_n1275_), .B(men_men_n1274_), .C(men_men_n1271_), .D(men_men_n1213_), .Y(men_men_n1276_));
  NA2        u1227(.A(men_men_n331_), .B(men_men_n340_), .Y(men_men_n1277_));
  AOI210     u1228(.A0(men_men_n1151_), .A1(men_men_n58_), .B0(men_men_n1277_), .Y(men_men_n1278_));
  NA4        u1229(.A(men_men_n1151_), .B(men_men_n683_), .C(men_men_n1083_), .D(men_men_n380_), .Y(men_men_n1279_));
  NO2        u1230(.A(men_men_n736_), .B(men_men_n53_), .Y(men_men_n1280_));
  NO2        u1231(.A(men_men_n761_), .B(men_men_n298_), .Y(men_men_n1281_));
  NA2        u1232(.A(men_men_n1281_), .B(men_men_n1280_), .Y(men_men_n1282_));
  NA2        u1233(.A(men_men_n1282_), .B(men_men_n1279_), .Y(men_men_n1283_));
  OAI210     u1234(.A0(men_men_n1283_), .A1(men_men_n1278_), .B0(men_men_n77_), .Y(men_men_n1284_));
  NA2        u1235(.A(men_men_n366_), .B(men_men_n686_), .Y(men_men_n1285_));
  NA2        u1236(.A(men_men_n555_), .B(men_men_n56_), .Y(men_men_n1286_));
  NA3        u1237(.A(men_men_n1286_), .B(men_men_n340_), .C(men_men_n111_), .Y(men_men_n1287_));
  AOI210     u1238(.A0(men_men_n1287_), .A1(men_men_n1285_), .B0(men_men_n491_), .Y(men_men_n1288_));
  NO3        u1239(.A(men_men_n786_), .B(men_men_n604_), .C(men_men_n201_), .Y(men_men_n1289_));
  OAI210     u1240(.A0(men_men_n1289_), .A1(men_men_n1288_), .B0(men_men_n484_), .Y(men_men_n1290_));
  NO2        u1241(.A(men_men_n852_), .B(men_men_n50_), .Y(men_men_n1291_));
  NO2        u1242(.A(men_men_n249_), .B(men_men_n64_), .Y(men_men_n1292_));
  OA210      u1243(.A0(men_men_n1292_), .A1(men_men_n1291_), .B0(men_men_n406_), .Y(men_men_n1293_));
  NA2        u1244(.A(men_men_n57_), .B(x3), .Y(men_men_n1294_));
  NO2        u1245(.A(men_men_n1294_), .B(men_men_n665_), .Y(men_men_n1295_));
  OAI210     u1246(.A0(men_men_n1295_), .A1(men_men_n1293_), .B0(men_men_n980_), .Y(men_men_n1296_));
  NA2        u1247(.A(men_men_n1255_), .B(men_men_n68_), .Y(men_men_n1297_));
  NO2        u1248(.A(men_men_n1203_), .B(x0), .Y(men_men_n1298_));
  AOI210     u1249(.A0(men_men_n1298_), .A1(men_men_n587_), .B0(x8), .Y(men_men_n1299_));
  NO2        u1250(.A(men_men_n426_), .B(men_men_n81_), .Y(men_men_n1300_));
  NO2        u1251(.A(men_men_n910_), .B(men_men_n71_), .Y(men_men_n1301_));
  NA2        u1252(.A(men_men_n1301_), .B(men_men_n1300_), .Y(men_men_n1302_));
  NO2        u1253(.A(men_men_n945_), .B(x6), .Y(men_men_n1303_));
  NA4        u1254(.A(men_men_n1303_), .B(men_men_n577_), .C(men_men_n160_), .D(men_men_n410_), .Y(men_men_n1304_));
  AN4        u1255(.A(men_men_n1304_), .B(men_men_n1302_), .C(men_men_n1299_), .D(men_men_n1297_), .Y(men_men_n1305_));
  NA4        u1256(.A(men_men_n1305_), .B(men_men_n1296_), .C(men_men_n1290_), .D(men_men_n1284_), .Y(men_men_n1306_));
  NA2        u1257(.A(men_men_n166_), .B(men_men_n720_), .Y(men_men_n1307_));
  NO2        u1258(.A(men_men_n632_), .B(x2), .Y(men_men_n1308_));
  OAI210     u1259(.A0(men_men_n68_), .A1(men_men_n53_), .B0(men_men_n145_), .Y(men_men_n1309_));
  OAI210     u1260(.A0(men_men_n1308_), .A1(men_men_n85_), .B0(men_men_n1309_), .Y(men_men_n1310_));
  AOI210     u1261(.A0(men_men_n1310_), .A1(men_men_n1307_), .B0(men_men_n318_), .Y(men_men_n1311_));
  NO3        u1262(.A(men_men_n1264_), .B(men_men_n268_), .C(men_men_n249_), .Y(men_men_n1312_));
  NA3        u1263(.A(men_men_n57_), .B(x1), .C(x0), .Y(men_men_n1313_));
  NA3        u1264(.A(men_men_n71_), .B(x5), .C(x2), .Y(men_men_n1314_));
  NA4        u1265(.A(x7), .B(x3), .C(men_men_n53_), .D(x0), .Y(men_men_n1315_));
  OAI220     u1266(.A0(men_men_n1315_), .A1(x6), .B0(men_men_n1314_), .B1(men_men_n1313_), .Y(men_men_n1316_));
  NO2        u1267(.A(men_men_n1316_), .B(men_men_n1312_), .Y(men_men_n1317_));
  NAi21      u1268(.An(men_men_n115_), .B(men_men_n730_), .Y(men_men_n1318_));
  NA4        u1269(.A(men_men_n1318_), .B(men_men_n316_), .C(men_men_n290_), .D(men_men_n607_), .Y(men_men_n1319_));
  OAI220     u1270(.A0(men_men_n321_), .A1(x7), .B0(men_men_n131_), .B1(men_men_n71_), .Y(men_men_n1320_));
  NA3        u1271(.A(men_men_n1320_), .B(men_men_n773_), .C(men_men_n1052_), .Y(men_men_n1321_));
  NA2        u1272(.A(men_men_n82_), .B(men_men_n50_), .Y(men_men_n1322_));
  AO210      u1273(.A0(men_men_n1322_), .A1(men_men_n311_), .B0(men_men_n158_), .Y(men_men_n1323_));
  NA4        u1274(.A(men_men_n1323_), .B(men_men_n1321_), .C(men_men_n1319_), .D(men_men_n1317_), .Y(men_men_n1324_));
  OAI210     u1275(.A0(men_men_n1324_), .A1(men_men_n1311_), .B0(men_men_n56_), .Y(men_men_n1325_));
  AOI210     u1276(.A0(men_men_n673_), .A1(x4), .B0(men_men_n929_), .Y(men_men_n1326_));
  OAI220     u1277(.A0(men_men_n1326_), .A1(men_men_n299_), .B0(men_men_n984_), .B1(men_men_n921_), .Y(men_men_n1327_));
  NA2        u1278(.A(men_men_n1327_), .B(x6), .Y(men_men_n1328_));
  NO2        u1279(.A(men_men_n57_), .B(men_men_n59_), .Y(men_men_n1329_));
  NO2        u1280(.A(x7), .B(x5), .Y(men_men_n1330_));
  AOI220     u1281(.A0(men_men_n836_), .A1(men_men_n1329_), .B0(men_men_n527_), .B1(men_men_n1330_), .Y(men_men_n1331_));
  NA2        u1282(.A(men_men_n746_), .B(men_men_n291_), .Y(men_men_n1332_));
  NA3        u1283(.A(men_men_n599_), .B(men_men_n293_), .C(men_men_n244_), .Y(men_men_n1333_));
  NA3        u1284(.A(men_men_n1333_), .B(men_men_n1332_), .C(men_men_n1331_), .Y(men_men_n1334_));
  NA2        u1285(.A(men_men_n1334_), .B(men_men_n421_), .Y(men_men_n1335_));
  AOI210     u1286(.A0(men_men_n376_), .A1(men_men_n338_), .B0(men_men_n55_), .Y(men_men_n1336_));
  NA4        u1287(.A(men_men_n1336_), .B(men_men_n1335_), .C(men_men_n1328_), .D(men_men_n1325_), .Y(men_men_n1337_));
  AO220      u1288(.A0(men_men_n1337_), .A1(men_men_n1306_), .B0(men_men_n1276_), .B1(men_men_n1270_), .Y(men16));
  NO2        u1289(.A(x4), .B(men_men_n59_), .Y(men_men_n1339_));
  NA2        u1290(.A(men_men_n646_), .B(men_men_n524_), .Y(men_men_n1340_));
  NA3        u1291(.A(men_men_n233_), .B(men_men_n427_), .C(men_men_n929_), .Y(men_men_n1341_));
  NA2        u1292(.A(men_men_n134_), .B(men_men_n210_), .Y(men_men_n1342_));
  AOI210     u1293(.A0(men_men_n1341_), .A1(men_men_n1340_), .B0(men_men_n1342_), .Y(men_men_n1343_));
  NO3        u1294(.A(x8), .B(x6), .C(men_men_n50_), .Y(men_men_n1344_));
  INV        u1295(.A(men_men_n188_), .Y(men_men_n1345_));
  OAI210     u1296(.A0(men_men_n1344_), .A1(men_men_n241_), .B0(men_men_n1345_), .Y(men_men_n1346_));
  NO2        u1297(.A(men_men_n162_), .B(x5), .Y(men_men_n1347_));
  NA2        u1298(.A(men_men_n1347_), .B(men_men_n1308_), .Y(men_men_n1348_));
  NA3        u1299(.A(men_men_n562_), .B(men_men_n526_), .C(men_men_n469_), .Y(men_men_n1349_));
  NA3        u1300(.A(men_men_n1349_), .B(men_men_n1348_), .C(men_men_n1346_), .Y(men_men_n1350_));
  OAI210     u1301(.A0(men_men_n1350_), .A1(men_men_n1343_), .B0(men_men_n1339_), .Y(men_men_n1351_));
  OAI210     u1302(.A0(men_men_n1224_), .A1(men_men_n903_), .B0(men_men_n418_), .Y(men_men_n1352_));
  NO2        u1303(.A(men_men_n318_), .B(x7), .Y(men_men_n1353_));
  NA2        u1304(.A(men_men_n1353_), .B(x0), .Y(men_men_n1354_));
  AOI210     u1305(.A0(men_men_n1354_), .A1(men_men_n1352_), .B0(men_men_n621_), .Y(men_men_n1355_));
  NA2        u1306(.A(men_men_n55_), .B(men_men_n107_), .Y(men_men_n1356_));
  NA2        u1307(.A(men_men_n375_), .B(men_men_n1039_), .Y(men_men_n1357_));
  OR2        u1308(.A(men_men_n1357_), .B(men_men_n55_), .Y(men_men_n1358_));
  OAI210     u1309(.A0(men_men_n1358_), .A1(men_men_n636_), .B0(men_men_n489_), .Y(men_men_n1359_));
  INV        u1310(.A(men_men_n980_), .Y(men_men_n1360_));
  NO2        u1311(.A(men_men_n1360_), .B(men_men_n62_), .Y(men_men_n1361_));
  AOI220     u1312(.A0(men_men_n1361_), .A1(men_men_n272_), .B0(men_men_n1209_), .B1(men_men_n127_), .Y(men_men_n1362_));
  AOI220     u1313(.A0(men_men_n620_), .A1(men_men_n360_), .B0(men_men_n607_), .B1(men_men_n88_), .Y(men_men_n1363_));
  NA3        u1314(.A(men_men_n458_), .B(men_men_n569_), .C(men_men_n195_), .Y(men_men_n1364_));
  OAI220     u1315(.A0(men_men_n1364_), .A1(men_men_n1363_), .B0(men_men_n1362_), .B1(men_men_n307_), .Y(men_men_n1365_));
  NO3        u1316(.A(men_men_n1365_), .B(men_men_n1359_), .C(men_men_n1355_), .Y(men_men_n1366_));
  NO3        u1317(.A(x6), .B(x4), .C(x3), .Y(men_men_n1367_));
  NA2        u1318(.A(men_men_n1367_), .B(men_men_n523_), .Y(men_men_n1368_));
  NA4        u1319(.A(men_men_n691_), .B(men_men_n188_), .C(men_men_n58_), .D(x6), .Y(men_men_n1369_));
  AOI210     u1320(.A0(men_men_n1369_), .A1(men_men_n1368_), .B0(men_men_n54_), .Y(men_men_n1370_));
  NO2        u1321(.A(men_men_n706_), .B(x3), .Y(men_men_n1371_));
  AOI210     u1322(.A0(men_men_n645_), .A1(men_men_n149_), .B0(men_men_n1021_), .Y(men_men_n1372_));
  OA210      u1323(.A0(men_men_n1371_), .A1(men_men_n421_), .B0(men_men_n1372_), .Y(men_men_n1373_));
  NO3        u1324(.A(men_men_n491_), .B(men_men_n222_), .C(men_men_n75_), .Y(men_men_n1374_));
  NO2        u1325(.A(men_men_n746_), .B(men_men_n500_), .Y(men_men_n1375_));
  NO3        u1326(.A(men_men_n1375_), .B(men_men_n262_), .C(men_men_n157_), .Y(men_men_n1376_));
  NO4        u1327(.A(men_men_n1376_), .B(men_men_n1374_), .C(men_men_n1373_), .D(men_men_n1370_), .Y(men_men_n1377_));
  NA2        u1328(.A(men_men_n404_), .B(men_men_n929_), .Y(men_men_n1378_));
  NA4        u1329(.A(men_men_n475_), .B(men_men_n368_), .C(men_men_n224_), .D(x6), .Y(men_men_n1379_));
  OAI210     u1330(.A0(men_men_n706_), .A1(men_men_n1378_), .B0(men_men_n1379_), .Y(men_men_n1380_));
  NA2        u1331(.A(men_men_n885_), .B(men_men_n1254_), .Y(men_men_n1381_));
  NA2        u1332(.A(men_men_n715_), .B(x7), .Y(men_men_n1382_));
  OAI210     u1333(.A0(men_men_n1382_), .A1(men_men_n387_), .B0(men_men_n1381_), .Y(men_men_n1383_));
  NA2        u1334(.A(men_men_n279_), .B(x2), .Y(men_men_n1384_));
  NO3        u1335(.A(men_men_n1384_), .B(men_men_n577_), .C(men_men_n72_), .Y(men_men_n1385_));
  OR2        u1336(.A(men_men_n1208_), .B(men_men_n58_), .Y(men_men_n1386_));
  AOI210     u1337(.A0(men_men_n562_), .A1(men_men_n50_), .B0(men_men_n572_), .Y(men_men_n1387_));
  OAI210     u1338(.A0(men_men_n904_), .A1(men_men_n920_), .B0(men_men_n382_), .Y(men_men_n1388_));
  OAI220     u1339(.A0(men_men_n1388_), .A1(men_men_n1387_), .B0(men_men_n1386_), .B1(men_men_n193_), .Y(men_men_n1389_));
  NO4        u1340(.A(men_men_n1389_), .B(men_men_n1385_), .C(men_men_n1383_), .D(men_men_n1380_), .Y(men_men_n1390_));
  OA220      u1341(.A0(men_men_n1390_), .A1(men_men_n439_), .B0(men_men_n1377_), .B1(men_men_n208_), .Y(men_men_n1391_));
  INV        u1342(.A(men_men_n415_), .Y(men_men_n1392_));
  NO3        u1343(.A(men_men_n930_), .B(men_men_n331_), .C(x8), .Y(men_men_n1393_));
  OAI210     u1344(.A0(men_men_n1393_), .A1(men_men_n415_), .B0(x6), .Y(men_men_n1394_));
  NA2        u1345(.A(men_men_n2550_), .B(men_men_n904_), .Y(men_men_n1395_));
  NA2        u1346(.A(men_men_n854_), .B(men_men_n71_), .Y(men_men_n1396_));
  AOI210     u1347(.A0(men_men_n491_), .A1(men_men_n57_), .B0(men_men_n615_), .Y(men_men_n1397_));
  NA3        u1348(.A(men_men_n230_), .B(men_men_n76_), .C(men_men_n71_), .Y(men_men_n1398_));
  OAI210     u1349(.A0(men_men_n895_), .A1(men_men_n233_), .B0(men_men_n1398_), .Y(men_men_n1399_));
  AOI210     u1350(.A0(men_men_n1397_), .A1(men_men_n2552_), .B0(men_men_n1399_), .Y(men_men_n1400_));
  NA3        u1351(.A(men_men_n1400_), .B(men_men_n1395_), .C(men_men_n1394_), .Y(men_men_n1401_));
  NO2        u1352(.A(men_men_n622_), .B(x6), .Y(men_men_n1402_));
  AN2        u1353(.A(men_men_n1402_), .B(men_men_n132_), .Y(men_men_n1403_));
  NO3        u1354(.A(men_men_n441_), .B(men_men_n385_), .C(x7), .Y(men_men_n1404_));
  NO3        u1355(.A(men_men_n162_), .B(men_men_n75_), .C(x2), .Y(men_men_n1405_));
  NO3        u1356(.A(men_men_n1405_), .B(men_men_n1404_), .C(men_men_n1403_), .Y(men_men_n1406_));
  NO2        u1357(.A(men_men_n233_), .B(x1), .Y(men_men_n1407_));
  OAI210     u1358(.A0(men_men_n1407_), .A1(men_men_n446_), .B0(men_men_n500_), .Y(men_men_n1408_));
  NO2        u1359(.A(men_men_n57_), .B(men_men_n107_), .Y(men_men_n1409_));
  NA2        u1360(.A(men_men_n1044_), .B(men_men_n1409_), .Y(men_men_n1410_));
  AOI210     u1361(.A0(men_men_n1410_), .A1(men_men_n1408_), .B0(men_men_n56_), .Y(men_men_n1411_));
  AOI220     u1362(.A0(men_men_n748_), .A1(men_men_n758_), .B0(men_men_n503_), .B1(men_men_n282_), .Y(men_men_n1412_));
  NO2        u1363(.A(men_men_n1412_), .B(men_men_n1254_), .Y(men_men_n1413_));
  NO3        u1364(.A(men_men_n523_), .B(men_men_n175_), .C(men_men_n1015_), .Y(men_men_n1414_));
  NA2        u1365(.A(men_men_n920_), .B(x4), .Y(men_men_n1415_));
  OAI220     u1366(.A0(men_men_n1415_), .A1(men_men_n672_), .B0(men_men_n630_), .B1(men_men_n593_), .Y(men_men_n1416_));
  NO4        u1367(.A(men_men_n1416_), .B(men_men_n1414_), .C(men_men_n1413_), .D(men_men_n1411_), .Y(men_men_n1417_));
  OAI210     u1368(.A0(men_men_n1406_), .A1(x5), .B0(men_men_n1417_), .Y(men_men_n1418_));
  AOI220     u1369(.A0(men_men_n1418_), .A1(men_men_n98_), .B0(men_men_n1401_), .B1(men_men_n338_), .Y(men_men_n1419_));
  NA4        u1370(.A(men_men_n1419_), .B(men_men_n1391_), .C(men_men_n1366_), .D(men_men_n1351_), .Y(men17));
  NO4        u1371(.A(men_men_n584_), .B(men_men_n685_), .C(men_men_n101_), .D(men_men_n100_), .Y(men_men_n1421_));
  NO2        u1372(.A(men_men_n125_), .B(men_men_n1118_), .Y(men_men_n1422_));
  AOI220     u1373(.A0(men_men_n1422_), .A1(men_men_n700_), .B0(men_men_n1421_), .B1(men_men_n494_), .Y(men_men_n1423_));
  NA2        u1374(.A(men_men_n166_), .B(men_men_n78_), .Y(men_men_n1424_));
  NOi21      u1375(.An(men_men_n380_), .B(men_men_n84_), .Y(men_men_n1425_));
  OAI210     u1376(.A0(men_men_n607_), .A1(men_men_n55_), .B0(men_men_n1425_), .Y(men_men_n1426_));
  NA2        u1377(.A(men_men_n1171_), .B(men_men_n976_), .Y(men_men_n1427_));
  NA4        u1378(.A(men_men_n1427_), .B(men_men_n1426_), .C(men_men_n718_), .D(men_men_n57_), .Y(men_men_n1428_));
  NA2        u1379(.A(x8), .B(men_men_n1254_), .Y(men_men_n1429_));
  NA3        u1380(.A(men_men_n1429_), .B(men_men_n1193_), .C(men_men_n397_), .Y(men_men_n1430_));
  NA2        u1381(.A(men_men_n393_), .B(men_men_n272_), .Y(men_men_n1431_));
  OA210      u1382(.A0(men_men_n1264_), .A1(men_men_n1112_), .B0(men_men_n738_), .Y(men_men_n1432_));
  NA4        u1383(.A(men_men_n1432_), .B(men_men_n1431_), .C(men_men_n1430_), .D(men_men_n1428_), .Y(men_men_n1433_));
  NA2        u1384(.A(men_men_n613_), .B(men_men_n1015_), .Y(men_men_n1434_));
  AOI210     u1385(.A0(men_men_n1041_), .A1(men_men_n303_), .B0(men_men_n59_), .Y(men_men_n1435_));
  NA2        u1386(.A(men_men_n1435_), .B(men_men_n1434_), .Y(men_men_n1436_));
  AOI210     u1387(.A0(men_men_n1433_), .A1(x1), .B0(men_men_n1436_), .Y(men_men_n1437_));
  NO2        u1388(.A(men_men_n947_), .B(men_men_n491_), .Y(men_men_n1438_));
  OAI210     u1389(.A0(men_men_n1438_), .A1(men_men_n1025_), .B0(men_men_n590_), .Y(men_men_n1439_));
  NO3        u1390(.A(men_men_n615_), .B(men_men_n541_), .C(men_men_n514_), .Y(men_men_n1440_));
  OAI210     u1391(.A0(men_men_n1440_), .A1(men_men_n884_), .B0(men_men_n1371_), .Y(men_men_n1441_));
  AOI210     u1392(.A0(men_men_n1441_), .A1(men_men_n1439_), .B0(x8), .Y(men_men_n1442_));
  NA3        u1393(.A(men_men_n615_), .B(men_men_n275_), .C(men_men_n122_), .Y(men_men_n1443_));
  NO2        u1394(.A(men_men_n145_), .B(men_men_n143_), .Y(men_men_n1444_));
  NO3        u1395(.A(men_men_n879_), .B(men_men_n758_), .C(men_men_n685_), .Y(men_men_n1445_));
  AOI210     u1396(.A0(men_men_n1445_), .A1(men_men_n1444_), .B0(x0), .Y(men_men_n1446_));
  OAI210     u1397(.A0(men_men_n1443_), .A1(men_men_n251_), .B0(men_men_n1446_), .Y(men_men_n1447_));
  NO2        u1398(.A(men_men_n1447_), .B(men_men_n1442_), .Y(men_men_n1448_));
  OAI220     u1399(.A0(men_men_n1448_), .A1(men_men_n1437_), .B0(men_men_n1424_), .B1(men_men_n1423_), .Y(men18));
  AOI210     u1400(.A0(x8), .A1(x0), .B0(x5), .Y(men_men_n1450_));
  NOi31      u1401(.An(men_men_n303_), .B(men_men_n1450_), .C(men_men_n1013_), .Y(men_men_n1451_));
  NA2        u1402(.A(men_men_n584_), .B(men_men_n59_), .Y(men_men_n1452_));
  NO2        u1403(.A(men_men_n349_), .B(men_men_n1452_), .Y(men_men_n1453_));
  NO2        u1404(.A(men_men_n600_), .B(men_men_n759_), .Y(men_men_n1454_));
  NO4        u1405(.A(men_men_n258_), .B(men_men_n796_), .C(men_men_n156_), .D(men_men_n70_), .Y(men_men_n1455_));
  NO4        u1406(.A(men_men_n1455_), .B(men_men_n1454_), .C(men_men_n1453_), .D(men_men_n1451_), .Y(men_men_n1456_));
  NO2        u1407(.A(men_men_n871_), .B(x5), .Y(men_men_n1457_));
  AOI210     u1408(.A0(men_men_n1099_), .A1(x5), .B0(men_men_n1457_), .Y(men_men_n1458_));
  OA220      u1409(.A0(men_men_n509_), .A1(men_men_n331_), .B0(men_men_n397_), .B1(x5), .Y(men_men_n1459_));
  OAI220     u1410(.A0(men_men_n1459_), .A1(men_men_n294_), .B0(men_men_n1458_), .B1(men_men_n216_), .Y(men_men_n1460_));
  AOI210     u1411(.A0(men_men_n386_), .A1(men_men_n293_), .B0(men_men_n1460_), .Y(men_men_n1461_));
  AOI210     u1412(.A0(men_men_n1461_), .A1(men_men_n1456_), .B0(x6), .Y(men_men_n1462_));
  NA3        u1413(.A(men_men_n513_), .B(men_men_n418_), .C(x2), .Y(men_men_n1463_));
  NA3        u1414(.A(men_men_n1013_), .B(men_men_n51_), .C(men_men_n57_), .Y(men_men_n1464_));
  AOI210     u1415(.A0(men_men_n1464_), .A1(men_men_n1463_), .B0(men_men_n773_), .Y(men_men_n1465_));
  AOI210     u1416(.A0(men_men_n422_), .A1(men_men_n139_), .B0(men_men_n771_), .Y(men_men_n1466_));
  NA2        u1417(.A(men_men_n272_), .B(x6), .Y(men_men_n1467_));
  OAI210     u1418(.A0(men_men_n181_), .A1(men_men_n109_), .B0(men_men_n1103_), .Y(men_men_n1468_));
  OAI220     u1419(.A0(men_men_n1468_), .A1(men_men_n1467_), .B0(men_men_n1466_), .B1(men_men_n730_), .Y(men_men_n1469_));
  OAI210     u1420(.A0(men_men_n1469_), .A1(men_men_n1465_), .B0(men_men_n53_), .Y(men_men_n1470_));
  NO2        u1421(.A(men_men_n268_), .B(x3), .Y(men_men_n1471_));
  AOI210     u1422(.A0(men_men_n1106_), .A1(men_men_n599_), .B0(x4), .Y(men_men_n1472_));
  OAI210     u1423(.A0(men_men_n541_), .A1(men_men_n584_), .B0(men_men_n59_), .Y(men_men_n1473_));
  OAI210     u1424(.A0(men_men_n607_), .A1(men_men_n632_), .B0(men_men_n1473_), .Y(men_men_n1474_));
  NA2        u1425(.A(men_men_n1474_), .B(men_men_n163_), .Y(men_men_n1475_));
  NA3        u1426(.A(men_men_n1475_), .B(men_men_n1472_), .C(men_men_n1470_), .Y(men_men_n1476_));
  NO3        u1427(.A(men_men_n1032_), .B(men_men_n132_), .C(men_men_n131_), .Y(men_men_n1477_));
  OAI210     u1428(.A0(men_men_n1477_), .A1(men_men_n637_), .B0(men_men_n107_), .Y(men_men_n1478_));
  NO2        u1429(.A(men_men_n1478_), .B(men_men_n773_), .Y(men_men_n1479_));
  NA3        u1430(.A(men_men_n1163_), .B(men_men_n193_), .C(men_men_n142_), .Y(men_men_n1480_));
  NA3        u1431(.A(men_men_n1035_), .B(men_men_n761_), .C(men_men_n342_), .Y(men_men_n1481_));
  INV        u1432(.A(men_men_n758_), .Y(men_men_n1482_));
  OAI210     u1433(.A0(men_men_n1482_), .A1(men_men_n1267_), .B0(men_men_n1481_), .Y(men_men_n1483_));
  AOI210     u1434(.A0(men_men_n1480_), .A1(men_men_n180_), .B0(men_men_n1483_), .Y(men_men_n1484_));
  OAI210     u1435(.A0(men_men_n1484_), .A1(men_men_n531_), .B0(x4), .Y(men_men_n1485_));
  OAI220     u1436(.A0(men_men_n1485_), .A1(men_men_n1479_), .B0(men_men_n1476_), .B1(men_men_n1462_), .Y(men_men_n1486_));
  NO2        u1437(.A(men_men_n148_), .B(men_men_n123_), .Y(men_men_n1487_));
  NO2        u1438(.A(men_men_n193_), .B(men_men_n788_), .Y(men_men_n1488_));
  AOI210     u1439(.A0(men_men_n585_), .A1(men_men_n500_), .B0(men_men_n1488_), .Y(men_men_n1489_));
  NO2        u1440(.A(men_men_n1489_), .B(x6), .Y(men_men_n1490_));
  NO2        u1441(.A(men_men_n385_), .B(men_men_n257_), .Y(men_men_n1491_));
  NO2        u1442(.A(men_men_n132_), .B(men_men_n720_), .Y(men_men_n1492_));
  NO2        u1443(.A(men_men_n930_), .B(men_men_n568_), .Y(men_men_n1493_));
  AO220      u1444(.A0(men_men_n1493_), .A1(men_men_n1492_), .B0(men_men_n1491_), .B1(men_men_n125_), .Y(men_men_n1494_));
  NO3        u1445(.A(men_men_n1494_), .B(men_men_n1490_), .C(men_men_n1487_), .Y(men_men_n1495_));
  NA2        u1446(.A(men_men_n1032_), .B(x3), .Y(men_men_n1496_));
  NA2        u1447(.A(men_men_n1303_), .B(men_men_n134_), .Y(men_men_n1497_));
  OAI220     u1448(.A0(men_men_n1497_), .A1(men_men_n1496_), .B0(men_men_n1495_), .B1(x3), .Y(men_men_n1498_));
  NO3        u1449(.A(men_men_n969_), .B(men_men_n671_), .C(men_men_n326_), .Y(men_men_n1499_));
  AO210      u1450(.A0(men_men_n993_), .A1(men_men_n298_), .B0(men_men_n1499_), .Y(men_men_n1500_));
  AOI220     u1451(.A0(men_men_n1500_), .A1(x8), .B0(men_men_n1303_), .B1(men_men_n432_), .Y(men_men_n1501_));
  NA2        u1452(.A(men_men_n734_), .B(men_men_n317_), .Y(men_men_n1502_));
  NO4        u1453(.A(men_men_n366_), .B(men_men_n206_), .C(men_men_n337_), .D(x2), .Y(men_men_n1503_));
  NA2        u1454(.A(men_men_n1356_), .B(men_men_n109_), .Y(men_men_n1504_));
  NO3        u1455(.A(men_men_n1165_), .B(men_men_n962_), .C(men_men_n1103_), .Y(men_men_n1505_));
  AOI210     u1456(.A0(men_men_n1505_), .A1(men_men_n1504_), .B0(men_men_n1503_), .Y(men_men_n1506_));
  OA220      u1457(.A0(men_men_n1506_), .A1(men_men_n930_), .B0(men_men_n1502_), .B1(men_men_n554_), .Y(men_men_n1507_));
  OAI210     u1458(.A0(men_men_n1501_), .A1(men_men_n407_), .B0(men_men_n1507_), .Y(men_men_n1508_));
  AOI210     u1459(.A0(men_men_n1498_), .A1(men_men_n139_), .B0(men_men_n1508_), .Y(men_men_n1509_));
  NA2        u1460(.A(men_men_n1509_), .B(men_men_n1486_), .Y(men19));
  NO2        u1461(.A(men_men_n1396_), .B(men_men_n261_), .Y(men_men_n1511_));
  NA2        u1462(.A(men_men_n632_), .B(x3), .Y(men_men_n1512_));
  OAI210     u1463(.A0(men_men_n156_), .A1(men_men_n108_), .B0(men_men_n81_), .Y(men_men_n1513_));
  NA3        u1464(.A(men_men_n1513_), .B(men_men_n1512_), .C(men_men_n244_), .Y(men_men_n1514_));
  NA2        u1465(.A(men_men_n1421_), .B(men_men_n352_), .Y(men_men_n1515_));
  AOI210     u1466(.A0(men_men_n1515_), .A1(men_men_n1514_), .B0(men_men_n56_), .Y(men_men_n1516_));
  INV        u1467(.A(men_men_n843_), .Y(men_men_n1517_));
  OAI210     u1468(.A0(men_men_n1516_), .A1(men_men_n1511_), .B0(men_men_n1517_), .Y(men_men_n1518_));
  NOi21      u1469(.An(men_men_n594_), .B(men_men_n636_), .Y(men_men_n1519_));
  AOI210     u1470(.A0(men_men_n352_), .A1(x6), .B0(men_men_n122_), .Y(men_men_n1520_));
  NO3        u1471(.A(men_men_n1520_), .B(men_men_n743_), .C(men_men_n127_), .Y(men_men_n1521_));
  NA2        u1472(.A(men_men_n1158_), .B(men_men_n123_), .Y(men_men_n1522_));
  NO4        u1473(.A(men_men_n1522_), .B(men_men_n969_), .C(men_men_n871_), .D(men_men_n77_), .Y(men_men_n1523_));
  NO2        u1474(.A(men_men_n1523_), .B(men_men_n1521_), .Y(men_men_n1524_));
  NO2        u1475(.A(men_men_n531_), .B(men_men_n603_), .Y(men_men_n1525_));
  NA2        u1476(.A(men_men_n1208_), .B(men_men_n50_), .Y(men_men_n1526_));
  NO3        u1477(.A(men_men_n507_), .B(men_men_n305_), .C(men_men_n64_), .Y(men_men_n1527_));
  AOI220     u1478(.A0(men_men_n1527_), .A1(men_men_n1526_), .B0(men_men_n1525_), .B1(men_men_n761_), .Y(men_men_n1528_));
  OAI210     u1479(.A0(men_men_n1524_), .A1(men_men_n57_), .B0(men_men_n1528_), .Y(men_men_n1529_));
  AOI210     u1480(.A0(men_men_n1529_), .A1(men_men_n758_), .B0(men_men_n1519_), .Y(men_men_n1530_));
  NA3        u1481(.A(men_men_n718_), .B(men_men_n260_), .C(x7), .Y(men_men_n1531_));
  AOI220     u1482(.A0(men_men_n1353_), .A1(men_men_n773_), .B0(men_men_n685_), .B1(men_men_n1118_), .Y(men_men_n1532_));
  AOI210     u1483(.A0(men_men_n1532_), .A1(men_men_n1531_), .B0(men_men_n492_), .Y(men_men_n1533_));
  NA2        u1484(.A(men_men_n1533_), .B(men_men_n796_), .Y(men_men_n1534_));
  NO2        u1485(.A(men_men_n730_), .B(men_men_n321_), .Y(men_men_n1535_));
  NO2        u1486(.A(men_men_n156_), .B(men_men_n990_), .Y(men_men_n1536_));
  AOI220     u1487(.A0(men_men_n1536_), .A1(men_men_n1224_), .B0(men_men_n1535_), .B1(men_men_n470_), .Y(men_men_n1537_));
  AO210      u1488(.A0(men_men_n1537_), .A1(men_men_n1534_), .B0(x1), .Y(men_men_n1538_));
  NA2        u1489(.A(men_men_n149_), .B(men_men_n110_), .Y(men_men_n1539_));
  NOi21      u1490(.An(x1), .B(x6), .Y(men_men_n1540_));
  NA2        u1491(.A(men_men_n1540_), .B(men_men_n84_), .Y(men_men_n1541_));
  NA2        u1492(.A(men_men_n1541_), .B(men_men_n1539_), .Y(men_men_n1542_));
  AOI220     u1493(.A0(men_men_n1542_), .A1(x3), .B0(men_men_n1166_), .B1(men_men_n381_), .Y(men_men_n1543_));
  NA3        u1494(.A(men_men_n1171_), .B(men_men_n783_), .C(men_men_n586_), .Y(men_men_n1544_));
  AOI220     u1495(.A0(men_men_n1212_), .A1(men_men_n122_), .B0(men_men_n899_), .B1(men_men_n798_), .Y(men_men_n1545_));
  AOI210     u1496(.A0(men_men_n1545_), .A1(men_men_n1544_), .B0(men_men_n321_), .Y(men_men_n1546_));
  NA2        u1497(.A(men_men_n920_), .B(men_men_n50_), .Y(men_men_n1547_));
  NA3        u1498(.A(men_men_n1158_), .B(men_men_n382_), .C(men_men_n109_), .Y(men_men_n1548_));
  AOI210     u1499(.A0(men_men_n1548_), .A1(men_men_n1547_), .B0(men_men_n938_), .Y(men_men_n1549_));
  NO3        u1500(.A(men_men_n601_), .B(men_men_n506_), .C(men_men_n1182_), .Y(men_men_n1550_));
  NO3        u1501(.A(men_men_n1550_), .B(men_men_n1549_), .C(men_men_n1546_), .Y(men_men_n1551_));
  OAI210     u1502(.A0(men_men_n1543_), .A1(men_men_n832_), .B0(men_men_n1551_), .Y(men_men_n1552_));
  NO2        u1503(.A(men_men_n54_), .B(men_men_n71_), .Y(men_men_n1553_));
  AO220      u1504(.A0(men_men_n1553_), .A1(men_men_n969_), .B0(men_men_n798_), .B1(men_men_n929_), .Y(men_men_n1554_));
  NA2        u1505(.A(men_men_n1141_), .B(men_men_n358_), .Y(men_men_n1555_));
  NO2        u1506(.A(men_men_n962_), .B(men_men_n1540_), .Y(men_men_n1556_));
  NA2        u1507(.A(men_men_n491_), .B(men_men_n715_), .Y(men_men_n1557_));
  OAI210     u1508(.A0(men_men_n1557_), .A1(men_men_n1556_), .B0(men_men_n1555_), .Y(men_men_n1558_));
  AOI210     u1509(.A0(men_men_n1554_), .A1(x2), .B0(men_men_n1558_), .Y(men_men_n1559_));
  NO2        u1510(.A(men_men_n1559_), .B(men_men_n156_), .Y(men_men_n1560_));
  OAI210     u1511(.A0(men_men_n1560_), .A1(men_men_n1552_), .B0(x8), .Y(men_men_n1561_));
  NA4        u1512(.A(men_men_n1561_), .B(men_men_n1538_), .C(men_men_n1530_), .D(men_men_n1518_), .Y(men20));
  NA4        u1513(.A(men_men_n392_), .B(men_men_n282_), .C(men_men_n380_), .D(men_men_n62_), .Y(men_men_n1563_));
  NA2        u1514(.A(men_men_n470_), .B(men_men_n411_), .Y(men_men_n1564_));
  AOI210     u1515(.A0(men_men_n1564_), .A1(men_men_n1563_), .B0(men_men_n87_), .Y(men_men_n1565_));
  AOI210     u1516(.A0(men_men_n1019_), .A1(men_men_n62_), .B0(men_men_n1525_), .Y(men_men_n1566_));
  AOI210     u1517(.A0(men_men_n956_), .A1(men_men_n348_), .B0(men_men_n1148_), .Y(men_men_n1567_));
  OAI210     u1518(.A0(men_men_n1566_), .A1(men_men_n667_), .B0(men_men_n1567_), .Y(men_men_n1568_));
  OAI210     u1519(.A0(men_men_n1568_), .A1(men_men_n1565_), .B0(men_men_n1067_), .Y(men_men_n1569_));
  NAi21      u1520(.An(men_men_n539_), .B(men_men_n399_), .Y(men_men_n1570_));
  NA3        u1521(.A(men_men_n1570_), .B(men_men_n954_), .C(men_men_n929_), .Y(men_men_n1571_));
  NO2        u1522(.A(men_men_n1571_), .B(men_men_n1254_), .Y(men_men_n1572_));
  NO2        u1523(.A(men_men_n734_), .B(men_men_n945_), .Y(men_men_n1573_));
  NOi31      u1524(.An(men_men_n1573_), .B(men_men_n1133_), .C(men_men_n519_), .Y(men_men_n1574_));
  OAI210     u1525(.A0(men_men_n1574_), .A1(men_men_n1572_), .B0(men_men_n326_), .Y(men_men_n1575_));
  NO4        u1526(.A(men_men_n535_), .B(men_men_n239_), .C(x5), .D(x2), .Y(men_men_n1576_));
  NA2        u1527(.A(men_men_n317_), .B(men_men_n92_), .Y(men_men_n1577_));
  NA2        u1528(.A(men_men_n327_), .B(men_men_n107_), .Y(men_men_n1578_));
  NA2        u1529(.A(men_men_n421_), .B(men_men_n52_), .Y(men_men_n1579_));
  OAI220     u1530(.A0(men_men_n1579_), .A1(men_men_n1578_), .B0(men_men_n1577_), .B1(men_men_n278_), .Y(men_men_n1580_));
  OAI210     u1531(.A0(men_men_n1580_), .A1(men_men_n1576_), .B0(men_men_n224_), .Y(men_men_n1581_));
  NO2        u1532(.A(men_men_n651_), .B(men_men_n590_), .Y(men_men_n1582_));
  NA2        u1533(.A(men_men_n930_), .B(men_men_n50_), .Y(men_men_n1583_));
  NO3        u1534(.A(men_men_n1583_), .B(men_men_n364_), .C(men_men_n232_), .Y(men_men_n1584_));
  NA3        u1535(.A(men_men_n338_), .B(men_men_n241_), .C(men_men_n64_), .Y(men_men_n1585_));
  OAI220     u1536(.A0(men_men_n1585_), .A1(men_men_n661_), .B0(men_men_n1415_), .B1(men_men_n1002_), .Y(men_men_n1586_));
  AOI210     u1537(.A0(men_men_n1584_), .A1(men_men_n1582_), .B0(men_men_n1586_), .Y(men_men_n1587_));
  NA4        u1538(.A(men_men_n1587_), .B(men_men_n1581_), .C(men_men_n1575_), .D(men_men_n1569_), .Y(men21));
  OAI210     u1539(.A0(men_men_n404_), .A1(men_men_n54_), .B0(x7), .Y(men_men_n1589_));
  OAI220     u1540(.A0(men_men_n1589_), .A1(men_men_n1243_), .B0(men_men_n1020_), .B1(men_men_n95_), .Y(men_men_n1590_));
  NA2        u1541(.A(men_men_n1590_), .B(men_men_n78_), .Y(men_men_n1591_));
  NA2        u1542(.A(men_men_n293_), .B(men_men_n841_), .Y(men_men_n1592_));
  NO2        u1543(.A(men_men_n307_), .B(men_men_n554_), .Y(men_men_n1593_));
  NA2        u1544(.A(men_men_n920_), .B(men_men_n277_), .Y(men_men_n1594_));
  NA2        u1545(.A(men_men_n527_), .B(men_men_n457_), .Y(men_men_n1595_));
  NA4        u1546(.A(men_men_n1595_), .B(men_men_n1594_), .C(men_men_n1332_), .D(men_men_n56_), .Y(men_men_n1596_));
  NO2        u1547(.A(men_men_n761_), .B(men_men_n431_), .Y(men_men_n1597_));
  NO3        u1548(.A(men_men_n1597_), .B(men_men_n707_), .C(men_men_n253_), .Y(men_men_n1598_));
  NOi31      u1549(.An(men_men_n196_), .B(men_men_n615_), .C(men_men_n1052_), .Y(men_men_n1599_));
  NO4        u1550(.A(men_men_n1599_), .B(men_men_n1598_), .C(men_men_n1596_), .D(men_men_n1593_), .Y(men_men_n1600_));
  NO2        u1551(.A(men_men_n431_), .B(men_men_n52_), .Y(men_men_n1601_));
  OA210      u1552(.A0(men_men_n1601_), .A1(men_men_n868_), .B0(x3), .Y(men_men_n1602_));
  OAI210     u1553(.A0(men_men_n772_), .A1(men_men_n572_), .B0(men_men_n340_), .Y(men_men_n1603_));
  NO2        u1554(.A(men_men_n70_), .B(x2), .Y(men_men_n1604_));
  OAI210     u1555(.A0(men_men_n180_), .A1(x0), .B0(men_men_n1604_), .Y(men_men_n1605_));
  NA2        u1556(.A(men_men_n146_), .B(men_men_n107_), .Y(men_men_n1606_));
  NA3        u1557(.A(men_men_n1606_), .B(men_men_n1605_), .C(men_men_n1603_), .Y(men_men_n1607_));
  OAI210     u1558(.A0(men_men_n1607_), .A1(men_men_n1602_), .B0(x8), .Y(men_men_n1608_));
  NO3        u1559(.A(men_men_n759_), .B(men_men_n604_), .C(men_men_n568_), .Y(men_men_n1609_));
  NA2        u1560(.A(men_men_n55_), .B(men_men_n50_), .Y(men_men_n1610_));
  OAI210     u1561(.A0(men_men_n628_), .A1(men_men_n567_), .B0(x4), .Y(men_men_n1611_));
  NO2        u1562(.A(men_men_n1611_), .B(men_men_n1609_), .Y(men_men_n1612_));
  AO220      u1563(.A0(men_men_n1612_), .A1(men_men_n1608_), .B0(men_men_n1600_), .B1(men_men_n1591_), .Y(men_men_n1613_));
  AO220      u1564(.A0(men_men_n616_), .A1(men_men_n321_), .B0(men_men_n573_), .B1(x8), .Y(men_men_n1614_));
  NO2        u1565(.A(men_men_n843_), .B(x0), .Y(men_men_n1615_));
  NO3        u1566(.A(men_men_n1615_), .B(men_men_n536_), .C(men_men_n88_), .Y(men_men_n1616_));
  NO2        u1567(.A(men_men_n162_), .B(x2), .Y(men_men_n1617_));
  NO3        u1568(.A(men_men_n377_), .B(men_men_n258_), .C(men_men_n188_), .Y(men_men_n1618_));
  AOI210     u1569(.A0(men_men_n1617_), .A1(men_men_n68_), .B0(men_men_n1618_), .Y(men_men_n1619_));
  OAI210     u1570(.A0(men_men_n1616_), .A1(men_men_n397_), .B0(men_men_n1619_), .Y(men_men_n1620_));
  AOI220     u1571(.A0(men_men_n1620_), .A1(x5), .B0(men_men_n1614_), .B1(men_men_n734_), .Y(men_men_n1621_));
  AOI210     u1572(.A0(men_men_n1621_), .A1(men_men_n1613_), .B0(men_men_n71_), .Y(men_men_n1622_));
  INV        u1573(.A(men_men_n889_), .Y(men_men_n1623_));
  NOi41      u1574(.An(men_men_n1384_), .B(men_men_n1450_), .C(men_men_n1117_), .D(men_men_n836_), .Y(men_men_n1624_));
  NA2        u1575(.A(men_men_n1624_), .B(men_men_n1623_), .Y(men_men_n1625_));
  NO2        u1576(.A(men_men_n78_), .B(x4), .Y(men_men_n1626_));
  OAI210     u1577(.A0(men_men_n291_), .A1(men_men_n160_), .B0(men_men_n1626_), .Y(men_men_n1627_));
  OAI210     u1578(.A0(men_men_n406_), .A1(men_men_n422_), .B0(men_men_n232_), .Y(men_men_n1628_));
  NO2        u1579(.A(men_men_n260_), .B(men_men_n50_), .Y(men_men_n1629_));
  NO2        u1580(.A(men_men_n1629_), .B(men_men_n57_), .Y(men_men_n1630_));
  NA2        u1581(.A(men_men_n1630_), .B(men_men_n1628_), .Y(men_men_n1631_));
  AOI210     u1582(.A0(men_men_n1627_), .A1(men_men_n1625_), .B0(men_men_n1631_), .Y(men_men_n1632_));
  NA2        u1583(.A(men_men_n746_), .B(men_men_n539_), .Y(men_men_n1633_));
  AO210      u1584(.A0(men_men_n1633_), .A1(men_men_n938_), .B0(men_men_n50_), .Y(men_men_n1634_));
  NO2        u1585(.A(men_men_n1570_), .B(men_men_n1176_), .Y(men_men_n1635_));
  AOI220     u1586(.A0(men_men_n1635_), .A1(men_men_n1126_), .B0(men_men_n1280_), .B1(men_men_n1013_), .Y(men_men_n1636_));
  AOI210     u1587(.A0(men_men_n1636_), .A1(men_men_n1634_), .B0(men_men_n109_), .Y(men_men_n1637_));
  NA2        u1588(.A(men_men_n298_), .B(men_men_n107_), .Y(men_men_n1638_));
  NA2        u1589(.A(men_men_n876_), .B(men_men_n55_), .Y(men_men_n1639_));
  NO2        u1590(.A(men_men_n1639_), .B(men_men_n1638_), .Y(men_men_n1640_));
  NO3        u1591(.A(men_men_n1640_), .B(men_men_n1637_), .C(men_men_n1632_), .Y(men_men_n1641_));
  NO2        u1592(.A(men_men_n1641_), .B(x6), .Y(men_men_n1642_));
  AOI210     u1593(.A0(men_men_n593_), .A1(men_men_n1021_), .B0(men_men_n1450_), .Y(men_men_n1643_));
  OAI210     u1594(.A0(men_men_n1643_), .A1(men_men_n674_), .B0(men_men_n56_), .Y(men_men_n1644_));
  NO2        u1595(.A(men_men_n736_), .B(men_men_n54_), .Y(men_men_n1645_));
  NO4        u1596(.A(men_men_n936_), .B(men_men_n281_), .C(men_men_n758_), .D(men_men_n743_), .Y(men_men_n1646_));
  NO2        u1597(.A(men_men_n848_), .B(x5), .Y(men_men_n1647_));
  NO4        u1598(.A(men_men_n1647_), .B(men_men_n1646_), .C(men_men_n1645_), .D(men_men_n926_), .Y(men_men_n1648_));
  AOI210     u1599(.A0(men_men_n1648_), .A1(men_men_n1644_), .B0(men_men_n50_), .Y(men_men_n1649_));
  NA2        u1600(.A(men_men_n162_), .B(men_men_n107_), .Y(men_men_n1650_));
  OA220      u1601(.A0(men_men_n1650_), .A1(men_men_n435_), .B0(men_men_n462_), .B1(men_men_n734_), .Y(men_men_n1651_));
  NA3        u1602(.A(men_men_n55_), .B(x2), .C(x0), .Y(men_men_n1652_));
  AOI220     u1603(.A0(men_men_n1652_), .A1(men_men_n173_), .B0(men_men_n848_), .B1(men_men_n158_), .Y(men_men_n1653_));
  NO2        u1604(.A(men_men_n667_), .B(men_men_n260_), .Y(men_men_n1654_));
  NO3        u1605(.A(men_men_n248_), .B(men_men_n230_), .C(men_men_n358_), .Y(men_men_n1655_));
  NO3        u1606(.A(men_men_n1655_), .B(men_men_n1654_), .C(men_men_n1653_), .Y(men_men_n1656_));
  OAI220     u1607(.A0(men_men_n1656_), .A1(men_men_n56_), .B0(men_men_n1651_), .B1(men_men_n683_), .Y(men_men_n1657_));
  OAI210     u1608(.A0(men_men_n1657_), .A1(men_men_n1649_), .B0(men_men_n115_), .Y(men_men_n1658_));
  NO2        u1609(.A(men_men_n598_), .B(men_men_n302_), .Y(men_men_n1659_));
  AOI210     u1610(.A0(men_men_n591_), .A1(x5), .B0(men_men_n1659_), .Y(men_men_n1660_));
  NO2        u1611(.A(men_men_n1660_), .B(men_men_n109_), .Y(men_men_n1661_));
  NA2        u1612(.A(men_men_n691_), .B(men_men_n81_), .Y(men_men_n1662_));
  NA3        u1613(.A(men_men_n1662_), .B(men_men_n428_), .C(men_men_n57_), .Y(men_men_n1663_));
  OAI210     u1614(.A0(men_men_n1639_), .A1(men_men_n1638_), .B0(men_men_n1663_), .Y(men_men_n1664_));
  OAI210     u1615(.A0(men_men_n1664_), .A1(men_men_n1661_), .B0(x1), .Y(men_men_n1665_));
  NO4        u1616(.A(men_men_n415_), .B(men_men_n78_), .C(men_men_n150_), .D(x3), .Y(men_men_n1666_));
  NO2        u1617(.A(men_men_n327_), .B(men_men_n111_), .Y(men_men_n1667_));
  OAI210     u1618(.A0(men_men_n1666_), .A1(men_men_n1255_), .B0(men_men_n1667_), .Y(men_men_n1668_));
  NO2        u1619(.A(men_men_n60_), .B(men_men_n107_), .Y(men_men_n1669_));
  NO4        u1620(.A(men_men_n1638_), .B(men_men_n936_), .C(men_men_n651_), .D(men_men_n50_), .Y(men_men_n1670_));
  AOI210     u1621(.A0(men_men_n1669_), .A1(men_men_n1488_), .B0(men_men_n1670_), .Y(men_men_n1671_));
  NA4        u1622(.A(men_men_n1671_), .B(men_men_n1668_), .C(men_men_n1665_), .D(men_men_n1658_), .Y(men_men_n1672_));
  NO3        u1623(.A(men_men_n1672_), .B(men_men_n1642_), .C(men_men_n1622_), .Y(men22));
  AOI210     u1624(.A0(men_men_n513_), .A1(men_men_n71_), .B0(men_men_n464_), .Y(men_men_n1674_));
  NO3        u1625(.A(men_men_n1153_), .B(men_men_n541_), .C(men_men_n685_), .Y(men_men_n1675_));
  AOI210     u1626(.A0(x5), .A1(x2), .B0(x8), .Y(men_men_n1676_));
  NA2        u1627(.A(men_men_n1676_), .B(men_men_n59_), .Y(men_men_n1677_));
  OAI220     u1628(.A0(men_men_n1677_), .A1(men_men_n1675_), .B0(men_men_n1674_), .B1(men_men_n397_), .Y(men_men_n1678_));
  NA2        u1629(.A(men_men_n567_), .B(men_men_n87_), .Y(men_men_n1679_));
  NA2        u1630(.A(men_men_n278_), .B(men_men_n77_), .Y(men_men_n1680_));
  OA220      u1631(.A0(men_men_n1680_), .A1(men_men_n1679_), .B0(men_men_n829_), .B1(men_men_n976_), .Y(men_men_n1681_));
  NO4        u1632(.A(men_men_n385_), .B(men_men_n222_), .C(men_men_n71_), .D(x3), .Y(men_men_n1682_));
  NO3        u1633(.A(men_men_n1203_), .B(men_men_n87_), .C(x0), .Y(men_men_n1683_));
  OAI210     u1634(.A0(men_men_n397_), .A1(men_men_n208_), .B0(x4), .Y(men_men_n1684_));
  NO3        u1635(.A(men_men_n1684_), .B(men_men_n1683_), .C(men_men_n1682_), .Y(men_men_n1685_));
  OAI210     u1636(.A0(men_men_n1681_), .A1(men_men_n201_), .B0(men_men_n1685_), .Y(men_men_n1686_));
  AOI210     u1637(.A0(men_men_n1678_), .A1(men_men_n53_), .B0(men_men_n1686_), .Y(men_men_n1687_));
  NA2        u1638(.A(men_men_n300_), .B(men_men_n305_), .Y(men_men_n1688_));
  NA3        u1639(.A(men_men_n1688_), .B(men_men_n224_), .C(men_men_n304_), .Y(men_men_n1689_));
  NA2        u1640(.A(men_men_n562_), .B(men_men_n247_), .Y(men_men_n1690_));
  NO3        u1641(.A(men_men_n491_), .B(men_men_n268_), .C(men_men_n216_), .Y(men_men_n1691_));
  NAi31      u1642(.An(men_men_n1691_), .B(men_men_n1690_), .C(men_men_n1689_), .Y(men_men_n1692_));
  NO2        u1643(.A(men_men_n462_), .B(men_men_n262_), .Y(men_men_n1693_));
  NO2        u1644(.A(men_men_n1203_), .B(x3), .Y(men_men_n1694_));
  AOI210     u1645(.A0(men_men_n1694_), .A1(men_men_n348_), .B0(men_men_n1693_), .Y(men_men_n1695_));
  OAI210     u1646(.A0(men_men_n1050_), .A1(men_men_n190_), .B0(men_men_n56_), .Y(men_men_n1696_));
  NA3        u1647(.A(men_men_n55_), .B(men_men_n71_), .C(x0), .Y(men_men_n1697_));
  NO2        u1648(.A(men_men_n1697_), .B(men_men_n1021_), .Y(men_men_n1698_));
  NO2        u1649(.A(men_men_n1698_), .B(men_men_n1696_), .Y(men_men_n1699_));
  OAI210     u1650(.A0(men_men_n1695_), .A1(men_men_n260_), .B0(men_men_n1699_), .Y(men_men_n1700_));
  AOI210     u1651(.A0(men_men_n1692_), .A1(men_men_n107_), .B0(men_men_n1700_), .Y(men_men_n1701_));
  AOI210     u1652(.A0(men_men_n928_), .A1(men_men_n760_), .B0(men_men_n852_), .Y(men_men_n1702_));
  NO2        u1653(.A(men_men_n790_), .B(men_men_n162_), .Y(men_men_n1703_));
  OAI210     u1654(.A0(men_men_n1703_), .A1(men_men_n1702_), .B0(men_men_n597_), .Y(men_men_n1704_));
  OA210      u1655(.A0(men_men_n1701_), .A1(men_men_n1687_), .B0(men_men_n1704_), .Y(men_men_n1705_));
  NA2        u1656(.A(men_men_n690_), .B(men_men_n678_), .Y(men_men_n1706_));
  NO2        u1657(.A(men_men_n353_), .B(x0), .Y(men_men_n1707_));
  NA3        u1658(.A(men_men_n1707_), .B(men_men_n348_), .C(men_men_n56_), .Y(men_men_n1708_));
  AOI210     u1659(.A0(men_men_n1708_), .A1(men_men_n1706_), .B0(men_men_n397_), .Y(men_men_n1709_));
  NA2        u1660(.A(men_men_n417_), .B(men_men_n109_), .Y(men_men_n1710_));
  NA2        u1661(.A(men_men_n142_), .B(men_men_n773_), .Y(men_men_n1711_));
  NA2        u1662(.A(men_men_n415_), .B(x3), .Y(men_men_n1712_));
  NAi31      u1663(.An(men_men_n1712_), .B(men_men_n1711_), .C(men_men_n1504_), .Y(men_men_n1713_));
  NO3        u1664(.A(men_men_n843_), .B(men_men_n461_), .C(men_men_n109_), .Y(men_men_n1714_));
  NO2        u1665(.A(men_men_n1051_), .B(men_men_n143_), .Y(men_men_n1715_));
  NO3        u1666(.A(men_men_n879_), .B(men_men_n411_), .C(men_men_n301_), .Y(men_men_n1716_));
  AOI220     u1667(.A0(men_men_n1716_), .A1(men_men_n1715_), .B0(men_men_n1714_), .B1(men_men_n1707_), .Y(men_men_n1717_));
  NA3        u1668(.A(men_men_n411_), .B(men_men_n92_), .C(men_men_n81_), .Y(men_men_n1718_));
  AOI210     u1669(.A0(men_men_n593_), .A1(men_men_n451_), .B0(men_men_n488_), .Y(men_men_n1719_));
  NA2        u1670(.A(men_men_n1137_), .B(x3), .Y(men_men_n1720_));
  OAI210     u1671(.A0(men_men_n1720_), .A1(men_men_n1719_), .B0(men_men_n1718_), .Y(men_men_n1721_));
  NA3        u1672(.A(men_men_n56_), .B(men_men_n50_), .C(x0), .Y(men_men_n1722_));
  NOi21      u1673(.An(men_men_n83_), .B(men_men_n718_), .Y(men_men_n1723_));
  NA3        u1674(.A(x6), .B(x4), .C(men_men_n50_), .Y(men_men_n1724_));
  NA3        u1675(.A(men_men_n1724_), .B(men_men_n962_), .C(men_men_n269_), .Y(men_men_n1725_));
  OAI220     u1676(.A0(men_men_n1725_), .A1(men_men_n1723_), .B0(men_men_n1024_), .B1(men_men_n1722_), .Y(men_men_n1726_));
  AOI220     u1677(.A0(men_men_n1726_), .A1(men_men_n1035_), .B0(men_men_n1721_), .B1(men_men_n348_), .Y(men_men_n1727_));
  NA4        u1678(.A(men_men_n1727_), .B(men_men_n1717_), .C(men_men_n1713_), .D(men_men_n1710_), .Y(men_men_n1728_));
  AOI210     u1679(.A0(men_men_n1728_), .A1(x7), .B0(men_men_n1709_), .Y(men_men_n1729_));
  OAI210     u1680(.A0(men_men_n1705_), .A1(x7), .B0(men_men_n1729_), .Y(men23));
  NA2        u1681(.A(men_men_n224_), .B(men_men_n1573_), .Y(men_men_n1731_));
  NO3        u1682(.A(men_men_n829_), .B(men_men_n576_), .C(men_men_n481_), .Y(men_men_n1732_));
  NO3        u1683(.A(men_men_n931_), .B(men_men_n151_), .C(men_men_n116_), .Y(men_men_n1733_));
  AOI210     u1684(.A0(men_men_n1733_), .A1(men_men_n996_), .B0(men_men_n1732_), .Y(men_men_n1734_));
  OAI210     u1685(.A0(men_men_n1731_), .A1(men_men_n156_), .B0(men_men_n1734_), .Y(men_men_n1735_));
  NA2        u1686(.A(men_men_n1735_), .B(men_men_n55_), .Y(men_men_n1736_));
  NO2        u1687(.A(men_men_n936_), .B(men_men_n505_), .Y(men_men_n1737_));
  AO220      u1688(.A0(men_men_n1239_), .A1(men_men_n184_), .B0(men_men_n969_), .B1(men_men_n734_), .Y(men_men_n1738_));
  OAI210     u1689(.A0(men_men_n1738_), .A1(men_men_n1737_), .B0(men_men_n573_), .Y(men_men_n1739_));
  NA2        u1690(.A(men_men_n181_), .B(men_men_n171_), .Y(men_men_n1740_));
  NA2        u1691(.A(men_men_n403_), .B(men_men_n163_), .Y(men_men_n1741_));
  AOI210     u1692(.A0(men_men_n1741_), .A1(men_men_n1740_), .B0(men_men_n239_), .Y(men_men_n1742_));
  NA3        u1693(.A(men_men_n852_), .B(men_men_n422_), .C(men_men_n260_), .Y(men_men_n1743_));
  NO2        u1694(.A(men_men_n1743_), .B(men_men_n382_), .Y(men_men_n1744_));
  OAI210     u1695(.A0(men_men_n1744_), .A1(men_men_n1742_), .B0(men_men_n298_), .Y(men_men_n1745_));
  NA3        u1696(.A(men_men_n57_), .B(x4), .C(x3), .Y(men_men_n1746_));
  NO3        u1697(.A(men_men_n1746_), .B(men_men_n731_), .C(men_men_n142_), .Y(men_men_n1747_));
  AOI210     u1698(.A0(men_men_n903_), .A1(men_men_n144_), .B0(men_men_n1747_), .Y(men_men_n1748_));
  NA4        u1699(.A(men_men_n1748_), .B(men_men_n1745_), .C(men_men_n1739_), .D(men_men_n1736_), .Y(men24));
  NO2        u1700(.A(men_men_n244_), .B(x1), .Y(men_men_n1750_));
  NA2        u1701(.A(men_men_n338_), .B(men_men_n485_), .Y(men_men_n1751_));
  NAi21      u1702(.An(men_men_n1750_), .B(men_men_n1751_), .Y(men_men_n1752_));
  NO3        u1703(.A(men_men_n531_), .B(men_men_n670_), .C(men_men_n158_), .Y(men_men_n1753_));
  AOI210     u1704(.A0(men_men_n1752_), .A1(men_men_n92_), .B0(men_men_n1753_), .Y(men_men_n1754_));
  NA2        u1705(.A(men_men_n101_), .B(x8), .Y(men_men_n1755_));
  NO2        u1706(.A(men_men_n1032_), .B(men_men_n1294_), .Y(men_men_n1756_));
  AOI210     u1707(.A0(men_men_n954_), .A1(men_men_n56_), .B0(men_men_n1402_), .Y(men_men_n1757_));
  AO220      u1708(.A0(men_men_n1757_), .A1(men_men_n1756_), .B0(men_men_n1226_), .B1(men_men_n326_), .Y(men_men_n1758_));
  NA2        u1709(.A(men_men_n451_), .B(x8), .Y(men_men_n1759_));
  NA2        u1710(.A(men_men_n652_), .B(men_men_n125_), .Y(men_men_n1760_));
  OAI220     u1711(.A0(men_men_n1760_), .A1(men_men_n1392_), .B0(men_men_n1759_), .B1(men_men_n827_), .Y(men_men_n1761_));
  AOI220     u1712(.A0(men_men_n1761_), .A1(men_men_n1629_), .B0(men_men_n1758_), .B1(men_men_n996_), .Y(men_men_n1762_));
  OAI210     u1713(.A0(men_men_n1755_), .A1(men_men_n1754_), .B0(men_men_n1762_), .Y(men25));
  NA2        u1714(.A(men_men_n327_), .B(men_men_n59_), .Y(men_men_n1764_));
  NO2        u1715(.A(men_men_n1764_), .B(men_men_n318_), .Y(men_men_n1765_));
  OAI210     u1716(.A0(men_men_n1765_), .A1(men_men_n1142_), .B0(men_men_n115_), .Y(men_men_n1766_));
  INV        u1717(.A(men_men_n1234_), .Y(men_men_n1767_));
  NO2        u1718(.A(men_men_n730_), .B(men_men_n55_), .Y(men_men_n1768_));
  AOI220     u1719(.A0(men_men_n1768_), .A1(men_men_n1767_), .B0(men_men_n1535_), .B1(men_men_n1143_), .Y(men_men_n1769_));
  AOI210     u1720(.A0(men_men_n1769_), .A1(men_men_n1766_), .B0(men_men_n665_), .Y(men_men_n1770_));
  NO3        u1721(.A(men_men_n1008_), .B(men_men_n145_), .C(men_men_n78_), .Y(men_men_n1771_));
  OAI210     u1722(.A0(men_men_n201_), .A1(men_men_n278_), .B0(men_men_n328_), .Y(men_men_n1772_));
  OAI210     u1723(.A0(men_men_n1772_), .A1(men_men_n1771_), .B0(men_men_n1141_), .Y(men_men_n1773_));
  NO2        u1724(.A(men_men_n1344_), .B(men_men_n445_), .Y(men_men_n1774_));
  NO3        u1725(.A(men_men_n1774_), .B(men_men_n523_), .C(men_men_n98_), .Y(men_men_n1775_));
  NA2        u1726(.A(men_men_n500_), .B(men_men_n55_), .Y(men_men_n1776_));
  OAI220     u1727(.A0(men_men_n1776_), .A1(men_men_n244_), .B0(men_men_n570_), .B1(men_men_n278_), .Y(men_men_n1777_));
  OAI210     u1728(.A0(men_men_n1777_), .A1(men_men_n1775_), .B0(men_men_n620_), .Y(men_men_n1778_));
  AOI220     u1729(.A0(men_men_n1693_), .A1(men_men_n1099_), .B0(men_men_n1444_), .B1(men_men_n378_), .Y(men_men_n1779_));
  NA3        u1730(.A(men_men_n1779_), .B(men_men_n1778_), .C(men_men_n1773_), .Y(men_men_n1780_));
  AO210      u1731(.A0(men_men_n1780_), .A1(men_men_n107_), .B0(men_men_n1770_), .Y(men26));
  NA2        u1732(.A(men_men_n758_), .B(men_men_n50_), .Y(men_men_n1782_));
  OAI220     u1733(.A0(men_men_n302_), .A1(men_men_n253_), .B0(men_men_n1782_), .B1(x7), .Y(men_men_n1783_));
  AOI220     u1734(.A0(men_men_n1783_), .A1(men_men_n92_), .B0(men_men_n1255_), .B1(men_men_n1103_), .Y(men_men_n1784_));
  NA2        u1735(.A(men_men_n608_), .B(men_men_n562_), .Y(men_men_n1785_));
  OAI210     u1736(.A0(men_men_n616_), .A1(men_men_n608_), .B0(men_men_n734_), .Y(men_men_n1786_));
  AOI210     u1737(.A0(men_men_n1785_), .A1(men_men_n1165_), .B0(men_men_n1786_), .Y(men_men_n1787_));
  NA2        u1738(.A(men_men_n988_), .B(men_men_n568_), .Y(men_men_n1788_));
  NO2        u1739(.A(men_men_n1788_), .B(men_men_n1208_), .Y(men_men_n1789_));
  AOI210     u1740(.A0(men_men_n1715_), .A1(men_men_n1409_), .B0(men_men_n1789_), .Y(men_men_n1790_));
  NO2        u1741(.A(men_men_n1051_), .B(men_men_n75_), .Y(men_men_n1791_));
  NA2        u1742(.A(men_men_n796_), .B(men_men_n180_), .Y(men_men_n1792_));
  NO2        u1743(.A(men_men_n1792_), .B(men_men_n528_), .Y(men_men_n1793_));
  AOI210     u1744(.A0(men_men_n1791_), .A1(men_men_n569_), .B0(men_men_n1793_), .Y(men_men_n1794_));
  OAI220     u1745(.A0(men_men_n1794_), .A1(men_men_n107_), .B0(men_men_n1790_), .B1(men_men_n53_), .Y(men_men_n1795_));
  NA2        u1746(.A(men_men_n585_), .B(men_men_n500_), .Y(men_men_n1796_));
  NO2        u1747(.A(men_men_n135_), .B(men_men_n132_), .Y(men_men_n1797_));
  NA2        u1748(.A(men_men_n1797_), .B(men_men_n122_), .Y(men_men_n1798_));
  NA2        u1749(.A(men_men_n734_), .B(x3), .Y(men_men_n1799_));
  AOI210     u1750(.A0(men_men_n1798_), .A1(men_men_n1796_), .B0(men_men_n1799_), .Y(men_men_n1800_));
  NA2        u1751(.A(men_men_n443_), .B(men_men_n107_), .Y(men_men_n1801_));
  NA3        u1752(.A(men_men_n555_), .B(men_men_n51_), .C(men_men_n56_), .Y(men_men_n1802_));
  AOI210     u1753(.A0(men_men_n1582_), .A1(men_men_n1025_), .B0(x0), .Y(men_men_n1803_));
  OAI210     u1754(.A0(men_men_n1802_), .A1(men_men_n1801_), .B0(men_men_n1803_), .Y(men_men_n1804_));
  NO4        u1755(.A(men_men_n1804_), .B(men_men_n1800_), .C(men_men_n1795_), .D(men_men_n1787_), .Y(men_men_n1805_));
  AOI210     u1756(.A0(x8), .A1(x6), .B0(x5), .Y(men_men_n1806_));
  AO220      u1757(.A0(men_men_n1806_), .A1(men_men_n147_), .B0(men_men_n576_), .B1(men_men_n142_), .Y(men_men_n1807_));
  NA2        u1758(.A(men_men_n1807_), .B(men_men_n444_), .Y(men_men_n1808_));
  NO2        u1759(.A(men_men_n744_), .B(men_men_n147_), .Y(men_men_n1809_));
  NA3        u1760(.A(men_men_n1809_), .B(men_men_n1604_), .C(men_men_n136_), .Y(men_men_n1810_));
  NO2        u1761(.A(men_men_n397_), .B(men_men_n1330_), .Y(men_men_n1811_));
  OAI210     u1762(.A0(men_men_n1811_), .A1(men_men_n1300_), .B0(men_men_n443_), .Y(men_men_n1812_));
  NA3        u1763(.A(men_men_n372_), .B(men_men_n841_), .C(men_men_n257_), .Y(men_men_n1813_));
  NA4        u1764(.A(men_men_n1813_), .B(men_men_n1812_), .C(men_men_n1810_), .D(men_men_n1808_), .Y(men_men_n1814_));
  AOI210     u1765(.A0(men_men_n226_), .A1(x2), .B0(men_men_n486_), .Y(men_men_n1815_));
  NO2        u1766(.A(men_men_n1815_), .B(men_men_n116_), .Y(men_men_n1816_));
  OAI220     u1767(.A0(men_men_n882_), .A1(men_men_n302_), .B0(men_men_n628_), .B1(men_men_n670_), .Y(men_men_n1817_));
  NO2        u1768(.A(men_men_n1817_), .B(men_men_n1816_), .Y(men_men_n1818_));
  NA3        u1769(.A(men_men_n652_), .B(men_men_n195_), .C(men_men_n929_), .Y(men_men_n1819_));
  NA2        u1770(.A(men_men_n1819_), .B(men_men_n628_), .Y(men_men_n1820_));
  INV        u1771(.A(men_men_n134_), .Y(men_men_n1821_));
  OAI210     u1772(.A0(men_men_n1821_), .A1(men_men_n1379_), .B0(x0), .Y(men_men_n1822_));
  AOI210     u1773(.A0(men_men_n1820_), .A1(men_men_n1367_), .B0(men_men_n1822_), .Y(men_men_n1823_));
  OAI210     u1774(.A0(men_men_n1818_), .A1(men_men_n53_), .B0(men_men_n1823_), .Y(men_men_n1824_));
  AOI210     u1775(.A0(men_men_n1814_), .A1(x4), .B0(men_men_n1824_), .Y(men_men_n1825_));
  OA220      u1776(.A0(men_men_n1825_), .A1(men_men_n1805_), .B0(men_men_n1784_), .B1(men_men_n108_), .Y(men27));
  NA2        u1777(.A(men_men_n1107_), .B(men_men_n443_), .Y(men_men_n1827_));
  NO2        u1778(.A(men_men_n1827_), .B(men_men_n299_), .Y(men_men_n1828_));
  NA3        u1779(.A(men_men_n804_), .B(men_men_n361_), .C(men_men_n990_), .Y(men_men_n1829_));
  NO2        u1780(.A(men_men_n1829_), .B(men_men_n218_), .Y(men_men_n1830_));
  OAI210     u1781(.A0(men_men_n1830_), .A1(men_men_n1828_), .B0(men_men_n686_), .Y(men_men_n1831_));
  XO2        u1782(.A(x8), .B(x4), .Y(men_men_n1832_));
  AN2        u1783(.A(men_men_n1209_), .B(men_men_n281_), .Y(men_men_n1833_));
  NO2        u1784(.A(men_men_n394_), .B(men_men_n167_), .Y(men_men_n1834_));
  OAI210     u1785(.A0(men_men_n1834_), .A1(men_men_n1833_), .B0(men_men_n1083_), .Y(men_men_n1835_));
  AOI210     u1786(.A0(men_men_n616_), .A1(men_men_n56_), .B0(men_men_n1791_), .Y(men_men_n1836_));
  OAI220     u1787(.A0(men_men_n1836_), .A1(men_men_n1208_), .B0(men_men_n1163_), .B1(men_men_n210_), .Y(men_men_n1837_));
  NO2        u1788(.A(men_men_n683_), .B(men_men_n145_), .Y(men_men_n1838_));
  NO2        u1789(.A(men_men_n1147_), .B(men_men_n260_), .Y(men_men_n1839_));
  AOI220     u1790(.A0(men_men_n1839_), .A1(men_men_n1838_), .B0(men_men_n1837_), .B1(men_men_n527_), .Y(men_men_n1840_));
  NA3        u1791(.A(men_men_n1840_), .B(men_men_n1835_), .C(men_men_n1831_), .Y(men28));
  NO3        u1792(.A(men_men_n1832_), .B(men_men_n1339_), .C(men_men_n149_), .Y(men_men_n1842_));
  OAI210     u1793(.A0(men_men_n1842_), .A1(men_men_n1227_), .B0(men_men_n568_), .Y(men_men_n1843_));
  NA3        u1794(.A(men_men_n1143_), .B(men_men_n876_), .C(x7), .Y(men_men_n1844_));
  NA3        u1795(.A(men_men_n488_), .B(men_men_n78_), .C(men_men_n590_), .Y(men_men_n1845_));
  NA3        u1796(.A(men_men_n1845_), .B(men_men_n1844_), .C(men_men_n1843_), .Y(men_men_n1846_));
  NA2        u1797(.A(men_men_n1203_), .B(men_men_n441_), .Y(men_men_n1847_));
  NA3        u1798(.A(men_men_n1847_), .B(men_men_n55_), .C(men_men_n410_), .Y(men_men_n1848_));
  NA2        u1799(.A(men_men_n1084_), .B(men_men_n660_), .Y(men_men_n1849_));
  NA2        u1800(.A(men_men_n1849_), .B(men_men_n1848_), .Y(men_men_n1850_));
  NO4        u1801(.A(x6), .B(men_men_n56_), .C(x2), .D(x0), .Y(men_men_n1851_));
  NA2        u1802(.A(men_men_n1851_), .B(men_men_n1013_), .Y(men_men_n1852_));
  NA2        u1803(.A(men_men_n1137_), .B(men_men_n107_), .Y(men_men_n1853_));
  INV        u1804(.A(men_men_n1049_), .Y(men_men_n1854_));
  OAI210     u1805(.A0(men_men_n1854_), .A1(men_men_n1853_), .B0(men_men_n1852_), .Y(men_men_n1855_));
  OAI210     u1806(.A0(men_men_n1855_), .A1(men_men_n1850_), .B0(x7), .Y(men_men_n1856_));
  NO2        u1807(.A(men_men_n385_), .B(x7), .Y(men_men_n1857_));
  NO3        u1808(.A(men_men_n397_), .B(men_men_n275_), .C(men_men_n123_), .Y(men_men_n1858_));
  OAI210     u1809(.A0(men_men_n852_), .A1(men_men_n262_), .B0(men_men_n81_), .Y(men_men_n1859_));
  OAI220     u1810(.A0(men_men_n1859_), .A1(men_men_n1858_), .B0(men_men_n1857_), .B1(men_men_n110_), .Y(men_men_n1860_));
  NA2        u1811(.A(men_men_n1724_), .B(men_men_n640_), .Y(men_men_n1861_));
  NO2        u1812(.A(men_men_n1776_), .B(men_men_n77_), .Y(men_men_n1862_));
  AOI220     u1813(.A0(men_men_n1862_), .A1(men_men_n1861_), .B0(men_men_n471_), .B1(men_men_n50_), .Y(men_men_n1863_));
  AOI210     u1814(.A0(men_men_n1863_), .A1(men_men_n1860_), .B0(men_men_n59_), .Y(men_men_n1864_));
  AOI220     u1815(.A0(men_men_n1344_), .A1(men_men_n658_), .B0(men_men_n409_), .B1(men_men_n451_), .Y(men_men_n1865_));
  OAI210     u1816(.A0(men_men_n1865_), .A1(men_men_n145_), .B0(x1), .Y(men_men_n1866_));
  NO2        u1817(.A(men_men_n1866_), .B(men_men_n1864_), .Y(men_men_n1867_));
  AOI210     u1818(.A0(men_men_n1522_), .A1(men_men_n397_), .B0(men_men_n650_), .Y(men_men_n1868_));
  NO2        u1819(.A(men_men_n397_), .B(x5), .Y(men_men_n1869_));
  NO2        u1820(.A(men_men_n1869_), .B(men_men_n230_), .Y(men_men_n1870_));
  NO2        u1821(.A(men_men_n1870_), .B(men_men_n1868_), .Y(men_men_n1871_));
  NOi21      u1822(.An(men_men_n691_), .B(men_men_n969_), .Y(men_men_n1872_));
  NA3        u1823(.A(men_men_n1872_), .B(men_men_n1049_), .C(men_men_n852_), .Y(men_men_n1873_));
  OAI210     u1824(.A0(men_men_n1314_), .A1(men_men_n1610_), .B0(men_men_n1873_), .Y(men_men_n1874_));
  OAI210     u1825(.A0(men_men_n1874_), .A1(men_men_n1871_), .B0(men_men_n1083_), .Y(men_men_n1875_));
  OAI210     u1826(.A0(men_men_n441_), .A1(men_men_n51_), .B0(men_men_n984_), .Y(men_men_n1876_));
  AOI220     u1827(.A0(men_men_n1876_), .A1(men_men_n457_), .B0(men_men_n441_), .B1(men_men_n386_), .Y(men_men_n1877_));
  NO2        u1828(.A(men_men_n1877_), .B(men_men_n156_), .Y(men_men_n1878_));
  NA2        u1829(.A(men_men_n165_), .B(men_men_n71_), .Y(men_men_n1879_));
  OAI210     u1830(.A0(men_men_n1788_), .A1(men_men_n1879_), .B0(men_men_n53_), .Y(men_men_n1880_));
  OAI220     u1831(.A0(men_men_n671_), .A1(men_men_n265_), .B0(men_men_n667_), .B1(x6), .Y(men_men_n1881_));
  NO2        u1832(.A(men_men_n300_), .B(x4), .Y(men_men_n1882_));
  AOI220     u1833(.A0(men_men_n1882_), .A1(men_men_n361_), .B0(men_men_n1881_), .B1(x4), .Y(men_men_n1883_));
  NO3        u1834(.A(men_men_n1883_), .B(men_men_n321_), .C(x5), .Y(men_men_n1884_));
  NO2        u1835(.A(men_men_n691_), .B(men_men_n57_), .Y(men_men_n1885_));
  OAI210     u1836(.A0(men_men_n1885_), .A1(men_men_n1838_), .B0(men_men_n443_), .Y(men_men_n1886_));
  AOI220     u1837(.A0(men_men_n648_), .A1(men_men_n720_), .B0(men_men_n486_), .B1(men_men_n240_), .Y(men_men_n1887_));
  AOI210     u1838(.A0(men_men_n1887_), .A1(men_men_n1886_), .B0(men_men_n260_), .Y(men_men_n1888_));
  NO4        u1839(.A(men_men_n1888_), .B(men_men_n1884_), .C(men_men_n1880_), .D(men_men_n1878_), .Y(men_men_n1889_));
  AOI220     u1840(.A0(men_men_n1889_), .A1(men_men_n1875_), .B0(men_men_n1867_), .B1(men_men_n1856_), .Y(men_men_n1890_));
  AOI210     u1841(.A0(men_men_n1846_), .A1(x3), .B0(men_men_n1890_), .Y(men29));
  NA2        u1842(.A(men_men_n736_), .B(men_men_n1013_), .Y(men_men_n1892_));
  AO210      u1843(.A0(men_men_n1119_), .A1(men_men_n1127_), .B0(men_men_n1892_), .Y(men_men_n1893_));
  AOI210     u1844(.A0(men_men_n185_), .A1(men_men_n169_), .B0(men_men_n691_), .Y(men_men_n1894_));
  AOI210     u1845(.A0(men_men_n1371_), .A1(men_men_n78_), .B0(men_men_n1894_), .Y(men_men_n1895_));
  NA2        u1846(.A(men_men_n1895_), .B(men_men_n1893_), .Y(men_men_n1896_));
  NO3        u1847(.A(men_men_n650_), .B(men_men_n1103_), .C(men_men_n50_), .Y(men_men_n1897_));
  NO3        u1848(.A(men_men_n1897_), .B(men_men_n1202_), .C(men_men_n542_), .Y(men_men_n1898_));
  NO2        u1849(.A(men_men_n439_), .B(men_men_n58_), .Y(men_men_n1899_));
  NA2        u1850(.A(men_men_n1899_), .B(men_men_n1165_), .Y(men_men_n1900_));
  OAI210     u1851(.A0(men_men_n1898_), .A1(men_men_n531_), .B0(men_men_n1900_), .Y(men_men_n1901_));
  AOI210     u1852(.A0(men_men_n1896_), .A1(x6), .B0(men_men_n1901_), .Y(men_men_n1902_));
  OAI210     u1853(.A0(x8), .A1(x4), .B0(x5), .Y(men_men_n1903_));
  NA2        u1854(.A(men_men_n1903_), .B(men_men_n111_), .Y(men_men_n1904_));
  NA2        u1855(.A(men_men_n300_), .B(men_men_n149_), .Y(men_men_n1905_));
  NA4        u1856(.A(men_men_n1905_), .B(men_men_n1904_), .C(men_men_n649_), .D(men_men_n64_), .Y(men_men_n1906_));
  AOI210     u1857(.A0(men_men_n1273_), .A1(men_men_n275_), .B0(men_men_n1659_), .Y(men_men_n1907_));
  AOI210     u1858(.A0(men_men_n1907_), .A1(men_men_n1906_), .B0(men_men_n871_), .Y(men_men_n1908_));
  NA3        u1859(.A(men_men_n650_), .B(men_men_n305_), .C(men_men_n169_), .Y(men_men_n1909_));
  NA3        u1860(.A(men_men_n614_), .B(men_men_n296_), .C(men_men_n788_), .Y(men_men_n1910_));
  AOI210     u1861(.A0(men_men_n1910_), .A1(men_men_n1909_), .B0(men_men_n1165_), .Y(men_men_n1911_));
  OAI210     u1862(.A0(men_men_n876_), .A1(x8), .B0(x7), .Y(men_men_n1912_));
  NO2        u1863(.A(men_men_n1912_), .B(men_men_n128_), .Y(men_men_n1913_));
  OAI220     u1864(.A0(men_men_n1903_), .A1(men_men_n570_), .B0(men_men_n1452_), .B1(men_men_n394_), .Y(men_men_n1914_));
  NO4        u1865(.A(men_men_n1914_), .B(men_men_n1913_), .C(men_men_n1911_), .D(men_men_n1908_), .Y(men_men_n1915_));
  OAI210     u1866(.A0(men_men_n1902_), .A1(x2), .B0(men_men_n1915_), .Y(men_men_n1916_));
  NA3        u1867(.A(x6), .B(men_men_n50_), .C(x2), .Y(men_men_n1917_));
  OAI210     u1868(.A0(men_men_n1182_), .A1(men_men_n352_), .B0(men_men_n1917_), .Y(men_men_n1918_));
  NO3        u1869(.A(men_men_n441_), .B(x3), .C(x0), .Y(men_men_n1919_));
  AO220      u1870(.A0(men_men_n1919_), .A1(x5), .B0(men_men_n1851_), .B1(men_men_n81_), .Y(men_men_n1920_));
  AOI210     u1871(.A0(men_men_n1918_), .A1(men_men_n342_), .B0(men_men_n1920_), .Y(men_men_n1921_));
  NO3        u1872(.A(men_men_n684_), .B(men_men_n362_), .C(men_men_n143_), .Y(men_men_n1922_));
  AOI210     u1873(.A0(men_men_n714_), .A1(men_men_n597_), .B0(men_men_n1922_), .Y(men_men_n1923_));
  OAI210     u1874(.A0(men_men_n1921_), .A1(x7), .B0(men_men_n1923_), .Y(men_men_n1924_));
  AOI210     u1875(.A0(men_men_n1053_), .A1(men_men_n397_), .B0(men_men_n1356_), .Y(men_men_n1925_));
  NO2        u1876(.A(men_men_n149_), .B(x2), .Y(men_men_n1926_));
  OA210      u1877(.A0(men_men_n1926_), .A1(men_men_n612_), .B0(men_men_n650_), .Y(men_men_n1927_));
  OAI210     u1878(.A0(men_men_n1927_), .A1(men_men_n1925_), .B0(men_men_n68_), .Y(men_men_n1928_));
  NO2        u1879(.A(men_men_n201_), .B(men_men_n85_), .Y(men_men_n1929_));
  OAI210     u1880(.A0(men_men_n1929_), .A1(men_men_n774_), .B0(men_men_n1062_), .Y(men_men_n1930_));
  NA3        u1881(.A(men_men_n1869_), .B(men_men_n233_), .C(men_men_n83_), .Y(men_men_n1931_));
  NA3        u1882(.A(men_men_n1931_), .B(men_men_n1930_), .C(men_men_n1928_), .Y(men_men_n1932_));
  AOI210     u1883(.A0(men_men_n1924_), .A1(x8), .B0(men_men_n1932_), .Y(men_men_n1933_));
  OAI210     u1884(.A0(men_men_n439_), .A1(men_men_n249_), .B0(men_men_n938_), .Y(men_men_n1934_));
  OAI210     u1885(.A0(men_men_n1934_), .A1(men_men_n1084_), .B0(men_men_n660_), .Y(men_men_n1935_));
  NO2        u1886(.A(men_men_n136_), .B(men_men_n92_), .Y(men_men_n1936_));
  NA2        u1887(.A(men_men_n1936_), .B(men_men_n571_), .Y(men_men_n1937_));
  NA2        u1888(.A(men_men_n175_), .B(x4), .Y(men_men_n1938_));
  NO3        u1889(.A(men_men_n1425_), .B(men_men_n244_), .C(men_men_n71_), .Y(men_men_n1939_));
  NA2        u1890(.A(men_men_n1939_), .B(men_men_n1938_), .Y(men_men_n1940_));
  NA3        u1891(.A(men_men_n1940_), .B(men_men_n1937_), .C(men_men_n1935_), .Y(men_men_n1941_));
  NO4        u1892(.A(men_men_n1158_), .B(men_men_n492_), .C(men_men_n1329_), .D(men_men_n107_), .Y(men_men_n1942_));
  NA2        u1893(.A(men_men_n1942_), .B(men_men_n109_), .Y(men_men_n1943_));
  AOI210     u1894(.A0(men_men_n304_), .A1(x4), .B0(men_men_n195_), .Y(men_men_n1944_));
  NA2        u1895(.A(men_men_n1944_), .B(men_men_n709_), .Y(men_men_n1945_));
  OR3        u1896(.A(men_men_n1680_), .B(men_men_n1382_), .C(men_men_n1050_), .Y(men_men_n1946_));
  NA2        u1897(.A(men_men_n1851_), .B(men_men_n795_), .Y(men_men_n1947_));
  OA220      u1898(.A0(men_men_n1947_), .A1(men_men_n249_), .B0(men_men_n563_), .B1(men_men_n1722_), .Y(men_men_n1948_));
  NA4        u1899(.A(men_men_n1948_), .B(men_men_n1946_), .C(men_men_n1945_), .D(men_men_n1943_), .Y(men_men_n1949_));
  AOI210     u1900(.A0(men_men_n1941_), .A1(men_men_n293_), .B0(men_men_n1949_), .Y(men_men_n1950_));
  OAI210     u1901(.A0(men_men_n1933_), .A1(x1), .B0(men_men_n1950_), .Y(men_men_n1951_));
  AO210      u1902(.A0(men_men_n1916_), .A1(x1), .B0(men_men_n1951_), .Y(men30));
  NO3        u1903(.A(men_men_n1707_), .B(men_men_n559_), .C(men_men_n98_), .Y(men_men_n1953_));
  NO3        u1904(.A(men_men_n1101_), .B(men_men_n139_), .C(men_men_n382_), .Y(men_men_n1954_));
  NO2        u1905(.A(men_men_n709_), .B(men_men_n1954_), .Y(men_men_n1955_));
  AOI210     u1906(.A0(men_men_n1955_), .A1(men_men_n1953_), .B0(men_men_n56_), .Y(men_men_n1956_));
  NA2        u1907(.A(men_men_n798_), .B(men_men_n340_), .Y(men_men_n1957_));
  NA2        u1908(.A(men_men_n1957_), .B(men_men_n1315_), .Y(men_men_n1958_));
  OAI210     u1909(.A0(men_men_n1958_), .A1(men_men_n1956_), .B0(men_men_n109_), .Y(men_men_n1959_));
  NA2        u1910(.A(men_men_n969_), .B(men_men_n660_), .Y(men_men_n1960_));
  AOI220     u1911(.A0(men_men_n444_), .A1(men_men_n920_), .B0(men_men_n326_), .B1(men_men_n451_), .Y(men_men_n1961_));
  AOI210     u1912(.A0(men_men_n1961_), .A1(men_men_n1960_), .B0(men_men_n260_), .Y(men_men_n1962_));
  NO3        u1913(.A(men_men_n283_), .B(men_men_n124_), .C(x0), .Y(men_men_n1963_));
  AOI210     u1914(.A0(men_men_n494_), .A1(x6), .B0(men_men_n1963_), .Y(men_men_n1964_));
  AOI220     u1915(.A0(men_men_n1099_), .A1(men_men_n421_), .B0(men_men_n748_), .B1(men_men_n91_), .Y(men_men_n1965_));
  OAI220     u1916(.A0(men_men_n1965_), .A1(men_men_n249_), .B0(men_men_n1964_), .B1(men_men_n54_), .Y(men_men_n1966_));
  NA3        u1917(.A(men_men_n322_), .B(men_men_n166_), .C(men_men_n71_), .Y(men_men_n1967_));
  AO210      u1918(.A0(men_men_n554_), .A1(men_men_n508_), .B0(x5), .Y(men_men_n1968_));
  AOI210     u1919(.A0(men_men_n1967_), .A1(men_men_n706_), .B0(men_men_n1968_), .Y(men_men_n1969_));
  AOI210     u1920(.A0(men_men_n1540_), .A1(men_men_n50_), .B0(men_men_n451_), .Y(men_men_n1970_));
  NA2        u1921(.A(men_men_n200_), .B(x2), .Y(men_men_n1971_));
  OA220      u1922(.A0(men_men_n1971_), .A1(men_men_n1970_), .B0(men_men_n279_), .B1(x6), .Y(men_men_n1972_));
  OAI210     u1923(.A0(x7), .A1(x6), .B0(x1), .Y(men_men_n1973_));
  NA3        u1924(.A(men_men_n57_), .B(x4), .C(men_men_n59_), .Y(men_men_n1974_));
  AOI220     u1925(.A0(men_men_n1974_), .A1(men_men_n1322_), .B0(men_men_n1973_), .B1(men_men_n1746_), .Y(men_men_n1975_));
  NO3        u1926(.A(men_men_n1318_), .B(men_men_n342_), .C(men_men_n990_), .Y(men_men_n1976_));
  NO2        u1927(.A(men_men_n506_), .B(men_men_n845_), .Y(men_men_n1977_));
  NOi21      u1928(.An(men_men_n1977_), .B(men_men_n832_), .Y(men_men_n1978_));
  NO3        u1929(.A(men_men_n1254_), .B(men_men_n235_), .C(men_men_n632_), .Y(men_men_n1979_));
  NO4        u1930(.A(men_men_n1979_), .B(men_men_n1978_), .C(men_men_n1976_), .D(men_men_n1975_), .Y(men_men_n1980_));
  OAI210     u1931(.A0(men_men_n1972_), .A1(men_men_n743_), .B0(men_men_n1980_), .Y(men_men_n1981_));
  NO4        u1932(.A(men_men_n1981_), .B(men_men_n1969_), .C(men_men_n1966_), .D(men_men_n1962_), .Y(men_men_n1982_));
  AOI210     u1933(.A0(men_men_n1982_), .A1(men_men_n1959_), .B0(x8), .Y(men_men_n1983_));
  NO3        u1934(.A(men_men_n484_), .B(men_men_n771_), .C(men_men_n53_), .Y(men_men_n1984_));
  OAI220     u1935(.A0(men_men_n1722_), .A1(men_men_n342_), .B0(men_men_n477_), .B1(men_men_n567_), .Y(men_men_n1985_));
  OAI210     u1936(.A0(men_men_n1985_), .A1(men_men_n1984_), .B0(x6), .Y(men_men_n1986_));
  OAI210     u1937(.A0(men_men_n1004_), .A1(men_men_n527_), .B0(men_men_n798_), .Y(men_men_n1987_));
  OAI210     u1938(.A0(men_men_n1669_), .A1(men_men_n329_), .B0(men_men_n127_), .Y(men_men_n1988_));
  AOI210     u1939(.A0(men_men_n377_), .A1(men_men_n232_), .B0(men_men_n72_), .Y(men_men_n1989_));
  AOI210     u1940(.A0(men_men_n969_), .A1(men_men_n734_), .B0(men_men_n1989_), .Y(men_men_n1990_));
  NA4        u1941(.A(men_men_n1990_), .B(men_men_n1988_), .C(men_men_n1987_), .D(men_men_n1986_), .Y(men_men_n1991_));
  NA2        u1942(.A(men_men_n1052_), .B(men_men_n59_), .Y(men_men_n1992_));
  NO2        u1943(.A(men_men_n1992_), .B(men_men_n476_), .Y(men_men_n1993_));
  AOI210     u1944(.A0(men_men_n1991_), .A1(x8), .B0(men_men_n1993_), .Y(men_men_n1994_));
  NO2        u1945(.A(men_men_n1994_), .B(men_men_n57_), .Y(men_men_n1995_));
  NA2        u1946(.A(men_men_n431_), .B(men_men_n832_), .Y(men_men_n1996_));
  NO2        u1947(.A(men_men_n903_), .B(men_men_n646_), .Y(men_men_n1997_));
  AOI210     u1948(.A0(men_men_n1997_), .A1(men_men_n1996_), .B0(men_men_n441_), .Y(men_men_n1998_));
  NO2        u1949(.A(men_men_n406_), .B(men_men_n1101_), .Y(men_men_n1999_));
  NO2        u1950(.A(men_men_n1999_), .B(men_men_n1208_), .Y(men_men_n2000_));
  AOI210     u1951(.A0(men_men_n301_), .A1(x1), .B0(men_men_n150_), .Y(men_men_n2001_));
  NO2        u1952(.A(men_men_n307_), .B(x5), .Y(men_men_n2002_));
  NO2        u1953(.A(men_men_n2002_), .B(men_men_n838_), .Y(men_men_n2003_));
  OAI220     u1954(.A0(men_men_n2003_), .A1(men_men_n1022_), .B0(men_men_n2001_), .B1(men_men_n210_), .Y(men_men_n2004_));
  NO3        u1955(.A(men_men_n2004_), .B(men_men_n2000_), .C(men_men_n1998_), .Y(men_men_n2005_));
  NA2        u1956(.A(men_men_n936_), .B(men_men_n82_), .Y(men_men_n2006_));
  AO210      u1957(.A0(men_men_n2006_), .A1(men_men_n1541_), .B0(x3), .Y(men_men_n2007_));
  NO2        u1958(.A(men_men_n221_), .B(men_men_n56_), .Y(men_men_n2008_));
  OAI220     u1959(.A0(men_men_n377_), .A1(men_men_n1208_), .B0(men_men_n353_), .B1(men_men_n235_), .Y(men_men_n2009_));
  AOI220     u1960(.A0(men_men_n2009_), .A1(x2), .B0(men_men_n2008_), .B1(men_men_n1553_), .Y(men_men_n2010_));
  AOI210     u1961(.A0(men_men_n2010_), .A1(men_men_n2007_), .B0(men_men_n265_), .Y(men_men_n2011_));
  NO2        u1962(.A(men_men_n301_), .B(men_men_n123_), .Y(men_men_n2012_));
  NO3        u1963(.A(men_men_n803_), .B(men_men_n685_), .C(men_men_n169_), .Y(men_men_n2013_));
  OAI210     u1964(.A0(men_men_n2013_), .A1(men_men_n2012_), .B0(men_men_n157_), .Y(men_men_n2014_));
  NA3        u1965(.A(x5), .B(x4), .C(men_men_n59_), .Y(men_men_n2015_));
  AOI210     u1966(.A0(men_men_n2015_), .A1(men_men_n1262_), .B0(men_men_n528_), .Y(men_men_n2016_));
  AOI210     u1967(.A0(men_men_n1280_), .A1(x2), .B0(men_men_n2016_), .Y(men_men_n2017_));
  AOI210     u1968(.A0(men_men_n2017_), .A1(men_men_n2014_), .B0(men_men_n50_), .Y(men_men_n2018_));
  NA3        u1969(.A(men_men_n1422_), .B(men_men_n1094_), .C(men_men_n469_), .Y(men_men_n2019_));
  AOI210     u1970(.A0(men_men_n2019_), .A1(men_men_n2006_), .B0(men_men_n593_), .Y(men_men_n2020_));
  AOI210     u1971(.A0(men_men_n990_), .A1(x1), .B0(men_men_n1273_), .Y(men_men_n2021_));
  OAI220     u1972(.A0(men_men_n305_), .A1(x4), .B0(men_men_n51_), .B1(x6), .Y(men_men_n2022_));
  NO2        u1973(.A(men_men_n122_), .B(men_men_n111_), .Y(men_men_n2023_));
  AOI220     u1974(.A0(men_men_n2023_), .A1(men_men_n2022_), .B0(men_men_n1121_), .B1(men_men_n607_), .Y(men_men_n2024_));
  OAI210     u1975(.A0(men_men_n2021_), .A1(men_men_n480_), .B0(men_men_n2024_), .Y(men_men_n2025_));
  NO4        u1976(.A(men_men_n2025_), .B(men_men_n2020_), .C(men_men_n2018_), .D(men_men_n2011_), .Y(men_men_n2026_));
  OAI210     u1977(.A0(men_men_n2005_), .A1(men_men_n136_), .B0(men_men_n2026_), .Y(men_men_n2027_));
  NO3        u1978(.A(men_men_n2027_), .B(men_men_n1995_), .C(men_men_n1983_), .Y(men31));
  NA2        u1979(.A(men_men_n954_), .B(men_men_n354_), .Y(men_men_n2029_));
  NO2        u1980(.A(men_men_n445_), .B(men_men_n660_), .Y(men_men_n2030_));
  AOI210     u1981(.A0(men_men_n2030_), .A1(men_men_n2029_), .B0(men_men_n58_), .Y(men_men_n2031_));
  NO2        u1982(.A(men_men_n773_), .B(men_men_n56_), .Y(men_men_n2032_));
  NA2        u1983(.A(men_men_n1947_), .B(men_men_n1785_), .Y(men_men_n2033_));
  OAI210     u1984(.A0(men_men_n2033_), .A1(men_men_n2031_), .B0(men_men_n53_), .Y(men_men_n2034_));
  NO2        u1985(.A(men_men_n428_), .B(men_men_n660_), .Y(men_men_n2035_));
  NO3        u1986(.A(men_men_n1882_), .B(men_men_n1851_), .C(men_men_n872_), .Y(men_men_n2036_));
  OA220      u1987(.A0(men_men_n2036_), .A1(men_men_n469_), .B0(men_men_n2035_), .B1(men_men_n1415_), .Y(men_men_n2037_));
  AOI210     u1988(.A0(men_men_n2037_), .A1(men_men_n2034_), .B0(men_men_n107_), .Y(men_men_n2038_));
  NO2        u1989(.A(men_men_n491_), .B(men_men_n75_), .Y(men_men_n2039_));
  NA2        u1990(.A(men_men_n441_), .B(men_men_n57_), .Y(men_men_n2040_));
  AOI210     u1991(.A0(men_men_n304_), .A1(men_men_n86_), .B0(men_men_n2040_), .Y(men_men_n2041_));
  OAI210     u1992(.A0(men_men_n2041_), .A1(men_men_n2039_), .B0(men_men_n758_), .Y(men_men_n2042_));
  NO4        u1993(.A(men_men_n1117_), .B(men_men_n362_), .C(men_men_n1540_), .D(men_men_n67_), .Y(men_men_n2043_));
  AOI210     u1994(.A0(men_men_n1577_), .A1(men_men_n1307_), .B0(men_men_n439_), .Y(men_men_n2044_));
  NO2        u1995(.A(men_men_n760_), .B(men_men_n116_), .Y(men_men_n2045_));
  NO3        u1996(.A(men_men_n2045_), .B(men_men_n2044_), .C(men_men_n2043_), .Y(men_men_n2046_));
  AOI210     u1997(.A0(men_men_n2046_), .A1(men_men_n2042_), .B0(x5), .Y(men_men_n2047_));
  NO2        u1998(.A(men_men_n563_), .B(men_men_n1182_), .Y(men_men_n2048_));
  AOI220     u1999(.A0(men_men_n937_), .A1(men_men_n720_), .B0(men_men_n1101_), .B1(men_men_n121_), .Y(men_men_n2049_));
  OAI220     u2000(.A0(men_men_n2049_), .A1(men_men_n385_), .B0(men_men_n476_), .B1(men_men_n759_), .Y(men_men_n2050_));
  NO4        u2001(.A(men_men_n2050_), .B(men_men_n2048_), .C(men_men_n2047_), .D(men_men_n2038_), .Y(men_men_n2051_));
  NO2        u2002(.A(men_men_n531_), .B(men_men_n142_), .Y(men_men_n2052_));
  OAI210     u2003(.A0(men_men_n103_), .A1(men_men_n278_), .B0(men_men_n1992_), .Y(men_men_n2053_));
  OAI210     u2004(.A0(men_men_n2053_), .A1(men_men_n2052_), .B0(x7), .Y(men_men_n2054_));
  NO3        u2005(.A(men_men_n377_), .B(men_men_n55_), .C(x7), .Y(men_men_n2055_));
  OA210      u2006(.A0(men_men_n2055_), .A1(men_men_n1272_), .B0(men_men_n100_), .Y(men_men_n2056_));
  NA2        u2007(.A(men_men_n1051_), .B(men_men_n91_), .Y(men_men_n2057_));
  AOI210     u2008(.A0(men_men_n882_), .A1(men_men_n111_), .B0(men_men_n2057_), .Y(men_men_n2058_));
  NA2        u2009(.A(men_men_n1491_), .B(x6), .Y(men_men_n2059_));
  AOI210     u2010(.A0(men_men_n2059_), .A1(men_men_n292_), .B0(men_men_n107_), .Y(men_men_n2060_));
  NA2        u2011(.A(men_men_n1143_), .B(men_men_n317_), .Y(men_men_n2061_));
  AOI210     u2012(.A0(men_men_n2061_), .A1(men_men_n628_), .B0(men_men_n53_), .Y(men_men_n2062_));
  NO4        u2013(.A(men_men_n2062_), .B(men_men_n2060_), .C(men_men_n2058_), .D(men_men_n2056_), .Y(men_men_n2063_));
  AOI210     u2014(.A0(men_men_n2063_), .A1(men_men_n2054_), .B0(men_men_n670_), .Y(men_men_n2064_));
  NOi21      u2015(.An(men_men_n1697_), .B(men_men_n1026_), .Y(men_men_n2065_));
  NO2        u2016(.A(men_men_n2065_), .B(men_men_n1853_), .Y(men_men_n2066_));
  NA2        u2017(.A(men_men_n2066_), .B(x3), .Y(men_men_n2067_));
  AOI220     u2018(.A0(men_men_n597_), .A1(men_men_n406_), .B0(men_men_n485_), .B1(men_men_n78_), .Y(men_men_n2068_));
  NA2        u2019(.A(men_men_n117_), .B(men_men_n519_), .Y(men_men_n2069_));
  OAI220     u2020(.A0(men_men_n2069_), .A1(men_men_n1853_), .B0(men_men_n2068_), .B1(x4), .Y(men_men_n2070_));
  INV        u2021(.A(men_men_n2070_), .Y(men_men_n2071_));
  AOI210     u2022(.A0(men_men_n2071_), .A1(men_men_n2067_), .B0(men_men_n188_), .Y(men_men_n2072_));
  NO4        u2023(.A(men_men_n598_), .B(men_men_n571_), .C(men_men_n686_), .D(men_men_n685_), .Y(men_men_n2073_));
  NA2        u2024(.A(men_men_n2073_), .B(x3), .Y(men_men_n2074_));
  NO4        u2025(.A(men_men_n791_), .B(men_men_n1182_), .C(men_men_n758_), .D(x5), .Y(men_men_n2075_));
  NO3        u2026(.A(x6), .B(men_men_n56_), .C(x1), .Y(men_men_n2076_));
  NA2        u2027(.A(men_men_n2076_), .B(men_men_n288_), .Y(men_men_n2077_));
  OAI210     u2028(.A0(men_men_n1827_), .A1(men_men_n377_), .B0(men_men_n2077_), .Y(men_men_n2078_));
  NA4        u2029(.A(men_men_n620_), .B(men_men_n181_), .C(x6), .D(men_men_n107_), .Y(men_men_n2079_));
  NO2        u2030(.A(men_men_n839_), .B(men_men_n253_), .Y(men_men_n2080_));
  NOi41      u2031(.An(men_men_n2079_), .B(men_men_n2080_), .C(men_men_n2078_), .D(men_men_n2075_), .Y(men_men_n2081_));
  AOI210     u2032(.A0(men_men_n2081_), .A1(men_men_n2074_), .B0(men_men_n523_), .Y(men_men_n2082_));
  OAI210     u2033(.A0(men_men_n597_), .A1(men_men_n464_), .B0(men_men_n920_), .Y(men_men_n2083_));
  NO3        u2034(.A(men_men_n372_), .B(men_men_n77_), .C(men_men_n53_), .Y(men_men_n2084_));
  NO3        u2035(.A(men_men_n457_), .B(men_men_n348_), .C(men_men_n50_), .Y(men_men_n2085_));
  OAI210     u2036(.A0(men_men_n2085_), .A1(men_men_n2084_), .B0(men_men_n1118_), .Y(men_men_n2086_));
  AOI210     u2037(.A0(men_men_n2086_), .A1(men_men_n2083_), .B0(men_men_n392_), .Y(men_men_n2087_));
  NO2        u2038(.A(men_men_n218_), .B(men_men_n528_), .Y(men_men_n2088_));
  OAI210     u2039(.A0(men_men_n139_), .A1(x2), .B0(men_men_n2088_), .Y(men_men_n2089_));
  NA3        u2040(.A(men_men_n406_), .B(men_men_n327_), .C(men_men_n77_), .Y(men_men_n2090_));
  OA210      u2041(.A0(men_men_n248_), .A1(men_men_n231_), .B0(men_men_n2090_), .Y(men_men_n2091_));
  AOI210     u2042(.A0(men_men_n2091_), .A1(men_men_n2089_), .B0(men_men_n64_), .Y(men_men_n2092_));
  NA2        u2043(.A(men_men_n122_), .B(men_men_n57_), .Y(men_men_n2093_));
  AOI220     u2044(.A0(men_men_n1522_), .A1(men_men_n889_), .B0(men_men_n277_), .B1(x4), .Y(men_men_n2094_));
  AOI220     u2045(.A0(men_men_n1570_), .A1(men_men_n599_), .B0(men_men_n707_), .B1(men_men_n758_), .Y(men_men_n2095_));
  OAI220     u2046(.A0(men_men_n2095_), .A1(men_men_n2093_), .B0(men_men_n2094_), .B1(men_men_n193_), .Y(men_men_n2096_));
  OR3        u2047(.A(men_men_n2096_), .B(men_men_n2092_), .C(men_men_n2087_), .Y(men_men_n2097_));
  NO4        u2048(.A(men_men_n2097_), .B(men_men_n2082_), .C(men_men_n2072_), .D(men_men_n2064_), .Y(men_men_n2098_));
  OAI210     u2049(.A0(men_men_n2051_), .A1(x3), .B0(men_men_n2098_), .Y(men32));
  OAI210     u2050(.A0(men_men_n548_), .A1(men_men_n53_), .B0(men_men_n411_), .Y(men_men_n2100_));
  NA2        u2051(.A(men_men_n503_), .B(x2), .Y(men_men_n2101_));
  AOI210     u2052(.A0(men_men_n2101_), .A1(men_men_n2100_), .B0(men_men_n57_), .Y(men_men_n2102_));
  OAI210     u2053(.A0(men_men_n2102_), .A1(men_men_n774_), .B0(men_men_n56_), .Y(men_men_n2103_));
  OAI210     u2054(.A0(men_men_n1639_), .A1(men_men_n1396_), .B0(men_men_n1424_), .Y(men_men_n2104_));
  AOI210     u2055(.A0(men_men_n2032_), .A1(men_men_n281_), .B0(men_men_n2104_), .Y(men_men_n2105_));
  AOI210     u2056(.A0(men_men_n2105_), .A1(men_men_n2103_), .B0(men_men_n50_), .Y(men_men_n2106_));
  NA3        u2057(.A(men_men_n1492_), .B(men_men_n789_), .C(men_men_n291_), .Y(men_men_n2107_));
  INV        u2058(.A(men_men_n731_), .Y(men_men_n2108_));
  OAI220     u2059(.A0(men_men_n1021_), .A1(men_men_n233_), .B0(men_men_n667_), .B1(men_men_n210_), .Y(men_men_n2109_));
  NO3        u2060(.A(men_men_n373_), .B(men_men_n556_), .C(men_men_n795_), .Y(men_men_n2110_));
  NO3        u2061(.A(men_men_n1318_), .B(men_men_n567_), .C(men_men_n275_), .Y(men_men_n2111_));
  NO4        u2062(.A(men_men_n2111_), .B(men_men_n2110_), .C(men_men_n2109_), .D(men_men_n2108_), .Y(men_men_n2112_));
  AOI210     u2063(.A0(men_men_n2112_), .A1(men_men_n2107_), .B0(men_men_n143_), .Y(men_men_n2113_));
  OAI220     u2064(.A0(men_men_n399_), .A1(x7), .B0(men_men_n300_), .B1(men_men_n296_), .Y(men_men_n2114_));
  NA2        u2065(.A(men_men_n2114_), .B(men_men_n936_), .Y(men_men_n2115_));
  NO2        u2066(.A(men_men_n539_), .B(men_men_n845_), .Y(men_men_n2116_));
  AOI220     u2067(.A0(men_men_n2116_), .A1(men_men_n1809_), .B0(men_men_n520_), .B1(men_men_n132_), .Y(men_men_n2117_));
  AOI210     u2068(.A0(men_men_n2117_), .A1(men_men_n2115_), .B0(men_men_n109_), .Y(men_men_n2118_));
  NA3        u2069(.A(men_men_n1272_), .B(men_men_n1103_), .C(men_men_n116_), .Y(men_men_n2119_));
  AOI220     u2070(.A0(men_men_n1308_), .A1(men_men_n686_), .B0(men_men_n1194_), .B1(men_men_n1011_), .Y(men_men_n2120_));
  AOI210     u2071(.A0(men_men_n2120_), .A1(men_men_n2119_), .B0(men_men_n56_), .Y(men_men_n2121_));
  NA2        u2072(.A(men_men_n936_), .B(men_men_n57_), .Y(men_men_n2122_));
  NOi21      u2073(.An(men_men_n2122_), .B(men_men_n132_), .Y(men_men_n2123_));
  NA2        u2074(.A(men_men_n980_), .B(men_men_n253_), .Y(men_men_n2124_));
  NO3        u2075(.A(men_men_n2124_), .B(men_men_n2123_), .C(men_men_n59_), .Y(men_men_n2125_));
  OR4        u2076(.A(men_men_n2125_), .B(men_men_n2121_), .C(men_men_n2118_), .D(men_men_n2113_), .Y(men_men_n2126_));
  OAI210     u2077(.A0(men_men_n2126_), .A1(men_men_n2106_), .B0(men_men_n107_), .Y(men_men_n2127_));
  NO3        u2078(.A(men_men_n1182_), .B(men_men_n147_), .C(men_men_n125_), .Y(men_men_n2128_));
  NO2        u2079(.A(men_men_n380_), .B(men_men_n55_), .Y(men_men_n2129_));
  NA2        u2080(.A(men_men_n2129_), .B(men_men_n115_), .Y(men_men_n2130_));
  OAI210     u2081(.A0(men_men_n616_), .A1(men_men_n573_), .B0(men_men_n798_), .Y(men_men_n2131_));
  NA2        u2082(.A(men_men_n2131_), .B(men_men_n2130_), .Y(men_men_n2132_));
  OAI210     u2083(.A0(men_men_n2132_), .A1(men_men_n2128_), .B0(x3), .Y(men_men_n2133_));
  NA2        u2084(.A(men_men_n275_), .B(men_men_n50_), .Y(men_men_n2134_));
  AOI210     u2085(.A0(men_men_n62_), .A1(men_men_n109_), .B0(men_men_n2134_), .Y(men_men_n2135_));
  OAI210     u2086(.A0(men_men_n2135_), .A1(men_men_n1791_), .B0(men_men_n685_), .Y(men_men_n2136_));
  NO3        u2087(.A(men_men_n302_), .B(men_men_n175_), .C(men_men_n123_), .Y(men_men_n2137_));
  NO3        u2088(.A(men_men_n789_), .B(men_men_n360_), .C(men_men_n143_), .Y(men_men_n2138_));
  OAI210     u2089(.A0(men_men_n2138_), .A1(men_men_n2137_), .B0(men_men_n59_), .Y(men_men_n2139_));
  NA2        u2090(.A(men_men_n1107_), .B(men_men_n71_), .Y(men_men_n2140_));
  NO2        u2091(.A(men_men_n1857_), .B(men_men_n573_), .Y(men_men_n2141_));
  NO2        u2092(.A(men_men_n2141_), .B(men_men_n2140_), .Y(men_men_n2142_));
  NO2        u2093(.A(men_men_n278_), .B(men_men_n57_), .Y(men_men_n2143_));
  NO3        u2094(.A(men_men_n1264_), .B(men_men_n218_), .C(men_men_n260_), .Y(men_men_n2144_));
  NO3        u2095(.A(men_men_n2144_), .B(men_men_n2142_), .C(x1), .Y(men_men_n2145_));
  NA4        u2096(.A(men_men_n2145_), .B(men_men_n2139_), .C(men_men_n2136_), .D(men_men_n2133_), .Y(men_men_n2146_));
  NA3        u2097(.A(men_men_n1832_), .B(men_men_n541_), .C(men_men_n278_), .Y(men_men_n2147_));
  NO2        u2098(.A(men_men_n2147_), .B(men_men_n302_), .Y(men_men_n2148_));
  NA4        u2099(.A(men_men_n1217_), .B(men_men_n517_), .C(men_men_n385_), .D(men_men_n233_), .Y(men_men_n2149_));
  NO2        u2100(.A(men_men_n1203_), .B(men_men_n383_), .Y(men_men_n2150_));
  NO2        u2101(.A(men_men_n1764_), .B(men_men_n64_), .Y(men_men_n2151_));
  NO3        u2102(.A(men_men_n2151_), .B(men_men_n2150_), .C(men_men_n53_), .Y(men_men_n2152_));
  NO3        u2103(.A(men_men_n461_), .B(men_men_n1051_), .C(men_men_n122_), .Y(men_men_n2153_));
  OAI220     u2104(.A0(men_men_n670_), .A1(men_men_n175_), .B0(men_men_n353_), .B1(men_men_n143_), .Y(men_men_n2154_));
  OAI210     u2105(.A0(men_men_n2154_), .A1(men_men_n2153_), .B0(men_men_n68_), .Y(men_men_n2155_));
  NO2        u2106(.A(men_men_n1903_), .B(men_men_n364_), .Y(men_men_n2156_));
  OAI210     u2107(.A0(men_men_n1797_), .A1(men_men_n591_), .B0(men_men_n2156_), .Y(men_men_n2157_));
  NA4        u2108(.A(men_men_n2157_), .B(men_men_n2155_), .C(men_men_n2152_), .D(men_men_n2149_), .Y(men_men_n2158_));
  OAI210     u2109(.A0(men_men_n2158_), .A1(men_men_n2148_), .B0(men_men_n2146_), .Y(men_men_n2159_));
  NO3        u2110(.A(x8), .B(men_men_n71_), .C(x2), .Y(men_men_n2160_));
  AOI220     u2111(.A0(men_men_n542_), .A1(men_men_n798_), .B0(men_men_n660_), .B1(men_men_n258_), .Y(men_men_n2161_));
  NO2        u2112(.A(men_men_n2161_), .B(men_men_n268_), .Y(men_men_n2162_));
  NA2        u2113(.A(men_men_n980_), .B(men_men_n1101_), .Y(men_men_n2163_));
  NO2        u2114(.A(men_men_n670_), .B(men_men_n2163_), .Y(men_men_n2164_));
  AOI210     u2115(.A0(men_men_n571_), .A1(men_men_n607_), .B0(men_men_n676_), .Y(men_men_n2165_));
  NO2        u2116(.A(men_men_n2165_), .B(men_men_n1746_), .Y(men_men_n2166_));
  NO2        u2117(.A(men_men_n446_), .B(men_men_n428_), .Y(men_men_n2167_));
  NOi31      u2118(.An(men_men_n1444_), .B(men_men_n2167_), .C(men_men_n571_), .Y(men_men_n2168_));
  NO4        u2119(.A(men_men_n2168_), .B(men_men_n2166_), .C(men_men_n2164_), .D(men_men_n2162_), .Y(men_men_n2169_));
  NA3        u2120(.A(men_men_n2169_), .B(men_men_n2159_), .C(men_men_n2127_), .Y(men33));
  OAI210     u2121(.A0(men_men_n2553_), .A1(x1), .B0(men_men_n204_), .Y(men_men_n2171_));
  OAI210     u2122(.A0(men_men_n2002_), .A1(men_men_n180_), .B0(men_men_n327_), .Y(men_men_n2172_));
  OAI220     u2123(.A0(men_men_n1039_), .A1(men_men_n795_), .B0(men_men_n1604_), .B1(men_men_n352_), .Y(men_men_n2173_));
  NA3        u2124(.A(men_men_n2173_), .B(men_men_n2172_), .C(men_men_n619_), .Y(men_men_n2174_));
  AOI210     u2125(.A0(men_men_n2171_), .A1(x5), .B0(men_men_n2174_), .Y(men_men_n2175_));
  NA2        u2126(.A(men_men_n232_), .B(men_men_n76_), .Y(men_men_n2176_));
  NA4        u2127(.A(men_men_n1676_), .B(men_men_n549_), .C(men_men_n249_), .D(x4), .Y(men_men_n2177_));
  AOI210     u2128(.A0(men_men_n2177_), .A1(men_men_n2176_), .B0(men_men_n352_), .Y(men_men_n2178_));
  OAI210     u2129(.A0(men_men_n431_), .A1(men_men_n272_), .B0(men_men_n53_), .Y(men_men_n2179_));
  AOI210     u2130(.A0(men_men_n2179_), .A1(men_men_n433_), .B0(men_men_n64_), .Y(men_men_n2180_));
  NA2        u2131(.A(men_men_n1592_), .B(men_men_n71_), .Y(men_men_n2181_));
  NO3        u2132(.A(men_men_n2181_), .B(men_men_n2180_), .C(men_men_n2178_), .Y(men_men_n2182_));
  OAI210     u2133(.A0(men_men_n2175_), .A1(x4), .B0(men_men_n2182_), .Y(men_men_n2183_));
  OAI210     u2134(.A0(men_men_n145_), .A1(x5), .B0(men_men_n242_), .Y(men_men_n2184_));
  NA2        u2135(.A(men_men_n188_), .B(x4), .Y(men_men_n2185_));
  NA2        u2136(.A(men_men_n307_), .B(men_men_n288_), .Y(men_men_n2186_));
  NO2        u2137(.A(men_men_n936_), .B(men_men_n230_), .Y(men_men_n2187_));
  NA2        u2138(.A(men_men_n622_), .B(x7), .Y(men_men_n2188_));
  OAI220     u2139(.A0(men_men_n2188_), .A1(men_men_n2187_), .B0(men_men_n2186_), .B1(men_men_n2185_), .Y(men_men_n2189_));
  AOI210     u2140(.A0(men_men_n2184_), .A1(men_men_n988_), .B0(men_men_n2189_), .Y(men_men_n2190_));
  NA2        u2141(.A(men_men_n215_), .B(men_men_n929_), .Y(men_men_n2191_));
  AOI210     u2142(.A0(men_men_n2191_), .A1(men_men_n2122_), .B0(men_men_n216_), .Y(men_men_n2192_));
  NO2        u2143(.A(men_men_n1578_), .B(men_men_n930_), .Y(men_men_n2193_));
  OAI210     u2144(.A0(men_men_n845_), .A1(men_men_n51_), .B0(x6), .Y(men_men_n2194_));
  NA3        u2145(.A(men_men_n899_), .B(men_men_n715_), .C(men_men_n55_), .Y(men_men_n2195_));
  OAI210     u2146(.A0(men_men_n601_), .A1(men_men_n494_), .B0(men_men_n2195_), .Y(men_men_n2196_));
  NO4        u2147(.A(men_men_n2196_), .B(men_men_n2194_), .C(men_men_n2193_), .D(men_men_n2192_), .Y(men_men_n2197_));
  OAI210     u2148(.A0(men_men_n2190_), .A1(men_men_n50_), .B0(men_men_n2197_), .Y(men_men_n2198_));
  NA3        u2149(.A(men_men_n2198_), .B(men_men_n2183_), .C(men_men_n59_), .Y(men_men_n2199_));
  NA2        u2150(.A(men_men_n524_), .B(men_men_n108_), .Y(men_men_n2200_));
  NO3        u2151(.A(men_men_n1504_), .B(men_men_n372_), .C(x4), .Y(men_men_n2201_));
  AOI210     u2152(.A0(men_men_n2201_), .A1(men_men_n2200_), .B0(men_men_n434_), .Y(men_men_n2202_));
  NA2        u2153(.A(men_men_n796_), .B(men_men_n107_), .Y(men_men_n2203_));
  NA2        u2154(.A(men_men_n2203_), .B(men_men_n456_), .Y(men_men_n2204_));
  NO2        u2155(.A(men_men_n691_), .B(men_men_n373_), .Y(men_men_n2205_));
  AOI210     u2156(.A0(men_men_n2205_), .A1(men_men_n2204_), .B0(x1), .Y(men_men_n2206_));
  OAI210     u2157(.A0(men_men_n2202_), .A1(men_men_n59_), .B0(men_men_n2206_), .Y(men_men_n2207_));
  AOI220     u2158(.A0(men_men_n670_), .A1(men_men_n239_), .B0(men_men_n385_), .B1(men_men_n233_), .Y(men_men_n2208_));
  NA2        u2159(.A(men_men_n716_), .B(men_men_n945_), .Y(men_men_n2209_));
  OAI210     u2160(.A0(men_men_n2209_), .A1(men_men_n2208_), .B0(men_men_n301_), .Y(men_men_n2210_));
  AOI210     u2161(.A0(men_men_n2032_), .A1(men_men_n217_), .B0(men_men_n53_), .Y(men_men_n2211_));
  NO2        u2162(.A(men_men_n143_), .B(men_men_n337_), .Y(men_men_n2212_));
  AOI220     u2163(.A0(men_men_n2212_), .A1(men_men_n962_), .B0(men_men_n655_), .B1(men_men_n352_), .Y(men_men_n2213_));
  NA2        u2164(.A(men_men_n441_), .B(men_men_n491_), .Y(men_men_n2214_));
  NO3        u2165(.A(men_men_n2214_), .B(men_men_n993_), .C(men_men_n185_), .Y(men_men_n2215_));
  AOI210     u2166(.A0(men_men_n1723_), .A1(men_men_n1143_), .B0(men_men_n2215_), .Y(men_men_n2216_));
  NA4        u2167(.A(men_men_n2216_), .B(men_men_n2213_), .C(men_men_n2211_), .D(men_men_n2210_), .Y(men_men_n2217_));
  NA3        u2168(.A(men_men_n2217_), .B(men_men_n2207_), .C(men_men_n57_), .Y(men_men_n2218_));
  INV        u2169(.A(men_men_n481_), .Y(men_men_n2219_));
  OAI210     u2170(.A0(men_men_n2212_), .A1(men_men_n1977_), .B0(x2), .Y(men_men_n2220_));
  INV        u2171(.A(men_men_n2220_), .Y(men_men_n2221_));
  AO220      u2172(.A0(men_men_n2221_), .A1(x0), .B0(men_men_n2219_), .B1(men_men_n140_), .Y(men_men_n2222_));
  NA3        u2173(.A(men_men_n758_), .B(men_men_n352_), .C(men_men_n60_), .Y(men_men_n2223_));
  NO2        u2174(.A(men_men_n2160_), .B(men_men_n410_), .Y(men_men_n2224_));
  NA2        u2175(.A(men_men_n620_), .B(men_men_n506_), .Y(men_men_n2225_));
  OAI220     u2176(.A0(men_men_n2225_), .A1(men_men_n2224_), .B0(men_men_n2223_), .B1(men_men_n71_), .Y(men_men_n2226_));
  OAI210     u2177(.A0(men_men_n1471_), .A1(men_men_n348_), .B0(men_men_n110_), .Y(men_men_n2227_));
  AOI210     u2178(.A0(men_men_n571_), .A1(men_men_n461_), .B0(men_men_n140_), .Y(men_men_n2228_));
  OAI210     u2179(.A0(men_men_n2228_), .A1(men_men_n385_), .B0(men_men_n2227_), .Y(men_men_n2229_));
  OAI210     u2180(.A0(men_men_n2229_), .A1(men_men_n2226_), .B0(men_men_n101_), .Y(men_men_n2230_));
  NA3        u2181(.A(men_men_n1163_), .B(men_men_n133_), .C(men_men_n380_), .Y(men_men_n2231_));
  NA2        u2182(.A(men_men_n2231_), .B(men_men_n1750_), .Y(men_men_n2232_));
  AOI220     u2183(.A0(men_men_n2129_), .A1(men_men_n295_), .B0(men_men_n1308_), .B1(men_men_n1124_), .Y(men_men_n2233_));
  NA3        u2184(.A(men_men_n2233_), .B(men_men_n2232_), .C(men_men_n2230_), .Y(men_men_n2234_));
  AOI210     u2185(.A0(men_men_n2222_), .A1(x7), .B0(men_men_n2234_), .Y(men_men_n2235_));
  NA3        u2186(.A(men_men_n2235_), .B(men_men_n2218_), .C(men_men_n2199_), .Y(men34));
  NO2        u2187(.A(men_men_n1882_), .B(men_men_n838_), .Y(men_men_n2237_));
  NO2        u2188(.A(men_men_n2237_), .B(men_men_n318_), .Y(men_men_n2238_));
  AOI210     u2189(.A0(men_men_n1957_), .A1(men_men_n531_), .B0(men_men_n142_), .Y(men_men_n2239_));
  NA2        u2190(.A(men_men_n1882_), .B(x0), .Y(men_men_n2240_));
  INV        u2191(.A(men_men_n2240_), .Y(men_men_n2241_));
  NO3        u2192(.A(men_men_n2241_), .B(men_men_n2239_), .C(men_men_n2238_), .Y(men_men_n2242_));
  NO2        u2193(.A(men_men_n2242_), .B(men_men_n469_), .Y(men_men_n2243_));
  NA2        u2194(.A(men_men_n718_), .B(x8), .Y(men_men_n2244_));
  AO210      u2195(.A0(men_men_n2244_), .A1(men_men_n479_), .B0(men_men_n645_), .Y(men_men_n2245_));
  NO2        u2196(.A(men_men_n2245_), .B(men_men_n268_), .Y(men_men_n2246_));
  NO2        u2197(.A(men_men_n1540_), .B(men_men_n58_), .Y(men_men_n2247_));
  NA3        u2198(.A(men_men_n2247_), .B(men_men_n338_), .C(x8), .Y(men_men_n2248_));
  NO3        u2199(.A(men_men_n961_), .B(men_men_n691_), .C(men_men_n450_), .Y(men_men_n2249_));
  AOI210     u2200(.A0(men_men_n1525_), .A1(men_men_n326_), .B0(men_men_n2249_), .Y(men_men_n2250_));
  NA2        u2201(.A(men_men_n649_), .B(men_men_n318_), .Y(men_men_n2251_));
  NA2        u2202(.A(men_men_n136_), .B(x0), .Y(men_men_n2252_));
  NAi31      u2203(.An(men_men_n2252_), .B(men_men_n2251_), .C(men_men_n783_), .Y(men_men_n2253_));
  NA3        u2204(.A(men_men_n1536_), .B(men_men_n1347_), .C(men_men_n50_), .Y(men_men_n2254_));
  NA4        u2205(.A(men_men_n2254_), .B(men_men_n2253_), .C(men_men_n2250_), .D(men_men_n2248_), .Y(men_men_n2255_));
  NA3        u2206(.A(men_men_n1066_), .B(men_men_n364_), .C(men_men_n734_), .Y(men_men_n2256_));
  NA3        u2207(.A(men_men_n1103_), .B(men_men_n169_), .C(men_men_n1052_), .Y(men_men_n2257_));
  AOI210     u2208(.A0(men_men_n2257_), .A1(men_men_n2256_), .B0(men_men_n744_), .Y(men_men_n2258_));
  AOI210     u2209(.A0(men_men_n1707_), .A1(men_men_n132_), .B0(men_men_n2258_), .Y(men_men_n2259_));
  AOI210     u2210(.A0(men_men_n542_), .A1(men_men_n798_), .B0(men_men_n257_), .Y(men_men_n2260_));
  OAI220     u2211(.A0(men_men_n2260_), .A1(men_men_n59_), .B0(men_men_n1076_), .B1(men_men_n55_), .Y(men_men_n2261_));
  NA3        u2212(.A(men_men_n2261_), .B(men_men_n718_), .C(men_men_n56_), .Y(men_men_n2262_));
  OAI210     u2213(.A0(men_men_n2259_), .A1(men_men_n143_), .B0(men_men_n2262_), .Y(men_men_n2263_));
  NO4        u2214(.A(men_men_n2263_), .B(men_men_n2255_), .C(men_men_n2246_), .D(men_men_n2243_), .Y(men_men_n2264_));
  NO2        u2215(.A(men_men_n308_), .B(men_men_n929_), .Y(men_men_n2265_));
  NO3        u2216(.A(men_men_n2265_), .B(men_men_n439_), .C(men_men_n326_), .Y(men_men_n2266_));
  NO3        u2217(.A(men_men_n2143_), .B(men_men_n301_), .C(men_men_n1052_), .Y(men_men_n2267_));
  NO2        u2218(.A(men_men_n2267_), .B(men_men_n1496_), .Y(men_men_n2268_));
  OAI210     u2219(.A0(men_men_n2268_), .A1(men_men_n2266_), .B0(x2), .Y(men_men_n2269_));
  OAI210     u2220(.A0(men_men_n848_), .A1(men_men_n368_), .B0(men_men_n2269_), .Y(men_men_n2270_));
  NA2        u2221(.A(men_men_n311_), .B(x4), .Y(men_men_n2271_));
  OAI220     u2222(.A0(men_men_n730_), .A1(men_men_n55_), .B0(men_men_n282_), .B1(men_men_n106_), .Y(men_men_n2272_));
  NO4        u2223(.A(men_men_n443_), .B(men_men_n77_), .C(x7), .D(x3), .Y(men_men_n2273_));
  NO2        u2224(.A(men_men_n1066_), .B(men_men_n289_), .Y(men_men_n2274_));
  NO4        u2225(.A(men_men_n2274_), .B(men_men_n2273_), .C(men_men_n2272_), .D(men_men_n2271_), .Y(men_men_n2275_));
  NA4        u2226(.A(men_men_n718_), .B(men_men_n181_), .C(men_men_n57_), .D(men_men_n107_), .Y(men_men_n2276_));
  NA3        u2227(.A(men_men_n1344_), .B(men_men_n260_), .C(x7), .Y(men_men_n2277_));
  NA2        u2228(.A(men_men_n2277_), .B(men_men_n2276_), .Y(men_men_n2278_));
  OAI210     u2229(.A0(men_men_n2278_), .A1(men_men_n2275_), .B0(men_men_n166_), .Y(men_men_n2279_));
  NA3        u2230(.A(men_men_n1107_), .B(men_men_n297_), .C(men_men_n569_), .Y(men_men_n2280_));
  NA2        u2231(.A(men_men_n1111_), .B(men_men_n660_), .Y(men_men_n2281_));
  OAI210     u2232(.A0(men_men_n2281_), .A1(men_men_n269_), .B0(men_men_n2079_), .Y(men_men_n2282_));
  AOI220     u2233(.A0(men_men_n2282_), .A1(x7), .B0(men_men_n979_), .B1(men_men_n646_), .Y(men_men_n2283_));
  OAI210     u2234(.A0(men_men_n1970_), .A1(men_men_n265_), .B0(men_men_n722_), .Y(men_men_n2284_));
  AOI220     u2235(.A0(men_men_n406_), .A1(x8), .B0(men_men_n91_), .B1(x2), .Y(men_men_n2285_));
  AOI210     u2236(.A0(men_men_n273_), .A1(men_men_n53_), .B0(men_men_n637_), .Y(men_men_n2286_));
  OAI220     u2237(.A0(men_men_n2286_), .A1(men_men_n96_), .B0(men_men_n2285_), .B1(men_men_n1294_), .Y(men_men_n2287_));
  AOI220     u2238(.A0(men_men_n2287_), .A1(men_men_n1273_), .B0(men_men_n2284_), .B1(men_men_n1457_), .Y(men_men_n2288_));
  NA4        u2239(.A(men_men_n2288_), .B(men_men_n2283_), .C(men_men_n2280_), .D(men_men_n2279_), .Y(men_men_n2289_));
  AOI210     u2240(.A0(men_men_n2270_), .A1(men_men_n798_), .B0(men_men_n2289_), .Y(men_men_n2290_));
  OAI210     u2241(.A0(men_men_n2264_), .A1(x2), .B0(men_men_n2290_), .Y(men35));
  NA2        u2242(.A(men_men_n494_), .B(men_men_n181_), .Y(men_men_n2292_));
  AOI220     u2243(.A0(men_men_n620_), .A1(men_men_n55_), .B0(men_men_n758_), .B1(men_men_n1176_), .Y(men_men_n2293_));
  AOI210     u2244(.A0(men_men_n2293_), .A1(men_men_n2292_), .B0(men_men_n71_), .Y(men_men_n2294_));
  NO3        u2245(.A(men_men_n502_), .B(men_men_n461_), .C(men_men_n337_), .Y(men_men_n2295_));
  OAI210     u2246(.A0(men_men_n2295_), .A1(men_men_n2294_), .B0(x2), .Y(men_men_n2296_));
  AOI210     u2247(.A0(men_men_n218_), .A1(x0), .B0(men_men_n277_), .Y(men_men_n2297_));
  OAI220     u2248(.A0(men_men_n2297_), .A1(men_men_n651_), .B0(men_men_n201_), .B1(x4), .Y(men_men_n2298_));
  NA2        u2249(.A(men_men_n2298_), .B(men_men_n140_), .Y(men_men_n2299_));
  NA3        u2250(.A(men_men_n406_), .B(x8), .C(men_men_n71_), .Y(men_men_n2300_));
  AOI210     u2251(.A0(men_men_n2300_), .A1(men_men_n1652_), .B0(men_men_n670_), .Y(men_men_n2301_));
  OAI210     u2252(.A0(men_men_n2223_), .A1(x6), .B0(men_men_n733_), .Y(men_men_n2302_));
  NO2        u2253(.A(men_men_n2302_), .B(men_men_n2301_), .Y(men_men_n2303_));
  NA3        u2254(.A(men_men_n2303_), .B(men_men_n2299_), .C(men_men_n2296_), .Y(men_men_n2304_));
  NAi21      u2255(.An(men_men_n1617_), .B(men_men_n1250_), .Y(men_men_n2305_));
  NA2        u2256(.A(men_men_n216_), .B(men_men_n556_), .Y(men_men_n2306_));
  NO2        u2257(.A(men_men_n428_), .B(men_men_n422_), .Y(men_men_n2307_));
  AOI220     u2258(.A0(men_men_n2307_), .A1(men_men_n2306_), .B0(men_men_n2305_), .B1(men_men_n56_), .Y(men_men_n2308_));
  NA2        u2259(.A(men_men_n748_), .B(men_men_n683_), .Y(men_men_n2309_));
  NO3        u2260(.A(men_men_n665_), .B(men_men_n55_), .C(x6), .Y(men_men_n2310_));
  OAI210     u2261(.A0(men_men_n2310_), .A1(men_men_n693_), .B0(men_men_n221_), .Y(men_men_n2311_));
  NA2        u2262(.A(men_men_n1280_), .B(men_men_n63_), .Y(men_men_n2312_));
  OAI210     u2263(.A0(men_men_n1035_), .A1(x6), .B0(men_men_n465_), .Y(men_men_n2313_));
  NA3        u2264(.A(men_men_n2313_), .B(men_men_n2312_), .C(men_men_n2311_), .Y(men_men_n2314_));
  NA3        u2265(.A(men_men_n1225_), .B(men_men_n736_), .C(x3), .Y(men_men_n2315_));
  NO3        u2266(.A(men_men_n2315_), .B(men_men_n667_), .C(men_men_n210_), .Y(men_men_n2316_));
  AOI210     u2267(.A0(men_men_n2314_), .A1(men_men_n50_), .B0(men_men_n2316_), .Y(men_men_n2317_));
  OAI210     u2268(.A0(men_men_n2309_), .A1(men_men_n2308_), .B0(men_men_n2317_), .Y(men_men_n2318_));
  AOI210     u2269(.A0(men_men_n2304_), .A1(men_men_n57_), .B0(men_men_n2318_), .Y(men_men_n2319_));
  NA2        u2270(.A(men_men_n936_), .B(men_men_n63_), .Y(men_men_n2320_));
  NO3        u2271(.A(men_men_n1035_), .B(men_men_n548_), .C(men_men_n123_), .Y(men_men_n2321_));
  OAI210     u2272(.A0(men_men_n159_), .A1(men_men_n67_), .B0(men_men_n2321_), .Y(men_men_n2322_));
  AOI210     u2273(.A0(men_men_n2322_), .A1(men_men_n2320_), .B0(men_men_n50_), .Y(men_men_n2323_));
  NA2        u2274(.A(men_men_n258_), .B(men_men_n737_), .Y(men_men_n2324_));
  OAI210     u2275(.A0(men_men_n258_), .A1(men_men_n568_), .B0(men_men_n2076_), .Y(men_men_n2325_));
  NA2        u2276(.A(men_men_n2325_), .B(men_men_n2324_), .Y(men_men_n2326_));
  OAI210     u2277(.A0(men_men_n2326_), .A1(men_men_n2323_), .B0(men_men_n59_), .Y(men_men_n2327_));
  NO4        u2278(.A(men_men_n930_), .B(men_men_n548_), .C(men_men_n360_), .D(men_men_n404_), .Y(men_men_n2328_));
  XN2        u2279(.A(x4), .B(x3), .Y(men_men_n2329_));
  NO3        u2280(.A(men_men_n2329_), .B(men_men_n650_), .C(men_men_n307_), .Y(men_men_n2330_));
  NO3        u2281(.A(men_men_n2330_), .B(men_men_n2328_), .C(men_men_n1405_), .Y(men_men_n2331_));
  OAI210     u2282(.A0(men_men_n523_), .A1(x3), .B0(men_men_n2331_), .Y(men_men_n2332_));
  NO3        u2283(.A(men_men_n730_), .B(men_men_n845_), .C(men_men_n278_), .Y(men_men_n2333_));
  OAI210     u2284(.A0(men_men_n2333_), .A1(men_men_n1405_), .B0(men_men_n50_), .Y(men_men_n2334_));
  NA3        u2285(.A(men_men_n1043_), .B(men_men_n796_), .C(men_men_n257_), .Y(men_men_n2335_));
  NA2        u2286(.A(men_men_n2335_), .B(men_men_n2334_), .Y(men_men_n2336_));
  AOI210     u2287(.A0(men_men_n2332_), .A1(men_men_n571_), .B0(men_men_n2336_), .Y(men_men_n2337_));
  OAI210     u2288(.A0(men_men_n1885_), .A1(men_men_n590_), .B0(men_men_n2160_), .Y(men_men_n2338_));
  OAI210     u2289(.A0(men_men_n2244_), .A1(x4), .B0(men_men_n2338_), .Y(men_men_n2339_));
  NA2        u2290(.A(men_men_n2339_), .B(men_men_n91_), .Y(men_men_n2340_));
  NO2        u2291(.A(x2), .B(men_men_n647_), .Y(men_men_n2341_));
  NO2        u2292(.A(men_men_n289_), .B(x6), .Y(men_men_n2342_));
  OAI210     u2293(.A0(men_men_n2341_), .A1(men_men_n1714_), .B0(men_men_n2342_), .Y(men_men_n2343_));
  NA4        u2294(.A(men_men_n2343_), .B(men_men_n2340_), .C(men_men_n2337_), .D(men_men_n2327_), .Y(men_men_n2344_));
  NA4        u2295(.A(men_men_n598_), .B(men_men_n670_), .C(men_men_n427_), .D(x6), .Y(men_men_n2345_));
  AOI210     u2296(.A0(men_men_n2345_), .A1(men_men_n423_), .B0(x1), .Y(men_men_n2346_));
  NO2        u2297(.A(men_men_n716_), .B(men_men_n667_), .Y(men_men_n2347_));
  OAI210     u2298(.A0(men_men_n461_), .A1(men_men_n170_), .B0(men_men_n780_), .Y(men_men_n2348_));
  AOI210     u2299(.A0(men_men_n2348_), .A1(men_men_n984_), .B0(men_men_n53_), .Y(men_men_n2349_));
  NO3        u2300(.A(men_men_n2349_), .B(men_men_n2347_), .C(men_men_n2346_), .Y(men_men_n2350_));
  NA3        u2301(.A(men_men_n1384_), .B(men_men_n1226_), .C(men_men_n802_), .Y(men_men_n2351_));
  AOI220     u2302(.A0(men_men_n1872_), .A1(men_men_n140_), .B0(men_men_n415_), .B1(men_men_n127_), .Y(men_men_n2352_));
  AOI210     u2303(.A0(men_men_n2352_), .A1(men_men_n2351_), .B0(men_men_n1452_), .Y(men_men_n2353_));
  NO2        u2304(.A(men_men_n620_), .B(x3), .Y(men_men_n2354_));
  NO3        u2305(.A(men_men_n678_), .B(men_men_n1540_), .C(x2), .Y(men_men_n2355_));
  AOI220     u2306(.A0(men_men_n2355_), .A1(men_men_n2354_), .B0(men_men_n1847_), .B1(men_men_n754_), .Y(men_men_n2356_));
  NA3        u2307(.A(x6), .B(x4), .C(x0), .Y(men_men_n2357_));
  OAI220     u2308(.A0(men_men_n2357_), .A1(men_men_n200_), .B0(men_men_n665_), .B1(men_men_n519_), .Y(men_men_n2358_));
  NO2        u2309(.A(men_men_n372_), .B(men_men_n351_), .Y(men_men_n2359_));
  AOI220     u2310(.A0(men_men_n2359_), .A1(men_men_n415_), .B0(men_men_n2358_), .B1(men_men_n898_), .Y(men_men_n2360_));
  OAI210     u2311(.A0(men_men_n2356_), .A1(men_men_n1119_), .B0(men_men_n2360_), .Y(men_men_n2361_));
  NO2        u2312(.A(men_men_n2361_), .B(men_men_n2353_), .Y(men_men_n2362_));
  OAI210     u2313(.A0(men_men_n2350_), .A1(men_men_n311_), .B0(men_men_n2362_), .Y(men_men_n2363_));
  AOI210     u2314(.A0(men_men_n2344_), .A1(x5), .B0(men_men_n2363_), .Y(men_men_n2364_));
  OAI210     u2315(.A0(men_men_n2319_), .A1(x5), .B0(men_men_n2364_), .Y(men36));
  OR4        u2316(.A(men_men_n931_), .B(men_men_n791_), .C(men_men_n375_), .D(men_men_n485_), .Y(men_men_n2366_));
  NA2        u2317(.A(men_men_n2129_), .B(men_men_n282_), .Y(men_men_n2367_));
  NA2        u2318(.A(men_men_n230_), .B(men_men_n121_), .Y(men_men_n2368_));
  NA3        u2319(.A(men_men_n2368_), .B(men_men_n2367_), .C(men_men_n2366_), .Y(men_men_n2369_));
  NO2        u2320(.A(men_men_n958_), .B(men_men_n528_), .Y(men_men_n2370_));
  AOI210     u2321(.A0(men_men_n1052_), .A1(x6), .B0(men_men_n419_), .Y(men_men_n2371_));
  NO2        u2322(.A(men_men_n2371_), .B(men_men_n359_), .Y(men_men_n2372_));
  OAI210     u2323(.A0(men_men_n2372_), .A1(men_men_n2370_), .B0(men_men_n461_), .Y(men_men_n2373_));
  NO2        u2324(.A(men_men_n634_), .B(men_men_n269_), .Y(men_men_n2374_));
  NO3        u2325(.A(men_men_n1806_), .B(men_men_n1539_), .C(men_men_n279_), .Y(men_men_n2375_));
  NO2        u2326(.A(men_men_n2320_), .B(men_men_n232_), .Y(men_men_n2376_));
  NO4        u2327(.A(men_men_n2376_), .B(men_men_n2375_), .C(men_men_n2374_), .D(men_men_n417_), .Y(men_men_n2377_));
  OAI210     u2328(.A0(men_men_n622_), .A1(men_men_n790_), .B0(men_men_n948_), .Y(men_men_n2378_));
  OAI220     u2329(.A0(men_men_n1583_), .A1(men_men_n1578_), .B0(men_men_n948_), .B1(men_men_n1052_), .Y(men_men_n2379_));
  AOI220     u2330(.A0(men_men_n2379_), .A1(men_men_n120_), .B0(men_men_n2378_), .B1(men_men_n612_), .Y(men_men_n2380_));
  NA3        u2331(.A(men_men_n2380_), .B(men_men_n2377_), .C(men_men_n2373_), .Y(men_men_n2381_));
  AOI210     u2332(.A0(men_men_n2369_), .A1(men_men_n338_), .B0(men_men_n2381_), .Y(men_men_n2382_));
  OAI210     u2333(.A0(men_men_n576_), .A1(men_men_n507_), .B0(men_men_n170_), .Y(men_men_n2383_));
  OAI210     u2334(.A0(men_men_n1917_), .A1(men_men_n70_), .B0(men_men_n2383_), .Y(men_men_n2384_));
  OAI210     u2335(.A0(men_men_n488_), .A1(men_men_n241_), .B0(men_men_n258_), .Y(men_men_n2385_));
  NO2        u2336(.A(men_men_n1926_), .B(men_men_n177_), .Y(men_men_n2386_));
  NA2        u2337(.A(men_men_n1165_), .B(men_men_n55_), .Y(men_men_n2387_));
  OAI210     u2338(.A0(men_men_n2387_), .A1(men_men_n2386_), .B0(men_men_n2385_), .Y(men_men_n2388_));
  OAI210     u2339(.A0(men_men_n2388_), .A1(men_men_n2384_), .B0(men_men_n876_), .Y(men_men_n2389_));
  AOI210     u2340(.A0(men_men_n106_), .A1(men_men_n109_), .B0(men_men_n340_), .Y(men_men_n2390_));
  NA2        u2341(.A(men_men_n655_), .B(men_men_n1540_), .Y(men_men_n2391_));
  OAI220     u2342(.A0(men_men_n2391_), .A1(men_men_n2390_), .B0(men_men_n733_), .B1(men_men_n1208_), .Y(men_men_n2392_));
  NO2        u2343(.A(men_men_n1347_), .B(men_men_n562_), .Y(men_men_n2393_));
  NO3        u2344(.A(men_men_n2393_), .B(men_men_n1722_), .C(men_men_n678_), .Y(men_men_n2394_));
  NOi31      u2345(.An(men_men_n1936_), .B(men_men_n2214_), .C(men_men_n743_), .Y(men_men_n2395_));
  NO3        u2346(.A(men_men_n2395_), .B(men_men_n2394_), .C(men_men_n2392_), .Y(men_men_n2396_));
  AOI210     u2347(.A0(men_men_n2396_), .A1(men_men_n2389_), .B0(x7), .Y(men_men_n2397_));
  NA2        u2348(.A(men_men_n139_), .B(men_men_n63_), .Y(men_men_n2398_));
  AOI210     u2349(.A0(men_men_n571_), .A1(men_men_n607_), .B0(men_men_n1143_), .Y(men_men_n2399_));
  NA4        u2350(.A(men_men_n2399_), .B(men_men_n2398_), .C(men_men_n961_), .D(men_men_n871_), .Y(men_men_n2400_));
  NA2        u2351(.A(men_men_n2400_), .B(men_men_n494_), .Y(men_men_n2401_));
  AOI220     u2352(.A0(men_men_n1676_), .A1(men_men_n261_), .B0(men_men_n1013_), .B1(men_men_n127_), .Y(men_men_n2402_));
  NO2        u2353(.A(men_men_n2402_), .B(men_men_n441_), .Y(men_men_n2403_));
  NO2        u2354(.A(men_men_n404_), .B(men_men_n230_), .Y(men_men_n2404_));
  NO3        u2355(.A(men_men_n2404_), .B(men_men_n1229_), .C(men_men_n59_), .Y(men_men_n2405_));
  AOI210     u2356(.A0(men_men_n1180_), .A1(men_men_n405_), .B0(x6), .Y(men_men_n2406_));
  NA3        u2357(.A(men_men_n1610_), .B(men_men_n282_), .C(men_men_n273_), .Y(men_men_n2407_));
  NA2        u2358(.A(men_men_n2407_), .B(men_men_n1564_), .Y(men_men_n2408_));
  NO4        u2359(.A(men_men_n2408_), .B(men_men_n2406_), .C(men_men_n2405_), .D(men_men_n2403_), .Y(men_men_n2409_));
  AOI210     u2360(.A0(men_men_n2409_), .A1(men_men_n2401_), .B0(men_men_n450_), .Y(men_men_n2410_));
  NO3        u2361(.A(men_men_n2329_), .B(men_men_n882_), .C(men_men_n493_), .Y(men_men_n2411_));
  AOI210     u2362(.A0(men_men_n1227_), .A1(men_men_n272_), .B0(men_men_n2411_), .Y(men_men_n2412_));
  NO2        u2363(.A(men_men_n852_), .B(men_men_n278_), .Y(men_men_n2413_));
  NA2        u2364(.A(men_men_n1165_), .B(men_men_n175_), .Y(men_men_n2414_));
  NO2        u2365(.A(men_men_n597_), .B(men_men_n109_), .Y(men_men_n2415_));
  AO210      u2366(.A0(men_men_n2415_), .A1(men_men_n2414_), .B0(men_men_n1693_), .Y(men_men_n2416_));
  NO2        u2367(.A(men_men_n457_), .B(men_men_n416_), .Y(men_men_n2417_));
  AOI220     u2368(.A0(men_men_n2417_), .A1(men_men_n2416_), .B0(men_men_n2413_), .B1(men_men_n295_), .Y(men_men_n2418_));
  OAI210     u2369(.A0(men_men_n2412_), .A1(x1), .B0(men_men_n2418_), .Y(men_men_n2419_));
  NO3        u2370(.A(men_men_n2419_), .B(men_men_n2410_), .C(men_men_n2397_), .Y(men_men_n2420_));
  OAI210     u2371(.A0(men_men_n2382_), .A1(men_men_n57_), .B0(men_men_n2420_), .Y(men37));
  NA3        u2372(.A(men_men_n1032_), .B(men_men_n142_), .C(x3), .Y(men_men_n2422_));
  NO2        u2373(.A(men_men_n2422_), .B(men_men_n671_), .Y(men_men_n2423_));
  NO3        u2374(.A(men_men_n1032_), .B(men_men_n375_), .C(men_men_n501_), .Y(men_men_n2424_));
  OAI210     u2375(.A0(men_men_n2424_), .A1(men_men_n2423_), .B0(men_men_n56_), .Y(men_men_n2425_));
  NA2        u2376(.A(men_men_n585_), .B(men_men_n734_), .Y(men_men_n2426_));
  AOI210     u2377(.A0(men_men_n2426_), .A1(men_men_n1014_), .B0(x3), .Y(men_men_n2427_));
  AOI220     u2378(.A0(men_men_n585_), .A1(men_men_n734_), .B0(men_men_n461_), .B1(men_men_n1013_), .Y(men_men_n2428_));
  NO2        u2379(.A(men_men_n650_), .B(men_men_n184_), .Y(men_men_n2429_));
  OAI220     u2380(.A0(men_men_n2429_), .A1(men_men_n823_), .B0(men_men_n2428_), .B1(men_men_n109_), .Y(men_men_n2430_));
  OAI210     u2381(.A0(men_men_n2430_), .A1(men_men_n2427_), .B0(men_men_n71_), .Y(men_men_n2431_));
  NA2        u2382(.A(men_men_n1145_), .B(men_men_n1035_), .Y(men_men_n2432_));
  OAI210     u2383(.A0(men_men_n1167_), .A1(men_men_n194_), .B0(men_men_n451_), .Y(men_men_n2433_));
  NA4        u2384(.A(men_men_n2433_), .B(men_men_n2432_), .C(men_men_n2431_), .D(men_men_n2425_), .Y(men_men_n2434_));
  NA2        u2385(.A(men_men_n422_), .B(men_men_n139_), .Y(men_men_n2435_));
  NO2        u2386(.A(men_men_n1639_), .B(men_men_n108_), .Y(men_men_n2436_));
  AOI210     u2387(.A0(men_men_n1905_), .A1(men_men_n846_), .B0(men_men_n2436_), .Y(men_men_n2437_));
  OAI220     u2388(.A0(men_men_n2437_), .A1(men_men_n51_), .B0(men_men_n1541_), .B1(men_men_n2435_), .Y(men_men_n2438_));
  AOI210     u2389(.A0(men_men_n2434_), .A1(men_men_n68_), .B0(men_men_n2438_), .Y(men_men_n2439_));
  OAI210     u2390(.A0(men_men_n273_), .A1(men_men_n1054_), .B0(men_men_n480_), .Y(men_men_n2440_));
  NA3        u2391(.A(men_men_n2440_), .B(men_men_n269_), .C(men_men_n1015_), .Y(men_men_n2441_));
  OAI210     u2392(.A0(men_men_n233_), .A1(men_men_n221_), .B0(men_men_n1652_), .Y(men_men_n2442_));
  NA2        u2393(.A(men_men_n346_), .B(men_men_n277_), .Y(men_men_n2443_));
  NA3        u2394(.A(men_men_n400_), .B(men_men_n802_), .C(men_men_n109_), .Y(men_men_n2444_));
  NO2        u2395(.A(men_men_n520_), .B(men_men_n56_), .Y(men_men_n2445_));
  NA3        u2396(.A(men_men_n2445_), .B(men_men_n2444_), .C(men_men_n2443_), .Y(men_men_n2446_));
  AOI210     u2397(.A0(men_men_n2442_), .A1(men_men_n501_), .B0(men_men_n2446_), .Y(men_men_n2447_));
  NO2        u2398(.A(men_men_n1136_), .B(men_men_n278_), .Y(men_men_n2448_));
  OAI210     u2399(.A0(men_men_n295_), .A1(men_men_n267_), .B0(men_men_n2448_), .Y(men_men_n2449_));
  OAI210     u2400(.A0(men_men_n652_), .A1(men_men_n140_), .B0(x3), .Y(men_men_n2450_));
  AOI210     u2401(.A0(men_men_n652_), .A1(men_men_n364_), .B0(men_men_n2450_), .Y(men_men_n2451_));
  AOI210     u2402(.A0(men_men_n1540_), .A1(men_men_n50_), .B0(men_men_n346_), .Y(men_men_n2452_));
  OAI210     u2403(.A0(men_men_n2452_), .A1(men_men_n399_), .B0(men_men_n56_), .Y(men_men_n2453_));
  NO2        u2404(.A(men_men_n2453_), .B(men_men_n2451_), .Y(men_men_n2454_));
  AOI220     u2405(.A0(men_men_n2454_), .A1(men_men_n2449_), .B0(men_men_n2447_), .B1(men_men_n2441_), .Y(men_men_n2455_));
  OAI210     u2406(.A0(men_men_n2455_), .A1(men_men_n1691_), .B0(men_men_n101_), .Y(men_men_n2456_));
  NA2        u2407(.A(men_men_n678_), .B(men_men_n1150_), .Y(men_men_n2457_));
  NOi21      u2408(.An(men_men_n1314_), .B(men_men_n110_), .Y(men_men_n2458_));
  AOI210     u2409(.A0(men_men_n2458_), .A1(men_men_n2457_), .B0(men_men_n431_), .Y(men_men_n2459_));
  NO2        u2410(.A(men_men_n2140_), .B(men_men_n55_), .Y(men_men_n2460_));
  OAI210     u2411(.A0(men_men_n2460_), .A1(men_men_n2459_), .B0(men_men_n1750_), .Y(men_men_n2461_));
  NA2        u2412(.A(men_men_n181_), .B(men_men_n107_), .Y(men_men_n2462_));
  NA2        u2413(.A(men_men_n670_), .B(x6), .Y(men_men_n2463_));
  AOI210     u2414(.A0(men_men_n2463_), .A1(men_men_n479_), .B0(men_men_n2462_), .Y(men_men_n2464_));
  AOI210     u2415(.A0(men_men_n353_), .A1(men_men_n142_), .B0(men_men_n143_), .Y(men_men_n2465_));
  OAI210     u2416(.A0(men_men_n2465_), .A1(men_men_n2464_), .B0(men_men_n346_), .Y(men_men_n2466_));
  AOI210     u2417(.A0(men_men_n598_), .A1(men_men_n431_), .B0(men_men_n1239_), .Y(men_men_n2467_));
  NO3        u2418(.A(men_men_n2467_), .B(men_men_n269_), .C(men_men_n63_), .Y(men_men_n2468_));
  OAI220     u2419(.A0(men_men_n2244_), .A1(men_men_n477_), .B0(men_men_n2015_), .B1(men_men_n385_), .Y(men_men_n2469_));
  OAI210     u2420(.A0(men_men_n2469_), .A1(men_men_n2468_), .B0(men_men_n53_), .Y(men_men_n2470_));
  NO3        u2421(.A(men_men_n2252_), .B(men_men_n916_), .C(men_men_n224_), .Y(men_men_n2471_));
  NO4        u2422(.A(men_men_n718_), .B(men_men_n586_), .C(men_men_n439_), .D(men_men_n1021_), .Y(men_men_n2472_));
  NO3        u2423(.A(men_men_n2472_), .B(men_men_n2471_), .C(men_men_n1027_), .Y(men_men_n2473_));
  NA4        u2424(.A(men_men_n2473_), .B(men_men_n2470_), .C(men_men_n2466_), .D(men_men_n2461_), .Y(men_men_n2474_));
  NO3        u2425(.A(men_men_n253_), .B(men_men_n352_), .C(men_men_n84_), .Y(men_men_n2475_));
  OAI210     u2426(.A0(men_men_n461_), .A1(men_men_n85_), .B0(men_men_n2475_), .Y(men_men_n2476_));
  NA2        u2427(.A(men_men_n1111_), .B(men_men_n177_), .Y(men_men_n2477_));
  OAI210     u2428(.A0(men_men_n2477_), .A1(x6), .B0(men_men_n2476_), .Y(men_men_n2478_));
  AOI220     u2429(.A0(men_men_n2478_), .A1(men_men_n1409_), .B0(men_men_n2474_), .B1(men_men_n57_), .Y(men_men_n2479_));
  NA3        u2430(.A(men_men_n2479_), .B(men_men_n2456_), .C(men_men_n2439_), .Y(men38));
  AOI210     u2431(.A0(men_men_n1595_), .A1(men_men_n190_), .B0(men_men_n945_), .Y(men_men_n2481_));
  AOI210     u2432(.A0(men_men_n1180_), .A1(men_men_n561_), .B0(men_men_n1051_), .Y(men_men_n2482_));
  NO3        u2433(.A(men_men_n1249_), .B(men_men_n318_), .C(x8), .Y(men_men_n2483_));
  NO3        u2434(.A(men_men_n2483_), .B(men_men_n2482_), .C(men_men_n2481_), .Y(men_men_n2484_));
  NO2        u2435(.A(men_men_n2484_), .B(x6), .Y(men_men_n2485_));
  NA4        u2436(.A(men_men_n377_), .B(men_men_n260_), .C(men_men_n193_), .D(x8), .Y(men_men_n2486_));
  NA2        u2437(.A(men_men_n398_), .B(men_men_n107_), .Y(men_men_n2487_));
  AOI210     u2438(.A0(men_men_n2487_), .A1(men_men_n2486_), .B0(men_men_n143_), .Y(men_men_n2488_));
  AOI210     u2439(.A0(men_men_n432_), .A1(men_men_n403_), .B0(men_men_n1662_), .Y(men_men_n2489_));
  NO2        u2440(.A(men_men_n796_), .B(men_men_n91_), .Y(men_men_n2490_));
  OAI210     u2441(.A0(men_men_n988_), .A1(men_men_n150_), .B0(men_men_n358_), .Y(men_men_n2491_));
  OAI220     u2442(.A0(men_men_n2491_), .A1(men_men_n2490_), .B0(men_men_n2489_), .B1(men_men_n193_), .Y(men_men_n2492_));
  OAI210     u2443(.A0(men_men_n2492_), .A1(men_men_n2488_), .B0(x6), .Y(men_men_n2493_));
  NO2        u2444(.A(men_men_n250_), .B(men_men_n758_), .Y(men_men_n2494_));
  NO3        u2445(.A(men_men_n2494_), .B(men_men_n1617_), .C(men_men_n260_), .Y(men_men_n2495_));
  NO3        u2446(.A(x3), .B(men_men_n53_), .C(x0), .Y(men_men_n2496_));
  OAI210     u2447(.A0(men_men_n513_), .A1(x2), .B0(men_men_n2496_), .Y(men_men_n2497_));
  NA2        u2448(.A(men_men_n431_), .B(men_men_n422_), .Y(men_men_n2498_));
  NA3        u2449(.A(men_men_n2498_), .B(men_men_n2497_), .C(men_men_n1740_), .Y(men_men_n2499_));
  OAI210     u2450(.A0(men_men_n2499_), .A1(men_men_n2495_), .B0(men_men_n798_), .Y(men_men_n2500_));
  NO2        u2451(.A(men_men_n586_), .B(men_men_n279_), .Y(men_men_n2501_));
  AN3        u2452(.A(men_men_n803_), .B(men_men_n768_), .C(x0), .Y(men_men_n2502_));
  OAI210     u2453(.A0(men_men_n2502_), .A1(men_men_n2501_), .B0(men_men_n327_), .Y(men_men_n2503_));
  OAI220     u2454(.A0(men_men_n586_), .A1(men_men_n279_), .B0(men_men_n802_), .B1(men_men_n92_), .Y(men_men_n2504_));
  OAI210     u2455(.A0(men_men_n670_), .A1(x0), .B0(men_men_n51_), .Y(men_men_n2505_));
  AOI210     u2456(.A0(men_men_n567_), .A1(x4), .B0(men_men_n231_), .Y(men_men_n2506_));
  AOI220     u2457(.A0(men_men_n2506_), .A1(men_men_n2505_), .B0(men_men_n2504_), .B1(men_men_n400_), .Y(men_men_n2507_));
  NA4        u2458(.A(men_men_n2507_), .B(men_men_n2503_), .C(men_men_n2500_), .D(men_men_n2493_), .Y(men_men_n2508_));
  OAI210     u2459(.A0(men_men_n2508_), .A1(men_men_n2485_), .B0(x7), .Y(men_men_n2509_));
  AOI210     u2460(.A0(men_men_n373_), .A1(x1), .B0(men_men_n1187_), .Y(men_men_n2510_));
  NO2        u2461(.A(men_men_n2510_), .B(men_men_n51_), .Y(men_men_n2511_));
  AOI210     u2462(.A0(men_men_n91_), .A1(men_men_n71_), .B0(men_men_n2160_), .Y(men_men_n2512_));
  NA2        u2463(.A(men_men_n385_), .B(x3), .Y(men_men_n2513_));
  NO2        u2464(.A(men_men_n1683_), .B(men_men_n520_), .Y(men_men_n2514_));
  OAI210     u2465(.A0(men_men_n2513_), .A1(men_men_n2512_), .B0(men_men_n2514_), .Y(men_men_n2515_));
  OAI210     u2466(.A0(men_men_n2515_), .A1(men_men_n2511_), .B0(x4), .Y(men_men_n2516_));
  NO2        u2467(.A(men_men_n1694_), .B(men_men_n455_), .Y(men_men_n2517_));
  NO3        u2468(.A(men_men_n2517_), .B(men_men_n399_), .C(men_men_n120_), .Y(men_men_n2518_));
  AOI210     u2469(.A0(men_men_n1021_), .A1(men_men_n244_), .B0(men_men_n394_), .Y(men_men_n2519_));
  AO210      u2470(.A0(men_men_n1255_), .A1(x6), .B0(men_men_n2519_), .Y(men_men_n2520_));
  NO2        u2471(.A(men_men_n1367_), .B(men_men_n140_), .Y(men_men_n2521_));
  NA2        u2472(.A(men_men_n1882_), .B(men_men_n321_), .Y(men_men_n2522_));
  OAI220     u2473(.A0(men_men_n2522_), .A1(men_men_n1040_), .B0(men_men_n2521_), .B1(men_men_n1764_), .Y(men_men_n2523_));
  NO3        u2474(.A(men_men_n2523_), .B(men_men_n2520_), .C(men_men_n2518_), .Y(men_men_n2524_));
  AOI210     u2475(.A0(men_men_n2524_), .A1(men_men_n2516_), .B0(men_men_n107_), .Y(men_men_n2525_));
  NA3        u2476(.A(men_men_n1872_), .B(men_men_n586_), .C(men_men_n166_), .Y(men_men_n2526_));
  AOI210     u2477(.A0(men_men_n2526_), .A1(men_men_n1378_), .B0(men_men_n233_), .Y(men_men_n2527_));
  AOI210     u2478(.A0(men_men_n494_), .A1(men_men_n485_), .B0(men_men_n666_), .Y(men_men_n2528_));
  NO2        u2479(.A(men_men_n2528_), .B(men_men_n462_), .Y(men_men_n2529_));
  OAI210     u2480(.A0(men_men_n2529_), .A1(men_men_n2527_), .B0(x0), .Y(men_men_n2530_));
  NA3        u2481(.A(men_men_n403_), .B(men_men_n802_), .C(men_men_n279_), .Y(men_men_n2531_));
  AOI210     u2482(.A0(men_men_n2531_), .A1(men_men_n701_), .B0(men_men_n2124_), .Y(men_men_n2532_));
  NA2        u2483(.A(men_men_n1085_), .B(men_men_n929_), .Y(men_men_n2533_));
  NA4        u2484(.A(men_men_n665_), .B(men_men_n586_), .C(men_men_n181_), .D(x3), .Y(men_men_n2534_));
  AOI210     u2485(.A0(men_men_n2534_), .A1(men_men_n2533_), .B0(men_men_n491_), .Y(men_men_n2535_));
  NO4        u2486(.A(men_men_n1360_), .B(men_men_n509_), .C(men_men_n1182_), .D(men_men_n758_), .Y(men_men_n2536_));
  OAI220     u2487(.A0(men_men_n1712_), .A1(men_men_n2203_), .B0(men_men_n231_), .B1(men_men_n152_), .Y(men_men_n2537_));
  NO4        u2488(.A(men_men_n2537_), .B(men_men_n2536_), .C(men_men_n2535_), .D(men_men_n2532_), .Y(men_men_n2538_));
  NA2        u2489(.A(men_men_n2538_), .B(men_men_n2530_), .Y(men_men_n2539_));
  OAI210     u2490(.A0(men_men_n2539_), .A1(men_men_n2525_), .B0(men_men_n57_), .Y(men_men_n2540_));
  AOI210     u2491(.A0(men_men_n1751_), .A1(men_men_n279_), .B0(men_men_n667_), .Y(men_men_n2541_));
  OAI210     u2492(.A0(men_men_n1690_), .A1(men_men_n216_), .B0(men_men_n487_), .Y(men_men_n2542_));
  OAI210     u2493(.A0(men_men_n2542_), .A1(men_men_n2541_), .B0(men_men_n614_), .Y(men_men_n2543_));
  OAI220     u2494(.A0(men_men_n1697_), .A1(men_men_n279_), .B0(men_men_n259_), .B1(men_men_n103_), .Y(men_men_n2544_));
  NO2        u2495(.A(men_men_n677_), .B(men_men_n152_), .Y(men_men_n2545_));
  AOI210     u2496(.A0(men_men_n2544_), .A1(men_men_n962_), .B0(men_men_n2545_), .Y(men_men_n2546_));
  NA4        u2497(.A(men_men_n2546_), .B(men_men_n2543_), .C(men_men_n2540_), .D(men_men_n2509_), .Y(men39));
  INV        u2498(.A(men_men_n87_), .Y(men_men_n2550_));
  INV        u2499(.A(x1), .Y(men_men_n2551_));
  INV        u2500(.A(men_men_n160_), .Y(men_men_n2552_));
  INV        u2501(.A(x3), .Y(men_men_n2553_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
  VOTADOR g14(.A(ori14), .B(mai14), .C(men14), .Y(z14));
  VOTADOR g15(.A(ori15), .B(mai15), .C(men15), .Y(z15));
  VOTADOR g16(.A(ori16), .B(mai16), .C(men16), .Y(z16));
  VOTADOR g17(.A(ori17), .B(mai17), .C(men17), .Y(z17));
  VOTADOR g18(.A(ori18), .B(mai18), .C(men18), .Y(z18));
  VOTADOR g19(.A(ori19), .B(mai19), .C(men19), .Y(z19));
  VOTADOR g20(.A(ori20), .B(mai20), .C(men20), .Y(z20));
  VOTADOR g21(.A(ori21), .B(mai21), .C(men21), .Y(z21));
  VOTADOR g22(.A(ori22), .B(mai22), .C(men22), .Y(z22));
  VOTADOR g23(.A(ori23), .B(mai23), .C(men23), .Y(z23));
  VOTADOR g24(.A(ori24), .B(mai24), .C(men24), .Y(z24));
  VOTADOR g25(.A(ori25), .B(mai25), .C(men25), .Y(z25));
  VOTADOR g26(.A(ori26), .B(mai26), .C(men26), .Y(z26));
  VOTADOR g27(.A(ori27), .B(mai27), .C(men27), .Y(z27));
  VOTADOR g28(.A(ori28), .B(mai28), .C(men28), .Y(z28));
  VOTADOR g29(.A(ori29), .B(mai29), .C(men29), .Y(z29));
  VOTADOR g30(.A(ori30), .B(mai30), .C(men30), .Y(z30));
  VOTADOR g31(.A(ori31), .B(mai31), .C(men31), .Y(z31));
  VOTADOR g32(.A(ori32), .B(mai32), .C(men32), .Y(z32));
  VOTADOR g33(.A(ori33), .B(mai33), .C(men33), .Y(z33));
  VOTADOR g34(.A(ori34), .B(mai34), .C(men34), .Y(z34));
  VOTADOR g35(.A(ori35), .B(mai35), .C(men35), .Y(z35));
  VOTADOR g36(.A(ori36), .B(mai36), .C(men36), .Y(z36));
  VOTADOR g37(.A(ori37), .B(mai37), .C(men37), .Y(z37));
  VOTADOR g38(.A(ori38), .B(mai38), .C(men38), .Y(z38));
  VOTADOR g39(.A(ori39), .B(mai39), .C(men39), .Y(z39));
endmodule