library verilog;
use verilog.vl_types.all;
entity tb_full_adder is
end tb_full_adder;
