library verilog;
use verilog.vl_types.all;
entity contadorprimo_vlg_vec_tst is
end contadorprimo_vlg_vec_tst;
