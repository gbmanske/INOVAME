//  Class: spi_vseqr
//
class spi_vseqr extends uvm_component;
  `uvm_component_utils(spi_vseqr)


  //  Group: Components


  //  Group: Variables


  //  Group: Functions

  //  Constructor: new
  function new(string name = "spi_vseqr", uvm_component parent);
    super.new(name, parent);
  endfunction: new


endclass: spi_vseqr
