// Benchmark "top" written by ABC on Fri Jun 21 17:49:28 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n139_,
    new_new_n140_, new_new_n141_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1042_, new_new_n1043_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g0062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g0063(.A(i_6_), .Y(new_new_n86_));
  OR4        g0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g0065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g0066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  NO2        g0067(.A(new_new_n88_), .B(new_new_n89_), .Y(new_new_n90_));
  OAI210     g0068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g0069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g0070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g0071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g0072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  INV        g0073(.A(new_new_n94_), .Y(new_new_n96_));
  AOI210     g0074(.A0(new_new_n96_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n97_));
  AN3        g0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g0076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g0077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NOi21      g0078(.An(new_new_n100_), .B(new_new_n99_), .Y(new_new_n101_));
  AOI220     g0079(.A0(new_new_n101_), .A1(new_new_n62_), .B0(new_new_n98_), .B1(new_new_n32_), .Y(new_new_n102_));
  INV        g0080(.A(i_7_), .Y(new_new_n103_));
  NA2        g0081(.A(new_new_n47_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g0082(.A(i_0_), .B(i_5_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(new_new_n86_), .Y(new_new_n106_));
  NA2        g0084(.A(i_12_), .B(i_3_), .Y(new_new_n107_));
  INV        g0085(.A(new_new_n107_), .Y(new_new_n108_));
  NA3        g0086(.A(new_new_n108_), .B(new_new_n106_), .C(new_new_n104_), .Y(new_new_n109_));
  NAi21      g0087(.An(i_7_), .B(i_11_), .Y(new_new_n110_));
  NO3        g0088(.A(new_new_n110_), .B(new_new_n92_), .C(new_new_n54_), .Y(new_new_n111_));
  AN2        g0089(.A(i_2_), .B(i_10_), .Y(new_new_n112_));
  NO2        g0090(.A(new_new_n112_), .B(i_7_), .Y(new_new_n113_));
  OR2        g0091(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n114_));
  NO2        g0092(.A(i_8_), .B(new_new_n103_), .Y(new_new_n115_));
  NO3        g0093(.A(new_new_n115_), .B(new_new_n114_), .C(new_new_n113_), .Y(new_new_n116_));
  NA2        g0094(.A(i_12_), .B(i_7_), .Y(new_new_n117_));
  NO2        g0095(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n118_));
  NA2        g0096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n1043_), .B(new_new_n116_), .Y(new_new_n120_));
  NAi41      g0098(.An(new_new_n111_), .B(new_new_n120_), .C(new_new_n109_), .D(new_new_n102_), .Y(new_new_n121_));
  NOi21      g0099(.An(i_1_), .B(i_5_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(i_11_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n124_));
  NA2        g0102(.A(i_7_), .B(new_new_n25_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(new_new_n124_), .Y(new_new_n126_));
  NO2        g0104(.A(new_new_n126_), .B(new_new_n47_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n128_));
  NAi21      g0106(.An(i_3_), .B(i_8_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n129_), .B(new_new_n62_), .Y(new_new_n130_));
  NOi31      g0108(.An(new_new_n130_), .B(new_new_n128_), .C(new_new_n127_), .Y(new_new_n131_));
  NO2        g0109(.A(i_1_), .B(new_new_n86_), .Y(new_new_n132_));
  NO2        g0110(.A(i_6_), .B(i_5_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(i_3_), .Y(new_new_n134_));
  AO210      g0112(.A0(new_new_n134_), .A1(new_new_n48_), .B0(new_new_n132_), .Y(new_new_n135_));
  OAI220     g0113(.A0(new_new_n135_), .A1(new_new_n110_), .B0(new_new_n131_), .B1(new_new_n123_), .Y(new_new_n136_));
  NO3        g0114(.A(new_new_n136_), .B(new_new_n121_), .C(new_new_n97_), .Y(new_new_n137_));
  NA3        g0115(.A(new_new_n137_), .B(new_new_n79_), .C(new_new_n56_), .Y(men2));
  NO2        g0116(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n139_));
  NA2        g0117(.A(i_6_), .B(new_new_n25_), .Y(new_new_n140_));
  NA2        g0118(.A(new_new_n140_), .B(new_new_n139_), .Y(new_new_n141_));
  NA4        g0119(.A(new_new_n141_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(men0));
  AN2        g0120(.A(i_8_), .B(i_7_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(i_6_), .Y(new_new_n144_));
  NO2        g0122(.A(i_12_), .B(i_13_), .Y(new_new_n145_));
  NAi21      g0123(.An(i_5_), .B(i_11_), .Y(new_new_n146_));
  NOi21      g0124(.An(new_new_n145_), .B(new_new_n146_), .Y(new_new_n147_));
  NO2        g0125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NA2        g0126(.A(i_2_), .B(i_3_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n149_), .B(i_4_), .Y(new_new_n150_));
  NA3        g0128(.A(new_new_n150_), .B(new_new_n148_), .C(new_new_n147_), .Y(new_new_n151_));
  AN2        g0129(.A(new_new_n145_), .B(new_new_n83_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(new_new_n27_), .Y(new_new_n153_));
  NA2        g0131(.A(i_1_), .B(i_5_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n155_));
  NA2        g0133(.A(new_new_n155_), .B(new_new_n36_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n156_), .B(new_new_n154_), .C(new_new_n153_), .Y(new_new_n157_));
  OR2        g0135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n159_));
  NAi32      g0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n160_));
  NAi21      g0138(.An(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NOi21      g0139(.An(i_4_), .B(i_10_), .Y(new_new_n162_));
  NA2        g0140(.A(new_new_n162_), .B(new_new_n40_), .Y(new_new_n163_));
  NO2        g0141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  NO3        g0142(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OAI210     g0144(.A0(new_new_n166_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n167_));
  NO2        g0145(.A(new_new_n167_), .B(new_new_n157_), .Y(new_new_n168_));
  AOI210     g0146(.A0(new_new_n168_), .A1(new_new_n151_), .B0(new_new_n144_), .Y(new_new_n169_));
  NA3        g0147(.A(new_new_n73_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n170_));
  NA2        g0148(.A(i_3_), .B(new_new_n49_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_4_), .B(i_9_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_11_), .B(i_13_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n173_), .B(new_new_n172_), .Y(new_new_n174_));
  NO2        g0152(.A(i_4_), .B(i_5_), .Y(new_new_n175_));
  NAi21      g0153(.An(i_12_), .B(i_11_), .Y(new_new_n176_));
  NO2        g0154(.A(new_new_n176_), .B(i_13_), .Y(new_new_n177_));
  NA3        g0155(.A(new_new_n177_), .B(new_new_n175_), .C(new_new_n83_), .Y(new_new_n178_));
  AOI210     g0156(.A0(new_new_n178_), .A1(new_new_n174_), .B0(new_new_n170_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n180_));
  NA2        g0158(.A(new_new_n180_), .B(new_new_n47_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n36_), .B(i_5_), .Y(new_new_n182_));
  NAi31      g0160(.An(new_new_n182_), .B(new_new_n152_), .C(i_11_), .Y(new_new_n183_));
  NA2        g0161(.A(i_3_), .B(i_5_), .Y(new_new_n184_));
  OR2        g0162(.A(new_new_n184_), .B(new_new_n174_), .Y(new_new_n185_));
  AOI210     g0163(.A0(new_new_n185_), .A1(new_new_n183_), .B0(new_new_n181_), .Y(new_new_n186_));
  NO2        g0164(.A(new_new_n73_), .B(i_5_), .Y(new_new_n187_));
  NO2        g0165(.A(i_13_), .B(i_10_), .Y(new_new_n188_));
  NA3        g0166(.A(new_new_n188_), .B(new_new_n187_), .C(new_new_n45_), .Y(new_new_n189_));
  NO2        g0167(.A(i_2_), .B(i_1_), .Y(new_new_n190_));
  NA2        g0168(.A(new_new_n190_), .B(i_3_), .Y(new_new_n191_));
  NAi21      g0169(.An(i_4_), .B(i_12_), .Y(new_new_n192_));
  NO4        g0170(.A(new_new_n192_), .B(new_new_n191_), .C(new_new_n189_), .D(new_new_n25_), .Y(new_new_n193_));
  NO3        g0171(.A(new_new_n193_), .B(new_new_n186_), .C(new_new_n179_), .Y(new_new_n194_));
  INV        g0172(.A(i_8_), .Y(new_new_n195_));
  NO2        g0173(.A(new_new_n195_), .B(i_7_), .Y(new_new_n196_));
  NA2        g0174(.A(new_new_n196_), .B(i_6_), .Y(new_new_n197_));
  NO3        g0175(.A(i_3_), .B(new_new_n86_), .C(new_new_n49_), .Y(new_new_n198_));
  NA2        g0176(.A(new_new_n198_), .B(new_new_n115_), .Y(new_new_n199_));
  NO3        g0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n200_));
  NA3        g0178(.A(new_new_n200_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n201_));
  NO3        g0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n202_));
  OAI210     g0180(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n202_), .Y(new_new_n203_));
  AOI210     g0181(.A0(new_new_n203_), .A1(new_new_n201_), .B0(new_new_n199_), .Y(new_new_n204_));
  NO2        g0182(.A(i_3_), .B(i_8_), .Y(new_new_n205_));
  NO3        g0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n206_));
  NO2        g0184(.A(new_new_n105_), .B(new_new_n58_), .Y(new_new_n207_));
  NO2        g0185(.A(i_13_), .B(i_9_), .Y(new_new_n208_));
  NA3        g0186(.A(new_new_n208_), .B(i_6_), .C(new_new_n195_), .Y(new_new_n209_));
  NAi21      g0187(.An(i_12_), .B(i_3_), .Y(new_new_n210_));
  NO2        g0188(.A(new_new_n45_), .B(i_5_), .Y(new_new_n211_));
  NO3        g0189(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n212_));
  NA3        g0190(.A(new_new_n212_), .B(new_new_n211_), .C(i_10_), .Y(new_new_n213_));
  NO2        g0191(.A(new_new_n213_), .B(new_new_n209_), .Y(new_new_n214_));
  AOI210     g0192(.A0(new_new_n214_), .A1(i_7_), .B0(new_new_n204_), .Y(new_new_n215_));
  OAI220     g0193(.A0(new_new_n215_), .A1(i_4_), .B0(new_new_n197_), .B1(new_new_n194_), .Y(new_new_n216_));
  NAi21      g0194(.An(i_12_), .B(i_7_), .Y(new_new_n217_));
  NA3        g0195(.A(i_13_), .B(new_new_n195_), .C(i_10_), .Y(new_new_n218_));
  NA2        g0196(.A(i_0_), .B(i_5_), .Y(new_new_n219_));
  NAi31      g0197(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n220_));
  NO2        g0198(.A(new_new_n36_), .B(i_13_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n223_));
  NA3        g0201(.A(new_new_n223_), .B(new_new_n222_), .C(new_new_n221_), .Y(new_new_n224_));
  INV        g0202(.A(i_13_), .Y(new_new_n225_));
  NO2        g0203(.A(i_12_), .B(new_new_n225_), .Y(new_new_n226_));
  NA3        g0204(.A(new_new_n226_), .B(new_new_n200_), .C(new_new_n198_), .Y(new_new_n227_));
  OAI210     g0205(.A0(new_new_n224_), .A1(new_new_n220_), .B0(new_new_n227_), .Y(new_new_n228_));
  NA2        g0206(.A(new_new_n228_), .B(new_new_n143_), .Y(new_new_n229_));
  NO2        g0207(.A(i_12_), .B(new_new_n37_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n184_), .B(i_4_), .Y(new_new_n231_));
  NA2        g0209(.A(new_new_n231_), .B(new_new_n230_), .Y(new_new_n232_));
  OR2        g0210(.A(i_8_), .B(i_7_), .Y(new_new_n233_));
  NO2        g0211(.A(new_new_n233_), .B(new_new_n86_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n54_), .B(i_1_), .Y(new_new_n235_));
  NA2        g0213(.A(new_new_n235_), .B(new_new_n234_), .Y(new_new_n236_));
  INV        g0214(.A(i_12_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n45_), .B(new_new_n237_), .Y(new_new_n238_));
  NO3        g0216(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n239_));
  NA2        g0217(.A(i_2_), .B(i_1_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n236_), .B(new_new_n232_), .Y(new_new_n241_));
  NO3        g0219(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n242_));
  NAi21      g0220(.An(i_4_), .B(i_3_), .Y(new_new_n243_));
  NO2        g0221(.A(i_0_), .B(i_6_), .Y(new_new_n244_));
  NOi41      g0222(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n245_));
  NA2        g0223(.A(new_new_n245_), .B(new_new_n244_), .Y(new_new_n246_));
  NO2        g0224(.A(new_new_n240_), .B(new_new_n184_), .Y(new_new_n247_));
  NAi21      g0225(.An(new_new_n246_), .B(new_new_n247_), .Y(new_new_n248_));
  INV        g0226(.A(new_new_n248_), .Y(new_new_n249_));
  AOI220     g0227(.A0(new_new_n249_), .A1(new_new_n40_), .B0(new_new_n241_), .B1(new_new_n208_), .Y(new_new_n250_));
  NO2        g0228(.A(i_11_), .B(new_new_n225_), .Y(new_new_n251_));
  NOi21      g0229(.An(i_1_), .B(i_6_), .Y(new_new_n252_));
  NAi21      g0230(.An(i_3_), .B(i_7_), .Y(new_new_n253_));
  NA2        g0231(.A(new_new_n237_), .B(i_9_), .Y(new_new_n254_));
  OR4        g0232(.A(new_new_n254_), .B(new_new_n253_), .C(new_new_n252_), .D(new_new_n187_), .Y(new_new_n255_));
  NO2        g0233(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n256_));
  NO2        g0234(.A(i_12_), .B(i_3_), .Y(new_new_n257_));
  NA2        g0235(.A(new_new_n73_), .B(i_5_), .Y(new_new_n258_));
  NA2        g0236(.A(i_3_), .B(i_9_), .Y(new_new_n259_));
  NAi21      g0237(.An(i_7_), .B(i_10_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n260_), .B(new_new_n259_), .Y(new_new_n261_));
  INV        g0239(.A(new_new_n255_), .Y(new_new_n262_));
  NA3        g0240(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n263_));
  INV        g0241(.A(new_new_n144_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n237_), .B(i_13_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n75_), .Y(new_new_n266_));
  AOI220     g0244(.A0(new_new_n266_), .A1(new_new_n264_), .B0(new_new_n262_), .B1(new_new_n251_), .Y(new_new_n267_));
  NO2        g0245(.A(new_new_n233_), .B(new_new_n37_), .Y(new_new_n268_));
  NA2        g0246(.A(i_12_), .B(i_6_), .Y(new_new_n269_));
  OR2        g0247(.A(i_13_), .B(i_9_), .Y(new_new_n270_));
  NO3        g0248(.A(new_new_n270_), .B(new_new_n269_), .C(new_new_n49_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n243_), .B(i_2_), .Y(new_new_n272_));
  NA3        g0250(.A(new_new_n272_), .B(new_new_n271_), .C(new_new_n45_), .Y(new_new_n273_));
  NA2        g0251(.A(new_new_n251_), .B(i_9_), .Y(new_new_n274_));
  NA2        g0252(.A(new_new_n258_), .B(new_new_n64_), .Y(new_new_n275_));
  OAI210     g0253(.A0(new_new_n275_), .A1(new_new_n274_), .B0(new_new_n273_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n155_), .B(new_new_n63_), .Y(new_new_n277_));
  NO3        g0255(.A(i_11_), .B(new_new_n225_), .C(new_new_n25_), .Y(new_new_n278_));
  NO2        g0256(.A(new_new_n253_), .B(i_8_), .Y(new_new_n279_));
  NO2        g0257(.A(i_6_), .B(new_new_n49_), .Y(new_new_n280_));
  NA3        g0258(.A(new_new_n280_), .B(new_new_n279_), .C(new_new_n278_), .Y(new_new_n281_));
  NO3        g0259(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n282_));
  NA3        g0260(.A(new_new_n282_), .B(new_new_n268_), .C(new_new_n226_), .Y(new_new_n283_));
  AOI210     g0261(.A0(new_new_n283_), .A1(new_new_n281_), .B0(new_new_n277_), .Y(new_new_n284_));
  AOI210     g0262(.A0(new_new_n276_), .A1(new_new_n268_), .B0(new_new_n284_), .Y(new_new_n285_));
  NA4        g0263(.A(new_new_n285_), .B(new_new_n267_), .C(new_new_n250_), .D(new_new_n229_), .Y(new_new_n286_));
  NO3        g0264(.A(i_12_), .B(new_new_n225_), .C(new_new_n37_), .Y(new_new_n287_));
  INV        g0265(.A(new_new_n287_), .Y(new_new_n288_));
  NA2        g0266(.A(i_8_), .B(new_new_n103_), .Y(new_new_n289_));
  NO3        g0267(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n240_), .B(i_0_), .Y(new_new_n291_));
  NA2        g0269(.A(i_0_), .B(i_1_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n292_), .B(i_2_), .Y(new_new_n293_));
  NO2        g0271(.A(new_new_n59_), .B(i_6_), .Y(new_new_n294_));
  NA3        g0272(.A(new_new_n294_), .B(new_new_n293_), .C(new_new_n164_), .Y(new_new_n295_));
  NO2        g0273(.A(i_3_), .B(i_10_), .Y(new_new_n296_));
  NA3        g0274(.A(new_new_n296_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n297_));
  NO2        g0275(.A(i_2_), .B(new_new_n103_), .Y(new_new_n298_));
  NA2        g0276(.A(i_1_), .B(new_new_n36_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n299_), .B(i_8_), .Y(new_new_n300_));
  NA2        g0278(.A(new_new_n300_), .B(new_new_n298_), .Y(new_new_n301_));
  AN2        g0279(.A(i_3_), .B(i_10_), .Y(new_new_n302_));
  NA4        g0280(.A(new_new_n302_), .B(new_new_n200_), .C(new_new_n177_), .D(new_new_n175_), .Y(new_new_n303_));
  NO2        g0281(.A(i_5_), .B(new_new_n37_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n305_));
  OR2        g0283(.A(new_new_n301_), .B(new_new_n297_), .Y(new_new_n306_));
  OAI220     g0284(.A0(new_new_n306_), .A1(i_6_), .B0(new_new_n295_), .B1(new_new_n288_), .Y(new_new_n307_));
  NO4        g0285(.A(new_new_n307_), .B(new_new_n286_), .C(new_new_n216_), .D(new_new_n169_), .Y(new_new_n308_));
  NO3        g0286(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n309_));
  NO2        g0287(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n310_));
  NA2        g0288(.A(new_new_n291_), .B(new_new_n310_), .Y(new_new_n311_));
  NO3        g0289(.A(i_6_), .B(new_new_n195_), .C(i_7_), .Y(new_new_n312_));
  NA2        g0290(.A(new_new_n312_), .B(new_new_n200_), .Y(new_new_n313_));
  AOI210     g0291(.A0(new_new_n313_), .A1(new_new_n311_), .B0(new_new_n171_), .Y(new_new_n314_));
  NO2        g0292(.A(i_2_), .B(i_3_), .Y(new_new_n315_));
  OR2        g0293(.A(i_0_), .B(i_5_), .Y(new_new_n316_));
  NA2        g0294(.A(new_new_n219_), .B(new_new_n316_), .Y(new_new_n317_));
  NO2        g0295(.A(i_8_), .B(i_6_), .Y(new_new_n318_));
  NO2        g0296(.A(new_new_n158_), .B(new_new_n47_), .Y(new_new_n319_));
  NA3        g0297(.A(new_new_n319_), .B(new_new_n318_), .C(new_new_n164_), .Y(new_new_n320_));
  INV        g0298(.A(new_new_n320_), .Y(new_new_n321_));
  OAI210     g0299(.A0(new_new_n321_), .A1(new_new_n314_), .B0(i_4_), .Y(new_new_n322_));
  NO2        g0300(.A(i_12_), .B(i_10_), .Y(new_new_n323_));
  NOi21      g0301(.An(i_5_), .B(i_0_), .Y(new_new_n324_));
  NO3        g0302(.A(new_new_n299_), .B(new_new_n324_), .C(new_new_n129_), .Y(new_new_n325_));
  NA4        g0303(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n326_));
  NA2        g0304(.A(new_new_n325_), .B(new_new_n323_), .Y(new_new_n327_));
  NO2        g0305(.A(i_6_), .B(i_8_), .Y(new_new_n328_));
  NOi21      g0306(.An(i_0_), .B(i_2_), .Y(new_new_n329_));
  AN2        g0307(.A(new_new_n329_), .B(new_new_n328_), .Y(new_new_n330_));
  NO2        g0308(.A(i_1_), .B(i_7_), .Y(new_new_n331_));
  AO220      g0309(.A0(new_new_n331_), .A1(new_new_n330_), .B0(new_new_n318_), .B1(new_new_n235_), .Y(new_new_n332_));
  NA3        g0310(.A(new_new_n332_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n333_));
  NA3        g0311(.A(new_new_n333_), .B(new_new_n327_), .C(new_new_n322_), .Y(new_new_n334_));
  NO3        g0312(.A(new_new_n233_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n335_));
  NO3        g0313(.A(i_8_), .B(i_2_), .C(i_1_), .Y(new_new_n336_));
  OAI210     g0314(.A0(new_new_n336_), .A1(new_new_n335_), .B0(i_6_), .Y(new_new_n337_));
  NO2        g0315(.A(new_new_n337_), .B(new_new_n317_), .Y(new_new_n338_));
  NOi21      g0316(.An(new_new_n154_), .B(new_new_n106_), .Y(new_new_n339_));
  NO2        g0317(.A(new_new_n339_), .B(new_new_n125_), .Y(new_new_n340_));
  OAI210     g0318(.A0(new_new_n340_), .A1(new_new_n338_), .B0(i_3_), .Y(new_new_n341_));
  INV        g0319(.A(new_new_n84_), .Y(new_new_n342_));
  NO2        g0320(.A(new_new_n292_), .B(new_new_n81_), .Y(new_new_n343_));
  NA2        g0321(.A(new_new_n343_), .B(new_new_n133_), .Y(new_new_n344_));
  NO2        g0322(.A(new_new_n95_), .B(new_new_n195_), .Y(new_new_n345_));
  NA2        g0323(.A(new_new_n345_), .B(new_new_n63_), .Y(new_new_n346_));
  AOI210     g0324(.A0(new_new_n346_), .A1(new_new_n344_), .B0(new_new_n342_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n195_), .B(i_9_), .Y(new_new_n348_));
  NA2        g0326(.A(new_new_n348_), .B(new_new_n207_), .Y(new_new_n349_));
  NO2        g0327(.A(new_new_n349_), .B(new_new_n47_), .Y(new_new_n350_));
  NO2        g0328(.A(new_new_n350_), .B(new_new_n347_), .Y(new_new_n351_));
  AOI210     g0329(.A0(new_new_n351_), .A1(new_new_n341_), .B0(new_new_n163_), .Y(new_new_n352_));
  AOI210     g0330(.A0(new_new_n334_), .A1(new_new_n309_), .B0(new_new_n352_), .Y(new_new_n353_));
  NOi32      g0331(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n354_));
  INV        g0332(.A(new_new_n354_), .Y(new_new_n355_));
  NAi21      g0333(.An(i_0_), .B(i_6_), .Y(new_new_n356_));
  NAi21      g0334(.An(i_1_), .B(i_5_), .Y(new_new_n357_));
  NA2        g0335(.A(new_new_n357_), .B(new_new_n356_), .Y(new_new_n358_));
  NA2        g0336(.A(new_new_n358_), .B(new_new_n25_), .Y(new_new_n359_));
  OAI210     g0337(.A0(new_new_n359_), .A1(new_new_n160_), .B0(new_new_n246_), .Y(new_new_n360_));
  NAi41      g0338(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n361_));
  AOI210     g0339(.A0(new_new_n361_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n362_));
  NOi32      g0340(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n363_));
  NO2        g0341(.A(i_1_), .B(new_new_n103_), .Y(new_new_n364_));
  NAi21      g0342(.An(i_3_), .B(i_4_), .Y(new_new_n365_));
  NO2        g0343(.A(new_new_n365_), .B(i_9_), .Y(new_new_n366_));
  AN2        g0344(.A(i_6_), .B(i_7_), .Y(new_new_n367_));
  OAI210     g0345(.A0(new_new_n367_), .A1(new_new_n364_), .B0(new_new_n366_), .Y(new_new_n368_));
  NA2        g0346(.A(i_2_), .B(i_7_), .Y(new_new_n369_));
  NO2        g0347(.A(new_new_n365_), .B(i_10_), .Y(new_new_n370_));
  NO2        g0348(.A(new_new_n368_), .B(new_new_n187_), .Y(new_new_n371_));
  AOI210     g0349(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n372_));
  OAI210     g0350(.A0(new_new_n372_), .A1(new_new_n190_), .B0(new_new_n370_), .Y(new_new_n373_));
  NO2        g0351(.A(new_new_n373_), .B(i_5_), .Y(new_new_n374_));
  NO4        g0352(.A(new_new_n374_), .B(new_new_n371_), .C(new_new_n362_), .D(new_new_n360_), .Y(new_new_n375_));
  NO2        g0353(.A(new_new_n375_), .B(new_new_n355_), .Y(new_new_n376_));
  NO2        g0354(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n377_));
  AN2        g0355(.A(i_12_), .B(i_5_), .Y(new_new_n378_));
  NO2        g0356(.A(i_4_), .B(new_new_n26_), .Y(new_new_n379_));
  NA2        g0357(.A(new_new_n379_), .B(new_new_n378_), .Y(new_new_n380_));
  NO2        g0358(.A(i_11_), .B(i_6_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n243_), .B(i_5_), .Y(new_new_n382_));
  NO2        g0360(.A(i_5_), .B(i_10_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n384_));
  NO3        g0362(.A(new_new_n86_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n385_));
  NO2        g0363(.A(i_3_), .B(new_new_n103_), .Y(new_new_n386_));
  NO2        g0364(.A(i_11_), .B(i_12_), .Y(new_new_n387_));
  NA2        g0365(.A(new_new_n383_), .B(new_new_n237_), .Y(new_new_n388_));
  NA3        g0366(.A(new_new_n115_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n389_));
  OAI220     g0367(.A0(new_new_n389_), .A1(new_new_n220_), .B0(new_new_n388_), .B1(new_new_n326_), .Y(new_new_n390_));
  NAi21      g0368(.An(i_13_), .B(i_0_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(new_new_n240_), .Y(new_new_n392_));
  NA2        g0370(.A(new_new_n390_), .B(new_new_n392_), .Y(new_new_n393_));
  INV        g0371(.A(new_new_n393_), .Y(new_new_n394_));
  NO3        g0372(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n395_));
  NO2        g0373(.A(i_0_), .B(i_11_), .Y(new_new_n396_));
  INV        g0374(.A(i_5_), .Y(new_new_n397_));
  AN2        g0375(.A(i_1_), .B(i_6_), .Y(new_new_n398_));
  NOi21      g0376(.An(i_2_), .B(i_12_), .Y(new_new_n399_));
  NA2        g0377(.A(new_new_n399_), .B(new_new_n398_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n400_), .B(new_new_n397_), .Y(new_new_n401_));
  NA2        g0379(.A(new_new_n143_), .B(i_9_), .Y(new_new_n402_));
  NO2        g0380(.A(new_new_n402_), .B(i_4_), .Y(new_new_n403_));
  NA2        g0381(.A(new_new_n401_), .B(new_new_n403_), .Y(new_new_n404_));
  NAi21      g0382(.An(i_9_), .B(i_4_), .Y(new_new_n405_));
  OR2        g0383(.A(i_13_), .B(i_10_), .Y(new_new_n406_));
  NO3        g0384(.A(new_new_n406_), .B(new_new_n119_), .C(new_new_n405_), .Y(new_new_n407_));
  OR2        g0385(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n103_), .B(new_new_n25_), .Y(new_new_n409_));
  NA2        g0387(.A(new_new_n287_), .B(new_new_n409_), .Y(new_new_n410_));
  NA2        g0388(.A(new_new_n280_), .B(new_new_n212_), .Y(new_new_n411_));
  OAI220     g0389(.A0(new_new_n411_), .A1(new_new_n408_), .B0(new_new_n410_), .B1(new_new_n339_), .Y(new_new_n412_));
  INV        g0390(.A(new_new_n412_), .Y(new_new_n413_));
  AOI210     g0391(.A0(new_new_n413_), .A1(new_new_n404_), .B0(new_new_n26_), .Y(new_new_n414_));
  AOI220     g0392(.A0(new_new_n294_), .A1(new_new_n290_), .B0(new_new_n291_), .B1(new_new_n310_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n415_), .B(new_new_n171_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n184_), .B(new_new_n86_), .Y(new_new_n417_));
  AOI220     g0395(.A0(new_new_n417_), .A1(new_new_n293_), .B0(new_new_n282_), .B1(new_new_n212_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n418_), .B(new_new_n289_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n419_), .B(new_new_n416_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n195_), .B(i_10_), .Y(new_new_n421_));
  NA3        g0399(.A(new_new_n258_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n422_));
  NA2        g0400(.A(new_new_n294_), .B(new_new_n235_), .Y(new_new_n423_));
  OAI220     g0401(.A0(new_new_n423_), .A1(new_new_n184_), .B0(new_new_n422_), .B1(new_new_n421_), .Y(new_new_n424_));
  NO2        g0402(.A(i_3_), .B(new_new_n49_), .Y(new_new_n425_));
  NA3        g0403(.A(new_new_n331_), .B(new_new_n330_), .C(new_new_n425_), .Y(new_new_n426_));
  NA2        g0404(.A(new_new_n312_), .B(new_new_n317_), .Y(new_new_n427_));
  OAI210     g0405(.A0(new_new_n427_), .A1(new_new_n191_), .B0(new_new_n426_), .Y(new_new_n428_));
  NO2        g0406(.A(new_new_n428_), .B(new_new_n424_), .Y(new_new_n429_));
  AOI210     g0407(.A0(new_new_n429_), .A1(new_new_n420_), .B0(new_new_n274_), .Y(new_new_n430_));
  NO4        g0408(.A(new_new_n430_), .B(new_new_n414_), .C(new_new_n394_), .D(new_new_n376_), .Y(new_new_n431_));
  NO2        g0409(.A(new_new_n63_), .B(i_4_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n73_), .B(i_13_), .Y(new_new_n433_));
  NO2        g0411(.A(i_10_), .B(i_9_), .Y(new_new_n434_));
  NAi21      g0412(.An(i_12_), .B(i_8_), .Y(new_new_n435_));
  NO2        g0413(.A(new_new_n435_), .B(i_3_), .Y(new_new_n436_));
  NA2        g0414(.A(new_new_n305_), .B(i_0_), .Y(new_new_n437_));
  NO3        g0415(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n269_), .B(new_new_n99_), .Y(new_new_n439_));
  NA2        g0417(.A(new_new_n439_), .B(new_new_n438_), .Y(new_new_n440_));
  NA2        g0418(.A(i_8_), .B(i_9_), .Y(new_new_n441_));
  AOI210     g0419(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n442_));
  OR2        g0420(.A(new_new_n442_), .B(new_new_n441_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n287_), .B(new_new_n207_), .Y(new_new_n444_));
  OAI220     g0422(.A0(new_new_n444_), .A1(new_new_n443_), .B0(new_new_n440_), .B1(new_new_n437_), .Y(new_new_n445_));
  NA2        g0423(.A(new_new_n251_), .B(new_new_n304_), .Y(new_new_n446_));
  NO3        g0424(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n447_));
  INV        g0425(.A(new_new_n447_), .Y(new_new_n448_));
  NA3        g0426(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n449_));
  NA4        g0427(.A(new_new_n146_), .B(new_new_n118_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n450_));
  OAI220     g0428(.A0(new_new_n450_), .A1(new_new_n449_), .B0(new_new_n448_), .B1(new_new_n446_), .Y(new_new_n451_));
  NO2        g0429(.A(new_new_n451_), .B(new_new_n445_), .Y(new_new_n452_));
  INV        g0430(.A(new_new_n293_), .Y(new_new_n453_));
  OR2        g0431(.A(new_new_n453_), .B(new_new_n209_), .Y(new_new_n454_));
  OA210      g0432(.A0(new_new_n349_), .A1(new_new_n103_), .B0(new_new_n295_), .Y(new_new_n455_));
  OA220      g0433(.A0(new_new_n455_), .A1(new_new_n163_), .B0(new_new_n454_), .B1(new_new_n232_), .Y(new_new_n456_));
  NA2        g0434(.A(new_new_n98_), .B(i_13_), .Y(new_new_n457_));
  NO2        g0435(.A(i_2_), .B(i_13_), .Y(new_new_n458_));
  NO3        g0436(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n459_));
  NO2        g0437(.A(i_6_), .B(i_7_), .Y(new_new_n460_));
  NA2        g0438(.A(new_new_n460_), .B(new_new_n459_), .Y(new_new_n461_));
  NO2        g0439(.A(i_11_), .B(i_1_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n73_), .B(i_3_), .Y(new_new_n463_));
  OR2        g0441(.A(i_11_), .B(i_8_), .Y(new_new_n464_));
  NOi21      g0442(.An(i_2_), .B(i_7_), .Y(new_new_n465_));
  NAi31      g0443(.An(new_new_n464_), .B(new_new_n465_), .C(new_new_n463_), .Y(new_new_n466_));
  NO2        g0444(.A(new_new_n406_), .B(i_6_), .Y(new_new_n467_));
  NA2        g0445(.A(new_new_n467_), .B(new_new_n432_), .Y(new_new_n468_));
  NO2        g0446(.A(new_new_n468_), .B(new_new_n466_), .Y(new_new_n469_));
  NO2        g0447(.A(i_3_), .B(new_new_n195_), .Y(new_new_n470_));
  NO2        g0448(.A(i_6_), .B(i_10_), .Y(new_new_n471_));
  NA4        g0449(.A(new_new_n471_), .B(new_new_n309_), .C(new_new_n470_), .D(new_new_n237_), .Y(new_new_n472_));
  NO2        g0450(.A(new_new_n472_), .B(new_new_n156_), .Y(new_new_n473_));
  NA3        g0451(.A(new_new_n245_), .B(new_new_n173_), .C(new_new_n133_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n158_), .B(i_3_), .Y(new_new_n476_));
  NAi31      g0454(.An(new_new_n475_), .B(new_new_n476_), .C(new_new_n226_), .Y(new_new_n477_));
  NA3        g0455(.A(new_new_n384_), .B(new_new_n180_), .C(new_new_n150_), .Y(new_new_n478_));
  NA3        g0456(.A(new_new_n478_), .B(new_new_n477_), .C(new_new_n474_), .Y(new_new_n479_));
  NO3        g0457(.A(new_new_n479_), .B(new_new_n473_), .C(new_new_n469_), .Y(new_new_n480_));
  NA2        g0458(.A(new_new_n438_), .B(new_new_n378_), .Y(new_new_n481_));
  NA2        g0459(.A(new_new_n447_), .B(new_new_n383_), .Y(new_new_n482_));
  NO2        g0460(.A(new_new_n482_), .B(new_new_n224_), .Y(new_new_n483_));
  NAi21      g0461(.An(new_new_n218_), .B(new_new_n387_), .Y(new_new_n484_));
  NA2        g0462(.A(new_new_n331_), .B(new_new_n219_), .Y(new_new_n485_));
  NO2        g0463(.A(new_new_n26_), .B(i_5_), .Y(new_new_n486_));
  NO2        g0464(.A(i_0_), .B(new_new_n86_), .Y(new_new_n487_));
  NA3        g0465(.A(new_new_n487_), .B(new_new_n486_), .C(new_new_n143_), .Y(new_new_n488_));
  OR3        g0466(.A(new_new_n299_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n489_));
  OAI220     g0467(.A0(new_new_n489_), .A1(new_new_n488_), .B0(new_new_n485_), .B1(new_new_n484_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n27_), .B(i_10_), .Y(new_new_n491_));
  NA2        g0469(.A(new_new_n309_), .B(new_new_n239_), .Y(new_new_n492_));
  OAI220     g0470(.A0(new_new_n492_), .A1(new_new_n422_), .B0(new_new_n491_), .B1(new_new_n457_), .Y(new_new_n493_));
  NA4        g0471(.A(new_new_n302_), .B(new_new_n223_), .C(new_new_n73_), .D(new_new_n237_), .Y(new_new_n494_));
  NO2        g0472(.A(new_new_n494_), .B(new_new_n461_), .Y(new_new_n495_));
  NO4        g0473(.A(new_new_n495_), .B(new_new_n493_), .C(new_new_n490_), .D(new_new_n483_), .Y(new_new_n496_));
  NA4        g0474(.A(new_new_n496_), .B(new_new_n480_), .C(new_new_n456_), .D(new_new_n452_), .Y(new_new_n497_));
  NA3        g0475(.A(new_new_n302_), .B(new_new_n177_), .C(new_new_n175_), .Y(new_new_n498_));
  OAI210     g0476(.A0(new_new_n297_), .A1(new_new_n182_), .B0(new_new_n498_), .Y(new_new_n499_));
  AN2        g0477(.A(new_new_n290_), .B(new_new_n234_), .Y(new_new_n500_));
  NA2        g0478(.A(new_new_n500_), .B(new_new_n499_), .Y(new_new_n501_));
  NA2        g0479(.A(new_new_n309_), .B(new_new_n165_), .Y(new_new_n502_));
  OAI210     g0480(.A0(new_new_n502_), .A1(new_new_n232_), .B0(new_new_n303_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n503_), .B(new_new_n318_), .Y(new_new_n504_));
  NA4        g0482(.A(new_new_n433_), .B(new_new_n432_), .C(new_new_n205_), .D(i_2_), .Y(new_new_n505_));
  INV        g0483(.A(new_new_n505_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n378_), .B(new_new_n225_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n354_), .B(new_new_n73_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n367_), .B(new_new_n363_), .Y(new_new_n509_));
  OR2        g0487(.A(new_new_n507_), .B(new_new_n509_), .Y(new_new_n510_));
  NO2        g0488(.A(new_new_n36_), .B(i_8_), .Y(new_new_n511_));
  NAi41      g0489(.An(new_new_n508_), .B(new_new_n471_), .C(new_new_n511_), .D(new_new_n47_), .Y(new_new_n512_));
  AOI210     g0490(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n407_), .Y(new_new_n513_));
  NA3        g0491(.A(new_new_n513_), .B(new_new_n512_), .C(new_new_n510_), .Y(new_new_n514_));
  AOI210     g0492(.A0(new_new_n506_), .A1(new_new_n206_), .B0(new_new_n514_), .Y(new_new_n515_));
  NO2        g0493(.A(i_7_), .B(new_new_n201_), .Y(new_new_n516_));
  OR2        g0494(.A(new_new_n184_), .B(i_4_), .Y(new_new_n517_));
  NO2        g0495(.A(new_new_n517_), .B(new_new_n86_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n518_), .B(new_new_n516_), .Y(new_new_n519_));
  NA4        g0497(.A(new_new_n519_), .B(new_new_n515_), .C(new_new_n504_), .D(new_new_n501_), .Y(new_new_n520_));
  NA2        g0498(.A(new_new_n382_), .B(new_new_n293_), .Y(new_new_n521_));
  OAI210     g0499(.A0(new_new_n380_), .A1(new_new_n170_), .B0(new_new_n521_), .Y(new_new_n522_));
  NO2        g0500(.A(i_12_), .B(new_new_n195_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n523_), .B(new_new_n225_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n471_), .B(new_new_n27_), .Y(new_new_n525_));
  NO2        g0503(.A(new_new_n525_), .B(new_new_n524_), .Y(new_new_n526_));
  NOi31      g0504(.An(new_new_n312_), .B(new_new_n406_), .C(new_new_n38_), .Y(new_new_n527_));
  OAI210     g0505(.A0(new_new_n527_), .A1(new_new_n526_), .B0(new_new_n522_), .Y(new_new_n528_));
  NO2        g0506(.A(i_8_), .B(i_7_), .Y(new_new_n529_));
  OAI210     g0507(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n530_), .B(new_new_n223_), .Y(new_new_n531_));
  AOI220     g0509(.A0(new_new_n319_), .A1(new_new_n40_), .B0(new_new_n235_), .B1(new_new_n208_), .Y(new_new_n532_));
  OAI220     g0510(.A0(new_new_n532_), .A1(new_new_n517_), .B0(new_new_n531_), .B1(new_new_n243_), .Y(new_new_n533_));
  NA2        g0511(.A(new_new_n45_), .B(i_10_), .Y(new_new_n534_));
  NO2        g0512(.A(new_new_n534_), .B(i_6_), .Y(new_new_n535_));
  NA3        g0513(.A(new_new_n535_), .B(new_new_n533_), .C(new_new_n529_), .Y(new_new_n536_));
  AOI220     g0514(.A0(new_new_n417_), .A1(new_new_n319_), .B0(new_new_n247_), .B1(new_new_n244_), .Y(new_new_n537_));
  OAI220     g0515(.A0(new_new_n537_), .A1(new_new_n265_), .B0(new_new_n457_), .B1(new_new_n134_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n538_), .B(new_new_n268_), .Y(new_new_n539_));
  NA3        g0517(.A(new_new_n539_), .B(new_new_n536_), .C(new_new_n528_), .Y(new_new_n540_));
  NA3        g0518(.A(new_new_n219_), .B(new_new_n71_), .C(new_new_n45_), .Y(new_new_n541_));
  NA2        g0519(.A(new_new_n287_), .B(new_new_n84_), .Y(new_new_n542_));
  AOI210     g0520(.A0(new_new_n541_), .A1(new_new_n344_), .B0(new_new_n542_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n434_), .B(new_new_n221_), .Y(new_new_n545_));
  NO2        g0523(.A(new_new_n544_), .B(new_new_n545_), .Y(new_new_n546_));
  NA2        g0524(.A(i_0_), .B(new_new_n49_), .Y(new_new_n547_));
  NO2        g0525(.A(new_new_n546_), .B(new_new_n543_), .Y(new_new_n548_));
  NO4        g0526(.A(new_new_n252_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n549_));
  NO3        g0527(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n550_));
  NO2        g0528(.A(new_new_n233_), .B(new_new_n36_), .Y(new_new_n551_));
  AN2        g0529(.A(new_new_n551_), .B(new_new_n550_), .Y(new_new_n552_));
  OA210      g0530(.A0(new_new_n552_), .A1(new_new_n549_), .B0(new_new_n354_), .Y(new_new_n553_));
  NO2        g0531(.A(new_new_n406_), .B(i_1_), .Y(new_new_n554_));
  NOi31      g0532(.An(new_new_n554_), .B(new_new_n439_), .C(new_new_n73_), .Y(new_new_n555_));
  AN4        g0533(.A(new_new_n555_), .B(new_new_n403_), .C(new_new_n486_), .D(i_2_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n415_), .B(new_new_n178_), .Y(new_new_n557_));
  NO3        g0535(.A(new_new_n557_), .B(new_new_n556_), .C(new_new_n553_), .Y(new_new_n558_));
  NOi21      g0536(.An(i_10_), .B(i_6_), .Y(new_new_n559_));
  NO2        g0537(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n560_));
  AOI220     g0538(.A0(new_new_n287_), .A1(new_new_n560_), .B0(new_new_n278_), .B1(new_new_n559_), .Y(new_new_n561_));
  NO2        g0539(.A(new_new_n561_), .B(new_new_n437_), .Y(new_new_n562_));
  NO2        g0540(.A(new_new_n117_), .B(new_new_n23_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n312_), .B(new_new_n165_), .Y(new_new_n564_));
  AOI220     g0542(.A0(new_new_n564_), .A1(new_new_n423_), .B0(new_new_n185_), .B1(new_new_n183_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n565_), .B(new_new_n562_), .Y(new_new_n566_));
  INV        g0544(.A(new_new_n315_), .Y(new_new_n567_));
  NO2        g0545(.A(i_12_), .B(new_new_n86_), .Y(new_new_n568_));
  NA3        g0546(.A(new_new_n568_), .B(new_new_n278_), .C(new_new_n547_), .Y(new_new_n569_));
  NA3        g0547(.A(new_new_n381_), .B(new_new_n287_), .C(new_new_n219_), .Y(new_new_n570_));
  AOI210     g0548(.A0(new_new_n570_), .A1(new_new_n569_), .B0(new_new_n567_), .Y(new_new_n571_));
  NA2        g0549(.A(new_new_n175_), .B(i_0_), .Y(new_new_n572_));
  NO3        g0550(.A(new_new_n572_), .B(new_new_n337_), .C(new_new_n297_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n573_), .B(new_new_n571_), .Y(new_new_n574_));
  NA4        g0552(.A(new_new_n574_), .B(new_new_n566_), .C(new_new_n558_), .D(new_new_n548_), .Y(new_new_n575_));
  NO4        g0553(.A(new_new_n575_), .B(new_new_n540_), .C(new_new_n520_), .D(new_new_n497_), .Y(new_new_n576_));
  NA4        g0554(.A(new_new_n576_), .B(new_new_n431_), .C(new_new_n353_), .D(new_new_n308_), .Y(men7));
  NO2        g0555(.A(new_new_n95_), .B(new_new_n55_), .Y(new_new_n578_));
  NO2        g0556(.A(new_new_n110_), .B(new_new_n92_), .Y(new_new_n579_));
  NA2        g0557(.A(new_new_n379_), .B(new_new_n579_), .Y(new_new_n580_));
  NA2        g0558(.A(new_new_n471_), .B(new_new_n84_), .Y(new_new_n581_));
  NA2        g0559(.A(i_11_), .B(new_new_n195_), .Y(new_new_n582_));
  NA2        g0560(.A(new_new_n145_), .B(new_new_n582_), .Y(new_new_n583_));
  OAI210     g0561(.A0(new_new_n583_), .A1(new_new_n581_), .B0(new_new_n580_), .Y(new_new_n584_));
  NA3        g0562(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n585_));
  NO2        g0563(.A(new_new_n237_), .B(i_4_), .Y(new_new_n586_));
  NA2        g0564(.A(new_new_n586_), .B(i_8_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n107_), .B(new_new_n585_), .Y(new_new_n588_));
  NA2        g0566(.A(i_2_), .B(new_new_n86_), .Y(new_new_n589_));
  OAI210     g0567(.A0(new_new_n89_), .A1(new_new_n205_), .B0(new_new_n206_), .Y(new_new_n590_));
  NO2        g0568(.A(i_7_), .B(new_new_n37_), .Y(new_new_n591_));
  NA2        g0569(.A(i_4_), .B(i_8_), .Y(new_new_n592_));
  AOI210     g0570(.A0(new_new_n592_), .A1(new_new_n302_), .B0(new_new_n591_), .Y(new_new_n593_));
  OAI220     g0571(.A0(new_new_n593_), .A1(new_new_n589_), .B0(new_new_n590_), .B1(i_13_), .Y(new_new_n594_));
  NO4        g0572(.A(new_new_n594_), .B(new_new_n588_), .C(new_new_n584_), .D(new_new_n578_), .Y(new_new_n595_));
  AOI210     g0573(.A0(new_new_n129_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n596_));
  AOI210     g0574(.A0(new_new_n596_), .A1(new_new_n237_), .B0(new_new_n162_), .Y(new_new_n597_));
  OR2        g0575(.A(i_6_), .B(i_10_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n598_), .B(new_new_n23_), .Y(new_new_n599_));
  OR3        g0577(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n600_));
  NO3        g0578(.A(new_new_n600_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n601_));
  INV        g0579(.A(new_new_n202_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n601_), .B(new_new_n599_), .Y(new_new_n603_));
  OA220      g0581(.A0(new_new_n603_), .A1(new_new_n567_), .B0(new_new_n597_), .B1(new_new_n270_), .Y(new_new_n604_));
  AOI210     g0582(.A0(new_new_n604_), .A1(new_new_n595_), .B0(new_new_n63_), .Y(new_new_n605_));
  NOi21      g0583(.An(i_11_), .B(i_7_), .Y(new_new_n606_));
  AO210      g0584(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n607_));
  NO2        g0585(.A(new_new_n607_), .B(new_new_n606_), .Y(new_new_n608_));
  NA2        g0586(.A(new_new_n608_), .B(new_new_n208_), .Y(new_new_n609_));
  NA3        g0587(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n610_));
  NAi31      g0588(.An(new_new_n610_), .B(new_new_n217_), .C(i_11_), .Y(new_new_n611_));
  AOI210     g0589(.A0(new_new_n611_), .A1(new_new_n609_), .B0(new_new_n63_), .Y(new_new_n612_));
  NA2        g0590(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n613_));
  OR2        g0591(.A(new_new_n613_), .B(new_new_n41_), .Y(new_new_n614_));
  NO3        g0592(.A(new_new_n260_), .B(new_new_n210_), .C(new_new_n582_), .Y(new_new_n615_));
  OAI210     g0593(.A0(new_new_n615_), .A1(new_new_n226_), .B0(new_new_n63_), .Y(new_new_n616_));
  NO2        g0594(.A(new_new_n63_), .B(i_9_), .Y(new_new_n617_));
  NO2        g0595(.A(i_1_), .B(i_12_), .Y(new_new_n618_));
  NA2        g0596(.A(new_new_n616_), .B(new_new_n614_), .Y(new_new_n619_));
  OAI210     g0597(.A0(new_new_n619_), .A1(new_new_n612_), .B0(i_6_), .Y(new_new_n620_));
  NO2        g0598(.A(new_new_n610_), .B(new_new_n110_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n621_), .B(new_new_n568_), .Y(new_new_n622_));
  NO2        g0600(.A(new_new_n237_), .B(new_new_n86_), .Y(new_new_n623_));
  NO2        g0601(.A(new_new_n623_), .B(i_11_), .Y(new_new_n624_));
  NA2        g0602(.A(new_new_n622_), .B(new_new_n440_), .Y(new_new_n625_));
  NO4        g0603(.A(new_new_n217_), .B(new_new_n129_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n626_));
  NA2        g0604(.A(new_new_n626_), .B(new_new_n617_), .Y(new_new_n627_));
  NA2        g0605(.A(new_new_n237_), .B(i_6_), .Y(new_new_n628_));
  NO3        g0606(.A(new_new_n598_), .B(new_new_n233_), .C(new_new_n23_), .Y(new_new_n629_));
  AOI210     g0607(.A0(i_1_), .A1(new_new_n261_), .B0(new_new_n629_), .Y(new_new_n630_));
  OAI210     g0608(.A0(new_new_n630_), .A1(new_new_n45_), .B0(new_new_n627_), .Y(new_new_n631_));
  INV        g0609(.A(i_2_), .Y(new_new_n632_));
  NA2        g0610(.A(new_new_n139_), .B(i_9_), .Y(new_new_n633_));
  NA3        g0611(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n634_));
  NO2        g0612(.A(new_new_n47_), .B(i_1_), .Y(new_new_n635_));
  NA3        g0613(.A(new_new_n635_), .B(new_new_n269_), .C(new_new_n45_), .Y(new_new_n636_));
  OAI220     g0614(.A0(new_new_n636_), .A1(new_new_n634_), .B0(new_new_n633_), .B1(new_new_n632_), .Y(new_new_n637_));
  NA3        g0615(.A(new_new_n617_), .B(new_new_n315_), .C(i_6_), .Y(new_new_n638_));
  NO2        g0616(.A(new_new_n638_), .B(new_new_n23_), .Y(new_new_n639_));
  AOI210     g0617(.A0(new_new_n462_), .A1(new_new_n409_), .B0(new_new_n242_), .Y(new_new_n640_));
  NO2        g0618(.A(new_new_n640_), .B(new_new_n589_), .Y(new_new_n641_));
  NA2        g0619(.A(new_new_n635_), .B(new_new_n269_), .Y(new_new_n642_));
  NO2        g0620(.A(i_11_), .B(new_new_n37_), .Y(new_new_n643_));
  NA2        g0621(.A(new_new_n643_), .B(new_new_n24_), .Y(new_new_n644_));
  NO2        g0622(.A(new_new_n644_), .B(new_new_n642_), .Y(new_new_n645_));
  OR4        g0623(.A(new_new_n645_), .B(new_new_n641_), .C(new_new_n639_), .D(new_new_n637_), .Y(new_new_n646_));
  NO3        g0624(.A(new_new_n646_), .B(new_new_n631_), .C(new_new_n625_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n237_), .B(new_new_n103_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n648_), .B(new_new_n606_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n649_), .B(i_1_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n650_), .B(new_new_n600_), .Y(new_new_n651_));
  NO2        g0629(.A(new_new_n405_), .B(new_new_n86_), .Y(new_new_n652_));
  NA2        g0630(.A(new_new_n651_), .B(new_new_n47_), .Y(new_new_n653_));
  NA2        g0631(.A(i_3_), .B(new_new_n195_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n654_), .B(new_new_n117_), .Y(new_new_n655_));
  AN2        g0633(.A(new_new_n655_), .B(new_new_n535_), .Y(new_new_n656_));
  NO2        g0634(.A(new_new_n233_), .B(new_new_n45_), .Y(new_new_n657_));
  NO3        g0635(.A(new_new_n657_), .B(new_new_n305_), .C(new_new_n238_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n119_), .B(new_new_n37_), .Y(new_new_n659_));
  NO2        g0637(.A(new_new_n659_), .B(i_6_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n86_), .B(i_9_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n661_), .B(new_new_n63_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n662_), .B(new_new_n618_), .Y(new_new_n663_));
  NO4        g0641(.A(new_new_n663_), .B(new_new_n660_), .C(new_new_n658_), .D(i_4_), .Y(new_new_n664_));
  NA2        g0642(.A(i_1_), .B(i_3_), .Y(new_new_n665_));
  NO2        g0643(.A(new_new_n441_), .B(new_new_n95_), .Y(new_new_n666_));
  AOI210     g0644(.A0(new_new_n657_), .A1(new_new_n559_), .B0(new_new_n666_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n667_), .B(new_new_n665_), .Y(new_new_n668_));
  NO3        g0646(.A(new_new_n668_), .B(new_new_n664_), .C(new_new_n656_), .Y(new_new_n669_));
  NA4        g0647(.A(new_new_n669_), .B(new_new_n653_), .C(new_new_n647_), .D(new_new_n620_), .Y(new_new_n670_));
  NO3        g0648(.A(new_new_n464_), .B(i_3_), .C(i_7_), .Y(new_new_n671_));
  NOi21      g0649(.An(new_new_n671_), .B(i_10_), .Y(new_new_n672_));
  OA210      g0650(.A0(new_new_n672_), .A1(new_new_n245_), .B0(new_new_n86_), .Y(new_new_n673_));
  NO3        g0651(.A(new_new_n465_), .B(new_new_n592_), .C(new_new_n86_), .Y(new_new_n674_));
  NA2        g0652(.A(new_new_n674_), .B(new_new_n25_), .Y(new_new_n675_));
  INV        g0653(.A(new_new_n675_), .Y(new_new_n676_));
  OAI210     g0654(.A0(new_new_n676_), .A1(new_new_n673_), .B0(i_1_), .Y(new_new_n677_));
  AOI210     g0655(.A0(new_new_n269_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n365_), .B(i_2_), .Y(new_new_n679_));
  NA2        g0657(.A(new_new_n679_), .B(new_new_n678_), .Y(new_new_n680_));
  OAI210     g0658(.A0(new_new_n638_), .A1(new_new_n435_), .B0(new_new_n680_), .Y(new_new_n681_));
  INV        g0659(.A(new_new_n681_), .Y(new_new_n682_));
  AOI210     g0660(.A0(new_new_n682_), .A1(new_new_n677_), .B0(i_13_), .Y(new_new_n683_));
  OR2        g0661(.A(i_11_), .B(i_7_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n55_), .B(i_12_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n465_), .B(new_new_n24_), .Y(new_new_n686_));
  AOI220     g0664(.A0(new_new_n686_), .A1(new_new_n652_), .B0(new_new_n245_), .B1(new_new_n132_), .Y(new_new_n687_));
  OAI220     g0665(.A0(new_new_n687_), .A1(new_new_n41_), .B0(new_new_n1042_), .B1(new_new_n95_), .Y(new_new_n688_));
  INV        g0666(.A(new_new_n688_), .Y(new_new_n689_));
  NA2        g0667(.A(new_new_n381_), .B(new_new_n635_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n690_), .B(new_new_n243_), .Y(new_new_n691_));
  AOI210     g0669(.A0(new_new_n435_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n692_));
  NOi31      g0670(.An(new_new_n692_), .B(new_new_n581_), .C(new_new_n45_), .Y(new_new_n693_));
  NA2        g0671(.A(new_new_n128_), .B(i_13_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n634_), .B(new_new_n117_), .Y(new_new_n695_));
  INV        g0673(.A(new_new_n695_), .Y(new_new_n696_));
  OAI220     g0674(.A0(new_new_n696_), .A1(new_new_n71_), .B0(new_new_n694_), .B1(new_new_n678_), .Y(new_new_n697_));
  NO3        g0675(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n103_), .Y(new_new_n698_));
  NA2        g0676(.A(new_new_n26_), .B(new_new_n195_), .Y(new_new_n699_));
  NA2        g0677(.A(new_new_n699_), .B(i_7_), .Y(new_new_n700_));
  NO3        g0678(.A(new_new_n465_), .B(new_new_n237_), .C(new_new_n86_), .Y(new_new_n701_));
  AOI210     g0679(.A0(new_new_n701_), .A1(new_new_n700_), .B0(new_new_n698_), .Y(new_new_n702_));
  AOI220     g0680(.A0(new_new_n381_), .A1(new_new_n635_), .B0(new_new_n94_), .B1(new_new_n104_), .Y(new_new_n703_));
  OAI220     g0681(.A0(new_new_n703_), .A1(new_new_n587_), .B0(new_new_n702_), .B1(new_new_n602_), .Y(new_new_n704_));
  NO4        g0682(.A(new_new_n704_), .B(new_new_n697_), .C(new_new_n693_), .D(new_new_n691_), .Y(new_new_n705_));
  OR2        g0683(.A(i_11_), .B(i_6_), .Y(new_new_n706_));
  NA3        g0684(.A(new_new_n586_), .B(new_new_n699_), .C(i_7_), .Y(new_new_n707_));
  AOI210     g0685(.A0(new_new_n707_), .A1(new_new_n696_), .B0(new_new_n706_), .Y(new_new_n708_));
  NA3        g0686(.A(new_new_n399_), .B(new_new_n591_), .C(new_new_n99_), .Y(new_new_n709_));
  NA2        g0687(.A(new_new_n624_), .B(i_13_), .Y(new_new_n710_));
  NA2        g0688(.A(new_new_n104_), .B(new_new_n699_), .Y(new_new_n711_));
  NAi21      g0689(.An(i_11_), .B(i_12_), .Y(new_new_n712_));
  NOi41      g0690(.An(new_new_n113_), .B(new_new_n712_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n713_));
  NO3        g0691(.A(new_new_n465_), .B(new_new_n568_), .C(new_new_n592_), .Y(new_new_n714_));
  AOI220     g0692(.A0(new_new_n714_), .A1(new_new_n309_), .B0(new_new_n713_), .B1(new_new_n711_), .Y(new_new_n715_));
  NA3        g0693(.A(new_new_n715_), .B(new_new_n710_), .C(new_new_n709_), .Y(new_new_n716_));
  OAI210     g0694(.A0(new_new_n716_), .A1(new_new_n708_), .B0(new_new_n63_), .Y(new_new_n717_));
  NO2        g0695(.A(i_2_), .B(i_12_), .Y(new_new_n718_));
  NA2        g0696(.A(new_new_n364_), .B(new_new_n718_), .Y(new_new_n719_));
  NA2        g0697(.A(i_8_), .B(new_new_n25_), .Y(new_new_n720_));
  NO3        g0698(.A(new_new_n720_), .B(new_new_n379_), .C(new_new_n586_), .Y(new_new_n721_));
  OAI210     g0699(.A0(new_new_n721_), .A1(new_new_n366_), .B0(new_new_n364_), .Y(new_new_n722_));
  NO2        g0700(.A(new_new_n129_), .B(i_2_), .Y(new_new_n723_));
  NA2        g0701(.A(new_new_n723_), .B(new_new_n618_), .Y(new_new_n724_));
  NA3        g0702(.A(new_new_n724_), .B(new_new_n722_), .C(new_new_n719_), .Y(new_new_n725_));
  NA3        g0703(.A(new_new_n725_), .B(new_new_n46_), .C(new_new_n225_), .Y(new_new_n726_));
  NA4        g0704(.A(new_new_n726_), .B(new_new_n717_), .C(new_new_n705_), .D(new_new_n689_), .Y(new_new_n727_));
  OR4        g0705(.A(new_new_n727_), .B(new_new_n683_), .C(new_new_n670_), .D(new_new_n605_), .Y(men5));
  NA2        g0706(.A(new_new_n649_), .B(new_new_n272_), .Y(new_new_n729_));
  AN2        g0707(.A(new_new_n24_), .B(i_10_), .Y(new_new_n730_));
  NA3        g0708(.A(new_new_n730_), .B(new_new_n718_), .C(new_new_n110_), .Y(new_new_n731_));
  NO2        g0709(.A(new_new_n587_), .B(i_11_), .Y(new_new_n732_));
  NA2        g0710(.A(new_new_n89_), .B(new_new_n732_), .Y(new_new_n733_));
  NA3        g0711(.A(new_new_n733_), .B(new_new_n731_), .C(new_new_n729_), .Y(new_new_n734_));
  NO3        g0712(.A(i_11_), .B(new_new_n237_), .C(i_13_), .Y(new_new_n735_));
  NO2        g0713(.A(new_new_n125_), .B(new_new_n23_), .Y(new_new_n736_));
  NA2        g0714(.A(i_12_), .B(i_8_), .Y(new_new_n737_));
  OAI210     g0715(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n737_), .Y(new_new_n738_));
  INV        g0716(.A(new_new_n434_), .Y(new_new_n739_));
  AOI220     g0717(.A0(new_new_n315_), .A1(new_new_n563_), .B0(new_new_n738_), .B1(new_new_n736_), .Y(new_new_n740_));
  INV        g0718(.A(new_new_n740_), .Y(new_new_n741_));
  NO2        g0719(.A(new_new_n741_), .B(new_new_n734_), .Y(new_new_n742_));
  INV        g0720(.A(new_new_n173_), .Y(new_new_n743_));
  INV        g0721(.A(new_new_n245_), .Y(new_new_n744_));
  OAI210     g0722(.A0(new_new_n679_), .A1(new_new_n436_), .B0(new_new_n113_), .Y(new_new_n745_));
  AOI210     g0723(.A0(new_new_n745_), .A1(new_new_n744_), .B0(new_new_n743_), .Y(new_new_n746_));
  NO2        g0724(.A(new_new_n441_), .B(new_new_n26_), .Y(new_new_n747_));
  NO2        g0725(.A(new_new_n747_), .B(new_new_n409_), .Y(new_new_n748_));
  NA2        g0726(.A(new_new_n748_), .B(i_2_), .Y(new_new_n749_));
  INV        g0727(.A(new_new_n749_), .Y(new_new_n750_));
  AOI210     g0728(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n406_), .Y(new_new_n751_));
  AOI210     g0729(.A0(new_new_n751_), .A1(new_new_n750_), .B0(new_new_n746_), .Y(new_new_n752_));
  NO2        g0730(.A(new_new_n192_), .B(new_new_n126_), .Y(new_new_n753_));
  OAI210     g0731(.A0(new_new_n753_), .A1(new_new_n736_), .B0(i_2_), .Y(new_new_n754_));
  INV        g0732(.A(new_new_n174_), .Y(new_new_n755_));
  NO3        g0733(.A(new_new_n607_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n756_));
  AOI210     g0734(.A0(new_new_n755_), .A1(new_new_n89_), .B0(new_new_n756_), .Y(new_new_n757_));
  AOI210     g0735(.A0(new_new_n757_), .A1(new_new_n754_), .B0(new_new_n195_), .Y(new_new_n758_));
  OA210      g0736(.A0(new_new_n608_), .A1(new_new_n127_), .B0(i_13_), .Y(new_new_n759_));
  NA2        g0737(.A(new_new_n202_), .B(new_new_n205_), .Y(new_new_n760_));
  NA2        g0738(.A(new_new_n152_), .B(new_new_n582_), .Y(new_new_n761_));
  AOI210     g0739(.A0(new_new_n761_), .A1(new_new_n760_), .B0(new_new_n369_), .Y(new_new_n762_));
  AOI210     g0740(.A0(new_new_n210_), .A1(new_new_n149_), .B0(new_new_n511_), .Y(new_new_n763_));
  NA2        g0741(.A(new_new_n763_), .B(new_new_n409_), .Y(new_new_n764_));
  NO2        g0742(.A(new_new_n104_), .B(new_new_n45_), .Y(new_new_n765_));
  INV        g0743(.A(new_new_n298_), .Y(new_new_n766_));
  NA4        g0744(.A(new_new_n766_), .B(new_new_n302_), .C(new_new_n125_), .D(new_new_n43_), .Y(new_new_n767_));
  OAI210     g0745(.A0(new_new_n767_), .A1(new_new_n765_), .B0(new_new_n764_), .Y(new_new_n768_));
  NO4        g0746(.A(new_new_n768_), .B(new_new_n762_), .C(new_new_n759_), .D(new_new_n758_), .Y(new_new_n769_));
  NA2        g0747(.A(new_new_n563_), .B(new_new_n28_), .Y(new_new_n770_));
  NA2        g0748(.A(new_new_n735_), .B(new_new_n279_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n771_), .B(new_new_n770_), .Y(new_new_n772_));
  NO2        g0750(.A(new_new_n62_), .B(i_12_), .Y(new_new_n773_));
  NO2        g0751(.A(new_new_n773_), .B(new_new_n127_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n774_), .B(new_new_n582_), .Y(new_new_n775_));
  AOI220     g0753(.A0(new_new_n775_), .A1(new_new_n36_), .B0(new_new_n772_), .B1(new_new_n47_), .Y(new_new_n776_));
  NA4        g0754(.A(new_new_n776_), .B(new_new_n769_), .C(new_new_n752_), .D(new_new_n742_), .Y(men6));
  NO3        g0755(.A(new_new_n256_), .B(new_new_n304_), .C(i_1_), .Y(new_new_n778_));
  NO2        g0756(.A(new_new_n187_), .B(new_new_n140_), .Y(new_new_n779_));
  OAI210     g0757(.A0(new_new_n779_), .A1(new_new_n778_), .B0(new_new_n723_), .Y(new_new_n780_));
  NA4        g0758(.A(new_new_n383_), .B(new_new_n470_), .C(new_new_n71_), .D(new_new_n103_), .Y(new_new_n781_));
  INV        g0759(.A(new_new_n781_), .Y(new_new_n782_));
  NO2        g0760(.A(new_new_n220_), .B(new_new_n475_), .Y(new_new_n783_));
  NO2        g0761(.A(i_11_), .B(i_9_), .Y(new_new_n784_));
  NO2        g0762(.A(new_new_n782_), .B(new_new_n324_), .Y(new_new_n785_));
  AO210      g0763(.A0(new_new_n785_), .A1(new_new_n780_), .B0(i_12_), .Y(new_new_n786_));
  NA2        g0764(.A(new_new_n370_), .B(new_new_n331_), .Y(new_new_n787_));
  NA2        g0765(.A(new_new_n568_), .B(new_new_n63_), .Y(new_new_n788_));
  NA2        g0766(.A(new_new_n672_), .B(new_new_n71_), .Y(new_new_n789_));
  BUFFER     g0767(.A(new_new_n613_), .Y(new_new_n790_));
  NA4        g0768(.A(new_new_n790_), .B(new_new_n789_), .C(new_new_n788_), .D(new_new_n787_), .Y(new_new_n791_));
  INV        g0769(.A(new_new_n199_), .Y(new_new_n792_));
  AOI220     g0770(.A0(new_new_n792_), .A1(new_new_n784_), .B0(new_new_n791_), .B1(new_new_n73_), .Y(new_new_n793_));
  INV        g0771(.A(new_new_n323_), .Y(new_new_n794_));
  NA2        g0772(.A(new_new_n75_), .B(new_new_n132_), .Y(new_new_n795_));
  INV        g0773(.A(new_new_n125_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n796_), .B(new_new_n47_), .Y(new_new_n797_));
  AOI210     g0775(.A0(new_new_n797_), .A1(new_new_n795_), .B0(new_new_n794_), .Y(new_new_n798_));
  NO2        g0776(.A(new_new_n252_), .B(i_9_), .Y(new_new_n799_));
  NA2        g0777(.A(new_new_n799_), .B(new_new_n773_), .Y(new_new_n800_));
  AOI210     g0778(.A0(new_new_n800_), .A1(new_new_n509_), .B0(new_new_n187_), .Y(new_new_n801_));
  NO2        g0779(.A(new_new_n32_), .B(i_11_), .Y(new_new_n802_));
  NA3        g0780(.A(new_new_n802_), .B(new_new_n460_), .C(new_new_n383_), .Y(new_new_n803_));
  NAi32      g0781(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n804_));
  NO2        g0782(.A(new_new_n706_), .B(new_new_n804_), .Y(new_new_n805_));
  OAI210     g0783(.A0(new_new_n671_), .A1(new_new_n551_), .B0(new_new_n550_), .Y(new_new_n806_));
  NAi31      g0784(.An(new_new_n805_), .B(new_new_n806_), .C(new_new_n803_), .Y(new_new_n807_));
  OR3        g0785(.A(new_new_n807_), .B(new_new_n801_), .C(new_new_n798_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n684_), .B(i_2_), .Y(new_new_n809_));
  NA2        g0787(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n810_));
  NO2        g0788(.A(new_new_n810_), .B(new_new_n398_), .Y(new_new_n811_));
  NA2        g0789(.A(new_new_n811_), .B(new_new_n809_), .Y(new_new_n812_));
  AO220      g0790(.A0(new_new_n358_), .A1(new_new_n348_), .B0(new_new_n385_), .B1(new_new_n582_), .Y(new_new_n813_));
  NA3        g0791(.A(new_new_n813_), .B(new_new_n257_), .C(i_7_), .Y(new_new_n814_));
  BUFFER     g0792(.A(new_new_n608_), .Y(new_new_n815_));
  NA3        g0793(.A(new_new_n815_), .B(new_new_n148_), .C(new_new_n69_), .Y(new_new_n816_));
  AO210      g0794(.A0(new_new_n482_), .A1(new_new_n739_), .B0(new_new_n36_), .Y(new_new_n817_));
  NA4        g0795(.A(new_new_n817_), .B(new_new_n816_), .C(new_new_n814_), .D(new_new_n812_), .Y(new_new_n818_));
  OAI210     g0796(.A0(new_new_n623_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n819_));
  AOI220     g0797(.A0(new_new_n819_), .A1(new_new_n550_), .B0(new_new_n783_), .B1(new_new_n700_), .Y(new_new_n820_));
  NA3        g0798(.A(new_new_n369_), .B(new_new_n239_), .C(new_new_n148_), .Y(new_new_n821_));
  NA2        g0799(.A(new_new_n385_), .B(new_new_n70_), .Y(new_new_n822_));
  NA4        g0800(.A(new_new_n822_), .B(new_new_n821_), .C(new_new_n820_), .D(new_new_n590_), .Y(new_new_n823_));
  AO210      g0801(.A0(new_new_n511_), .A1(new_new_n47_), .B0(new_new_n88_), .Y(new_new_n824_));
  NA3        g0802(.A(new_new_n824_), .B(new_new_n471_), .C(new_new_n219_), .Y(new_new_n825_));
  AOI210     g0803(.A0(new_new_n436_), .A1(new_new_n434_), .B0(new_new_n549_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n598_), .B(new_new_n104_), .Y(new_new_n827_));
  OAI210     g0805(.A0(new_new_n827_), .A1(new_new_n114_), .B0(new_new_n396_), .Y(new_new_n828_));
  NA3        g0806(.A(new_new_n828_), .B(new_new_n826_), .C(new_new_n825_), .Y(new_new_n829_));
  NO4        g0807(.A(new_new_n829_), .B(new_new_n823_), .C(new_new_n818_), .D(new_new_n808_), .Y(new_new_n830_));
  NA4        g0808(.A(new_new_n830_), .B(new_new_n793_), .C(new_new_n786_), .D(new_new_n375_), .Y(men3));
  NA2        g0809(.A(i_6_), .B(i_7_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n832_), .B(i_0_), .Y(new_new_n833_));
  NO2        g0811(.A(i_11_), .B(new_new_n237_), .Y(new_new_n834_));
  OAI210     g0812(.A0(new_new_n833_), .A1(new_new_n291_), .B0(new_new_n834_), .Y(new_new_n835_));
  NO2        g0813(.A(new_new_n835_), .B(new_new_n195_), .Y(new_new_n836_));
  NO3        g0814(.A(new_new_n437_), .B(new_new_n92_), .C(new_new_n45_), .Y(new_new_n837_));
  OA210      g0815(.A0(new_new_n837_), .A1(new_new_n836_), .B0(new_new_n175_), .Y(new_new_n838_));
  NA2        g0816(.A(new_new_n821_), .B(new_new_n368_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n839_), .B(new_new_n40_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n399_), .B(new_new_n46_), .Y(new_new_n841_));
  NO2        g0819(.A(new_new_n840_), .B(new_new_n49_), .Y(new_new_n842_));
  NO4        g0820(.A(new_new_n372_), .B(new_new_n378_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n187_), .B(new_new_n559_), .Y(new_new_n844_));
  NOi21      g0822(.An(new_new_n844_), .B(new_new_n843_), .Y(new_new_n845_));
  NA2        g0823(.A(new_new_n692_), .B(new_new_n661_), .Y(new_new_n846_));
  NA2        g0824(.A(new_new_n329_), .B(new_new_n425_), .Y(new_new_n847_));
  OAI220     g0825(.A0(new_new_n847_), .A1(new_new_n846_), .B0(new_new_n845_), .B1(new_new_n63_), .Y(new_new_n848_));
  NOi21      g0826(.An(i_5_), .B(i_9_), .Y(new_new_n849_));
  NA2        g0827(.A(new_new_n849_), .B(new_new_n433_), .Y(new_new_n850_));
  BUFFER     g0828(.A(new_new_n269_), .Y(new_new_n851_));
  AOI210     g0829(.A0(new_new_n851_), .A1(new_new_n462_), .B0(new_new_n674_), .Y(new_new_n852_));
  NO3        g0830(.A(new_new_n402_), .B(new_new_n269_), .C(new_new_n73_), .Y(new_new_n853_));
  NO2        g0831(.A(new_new_n176_), .B(new_new_n149_), .Y(new_new_n854_));
  AOI210     g0832(.A0(new_new_n854_), .A1(new_new_n244_), .B0(new_new_n853_), .Y(new_new_n855_));
  OAI220     g0833(.A0(new_new_n855_), .A1(new_new_n182_), .B0(new_new_n852_), .B1(new_new_n850_), .Y(new_new_n856_));
  NO4        g0834(.A(new_new_n856_), .B(new_new_n848_), .C(new_new_n842_), .D(new_new_n838_), .Y(new_new_n857_));
  NA2        g0835(.A(new_new_n187_), .B(new_new_n24_), .Y(new_new_n858_));
  NO2        g0836(.A(new_new_n659_), .B(new_new_n579_), .Y(new_new_n859_));
  NO2        g0837(.A(new_new_n859_), .B(new_new_n858_), .Y(new_new_n860_));
  NA2        g0838(.A(new_new_n309_), .B(new_new_n130_), .Y(new_new_n861_));
  NO2        g0839(.A(new_new_n861_), .B(new_new_n388_), .Y(new_new_n862_));
  NO2        g0840(.A(new_new_n862_), .B(new_new_n860_), .Y(new_new_n863_));
  NO2        g0841(.A(new_new_n383_), .B(new_new_n292_), .Y(new_new_n864_));
  NA2        g0842(.A(new_new_n864_), .B(new_new_n695_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n560_), .B(i_0_), .Y(new_new_n866_));
  NO3        g0844(.A(new_new_n866_), .B(new_new_n380_), .C(new_new_n89_), .Y(new_new_n867_));
  INV        g0845(.A(new_new_n867_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n735_), .B(new_new_n324_), .Y(new_new_n869_));
  AOI210     g0847(.A0(new_new_n471_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n870_));
  OAI220     g0848(.A0(new_new_n870_), .A1(new_new_n869_), .B0(new_new_n644_), .B1(new_new_n531_), .Y(new_new_n871_));
  NO2        g0849(.A(new_new_n254_), .B(new_new_n154_), .Y(new_new_n872_));
  NA2        g0850(.A(i_0_), .B(i_10_), .Y(new_new_n873_));
  AN2        g0851(.A(new_new_n872_), .B(i_6_), .Y(new_new_n874_));
  AOI220     g0852(.A0(new_new_n329_), .A1(new_new_n100_), .B0(new_new_n187_), .B1(new_new_n84_), .Y(new_new_n875_));
  NA2        g0853(.A(new_new_n554_), .B(i_4_), .Y(new_new_n876_));
  NA2        g0854(.A(new_new_n190_), .B(new_new_n205_), .Y(new_new_n877_));
  OAI220     g0855(.A0(new_new_n877_), .A1(new_new_n869_), .B0(new_new_n876_), .B1(new_new_n875_), .Y(new_new_n878_));
  NO3        g0856(.A(new_new_n878_), .B(new_new_n874_), .C(new_new_n871_), .Y(new_new_n879_));
  NA4        g0857(.A(new_new_n879_), .B(new_new_n868_), .C(new_new_n865_), .D(new_new_n863_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n881_));
  NA2        g0859(.A(i_11_), .B(i_9_), .Y(new_new_n882_));
  NO3        g0860(.A(i_12_), .B(new_new_n882_), .C(new_new_n589_), .Y(new_new_n883_));
  AN2        g0861(.A(new_new_n883_), .B(new_new_n881_), .Y(new_new_n884_));
  NO2        g0862(.A(new_new_n49_), .B(i_7_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n384_), .B(new_new_n180_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n886_), .B(new_new_n161_), .Y(new_new_n887_));
  NO2        g0865(.A(new_new_n176_), .B(i_0_), .Y(new_new_n888_));
  AOI210     g0866(.A0(new_new_n367_), .A1(new_new_n42_), .B0(new_new_n395_), .Y(new_new_n889_));
  NO2        g0867(.A(new_new_n889_), .B(new_new_n850_), .Y(new_new_n890_));
  NO3        g0868(.A(new_new_n890_), .B(new_new_n887_), .C(new_new_n884_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n643_), .B(new_new_n122_), .Y(new_new_n892_));
  NO2        g0870(.A(i_6_), .B(new_new_n892_), .Y(new_new_n893_));
  AOI210     g0871(.A0(new_new_n435_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n894_));
  NA2        g0872(.A(new_new_n173_), .B(new_new_n105_), .Y(new_new_n895_));
  NOi32      g0873(.An(new_new_n894_), .Bn(new_new_n190_), .C(new_new_n895_), .Y(new_new_n896_));
  NA2        g0874(.A(new_new_n591_), .B(new_new_n324_), .Y(new_new_n897_));
  NO2        g0875(.A(new_new_n897_), .B(new_new_n841_), .Y(new_new_n898_));
  NO3        g0876(.A(new_new_n898_), .B(new_new_n896_), .C(new_new_n893_), .Y(new_new_n899_));
  NOi21      g0877(.An(i_7_), .B(i_5_), .Y(new_new_n900_));
  NOi31      g0878(.An(new_new_n900_), .B(i_0_), .C(new_new_n712_), .Y(new_new_n901_));
  NA3        g0879(.A(new_new_n901_), .B(new_new_n379_), .C(i_6_), .Y(new_new_n902_));
  BUFFER     g0880(.A(new_new_n902_), .Y(new_new_n903_));
  NO3        g0881(.A(new_new_n391_), .B(new_new_n361_), .C(new_new_n357_), .Y(new_new_n904_));
  NO2        g0882(.A(new_new_n263_), .B(new_new_n316_), .Y(new_new_n905_));
  NO2        g0883(.A(new_new_n712_), .B(new_new_n259_), .Y(new_new_n906_));
  AOI210     g0884(.A0(new_new_n906_), .A1(new_new_n905_), .B0(new_new_n904_), .Y(new_new_n907_));
  NA4        g0885(.A(new_new_n907_), .B(new_new_n903_), .C(new_new_n899_), .D(new_new_n891_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n858_), .B(new_new_n240_), .Y(new_new_n909_));
  AN2        g0887(.A(new_new_n328_), .B(new_new_n324_), .Y(new_new_n910_));
  AN2        g0888(.A(new_new_n910_), .B(new_new_n854_), .Y(new_new_n911_));
  OAI210     g0889(.A0(new_new_n911_), .A1(new_new_n909_), .B0(i_10_), .Y(new_new_n912_));
  OA210      g0890(.A0(new_new_n460_), .A1(new_new_n223_), .B0(new_new_n459_), .Y(new_new_n913_));
  NO2        g0891(.A(new_new_n257_), .B(new_new_n47_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n914_), .B(new_new_n189_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n915_), .B(new_new_n460_), .Y(new_new_n916_));
  NA3        g0894(.A(new_new_n810_), .B(new_new_n377_), .C(new_new_n623_), .Y(new_new_n917_));
  NA2        g0895(.A(new_new_n95_), .B(new_new_n45_), .Y(new_new_n918_));
  NO2        g0896(.A(new_new_n75_), .B(new_new_n737_), .Y(new_new_n919_));
  AOI220     g0897(.A0(new_new_n919_), .A1(new_new_n918_), .B0(new_new_n175_), .B1(new_new_n579_), .Y(new_new_n920_));
  AOI210     g0898(.A0(new_new_n920_), .A1(new_new_n917_), .B0(new_new_n48_), .Y(new_new_n921_));
  NO3        g0899(.A(i_5_), .B(new_new_n356_), .C(new_new_n24_), .Y(new_new_n922_));
  INV        g0900(.A(new_new_n922_), .Y(new_new_n923_));
  NAi21      g0901(.An(i_9_), .B(i_5_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n924_), .B(new_new_n391_), .Y(new_new_n925_));
  NO2        g0903(.A(new_new_n585_), .B(new_new_n107_), .Y(new_new_n926_));
  AOI220     g0904(.A0(new_new_n926_), .A1(i_0_), .B0(new_new_n925_), .B1(new_new_n608_), .Y(new_new_n927_));
  OAI220     g0905(.A0(new_new_n927_), .A1(new_new_n86_), .B0(new_new_n923_), .B1(new_new_n174_), .Y(new_new_n928_));
  NO3        g0906(.A(new_new_n928_), .B(new_new_n921_), .C(new_new_n514_), .Y(new_new_n929_));
  NA3        g0907(.A(new_new_n929_), .B(new_new_n916_), .C(new_new_n912_), .Y(new_new_n930_));
  NO3        g0908(.A(new_new_n930_), .B(new_new_n908_), .C(new_new_n880_), .Y(new_new_n931_));
  NO2        g0909(.A(i_0_), .B(new_new_n712_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n933_));
  INV        g0911(.A(new_new_n933_), .Y(new_new_n934_));
  NO3        g0912(.A(new_new_n107_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n935_));
  AO220      g0913(.A0(new_new_n935_), .A1(new_new_n934_), .B0(new_new_n932_), .B1(new_new_n175_), .Y(new_new_n936_));
  NO2        g0914(.A(new_new_n788_), .B(new_new_n895_), .Y(new_new_n937_));
  AOI210     g0915(.A0(new_new_n936_), .A1(new_new_n345_), .B0(new_new_n937_), .Y(new_new_n938_));
  NA2        g0916(.A(new_new_n723_), .B(new_new_n147_), .Y(new_new_n939_));
  INV        g0917(.A(new_new_n939_), .Y(new_new_n940_));
  NA3        g0918(.A(new_new_n940_), .B(new_new_n661_), .C(new_new_n73_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n806_), .B(new_new_n391_), .Y(new_new_n942_));
  NA3        g0920(.A(new_new_n833_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n943_));
  NA2        g0921(.A(new_new_n834_), .B(i_9_), .Y(new_new_n944_));
  AOI210     g0922(.A0(new_new_n943_), .A1(new_new_n488_), .B0(new_new_n944_), .Y(new_new_n945_));
  OAI210     g0923(.A0(new_new_n244_), .A1(i_9_), .B0(new_new_n230_), .Y(new_new_n946_));
  AOI210     g0924(.A0(new_new_n946_), .A1(new_new_n866_), .B0(new_new_n154_), .Y(new_new_n947_));
  NO3        g0925(.A(new_new_n947_), .B(new_new_n945_), .C(new_new_n942_), .Y(new_new_n948_));
  NA3        g0926(.A(new_new_n948_), .B(new_new_n941_), .C(new_new_n938_), .Y(new_new_n949_));
  NA2        g0927(.A(new_new_n910_), .B(new_new_n369_), .Y(new_new_n950_));
  AOI210     g0928(.A0(new_new_n297_), .A1(new_new_n163_), .B0(new_new_n950_), .Y(new_new_n951_));
  NA3        g0929(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n952_));
  NA2        g0930(.A(new_new_n885_), .B(new_new_n476_), .Y(new_new_n953_));
  AOI210     g0931(.A0(new_new_n952_), .A1(new_new_n163_), .B0(new_new_n953_), .Y(new_new_n954_));
  NO2        g0932(.A(new_new_n954_), .B(new_new_n951_), .Y(new_new_n955_));
  NO3        g0933(.A(new_new_n873_), .B(new_new_n849_), .C(new_new_n192_), .Y(new_new_n956_));
  AOI220     g0934(.A0(new_new_n956_), .A1(i_11_), .B0(new_new_n555_), .B1(new_new_n75_), .Y(new_new_n957_));
  NO3        g0935(.A(new_new_n211_), .B(new_new_n378_), .C(i_0_), .Y(new_new_n958_));
  OAI210     g0936(.A0(new_new_n958_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n959_));
  INV        g0937(.A(new_new_n219_), .Y(new_new_n960_));
  OAI220     g0938(.A0(new_new_n524_), .A1(new_new_n140_), .B0(new_new_n628_), .B1(new_new_n602_), .Y(new_new_n961_));
  NA3        g0939(.A(new_new_n961_), .B(new_new_n386_), .C(new_new_n960_), .Y(new_new_n962_));
  NA4        g0940(.A(new_new_n962_), .B(new_new_n959_), .C(new_new_n957_), .D(new_new_n955_), .Y(new_new_n963_));
  NO2        g0941(.A(new_new_n243_), .B(new_new_n95_), .Y(new_new_n964_));
  AOI210     g0942(.A0(new_new_n964_), .A1(new_new_n932_), .B0(new_new_n111_), .Y(new_new_n965_));
  AOI220     g0943(.A0(new_new_n900_), .A1(new_new_n476_), .B0(new_new_n833_), .B1(new_new_n164_), .Y(new_new_n966_));
  NA2        g0944(.A(new_new_n348_), .B(new_new_n177_), .Y(new_new_n967_));
  OA220      g0945(.A0(new_new_n967_), .A1(new_new_n966_), .B0(new_new_n965_), .B1(i_5_), .Y(new_new_n968_));
  AOI210     g0946(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n176_), .Y(new_new_n969_));
  NA2        g0947(.A(new_new_n969_), .B(new_new_n913_), .Y(new_new_n970_));
  NA3        g0948(.A(new_new_n599_), .B(new_new_n187_), .C(new_new_n84_), .Y(new_new_n971_));
  INV        g0949(.A(new_new_n971_), .Y(new_new_n972_));
  NO3        g0950(.A(new_new_n841_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n973_));
  NA2        g0951(.A(new_new_n481_), .B(new_new_n474_), .Y(new_new_n974_));
  NO3        g0952(.A(new_new_n974_), .B(new_new_n973_), .C(new_new_n972_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n885_), .B(new_new_n291_), .C(new_new_n230_), .Y(new_new_n976_));
  INV        g0954(.A(new_new_n976_), .Y(new_new_n977_));
  NO3        g0955(.A(new_new_n882_), .B(new_new_n219_), .C(new_new_n192_), .Y(new_new_n978_));
  NO2        g0956(.A(new_new_n978_), .B(new_new_n977_), .Y(new_new_n979_));
  NA4        g0957(.A(new_new_n979_), .B(new_new_n975_), .C(new_new_n970_), .D(new_new_n968_), .Y(new_new_n980_));
  INV        g0958(.A(new_new_n601_), .Y(new_new_n981_));
  NO3        g0959(.A(new_new_n981_), .B(new_new_n547_), .C(new_new_n342_), .Y(new_new_n982_));
  INV        g0960(.A(new_new_n982_), .Y(new_new_n983_));
  NA2        g0961(.A(new_new_n302_), .B(i_5_), .Y(new_new_n984_));
  NA2        g0962(.A(new_new_n984_), .B(new_new_n243_), .Y(new_new_n985_));
  NO4        g0963(.A(new_new_n240_), .B(new_new_n211_), .C(i_0_), .D(i_12_), .Y(new_new_n986_));
  AOI220     g0964(.A0(new_new_n986_), .A1(new_new_n985_), .B0(new_new_n782_), .B1(new_new_n177_), .Y(new_new_n987_));
  NA3        g0965(.A(new_new_n100_), .B(new_new_n559_), .C(i_11_), .Y(new_new_n988_));
  NO2        g0966(.A(new_new_n988_), .B(new_new_n156_), .Y(new_new_n989_));
  NA2        g0967(.A(new_new_n900_), .B(new_new_n458_), .Y(new_new_n990_));
  NA2        g0968(.A(new_new_n64_), .B(new_new_n103_), .Y(new_new_n991_));
  OAI220     g0969(.A0(new_new_n991_), .A1(new_new_n984_), .B0(new_new_n990_), .B1(new_new_n662_), .Y(new_new_n992_));
  AOI210     g0970(.A0(new_new_n992_), .A1(new_new_n888_), .B0(new_new_n989_), .Y(new_new_n993_));
  NA3        g0971(.A(new_new_n993_), .B(new_new_n987_), .C(new_new_n983_), .Y(new_new_n994_));
  NO4        g0972(.A(new_new_n994_), .B(new_new_n980_), .C(new_new_n963_), .D(new_new_n949_), .Y(new_new_n995_));
  OAI210     g0973(.A0(new_new_n809_), .A1(new_new_n802_), .B0(new_new_n37_), .Y(new_new_n996_));
  NA3        g0974(.A(new_new_n894_), .B(new_new_n364_), .C(i_5_), .Y(new_new_n997_));
  NA3        g0975(.A(new_new_n997_), .B(new_new_n996_), .C(new_new_n597_), .Y(new_new_n998_));
  NA2        g0976(.A(new_new_n998_), .B(new_new_n208_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n188_), .B(new_new_n190_), .Y(new_new_n1000_));
  AO210      g0978(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n1000_), .Y(new_new_n1001_));
  OAI210     g0979(.A0(new_new_n601_), .A1(new_new_n599_), .B0(new_new_n315_), .Y(new_new_n1002_));
  NAi31      g0980(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1003_));
  NO2        g0981(.A(new_new_n70_), .B(new_new_n1003_), .Y(new_new_n1004_));
  NO2        g0982(.A(new_new_n1004_), .B(new_new_n629_), .Y(new_new_n1005_));
  NA3        g0983(.A(new_new_n1005_), .B(new_new_n1002_), .C(new_new_n1001_), .Y(new_new_n1006_));
  NO2        g0984(.A(new_new_n449_), .B(new_new_n269_), .Y(new_new_n1007_));
  NO4        g0985(.A(new_new_n233_), .B(new_new_n146_), .C(new_new_n665_), .D(new_new_n37_), .Y(new_new_n1008_));
  NO2        g0986(.A(new_new_n1008_), .B(new_new_n1007_), .Y(new_new_n1009_));
  OAI210     g0987(.A0(new_new_n988_), .A1(new_new_n149_), .B0(new_new_n1009_), .Y(new_new_n1010_));
  AOI210     g0988(.A0(new_new_n1006_), .A1(new_new_n49_), .B0(new_new_n1010_), .Y(new_new_n1011_));
  AOI210     g0989(.A0(new_new_n1011_), .A1(new_new_n999_), .B0(new_new_n73_), .Y(new_new_n1012_));
  NO2        g0990(.A(new_new_n552_), .B(new_new_n374_), .Y(new_new_n1013_));
  NO2        g0991(.A(new_new_n1013_), .B(new_new_n743_), .Y(new_new_n1014_));
  INV        g0992(.A(new_new_n76_), .Y(new_new_n1015_));
  AOI210     g0993(.A0(new_new_n969_), .A1(new_new_n885_), .B0(new_new_n901_), .Y(new_new_n1016_));
  AOI210     g0994(.A0(new_new_n1016_), .A1(new_new_n1015_), .B0(new_new_n665_), .Y(new_new_n1017_));
  NA2        g0995(.A(new_new_n263_), .B(new_new_n57_), .Y(new_new_n1018_));
  AOI220     g0996(.A0(new_new_n1018_), .A1(new_new_n76_), .B0(new_new_n343_), .B1(new_new_n256_), .Y(new_new_n1019_));
  NO2        g0997(.A(new_new_n1019_), .B(new_new_n237_), .Y(new_new_n1020_));
  NA3        g0998(.A(new_new_n98_), .B(new_new_n304_), .C(new_new_n31_), .Y(new_new_n1021_));
  INV        g0999(.A(new_new_n1021_), .Y(new_new_n1022_));
  NO3        g1000(.A(new_new_n1022_), .B(new_new_n1020_), .C(new_new_n1017_), .Y(new_new_n1023_));
  OAI210     g1001(.A0(new_new_n271_), .A1(new_new_n159_), .B0(new_new_n89_), .Y(new_new_n1024_));
  NO2        g1002(.A(new_new_n1024_), .B(i_11_), .Y(new_new_n1025_));
  NA2        g1003(.A(new_new_n592_), .B(new_new_n217_), .Y(new_new_n1026_));
  OAI210     g1004(.A0(new_new_n1026_), .A1(new_new_n894_), .B0(new_new_n208_), .Y(new_new_n1027_));
  NA2        g1005(.A(new_new_n165_), .B(i_5_), .Y(new_new_n1028_));
  NO2        g1006(.A(new_new_n1027_), .B(new_new_n1028_), .Y(new_new_n1029_));
  NO3        g1007(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1030_));
  OAI210     g1008(.A0(new_new_n905_), .A1(new_new_n304_), .B0(new_new_n1030_), .Y(new_new_n1031_));
  NO2        g1009(.A(new_new_n1031_), .B(new_new_n712_), .Y(new_new_n1032_));
  NO4        g1010(.A(new_new_n924_), .B(new_new_n464_), .C(new_new_n253_), .D(new_new_n252_), .Y(new_new_n1033_));
  NO2        g1011(.A(new_new_n1033_), .B(new_new_n549_), .Y(new_new_n1034_));
  NO2        g1012(.A(new_new_n1034_), .B(new_new_n41_), .Y(new_new_n1035_));
  NO4        g1013(.A(new_new_n1035_), .B(new_new_n1032_), .C(new_new_n1029_), .D(new_new_n1025_), .Y(new_new_n1036_));
  OAI210     g1014(.A0(new_new_n1023_), .A1(i_4_), .B0(new_new_n1036_), .Y(new_new_n1037_));
  NO3        g1015(.A(new_new_n1037_), .B(new_new_n1014_), .C(new_new_n1012_), .Y(new_new_n1038_));
  NA4        g1016(.A(new_new_n1038_), .B(new_new_n995_), .C(new_new_n931_), .D(new_new_n857_), .Y(men4));
  INV        g1017(.A(new_new_n685_), .Y(new_new_n1042_));
  INV        g1018(.A(new_new_n119_), .Y(new_new_n1043_));
endmodule


