//Benchmark atmr_9sym_175_0.5

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, ori00, mai00, men00;
  ONE        o0(.Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  INV        m002(.A(i_5_), .Y(mai_mai_n13_));
  NOi21      m003(.An(i_3_), .B(i_7_), .Y(mai_mai_n14_));
  INV        m004(.A(i_0_), .Y(mai_mai_n15_));
  NOi21      m005(.An(i_1_), .B(i_3_), .Y(mai_mai_n16_));
  INV        m006(.A(i_4_), .Y(mai_mai_n17_));
  NA2        m007(.A(i_0_), .B(mai_mai_n17_), .Y(mai_mai_n18_));
  INV        m008(.A(i_7_), .Y(mai_mai_n19_));
  NA3        m009(.A(i_6_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n20_));
  NOi21      m010(.An(i_8_), .B(i_6_), .Y(mai_mai_n21_));
  NO2        m011(.A(mai_mai_n20_), .B(mai_mai_n18_), .Y(mai_mai_n22_));
  NA2        m012(.A(mai_mai_n22_), .B(mai_mai_n11_), .Y(mai_mai_n23_));
  NA2        m013(.A(i_0_), .B(mai_mai_n13_), .Y(mai_mai_n24_));
  NA2        m014(.A(mai_mai_n15_), .B(i_5_), .Y(mai_mai_n25_));
  NO2        m015(.A(i_2_), .B(i_4_), .Y(mai_mai_n26_));
  NA3        m016(.A(mai_mai_n26_), .B(i_6_), .C(i_8_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n27_), .Y(mai_mai_n28_));
  INV        m018(.A(i_2_), .Y(mai_mai_n29_));
  NOi21      m019(.An(i_5_), .B(i_0_), .Y(mai_mai_n30_));
  NOi21      m020(.An(i_6_), .B(i_8_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_7_), .B(i_1_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_5_), .B(i_6_), .Y(mai_mai_n33_));
  AOI220     m023(.A0(mai_mai_n33_), .A1(mai_mai_n32_), .B0(mai_mai_n31_), .B1(mai_mai_n30_), .Y(mai_mai_n34_));
  NO3        m024(.A(mai_mai_n34_), .B(mai_mai_n29_), .C(i_4_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_0_), .B(i_4_), .Y(mai_mai_n36_));
  XO2        m026(.A(i_1_), .B(i_3_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_7_), .B(i_5_), .Y(mai_mai_n38_));
  AN3        m028(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n36_), .Y(mai_mai_n39_));
  INV        m029(.A(i_1_), .Y(mai_mai_n40_));
  NOi21      m030(.An(i_3_), .B(i_0_), .Y(mai_mai_n41_));
  NA2        m031(.A(mai_mai_n41_), .B(mai_mai_n40_), .Y(mai_mai_n42_));
  NA3        m032(.A(i_6_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n43_));
  AOI210     m033(.A0(mai_mai_n43_), .A1(mai_mai_n20_), .B0(mai_mai_n42_), .Y(mai_mai_n44_));
  NO4        m034(.A(mai_mai_n44_), .B(mai_mai_n39_), .C(mai_mai_n35_), .D(mai_mai_n28_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_4_), .B(i_0_), .Y(mai_mai_n46_));
  AOI210     m036(.A0(mai_mai_n46_), .A1(mai_mai_n21_), .B0(mai_mai_n14_), .Y(mai_mai_n47_));
  NA2        m037(.A(i_1_), .B(mai_mai_n13_), .Y(mai_mai_n48_));
  NOi21      m038(.An(i_2_), .B(i_8_), .Y(mai_mai_n49_));
  NO3        m039(.A(mai_mai_n49_), .B(mai_mai_n46_), .C(mai_mai_n36_), .Y(mai_mai_n50_));
  NO3        m040(.A(mai_mai_n50_), .B(mai_mai_n48_), .C(mai_mai_n47_), .Y(mai_mai_n51_));
  INV        m041(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_4_), .B(i_3_), .Y(mai_mai_n53_));
  NOi21      m043(.An(i_1_), .B(i_4_), .Y(mai_mai_n54_));
  OAI210     m044(.A0(mai_mai_n54_), .A1(mai_mai_n53_), .B0(mai_mai_n49_), .Y(mai_mai_n55_));
  INV        m045(.A(mai_mai_n55_), .Y(mai_mai_n56_));
  AN2        m046(.A(i_8_), .B(i_7_), .Y(mai_mai_n57_));
  NA2        m047(.A(mai_mai_n57_), .B(mai_mai_n12_), .Y(mai_mai_n58_));
  NOi21      m048(.An(i_8_), .B(i_7_), .Y(mai_mai_n59_));
  NA3        m049(.A(mai_mai_n59_), .B(mai_mai_n53_), .C(i_6_), .Y(mai_mai_n60_));
  OAI210     m050(.A0(mai_mai_n58_), .A1(mai_mai_n48_), .B0(mai_mai_n60_), .Y(mai_mai_n61_));
  AOI220     m051(.A0(mai_mai_n61_), .A1(mai_mai_n29_), .B0(mai_mai_n56_), .B1(mai_mai_n33_), .Y(mai_mai_n62_));
  NA4        m052(.A(mai_mai_n62_), .B(mai_mai_n52_), .C(mai_mai_n45_), .D(mai_mai_n23_), .Y(mai_mai_n63_));
  NA2        m053(.A(i_8_), .B(mai_mai_n19_), .Y(mai_mai_n64_));
  AOI220     m054(.A0(mai_mai_n41_), .A1(i_1_), .B0(mai_mai_n37_), .B1(i_2_), .Y(mai_mai_n65_));
  NOi21      m055(.An(i_1_), .B(i_2_), .Y(mai_mai_n66_));
  NA3        m056(.A(mai_mai_n66_), .B(mai_mai_n46_), .C(i_6_), .Y(mai_mai_n67_));
  OAI210     m057(.A0(mai_mai_n65_), .A1(mai_mai_n64_), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  NA2        m058(.A(mai_mai_n68_), .B(mai_mai_n13_), .Y(mai_mai_n69_));
  NA3        m059(.A(mai_mai_n59_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n70_));
  INV        m060(.A(mai_mai_n70_), .Y(mai_mai_n71_));
  NA2        m061(.A(mai_mai_n71_), .B(mai_mai_n53_), .Y(mai_mai_n72_));
  NA2        m062(.A(mai_mai_n72_), .B(mai_mai_n69_), .Y(mai_mai_n73_));
  NA2        m063(.A(mai_mai_n31_), .B(mai_mai_n30_), .Y(mai_mai_n74_));
  NOi21      m064(.An(i_7_), .B(i_8_), .Y(mai_mai_n75_));
  INV        m065(.A(mai_mai_n74_), .Y(mai_mai_n76_));
  NA2        m066(.A(mai_mai_n76_), .B(mai_mai_n66_), .Y(mai_mai_n77_));
  AOI220     m067(.A0(mai_mai_n41_), .A1(mai_mai_n40_), .B0(mai_mai_n16_), .B1(mai_mai_n29_), .Y(mai_mai_n78_));
  NA3        m068(.A(mai_mai_n17_), .B(i_5_), .C(i_7_), .Y(mai_mai_n79_));
  NO2        m069(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  INV        m070(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NA3        m071(.A(mai_mai_n59_), .B(mai_mai_n29_), .C(i_3_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n40_), .B(i_6_), .Y(mai_mai_n83_));
  AOI210     m073(.A0(mai_mai_n83_), .A1(mai_mai_n18_), .B0(mai_mai_n82_), .Y(mai_mai_n84_));
  NAi21      m074(.An(i_6_), .B(i_0_), .Y(mai_mai_n85_));
  NA3        m075(.A(mai_mai_n54_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n86_));
  NOi21      m076(.An(i_4_), .B(i_6_), .Y(mai_mai_n87_));
  NOi21      m077(.An(i_5_), .B(i_3_), .Y(mai_mai_n88_));
  NA3        m078(.A(mai_mai_n88_), .B(mai_mai_n66_), .C(mai_mai_n87_), .Y(mai_mai_n89_));
  OAI210     m079(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NA2        m080(.A(mai_mai_n66_), .B(mai_mai_n31_), .Y(mai_mai_n91_));
  NOi21      m081(.An(mai_mai_n38_), .B(mai_mai_n91_), .Y(mai_mai_n92_));
  NO3        m082(.A(mai_mai_n92_), .B(mai_mai_n90_), .C(mai_mai_n84_), .Y(mai_mai_n93_));
  NOi21      m083(.An(i_6_), .B(i_1_), .Y(mai_mai_n94_));
  AOI220     m084(.A0(mai_mai_n94_), .A1(i_7_), .B0(mai_mai_n21_), .B1(i_5_), .Y(mai_mai_n95_));
  NOi31      m085(.An(mai_mai_n46_), .B(mai_mai_n95_), .C(i_2_), .Y(mai_mai_n96_));
  INV        m086(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NA4        m087(.A(mai_mai_n97_), .B(mai_mai_n93_), .C(mai_mai_n81_), .D(mai_mai_n77_), .Y(mai_mai_n98_));
  NA3        m088(.A(mai_mai_n31_), .B(i_2_), .C(mai_mai_n13_), .Y(mai_mai_n99_));
  INV        m089(.A(mai_mai_n99_), .Y(mai_mai_n100_));
  NA2        m090(.A(mai_mai_n100_), .B(mai_mai_n36_), .Y(mai_mai_n101_));
  NA2        m091(.A(mai_mai_n53_), .B(mai_mai_n32_), .Y(mai_mai_n102_));
  AOI210     m092(.A0(mai_mai_n102_), .A1(mai_mai_n70_), .B0(mai_mai_n25_), .Y(mai_mai_n103_));
  NOi21      m093(.An(i_0_), .B(i_2_), .Y(mai_mai_n104_));
  NA3        m094(.A(mai_mai_n104_), .B(mai_mai_n32_), .C(mai_mai_n87_), .Y(mai_mai_n105_));
  NA3        m095(.A(mai_mai_n46_), .B(mai_mai_n38_), .C(mai_mai_n16_), .Y(mai_mai_n106_));
  NA3        m096(.A(mai_mai_n104_), .B(mai_mai_n53_), .C(mai_mai_n31_), .Y(mai_mai_n107_));
  NA3        m097(.A(mai_mai_n107_), .B(mai_mai_n106_), .C(mai_mai_n105_), .Y(mai_mai_n108_));
  NO2        m098(.A(mai_mai_n108_), .B(mai_mai_n103_), .Y(mai_mai_n109_));
  NA2        m099(.A(mai_mai_n75_), .B(mai_mai_n12_), .Y(mai_mai_n110_));
  NA3        m100(.A(i_2_), .B(i_1_), .C(mai_mai_n13_), .Y(mai_mai_n111_));
  NA2        m101(.A(mai_mai_n46_), .B(i_3_), .Y(mai_mai_n112_));
  AOI210     m102(.A0(mai_mai_n112_), .A1(mai_mai_n111_), .B0(mai_mai_n110_), .Y(mai_mai_n113_));
  NA3        m103(.A(mai_mai_n104_), .B(mai_mai_n59_), .C(mai_mai_n87_), .Y(mai_mai_n114_));
  OAI210     m104(.A0(mai_mai_n82_), .A1(mai_mai_n25_), .B0(mai_mai_n114_), .Y(mai_mai_n115_));
  NA4        m105(.A(mai_mai_n88_), .B(mai_mai_n57_), .C(mai_mai_n40_), .D(mai_mai_n17_), .Y(mai_mai_n116_));
  NA3        m106(.A(mai_mai_n49_), .B(mai_mai_n30_), .C(mai_mai_n14_), .Y(mai_mai_n117_));
  NA2        m107(.A(mai_mai_n117_), .B(mai_mai_n116_), .Y(mai_mai_n118_));
  NO3        m108(.A(mai_mai_n118_), .B(mai_mai_n115_), .C(mai_mai_n113_), .Y(mai_mai_n119_));
  NA3        m109(.A(mai_mai_n119_), .B(mai_mai_n109_), .C(mai_mai_n101_), .Y(mai_mai_n120_));
  OR4        m110(.A(mai_mai_n120_), .B(mai_mai_n98_), .C(mai_mai_n73_), .D(mai_mai_n63_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  NOi21      u014(.An(i_1_), .B(i_8_), .Y(men_men_n25_));
  AOI220     u015(.A0(men_men_n25_), .A1(i_2_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n26_));
  NO2        u016(.A(men_men_n26_), .B(men_men_n22_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n28_));
  NA2        u018(.A(i_0_), .B(men_men_n14_), .Y(men_men_n29_));
  NO2        u019(.A(i_2_), .B(i_4_), .Y(men_men_n30_));
  INV        u020(.A(i_2_), .Y(men_men_n31_));
  NOi21      u021(.An(i_6_), .B(i_8_), .Y(men_men_n32_));
  NOi21      u022(.An(i_5_), .B(i_6_), .Y(men_men_n33_));
  NOi21      u023(.An(i_0_), .B(i_4_), .Y(men_men_n34_));
  INV        u024(.A(i_1_), .Y(men_men_n35_));
  NOi21      u025(.An(i_3_), .B(i_0_), .Y(men_men_n36_));
  INV        u026(.A(i_8_), .Y(men_men_n37_));
  NA2        u027(.A(i_1_), .B(men_men_n11_), .Y(men_men_n38_));
  NO4        u028(.A(men_men_n38_), .B(men_men_n29_), .C(i_2_), .D(men_men_n37_), .Y(men_men_n39_));
  NOi21      u029(.An(i_4_), .B(i_0_), .Y(men_men_n40_));
  NOi21      u030(.An(i_2_), .B(i_8_), .Y(men_men_n41_));
  INV        u031(.A(men_men_n39_), .Y(men_men_n42_));
  NOi31      u032(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n43_));
  NA2        u033(.A(men_men_n43_), .B(i_0_), .Y(men_men_n44_));
  NOi21      u034(.An(i_4_), .B(i_3_), .Y(men_men_n45_));
  NOi21      u035(.An(i_1_), .B(i_4_), .Y(men_men_n46_));
  INV        u036(.A(men_men_n44_), .Y(men_men_n47_));
  AN2        u037(.A(i_8_), .B(i_7_), .Y(men_men_n48_));
  NOi21      u038(.An(i_8_), .B(i_7_), .Y(men_men_n49_));
  NA2        u039(.A(men_men_n47_), .B(men_men_n33_), .Y(men_men_n50_));
  NA3        u040(.A(men_men_n50_), .B(men_men_n42_), .C(men_men_n28_), .Y(men_men_n51_));
  NA2        u041(.A(i_8_), .B(i_7_), .Y(men_men_n52_));
  NO3        u042(.A(men_men_n52_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n53_));
  NOi21      u043(.An(i_1_), .B(i_2_), .Y(men_men_n54_));
  NA2        u044(.A(men_men_n53_), .B(men_men_n14_), .Y(men_men_n55_));
  NA3        u045(.A(men_men_n25_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n56_));
  INV        u046(.A(men_men_n56_), .Y(men_men_n57_));
  NOi32      u047(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n58_), .B(i_3_), .Y(men_men_n59_));
  NA3        u049(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n60_));
  NA2        u050(.A(men_men_n60_), .B(men_men_n59_), .Y(men_men_n61_));
  NO2        u051(.A(i_0_), .B(i_4_), .Y(men_men_n62_));
  AOI220     u052(.A0(men_men_n62_), .A1(men_men_n61_), .B0(men_men_n57_), .B1(men_men_n45_), .Y(men_men_n63_));
  NA2        u053(.A(men_men_n63_), .B(men_men_n55_), .Y(men_men_n64_));
  NAi21      u054(.An(i_3_), .B(i_6_), .Y(men_men_n65_));
  NO3        u055(.A(men_men_n65_), .B(i_0_), .C(men_men_n37_), .Y(men_men_n66_));
  NOi21      u056(.An(i_7_), .B(i_8_), .Y(men_men_n67_));
  NOi31      u057(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n68_));
  AOI210     u058(.A0(men_men_n67_), .A1(men_men_n12_), .B0(men_men_n68_), .Y(men_men_n69_));
  NO2        u059(.A(men_men_n69_), .B(men_men_n11_), .Y(men_men_n70_));
  OAI210     u060(.A0(men_men_n70_), .A1(men_men_n66_), .B0(men_men_n54_), .Y(men_men_n71_));
  NA3        u061(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n72_));
  AOI210     u062(.A0(men_men_n22_), .A1(men_men_n38_), .B0(men_men_n72_), .Y(men_men_n73_));
  OAI210     u063(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n74_));
  NA3        u064(.A(men_men_n52_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n75_));
  NO2        u065(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  NO2        u066(.A(men_men_n76_), .B(men_men_n73_), .Y(men_men_n77_));
  NA2        u067(.A(men_men_n35_), .B(i_6_), .Y(men_men_n78_));
  NOi21      u068(.An(i_2_), .B(i_1_), .Y(men_men_n79_));
  AN3        u069(.A(men_men_n67_), .B(men_men_n79_), .C(men_men_n40_), .Y(men_men_n80_));
  NAi21      u070(.An(i_6_), .B(i_0_), .Y(men_men_n81_));
  NOi21      u071(.An(i_4_), .B(i_6_), .Y(men_men_n82_));
  NA2        u072(.A(men_men_n54_), .B(men_men_n32_), .Y(men_men_n83_));
  INV        u073(.A(men_men_n80_), .Y(men_men_n84_));
  NA2        u074(.A(men_men_n49_), .B(men_men_n12_), .Y(men_men_n85_));
  NA2        u075(.A(men_men_n32_), .B(men_men_n14_), .Y(men_men_n86_));
  NOi21      u076(.An(i_3_), .B(i_1_), .Y(men_men_n87_));
  NA2        u077(.A(men_men_n87_), .B(i_4_), .Y(men_men_n88_));
  AOI210     u078(.A0(men_men_n86_), .A1(men_men_n85_), .B0(men_men_n88_), .Y(men_men_n89_));
  AOI220     u079(.A0(men_men_n67_), .A1(men_men_n14_), .B0(men_men_n82_), .B1(men_men_n23_), .Y(men_men_n90_));
  NOi31      u080(.An(men_men_n36_), .B(men_men_n90_), .C(men_men_n31_), .Y(men_men_n91_));
  NO2        u081(.A(men_men_n91_), .B(men_men_n89_), .Y(men_men_n92_));
  NA4        u082(.A(men_men_n92_), .B(men_men_n84_), .C(men_men_n77_), .D(men_men_n71_), .Y(men_men_n93_));
  NA2        u083(.A(men_men_n41_), .B(men_men_n15_), .Y(men_men_n94_));
  NOi31      u084(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n95_));
  NOi31      u085(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n96_));
  OAI210     u086(.A0(men_men_n96_), .A1(men_men_n95_), .B0(i_7_), .Y(men_men_n97_));
  NA3        u087(.A(men_men_n97_), .B(men_men_n94_), .C(men_men_n83_), .Y(men_men_n98_));
  NA2        u088(.A(men_men_n98_), .B(men_men_n34_), .Y(men_men_n99_));
  NA4        u089(.A(men_men_n48_), .B(men_men_n79_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n100_));
  NAi31      u090(.An(men_men_n81_), .B(men_men_n67_), .C(men_men_n79_), .Y(men_men_n101_));
  NA3        u091(.A(men_men_n49_), .B(men_men_n43_), .C(i_6_), .Y(men_men_n102_));
  NA3        u092(.A(men_men_n102_), .B(men_men_n101_), .C(men_men_n100_), .Y(men_men_n103_));
  NOi32      u093(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n104_));
  NA2        u094(.A(men_men_n104_), .B(men_men_n95_), .Y(men_men_n105_));
  INV        u095(.A(men_men_n105_), .Y(men_men_n106_));
  NA4        u096(.A(men_men_n43_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n107_));
  NA4        u097(.A(men_men_n46_), .B(men_men_n33_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n108_));
  NA4        u098(.A(men_men_n46_), .B(men_men_n36_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n109_));
  NA3        u099(.A(men_men_n109_), .B(men_men_n108_), .C(men_men_n107_), .Y(men_men_n110_));
  NO3        u100(.A(men_men_n110_), .B(men_men_n106_), .C(men_men_n103_), .Y(men_men_n111_));
  NOi21      u101(.An(i_5_), .B(i_2_), .Y(men_men_n112_));
  AOI220     u102(.A0(men_men_n112_), .A1(men_men_n67_), .B0(men_men_n48_), .B1(men_men_n30_), .Y(men_men_n113_));
  AOI210     u103(.A0(men_men_n113_), .A1(men_men_n94_), .B0(men_men_n78_), .Y(men_men_n114_));
  NO4        u104(.A(i_2_), .B(men_men_n21_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n115_));
  NA2        u105(.A(i_2_), .B(i_4_), .Y(men_men_n116_));
  AOI210     u106(.A0(men_men_n81_), .A1(men_men_n65_), .B0(men_men_n116_), .Y(men_men_n117_));
  NO2        u107(.A(i_8_), .B(i_7_), .Y(men_men_n118_));
  OA210      u108(.A0(men_men_n117_), .A1(men_men_n115_), .B0(men_men_n118_), .Y(men_men_n119_));
  NA4        u109(.A(men_men_n87_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n120_));
  NO2        u110(.A(men_men_n120_), .B(i_4_), .Y(men_men_n121_));
  NO3        u111(.A(men_men_n121_), .B(men_men_n119_), .C(men_men_n114_), .Y(men_men_n122_));
  NA3        u112(.A(men_men_n68_), .B(men_men_n87_), .C(i_0_), .Y(men_men_n123_));
  NOi31      u113(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n124_));
  OAI210     u114(.A0(men_men_n104_), .A1(men_men_n58_), .B0(men_men_n124_), .Y(men_men_n125_));
  NA2        u115(.A(men_men_n125_), .B(men_men_n123_), .Y(men_men_n126_));
  INV        u116(.A(men_men_n126_), .Y(men_men_n127_));
  NA4        u117(.A(men_men_n127_), .B(men_men_n122_), .C(men_men_n111_), .D(men_men_n99_), .Y(men_men_n128_));
  OR4        u118(.A(men_men_n128_), .B(men_men_n93_), .C(men_men_n64_), .D(men_men_n51_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule