// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n141_, new_new_n142_, new_new_n143_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1009_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g040(.A(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g063(.A(i_6_), .Y(new_new_n86_));
  OR4        g064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  NO2        g067(.A(new_new_n88_), .B(new_new_n89_), .Y(new_new_n90_));
  OAI210     g068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  NO3        g073(.A(new_new_n95_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n96_));
  NO2        g074(.A(new_new_n96_), .B(new_new_n94_), .Y(new_new_n97_));
  AOI210     g075(.A0(new_new_n97_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n98_));
  AN3        g076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n99_));
  NAi21      g077(.An(i_6_), .B(i_11_), .Y(new_new_n100_));
  NO2        g078(.A(i_5_), .B(i_8_), .Y(new_new_n101_));
  NOi21      g079(.An(new_new_n101_), .B(new_new_n100_), .Y(new_new_n102_));
  AOI220     g080(.A0(new_new_n102_), .A1(new_new_n62_), .B0(new_new_n99_), .B1(new_new_n32_), .Y(new_new_n103_));
  INV        g081(.A(i_7_), .Y(new_new_n104_));
  NA2        g082(.A(new_new_n46_), .B(new_new_n104_), .Y(new_new_n105_));
  NO2        g083(.A(i_0_), .B(i_5_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(new_new_n86_), .Y(new_new_n107_));
  NA2        g085(.A(i_12_), .B(i_3_), .Y(new_new_n108_));
  INV        g086(.A(new_new_n108_), .Y(new_new_n109_));
  NA3        g087(.A(new_new_n109_), .B(new_new_n107_), .C(new_new_n105_), .Y(new_new_n110_));
  NAi21      g088(.An(i_7_), .B(i_11_), .Y(new_new_n111_));
  NO3        g089(.A(new_new_n111_), .B(new_new_n92_), .C(new_new_n53_), .Y(new_new_n112_));
  AN2        g090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g092(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n115_));
  NO2        g093(.A(i_8_), .B(new_new_n104_), .Y(new_new_n116_));
  NO3        g094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g096(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g097(.A(i_11_), .B(i_12_), .Y(new_new_n120_));
  INV        g098(.A(new_new_n120_), .Y(new_new_n121_));
  NO2        g099(.A(new_new_n121_), .B(new_new_n117_), .Y(new_new_n122_));
  NAi41      g100(.An(new_new_n112_), .B(new_new_n122_), .C(new_new_n110_), .D(new_new_n103_), .Y(new_new_n123_));
  NOi21      g101(.An(i_1_), .B(i_5_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(i_11_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n126_));
  NA2        g104(.A(i_7_), .B(new_new_n25_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(new_new_n126_), .Y(new_new_n128_));
  NO2        g106(.A(new_new_n128_), .B(new_new_n46_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n130_));
  NAi21      g108(.An(i_3_), .B(i_8_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(new_new_n62_), .Y(new_new_n132_));
  NOi31      g110(.An(new_new_n132_), .B(new_new_n130_), .C(new_new_n129_), .Y(new_new_n133_));
  NO2        g111(.A(i_1_), .B(new_new_n86_), .Y(new_new_n134_));
  NO2        g112(.A(i_6_), .B(i_5_), .Y(new_new_n135_));
  NA2        g113(.A(new_new_n135_), .B(i_3_), .Y(new_new_n136_));
  AO210      g114(.A0(new_new_n136_), .A1(new_new_n47_), .B0(new_new_n134_), .Y(new_new_n137_));
  OAI220     g115(.A0(new_new_n137_), .A1(new_new_n111_), .B0(new_new_n133_), .B1(new_new_n125_), .Y(new_new_n138_));
  NO3        g116(.A(new_new_n138_), .B(new_new_n123_), .C(new_new_n98_), .Y(new_new_n139_));
  NA3        g117(.A(new_new_n139_), .B(new_new_n79_), .C(new_new_n56_), .Y(ori2));
  NO2        g118(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n141_));
  NA2        g119(.A(i_6_), .B(new_new_n25_), .Y(new_new_n142_));
  NA2        g120(.A(new_new_n142_), .B(new_new_n141_), .Y(new_new_n143_));
  NA4        g121(.A(new_new_n143_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(ori0));
  AN2        g122(.A(i_8_), .B(i_7_), .Y(new_new_n145_));
  NA2        g123(.A(new_new_n145_), .B(i_6_), .Y(new_new_n146_));
  NO2        g124(.A(i_12_), .B(i_13_), .Y(new_new_n147_));
  NAi21      g125(.An(i_5_), .B(i_11_), .Y(new_new_n148_));
  NOi21      g126(.An(new_new_n147_), .B(new_new_n148_), .Y(new_new_n149_));
  NO2        g127(.A(i_0_), .B(i_1_), .Y(new_new_n150_));
  NA2        g128(.A(i_2_), .B(i_3_), .Y(new_new_n151_));
  NO2        g129(.A(new_new_n151_), .B(i_4_), .Y(new_new_n152_));
  NA3        g130(.A(new_new_n152_), .B(new_new_n150_), .C(new_new_n149_), .Y(new_new_n153_));
  AN2        g131(.A(new_new_n147_), .B(new_new_n83_), .Y(new_new_n154_));
  NO2        g132(.A(new_new_n154_), .B(new_new_n27_), .Y(new_new_n155_));
  NA2        g133(.A(i_1_), .B(i_5_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n73_), .B(new_new_n46_), .Y(new_new_n157_));
  NA2        g135(.A(new_new_n157_), .B(new_new_n36_), .Y(new_new_n158_));
  NO3        g136(.A(new_new_n158_), .B(new_new_n156_), .C(new_new_n155_), .Y(new_new_n159_));
  OR2        g137(.A(i_0_), .B(i_1_), .Y(new_new_n160_));
  NO3        g138(.A(new_new_n160_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n161_));
  NAi32      g139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n162_));
  NAi21      g140(.An(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  NOi21      g141(.An(i_4_), .B(i_10_), .Y(new_new_n164_));
  NA2        g142(.A(new_new_n164_), .B(new_new_n40_), .Y(new_new_n165_));
  NO2        g143(.A(i_3_), .B(i_5_), .Y(new_new_n166_));
  NO3        g144(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n167_));
  NA2        g145(.A(new_new_n167_), .B(new_new_n166_), .Y(new_new_n168_));
  OAI210     g146(.A0(new_new_n168_), .A1(new_new_n165_), .B0(new_new_n163_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n169_), .B(new_new_n159_), .Y(new_new_n170_));
  AOI210     g148(.A0(new_new_n170_), .A1(new_new_n153_), .B0(new_new_n146_), .Y(new_new_n171_));
  NA2        g149(.A(i_3_), .B(new_new_n48_), .Y(new_new_n172_));
  NOi21      g150(.An(i_4_), .B(i_9_), .Y(new_new_n173_));
  NOi21      g151(.An(i_11_), .B(i_13_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n174_), .B(new_new_n173_), .Y(new_new_n175_));
  OR2        g153(.A(new_new_n175_), .B(new_new_n172_), .Y(new_new_n176_));
  NO2        g154(.A(i_4_), .B(i_5_), .Y(new_new_n177_));
  NAi21      g155(.An(i_12_), .B(i_11_), .Y(new_new_n178_));
  NO2        g156(.A(new_new_n178_), .B(i_13_), .Y(new_new_n179_));
  NA3        g157(.A(new_new_n179_), .B(new_new_n177_), .C(new_new_n83_), .Y(new_new_n180_));
  NO2        g158(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n181_));
  NA2        g159(.A(new_new_n181_), .B(new_new_n46_), .Y(new_new_n182_));
  NAi31      g160(.An(i_4_), .B(new_new_n154_), .C(i_11_), .Y(new_new_n183_));
  NA2        g161(.A(i_3_), .B(i_5_), .Y(new_new_n184_));
  OR2        g162(.A(new_new_n184_), .B(new_new_n175_), .Y(new_new_n185_));
  AOI210     g163(.A0(new_new_n185_), .A1(new_new_n183_), .B0(new_new_n182_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n73_), .B(i_5_), .Y(new_new_n187_));
  NO2        g165(.A(i_13_), .B(i_10_), .Y(new_new_n188_));
  NO2        g166(.A(i_2_), .B(i_1_), .Y(new_new_n189_));
  NA2        g167(.A(new_new_n189_), .B(i_3_), .Y(new_new_n190_));
  NAi21      g168(.An(i_4_), .B(i_12_), .Y(new_new_n191_));
  INV        g169(.A(new_new_n186_), .Y(new_new_n192_));
  INV        g170(.A(i_8_), .Y(new_new_n193_));
  NO2        g171(.A(new_new_n193_), .B(i_7_), .Y(new_new_n194_));
  NA2        g172(.A(new_new_n194_), .B(i_6_), .Y(new_new_n195_));
  NO3        g173(.A(i_3_), .B(new_new_n86_), .C(new_new_n48_), .Y(new_new_n196_));
  NA2        g174(.A(new_new_n196_), .B(new_new_n116_), .Y(new_new_n197_));
  NO3        g175(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n198_));
  NA3        g176(.A(new_new_n198_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n199_));
  NO3        g177(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n200_));
  OAI210     g178(.A0(new_new_n99_), .A1(i_12_), .B0(new_new_n200_), .Y(new_new_n201_));
  AOI210     g179(.A0(new_new_n201_), .A1(new_new_n199_), .B0(new_new_n197_), .Y(new_new_n202_));
  NO2        g180(.A(i_3_), .B(i_8_), .Y(new_new_n203_));
  NO3        g181(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n204_));
  NA3        g182(.A(new_new_n204_), .B(new_new_n203_), .C(new_new_n40_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n106_), .B(new_new_n58_), .Y(new_new_n206_));
  INV        g184(.A(new_new_n206_), .Y(new_new_n207_));
  NO2        g185(.A(i_13_), .B(i_9_), .Y(new_new_n208_));
  NAi21      g186(.An(i_12_), .B(i_3_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n44_), .B(i_5_), .Y(new_new_n210_));
  NO3        g188(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n207_), .B(new_new_n205_), .Y(new_new_n212_));
  AOI210     g190(.A0(new_new_n212_), .A1(i_7_), .B0(new_new_n202_), .Y(new_new_n213_));
  OAI220     g191(.A0(new_new_n213_), .A1(i_4_), .B0(new_new_n195_), .B1(new_new_n192_), .Y(new_new_n214_));
  NAi21      g192(.An(i_12_), .B(i_7_), .Y(new_new_n215_));
  NA3        g193(.A(i_13_), .B(new_new_n193_), .C(i_10_), .Y(new_new_n216_));
  NA2        g194(.A(i_0_), .B(i_5_), .Y(new_new_n217_));
  NAi31      g195(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n36_), .B(i_13_), .Y(new_new_n219_));
  NO2        g197(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n221_));
  INV        g199(.A(i_13_), .Y(new_new_n222_));
  NO2        g200(.A(i_12_), .B(new_new_n222_), .Y(new_new_n223_));
  NO2        g201(.A(i_12_), .B(new_new_n37_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n184_), .B(i_4_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  OR2        g204(.A(i_8_), .B(i_7_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n86_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n53_), .B(i_1_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n230_));
  INV        g208(.A(i_12_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n44_), .B(new_new_n231_), .Y(new_new_n232_));
  NO3        g210(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n233_));
  NA2        g211(.A(i_2_), .B(i_1_), .Y(new_new_n234_));
  NO2        g212(.A(new_new_n230_), .B(new_new_n226_), .Y(new_new_n235_));
  NO3        g213(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n236_));
  NAi21      g214(.An(i_4_), .B(i_3_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n237_), .B(new_new_n75_), .Y(new_new_n238_));
  NO2        g216(.A(i_0_), .B(i_6_), .Y(new_new_n239_));
  NOi41      g217(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n240_));
  NO2        g218(.A(new_new_n234_), .B(new_new_n184_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n235_), .B(new_new_n208_), .Y(new_new_n242_));
  NO2        g220(.A(i_11_), .B(new_new_n222_), .Y(new_new_n243_));
  NOi21      g221(.An(i_1_), .B(i_6_), .Y(new_new_n244_));
  NAi21      g222(.An(i_3_), .B(i_7_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n231_), .B(i_9_), .Y(new_new_n246_));
  OR4        g224(.A(new_new_n246_), .B(new_new_n245_), .C(new_new_n244_), .D(new_new_n187_), .Y(new_new_n247_));
  NO2        g225(.A(i_12_), .B(i_3_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n73_), .B(i_5_), .Y(new_new_n249_));
  NA2        g227(.A(i_3_), .B(i_9_), .Y(new_new_n250_));
  NAi21      g228(.An(i_7_), .B(i_10_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n251_), .B(new_new_n250_), .Y(new_new_n252_));
  NA3        g230(.A(new_new_n252_), .B(new_new_n249_), .C(new_new_n64_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n253_), .B(new_new_n247_), .Y(new_new_n254_));
  INV        g232(.A(new_new_n146_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n231_), .B(i_13_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n256_), .B(new_new_n75_), .Y(new_new_n257_));
  AOI220     g235(.A0(new_new_n257_), .A1(new_new_n255_), .B0(new_new_n254_), .B1(new_new_n243_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n227_), .B(new_new_n37_), .Y(new_new_n259_));
  NA2        g237(.A(i_12_), .B(i_6_), .Y(new_new_n260_));
  OR2        g238(.A(i_13_), .B(i_9_), .Y(new_new_n261_));
  NO3        g239(.A(new_new_n261_), .B(new_new_n260_), .C(new_new_n48_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n237_), .B(i_2_), .Y(new_new_n263_));
  NA2        g241(.A(new_new_n243_), .B(i_9_), .Y(new_new_n264_));
  NA2        g242(.A(new_new_n157_), .B(new_new_n63_), .Y(new_new_n265_));
  NO3        g243(.A(i_11_), .B(new_new_n222_), .C(new_new_n25_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n245_), .B(i_8_), .Y(new_new_n267_));
  NO2        g245(.A(i_6_), .B(new_new_n48_), .Y(new_new_n268_));
  NA3        g246(.A(new_new_n268_), .B(new_new_n267_), .C(new_new_n266_), .Y(new_new_n269_));
  NO3        g247(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n270_));
  NA3        g248(.A(new_new_n270_), .B(new_new_n259_), .C(new_new_n223_), .Y(new_new_n271_));
  AOI210     g249(.A0(new_new_n271_), .A1(new_new_n269_), .B0(new_new_n265_), .Y(new_new_n272_));
  INV        g250(.A(new_new_n272_), .Y(new_new_n273_));
  NA3        g251(.A(new_new_n273_), .B(new_new_n258_), .C(new_new_n242_), .Y(new_new_n274_));
  NO3        g252(.A(i_12_), .B(new_new_n222_), .C(new_new_n37_), .Y(new_new_n275_));
  INV        g253(.A(new_new_n275_), .Y(new_new_n276_));
  NA2        g254(.A(i_8_), .B(new_new_n104_), .Y(new_new_n277_));
  NOi21      g255(.An(new_new_n166_), .B(new_new_n86_), .Y(new_new_n278_));
  NO3        g256(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n279_));
  AOI220     g257(.A0(new_new_n279_), .A1(new_new_n196_), .B0(new_new_n278_), .B1(new_new_n229_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(new_new_n277_), .Y(new_new_n281_));
  NO3        g259(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n234_), .B(i_0_), .Y(new_new_n283_));
  AOI220     g261(.A0(new_new_n283_), .A1(new_new_n194_), .B0(new_new_n282_), .B1(new_new_n145_), .Y(new_new_n284_));
  NA2        g262(.A(new_new_n268_), .B(new_new_n26_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n285_), .B(new_new_n284_), .Y(new_new_n286_));
  NA2        g264(.A(i_0_), .B(i_1_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n287_), .B(i_2_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n59_), .B(i_6_), .Y(new_new_n289_));
  NA3        g267(.A(new_new_n289_), .B(new_new_n288_), .C(new_new_n166_), .Y(new_new_n290_));
  OAI210     g268(.A0(new_new_n168_), .A1(new_new_n146_), .B0(new_new_n290_), .Y(new_new_n291_));
  NO3        g269(.A(new_new_n291_), .B(new_new_n286_), .C(new_new_n281_), .Y(new_new_n292_));
  NO2        g270(.A(i_2_), .B(new_new_n104_), .Y(new_new_n293_));
  NA2        g271(.A(i_1_), .B(new_new_n36_), .Y(new_new_n294_));
  BUFFER     g272(.A(new_new_n217_), .Y(new_new_n295_));
  AN2        g273(.A(i_3_), .B(i_10_), .Y(new_new_n296_));
  NO2        g274(.A(i_5_), .B(new_new_n37_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n292_), .B(new_new_n276_), .Y(new_new_n299_));
  NO4        g277(.A(new_new_n299_), .B(new_new_n274_), .C(new_new_n214_), .D(new_new_n171_), .Y(new_new_n300_));
  NO3        g278(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n283_), .B(new_new_n302_), .Y(new_new_n303_));
  NO3        g281(.A(i_6_), .B(new_new_n193_), .C(i_7_), .Y(new_new_n304_));
  NA2        g282(.A(new_new_n304_), .B(new_new_n198_), .Y(new_new_n305_));
  AOI210     g283(.A0(new_new_n305_), .A1(new_new_n303_), .B0(new_new_n172_), .Y(new_new_n306_));
  NO2        g284(.A(i_2_), .B(i_3_), .Y(new_new_n307_));
  OR2        g285(.A(i_0_), .B(i_5_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n217_), .B(new_new_n308_), .Y(new_new_n309_));
  NA4        g287(.A(new_new_n309_), .B(new_new_n228_), .C(new_new_n307_), .D(i_1_), .Y(new_new_n310_));
  NA3        g288(.A(new_new_n283_), .B(new_new_n278_), .C(new_new_n116_), .Y(new_new_n311_));
  NAi21      g289(.An(i_8_), .B(i_7_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n160_), .B(new_new_n46_), .Y(new_new_n313_));
  NA2        g291(.A(new_new_n311_), .B(new_new_n310_), .Y(new_new_n314_));
  OAI210     g292(.A0(new_new_n314_), .A1(new_new_n306_), .B0(i_4_), .Y(new_new_n315_));
  NO2        g293(.A(i_12_), .B(i_10_), .Y(new_new_n316_));
  NOi21      g294(.An(i_5_), .B(i_0_), .Y(new_new_n317_));
  AOI210     g295(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n104_), .Y(new_new_n318_));
  NO4        g296(.A(new_new_n318_), .B(new_new_n294_), .C(new_new_n317_), .D(new_new_n131_), .Y(new_new_n319_));
  NA4        g297(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n319_), .B(new_new_n316_), .Y(new_new_n321_));
  NO2        g299(.A(i_6_), .B(i_8_), .Y(new_new_n322_));
  NOi21      g300(.An(i_0_), .B(i_2_), .Y(new_new_n323_));
  AN2        g301(.A(new_new_n323_), .B(new_new_n322_), .Y(new_new_n324_));
  NO2        g302(.A(i_1_), .B(i_7_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n321_), .B(new_new_n315_), .Y(new_new_n326_));
  NOi21      g304(.An(new_new_n156_), .B(new_new_n107_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n327_), .B(new_new_n127_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n328_), .B(i_3_), .Y(new_new_n329_));
  INV        g307(.A(new_new_n84_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n287_), .B(new_new_n81_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n331_), .B(new_new_n135_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n95_), .B(new_new_n193_), .Y(new_new_n333_));
  NA3        g311(.A(new_new_n295_), .B(new_new_n333_), .C(new_new_n63_), .Y(new_new_n334_));
  AOI210     g312(.A0(new_new_n334_), .A1(new_new_n332_), .B0(new_new_n330_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n193_), .B(i_9_), .Y(new_new_n336_));
  NA2        g314(.A(new_new_n336_), .B(new_new_n206_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n337_), .B(new_new_n46_), .Y(new_new_n338_));
  NO3        g316(.A(new_new_n338_), .B(new_new_n335_), .C(new_new_n286_), .Y(new_new_n339_));
  AOI210     g317(.A0(new_new_n339_), .A1(new_new_n329_), .B0(new_new_n165_), .Y(new_new_n340_));
  AOI210     g318(.A0(new_new_n326_), .A1(new_new_n301_), .B0(new_new_n340_), .Y(new_new_n341_));
  NOi32      g319(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n342_));
  INV        g320(.A(new_new_n342_), .Y(new_new_n343_));
  NAi21      g321(.An(i_0_), .B(i_6_), .Y(new_new_n344_));
  NAi21      g322(.An(i_1_), .B(i_5_), .Y(new_new_n345_));
  NA2        g323(.A(new_new_n345_), .B(new_new_n344_), .Y(new_new_n346_));
  NA2        g324(.A(new_new_n346_), .B(new_new_n25_), .Y(new_new_n347_));
  NO2        g325(.A(new_new_n347_), .B(new_new_n162_), .Y(new_new_n348_));
  NAi41      g326(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n349_));
  OAI220     g327(.A0(new_new_n349_), .A1(new_new_n345_), .B0(new_new_n218_), .B1(new_new_n162_), .Y(new_new_n350_));
  AOI210     g328(.A0(new_new_n349_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n351_));
  NOi32      g329(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n352_));
  NAi21      g330(.An(i_6_), .B(i_1_), .Y(new_new_n353_));
  NA3        g331(.A(new_new_n353_), .B(new_new_n352_), .C(new_new_n46_), .Y(new_new_n354_));
  NO2        g332(.A(new_new_n354_), .B(i_0_), .Y(new_new_n355_));
  OR3        g333(.A(new_new_n355_), .B(new_new_n351_), .C(new_new_n350_), .Y(new_new_n356_));
  NO2        g334(.A(i_1_), .B(new_new_n104_), .Y(new_new_n357_));
  NAi21      g335(.An(i_3_), .B(i_4_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n358_), .B(i_9_), .Y(new_new_n359_));
  AN2        g337(.A(i_6_), .B(i_7_), .Y(new_new_n360_));
  OAI210     g338(.A0(new_new_n360_), .A1(new_new_n357_), .B0(new_new_n359_), .Y(new_new_n361_));
  NA2        g339(.A(i_2_), .B(i_7_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n358_), .B(i_10_), .Y(new_new_n363_));
  NA3        g341(.A(new_new_n363_), .B(new_new_n362_), .C(new_new_n239_), .Y(new_new_n364_));
  AOI210     g342(.A0(new_new_n364_), .A1(new_new_n361_), .B0(new_new_n187_), .Y(new_new_n365_));
  AOI210     g343(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n366_));
  OAI210     g344(.A0(new_new_n366_), .A1(new_new_n189_), .B0(new_new_n363_), .Y(new_new_n367_));
  AOI220     g345(.A0(new_new_n363_), .A1(new_new_n325_), .B0(new_new_n233_), .B1(new_new_n189_), .Y(new_new_n368_));
  AOI210     g346(.A0(new_new_n368_), .A1(new_new_n367_), .B0(i_5_), .Y(new_new_n369_));
  NO4        g347(.A(new_new_n369_), .B(new_new_n365_), .C(new_new_n356_), .D(new_new_n348_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n370_), .B(new_new_n343_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n372_));
  AN2        g350(.A(i_12_), .B(i_5_), .Y(new_new_n373_));
  NO2        g351(.A(i_4_), .B(new_new_n26_), .Y(new_new_n374_));
  NA2        g352(.A(new_new_n374_), .B(new_new_n373_), .Y(new_new_n375_));
  NO2        g353(.A(i_11_), .B(i_6_), .Y(new_new_n376_));
  NA3        g354(.A(new_new_n376_), .B(new_new_n313_), .C(new_new_n222_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n377_), .B(new_new_n375_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n237_), .B(i_5_), .Y(new_new_n379_));
  NO2        g357(.A(i_5_), .B(i_10_), .Y(new_new_n380_));
  AOI220     g358(.A0(new_new_n380_), .A1(new_new_n263_), .B0(new_new_n379_), .B1(new_new_n198_), .Y(new_new_n381_));
  NA2        g359(.A(new_new_n147_), .B(new_new_n45_), .Y(new_new_n382_));
  NO2        g360(.A(new_new_n382_), .B(new_new_n381_), .Y(new_new_n383_));
  OAI210     g361(.A0(new_new_n383_), .A1(new_new_n378_), .B0(new_new_n372_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n153_), .B(new_new_n86_), .Y(new_new_n386_));
  OAI210     g364(.A0(new_new_n386_), .A1(new_new_n378_), .B0(new_new_n385_), .Y(new_new_n387_));
  NO3        g365(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n388_));
  NO2        g366(.A(i_3_), .B(new_new_n104_), .Y(new_new_n389_));
  NO2        g367(.A(i_11_), .B(i_12_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n380_), .B(new_new_n231_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n387_), .B(new_new_n384_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n44_), .B(new_new_n222_), .Y(new_new_n393_));
  NO3        g371(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n394_));
  NO2        g372(.A(i_0_), .B(i_11_), .Y(new_new_n395_));
  INV        g373(.A(i_5_), .Y(new_new_n396_));
  AN2        g374(.A(i_1_), .B(i_6_), .Y(new_new_n397_));
  NOi21      g375(.An(i_2_), .B(i_12_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n398_), .B(new_new_n397_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(new_new_n396_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n145_), .B(i_9_), .Y(new_new_n401_));
  NO2        g379(.A(new_new_n401_), .B(i_4_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n400_), .B(new_new_n402_), .Y(new_new_n403_));
  NAi21      g381(.An(i_9_), .B(i_4_), .Y(new_new_n404_));
  OR2        g382(.A(i_13_), .B(i_10_), .Y(new_new_n405_));
  NO3        g383(.A(new_new_n405_), .B(new_new_n120_), .C(new_new_n404_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n175_), .B(new_new_n126_), .Y(new_new_n407_));
  OR2        g385(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n104_), .B(new_new_n25_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n275_), .B(new_new_n409_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n268_), .B(new_new_n211_), .Y(new_new_n411_));
  OAI220     g389(.A0(new_new_n411_), .A1(new_new_n408_), .B0(new_new_n410_), .B1(new_new_n327_), .Y(new_new_n412_));
  INV        g390(.A(new_new_n412_), .Y(new_new_n413_));
  AOI210     g391(.A0(new_new_n413_), .A1(new_new_n403_), .B0(new_new_n26_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n311_), .B(new_new_n310_), .Y(new_new_n415_));
  AOI220     g393(.A0(new_new_n289_), .A1(new_new_n279_), .B0(new_new_n283_), .B1(new_new_n302_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n416_), .B(new_new_n172_), .Y(new_new_n417_));
  NO2        g395(.A(new_new_n184_), .B(new_new_n86_), .Y(new_new_n418_));
  AOI220     g396(.A0(new_new_n418_), .A1(new_new_n288_), .B0(new_new_n270_), .B1(new_new_n211_), .Y(new_new_n419_));
  NO2        g397(.A(new_new_n419_), .B(new_new_n277_), .Y(new_new_n420_));
  NO3        g398(.A(new_new_n420_), .B(new_new_n417_), .C(new_new_n415_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n196_), .B(new_new_n99_), .Y(new_new_n422_));
  NA3        g400(.A(new_new_n313_), .B(new_new_n166_), .C(new_new_n86_), .Y(new_new_n423_));
  AOI210     g401(.A0(new_new_n423_), .A1(new_new_n422_), .B0(new_new_n312_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n193_), .B(i_10_), .Y(new_new_n425_));
  NA3        g403(.A(new_new_n249_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n289_), .B(new_new_n229_), .Y(new_new_n427_));
  OAI220     g405(.A0(new_new_n427_), .A1(new_new_n184_), .B0(new_new_n426_), .B1(new_new_n425_), .Y(new_new_n428_));
  NO2        g406(.A(i_3_), .B(new_new_n48_), .Y(new_new_n429_));
  NA3        g407(.A(new_new_n325_), .B(new_new_n324_), .C(new_new_n429_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n304_), .B(new_new_n309_), .Y(new_new_n431_));
  OAI210     g409(.A0(new_new_n431_), .A1(new_new_n190_), .B0(new_new_n430_), .Y(new_new_n432_));
  NO3        g410(.A(new_new_n432_), .B(new_new_n428_), .C(new_new_n424_), .Y(new_new_n433_));
  AOI210     g411(.A0(new_new_n433_), .A1(new_new_n421_), .B0(new_new_n264_), .Y(new_new_n434_));
  NO4        g412(.A(new_new_n434_), .B(new_new_n414_), .C(new_new_n392_), .D(new_new_n371_), .Y(new_new_n435_));
  NO2        g413(.A(new_new_n63_), .B(i_4_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n73_), .B(i_13_), .Y(new_new_n437_));
  NA3        g415(.A(new_new_n437_), .B(new_new_n436_), .C(i_2_), .Y(new_new_n438_));
  NO2        g416(.A(i_10_), .B(i_9_), .Y(new_new_n439_));
  NAi21      g417(.An(i_12_), .B(i_8_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n440_), .B(i_3_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n441_), .B(new_new_n439_), .Y(new_new_n442_));
  NO2        g420(.A(new_new_n46_), .B(i_4_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n443_), .B(new_new_n107_), .Y(new_new_n444_));
  OAI220     g422(.A0(new_new_n444_), .A1(new_new_n205_), .B0(new_new_n442_), .B1(new_new_n438_), .Y(new_new_n445_));
  NO3        g423(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n446_));
  NA2        g424(.A(new_new_n260_), .B(new_new_n100_), .Y(new_new_n447_));
  NA2        g425(.A(new_new_n447_), .B(new_new_n446_), .Y(new_new_n448_));
  NA2        g426(.A(i_8_), .B(i_9_), .Y(new_new_n449_));
  AOI210     g427(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n450_));
  OR2        g428(.A(new_new_n450_), .B(new_new_n449_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n275_), .B(new_new_n206_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n452_), .B(new_new_n451_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n243_), .B(new_new_n297_), .Y(new_new_n454_));
  NO3        g432(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n455_));
  INV        g433(.A(new_new_n455_), .Y(new_new_n456_));
  NA3        g434(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n457_));
  NA4        g435(.A(new_new_n148_), .B(new_new_n119_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n458_));
  OAI220     g436(.A0(new_new_n458_), .A1(new_new_n457_), .B0(new_new_n456_), .B1(new_new_n454_), .Y(new_new_n459_));
  NO3        g437(.A(new_new_n459_), .B(new_new_n453_), .C(new_new_n445_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n99_), .B(i_13_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n418_), .B(new_new_n372_), .Y(new_new_n462_));
  NO2        g440(.A(i_2_), .B(i_13_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n462_), .B(new_new_n461_), .Y(new_new_n464_));
  NO3        g442(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n465_));
  NO2        g443(.A(i_6_), .B(i_7_), .Y(new_new_n466_));
  NO2        g444(.A(i_11_), .B(i_1_), .Y(new_new_n467_));
  NOi21      g445(.An(i_2_), .B(i_7_), .Y(new_new_n468_));
  NO2        g446(.A(i_3_), .B(new_new_n193_), .Y(new_new_n469_));
  NO2        g447(.A(i_6_), .B(i_10_), .Y(new_new_n470_));
  NA4        g448(.A(new_new_n470_), .B(new_new_n301_), .C(new_new_n469_), .D(new_new_n231_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n471_), .B(new_new_n158_), .Y(new_new_n472_));
  NA3        g450(.A(new_new_n240_), .B(new_new_n174_), .C(new_new_n135_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n160_), .B(i_3_), .Y(new_new_n475_));
  NAi31      g453(.An(new_new_n474_), .B(new_new_n475_), .C(new_new_n223_), .Y(new_new_n476_));
  NA3        g454(.A(new_new_n385_), .B(new_new_n181_), .C(new_new_n152_), .Y(new_new_n477_));
  NA3        g455(.A(new_new_n477_), .B(new_new_n476_), .C(new_new_n473_), .Y(new_new_n478_));
  NO3        g456(.A(new_new_n478_), .B(new_new_n472_), .C(new_new_n464_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n446_), .B(new_new_n373_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n455_), .B(new_new_n380_), .Y(new_new_n481_));
  NAi21      g459(.An(new_new_n216_), .B(new_new_n390_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n325_), .B(new_new_n217_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n26_), .B(i_5_), .Y(new_new_n484_));
  NO2        g462(.A(i_0_), .B(new_new_n86_), .Y(new_new_n485_));
  NA3        g463(.A(new_new_n485_), .B(new_new_n484_), .C(new_new_n145_), .Y(new_new_n486_));
  OR3        g464(.A(new_new_n294_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n487_));
  OAI220     g465(.A0(new_new_n487_), .A1(new_new_n486_), .B0(new_new_n483_), .B1(new_new_n482_), .Y(new_new_n488_));
  NA2        g466(.A(new_new_n27_), .B(i_10_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n301_), .B(new_new_n233_), .Y(new_new_n490_));
  OAI220     g468(.A0(new_new_n490_), .A1(new_new_n426_), .B0(new_new_n489_), .B1(new_new_n461_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n491_), .B(new_new_n488_), .Y(new_new_n492_));
  NA3        g470(.A(new_new_n492_), .B(new_new_n479_), .C(new_new_n460_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n125_), .B(new_new_n115_), .Y(new_new_n494_));
  AN2        g472(.A(new_new_n494_), .B(new_new_n446_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n495_), .B(new_new_n298_), .Y(new_new_n496_));
  NA4        g474(.A(new_new_n437_), .B(new_new_n436_), .C(new_new_n203_), .D(i_2_), .Y(new_new_n497_));
  INV        g475(.A(new_new_n497_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n373_), .B(new_new_n222_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n342_), .B(new_new_n73_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n360_), .B(new_new_n352_), .Y(new_new_n501_));
  OR2        g479(.A(new_new_n499_), .B(new_new_n501_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n36_), .B(i_8_), .Y(new_new_n503_));
  AOI210     g481(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n406_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n504_), .B(new_new_n502_), .Y(new_new_n505_));
  AOI210     g483(.A0(new_new_n498_), .A1(new_new_n204_), .B0(new_new_n505_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n249_), .B(new_new_n64_), .Y(new_new_n507_));
  OAI210     g485(.A0(i_8_), .A1(new_new_n507_), .B0(new_new_n137_), .Y(new_new_n508_));
  AOI210     g486(.A0(new_new_n194_), .A1(i_9_), .B0(new_new_n259_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n509_), .B(new_new_n199_), .Y(new_new_n510_));
  OR2        g488(.A(new_new_n184_), .B(i_4_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n511_), .B(new_new_n86_), .Y(new_new_n512_));
  AOI220     g490(.A0(new_new_n512_), .A1(new_new_n510_), .B0(new_new_n508_), .B1(new_new_n407_), .Y(new_new_n513_));
  NA3        g491(.A(new_new_n513_), .B(new_new_n506_), .C(new_new_n496_), .Y(new_new_n514_));
  NO2        g492(.A(i_12_), .B(new_new_n193_), .Y(new_new_n515_));
  NA2        g493(.A(new_new_n515_), .B(new_new_n222_), .Y(new_new_n516_));
  NO2        g494(.A(i_8_), .B(i_7_), .Y(new_new_n517_));
  OAI210     g495(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n518_), .B(new_new_n221_), .Y(new_new_n519_));
  AOI220     g497(.A0(new_new_n313_), .A1(new_new_n40_), .B0(new_new_n229_), .B1(new_new_n208_), .Y(new_new_n520_));
  OAI220     g498(.A0(new_new_n520_), .A1(new_new_n511_), .B0(new_new_n519_), .B1(new_new_n237_), .Y(new_new_n521_));
  NA2        g499(.A(new_new_n44_), .B(i_10_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n522_), .B(i_6_), .Y(new_new_n523_));
  NA3        g501(.A(new_new_n523_), .B(new_new_n521_), .C(new_new_n517_), .Y(new_new_n524_));
  AOI220     g502(.A0(new_new_n418_), .A1(new_new_n313_), .B0(new_new_n241_), .B1(new_new_n239_), .Y(new_new_n525_));
  OAI220     g503(.A0(new_new_n525_), .A1(new_new_n256_), .B0(new_new_n461_), .B1(new_new_n136_), .Y(new_new_n526_));
  NA2        g504(.A(new_new_n526_), .B(new_new_n259_), .Y(new_new_n527_));
  NA3        g505(.A(new_new_n296_), .B(new_new_n177_), .C(new_new_n99_), .Y(new_new_n528_));
  NO2        g506(.A(new_new_n219_), .B(new_new_n44_), .Y(new_new_n529_));
  NO2        g507(.A(new_new_n160_), .B(i_5_), .Y(new_new_n530_));
  NA3        g508(.A(new_new_n530_), .B(new_new_n393_), .C(new_new_n307_), .Y(new_new_n531_));
  OAI210     g509(.A0(new_new_n531_), .A1(new_new_n529_), .B0(new_new_n528_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n532_), .B(new_new_n455_), .Y(new_new_n533_));
  NA3        g511(.A(new_new_n533_), .B(new_new_n527_), .C(new_new_n524_), .Y(new_new_n534_));
  NA3        g512(.A(new_new_n217_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n535_));
  NA2        g513(.A(new_new_n275_), .B(new_new_n84_), .Y(new_new_n536_));
  AOI210     g514(.A0(new_new_n535_), .A1(new_new_n332_), .B0(new_new_n536_), .Y(new_new_n537_));
  NA2        g515(.A(new_new_n289_), .B(new_new_n279_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n538_), .B(new_new_n176_), .Y(new_new_n539_));
  NA2        g517(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n540_));
  NA2        g518(.A(new_new_n439_), .B(new_new_n219_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n540_), .B(new_new_n541_), .Y(new_new_n542_));
  AOI210     g520(.A0(new_new_n353_), .A1(new_new_n46_), .B0(new_new_n357_), .Y(new_new_n543_));
  NA2        g521(.A(i_0_), .B(new_new_n48_), .Y(new_new_n544_));
  NA3        g522(.A(new_new_n515_), .B(new_new_n266_), .C(new_new_n544_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n543_), .B(new_new_n545_), .Y(new_new_n546_));
  NO4        g524(.A(new_new_n546_), .B(new_new_n542_), .C(new_new_n539_), .D(new_new_n537_), .Y(new_new_n547_));
  NO4        g525(.A(new_new_n244_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n548_));
  NO3        g526(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n405_), .B(i_1_), .Y(new_new_n550_));
  NOi31      g528(.An(new_new_n550_), .B(new_new_n447_), .C(new_new_n73_), .Y(new_new_n551_));
  AN4        g529(.A(new_new_n551_), .B(new_new_n402_), .C(new_new_n484_), .D(i_2_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n416_), .B(new_new_n180_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n553_), .B(new_new_n552_), .Y(new_new_n554_));
  NOi21      g532(.An(i_10_), .B(i_6_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n556_));
  NO2        g534(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n557_));
  NA2        g535(.A(new_new_n304_), .B(new_new_n167_), .Y(new_new_n558_));
  AOI220     g536(.A0(new_new_n558_), .A1(new_new_n427_), .B0(new_new_n185_), .B1(new_new_n183_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n198_), .B(new_new_n37_), .Y(new_new_n560_));
  NOi31      g538(.An(new_new_n149_), .B(new_new_n560_), .C(new_new_n320_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n561_), .B(new_new_n559_), .Y(new_new_n562_));
  NO2        g540(.A(new_new_n500_), .B(new_new_n368_), .Y(new_new_n563_));
  INV        g541(.A(new_new_n307_), .Y(new_new_n564_));
  NO2        g542(.A(i_12_), .B(new_new_n86_), .Y(new_new_n565_));
  OR2        g543(.A(i_2_), .B(i_5_), .Y(new_new_n566_));
  OR2        g544(.A(new_new_n566_), .B(new_new_n397_), .Y(new_new_n567_));
  AOI210     g545(.A0(new_new_n362_), .A1(new_new_n239_), .B0(new_new_n198_), .Y(new_new_n568_));
  AOI210     g546(.A0(new_new_n568_), .A1(new_new_n567_), .B0(new_new_n482_), .Y(new_new_n569_));
  NO2        g547(.A(new_new_n569_), .B(new_new_n563_), .Y(new_new_n570_));
  NA4        g548(.A(new_new_n570_), .B(new_new_n562_), .C(new_new_n554_), .D(new_new_n547_), .Y(new_new_n571_));
  NO4        g549(.A(new_new_n571_), .B(new_new_n534_), .C(new_new_n514_), .D(new_new_n493_), .Y(new_new_n572_));
  NA4        g550(.A(new_new_n572_), .B(new_new_n435_), .C(new_new_n341_), .D(new_new_n300_), .Y(ori7));
  NO2        g551(.A(new_new_n95_), .B(new_new_n54_), .Y(new_new_n574_));
  NO2        g552(.A(new_new_n111_), .B(new_new_n92_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n374_), .B(new_new_n575_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n470_), .B(new_new_n84_), .Y(new_new_n577_));
  NA2        g555(.A(i_11_), .B(new_new_n193_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n147_), .B(new_new_n578_), .Y(new_new_n579_));
  OAI210     g557(.A0(new_new_n579_), .A1(new_new_n577_), .B0(new_new_n576_), .Y(new_new_n580_));
  NA3        g558(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n231_), .B(i_4_), .Y(new_new_n582_));
  NA2        g560(.A(new_new_n582_), .B(i_8_), .Y(new_new_n583_));
  NO2        g561(.A(new_new_n108_), .B(new_new_n581_), .Y(new_new_n584_));
  NA2        g562(.A(i_2_), .B(new_new_n86_), .Y(new_new_n585_));
  OAI210     g563(.A0(new_new_n89_), .A1(new_new_n203_), .B0(new_new_n204_), .Y(new_new_n586_));
  NO2        g564(.A(i_7_), .B(new_new_n37_), .Y(new_new_n587_));
  NA2        g565(.A(i_4_), .B(i_8_), .Y(new_new_n588_));
  AOI210     g566(.A0(new_new_n588_), .A1(new_new_n296_), .B0(new_new_n587_), .Y(new_new_n589_));
  OAI220     g567(.A0(new_new_n589_), .A1(new_new_n585_), .B0(new_new_n586_), .B1(i_13_), .Y(new_new_n590_));
  NO4        g568(.A(new_new_n590_), .B(new_new_n584_), .C(new_new_n580_), .D(new_new_n574_), .Y(new_new_n591_));
  AOI210     g569(.A0(new_new_n131_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n592_));
  AOI210     g570(.A0(new_new_n592_), .A1(new_new_n231_), .B0(new_new_n164_), .Y(new_new_n593_));
  OR2        g571(.A(i_6_), .B(i_10_), .Y(new_new_n594_));
  NO2        g572(.A(new_new_n594_), .B(new_new_n23_), .Y(new_new_n595_));
  OR3        g573(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n596_));
  INV        g574(.A(new_new_n200_), .Y(new_new_n597_));
  INV        g575(.A(new_new_n595_), .Y(new_new_n598_));
  OA220      g576(.A0(new_new_n598_), .A1(new_new_n564_), .B0(new_new_n593_), .B1(new_new_n261_), .Y(new_new_n599_));
  AOI210     g577(.A0(new_new_n599_), .A1(new_new_n591_), .B0(new_new_n63_), .Y(new_new_n600_));
  NOi21      g578(.An(i_11_), .B(i_7_), .Y(new_new_n601_));
  AO210      g579(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n602_), .B(new_new_n601_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n603_), .B(new_new_n208_), .Y(new_new_n604_));
  NA3        g582(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n605_));
  NAi31      g583(.An(new_new_n605_), .B(new_new_n215_), .C(i_11_), .Y(new_new_n606_));
  AOI210     g584(.A0(new_new_n606_), .A1(new_new_n604_), .B0(new_new_n63_), .Y(new_new_n607_));
  NA2        g585(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n608_));
  AO210      g586(.A0(new_new_n608_), .A1(new_new_n368_), .B0(new_new_n41_), .Y(new_new_n609_));
  NO3        g587(.A(new_new_n251_), .B(new_new_n209_), .C(new_new_n578_), .Y(new_new_n610_));
  OAI210     g588(.A0(new_new_n610_), .A1(new_new_n223_), .B0(new_new_n63_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n398_), .B(new_new_n31_), .Y(new_new_n612_));
  OR2        g590(.A(new_new_n209_), .B(new_new_n111_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n613_), .B(new_new_n612_), .Y(new_new_n614_));
  NO2        g592(.A(new_new_n63_), .B(i_9_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n615_), .B(i_4_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n616_), .B(new_new_n614_), .Y(new_new_n617_));
  NO2        g595(.A(i_1_), .B(i_12_), .Y(new_new_n618_));
  NA3        g596(.A(new_new_n618_), .B(new_new_n113_), .C(new_new_n24_), .Y(new_new_n619_));
  BUFFER     g597(.A(new_new_n619_), .Y(new_new_n620_));
  NA4        g598(.A(new_new_n620_), .B(new_new_n617_), .C(new_new_n611_), .D(new_new_n609_), .Y(new_new_n621_));
  OAI210     g599(.A0(new_new_n621_), .A1(new_new_n607_), .B0(i_6_), .Y(new_new_n622_));
  NO2        g600(.A(new_new_n605_), .B(new_new_n111_), .Y(new_new_n623_));
  NA2        g601(.A(new_new_n623_), .B(new_new_n565_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n231_), .B(new_new_n86_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(i_11_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n624_), .B(new_new_n448_), .Y(new_new_n627_));
  NO4        g605(.A(new_new_n215_), .B(new_new_n131_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n628_));
  NA2        g606(.A(new_new_n628_), .B(new_new_n615_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n231_), .B(i_6_), .Y(new_new_n630_));
  NO3        g608(.A(new_new_n594_), .B(new_new_n227_), .C(new_new_n23_), .Y(new_new_n631_));
  AOI210     g609(.A0(i_1_), .A1(new_new_n252_), .B0(new_new_n631_), .Y(new_new_n632_));
  OAI210     g610(.A0(new_new_n632_), .A1(new_new_n44_), .B0(new_new_n629_), .Y(new_new_n633_));
  INV        g611(.A(i_2_), .Y(new_new_n634_));
  NA2        g612(.A(new_new_n141_), .B(i_9_), .Y(new_new_n635_));
  NA3        g613(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n46_), .B(i_1_), .Y(new_new_n637_));
  NA3        g615(.A(new_new_n637_), .B(new_new_n260_), .C(new_new_n44_), .Y(new_new_n638_));
  OAI220     g616(.A0(new_new_n638_), .A1(new_new_n636_), .B0(new_new_n635_), .B1(new_new_n634_), .Y(new_new_n639_));
  NA3        g617(.A(new_new_n615_), .B(new_new_n307_), .C(i_6_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n640_), .B(new_new_n23_), .Y(new_new_n641_));
  AOI210     g619(.A0(new_new_n467_), .A1(new_new_n409_), .B0(new_new_n236_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n642_), .B(new_new_n585_), .Y(new_new_n643_));
  NA2        g621(.A(new_new_n637_), .B(new_new_n260_), .Y(new_new_n644_));
  NO2        g622(.A(i_11_), .B(new_new_n37_), .Y(new_new_n645_));
  NA2        g623(.A(new_new_n645_), .B(new_new_n24_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n646_), .B(new_new_n644_), .Y(new_new_n647_));
  OR4        g625(.A(new_new_n647_), .B(new_new_n643_), .C(new_new_n641_), .D(new_new_n639_), .Y(new_new_n648_));
  NO3        g626(.A(new_new_n648_), .B(new_new_n633_), .C(new_new_n627_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n231_), .B(new_new_n104_), .Y(new_new_n650_));
  NO2        g628(.A(new_new_n650_), .B(new_new_n601_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n651_), .B(i_1_), .Y(new_new_n652_));
  NO2        g630(.A(new_new_n652_), .B(new_new_n596_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n404_), .B(new_new_n86_), .Y(new_new_n654_));
  NA2        g632(.A(new_new_n653_), .B(new_new_n46_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n227_), .B(new_new_n44_), .Y(new_new_n656_));
  NO3        g634(.A(new_new_n656_), .B(new_new_n298_), .C(new_new_n232_), .Y(new_new_n657_));
  NO2        g635(.A(new_new_n120_), .B(new_new_n37_), .Y(new_new_n658_));
  NO2        g636(.A(new_new_n658_), .B(i_6_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n86_), .B(i_9_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n660_), .B(new_new_n63_), .Y(new_new_n661_));
  NO2        g639(.A(new_new_n661_), .B(new_new_n618_), .Y(new_new_n662_));
  NO4        g640(.A(new_new_n662_), .B(new_new_n659_), .C(new_new_n657_), .D(i_4_), .Y(new_new_n663_));
  NA2        g641(.A(i_1_), .B(i_3_), .Y(new_new_n664_));
  INV        g642(.A(new_new_n663_), .Y(new_new_n665_));
  NA4        g643(.A(new_new_n665_), .B(new_new_n655_), .C(new_new_n649_), .D(new_new_n622_), .Y(new_new_n666_));
  NO3        g644(.A(new_new_n468_), .B(new_new_n588_), .C(new_new_n86_), .Y(new_new_n667_));
  NA2        g645(.A(new_new_n667_), .B(new_new_n25_), .Y(new_new_n668_));
  NA3        g646(.A(new_new_n164_), .B(new_new_n84_), .C(new_new_n86_), .Y(new_new_n669_));
  NA2        g647(.A(new_new_n669_), .B(new_new_n668_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n670_), .B(i_1_), .Y(new_new_n671_));
  AOI210     g649(.A0(new_new_n260_), .A1(new_new_n100_), .B0(i_1_), .Y(new_new_n672_));
  NO2        g650(.A(new_new_n358_), .B(i_2_), .Y(new_new_n673_));
  NA2        g651(.A(new_new_n673_), .B(new_new_n672_), .Y(new_new_n674_));
  OAI210     g652(.A0(new_new_n640_), .A1(new_new_n440_), .B0(new_new_n674_), .Y(new_new_n675_));
  INV        g653(.A(new_new_n675_), .Y(new_new_n676_));
  AOI210     g654(.A0(new_new_n676_), .A1(new_new_n671_), .B0(i_13_), .Y(new_new_n677_));
  OR2        g655(.A(i_11_), .B(i_7_), .Y(new_new_n678_));
  NA3        g656(.A(new_new_n678_), .B(new_new_n109_), .C(new_new_n141_), .Y(new_new_n679_));
  AOI220     g657(.A0(new_new_n463_), .A1(new_new_n164_), .B0(new_new_n443_), .B1(new_new_n141_), .Y(new_new_n680_));
  OAI210     g658(.A0(new_new_n680_), .A1(new_new_n44_), .B0(new_new_n679_), .Y(new_new_n681_));
  AOI210     g659(.A0(new_new_n636_), .A1(new_new_n54_), .B0(i_12_), .Y(new_new_n682_));
  NO2        g660(.A(new_new_n468_), .B(new_new_n24_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n683_), .B(new_new_n654_), .Y(new_new_n684_));
  OAI220     g662(.A0(new_new_n684_), .A1(new_new_n41_), .B0(new_new_n1009_), .B1(new_new_n95_), .Y(new_new_n685_));
  AOI210     g663(.A0(new_new_n681_), .A1(new_new_n322_), .B0(new_new_n685_), .Y(new_new_n686_));
  INV        g664(.A(new_new_n118_), .Y(new_new_n687_));
  AOI220     g665(.A0(new_new_n687_), .A1(new_new_n72_), .B0(new_new_n376_), .B1(new_new_n637_), .Y(new_new_n688_));
  NO2        g666(.A(new_new_n688_), .B(new_new_n237_), .Y(new_new_n689_));
  AOI210     g667(.A0(new_new_n440_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n690_));
  NOi31      g668(.An(new_new_n690_), .B(new_new_n577_), .C(new_new_n44_), .Y(new_new_n691_));
  NA2        g669(.A(new_new_n130_), .B(i_13_), .Y(new_new_n692_));
  NO2        g670(.A(new_new_n636_), .B(new_new_n118_), .Y(new_new_n693_));
  INV        g671(.A(new_new_n693_), .Y(new_new_n694_));
  OAI220     g672(.A0(new_new_n694_), .A1(new_new_n71_), .B0(new_new_n692_), .B1(new_new_n672_), .Y(new_new_n695_));
  NO3        g673(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n104_), .Y(new_new_n696_));
  NA2        g674(.A(new_new_n26_), .B(new_new_n193_), .Y(new_new_n697_));
  NA2        g675(.A(new_new_n697_), .B(i_7_), .Y(new_new_n698_));
  NO3        g676(.A(new_new_n468_), .B(new_new_n231_), .C(new_new_n86_), .Y(new_new_n699_));
  AOI210     g677(.A0(new_new_n699_), .A1(new_new_n698_), .B0(new_new_n696_), .Y(new_new_n700_));
  AOI220     g678(.A0(new_new_n376_), .A1(new_new_n637_), .B0(new_new_n94_), .B1(new_new_n105_), .Y(new_new_n701_));
  OAI220     g679(.A0(new_new_n701_), .A1(new_new_n583_), .B0(new_new_n700_), .B1(new_new_n597_), .Y(new_new_n702_));
  NO4        g680(.A(new_new_n702_), .B(new_new_n695_), .C(new_new_n691_), .D(new_new_n689_), .Y(new_new_n703_));
  OR2        g681(.A(i_11_), .B(i_6_), .Y(new_new_n704_));
  NA3        g682(.A(new_new_n582_), .B(new_new_n697_), .C(i_7_), .Y(new_new_n705_));
  AOI210     g683(.A0(new_new_n705_), .A1(new_new_n694_), .B0(new_new_n704_), .Y(new_new_n706_));
  NA3        g684(.A(new_new_n398_), .B(new_new_n587_), .C(new_new_n100_), .Y(new_new_n707_));
  NA2        g685(.A(new_new_n626_), .B(i_13_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n105_), .B(new_new_n697_), .Y(new_new_n709_));
  NAi21      g687(.An(i_11_), .B(i_12_), .Y(new_new_n710_));
  NOi41      g688(.An(new_new_n114_), .B(new_new_n710_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n711_), .B(new_new_n709_), .Y(new_new_n712_));
  NA3        g690(.A(new_new_n712_), .B(new_new_n708_), .C(new_new_n707_), .Y(new_new_n713_));
  OAI210     g691(.A0(new_new_n713_), .A1(new_new_n706_), .B0(new_new_n63_), .Y(new_new_n714_));
  NO2        g692(.A(i_2_), .B(i_12_), .Y(new_new_n715_));
  NA2        g693(.A(new_new_n357_), .B(new_new_n715_), .Y(new_new_n716_));
  NA2        g694(.A(i_8_), .B(new_new_n25_), .Y(new_new_n717_));
  NO3        g695(.A(new_new_n717_), .B(new_new_n374_), .C(new_new_n582_), .Y(new_new_n718_));
  OAI210     g696(.A0(new_new_n718_), .A1(new_new_n359_), .B0(new_new_n357_), .Y(new_new_n719_));
  NO2        g697(.A(new_new_n131_), .B(i_2_), .Y(new_new_n720_));
  NA2        g698(.A(new_new_n720_), .B(new_new_n618_), .Y(new_new_n721_));
  NA3        g699(.A(new_new_n721_), .B(new_new_n719_), .C(new_new_n716_), .Y(new_new_n722_));
  NA3        g700(.A(new_new_n722_), .B(new_new_n45_), .C(new_new_n222_), .Y(new_new_n723_));
  NA4        g701(.A(new_new_n723_), .B(new_new_n714_), .C(new_new_n703_), .D(new_new_n686_), .Y(new_new_n724_));
  OR4        g702(.A(new_new_n724_), .B(new_new_n677_), .C(new_new_n666_), .D(new_new_n600_), .Y(ori5));
  NA2        g703(.A(new_new_n651_), .B(new_new_n263_), .Y(new_new_n726_));
  AN2        g704(.A(new_new_n24_), .B(i_10_), .Y(new_new_n727_));
  NA3        g705(.A(new_new_n727_), .B(new_new_n715_), .C(new_new_n111_), .Y(new_new_n728_));
  NO2        g706(.A(new_new_n583_), .B(i_11_), .Y(new_new_n729_));
  NA2        g707(.A(new_new_n89_), .B(new_new_n729_), .Y(new_new_n730_));
  NA3        g708(.A(new_new_n730_), .B(new_new_n728_), .C(new_new_n726_), .Y(new_new_n731_));
  NO3        g709(.A(i_11_), .B(new_new_n231_), .C(i_13_), .Y(new_new_n732_));
  NO2        g710(.A(new_new_n127_), .B(new_new_n23_), .Y(new_new_n733_));
  NA2        g711(.A(i_12_), .B(i_8_), .Y(new_new_n734_));
  OAI210     g712(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n734_), .Y(new_new_n735_));
  INV        g713(.A(new_new_n439_), .Y(new_new_n736_));
  AOI220     g714(.A0(new_new_n307_), .A1(new_new_n557_), .B0(new_new_n735_), .B1(new_new_n733_), .Y(new_new_n737_));
  INV        g715(.A(new_new_n737_), .Y(new_new_n738_));
  NO2        g716(.A(new_new_n738_), .B(new_new_n731_), .Y(new_new_n739_));
  INV        g717(.A(new_new_n174_), .Y(new_new_n740_));
  INV        g718(.A(new_new_n240_), .Y(new_new_n741_));
  OAI210     g719(.A0(new_new_n673_), .A1(new_new_n441_), .B0(new_new_n114_), .Y(new_new_n742_));
  AOI210     g720(.A0(new_new_n742_), .A1(new_new_n741_), .B0(new_new_n740_), .Y(new_new_n743_));
  NO2        g721(.A(new_new_n449_), .B(new_new_n26_), .Y(new_new_n744_));
  NO2        g722(.A(new_new_n744_), .B(new_new_n409_), .Y(new_new_n745_));
  NA2        g723(.A(new_new_n745_), .B(i_2_), .Y(new_new_n746_));
  INV        g724(.A(new_new_n746_), .Y(new_new_n747_));
  AOI210     g725(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n405_), .Y(new_new_n748_));
  AOI210     g726(.A0(new_new_n748_), .A1(new_new_n747_), .B0(new_new_n743_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n191_), .B(new_new_n128_), .Y(new_new_n750_));
  OAI210     g728(.A0(new_new_n750_), .A1(new_new_n733_), .B0(i_2_), .Y(new_new_n751_));
  INV        g729(.A(new_new_n175_), .Y(new_new_n752_));
  NO3        g730(.A(new_new_n602_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n753_));
  AOI210     g731(.A0(new_new_n752_), .A1(new_new_n89_), .B0(new_new_n753_), .Y(new_new_n754_));
  AOI210     g732(.A0(new_new_n754_), .A1(new_new_n751_), .B0(new_new_n193_), .Y(new_new_n755_));
  OA210      g733(.A0(new_new_n603_), .A1(new_new_n129_), .B0(i_13_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n200_), .B(new_new_n203_), .Y(new_new_n757_));
  NA2        g735(.A(new_new_n154_), .B(new_new_n578_), .Y(new_new_n758_));
  AOI210     g736(.A0(new_new_n758_), .A1(new_new_n757_), .B0(new_new_n362_), .Y(new_new_n759_));
  AOI210     g737(.A0(new_new_n209_), .A1(new_new_n151_), .B0(new_new_n503_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n760_), .B(new_new_n409_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n105_), .B(new_new_n44_), .Y(new_new_n762_));
  INV        g740(.A(new_new_n293_), .Y(new_new_n763_));
  NA4        g741(.A(new_new_n763_), .B(new_new_n296_), .C(new_new_n127_), .D(new_new_n42_), .Y(new_new_n764_));
  OAI210     g742(.A0(new_new_n764_), .A1(new_new_n762_), .B0(new_new_n761_), .Y(new_new_n765_));
  NO4        g743(.A(new_new_n765_), .B(new_new_n759_), .C(new_new_n756_), .D(new_new_n755_), .Y(new_new_n766_));
  NA2        g744(.A(new_new_n557_), .B(new_new_n28_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n732_), .B(new_new_n267_), .Y(new_new_n768_));
  NA2        g746(.A(new_new_n768_), .B(new_new_n767_), .Y(new_new_n769_));
  NO2        g747(.A(new_new_n62_), .B(i_12_), .Y(new_new_n770_));
  NO2        g748(.A(new_new_n770_), .B(new_new_n129_), .Y(new_new_n771_));
  NO2        g749(.A(new_new_n771_), .B(new_new_n578_), .Y(new_new_n772_));
  AOI220     g750(.A0(new_new_n772_), .A1(new_new_n36_), .B0(new_new_n769_), .B1(new_new_n46_), .Y(new_new_n773_));
  NA4        g751(.A(new_new_n773_), .B(new_new_n766_), .C(new_new_n749_), .D(new_new_n739_), .Y(ori6));
  NO3        g752(.A(i_9_), .B(new_new_n297_), .C(i_1_), .Y(new_new_n775_));
  NO2        g753(.A(new_new_n187_), .B(new_new_n142_), .Y(new_new_n776_));
  OAI210     g754(.A0(new_new_n776_), .A1(new_new_n775_), .B0(new_new_n720_), .Y(new_new_n777_));
  NA4        g755(.A(new_new_n380_), .B(new_new_n469_), .C(new_new_n71_), .D(new_new_n104_), .Y(new_new_n778_));
  INV        g756(.A(new_new_n778_), .Y(new_new_n779_));
  NO2        g757(.A(new_new_n218_), .B(new_new_n474_), .Y(new_new_n780_));
  NO2        g758(.A(new_new_n779_), .B(new_new_n317_), .Y(new_new_n781_));
  AO210      g759(.A0(new_new_n781_), .A1(new_new_n777_), .B0(i_12_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n565_), .B(new_new_n63_), .Y(new_new_n783_));
  BUFFER     g761(.A(new_new_n608_), .Y(new_new_n784_));
  NA2        g762(.A(new_new_n784_), .B(new_new_n783_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n785_), .B(new_new_n73_), .Y(new_new_n786_));
  INV        g764(.A(new_new_n316_), .Y(new_new_n787_));
  NA2        g765(.A(new_new_n75_), .B(new_new_n134_), .Y(new_new_n788_));
  INV        g766(.A(new_new_n127_), .Y(new_new_n789_));
  NA2        g767(.A(new_new_n789_), .B(new_new_n46_), .Y(new_new_n790_));
  AOI210     g768(.A0(new_new_n790_), .A1(new_new_n788_), .B0(new_new_n787_), .Y(new_new_n791_));
  NO3        g769(.A(new_new_n244_), .B(new_new_n135_), .C(i_9_), .Y(new_new_n792_));
  NA2        g770(.A(new_new_n792_), .B(new_new_n770_), .Y(new_new_n793_));
  AOI210     g771(.A0(new_new_n793_), .A1(new_new_n501_), .B0(new_new_n187_), .Y(new_new_n794_));
  NO2        g772(.A(new_new_n32_), .B(i_11_), .Y(new_new_n795_));
  NAi32      g773(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n796_));
  NO2        g774(.A(new_new_n704_), .B(new_new_n796_), .Y(new_new_n797_));
  OR3        g775(.A(new_new_n797_), .B(new_new_n794_), .C(new_new_n791_), .Y(new_new_n798_));
  NO2        g776(.A(new_new_n678_), .B(i_2_), .Y(new_new_n799_));
  NA2        g777(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n800_), .B(new_new_n397_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n801_), .B(new_new_n799_), .Y(new_new_n802_));
  AO220      g780(.A0(new_new_n346_), .A1(new_new_n336_), .B0(new_new_n388_), .B1(new_new_n578_), .Y(new_new_n803_));
  NA3        g781(.A(new_new_n803_), .B(new_new_n248_), .C(i_7_), .Y(new_new_n804_));
  OR2        g782(.A(new_new_n603_), .B(new_new_n441_), .Y(new_new_n805_));
  NA3        g783(.A(new_new_n805_), .B(new_new_n150_), .C(new_new_n69_), .Y(new_new_n806_));
  AO210      g784(.A0(new_new_n481_), .A1(new_new_n736_), .B0(new_new_n36_), .Y(new_new_n807_));
  NA4        g785(.A(new_new_n807_), .B(new_new_n806_), .C(new_new_n804_), .D(new_new_n802_), .Y(new_new_n808_));
  OAI210     g786(.A0(new_new_n625_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n809_));
  AOI220     g787(.A0(new_new_n809_), .A1(new_new_n549_), .B0(new_new_n780_), .B1(new_new_n698_), .Y(new_new_n810_));
  NA3        g788(.A(new_new_n362_), .B(new_new_n233_), .C(new_new_n150_), .Y(new_new_n811_));
  NA2        g789(.A(new_new_n388_), .B(new_new_n70_), .Y(new_new_n812_));
  NA4        g790(.A(new_new_n812_), .B(new_new_n811_), .C(new_new_n810_), .D(new_new_n586_), .Y(new_new_n813_));
  AOI210     g791(.A0(new_new_n441_), .A1(new_new_n439_), .B0(new_new_n548_), .Y(new_new_n814_));
  NO2        g792(.A(new_new_n594_), .B(new_new_n105_), .Y(new_new_n815_));
  OAI210     g793(.A0(new_new_n815_), .A1(new_new_n115_), .B0(new_new_n395_), .Y(new_new_n816_));
  NA2        g794(.A(new_new_n239_), .B(new_new_n46_), .Y(new_new_n817_));
  INV        g795(.A(new_new_n567_), .Y(new_new_n818_));
  NA3        g796(.A(new_new_n818_), .B(new_new_n316_), .C(i_7_), .Y(new_new_n819_));
  NA3        g797(.A(new_new_n819_), .B(new_new_n816_), .C(new_new_n814_), .Y(new_new_n820_));
  NO4        g798(.A(new_new_n820_), .B(new_new_n813_), .C(new_new_n808_), .D(new_new_n798_), .Y(new_new_n821_));
  NA4        g799(.A(new_new_n821_), .B(new_new_n786_), .C(new_new_n782_), .D(new_new_n370_), .Y(ori3));
  NA2        g800(.A(i_12_), .B(i_10_), .Y(new_new_n823_));
  NA2        g801(.A(i_6_), .B(i_7_), .Y(new_new_n824_));
  NO2        g802(.A(new_new_n824_), .B(i_0_), .Y(new_new_n825_));
  NO2        g803(.A(i_11_), .B(new_new_n231_), .Y(new_new_n826_));
  NA3        g804(.A(new_new_n811_), .B(new_new_n586_), .C(new_new_n361_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n827_), .B(new_new_n40_), .Y(new_new_n828_));
  NOi21      g806(.An(new_new_n99_), .B(new_new_n745_), .Y(new_new_n829_));
  NO3        g807(.A(new_new_n613_), .B(new_new_n449_), .C(new_new_n134_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n398_), .B(new_new_n45_), .Y(new_new_n831_));
  AN2        g809(.A(new_new_n447_), .B(new_new_n55_), .Y(new_new_n832_));
  NO3        g810(.A(new_new_n832_), .B(new_new_n830_), .C(new_new_n829_), .Y(new_new_n833_));
  AOI210     g811(.A0(new_new_n833_), .A1(new_new_n828_), .B0(new_new_n48_), .Y(new_new_n834_));
  NO4        g812(.A(new_new_n366_), .B(new_new_n373_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n187_), .B(new_new_n555_), .Y(new_new_n836_));
  NOi21      g814(.An(new_new_n836_), .B(new_new_n835_), .Y(new_new_n837_));
  NA2        g815(.A(new_new_n690_), .B(new_new_n660_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n323_), .B(new_new_n429_), .Y(new_new_n839_));
  OAI220     g817(.A0(new_new_n839_), .A1(new_new_n838_), .B0(new_new_n837_), .B1(new_new_n63_), .Y(new_new_n840_));
  NOi21      g818(.An(i_5_), .B(i_9_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n841_), .B(new_new_n437_), .Y(new_new_n842_));
  BUFFER     g820(.A(new_new_n260_), .Y(new_new_n843_));
  AOI210     g821(.A0(new_new_n843_), .A1(new_new_n467_), .B0(new_new_n667_), .Y(new_new_n844_));
  NO2        g822(.A(new_new_n844_), .B(new_new_n842_), .Y(new_new_n845_));
  NO3        g823(.A(new_new_n845_), .B(new_new_n840_), .C(new_new_n834_), .Y(new_new_n846_));
  NA2        g824(.A(new_new_n187_), .B(new_new_n24_), .Y(new_new_n847_));
  NO2        g825(.A(new_new_n658_), .B(new_new_n575_), .Y(new_new_n848_));
  NO2        g826(.A(new_new_n848_), .B(new_new_n847_), .Y(new_new_n849_));
  NA2        g827(.A(new_new_n301_), .B(new_new_n132_), .Y(new_new_n850_));
  NAi21      g828(.An(new_new_n165_), .B(new_new_n429_), .Y(new_new_n851_));
  OAI220     g829(.A0(new_new_n851_), .A1(new_new_n817_), .B0(new_new_n850_), .B1(new_new_n391_), .Y(new_new_n852_));
  NO2        g830(.A(new_new_n852_), .B(new_new_n849_), .Y(new_new_n853_));
  NA2        g831(.A(new_new_n556_), .B(i_0_), .Y(new_new_n854_));
  NO4        g832(.A(new_new_n566_), .B(new_new_n215_), .C(new_new_n405_), .D(new_new_n397_), .Y(new_new_n855_));
  NA2        g833(.A(new_new_n855_), .B(i_11_), .Y(new_new_n856_));
  INV        g834(.A(new_new_n466_), .Y(new_new_n857_));
  AN2        g835(.A(new_new_n99_), .B(new_new_n238_), .Y(new_new_n858_));
  NA2        g836(.A(new_new_n732_), .B(new_new_n317_), .Y(new_new_n859_));
  AOI210     g837(.A0(new_new_n470_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n860_));
  OAI220     g838(.A0(new_new_n860_), .A1(new_new_n859_), .B0(new_new_n646_), .B1(new_new_n519_), .Y(new_new_n861_));
  NO2        g839(.A(new_new_n246_), .B(new_new_n156_), .Y(new_new_n862_));
  NA2        g840(.A(i_0_), .B(i_10_), .Y(new_new_n863_));
  AN2        g841(.A(new_new_n862_), .B(i_6_), .Y(new_new_n864_));
  AOI220     g842(.A0(new_new_n323_), .A1(new_new_n101_), .B0(new_new_n187_), .B1(new_new_n84_), .Y(new_new_n865_));
  NA2        g843(.A(new_new_n550_), .B(i_4_), .Y(new_new_n866_));
  NA2        g844(.A(new_new_n189_), .B(new_new_n203_), .Y(new_new_n867_));
  OAI220     g845(.A0(new_new_n867_), .A1(new_new_n859_), .B0(new_new_n866_), .B1(new_new_n865_), .Y(new_new_n868_));
  NO4        g846(.A(new_new_n868_), .B(new_new_n864_), .C(new_new_n861_), .D(new_new_n858_), .Y(new_new_n869_));
  NA3        g847(.A(new_new_n869_), .B(new_new_n856_), .C(new_new_n853_), .Y(new_new_n870_));
  NO2        g848(.A(new_new_n106_), .B(new_new_n37_), .Y(new_new_n871_));
  NA2        g849(.A(i_11_), .B(i_9_), .Y(new_new_n872_));
  NO3        g850(.A(i_12_), .B(new_new_n872_), .C(new_new_n585_), .Y(new_new_n873_));
  AN2        g851(.A(new_new_n873_), .B(new_new_n871_), .Y(new_new_n874_));
  NO2        g852(.A(new_new_n48_), .B(i_7_), .Y(new_new_n875_));
  NA2        g853(.A(new_new_n385_), .B(new_new_n181_), .Y(new_new_n876_));
  NA2        g854(.A(new_new_n876_), .B(new_new_n163_), .Y(new_new_n877_));
  NO2        g855(.A(new_new_n872_), .B(new_new_n73_), .Y(new_new_n878_));
  NO2        g856(.A(new_new_n178_), .B(i_0_), .Y(new_new_n879_));
  INV        g857(.A(new_new_n879_), .Y(new_new_n880_));
  NA2        g858(.A(new_new_n466_), .B(new_new_n225_), .Y(new_new_n881_));
  INV        g859(.A(new_new_n394_), .Y(new_new_n882_));
  OAI220     g860(.A0(new_new_n882_), .A1(new_new_n842_), .B0(new_new_n881_), .B1(new_new_n880_), .Y(new_new_n883_));
  NO3        g861(.A(new_new_n883_), .B(new_new_n877_), .C(new_new_n874_), .Y(new_new_n884_));
  NA2        g862(.A(new_new_n645_), .B(new_new_n124_), .Y(new_new_n885_));
  NO2        g863(.A(i_6_), .B(new_new_n885_), .Y(new_new_n886_));
  AOI210     g864(.A0(new_new_n440_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n887_));
  NA2        g865(.A(new_new_n174_), .B(new_new_n106_), .Y(new_new_n888_));
  NOi32      g866(.An(new_new_n887_), .Bn(new_new_n189_), .C(new_new_n888_), .Y(new_new_n889_));
  NO2        g867(.A(new_new_n889_), .B(new_new_n886_), .Y(new_new_n890_));
  NOi21      g868(.An(i_7_), .B(i_5_), .Y(new_new_n891_));
  NOi31      g869(.An(new_new_n891_), .B(i_0_), .C(new_new_n710_), .Y(new_new_n892_));
  NA3        g870(.A(new_new_n892_), .B(new_new_n374_), .C(i_6_), .Y(new_new_n893_));
  OA210      g871(.A0(new_new_n888_), .A1(new_new_n501_), .B0(new_new_n893_), .Y(new_new_n894_));
  INV        g872(.A(new_new_n308_), .Y(new_new_n895_));
  NA3        g873(.A(new_new_n894_), .B(new_new_n890_), .C(new_new_n884_), .Y(new_new_n896_));
  NO2        g874(.A(new_new_n823_), .B(new_new_n307_), .Y(new_new_n897_));
  OA210      g875(.A0(new_new_n466_), .A1(new_new_n221_), .B0(new_new_n465_), .Y(new_new_n898_));
  NA2        g876(.A(new_new_n897_), .B(new_new_n878_), .Y(new_new_n899_));
  NA3        g877(.A(new_new_n465_), .B(new_new_n398_), .C(new_new_n45_), .Y(new_new_n900_));
  OAI210     g878(.A0(new_new_n851_), .A1(new_new_n857_), .B0(new_new_n900_), .Y(new_new_n901_));
  NA2        g879(.A(new_new_n901_), .B(new_new_n73_), .Y(new_new_n902_));
  NA3        g880(.A(new_new_n800_), .B(new_new_n372_), .C(new_new_n625_), .Y(new_new_n903_));
  NA2        g881(.A(new_new_n95_), .B(new_new_n44_), .Y(new_new_n904_));
  NO2        g882(.A(new_new_n75_), .B(new_new_n734_), .Y(new_new_n905_));
  AOI220     g883(.A0(new_new_n905_), .A1(new_new_n904_), .B0(new_new_n177_), .B1(new_new_n575_), .Y(new_new_n906_));
  AOI210     g884(.A0(new_new_n906_), .A1(new_new_n903_), .B0(new_new_n47_), .Y(new_new_n907_));
  NO3        g885(.A(new_new_n566_), .B(new_new_n344_), .C(new_new_n24_), .Y(new_new_n908_));
  AOI210     g886(.A0(new_new_n683_), .A1(new_new_n530_), .B0(new_new_n908_), .Y(new_new_n909_));
  NO2        g887(.A(new_new_n581_), .B(new_new_n108_), .Y(new_new_n910_));
  NA2        g888(.A(new_new_n910_), .B(i_0_), .Y(new_new_n911_));
  OAI220     g889(.A0(new_new_n911_), .A1(new_new_n86_), .B0(new_new_n909_), .B1(new_new_n175_), .Y(new_new_n912_));
  NO3        g890(.A(new_new_n912_), .B(new_new_n907_), .C(new_new_n505_), .Y(new_new_n913_));
  NA3        g891(.A(new_new_n913_), .B(new_new_n902_), .C(new_new_n899_), .Y(new_new_n914_));
  NO3        g892(.A(new_new_n914_), .B(new_new_n896_), .C(new_new_n870_), .Y(new_new_n915_));
  NO2        g893(.A(i_0_), .B(new_new_n710_), .Y(new_new_n916_));
  NA2        g894(.A(new_new_n73_), .B(new_new_n44_), .Y(new_new_n917_));
  NO2        g895(.A(new_new_n783_), .B(new_new_n888_), .Y(new_new_n918_));
  INV        g896(.A(new_new_n918_), .Y(new_new_n919_));
  NA3        g897(.A(new_new_n825_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n920_));
  NA2        g898(.A(new_new_n826_), .B(i_9_), .Y(new_new_n921_));
  AOI210     g899(.A0(new_new_n920_), .A1(new_new_n486_), .B0(new_new_n921_), .Y(new_new_n922_));
  OAI210     g900(.A0(new_new_n239_), .A1(i_9_), .B0(new_new_n224_), .Y(new_new_n923_));
  AOI210     g901(.A0(new_new_n923_), .A1(new_new_n854_), .B0(new_new_n156_), .Y(new_new_n924_));
  NO2        g902(.A(new_new_n924_), .B(new_new_n922_), .Y(new_new_n925_));
  NA2        g903(.A(new_new_n925_), .B(new_new_n919_), .Y(new_new_n926_));
  NO3        g904(.A(new_new_n863_), .B(new_new_n841_), .C(new_new_n191_), .Y(new_new_n927_));
  AOI220     g905(.A0(new_new_n927_), .A1(i_11_), .B0(new_new_n551_), .B1(new_new_n75_), .Y(new_new_n928_));
  NO3        g906(.A(new_new_n210_), .B(new_new_n373_), .C(i_0_), .Y(new_new_n929_));
  OAI210     g907(.A0(new_new_n929_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n930_));
  INV        g908(.A(new_new_n217_), .Y(new_new_n931_));
  OAI220     g909(.A0(new_new_n516_), .A1(new_new_n142_), .B0(new_new_n630_), .B1(new_new_n597_), .Y(new_new_n932_));
  NA3        g910(.A(new_new_n932_), .B(new_new_n389_), .C(new_new_n931_), .Y(new_new_n933_));
  NA3        g911(.A(new_new_n933_), .B(new_new_n930_), .C(new_new_n928_), .Y(new_new_n934_));
  NO2        g912(.A(new_new_n237_), .B(new_new_n95_), .Y(new_new_n935_));
  AOI210     g913(.A0(new_new_n935_), .A1(new_new_n916_), .B0(new_new_n112_), .Y(new_new_n936_));
  AOI220     g914(.A0(new_new_n891_), .A1(new_new_n475_), .B0(new_new_n825_), .B1(new_new_n166_), .Y(new_new_n937_));
  NA2        g915(.A(new_new_n336_), .B(new_new_n179_), .Y(new_new_n938_));
  OA220      g916(.A0(new_new_n938_), .A1(new_new_n937_), .B0(new_new_n936_), .B1(i_5_), .Y(new_new_n939_));
  AOI210     g917(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n178_), .Y(new_new_n940_));
  NA2        g918(.A(new_new_n940_), .B(new_new_n898_), .Y(new_new_n941_));
  NA3        g919(.A(new_new_n595_), .B(new_new_n187_), .C(new_new_n84_), .Y(new_new_n942_));
  NA2        g920(.A(new_new_n942_), .B(new_new_n528_), .Y(new_new_n943_));
  NO3        g921(.A(new_new_n831_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n944_));
  NA2        g922(.A(new_new_n480_), .B(new_new_n473_), .Y(new_new_n945_));
  NO3        g923(.A(new_new_n945_), .B(new_new_n944_), .C(new_new_n943_), .Y(new_new_n946_));
  NA3        g924(.A(new_new_n380_), .B(new_new_n174_), .C(new_new_n173_), .Y(new_new_n947_));
  NA3        g925(.A(new_new_n875_), .B(new_new_n283_), .C(new_new_n224_), .Y(new_new_n948_));
  NA2        g926(.A(new_new_n948_), .B(new_new_n947_), .Y(new_new_n949_));
  NA3        g927(.A(new_new_n380_), .B(new_new_n324_), .C(new_new_n219_), .Y(new_new_n950_));
  INV        g928(.A(new_new_n950_), .Y(new_new_n951_));
  NOi31      g929(.An(new_new_n379_), .B(new_new_n917_), .C(new_new_n234_), .Y(new_new_n952_));
  NO3        g930(.A(new_new_n872_), .B(new_new_n217_), .C(new_new_n191_), .Y(new_new_n953_));
  NO4        g931(.A(new_new_n953_), .B(new_new_n952_), .C(new_new_n951_), .D(new_new_n949_), .Y(new_new_n954_));
  NA4        g932(.A(new_new_n954_), .B(new_new_n946_), .C(new_new_n941_), .D(new_new_n939_), .Y(new_new_n955_));
  NO2        g933(.A(new_new_n86_), .B(i_5_), .Y(new_new_n956_));
  NA3        g934(.A(new_new_n826_), .B(new_new_n113_), .C(new_new_n127_), .Y(new_new_n957_));
  INV        g935(.A(new_new_n957_), .Y(new_new_n958_));
  NA2        g936(.A(new_new_n958_), .B(new_new_n956_), .Y(new_new_n959_));
  NA3        g937(.A(new_new_n296_), .B(i_5_), .C(new_new_n193_), .Y(new_new_n960_));
  NAi31      g938(.An(new_new_n236_), .B(new_new_n960_), .C(new_new_n237_), .Y(new_new_n961_));
  NO4        g939(.A(new_new_n234_), .B(new_new_n210_), .C(i_0_), .D(i_12_), .Y(new_new_n962_));
  AOI220     g940(.A0(new_new_n962_), .A1(new_new_n961_), .B0(new_new_n779_), .B1(new_new_n179_), .Y(new_new_n963_));
  NA3        g941(.A(new_new_n101_), .B(new_new_n555_), .C(i_11_), .Y(new_new_n964_));
  NO2        g942(.A(new_new_n964_), .B(new_new_n158_), .Y(new_new_n965_));
  NA2        g943(.A(new_new_n891_), .B(new_new_n463_), .Y(new_new_n966_));
  NA2        g944(.A(new_new_n64_), .B(new_new_n104_), .Y(new_new_n967_));
  OAI220     g945(.A0(new_new_n967_), .A1(new_new_n960_), .B0(new_new_n966_), .B1(new_new_n661_), .Y(new_new_n968_));
  AOI210     g946(.A0(new_new_n968_), .A1(new_new_n879_), .B0(new_new_n965_), .Y(new_new_n969_));
  NA3        g947(.A(new_new_n969_), .B(new_new_n963_), .C(new_new_n959_), .Y(new_new_n970_));
  NO4        g948(.A(new_new_n970_), .B(new_new_n955_), .C(new_new_n934_), .D(new_new_n926_), .Y(new_new_n971_));
  OAI210     g949(.A0(new_new_n799_), .A1(new_new_n795_), .B0(new_new_n37_), .Y(new_new_n972_));
  NA3        g950(.A(new_new_n887_), .B(new_new_n357_), .C(i_5_), .Y(new_new_n973_));
  NA3        g951(.A(new_new_n973_), .B(new_new_n972_), .C(new_new_n593_), .Y(new_new_n974_));
  NA2        g952(.A(new_new_n974_), .B(new_new_n208_), .Y(new_new_n975_));
  AN2        g953(.A(new_new_n678_), .B(new_new_n358_), .Y(new_new_n976_));
  NA2        g954(.A(new_new_n188_), .B(new_new_n189_), .Y(new_new_n977_));
  AO210      g955(.A0(new_new_n976_), .A1(new_new_n33_), .B0(new_new_n977_), .Y(new_new_n978_));
  NAi31      g956(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n979_));
  NO2        g957(.A(new_new_n70_), .B(new_new_n979_), .Y(new_new_n980_));
  INV        g958(.A(new_new_n980_), .Y(new_new_n981_));
  NA2        g959(.A(new_new_n981_), .B(new_new_n978_), .Y(new_new_n982_));
  NO2        g960(.A(new_new_n457_), .B(new_new_n260_), .Y(new_new_n983_));
  NO2        g961(.A(new_new_n983_), .B(new_new_n855_), .Y(new_new_n984_));
  OAI210     g962(.A0(new_new_n964_), .A1(new_new_n151_), .B0(new_new_n984_), .Y(new_new_n985_));
  AOI210     g963(.A0(new_new_n982_), .A1(new_new_n48_), .B0(new_new_n985_), .Y(new_new_n986_));
  AOI210     g964(.A0(new_new_n986_), .A1(new_new_n975_), .B0(new_new_n73_), .Y(new_new_n987_));
  INV        g965(.A(new_new_n369_), .Y(new_new_n988_));
  NO2        g966(.A(new_new_n988_), .B(new_new_n740_), .Y(new_new_n989_));
  OAI210     g967(.A0(new_new_n80_), .A1(new_new_n54_), .B0(new_new_n111_), .Y(new_new_n990_));
  NA2        g968(.A(new_new_n990_), .B(new_new_n76_), .Y(new_new_n991_));
  AOI210     g969(.A0(new_new_n940_), .A1(new_new_n875_), .B0(new_new_n892_), .Y(new_new_n992_));
  AOI210     g970(.A0(new_new_n992_), .A1(new_new_n991_), .B0(new_new_n664_), .Y(new_new_n993_));
  INV        g971(.A(new_new_n993_), .Y(new_new_n994_));
  OAI210     g972(.A0(new_new_n262_), .A1(new_new_n161_), .B0(new_new_n89_), .Y(new_new_n995_));
  NA3        g973(.A(new_new_n744_), .B(new_new_n283_), .C(new_new_n80_), .Y(new_new_n996_));
  AOI210     g974(.A0(new_new_n996_), .A1(new_new_n995_), .B0(i_11_), .Y(new_new_n997_));
  NO3        g975(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n998_));
  OAI210     g976(.A0(new_new_n895_), .A1(new_new_n297_), .B0(new_new_n998_), .Y(new_new_n999_));
  NO2        g977(.A(new_new_n999_), .B(new_new_n710_), .Y(new_new_n1000_));
  INV        g978(.A(new_new_n350_), .Y(new_new_n1001_));
  NO2        g979(.A(new_new_n1001_), .B(new_new_n41_), .Y(new_new_n1002_));
  NO3        g980(.A(new_new_n1002_), .B(new_new_n1000_), .C(new_new_n997_), .Y(new_new_n1003_));
  OAI210     g981(.A0(new_new_n994_), .A1(i_4_), .B0(new_new_n1003_), .Y(new_new_n1004_));
  NO3        g982(.A(new_new_n1004_), .B(new_new_n989_), .C(new_new_n987_), .Y(new_new_n1005_));
  NA4        g983(.A(new_new_n1005_), .B(new_new_n971_), .C(new_new_n915_), .D(new_new_n846_), .Y(ori4));
  INV        g984(.A(new_new_n682_), .Y(new_new_n1009_));
endmodule


