//Benchmark atmr_max1024_476_0.0625

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n438_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n444_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(x8), .B(x7), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n61_));
  INV        o045(.A(x9), .Y(ori_ori_n62_));
  NO2        o046(.A(ori_ori_n62_), .B(ori_ori_n36_), .Y(ori_ori_n63_));
  NO2        o047(.A(x7), .B(x6), .Y(ori_ori_n64_));
  NO2        o048(.A(ori_ori_n61_), .B(x5), .Y(ori_ori_n65_));
  NO2        o049(.A(x8), .B(x2), .Y(ori_ori_n66_));
  INV        o050(.A(ori_ori_n66_), .Y(ori_ori_n67_));
  AN2        o051(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n68_));
  OAI210     o052(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n69_), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n70_), .B(ori_ori_n68_), .Y(ori_ori_n71_));
  NA2        o055(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n73_));
  OAI210     o057(.A0(ori_ori_n73_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n74_));
  NA2        o058(.A(x5), .B(x3), .Y(ori_ori_n75_));
  NO2        o059(.A(x8), .B(x6), .Y(ori_ori_n76_));
  NO4        o060(.A(ori_ori_n76_), .B(ori_ori_n75_), .C(ori_ori_n64_), .D(ori_ori_n54_), .Y(ori_ori_n77_));
  NAi21      o061(.An(x4), .B(x3), .Y(ori_ori_n78_));
  INV        o062(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NO2        o063(.A(ori_ori_n79_), .B(ori_ori_n22_), .Y(ori_ori_n80_));
  NO2        o064(.A(x4), .B(x2), .Y(ori_ori_n81_));
  NO2        o065(.A(ori_ori_n81_), .B(x3), .Y(ori_ori_n82_));
  NO3        o066(.A(ori_ori_n82_), .B(ori_ori_n80_), .C(ori_ori_n18_), .Y(ori_ori_n83_));
  NO3        o067(.A(ori_ori_n83_), .B(ori_ori_n77_), .C(ori_ori_n74_), .Y(ori_ori_n84_));
  NA2        o068(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n85_));
  NO2        o069(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n86_));
  INV        o070(.A(x8), .Y(ori_ori_n87_));
  NA2        o071(.A(x2), .B(x1), .Y(ori_ori_n88_));
  NO2        o072(.A(ori_ori_n88_), .B(ori_ori_n87_), .Y(ori_ori_n89_));
  NO2        o073(.A(ori_ori_n89_), .B(ori_ori_n86_), .Y(ori_ori_n90_));
  NO2        o074(.A(ori_ori_n90_), .B(ori_ori_n26_), .Y(ori_ori_n91_));
  AOI210     o075(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n92_));
  OAI210     o076(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n93_));
  NO3        o077(.A(ori_ori_n93_), .B(ori_ori_n92_), .C(ori_ori_n91_), .Y(ori_ori_n94_));
  NA2        o078(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n95_));
  NO2        o079(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n96_));
  OAI210     o080(.A0(ori_ori_n96_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n97_));
  AOI210     o081(.A0(ori_ori_n95_), .A1(ori_ori_n52_), .B0(ori_ori_n97_), .Y(ori_ori_n98_));
  NO2        o082(.A(x3), .B(x2), .Y(ori_ori_n99_));
  NA3        o083(.A(ori_ori_n99_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n100_));
  INV        o084(.A(ori_ori_n100_), .Y(ori_ori_n101_));
  NA2        o085(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n102_));
  OAI210     o086(.A0(ori_ori_n102_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n103_));
  NO4        o087(.A(ori_ori_n103_), .B(ori_ori_n101_), .C(ori_ori_n98_), .D(ori_ori_n94_), .Y(ori_ori_n104_));
  AO210      o088(.A0(ori_ori_n84_), .A1(ori_ori_n72_), .B0(ori_ori_n104_), .Y(ori02));
  NO2        o089(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n106_));
  NO2        o090(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n107_));
  NA2        o091(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n108_));
  NA2        o092(.A(ori_ori_n106_), .B(x4), .Y(ori_ori_n109_));
  NO3        o093(.A(ori_ori_n109_), .B(x7), .C(x5), .Y(ori_ori_n110_));
  NA2        o094(.A(x9), .B(x2), .Y(ori_ori_n111_));
  OR2        o095(.A(x8), .B(x0), .Y(ori_ori_n112_));
  INV        o096(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  NAi21      o097(.An(x2), .B(x8), .Y(ori_ori_n114_));
  NO2        o098(.A(x4), .B(x1), .Y(ori_ori_n115_));
  NA2        o099(.A(ori_ori_n115_), .B(x2), .Y(ori_ori_n116_));
  NOi21      o100(.An(x0), .B(x1), .Y(ori_ori_n117_));
  NO3        o101(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n118_));
  NOi21      o102(.An(x0), .B(x4), .Y(ori_ori_n119_));
  NAi21      o103(.An(x8), .B(x7), .Y(ori_ori_n120_));
  NO2        o104(.A(ori_ori_n120_), .B(ori_ori_n62_), .Y(ori_ori_n121_));
  AOI220     o105(.A0(ori_ori_n121_), .A1(ori_ori_n119_), .B0(ori_ori_n118_), .B1(ori_ori_n117_), .Y(ori_ori_n122_));
  AOI210     o106(.A0(ori_ori_n122_), .A1(ori_ori_n116_), .B0(ori_ori_n75_), .Y(ori_ori_n123_));
  NO2        o107(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n124_));
  NA2        o108(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n125_));
  AOI210     o109(.A0(ori_ori_n125_), .A1(ori_ori_n102_), .B0(ori_ori_n108_), .Y(ori_ori_n126_));
  OAI210     o110(.A0(ori_ori_n126_), .A1(ori_ori_n35_), .B0(ori_ori_n124_), .Y(ori_ori_n127_));
  NAi21      o111(.An(x0), .B(x4), .Y(ori_ori_n128_));
  NO2        o112(.A(ori_ori_n128_), .B(x1), .Y(ori_ori_n129_));
  NO2        o113(.A(x7), .B(x0), .Y(ori_ori_n130_));
  NO2        o114(.A(ori_ori_n81_), .B(ori_ori_n96_), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n131_), .B(x3), .Y(ori_ori_n132_));
  OAI210     o116(.A0(ori_ori_n130_), .A1(ori_ori_n129_), .B0(ori_ori_n132_), .Y(ori_ori_n133_));
  NO2        o117(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n134_));
  NA2        o118(.A(x5), .B(x0), .Y(ori_ori_n135_));
  NO2        o119(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n136_));
  NA3        o120(.A(ori_ori_n136_), .B(ori_ori_n135_), .C(ori_ori_n134_), .Y(ori_ori_n137_));
  NA4        o121(.A(ori_ori_n137_), .B(ori_ori_n133_), .C(ori_ori_n127_), .D(ori_ori_n36_), .Y(ori_ori_n138_));
  NO3        o122(.A(ori_ori_n138_), .B(ori_ori_n123_), .C(ori_ori_n110_), .Y(ori_ori_n139_));
  NO3        o123(.A(ori_ori_n75_), .B(ori_ori_n73_), .C(ori_ori_n24_), .Y(ori_ori_n140_));
  NO2        o124(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n141_));
  AOI220     o125(.A0(ori_ori_n117_), .A1(ori_ori_n141_), .B0(ori_ori_n65_), .B1(ori_ori_n17_), .Y(ori_ori_n142_));
  NO2        o126(.A(ori_ori_n142_), .B(ori_ori_n60_), .Y(ori_ori_n143_));
  NA2        o127(.A(x7), .B(x3), .Y(ori_ori_n144_));
  NO2        o128(.A(ori_ori_n95_), .B(x5), .Y(ori_ori_n145_));
  NO2        o129(.A(x9), .B(x7), .Y(ori_ori_n146_));
  NOi21      o130(.An(x8), .B(x0), .Y(ori_ori_n147_));
  NO2        o131(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n148_));
  INV        o132(.A(x7), .Y(ori_ori_n149_));
  NA2        o133(.A(ori_ori_n149_), .B(ori_ori_n18_), .Y(ori_ori_n150_));
  AOI220     o134(.A0(ori_ori_n150_), .A1(ori_ori_n148_), .B0(ori_ori_n106_), .B1(ori_ori_n38_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n152_));
  NO2        o136(.A(ori_ori_n152_), .B(ori_ori_n119_), .Y(ori_ori_n153_));
  NO2        o137(.A(ori_ori_n153_), .B(ori_ori_n151_), .Y(ori_ori_n154_));
  INV        o138(.A(ori_ori_n154_), .Y(ori_ori_n155_));
  OAI210     o139(.A0(ori_ori_n144_), .A1(ori_ori_n50_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NA2        o140(.A(x5), .B(x1), .Y(ori_ori_n157_));
  INV        o141(.A(ori_ori_n157_), .Y(ori_ori_n158_));
  AOI210     o142(.A0(ori_ori_n158_), .A1(ori_ori_n119_), .B0(ori_ori_n36_), .Y(ori_ori_n159_));
  NAi21      o143(.An(x2), .B(x7), .Y(ori_ori_n160_));
  NO2        o144(.A(ori_ori_n160_), .B(ori_ori_n48_), .Y(ori_ori_n161_));
  NA2        o145(.A(ori_ori_n161_), .B(ori_ori_n65_), .Y(ori_ori_n162_));
  NAi31      o146(.An(ori_ori_n75_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n163_));
  NA3        o147(.A(ori_ori_n163_), .B(ori_ori_n162_), .C(ori_ori_n159_), .Y(ori_ori_n164_));
  NO4        o148(.A(ori_ori_n164_), .B(ori_ori_n156_), .C(ori_ori_n143_), .D(ori_ori_n140_), .Y(ori_ori_n165_));
  NO2        o149(.A(ori_ori_n165_), .B(ori_ori_n139_), .Y(ori_ori_n166_));
  NO2        o150(.A(ori_ori_n135_), .B(ori_ori_n131_), .Y(ori_ori_n167_));
  NA2        o151(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n168_));
  NA2        o152(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n169_));
  NA3        o153(.A(ori_ori_n169_), .B(ori_ori_n168_), .C(ori_ori_n24_), .Y(ori_ori_n170_));
  AN2        o154(.A(ori_ori_n170_), .B(ori_ori_n136_), .Y(ori_ori_n171_));
  NA2        o155(.A(x8), .B(x0), .Y(ori_ori_n172_));
  NO2        o156(.A(ori_ori_n149_), .B(ori_ori_n25_), .Y(ori_ori_n173_));
  NA2        o157(.A(x2), .B(x0), .Y(ori_ori_n174_));
  NA2        o158(.A(x4), .B(x1), .Y(ori_ori_n175_));
  NAi21      o159(.An(ori_ori_n115_), .B(ori_ori_n175_), .Y(ori_ori_n176_));
  NOi31      o160(.An(ori_ori_n176_), .B(ori_ori_n152_), .C(ori_ori_n174_), .Y(ori_ori_n177_));
  NO3        o161(.A(ori_ori_n177_), .B(ori_ori_n171_), .C(ori_ori_n167_), .Y(ori_ori_n178_));
  NO2        o162(.A(ori_ori_n178_), .B(ori_ori_n43_), .Y(ori_ori_n179_));
  NO2        o163(.A(ori_ori_n170_), .B(ori_ori_n73_), .Y(ori_ori_n180_));
  INV        o164(.A(ori_ori_n124_), .Y(ori_ori_n181_));
  NO2        o165(.A(ori_ori_n102_), .B(ori_ori_n17_), .Y(ori_ori_n182_));
  AOI210     o166(.A0(ori_ori_n35_), .A1(ori_ori_n87_), .B0(ori_ori_n182_), .Y(ori_ori_n183_));
  NO3        o167(.A(ori_ori_n183_), .B(ori_ori_n181_), .C(x7), .Y(ori_ori_n184_));
  NA3        o168(.A(ori_ori_n176_), .B(ori_ori_n181_), .C(ori_ori_n42_), .Y(ori_ori_n185_));
  OAI210     o169(.A0(ori_ori_n169_), .A1(ori_ori_n131_), .B0(ori_ori_n185_), .Y(ori_ori_n186_));
  NO3        o170(.A(ori_ori_n186_), .B(ori_ori_n184_), .C(ori_ori_n180_), .Y(ori_ori_n187_));
  NO2        o171(.A(ori_ori_n187_), .B(x3), .Y(ori_ori_n188_));
  NO3        o172(.A(ori_ori_n188_), .B(ori_ori_n179_), .C(ori_ori_n166_), .Y(ori03));
  NO2        o173(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n190_));
  NO2        o174(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n191_));
  NO2        o175(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n192_));
  OAI210     o176(.A0(ori_ori_n192_), .A1(ori_ori_n25_), .B0(ori_ori_n63_), .Y(ori_ori_n193_));
  NO2        o177(.A(ori_ori_n193_), .B(ori_ori_n17_), .Y(ori_ori_n194_));
  NA2        o178(.A(ori_ori_n194_), .B(ori_ori_n190_), .Y(ori_ori_n195_));
  NA2        o179(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n196_));
  NO2        o180(.A(ori_ori_n196_), .B(x4), .Y(ori_ori_n197_));
  NO2        o181(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n198_));
  NA2        o182(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n199_));
  NO2        o183(.A(ori_ori_n199_), .B(ori_ori_n196_), .Y(ori_ori_n200_));
  NA2        o184(.A(x9), .B(ori_ori_n54_), .Y(ori_ori_n201_));
  NA2        o185(.A(ori_ori_n201_), .B(x4), .Y(ori_ori_n202_));
  NA2        o186(.A(ori_ori_n196_), .B(ori_ori_n78_), .Y(ori_ori_n203_));
  AOI210     o187(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n174_), .Y(ori_ori_n204_));
  AOI220     o188(.A0(ori_ori_n204_), .A1(ori_ori_n203_), .B0(ori_ori_n202_), .B1(ori_ori_n200_), .Y(ori_ori_n205_));
  NO2        o189(.A(x5), .B(x1), .Y(ori_ori_n206_));
  NO2        o190(.A(ori_ori_n199_), .B(ori_ori_n168_), .Y(ori_ori_n207_));
  NO3        o191(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n208_));
  NO2        o192(.A(ori_ori_n208_), .B(ori_ori_n207_), .Y(ori_ori_n209_));
  INV        o193(.A(ori_ori_n209_), .Y(ori_ori_n210_));
  NA2        o194(.A(ori_ori_n210_), .B(ori_ori_n48_), .Y(ori_ori_n211_));
  NA3        o195(.A(ori_ori_n211_), .B(ori_ori_n205_), .C(ori_ori_n195_), .Y(ori_ori_n212_));
  NO2        o196(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n213_));
  NA2        o197(.A(ori_ori_n213_), .B(ori_ori_n19_), .Y(ori_ori_n214_));
  NO2        o198(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n215_));
  NO2        o199(.A(ori_ori_n215_), .B(x6), .Y(ori_ori_n216_));
  NOi21      o200(.An(ori_ori_n81_), .B(ori_ori_n216_), .Y(ori_ori_n217_));
  NA2        o201(.A(ori_ori_n62_), .B(ori_ori_n87_), .Y(ori_ori_n218_));
  NA3        o202(.A(ori_ori_n218_), .B(ori_ori_n215_), .C(x6), .Y(ori_ori_n219_));
  AOI210     o203(.A0(ori_ori_n219_), .A1(ori_ori_n217_), .B0(ori_ori_n149_), .Y(ori_ori_n220_));
  AO210      o204(.A0(ori_ori_n220_), .A1(ori_ori_n214_), .B0(ori_ori_n173_), .Y(ori_ori_n221_));
  NA2        o205(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n222_));
  OAI210     o206(.A0(ori_ori_n222_), .A1(ori_ori_n25_), .B0(ori_ori_n169_), .Y(ori_ori_n223_));
  NO2        o207(.A(ori_ori_n175_), .B(x6), .Y(ori_ori_n224_));
  AOI220     o208(.A0(ori_ori_n224_), .A1(ori_ori_n223_), .B0(ori_ori_n136_), .B1(ori_ori_n86_), .Y(ori_ori_n225_));
  NA2        o209(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n226_));
  OAI210     o210(.A0(ori_ori_n113_), .A1(ori_ori_n76_), .B0(x4), .Y(ori_ori_n227_));
  AOI210     o211(.A0(ori_ori_n227_), .A1(ori_ori_n226_), .B0(ori_ori_n75_), .Y(ori_ori_n228_));
  NO2        o212(.A(ori_ori_n157_), .B(ori_ori_n43_), .Y(ori_ori_n229_));
  OAI210     o213(.A0(ori_ori_n229_), .A1(ori_ori_n207_), .B0(ori_ori_n438_), .Y(ori_ori_n230_));
  NA2        o214(.A(ori_ori_n191_), .B(ori_ori_n129_), .Y(ori_ori_n231_));
  NA3        o215(.A(ori_ori_n199_), .B(ori_ori_n124_), .C(x6), .Y(ori_ori_n232_));
  OAI210     o216(.A0(ori_ori_n87_), .A1(ori_ori_n36_), .B0(ori_ori_n65_), .Y(ori_ori_n233_));
  NA4        o217(.A(ori_ori_n233_), .B(ori_ori_n232_), .C(ori_ori_n231_), .D(ori_ori_n230_), .Y(ori_ori_n234_));
  OAI210     o218(.A0(ori_ori_n234_), .A1(ori_ori_n228_), .B0(x2), .Y(ori_ori_n235_));
  NA3        o219(.A(ori_ori_n235_), .B(ori_ori_n225_), .C(ori_ori_n221_), .Y(ori_ori_n236_));
  AOI210     o220(.A0(ori_ori_n212_), .A1(x8), .B0(ori_ori_n236_), .Y(ori_ori_n237_));
  NO2        o221(.A(ori_ori_n87_), .B(x3), .Y(ori_ori_n238_));
  NA2        o222(.A(ori_ori_n238_), .B(ori_ori_n197_), .Y(ori_ori_n239_));
  NO2        o223(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n240_));
  AOI210     o224(.A0(ori_ori_n216_), .A1(ori_ori_n152_), .B0(ori_ori_n240_), .Y(ori_ori_n241_));
  AOI210     o225(.A0(ori_ori_n241_), .A1(ori_ori_n239_), .B0(x2), .Y(ori_ori_n242_));
  NO2        o226(.A(x4), .B(ori_ori_n54_), .Y(ori_ori_n243_));
  AOI220     o227(.A0(ori_ori_n197_), .A1(ori_ori_n182_), .B0(ori_ori_n243_), .B1(ori_ori_n65_), .Y(ori_ori_n244_));
  NA2        o228(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n245_));
  NA3        o229(.A(ori_ori_n25_), .B(x3), .C(x2), .Y(ori_ori_n246_));
  AOI210     o230(.A0(ori_ori_n246_), .A1(ori_ori_n135_), .B0(ori_ori_n245_), .Y(ori_ori_n247_));
  NA2        o231(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n248_));
  NO2        o232(.A(ori_ori_n248_), .B(ori_ori_n25_), .Y(ori_ori_n249_));
  OAI210     o233(.A0(ori_ori_n249_), .A1(ori_ori_n247_), .B0(ori_ori_n115_), .Y(ori_ori_n250_));
  NA2        o234(.A(ori_ori_n199_), .B(x6), .Y(ori_ori_n251_));
  NO2        o235(.A(ori_ori_n199_), .B(x6), .Y(ori_ori_n252_));
  INV        o236(.A(ori_ori_n252_), .Y(ori_ori_n253_));
  NA3        o237(.A(ori_ori_n253_), .B(ori_ori_n251_), .C(ori_ori_n141_), .Y(ori_ori_n254_));
  NA4        o238(.A(ori_ori_n254_), .B(ori_ori_n250_), .C(ori_ori_n244_), .D(ori_ori_n149_), .Y(ori_ori_n255_));
  NA2        o239(.A(ori_ori_n191_), .B(ori_ori_n215_), .Y(ori_ori_n256_));
  NO2        o240(.A(x9), .B(x6), .Y(ori_ori_n257_));
  NO2        o241(.A(ori_ori_n135_), .B(ori_ori_n18_), .Y(ori_ori_n258_));
  NAi21      o242(.An(ori_ori_n258_), .B(ori_ori_n246_), .Y(ori_ori_n259_));
  NAi21      o243(.An(x1), .B(x4), .Y(ori_ori_n260_));
  AOI210     o244(.A0(x3), .A1(x2), .B0(ori_ori_n48_), .Y(ori_ori_n261_));
  OAI210     o245(.A0(ori_ori_n135_), .A1(x3), .B0(ori_ori_n261_), .Y(ori_ori_n262_));
  AOI220     o246(.A0(ori_ori_n262_), .A1(ori_ori_n260_), .B0(ori_ori_n259_), .B1(ori_ori_n257_), .Y(ori_ori_n263_));
  NA2        o247(.A(ori_ori_n263_), .B(ori_ori_n256_), .Y(ori_ori_n264_));
  NA2        o248(.A(ori_ori_n62_), .B(x2), .Y(ori_ori_n265_));
  NO2        o249(.A(ori_ori_n265_), .B(ori_ori_n256_), .Y(ori_ori_n266_));
  NA2        o250(.A(x6), .B(x2), .Y(ori_ori_n267_));
  OAI210     o251(.A0(x4), .A1(ori_ori_n266_), .B0(ori_ori_n264_), .Y(ori_ori_n268_));
  NO2        o252(.A(x3), .B(ori_ori_n196_), .Y(ori_ori_n269_));
  NA2        o253(.A(x4), .B(x0), .Y(ori_ori_n270_));
  NA2        o254(.A(ori_ori_n269_), .B(ori_ori_n42_), .Y(ori_ori_n271_));
  AOI210     o255(.A0(ori_ori_n271_), .A1(ori_ori_n268_), .B0(x8), .Y(ori_ori_n272_));
  INV        o256(.A(ori_ori_n245_), .Y(ori_ori_n273_));
  NA2        o257(.A(ori_ori_n258_), .B(ori_ori_n273_), .Y(ori_ori_n274_));
  INV        o258(.A(ori_ori_n172_), .Y(ori_ori_n275_));
  OAI210     o259(.A0(ori_ori_n275_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n276_));
  AOI210     o260(.A0(ori_ori_n276_), .A1(ori_ori_n274_), .B0(ori_ori_n222_), .Y(ori_ori_n277_));
  NO4        o261(.A(ori_ori_n277_), .B(ori_ori_n272_), .C(ori_ori_n255_), .D(ori_ori_n242_), .Y(ori_ori_n278_));
  INV        o262(.A(x1), .Y(ori_ori_n279_));
  NO3        o263(.A(ori_ori_n279_), .B(x3), .C(ori_ori_n36_), .Y(ori_ori_n280_));
  OAI210     o264(.A0(ori_ori_n280_), .A1(ori_ori_n252_), .B0(x2), .Y(ori_ori_n281_));
  OAI210     o265(.A0(ori_ori_n275_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n282_));
  AOI210     o266(.A0(ori_ori_n282_), .A1(ori_ori_n281_), .B0(ori_ori_n181_), .Y(ori_ori_n283_));
  NOi21      o267(.An(ori_ori_n267_), .B(ori_ori_n17_), .Y(ori_ori_n284_));
  NA3        o268(.A(ori_ori_n284_), .B(ori_ori_n206_), .C(ori_ori_n40_), .Y(ori_ori_n285_));
  AOI210     o269(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n286_));
  NA3        o270(.A(ori_ori_n286_), .B(ori_ori_n158_), .C(ori_ori_n32_), .Y(ori_ori_n287_));
  NA2        o271(.A(x3), .B(x2), .Y(ori_ori_n288_));
  AOI220     o272(.A0(ori_ori_n288_), .A1(ori_ori_n222_), .B0(ori_ori_n287_), .B1(ori_ori_n285_), .Y(ori_ori_n289_));
  NAi21      o273(.An(x4), .B(x0), .Y(ori_ori_n290_));
  NO3        o274(.A(ori_ori_n290_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n291_));
  OAI210     o275(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n291_), .Y(ori_ori_n292_));
  OAI220     o276(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n293_));
  NO2        o277(.A(x9), .B(x8), .Y(ori_ori_n294_));
  NA3        o278(.A(ori_ori_n294_), .B(ori_ori_n36_), .C(ori_ori_n54_), .Y(ori_ori_n295_));
  OAI210     o279(.A0(ori_ori_n286_), .A1(ori_ori_n284_), .B0(ori_ori_n295_), .Y(ori_ori_n296_));
  AOI220     o280(.A0(ori_ori_n296_), .A1(ori_ori_n79_), .B0(ori_ori_n293_), .B1(ori_ori_n31_), .Y(ori_ori_n297_));
  AOI210     o281(.A0(ori_ori_n297_), .A1(ori_ori_n292_), .B0(ori_ori_n25_), .Y(ori_ori_n298_));
  NA3        o282(.A(ori_ori_n36_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n299_));
  OAI210     o283(.A0(ori_ori_n286_), .A1(ori_ori_n284_), .B0(ori_ori_n299_), .Y(ori_ori_n300_));
  INV        o284(.A(ori_ori_n207_), .Y(ori_ori_n301_));
  NA2        o285(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n302_));
  OR2        o286(.A(ori_ori_n302_), .B(ori_ori_n270_), .Y(ori_ori_n303_));
  OAI220     o287(.A0(ori_ori_n303_), .A1(ori_ori_n157_), .B0(ori_ori_n226_), .B1(ori_ori_n301_), .Y(ori_ori_n304_));
  AO210      o288(.A0(ori_ori_n300_), .A1(ori_ori_n145_), .B0(ori_ori_n304_), .Y(ori_ori_n305_));
  NO4        o289(.A(ori_ori_n305_), .B(ori_ori_n298_), .C(ori_ori_n289_), .D(ori_ori_n283_), .Y(ori_ori_n306_));
  OAI210     o290(.A0(ori_ori_n278_), .A1(ori_ori_n237_), .B0(ori_ori_n306_), .Y(ori04));
  NO2        o291(.A(x2), .B(x1), .Y(ori_ori_n308_));
  OAI210     o292(.A0(ori_ori_n248_), .A1(ori_ori_n308_), .B0(ori_ori_n36_), .Y(ori_ori_n309_));
  NO2        o293(.A(ori_ori_n308_), .B(ori_ori_n290_), .Y(ori_ori_n310_));
  OAI210     o294(.A0(ori_ori_n54_), .A1(ori_ori_n310_), .B0(ori_ori_n238_), .Y(ori_ori_n311_));
  NO2        o295(.A(ori_ori_n265_), .B(ori_ori_n85_), .Y(ori_ori_n312_));
  NO2        o296(.A(ori_ori_n312_), .B(ori_ori_n36_), .Y(ori_ori_n313_));
  NO2        o297(.A(ori_ori_n288_), .B(ori_ori_n198_), .Y(ori_ori_n314_));
  NA2        o298(.A(ori_ori_n314_), .B(ori_ori_n87_), .Y(ori_ori_n315_));
  NA3        o299(.A(ori_ori_n315_), .B(ori_ori_n313_), .C(ori_ori_n311_), .Y(ori_ori_n316_));
  NA2        o300(.A(ori_ori_n316_), .B(ori_ori_n309_), .Y(ori_ori_n317_));
  OAI210     o301(.A0(ori_ori_n112_), .A1(ori_ori_n102_), .B0(ori_ori_n172_), .Y(ori_ori_n318_));
  NA3        o302(.A(ori_ori_n318_), .B(x6), .C(x3), .Y(ori_ori_n319_));
  NOi21      o303(.An(ori_ori_n147_), .B(ori_ori_n125_), .Y(ori_ori_n320_));
  AOI210     o304(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n321_));
  OAI220     o305(.A0(ori_ori_n321_), .A1(ori_ori_n302_), .B0(ori_ori_n265_), .B1(ori_ori_n299_), .Y(ori_ori_n322_));
  AOI210     o306(.A0(ori_ori_n320_), .A1(ori_ori_n63_), .B0(ori_ori_n322_), .Y(ori_ori_n323_));
  NA2        o307(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n324_));
  OAI210     o308(.A0(ori_ori_n102_), .A1(ori_ori_n17_), .B0(ori_ori_n324_), .Y(ori_ori_n325_));
  AOI220     o309(.A0(ori_ori_n325_), .A1(ori_ori_n76_), .B0(ori_ori_n312_), .B1(ori_ori_n87_), .Y(ori_ori_n326_));
  NA3        o310(.A(ori_ori_n326_), .B(ori_ori_n323_), .C(ori_ori_n319_), .Y(ori_ori_n327_));
  OAI210     o311(.A0(ori_ori_n107_), .A1(x3), .B0(ori_ori_n291_), .Y(ori_ori_n328_));
  NA2        o312(.A(ori_ori_n328_), .B(ori_ori_n149_), .Y(ori_ori_n329_));
  AOI210     o313(.A0(ori_ori_n327_), .A1(x4), .B0(ori_ori_n329_), .Y(ori_ori_n330_));
  NA3        o314(.A(ori_ori_n310_), .B(ori_ori_n201_), .C(ori_ori_n87_), .Y(ori_ori_n331_));
  XO2        o315(.A(x4), .B(x0), .Y(ori_ori_n332_));
  OAI210     o316(.A0(ori_ori_n332_), .A1(ori_ori_n111_), .B0(ori_ori_n260_), .Y(ori_ori_n333_));
  AOI220     o317(.A0(ori_ori_n333_), .A1(x8), .B0(x4), .B1(ori_ori_n88_), .Y(ori_ori_n334_));
  AOI210     o318(.A0(ori_ori_n334_), .A1(ori_ori_n331_), .B0(x3), .Y(ori_ori_n335_));
  INV        o319(.A(ori_ori_n88_), .Y(ori_ori_n336_));
  NO2        o320(.A(ori_ori_n87_), .B(x4), .Y(ori_ori_n337_));
  AOI220     o321(.A0(ori_ori_n337_), .A1(ori_ori_n44_), .B0(ori_ori_n119_), .B1(ori_ori_n336_), .Y(ori_ori_n338_));
  NO2        o322(.A(ori_ori_n332_), .B(x2), .Y(ori_ori_n339_));
  NO3        o323(.A(ori_ori_n218_), .B(ori_ori_n28_), .C(ori_ori_n24_), .Y(ori_ori_n340_));
  NO2        o324(.A(ori_ori_n340_), .B(ori_ori_n339_), .Y(ori_ori_n341_));
  NA4        o325(.A(ori_ori_n341_), .B(ori_ori_n338_), .C(ori_ori_n214_), .D(x6), .Y(ori_ori_n342_));
  OAI220     o326(.A0(ori_ori_n290_), .A1(ori_ori_n85_), .B0(ori_ori_n174_), .B1(ori_ori_n87_), .Y(ori_ori_n343_));
  NO2        o327(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n344_));
  OR2        o328(.A(ori_ori_n337_), .B(ori_ori_n344_), .Y(ori_ori_n345_));
  NO2        o329(.A(ori_ori_n147_), .B(ori_ori_n102_), .Y(ori_ori_n346_));
  AOI220     o330(.A0(ori_ori_n346_), .A1(ori_ori_n345_), .B0(ori_ori_n343_), .B1(ori_ori_n61_), .Y(ori_ori_n347_));
  NO2        o331(.A(ori_ori_n147_), .B(ori_ori_n78_), .Y(ori_ori_n348_));
  NO2        o332(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n349_));
  NOi21      o333(.An(ori_ori_n115_), .B(ori_ori_n27_), .Y(ori_ori_n350_));
  AOI210     o334(.A0(ori_ori_n349_), .A1(ori_ori_n348_), .B0(ori_ori_n350_), .Y(ori_ori_n351_));
  OAI210     o335(.A0(ori_ori_n347_), .A1(ori_ori_n62_), .B0(ori_ori_n351_), .Y(ori_ori_n352_));
  OAI220     o336(.A0(ori_ori_n352_), .A1(x6), .B0(ori_ori_n342_), .B1(ori_ori_n335_), .Y(ori_ori_n353_));
  OAI210     o337(.A0(ori_ori_n63_), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n354_));
  OAI210     o338(.A0(ori_ori_n354_), .A1(ori_ori_n87_), .B0(ori_ori_n303_), .Y(ori_ori_n355_));
  AOI210     o339(.A0(ori_ori_n355_), .A1(ori_ori_n18_), .B0(ori_ori_n149_), .Y(ori_ori_n356_));
  AO220      o340(.A0(ori_ori_n356_), .A1(ori_ori_n353_), .B0(ori_ori_n330_), .B1(ori_ori_n317_), .Y(ori_ori_n357_));
  NA2        o341(.A(ori_ori_n208_), .B(ori_ori_n49_), .Y(ori_ori_n358_));
  NA2        o342(.A(ori_ori_n358_), .B(ori_ori_n357_), .Y(ori_ori_n359_));
  AOI210     o343(.A0(ori_ori_n192_), .A1(x8), .B0(ori_ori_n107_), .Y(ori_ori_n360_));
  NA2        o344(.A(ori_ori_n360_), .B(ori_ori_n324_), .Y(ori_ori_n361_));
  NA3        o345(.A(ori_ori_n361_), .B(ori_ori_n190_), .C(ori_ori_n149_), .Y(ori_ori_n362_));
  NA3        o346(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n363_));
  NA2        o347(.A(ori_ori_n213_), .B(x0), .Y(ori_ori_n364_));
  OAI220     o348(.A0(ori_ori_n364_), .A1(ori_ori_n201_), .B0(ori_ori_n363_), .B1(ori_ori_n336_), .Y(ori_ori_n365_));
  INV        o349(.A(ori_ori_n365_), .Y(ori_ori_n366_));
  AOI210     o350(.A0(ori_ori_n366_), .A1(ori_ori_n362_), .B0(ori_ori_n25_), .Y(ori_ori_n367_));
  OAI210     o351(.A0(ori_ori_n190_), .A1(ori_ori_n66_), .B0(ori_ori_n198_), .Y(ori_ori_n368_));
  NA3        o352(.A(ori_ori_n192_), .B(ori_ori_n215_), .C(x8), .Y(ori_ori_n369_));
  AOI210     o353(.A0(ori_ori_n369_), .A1(ori_ori_n368_), .B0(ori_ori_n25_), .Y(ori_ori_n370_));
  AOI210     o354(.A0(ori_ori_n114_), .A1(ori_ori_n112_), .B0(ori_ori_n42_), .Y(ori_ori_n371_));
  NOi31      o355(.An(ori_ori_n371_), .B(ori_ori_n344_), .C(ori_ori_n175_), .Y(ori_ori_n372_));
  OAI210     o356(.A0(ori_ori_n372_), .A1(ori_ori_n370_), .B0(ori_ori_n146_), .Y(ori_ori_n373_));
  INV        o357(.A(ori_ori_n373_), .Y(ori_ori_n374_));
  OAI210     o358(.A0(ori_ori_n374_), .A1(ori_ori_n367_), .B0(x6), .Y(ori_ori_n375_));
  NA2        o359(.A(ori_ori_n48_), .B(ori_ori_n130_), .Y(ori_ori_n376_));
  NA3        o360(.A(ori_ori_n55_), .B(ori_ori_n38_), .C(ori_ori_n31_), .Y(ori_ori_n377_));
  AOI220     o361(.A0(ori_ori_n377_), .A1(ori_ori_n376_), .B0(ori_ori_n40_), .B1(ori_ori_n32_), .Y(ori_ori_n378_));
  NO2        o362(.A(ori_ori_n149_), .B(x0), .Y(ori_ori_n379_));
  AOI220     o363(.A0(ori_ori_n379_), .A1(ori_ori_n213_), .B0(ori_ori_n190_), .B1(ori_ori_n149_), .Y(ori_ori_n380_));
  AOI210     o364(.A0(ori_ori_n121_), .A1(ori_ori_n243_), .B0(x1), .Y(ori_ori_n381_));
  OAI210     o365(.A0(ori_ori_n380_), .A1(x8), .B0(ori_ori_n381_), .Y(ori_ori_n382_));
  NAi31      o366(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n383_));
  OAI210     o367(.A0(ori_ori_n383_), .A1(x4), .B0(ori_ori_n160_), .Y(ori_ori_n384_));
  NA3        o368(.A(ori_ori_n384_), .B(ori_ori_n144_), .C(x9), .Y(ori_ori_n385_));
  NO4        o369(.A(ori_ori_n120_), .B(ori_ori_n290_), .C(x9), .D(x2), .Y(ori_ori_n386_));
  NOi21      o370(.An(ori_ori_n118_), .B(ori_ori_n174_), .Y(ori_ori_n387_));
  NO3        o371(.A(ori_ori_n387_), .B(ori_ori_n386_), .C(ori_ori_n18_), .Y(ori_ori_n388_));
  NO3        o372(.A(x9), .B(ori_ori_n149_), .C(x0), .Y(ori_ori_n389_));
  AOI220     o373(.A0(ori_ori_n389_), .A1(ori_ori_n238_), .B0(ori_ori_n348_), .B1(ori_ori_n149_), .Y(ori_ori_n390_));
  NA4        o374(.A(ori_ori_n390_), .B(ori_ori_n388_), .C(ori_ori_n385_), .D(ori_ori_n50_), .Y(ori_ori_n391_));
  OAI210     o375(.A0(ori_ori_n382_), .A1(ori_ori_n378_), .B0(ori_ori_n391_), .Y(ori_ori_n392_));
  NOi31      o376(.An(ori_ori_n379_), .B(ori_ori_n32_), .C(x8), .Y(ori_ori_n393_));
  AOI210     o377(.A0(ori_ori_n38_), .A1(x9), .B0(ori_ori_n128_), .Y(ori_ori_n394_));
  NO3        o378(.A(ori_ori_n394_), .B(ori_ori_n118_), .C(ori_ori_n43_), .Y(ori_ori_n395_));
  AOI210     o379(.A0(ori_ori_n260_), .A1(ori_ori_n60_), .B0(ori_ori_n117_), .Y(ori_ori_n396_));
  NO2        o380(.A(ori_ori_n396_), .B(x3), .Y(ori_ori_n397_));
  NO3        o381(.A(ori_ori_n397_), .B(ori_ori_n395_), .C(x2), .Y(ori_ori_n398_));
  OAI220     o382(.A0(ori_ori_n332_), .A1(ori_ori_n294_), .B0(ori_ori_n290_), .B1(ori_ori_n43_), .Y(ori_ori_n399_));
  AOI210     o383(.A0(x9), .A1(ori_ori_n48_), .B0(ori_ori_n363_), .Y(ori_ori_n400_));
  AOI220     o384(.A0(ori_ori_n400_), .A1(ori_ori_n87_), .B0(ori_ori_n399_), .B1(ori_ori_n149_), .Y(ori_ori_n401_));
  NO2        o385(.A(ori_ori_n401_), .B(ori_ori_n54_), .Y(ori_ori_n402_));
  NO3        o386(.A(ori_ori_n402_), .B(ori_ori_n398_), .C(ori_ori_n393_), .Y(ori_ori_n403_));
  AOI210     o387(.A0(ori_ori_n403_), .A1(ori_ori_n392_), .B0(ori_ori_n25_), .Y(ori_ori_n404_));
  NA4        o388(.A(ori_ori_n31_), .B(ori_ori_n87_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n405_));
  NO3        o389(.A(ori_ori_n62_), .B(x4), .C(x1), .Y(ori_ori_n406_));
  NO3        o390(.A(ori_ori_n66_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n407_));
  AOI220     o391(.A0(ori_ori_n407_), .A1(ori_ori_n261_), .B0(ori_ori_n406_), .B1(ori_ori_n371_), .Y(ori_ori_n408_));
  NO2        o392(.A(ori_ori_n408_), .B(ori_ori_n99_), .Y(ori_ori_n409_));
  NO3        o393(.A(ori_ori_n265_), .B(ori_ori_n172_), .C(ori_ori_n40_), .Y(ori_ori_n410_));
  OAI210     o394(.A0(ori_ori_n410_), .A1(ori_ori_n409_), .B0(x7), .Y(ori_ori_n411_));
  NA2        o395(.A(ori_ori_n218_), .B(x7), .Y(ori_ori_n412_));
  NA3        o396(.A(ori_ori_n412_), .B(ori_ori_n148_), .C(ori_ori_n129_), .Y(ori_ori_n413_));
  NA3        o397(.A(ori_ori_n413_), .B(ori_ori_n411_), .C(ori_ori_n405_), .Y(ori_ori_n414_));
  OAI210     o398(.A0(ori_ori_n414_), .A1(ori_ori_n404_), .B0(ori_ori_n36_), .Y(ori_ori_n415_));
  NO2        o399(.A(ori_ori_n389_), .B(ori_ori_n198_), .Y(ori_ori_n416_));
  NO4        o400(.A(ori_ori_n416_), .B(ori_ori_n75_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n417_));
  NA2        o401(.A(ori_ori_n248_), .B(ori_ori_n21_), .Y(ori_ori_n418_));
  NO2        o402(.A(ori_ori_n157_), .B(ori_ori_n130_), .Y(ori_ori_n419_));
  NA2        o403(.A(ori_ori_n419_), .B(ori_ori_n418_), .Y(ori_ori_n420_));
  AOI210     o404(.A0(ori_ori_n420_), .A1(ori_ori_n163_), .B0(ori_ori_n28_), .Y(ori_ori_n421_));
  AOI220     o405(.A0(ori_ori_n344_), .A1(ori_ori_n87_), .B0(ori_ori_n147_), .B1(ori_ori_n192_), .Y(ori_ori_n422_));
  NA3        o406(.A(ori_ori_n422_), .B(ori_ori_n383_), .C(ori_ori_n85_), .Y(ori_ori_n423_));
  NA2        o407(.A(ori_ori_n423_), .B(ori_ori_n173_), .Y(ori_ori_n424_));
  OAI220     o408(.A0(x3), .A1(ori_ori_n67_), .B0(ori_ori_n157_), .B1(ori_ori_n43_), .Y(ori_ori_n425_));
  NA2        o409(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n426_));
  OAI210     o410(.A0(ori_ori_n146_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n427_));
  NO2        o411(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n428_));
  NA2        o412(.A(ori_ori_n428_), .B(ori_ori_n427_), .Y(ori_ori_n429_));
  OAI210     o413(.A0(ori_ori_n150_), .A1(ori_ori_n426_), .B0(ori_ori_n429_), .Y(ori_ori_n430_));
  AOI220     o414(.A0(ori_ori_n430_), .A1(x0), .B0(ori_ori_n425_), .B1(ori_ori_n130_), .Y(ori_ori_n431_));
  AOI210     o415(.A0(ori_ori_n431_), .A1(ori_ori_n424_), .B0(ori_ori_n226_), .Y(ori_ori_n432_));
  NO3        o416(.A(ori_ori_n432_), .B(ori_ori_n421_), .C(ori_ori_n417_), .Y(ori_ori_n433_));
  NA3        o417(.A(ori_ori_n433_), .B(ori_ori_n415_), .C(ori_ori_n375_), .Y(ori_ori_n434_));
  AOI210     o418(.A0(ori_ori_n359_), .A1(ori_ori_n25_), .B0(ori_ori_n434_), .Y(ori05));
  INV        o419(.A(x6), .Y(ori_ori_n438_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  INV        m005(.A(mai_mai_n19_), .Y(mai_mai_n22_));
  NA2        m006(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n23_));
  INV        m007(.A(x5), .Y(mai_mai_n24_));
  NA2        m008(.A(x7), .B(x6), .Y(mai_mai_n25_));
  NA2        m009(.A(x8), .B(x3), .Y(mai_mai_n26_));
  NA2        m010(.A(x4), .B(x2), .Y(mai_mai_n27_));
  INV        m011(.A(mai_mai_n23_), .Y(mai_mai_n28_));
  NO2        m012(.A(x4), .B(x3), .Y(mai_mai_n29_));
  INV        m013(.A(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m014(.An(mai_mai_n22_), .B(mai_mai_n28_), .Y(mai00));
  NO2        m015(.A(x1), .B(x0), .Y(mai_mai_n32_));
  INV        m016(.A(x6), .Y(mai_mai_n33_));
  NO2        m017(.A(mai_mai_n33_), .B(mai_mai_n24_), .Y(mai_mai_n34_));
  AN2        m018(.A(x8), .B(x7), .Y(mai_mai_n35_));
  NA3        m019(.A(mai_mai_n35_), .B(mai_mai_n34_), .C(mai_mai_n32_), .Y(mai_mai_n36_));
  NA2        m020(.A(x4), .B(x3), .Y(mai_mai_n37_));
  AOI210     m021(.A0(mai_mai_n36_), .A1(mai_mai_n22_), .B0(mai_mai_n37_), .Y(mai_mai_n38_));
  NO2        m022(.A(x2), .B(x0), .Y(mai_mai_n39_));
  INV        m023(.A(x3), .Y(mai_mai_n40_));
  NO2        m024(.A(mai_mai_n40_), .B(mai_mai_n18_), .Y(mai_mai_n41_));
  INV        m025(.A(mai_mai_n41_), .Y(mai_mai_n42_));
  NO2        m026(.A(mai_mai_n34_), .B(x4), .Y(mai_mai_n43_));
  OAI210     m027(.A0(mai_mai_n43_), .A1(mai_mai_n42_), .B0(mai_mai_n39_), .Y(mai_mai_n44_));
  INV        m028(.A(x4), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n45_), .B(mai_mai_n17_), .Y(mai_mai_n46_));
  NA2        m030(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n47_));
  OAI210     m031(.A0(mai_mai_n47_), .A1(mai_mai_n20_), .B0(mai_mai_n44_), .Y(mai_mai_n48_));
  NA2        m032(.A(mai_mai_n35_), .B(mai_mai_n34_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(mai_mai_n32_), .Y(mai_mai_n50_));
  INV        m034(.A(x2), .Y(mai_mai_n51_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n17_), .Y(mai_mai_n52_));
  NA2        m036(.A(mai_mai_n40_), .B(mai_mai_n18_), .Y(mai_mai_n53_));
  NA2        m037(.A(mai_mai_n53_), .B(mai_mai_n52_), .Y(mai_mai_n54_));
  OAI210     m038(.A0(mai_mai_n50_), .A1(mai_mai_n30_), .B0(mai_mai_n54_), .Y(mai_mai_n55_));
  NO3        m039(.A(mai_mai_n55_), .B(mai_mai_n48_), .C(mai_mai_n38_), .Y(mai01));
  NA2        m040(.A(x8), .B(x7), .Y(mai_mai_n57_));
  NA2        m041(.A(mai_mai_n40_), .B(x1), .Y(mai_mai_n58_));
  INV        m042(.A(x9), .Y(mai_mai_n59_));
  NO2        m043(.A(mai_mai_n59_), .B(mai_mai_n33_), .Y(mai_mai_n60_));
  INV        m044(.A(mai_mai_n60_), .Y(mai_mai_n61_));
  NO3        m045(.A(mai_mai_n61_), .B(mai_mai_n58_), .C(mai_mai_n57_), .Y(mai_mai_n62_));
  NO2        m046(.A(x7), .B(x6), .Y(mai_mai_n63_));
  NO2        m047(.A(mai_mai_n58_), .B(x5), .Y(mai_mai_n64_));
  NO2        m048(.A(x8), .B(x2), .Y(mai_mai_n65_));
  OA210      m049(.A0(mai_mai_n65_), .A1(mai_mai_n64_), .B0(mai_mai_n63_), .Y(mai_mai_n66_));
  OAI210     m050(.A0(mai_mai_n41_), .A1(mai_mai_n24_), .B0(mai_mai_n51_), .Y(mai_mai_n67_));
  OAI210     m051(.A0(mai_mai_n53_), .A1(mai_mai_n20_), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  NAi31      m052(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n69_));
  OAI220     m053(.A0(mai_mai_n69_), .A1(mai_mai_n40_), .B0(mai_mai_n68_), .B1(mai_mai_n66_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n70_), .A1(mai_mai_n62_), .B0(x4), .Y(mai_mai_n71_));
  NA2        m055(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n72_));
  OAI210     m056(.A0(mai_mai_n72_), .A1(mai_mai_n53_), .B0(x0), .Y(mai_mai_n73_));
  NA2        m057(.A(x5), .B(x3), .Y(mai_mai_n74_));
  NO2        m058(.A(x8), .B(x6), .Y(mai_mai_n75_));
  NO4        m059(.A(mai_mai_n75_), .B(mai_mai_n74_), .C(mai_mai_n63_), .D(mai_mai_n51_), .Y(mai_mai_n76_));
  NAi21      m060(.An(x4), .B(x3), .Y(mai_mai_n77_));
  INV        m061(.A(mai_mai_n77_), .Y(mai_mai_n78_));
  NO2        m062(.A(x4), .B(x2), .Y(mai_mai_n79_));
  NO2        m063(.A(mai_mai_n79_), .B(x3), .Y(mai_mai_n80_));
  NO2        m064(.A(mai_mai_n77_), .B(mai_mai_n18_), .Y(mai_mai_n81_));
  NO3        m065(.A(mai_mai_n81_), .B(mai_mai_n76_), .C(mai_mai_n73_), .Y(mai_mai_n82_));
  NO4        m066(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n40_), .D(x1), .Y(mai_mai_n83_));
  NA2        m067(.A(mai_mai_n83_), .B(mai_mai_n45_), .Y(mai_mai_n84_));
  NA2        m068(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n85_));
  NO2        m069(.A(mai_mai_n85_), .B(mai_mai_n24_), .Y(mai_mai_n86_));
  INV        m070(.A(x8), .Y(mai_mai_n87_));
  NA2        m071(.A(x2), .B(x1), .Y(mai_mai_n88_));
  INV        m072(.A(mai_mai_n86_), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n89_), .B(mai_mai_n25_), .Y(mai_mai_n90_));
  AOI210     m074(.A0(mai_mai_n53_), .A1(mai_mai_n24_), .B0(mai_mai_n51_), .Y(mai_mai_n91_));
  OAI210     m075(.A0(mai_mai_n42_), .A1(mai_mai_n34_), .B0(mai_mai_n45_), .Y(mai_mai_n92_));
  NO3        m076(.A(mai_mai_n92_), .B(mai_mai_n91_), .C(mai_mai_n90_), .Y(mai_mai_n93_));
  NA2        m077(.A(x4), .B(mai_mai_n40_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n45_), .B(mai_mai_n51_), .Y(mai_mai_n95_));
  OAI210     m079(.A0(mai_mai_n95_), .A1(mai_mai_n40_), .B0(mai_mai_n18_), .Y(mai_mai_n96_));
  AOI210     m080(.A0(mai_mai_n94_), .A1(mai_mai_n49_), .B0(mai_mai_n96_), .Y(mai_mai_n97_));
  NO2        m081(.A(x3), .B(x2), .Y(mai_mai_n98_));
  NA3        m082(.A(mai_mai_n98_), .B(mai_mai_n25_), .C(mai_mai_n24_), .Y(mai_mai_n99_));
  AOI210     m083(.A0(x8), .A1(x6), .B0(mai_mai_n99_), .Y(mai_mai_n100_));
  NA2        m084(.A(mai_mai_n51_), .B(x1), .Y(mai_mai_n101_));
  OAI210     m085(.A0(mai_mai_n101_), .A1(mai_mai_n37_), .B0(mai_mai_n17_), .Y(mai_mai_n102_));
  NO4        m086(.A(mai_mai_n102_), .B(mai_mai_n100_), .C(mai_mai_n97_), .D(mai_mai_n93_), .Y(mai_mai_n103_));
  AO220      m087(.A0(mai_mai_n103_), .A1(mai_mai_n84_), .B0(mai_mai_n82_), .B1(mai_mai_n71_), .Y(mai02));
  NO2        m088(.A(x3), .B(mai_mai_n51_), .Y(mai_mai_n105_));
  NO2        m089(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n106_));
  NA2        m090(.A(mai_mai_n51_), .B(mai_mai_n17_), .Y(mai_mai_n107_));
  NA2        m091(.A(mai_mai_n40_), .B(x0), .Y(mai_mai_n108_));
  OAI210     m092(.A0(x9), .A1(mai_mai_n107_), .B0(mai_mai_n108_), .Y(mai_mai_n109_));
  AOI220     m093(.A0(mai_mai_n109_), .A1(mai_mai_n106_), .B0(mai_mai_n105_), .B1(x4), .Y(mai_mai_n110_));
  NO3        m094(.A(mai_mai_n110_), .B(x7), .C(x5), .Y(mai_mai_n111_));
  OR2        m095(.A(x8), .B(x0), .Y(mai_mai_n112_));
  INV        m096(.A(mai_mai_n112_), .Y(mai_mai_n113_));
  NAi21      m097(.An(x2), .B(x8), .Y(mai_mai_n114_));
  INV        m098(.A(mai_mai_n114_), .Y(mai_mai_n115_));
  NO2        m099(.A(mai_mai_n115_), .B(mai_mai_n113_), .Y(mai_mai_n116_));
  NO2        m100(.A(x4), .B(x1), .Y(mai_mai_n117_));
  NA3        m101(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(mai_mai_n57_), .Y(mai_mai_n118_));
  NOi21      m102(.An(x0), .B(x1), .Y(mai_mai_n119_));
  NO3        m103(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n120_));
  NOi21      m104(.An(x0), .B(x4), .Y(mai_mai_n121_));
  NO2        m105(.A(mai_mai_n118_), .B(mai_mai_n74_), .Y(mai_mai_n122_));
  NO2        m106(.A(x5), .B(mai_mai_n45_), .Y(mai_mai_n123_));
  NA2        m107(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n124_));
  AOI210     m108(.A0(mai_mai_n124_), .A1(mai_mai_n101_), .B0(mai_mai_n108_), .Y(mai_mai_n125_));
  OAI210     m109(.A0(mai_mai_n125_), .A1(mai_mai_n32_), .B0(mai_mai_n123_), .Y(mai_mai_n126_));
  NAi21      m110(.An(x0), .B(x4), .Y(mai_mai_n127_));
  NO2        m111(.A(mai_mai_n127_), .B(x1), .Y(mai_mai_n128_));
  NO2        m112(.A(x7), .B(x0), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n79_), .B(mai_mai_n95_), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n130_), .B(x3), .Y(mai_mai_n131_));
  OAI210     m115(.A0(mai_mai_n129_), .A1(mai_mai_n128_), .B0(mai_mai_n131_), .Y(mai_mai_n132_));
  NA2        m116(.A(x5), .B(x0), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n134_));
  NA3        m118(.A(mai_mai_n132_), .B(mai_mai_n126_), .C(mai_mai_n33_), .Y(mai_mai_n135_));
  NO3        m119(.A(mai_mai_n135_), .B(mai_mai_n122_), .C(mai_mai_n111_), .Y(mai_mai_n136_));
  NO3        m120(.A(mai_mai_n74_), .B(mai_mai_n72_), .C(mai_mai_n23_), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n27_), .B(mai_mai_n24_), .Y(mai_mai_n138_));
  NA2        m122(.A(x7), .B(x3), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n94_), .B(x5), .Y(mai_mai_n140_));
  NO2        m124(.A(x9), .B(x7), .Y(mai_mai_n141_));
  NOi21      m125(.An(x8), .B(x0), .Y(mai_mai_n142_));
  OA210      m126(.A0(mai_mai_n141_), .A1(x1), .B0(mai_mai_n142_), .Y(mai_mai_n143_));
  NO2        m127(.A(mai_mai_n40_), .B(x2), .Y(mai_mai_n144_));
  INV        m128(.A(x7), .Y(mai_mai_n145_));
  NA2        m129(.A(mai_mai_n145_), .B(mai_mai_n18_), .Y(mai_mai_n146_));
  AOI220     m130(.A0(mai_mai_n146_), .A1(mai_mai_n144_), .B0(mai_mai_n105_), .B1(mai_mai_n35_), .Y(mai_mai_n147_));
  NO2        m131(.A(mai_mai_n24_), .B(x4), .Y(mai_mai_n148_));
  NO2        m132(.A(mai_mai_n148_), .B(mai_mai_n121_), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n149_), .B(mai_mai_n147_), .Y(mai_mai_n150_));
  AOI210     m134(.A0(mai_mai_n143_), .A1(mai_mai_n140_), .B0(mai_mai_n150_), .Y(mai_mai_n151_));
  OAI210     m135(.A0(mai_mai_n139_), .A1(mai_mai_n47_), .B0(mai_mai_n151_), .Y(mai_mai_n152_));
  NA2        m136(.A(x5), .B(x1), .Y(mai_mai_n153_));
  INV        m137(.A(mai_mai_n153_), .Y(mai_mai_n154_));
  AOI210     m138(.A0(mai_mai_n154_), .A1(mai_mai_n121_), .B0(mai_mai_n33_), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n59_), .B(mai_mai_n87_), .Y(mai_mai_n156_));
  NAi21      m140(.An(x2), .B(x7), .Y(mai_mai_n157_));
  NO3        m141(.A(mai_mai_n157_), .B(mai_mai_n156_), .C(mai_mai_n45_), .Y(mai_mai_n158_));
  NA2        m142(.A(mai_mai_n158_), .B(mai_mai_n64_), .Y(mai_mai_n159_));
  NAi31      m143(.An(mai_mai_n74_), .B(mai_mai_n35_), .C(mai_mai_n32_), .Y(mai_mai_n160_));
  NA3        m144(.A(mai_mai_n160_), .B(mai_mai_n159_), .C(mai_mai_n155_), .Y(mai_mai_n161_));
  NO3        m145(.A(mai_mai_n161_), .B(mai_mai_n152_), .C(mai_mai_n137_), .Y(mai_mai_n162_));
  NO2        m146(.A(mai_mai_n162_), .B(mai_mai_n136_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n133_), .B(mai_mai_n130_), .Y(mai_mai_n164_));
  NA2        m148(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n165_));
  NA2        m149(.A(mai_mai_n24_), .B(mai_mai_n17_), .Y(mai_mai_n166_));
  NA3        m150(.A(mai_mai_n166_), .B(mai_mai_n165_), .C(mai_mai_n23_), .Y(mai_mai_n167_));
  AN2        m151(.A(mai_mai_n167_), .B(mai_mai_n134_), .Y(mai_mai_n168_));
  NA2        m152(.A(x8), .B(x0), .Y(mai_mai_n169_));
  NO2        m153(.A(mai_mai_n145_), .B(mai_mai_n24_), .Y(mai_mai_n170_));
  NO2        m154(.A(mai_mai_n119_), .B(x4), .Y(mai_mai_n171_));
  NA2        m155(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  AOI210     m156(.A0(mai_mai_n169_), .A1(mai_mai_n124_), .B0(mai_mai_n172_), .Y(mai_mai_n173_));
  NA2        m157(.A(x2), .B(x0), .Y(mai_mai_n174_));
  NA2        m158(.A(x4), .B(x1), .Y(mai_mai_n175_));
  NAi21      m159(.An(mai_mai_n117_), .B(mai_mai_n175_), .Y(mai_mai_n176_));
  NOi31      m160(.An(mai_mai_n176_), .B(mai_mai_n148_), .C(mai_mai_n174_), .Y(mai_mai_n177_));
  NO4        m161(.A(mai_mai_n177_), .B(mai_mai_n173_), .C(mai_mai_n168_), .D(mai_mai_n164_), .Y(mai_mai_n178_));
  NO2        m162(.A(mai_mai_n178_), .B(mai_mai_n40_), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n167_), .B(mai_mai_n72_), .Y(mai_mai_n180_));
  INV        m164(.A(mai_mai_n123_), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n101_), .B(mai_mai_n17_), .Y(mai_mai_n182_));
  AOI210     m166(.A0(mai_mai_n32_), .A1(mai_mai_n87_), .B0(mai_mai_n182_), .Y(mai_mai_n183_));
  NO3        m167(.A(mai_mai_n183_), .B(mai_mai_n181_), .C(x7), .Y(mai_mai_n184_));
  NA3        m168(.A(mai_mai_n176_), .B(mai_mai_n181_), .C(mai_mai_n39_), .Y(mai_mai_n185_));
  OAI210     m169(.A0(mai_mai_n166_), .A1(mai_mai_n130_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  NO3        m170(.A(mai_mai_n186_), .B(mai_mai_n184_), .C(mai_mai_n180_), .Y(mai_mai_n187_));
  NO2        m171(.A(mai_mai_n187_), .B(x3), .Y(mai_mai_n188_));
  NO3        m172(.A(mai_mai_n188_), .B(mai_mai_n179_), .C(mai_mai_n163_), .Y(mai03));
  NO2        m173(.A(mai_mai_n45_), .B(x3), .Y(mai_mai_n190_));
  NO2        m174(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n191_));
  INV        m175(.A(mai_mai_n191_), .Y(mai_mai_n192_));
  NO2        m176(.A(mai_mai_n51_), .B(x1), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n192_), .B(mai_mai_n101_), .Y(mai_mai_n194_));
  NA2        m178(.A(mai_mai_n194_), .B(mai_mai_n190_), .Y(mai_mai_n195_));
  NO2        m179(.A(mai_mai_n74_), .B(x6), .Y(mai_mai_n196_));
  NA2        m180(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n197_));
  NO2        m181(.A(mai_mai_n197_), .B(x4), .Y(mai_mai_n198_));
  NO2        m182(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n199_));
  AO220      m183(.A0(mai_mai_n199_), .A1(mai_mai_n198_), .B0(mai_mai_n196_), .B1(mai_mai_n52_), .Y(mai_mai_n200_));
  INV        m184(.A(mai_mai_n200_), .Y(mai_mai_n201_));
  NA2        m185(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n202_));
  NO2        m186(.A(mai_mai_n202_), .B(mai_mai_n197_), .Y(mai_mai_n203_));
  NA2        m187(.A(x9), .B(mai_mai_n51_), .Y(mai_mai_n204_));
  INV        m188(.A(mai_mai_n197_), .Y(mai_mai_n205_));
  AOI210     m189(.A0(mai_mai_n24_), .A1(x3), .B0(mai_mai_n174_), .Y(mai_mai_n206_));
  AOI220     m190(.A0(mai_mai_n206_), .A1(mai_mai_n205_), .B0(x9), .B1(mai_mai_n203_), .Y(mai_mai_n207_));
  NO3        m191(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n208_));
  NO2        m192(.A(x5), .B(x1), .Y(mai_mai_n209_));
  AOI220     m193(.A0(mai_mai_n209_), .A1(mai_mai_n17_), .B0(mai_mai_n98_), .B1(x5), .Y(mai_mai_n210_));
  NO2        m194(.A(mai_mai_n202_), .B(mai_mai_n165_), .Y(mai_mai_n211_));
  NO3        m195(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n212_));
  NO2        m196(.A(mai_mai_n212_), .B(mai_mai_n211_), .Y(mai_mai_n213_));
  OAI210     m197(.A0(mai_mai_n210_), .A1(mai_mai_n61_), .B0(mai_mai_n213_), .Y(mai_mai_n214_));
  AOI220     m198(.A0(mai_mai_n214_), .A1(mai_mai_n45_), .B0(mai_mai_n208_), .B1(mai_mai_n123_), .Y(mai_mai_n215_));
  NA4        m199(.A(mai_mai_n215_), .B(mai_mai_n207_), .C(mai_mai_n201_), .D(mai_mai_n195_), .Y(mai_mai_n216_));
  NO2        m200(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n217_));
  NA2        m201(.A(mai_mai_n217_), .B(mai_mai_n19_), .Y(mai_mai_n218_));
  NO2        m202(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n219_));
  NO2        m203(.A(mai_mai_n219_), .B(x6), .Y(mai_mai_n220_));
  NOi21      m204(.An(mai_mai_n79_), .B(mai_mai_n220_), .Y(mai_mai_n221_));
  NA2        m205(.A(mai_mai_n59_), .B(mai_mai_n87_), .Y(mai_mai_n222_));
  NA3        m206(.A(mai_mai_n222_), .B(mai_mai_n219_), .C(x6), .Y(mai_mai_n223_));
  AOI210     m207(.A0(mai_mai_n223_), .A1(mai_mai_n221_), .B0(mai_mai_n145_), .Y(mai_mai_n224_));
  OR2        m208(.A(mai_mai_n224_), .B(mai_mai_n170_), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n40_), .B(mai_mai_n51_), .Y(mai_mai_n226_));
  NA2        m210(.A(mai_mai_n134_), .B(mai_mai_n86_), .Y(mai_mai_n227_));
  NA2        m211(.A(x6), .B(mai_mai_n45_), .Y(mai_mai_n228_));
  OAI210     m212(.A0(mai_mai_n113_), .A1(mai_mai_n75_), .B0(x4), .Y(mai_mai_n229_));
  AOI210     m213(.A0(mai_mai_n229_), .A1(mai_mai_n228_), .B0(mai_mai_n74_), .Y(mai_mai_n230_));
  NA2        m214(.A(mai_mai_n191_), .B(mai_mai_n128_), .Y(mai_mai_n231_));
  NA3        m215(.A(mai_mai_n202_), .B(mai_mai_n123_), .C(x6), .Y(mai_mai_n232_));
  OAI210     m216(.A0(mai_mai_n87_), .A1(mai_mai_n33_), .B0(mai_mai_n64_), .Y(mai_mai_n233_));
  NA3        m217(.A(mai_mai_n233_), .B(mai_mai_n232_), .C(mai_mai_n231_), .Y(mai_mai_n234_));
  OAI210     m218(.A0(mai_mai_n234_), .A1(mai_mai_n230_), .B0(x2), .Y(mai_mai_n235_));
  NA3        m219(.A(mai_mai_n235_), .B(mai_mai_n227_), .C(mai_mai_n225_), .Y(mai_mai_n236_));
  AOI210     m220(.A0(mai_mai_n216_), .A1(x8), .B0(mai_mai_n236_), .Y(mai_mai_n237_));
  NO2        m221(.A(mai_mai_n87_), .B(x3), .Y(mai_mai_n238_));
  NA2        m222(.A(mai_mai_n238_), .B(mai_mai_n198_), .Y(mai_mai_n239_));
  NO3        m223(.A(mai_mai_n85_), .B(mai_mai_n75_), .C(mai_mai_n24_), .Y(mai_mai_n240_));
  AOI210     m224(.A0(mai_mai_n220_), .A1(mai_mai_n148_), .B0(mai_mai_n240_), .Y(mai_mai_n241_));
  AOI210     m225(.A0(mai_mai_n241_), .A1(mai_mai_n239_), .B0(x2), .Y(mai_mai_n242_));
  NO2        m226(.A(x4), .B(mai_mai_n51_), .Y(mai_mai_n243_));
  AOI220     m227(.A0(mai_mai_n198_), .A1(mai_mai_n182_), .B0(mai_mai_n243_), .B1(mai_mai_n64_), .Y(mai_mai_n244_));
  NA2        m228(.A(mai_mai_n59_), .B(x6), .Y(mai_mai_n245_));
  NA3        m229(.A(mai_mai_n24_), .B(x3), .C(x2), .Y(mai_mai_n246_));
  AOI210     m230(.A0(mai_mai_n246_), .A1(mai_mai_n133_), .B0(mai_mai_n245_), .Y(mai_mai_n247_));
  NA2        m231(.A(mai_mai_n40_), .B(mai_mai_n17_), .Y(mai_mai_n248_));
  NO2        m232(.A(mai_mai_n248_), .B(mai_mai_n24_), .Y(mai_mai_n249_));
  OAI210     m233(.A0(mai_mai_n249_), .A1(mai_mai_n247_), .B0(mai_mai_n117_), .Y(mai_mai_n250_));
  NA2        m234(.A(mai_mai_n202_), .B(x6), .Y(mai_mai_n251_));
  NO2        m235(.A(mai_mai_n202_), .B(x6), .Y(mai_mai_n252_));
  NAi21      m236(.An(mai_mai_n156_), .B(mai_mai_n252_), .Y(mai_mai_n253_));
  NA3        m237(.A(mai_mai_n253_), .B(mai_mai_n251_), .C(mai_mai_n138_), .Y(mai_mai_n254_));
  NA4        m238(.A(mai_mai_n254_), .B(mai_mai_n250_), .C(mai_mai_n244_), .D(mai_mai_n145_), .Y(mai_mai_n255_));
  NO2        m239(.A(x9), .B(x6), .Y(mai_mai_n256_));
  NO2        m240(.A(mai_mai_n133_), .B(mai_mai_n18_), .Y(mai_mai_n257_));
  NAi21      m241(.An(mai_mai_n257_), .B(mai_mai_n246_), .Y(mai_mai_n258_));
  NAi21      m242(.An(x1), .B(x4), .Y(mai_mai_n259_));
  AOI210     m243(.A0(x3), .A1(x2), .B0(mai_mai_n45_), .Y(mai_mai_n260_));
  OAI210     m244(.A0(mai_mai_n133_), .A1(x3), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  AOI220     m245(.A0(mai_mai_n261_), .A1(mai_mai_n259_), .B0(mai_mai_n258_), .B1(mai_mai_n256_), .Y(mai_mai_n262_));
  INV        m246(.A(mai_mai_n262_), .Y(mai_mai_n263_));
  NO3        m247(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n264_));
  NA2        m248(.A(mai_mai_n101_), .B(mai_mai_n24_), .Y(mai_mai_n265_));
  NA2        m249(.A(x6), .B(x2), .Y(mai_mai_n266_));
  NO2        m250(.A(mai_mai_n266_), .B(mai_mai_n165_), .Y(mai_mai_n267_));
  AOI210     m251(.A0(mai_mai_n265_), .A1(mai_mai_n264_), .B0(mai_mai_n267_), .Y(mai_mai_n268_));
  OAI220     m252(.A0(mai_mai_n268_), .A1(mai_mai_n40_), .B0(mai_mai_n171_), .B1(mai_mai_n43_), .Y(mai_mai_n269_));
  NA2        m253(.A(mai_mai_n269_), .B(mai_mai_n263_), .Y(mai_mai_n270_));
  OR2        m254(.A(mai_mai_n196_), .B(mai_mai_n140_), .Y(mai_mai_n271_));
  NA2        m255(.A(x4), .B(x0), .Y(mai_mai_n272_));
  NO3        m256(.A(mai_mai_n69_), .B(mai_mai_n272_), .C(x6), .Y(mai_mai_n273_));
  AOI210     m257(.A0(mai_mai_n271_), .A1(mai_mai_n39_), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  AOI210     m258(.A0(mai_mai_n274_), .A1(mai_mai_n270_), .B0(x8), .Y(mai_mai_n275_));
  INV        m259(.A(mai_mai_n245_), .Y(mai_mai_n276_));
  OAI210     m260(.A0(mai_mai_n257_), .A1(mai_mai_n209_), .B0(mai_mai_n276_), .Y(mai_mai_n277_));
  OAI210     m261(.A0(x0), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n278_));
  AOI210     m262(.A0(mai_mai_n278_), .A1(mai_mai_n277_), .B0(mai_mai_n226_), .Y(mai_mai_n279_));
  NO4        m263(.A(mai_mai_n279_), .B(mai_mai_n275_), .C(mai_mai_n255_), .D(mai_mai_n242_), .Y(mai_mai_n280_));
  NO2        m264(.A(mai_mai_n156_), .B(x1), .Y(mai_mai_n281_));
  NO3        m265(.A(mai_mai_n281_), .B(x3), .C(mai_mai_n33_), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n282_), .A1(mai_mai_n252_), .B0(x2), .Y(mai_mai_n283_));
  OAI210     m267(.A0(x0), .A1(x6), .B0(mai_mai_n41_), .Y(mai_mai_n284_));
  AOI210     m268(.A0(mai_mai_n284_), .A1(mai_mai_n283_), .B0(mai_mai_n181_), .Y(mai_mai_n285_));
  NOi21      m269(.An(mai_mai_n266_), .B(mai_mai_n17_), .Y(mai_mai_n286_));
  NA3        m270(.A(mai_mai_n286_), .B(mai_mai_n209_), .C(mai_mai_n37_), .Y(mai_mai_n287_));
  AOI210     m271(.A0(mai_mai_n33_), .A1(mai_mai_n51_), .B0(x0), .Y(mai_mai_n288_));
  NA3        m272(.A(mai_mai_n288_), .B(mai_mai_n154_), .C(mai_mai_n30_), .Y(mai_mai_n289_));
  NA2        m273(.A(x3), .B(x2), .Y(mai_mai_n290_));
  AOI220     m274(.A0(mai_mai_n290_), .A1(mai_mai_n226_), .B0(mai_mai_n289_), .B1(mai_mai_n287_), .Y(mai_mai_n291_));
  NAi21      m275(.An(x4), .B(x0), .Y(mai_mai_n292_));
  NO3        m276(.A(mai_mai_n292_), .B(mai_mai_n41_), .C(x2), .Y(mai_mai_n293_));
  OAI210     m277(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n293_), .Y(mai_mai_n294_));
  OAI220     m278(.A0(mai_mai_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n295_));
  NO2        m279(.A(mai_mai_n288_), .B(mai_mai_n286_), .Y(mai_mai_n296_));
  AOI220     m280(.A0(mai_mai_n296_), .A1(mai_mai_n78_), .B0(mai_mai_n295_), .B1(mai_mai_n29_), .Y(mai_mai_n297_));
  AOI210     m281(.A0(mai_mai_n297_), .A1(mai_mai_n294_), .B0(mai_mai_n24_), .Y(mai_mai_n298_));
  NA3        m282(.A(mai_mai_n33_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n299_));
  OAI210     m283(.A0(mai_mai_n288_), .A1(mai_mai_n286_), .B0(mai_mai_n299_), .Y(mai_mai_n300_));
  INV        m284(.A(mai_mai_n211_), .Y(mai_mai_n301_));
  NA2        m285(.A(mai_mai_n33_), .B(mai_mai_n40_), .Y(mai_mai_n302_));
  OR2        m286(.A(mai_mai_n302_), .B(mai_mai_n272_), .Y(mai_mai_n303_));
  OAI220     m287(.A0(mai_mai_n303_), .A1(mai_mai_n153_), .B0(mai_mai_n228_), .B1(mai_mai_n301_), .Y(mai_mai_n304_));
  AO210      m288(.A0(mai_mai_n300_), .A1(mai_mai_n140_), .B0(mai_mai_n304_), .Y(mai_mai_n305_));
  NO4        m289(.A(mai_mai_n305_), .B(mai_mai_n298_), .C(mai_mai_n291_), .D(mai_mai_n285_), .Y(mai_mai_n306_));
  OAI210     m290(.A0(mai_mai_n280_), .A1(mai_mai_n237_), .B0(mai_mai_n306_), .Y(mai04));
  OAI210     m291(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n308_));
  NA3        m292(.A(mai_mai_n308_), .B(mai_mai_n264_), .C(mai_mai_n80_), .Y(mai_mai_n309_));
  NO2        m293(.A(x2), .B(x1), .Y(mai_mai_n310_));
  OAI210     m294(.A0(mai_mai_n248_), .A1(mai_mai_n310_), .B0(mai_mai_n33_), .Y(mai_mai_n311_));
  NO2        m295(.A(mai_mai_n310_), .B(mai_mai_n292_), .Y(mai_mai_n312_));
  AOI210     m296(.A0(mai_mai_n59_), .A1(x4), .B0(mai_mai_n107_), .Y(mai_mai_n313_));
  OAI210     m297(.A0(mai_mai_n313_), .A1(mai_mai_n312_), .B0(mai_mai_n238_), .Y(mai_mai_n314_));
  NO2        m298(.A(mai_mai_n444_), .B(mai_mai_n85_), .Y(mai_mai_n315_));
  NO2        m299(.A(mai_mai_n315_), .B(mai_mai_n33_), .Y(mai_mai_n316_));
  NO2        m300(.A(mai_mai_n290_), .B(mai_mai_n199_), .Y(mai_mai_n317_));
  NA2        m301(.A(x9), .B(x0), .Y(mai_mai_n318_));
  AOI210     m302(.A0(mai_mai_n85_), .A1(mai_mai_n72_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  OAI210     m303(.A0(mai_mai_n319_), .A1(mai_mai_n317_), .B0(mai_mai_n87_), .Y(mai_mai_n320_));
  NA3        m304(.A(mai_mai_n320_), .B(mai_mai_n316_), .C(mai_mai_n314_), .Y(mai_mai_n321_));
  NA2        m305(.A(mai_mai_n321_), .B(mai_mai_n311_), .Y(mai_mai_n322_));
  NO2        m306(.A(mai_mai_n204_), .B(mai_mai_n108_), .Y(mai_mai_n323_));
  NO3        m307(.A(mai_mai_n245_), .B(mai_mai_n114_), .C(mai_mai_n18_), .Y(mai_mai_n324_));
  NO2        m308(.A(mai_mai_n324_), .B(mai_mai_n323_), .Y(mai_mai_n325_));
  NOi21      m309(.An(mai_mai_n142_), .B(mai_mai_n124_), .Y(mai_mai_n326_));
  AOI210     m310(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n327_));
  OAI220     m311(.A0(mai_mai_n327_), .A1(mai_mai_n302_), .B0(mai_mai_n444_), .B1(mai_mai_n299_), .Y(mai_mai_n328_));
  AOI210     m312(.A0(mai_mai_n326_), .A1(mai_mai_n60_), .B0(mai_mai_n328_), .Y(mai_mai_n329_));
  NA2        m313(.A(mai_mai_n315_), .B(mai_mai_n87_), .Y(mai_mai_n330_));
  NA3        m314(.A(mai_mai_n330_), .B(mai_mai_n329_), .C(mai_mai_n325_), .Y(mai_mai_n331_));
  OAI210     m315(.A0(mai_mai_n106_), .A1(x3), .B0(mai_mai_n293_), .Y(mai_mai_n332_));
  NA3        m316(.A(mai_mai_n222_), .B(mai_mai_n208_), .C(mai_mai_n79_), .Y(mai_mai_n333_));
  NA3        m317(.A(mai_mai_n333_), .B(mai_mai_n332_), .C(mai_mai_n145_), .Y(mai_mai_n334_));
  AOI210     m318(.A0(mai_mai_n331_), .A1(x4), .B0(mai_mai_n334_), .Y(mai_mai_n335_));
  NA3        m319(.A(mai_mai_n312_), .B(mai_mai_n204_), .C(mai_mai_n87_), .Y(mai_mai_n336_));
  NOi21      m320(.An(x4), .B(x0), .Y(mai_mai_n337_));
  XO2        m321(.A(x4), .B(x0), .Y(mai_mai_n338_));
  NA2        m322(.A(mai_mai_n337_), .B(mai_mai_n88_), .Y(mai_mai_n339_));
  AOI210     m323(.A0(mai_mai_n339_), .A1(mai_mai_n336_), .B0(x3), .Y(mai_mai_n340_));
  INV        m324(.A(mai_mai_n88_), .Y(mai_mai_n341_));
  NO2        m325(.A(mai_mai_n87_), .B(x4), .Y(mai_mai_n342_));
  AOI220     m326(.A0(mai_mai_n342_), .A1(mai_mai_n41_), .B0(mai_mai_n121_), .B1(mai_mai_n341_), .Y(mai_mai_n343_));
  NO3        m327(.A(mai_mai_n338_), .B(mai_mai_n156_), .C(x2), .Y(mai_mai_n344_));
  NO3        m328(.A(mai_mai_n222_), .B(mai_mai_n27_), .C(mai_mai_n23_), .Y(mai_mai_n345_));
  NO2        m329(.A(mai_mai_n345_), .B(mai_mai_n344_), .Y(mai_mai_n346_));
  NA4        m330(.A(mai_mai_n346_), .B(mai_mai_n343_), .C(mai_mai_n218_), .D(x6), .Y(mai_mai_n347_));
  NO2        m331(.A(mai_mai_n174_), .B(mai_mai_n87_), .Y(mai_mai_n348_));
  NO2        m332(.A(mai_mai_n40_), .B(x0), .Y(mai_mai_n349_));
  NA2        m333(.A(mai_mai_n348_), .B(mai_mai_n58_), .Y(mai_mai_n350_));
  NO2        m334(.A(mai_mai_n142_), .B(mai_mai_n77_), .Y(mai_mai_n351_));
  NO2        m335(.A(mai_mai_n32_), .B(x2), .Y(mai_mai_n352_));
  NA2        m336(.A(mai_mai_n352_), .B(mai_mai_n351_), .Y(mai_mai_n353_));
  NA2        m337(.A(mai_mai_n350_), .B(mai_mai_n353_), .Y(mai_mai_n354_));
  OAI220     m338(.A0(mai_mai_n354_), .A1(x6), .B0(mai_mai_n347_), .B1(mai_mai_n340_), .Y(mai_mai_n355_));
  OAI210     m339(.A0(mai_mai_n60_), .A1(mai_mai_n45_), .B0(mai_mai_n39_), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n356_), .A1(mai_mai_n87_), .B0(mai_mai_n303_), .Y(mai_mai_n357_));
  AOI210     m341(.A0(mai_mai_n357_), .A1(mai_mai_n18_), .B0(mai_mai_n145_), .Y(mai_mai_n358_));
  AO220      m342(.A0(mai_mai_n358_), .A1(mai_mai_n355_), .B0(mai_mai_n335_), .B1(mai_mai_n322_), .Y(mai_mai_n359_));
  NA2        m343(.A(mai_mai_n352_), .B(x6), .Y(mai_mai_n360_));
  AOI210     m344(.A0(x6), .A1(x1), .B0(mai_mai_n144_), .Y(mai_mai_n361_));
  NA2        m345(.A(mai_mai_n342_), .B(x0), .Y(mai_mai_n362_));
  NA2        m346(.A(mai_mai_n79_), .B(x6), .Y(mai_mai_n363_));
  OAI210     m347(.A0(mai_mai_n362_), .A1(mai_mai_n361_), .B0(mai_mai_n363_), .Y(mai_mai_n364_));
  AOI220     m348(.A0(mai_mai_n364_), .A1(mai_mai_n360_), .B0(mai_mai_n212_), .B1(mai_mai_n46_), .Y(mai_mai_n365_));
  NA3        m349(.A(mai_mai_n365_), .B(mai_mai_n359_), .C(mai_mai_n309_), .Y(mai_mai_n366_));
  OAI210     m350(.A0(mai_mai_n27_), .A1(x1), .B0(mai_mai_n226_), .Y(mai_mai_n367_));
  AO220      m351(.A0(mai_mai_n367_), .A1(mai_mai_n141_), .B0(mai_mai_n105_), .B1(x4), .Y(mai_mai_n368_));
  NA3        m352(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n369_));
  NO2        m353(.A(mai_mai_n369_), .B(mai_mai_n341_), .Y(mai_mai_n370_));
  AOI210     m354(.A0(mai_mai_n368_), .A1(mai_mai_n113_), .B0(mai_mai_n370_), .Y(mai_mai_n371_));
  NO2        m355(.A(mai_mai_n371_), .B(mai_mai_n24_), .Y(mai_mai_n372_));
  NA3        m356(.A(mai_mai_n115_), .B(mai_mai_n217_), .C(x0), .Y(mai_mai_n373_));
  OAI210     m357(.A0(mai_mai_n190_), .A1(mai_mai_n65_), .B0(mai_mai_n199_), .Y(mai_mai_n374_));
  NA3        m358(.A(mai_mai_n193_), .B(mai_mai_n219_), .C(x8), .Y(mai_mai_n375_));
  AOI210     m359(.A0(mai_mai_n375_), .A1(mai_mai_n374_), .B0(mai_mai_n24_), .Y(mai_mai_n376_));
  AOI210     m360(.A0(mai_mai_n114_), .A1(mai_mai_n112_), .B0(mai_mai_n39_), .Y(mai_mai_n377_));
  NOi31      m361(.An(mai_mai_n377_), .B(mai_mai_n349_), .C(mai_mai_n175_), .Y(mai_mai_n378_));
  OAI210     m362(.A0(mai_mai_n378_), .A1(mai_mai_n376_), .B0(mai_mai_n141_), .Y(mai_mai_n379_));
  NAi31      m363(.An(mai_mai_n47_), .B(mai_mai_n281_), .C(mai_mai_n170_), .Y(mai_mai_n380_));
  NA3        m364(.A(mai_mai_n380_), .B(mai_mai_n379_), .C(mai_mai_n373_), .Y(mai_mai_n381_));
  OAI210     m365(.A0(mai_mai_n381_), .A1(mai_mai_n372_), .B0(x6), .Y(mai_mai_n382_));
  OAI210     m366(.A0(mai_mai_n156_), .A1(mai_mai_n45_), .B0(mai_mai_n129_), .Y(mai_mai_n383_));
  NA2        m367(.A(mai_mai_n52_), .B(mai_mai_n35_), .Y(mai_mai_n384_));
  AOI220     m368(.A0(mai_mai_n384_), .A1(mai_mai_n383_), .B0(mai_mai_n37_), .B1(mai_mai_n30_), .Y(mai_mai_n385_));
  NO2        m369(.A(mai_mai_n145_), .B(x0), .Y(mai_mai_n386_));
  AOI220     m370(.A0(mai_mai_n386_), .A1(mai_mai_n217_), .B0(mai_mai_n190_), .B1(mai_mai_n145_), .Y(mai_mai_n387_));
  INV        m371(.A(x1), .Y(mai_mai_n388_));
  OAI210     m372(.A0(mai_mai_n387_), .A1(x8), .B0(mai_mai_n388_), .Y(mai_mai_n389_));
  NAi31      m373(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n390_));
  OAI210     m374(.A0(mai_mai_n390_), .A1(x4), .B0(mai_mai_n157_), .Y(mai_mai_n391_));
  NA3        m375(.A(mai_mai_n391_), .B(mai_mai_n139_), .C(x9), .Y(mai_mai_n392_));
  NA2        m376(.A(mai_mai_n351_), .B(mai_mai_n145_), .Y(mai_mai_n393_));
  NA4        m377(.A(mai_mai_n393_), .B(x1), .C(mai_mai_n392_), .D(mai_mai_n47_), .Y(mai_mai_n394_));
  OAI210     m378(.A0(mai_mai_n389_), .A1(mai_mai_n385_), .B0(mai_mai_n394_), .Y(mai_mai_n395_));
  NOi31      m379(.An(mai_mai_n386_), .B(mai_mai_n30_), .C(x8), .Y(mai_mai_n396_));
  AOI210     m380(.A0(mai_mai_n35_), .A1(x9), .B0(mai_mai_n127_), .Y(mai_mai_n397_));
  NO3        m381(.A(mai_mai_n397_), .B(mai_mai_n120_), .C(mai_mai_n40_), .Y(mai_mai_n398_));
  NOi31      m382(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n399_));
  AOI220     m383(.A0(mai_mai_n399_), .A1(mai_mai_n337_), .B0(mai_mai_n121_), .B1(x3), .Y(mai_mai_n400_));
  AOI210     m384(.A0(mai_mai_n259_), .A1(mai_mai_n57_), .B0(mai_mai_n119_), .Y(mai_mai_n401_));
  OAI210     m385(.A0(mai_mai_n401_), .A1(x3), .B0(mai_mai_n400_), .Y(mai_mai_n402_));
  NO3        m386(.A(mai_mai_n402_), .B(mai_mai_n398_), .C(x2), .Y(mai_mai_n403_));
  OAI210     m387(.A0(mai_mai_n292_), .A1(mai_mai_n40_), .B0(mai_mai_n338_), .Y(mai_mai_n404_));
  INV        m388(.A(mai_mai_n369_), .Y(mai_mai_n405_));
  AOI220     m389(.A0(mai_mai_n405_), .A1(mai_mai_n87_), .B0(mai_mai_n404_), .B1(mai_mai_n145_), .Y(mai_mai_n406_));
  NO2        m390(.A(mai_mai_n406_), .B(mai_mai_n51_), .Y(mai_mai_n407_));
  NO3        m391(.A(mai_mai_n407_), .B(mai_mai_n403_), .C(mai_mai_n396_), .Y(mai_mai_n408_));
  AOI210     m392(.A0(mai_mai_n408_), .A1(mai_mai_n395_), .B0(mai_mai_n24_), .Y(mai_mai_n409_));
  NO3        m393(.A(mai_mai_n59_), .B(x4), .C(x1), .Y(mai_mai_n410_));
  NO3        m394(.A(mai_mai_n65_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n411_));
  AOI220     m395(.A0(mai_mai_n411_), .A1(mai_mai_n260_), .B0(mai_mai_n410_), .B1(mai_mai_n377_), .Y(mai_mai_n412_));
  NO2        m396(.A(mai_mai_n412_), .B(mai_mai_n98_), .Y(mai_mai_n413_));
  NA2        m397(.A(mai_mai_n413_), .B(x7), .Y(mai_mai_n414_));
  NA2        m398(.A(mai_mai_n222_), .B(x7), .Y(mai_mai_n415_));
  NA3        m399(.A(mai_mai_n415_), .B(mai_mai_n144_), .C(mai_mai_n128_), .Y(mai_mai_n416_));
  NA2        m400(.A(mai_mai_n416_), .B(mai_mai_n414_), .Y(mai_mai_n417_));
  OAI210     m401(.A0(mai_mai_n417_), .A1(mai_mai_n409_), .B0(mai_mai_n33_), .Y(mai_mai_n418_));
  INV        m402(.A(mai_mai_n199_), .Y(mai_mai_n419_));
  NO4        m403(.A(mai_mai_n419_), .B(mai_mai_n74_), .C(x4), .D(mai_mai_n51_), .Y(mai_mai_n420_));
  NA2        m404(.A(mai_mai_n248_), .B(mai_mai_n21_), .Y(mai_mai_n421_));
  NO2        m405(.A(mai_mai_n153_), .B(mai_mai_n129_), .Y(mai_mai_n422_));
  NA2        m406(.A(mai_mai_n422_), .B(mai_mai_n421_), .Y(mai_mai_n423_));
  AOI210     m407(.A0(mai_mai_n423_), .A1(mai_mai_n160_), .B0(mai_mai_n27_), .Y(mai_mai_n424_));
  AOI220     m408(.A0(mai_mai_n349_), .A1(mai_mai_n87_), .B0(mai_mai_n142_), .B1(mai_mai_n193_), .Y(mai_mai_n425_));
  NA3        m409(.A(mai_mai_n425_), .B(mai_mai_n390_), .C(mai_mai_n85_), .Y(mai_mai_n426_));
  NA2        m410(.A(mai_mai_n426_), .B(mai_mai_n170_), .Y(mai_mai_n427_));
  NO2        m411(.A(mai_mai_n153_), .B(mai_mai_n40_), .Y(mai_mai_n428_));
  NA2        m412(.A(x3), .B(mai_mai_n51_), .Y(mai_mai_n429_));
  AOI210     m413(.A0(mai_mai_n157_), .A1(mai_mai_n26_), .B0(mai_mai_n69_), .Y(mai_mai_n430_));
  OAI210     m414(.A0(mai_mai_n141_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n431_));
  NO3        m415(.A(mai_mai_n399_), .B(x3), .C(mai_mai_n51_), .Y(mai_mai_n432_));
  AOI210     m416(.A0(mai_mai_n432_), .A1(mai_mai_n431_), .B0(mai_mai_n430_), .Y(mai_mai_n433_));
  OAI210     m417(.A0(mai_mai_n146_), .A1(mai_mai_n429_), .B0(mai_mai_n433_), .Y(mai_mai_n434_));
  AOI220     m418(.A0(mai_mai_n434_), .A1(x0), .B0(mai_mai_n428_), .B1(mai_mai_n129_), .Y(mai_mai_n435_));
  AOI210     m419(.A0(mai_mai_n435_), .A1(mai_mai_n427_), .B0(mai_mai_n228_), .Y(mai_mai_n436_));
  NA2        m420(.A(x9), .B(x5), .Y(mai_mai_n437_));
  NO4        m421(.A(mai_mai_n101_), .B(mai_mai_n437_), .C(mai_mai_n57_), .D(mai_mai_n30_), .Y(mai_mai_n438_));
  NO4        m422(.A(mai_mai_n438_), .B(mai_mai_n436_), .C(mai_mai_n424_), .D(mai_mai_n420_), .Y(mai_mai_n439_));
  NA3        m423(.A(mai_mai_n439_), .B(mai_mai_n418_), .C(mai_mai_n382_), .Y(mai_mai_n440_));
  AOI210     m424(.A0(mai_mai_n366_), .A1(mai_mai_n24_), .B0(mai_mai_n440_), .Y(mai05));
  INV        m425(.A(x2), .Y(mai_mai_n444_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  NO2        u022(.A(men_men_n23_), .B(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n37_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  AOI210     u033(.A0(men_men_n22_), .A1(men_men_n19_), .B0(men_men_n35_), .Y(men_men_n50_));
  INV        u034(.A(x2), .Y(men_men_n51_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n17_), .Y(men_men_n52_));
  NA2        u036(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n53_), .B(men_men_n52_), .Y(men_men_n54_));
  OAI210     u038(.A0(men_men_n50_), .A1(men_men_n32_), .B0(men_men_n54_), .Y(men_men_n55_));
  NO3        u039(.A(men_men_n55_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u040(.A(x8), .B(x7), .Y(men_men_n57_));
  NA2        u041(.A(men_men_n41_), .B(x1), .Y(men_men_n58_));
  INV        u042(.A(x9), .Y(men_men_n59_));
  NO2        u043(.A(men_men_n59_), .B(men_men_n36_), .Y(men_men_n60_));
  INV        u044(.A(men_men_n60_), .Y(men_men_n61_));
  NO3        u045(.A(men_men_n61_), .B(men_men_n58_), .C(men_men_n57_), .Y(men_men_n62_));
  NO2        u046(.A(x7), .B(x6), .Y(men_men_n63_));
  NO2        u047(.A(men_men_n58_), .B(x5), .Y(men_men_n64_));
  NO2        u048(.A(x8), .B(x2), .Y(men_men_n65_));
  INV        u049(.A(men_men_n65_), .Y(men_men_n66_));
  NO2        u050(.A(men_men_n66_), .B(x1), .Y(men_men_n67_));
  OA210      u051(.A0(men_men_n67_), .A1(men_men_n64_), .B0(men_men_n63_), .Y(men_men_n68_));
  OAI210     u052(.A0(men_men_n42_), .A1(men_men_n25_), .B0(men_men_n51_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n53_), .A1(men_men_n20_), .B0(men_men_n69_), .Y(men_men_n70_));
  NAi31      u054(.An(x1), .B(x9), .C(x5), .Y(men_men_n71_));
  OAI220     u055(.A0(men_men_n71_), .A1(men_men_n41_), .B0(men_men_n70_), .B1(men_men_n68_), .Y(men_men_n72_));
  OAI210     u056(.A0(men_men_n72_), .A1(men_men_n62_), .B0(x4), .Y(men_men_n73_));
  NA2        u057(.A(men_men_n46_), .B(x2), .Y(men_men_n74_));
  OAI210     u058(.A0(men_men_n74_), .A1(men_men_n53_), .B0(x0), .Y(men_men_n75_));
  NA2        u059(.A(x5), .B(x3), .Y(men_men_n76_));
  NO2        u060(.A(x8), .B(x6), .Y(men_men_n77_));
  NO4        u061(.A(men_men_n77_), .B(men_men_n76_), .C(men_men_n63_), .D(men_men_n51_), .Y(men_men_n78_));
  NAi21      u062(.An(x4), .B(x3), .Y(men_men_n79_));
  INV        u063(.A(men_men_n79_), .Y(men_men_n80_));
  NO2        u064(.A(men_men_n80_), .B(men_men_n22_), .Y(men_men_n81_));
  NO2        u065(.A(x4), .B(x2), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(x3), .Y(men_men_n83_));
  NO3        u067(.A(men_men_n83_), .B(men_men_n81_), .C(men_men_n18_), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n78_), .C(men_men_n75_), .Y(men_men_n85_));
  NO4        u069(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n86_));
  NA2        u070(.A(men_men_n59_), .B(men_men_n46_), .Y(men_men_n87_));
  INV        u071(.A(men_men_n87_), .Y(men_men_n88_));
  OAI210     u072(.A0(men_men_n86_), .A1(men_men_n64_), .B0(men_men_n88_), .Y(men_men_n89_));
  NA2        u073(.A(x3), .B(men_men_n18_), .Y(men_men_n90_));
  NO2        u074(.A(men_men_n90_), .B(men_men_n25_), .Y(men_men_n91_));
  INV        u075(.A(x8), .Y(men_men_n92_));
  NA2        u076(.A(x2), .B(x1), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n91_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n26_), .Y(men_men_n96_));
  AOI210     u080(.A0(men_men_n53_), .A1(men_men_n25_), .B0(men_men_n51_), .Y(men_men_n97_));
  OAI210     u081(.A0(men_men_n43_), .A1(men_men_n37_), .B0(men_men_n46_), .Y(men_men_n98_));
  NO3        u082(.A(men_men_n98_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n99_));
  NA2        u083(.A(x4), .B(men_men_n41_), .Y(men_men_n100_));
  NO2        u084(.A(men_men_n46_), .B(men_men_n51_), .Y(men_men_n101_));
  NO2        u085(.A(men_men_n100_), .B(x1), .Y(men_men_n102_));
  NO2        u086(.A(x3), .B(x2), .Y(men_men_n103_));
  NA3        u087(.A(men_men_n103_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n104_));
  AOI210     u088(.A0(x8), .A1(x6), .B0(men_men_n104_), .Y(men_men_n105_));
  NA2        u089(.A(men_men_n51_), .B(x1), .Y(men_men_n106_));
  OAI210     u090(.A0(men_men_n106_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n107_));
  NO4        u091(.A(men_men_n107_), .B(men_men_n105_), .C(men_men_n102_), .D(men_men_n99_), .Y(men_men_n108_));
  AO220      u092(.A0(men_men_n108_), .A1(men_men_n89_), .B0(men_men_n85_), .B1(men_men_n73_), .Y(men02));
  NO2        u093(.A(x3), .B(men_men_n51_), .Y(men_men_n110_));
  NO2        u094(.A(x8), .B(men_men_n18_), .Y(men_men_n111_));
  NA2        u095(.A(men_men_n51_), .B(men_men_n17_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n41_), .B(x0), .Y(men_men_n113_));
  OAI210     u097(.A0(men_men_n87_), .A1(men_men_n112_), .B0(men_men_n113_), .Y(men_men_n114_));
  AOI220     u098(.A0(men_men_n114_), .A1(men_men_n111_), .B0(men_men_n110_), .B1(x4), .Y(men_men_n115_));
  NO3        u099(.A(men_men_n115_), .B(x7), .C(x5), .Y(men_men_n116_));
  NA2        u100(.A(x9), .B(x2), .Y(men_men_n117_));
  OR2        u101(.A(x8), .B(x0), .Y(men_men_n118_));
  INV        u102(.A(men_men_n118_), .Y(men_men_n119_));
  NAi21      u103(.An(x2), .B(x8), .Y(men_men_n120_));
  INV        u104(.A(men_men_n120_), .Y(men_men_n121_));
  OAI220     u105(.A0(men_men_n121_), .A1(men_men_n119_), .B0(men_men_n117_), .B1(x7), .Y(men_men_n122_));
  NO2        u106(.A(x4), .B(x1), .Y(men_men_n123_));
  NA3        u107(.A(men_men_n123_), .B(men_men_n122_), .C(men_men_n57_), .Y(men_men_n124_));
  NOi21      u108(.An(x0), .B(x1), .Y(men_men_n125_));
  NO3        u109(.A(x9), .B(x8), .C(x7), .Y(men_men_n126_));
  NOi21      u110(.An(x0), .B(x4), .Y(men_men_n127_));
  NAi21      u111(.An(x8), .B(x7), .Y(men_men_n128_));
  NO2        u112(.A(men_men_n128_), .B(men_men_n59_), .Y(men_men_n129_));
  AOI220     u113(.A0(men_men_n129_), .A1(men_men_n127_), .B0(men_men_n126_), .B1(men_men_n125_), .Y(men_men_n130_));
  AOI210     u114(.A0(men_men_n130_), .A1(men_men_n124_), .B0(men_men_n76_), .Y(men_men_n131_));
  NO2        u115(.A(x5), .B(men_men_n46_), .Y(men_men_n132_));
  NA2        u116(.A(x2), .B(men_men_n18_), .Y(men_men_n133_));
  AOI210     u117(.A0(men_men_n133_), .A1(men_men_n106_), .B0(men_men_n113_), .Y(men_men_n134_));
  OAI210     u118(.A0(men_men_n134_), .A1(men_men_n35_), .B0(men_men_n132_), .Y(men_men_n135_));
  NAi21      u119(.An(x0), .B(x4), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n136_), .B(x1), .Y(men_men_n137_));
  NO2        u121(.A(x7), .B(x0), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n82_), .B(men_men_n101_), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n139_), .B(x3), .Y(men_men_n140_));
  OAI210     u124(.A0(men_men_n138_), .A1(men_men_n137_), .B0(men_men_n140_), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n21_), .B(men_men_n41_), .Y(men_men_n142_));
  NA2        u126(.A(x5), .B(x0), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n46_), .B(x2), .Y(men_men_n144_));
  NA3        u128(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n142_), .Y(men_men_n145_));
  NA4        u129(.A(men_men_n145_), .B(men_men_n141_), .C(men_men_n135_), .D(men_men_n36_), .Y(men_men_n146_));
  NO3        u130(.A(men_men_n146_), .B(men_men_n131_), .C(men_men_n116_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n76_), .B(men_men_n74_), .C(men_men_n24_), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n149_));
  AOI220     u133(.A0(men_men_n125_), .A1(men_men_n149_), .B0(men_men_n64_), .B1(men_men_n17_), .Y(men_men_n150_));
  NO3        u134(.A(men_men_n150_), .B(men_men_n57_), .C(men_men_n59_), .Y(men_men_n151_));
  NA2        u135(.A(x7), .B(x3), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n100_), .B(x5), .Y(men_men_n153_));
  NO2        u137(.A(x9), .B(x7), .Y(men_men_n154_));
  NOi21      u138(.An(x8), .B(x0), .Y(men_men_n155_));
  BUFFER     u139(.A(men_men_n155_), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n41_), .B(x2), .Y(men_men_n157_));
  INV        u141(.A(x7), .Y(men_men_n158_));
  NA2        u142(.A(men_men_n158_), .B(men_men_n18_), .Y(men_men_n159_));
  NA2        u143(.A(men_men_n159_), .B(men_men_n157_), .Y(men_men_n160_));
  NO2        u144(.A(men_men_n25_), .B(x4), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n161_), .B(men_men_n127_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n162_), .B(men_men_n160_), .Y(men_men_n163_));
  AOI210     u147(.A0(men_men_n156_), .A1(men_men_n153_), .B0(men_men_n163_), .Y(men_men_n164_));
  OAI210     u148(.A0(men_men_n152_), .A1(men_men_n48_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u149(.A(x5), .B(x1), .Y(men_men_n166_));
  INV        u150(.A(men_men_n166_), .Y(men_men_n167_));
  AOI210     u151(.A0(men_men_n167_), .A1(men_men_n127_), .B0(men_men_n36_), .Y(men_men_n168_));
  NO2        u152(.A(men_men_n59_), .B(men_men_n92_), .Y(men_men_n169_));
  NAi21      u153(.An(x2), .B(x7), .Y(men_men_n170_));
  NO3        u154(.A(men_men_n170_), .B(men_men_n169_), .C(men_men_n46_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n171_), .B(men_men_n64_), .Y(men_men_n172_));
  NA2        u156(.A(men_men_n172_), .B(men_men_n168_), .Y(men_men_n173_));
  NO4        u157(.A(men_men_n173_), .B(men_men_n165_), .C(men_men_n151_), .D(men_men_n148_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n174_), .B(men_men_n147_), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n143_), .B(men_men_n139_), .Y(men_men_n176_));
  NA2        u160(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n177_));
  NA2        u161(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n178_));
  NA3        u162(.A(men_men_n178_), .B(men_men_n177_), .C(men_men_n24_), .Y(men_men_n179_));
  AN2        u163(.A(men_men_n179_), .B(men_men_n144_), .Y(men_men_n180_));
  NA2        u164(.A(x8), .B(x0), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n158_), .B(men_men_n25_), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n125_), .B(x4), .Y(men_men_n183_));
  NA2        u167(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  AOI210     u168(.A0(men_men_n181_), .A1(men_men_n133_), .B0(men_men_n184_), .Y(men_men_n185_));
  NA2        u169(.A(x2), .B(x0), .Y(men_men_n186_));
  NA2        u170(.A(x4), .B(x1), .Y(men_men_n187_));
  NAi21      u171(.An(men_men_n123_), .B(men_men_n187_), .Y(men_men_n188_));
  NOi31      u172(.An(men_men_n188_), .B(men_men_n161_), .C(men_men_n186_), .Y(men_men_n189_));
  NO4        u173(.A(men_men_n189_), .B(men_men_n185_), .C(men_men_n180_), .D(men_men_n176_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n190_), .B(men_men_n41_), .Y(men_men_n191_));
  NO2        u175(.A(men_men_n179_), .B(men_men_n74_), .Y(men_men_n192_));
  INV        u176(.A(men_men_n132_), .Y(men_men_n193_));
  NO2        u177(.A(men_men_n106_), .B(men_men_n17_), .Y(men_men_n194_));
  NA3        u178(.A(men_men_n188_), .B(men_men_n193_), .C(men_men_n40_), .Y(men_men_n195_));
  OAI210     u179(.A0(men_men_n178_), .A1(men_men_n139_), .B0(men_men_n195_), .Y(men_men_n196_));
  NO2        u180(.A(men_men_n196_), .B(men_men_n192_), .Y(men_men_n197_));
  NO2        u181(.A(men_men_n197_), .B(x3), .Y(men_men_n198_));
  NO3        u182(.A(men_men_n198_), .B(men_men_n191_), .C(men_men_n175_), .Y(men03));
  NO2        u183(.A(men_men_n46_), .B(x3), .Y(men_men_n200_));
  NO2        u184(.A(x6), .B(men_men_n25_), .Y(men_men_n201_));
  INV        u185(.A(men_men_n201_), .Y(men_men_n202_));
  NO2        u186(.A(men_men_n51_), .B(x1), .Y(men_men_n203_));
  OAI210     u187(.A0(men_men_n203_), .A1(men_men_n25_), .B0(men_men_n60_), .Y(men_men_n204_));
  OAI220     u188(.A0(men_men_n204_), .A1(men_men_n17_), .B0(men_men_n202_), .B1(men_men_n106_), .Y(men_men_n205_));
  NA2        u189(.A(men_men_n205_), .B(men_men_n200_), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n76_), .B(x6), .Y(men_men_n207_));
  NA2        u191(.A(x6), .B(men_men_n25_), .Y(men_men_n208_));
  NO2        u192(.A(men_men_n208_), .B(x4), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n18_), .B(x0), .Y(men_men_n210_));
  AO220      u194(.A0(men_men_n210_), .A1(men_men_n209_), .B0(men_men_n207_), .B1(men_men_n52_), .Y(men_men_n211_));
  NA2        u195(.A(men_men_n211_), .B(men_men_n59_), .Y(men_men_n212_));
  NA2        u196(.A(x3), .B(men_men_n17_), .Y(men_men_n213_));
  NO3        u197(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n214_));
  NO2        u198(.A(x5), .B(x1), .Y(men_men_n215_));
  AOI220     u199(.A0(men_men_n215_), .A1(men_men_n17_), .B0(men_men_n103_), .B1(x5), .Y(men_men_n216_));
  NO2        u200(.A(men_men_n213_), .B(men_men_n177_), .Y(men_men_n217_));
  INV        u201(.A(men_men_n217_), .Y(men_men_n218_));
  OAI210     u202(.A0(men_men_n216_), .A1(men_men_n61_), .B0(men_men_n218_), .Y(men_men_n219_));
  AOI220     u203(.A0(men_men_n219_), .A1(men_men_n46_), .B0(men_men_n214_), .B1(men_men_n132_), .Y(men_men_n220_));
  NA3        u204(.A(men_men_n220_), .B(men_men_n212_), .C(men_men_n206_), .Y(men_men_n221_));
  NO2        u205(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n222_));
  NA2        u206(.A(men_men_n222_), .B(men_men_n19_), .Y(men_men_n223_));
  NO2        u207(.A(x3), .B(men_men_n17_), .Y(men_men_n224_));
  NO2        u208(.A(men_men_n224_), .B(x6), .Y(men_men_n225_));
  NOi21      u209(.An(men_men_n82_), .B(men_men_n225_), .Y(men_men_n226_));
  NA2        u210(.A(men_men_n59_), .B(men_men_n92_), .Y(men_men_n227_));
  NA2        u211(.A(men_men_n224_), .B(x6), .Y(men_men_n228_));
  AOI210     u212(.A0(men_men_n228_), .A1(men_men_n226_), .B0(men_men_n158_), .Y(men_men_n229_));
  AO210      u213(.A0(men_men_n229_), .A1(men_men_n223_), .B0(men_men_n182_), .Y(men_men_n230_));
  NA2        u214(.A(men_men_n41_), .B(men_men_n51_), .Y(men_men_n231_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n25_), .B0(men_men_n178_), .Y(men_men_n232_));
  NO3        u216(.A(men_men_n187_), .B(men_men_n59_), .C(x6), .Y(men_men_n233_));
  AOI220     u217(.A0(men_men_n233_), .A1(men_men_n232_), .B0(men_men_n144_), .B1(men_men_n91_), .Y(men_men_n234_));
  NA2        u218(.A(x6), .B(men_men_n46_), .Y(men_men_n235_));
  OAI210     u219(.A0(men_men_n119_), .A1(men_men_n77_), .B0(x4), .Y(men_men_n236_));
  AOI210     u220(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n76_), .Y(men_men_n237_));
  NO2        u221(.A(men_men_n59_), .B(x6), .Y(men_men_n238_));
  NO2        u222(.A(men_men_n166_), .B(men_men_n41_), .Y(men_men_n239_));
  OAI210     u223(.A0(men_men_n239_), .A1(men_men_n217_), .B0(men_men_n238_), .Y(men_men_n240_));
  NA2        u224(.A(men_men_n201_), .B(men_men_n137_), .Y(men_men_n241_));
  NA3        u225(.A(men_men_n213_), .B(men_men_n132_), .C(x6), .Y(men_men_n242_));
  OAI210     u226(.A0(men_men_n92_), .A1(men_men_n36_), .B0(men_men_n64_), .Y(men_men_n243_));
  NA4        u227(.A(men_men_n243_), .B(men_men_n242_), .C(men_men_n241_), .D(men_men_n240_), .Y(men_men_n244_));
  OAI210     u228(.A0(men_men_n244_), .A1(men_men_n237_), .B0(x2), .Y(men_men_n245_));
  NA3        u229(.A(men_men_n245_), .B(men_men_n234_), .C(men_men_n230_), .Y(men_men_n246_));
  AOI210     u230(.A0(men_men_n221_), .A1(x8), .B0(men_men_n246_), .Y(men_men_n247_));
  NO2        u231(.A(men_men_n92_), .B(x3), .Y(men_men_n248_));
  NO3        u232(.A(men_men_n90_), .B(men_men_n77_), .C(men_men_n25_), .Y(men_men_n249_));
  AOI210     u233(.A0(men_men_n225_), .A1(men_men_n161_), .B0(men_men_n249_), .Y(men_men_n250_));
  NO2        u234(.A(men_men_n250_), .B(x2), .Y(men_men_n251_));
  NO2        u235(.A(x4), .B(men_men_n51_), .Y(men_men_n252_));
  AOI220     u236(.A0(men_men_n209_), .A1(men_men_n194_), .B0(men_men_n252_), .B1(men_men_n64_), .Y(men_men_n253_));
  NA2        u237(.A(men_men_n59_), .B(x6), .Y(men_men_n254_));
  NA2        u238(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n255_));
  NO2        u239(.A(men_men_n255_), .B(men_men_n25_), .Y(men_men_n256_));
  NA2        u240(.A(men_men_n256_), .B(men_men_n123_), .Y(men_men_n257_));
  NA2        u241(.A(men_men_n213_), .B(x6), .Y(men_men_n258_));
  NO2        u242(.A(men_men_n213_), .B(x6), .Y(men_men_n259_));
  NA2        u243(.A(men_men_n258_), .B(men_men_n149_), .Y(men_men_n260_));
  NA4        u244(.A(men_men_n260_), .B(men_men_n257_), .C(men_men_n253_), .D(men_men_n158_), .Y(men_men_n261_));
  NA2        u245(.A(men_men_n201_), .B(men_men_n224_), .Y(men_men_n262_));
  NAi21      u246(.An(x1), .B(x4), .Y(men_men_n263_));
  AOI210     u247(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n264_));
  OAI210     u248(.A0(men_men_n143_), .A1(x3), .B0(men_men_n264_), .Y(men_men_n265_));
  NA2        u249(.A(men_men_n265_), .B(men_men_n263_), .Y(men_men_n266_));
  NA2        u250(.A(men_men_n266_), .B(men_men_n262_), .Y(men_men_n267_));
  NA2        u251(.A(men_men_n59_), .B(x2), .Y(men_men_n268_));
  NO2        u252(.A(men_men_n268_), .B(men_men_n262_), .Y(men_men_n269_));
  NO3        u253(.A(x9), .B(x6), .C(x0), .Y(men_men_n270_));
  NA2        u254(.A(men_men_n106_), .B(men_men_n25_), .Y(men_men_n271_));
  NA2        u255(.A(x6), .B(x2), .Y(men_men_n272_));
  NO2        u256(.A(men_men_n272_), .B(men_men_n177_), .Y(men_men_n273_));
  AOI210     u257(.A0(men_men_n271_), .A1(men_men_n270_), .B0(men_men_n273_), .Y(men_men_n274_));
  OAI220     u258(.A0(men_men_n274_), .A1(men_men_n41_), .B0(men_men_n183_), .B1(men_men_n44_), .Y(men_men_n275_));
  OAI210     u259(.A0(men_men_n275_), .A1(men_men_n269_), .B0(men_men_n267_), .Y(men_men_n276_));
  NA2        u260(.A(x9), .B(men_men_n41_), .Y(men_men_n277_));
  NO2        u261(.A(men_men_n277_), .B(men_men_n208_), .Y(men_men_n278_));
  OR3        u262(.A(men_men_n278_), .B(men_men_n207_), .C(men_men_n153_), .Y(men_men_n279_));
  NA2        u263(.A(x4), .B(x0), .Y(men_men_n280_));
  NO3        u264(.A(men_men_n71_), .B(men_men_n280_), .C(x6), .Y(men_men_n281_));
  AOI210     u265(.A0(men_men_n279_), .A1(men_men_n40_), .B0(men_men_n281_), .Y(men_men_n282_));
  AOI210     u266(.A0(men_men_n282_), .A1(men_men_n276_), .B0(x8), .Y(men_men_n283_));
  NA2        u267(.A(men_men_n215_), .B(x6), .Y(men_men_n284_));
  INV        u268(.A(men_men_n181_), .Y(men_men_n285_));
  OAI210     u269(.A0(men_men_n285_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n286_));
  AOI210     u270(.A0(men_men_n286_), .A1(men_men_n284_), .B0(men_men_n231_), .Y(men_men_n287_));
  NO4        u271(.A(men_men_n287_), .B(men_men_n283_), .C(men_men_n261_), .D(men_men_n251_), .Y(men_men_n288_));
  NO2        u272(.A(men_men_n169_), .B(x1), .Y(men_men_n289_));
  NO3        u273(.A(men_men_n289_), .B(x3), .C(men_men_n36_), .Y(men_men_n290_));
  OAI210     u274(.A0(men_men_n290_), .A1(men_men_n259_), .B0(x2), .Y(men_men_n291_));
  OAI210     u275(.A0(men_men_n285_), .A1(x6), .B0(men_men_n42_), .Y(men_men_n292_));
  AOI210     u276(.A0(men_men_n292_), .A1(men_men_n291_), .B0(men_men_n193_), .Y(men_men_n293_));
  NOi21      u277(.An(men_men_n272_), .B(men_men_n17_), .Y(men_men_n294_));
  NA3        u278(.A(men_men_n294_), .B(men_men_n215_), .C(men_men_n38_), .Y(men_men_n295_));
  AOI210     u279(.A0(men_men_n36_), .A1(men_men_n51_), .B0(x0), .Y(men_men_n296_));
  NA3        u280(.A(men_men_n296_), .B(men_men_n167_), .C(men_men_n32_), .Y(men_men_n297_));
  NA2        u281(.A(x3), .B(x2), .Y(men_men_n298_));
  AOI220     u282(.A0(men_men_n298_), .A1(men_men_n231_), .B0(men_men_n297_), .B1(men_men_n295_), .Y(men_men_n299_));
  NAi21      u283(.An(x4), .B(x0), .Y(men_men_n300_));
  NO3        u284(.A(men_men_n300_), .B(men_men_n42_), .C(x2), .Y(men_men_n301_));
  OAI210     u285(.A0(x6), .A1(men_men_n18_), .B0(men_men_n301_), .Y(men_men_n302_));
  OAI220     u286(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n303_));
  NO2        u287(.A(x9), .B(x8), .Y(men_men_n304_));
  NA3        u288(.A(men_men_n304_), .B(men_men_n36_), .C(men_men_n51_), .Y(men_men_n305_));
  OAI210     u289(.A0(men_men_n296_), .A1(men_men_n294_), .B0(men_men_n305_), .Y(men_men_n306_));
  AOI220     u290(.A0(men_men_n306_), .A1(men_men_n80_), .B0(men_men_n303_), .B1(men_men_n31_), .Y(men_men_n307_));
  AOI210     u291(.A0(men_men_n307_), .A1(men_men_n302_), .B0(men_men_n25_), .Y(men_men_n308_));
  NA3        u292(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n309_));
  OAI210     u293(.A0(men_men_n296_), .A1(men_men_n294_), .B0(men_men_n309_), .Y(men_men_n310_));
  INV        u294(.A(men_men_n217_), .Y(men_men_n311_));
  NA2        u295(.A(men_men_n36_), .B(men_men_n41_), .Y(men_men_n312_));
  OR2        u296(.A(men_men_n312_), .B(men_men_n280_), .Y(men_men_n313_));
  OAI220     u297(.A0(men_men_n313_), .A1(men_men_n166_), .B0(men_men_n235_), .B1(men_men_n311_), .Y(men_men_n314_));
  AO210      u298(.A0(men_men_n310_), .A1(men_men_n153_), .B0(men_men_n314_), .Y(men_men_n315_));
  NO4        u299(.A(men_men_n315_), .B(men_men_n308_), .C(men_men_n299_), .D(men_men_n293_), .Y(men_men_n316_));
  OAI210     u300(.A0(men_men_n288_), .A1(men_men_n247_), .B0(men_men_n316_), .Y(men04));
  OAI210     u301(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n318_));
  NA3        u302(.A(men_men_n318_), .B(men_men_n270_), .C(men_men_n83_), .Y(men_men_n319_));
  NO2        u303(.A(x2), .B(x1), .Y(men_men_n320_));
  OAI210     u304(.A0(men_men_n255_), .A1(men_men_n320_), .B0(men_men_n36_), .Y(men_men_n321_));
  NO2        u305(.A(men_men_n320_), .B(men_men_n300_), .Y(men_men_n322_));
  AOI210     u306(.A0(men_men_n59_), .A1(x4), .B0(men_men_n112_), .Y(men_men_n323_));
  OAI210     u307(.A0(men_men_n323_), .A1(men_men_n322_), .B0(men_men_n248_), .Y(men_men_n324_));
  NO2        u308(.A(men_men_n298_), .B(men_men_n210_), .Y(men_men_n325_));
  NA2        u309(.A(x9), .B(x0), .Y(men_men_n326_));
  AOI210     u310(.A0(men_men_n90_), .A1(men_men_n74_), .B0(men_men_n326_), .Y(men_men_n327_));
  OAI210     u311(.A0(men_men_n327_), .A1(men_men_n325_), .B0(men_men_n92_), .Y(men_men_n328_));
  NA3        u312(.A(men_men_n328_), .B(x6), .C(men_men_n324_), .Y(men_men_n329_));
  NA2        u313(.A(men_men_n329_), .B(men_men_n321_), .Y(men_men_n330_));
  NO2        u314(.A(x2), .B(men_men_n113_), .Y(men_men_n331_));
  NO3        u315(.A(men_men_n254_), .B(men_men_n120_), .C(men_men_n18_), .Y(men_men_n332_));
  NO2        u316(.A(men_men_n332_), .B(men_men_n331_), .Y(men_men_n333_));
  OAI210     u317(.A0(men_men_n118_), .A1(men_men_n106_), .B0(men_men_n181_), .Y(men_men_n334_));
  NA3        u318(.A(men_men_n334_), .B(x6), .C(x3), .Y(men_men_n335_));
  AOI210     u319(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n336_));
  NO2        u320(.A(men_men_n336_), .B(men_men_n312_), .Y(men_men_n337_));
  INV        u321(.A(men_men_n337_), .Y(men_men_n338_));
  NA2        u322(.A(x2), .B(men_men_n17_), .Y(men_men_n339_));
  OAI210     u323(.A0(men_men_n106_), .A1(men_men_n17_), .B0(men_men_n339_), .Y(men_men_n340_));
  NA2        u324(.A(men_men_n340_), .B(men_men_n77_), .Y(men_men_n341_));
  NA4        u325(.A(men_men_n341_), .B(men_men_n338_), .C(men_men_n335_), .D(men_men_n333_), .Y(men_men_n342_));
  OAI210     u326(.A0(men_men_n111_), .A1(x3), .B0(men_men_n301_), .Y(men_men_n343_));
  NA3        u327(.A(men_men_n227_), .B(men_men_n214_), .C(men_men_n82_), .Y(men_men_n344_));
  NA3        u328(.A(men_men_n344_), .B(men_men_n343_), .C(men_men_n158_), .Y(men_men_n345_));
  AOI210     u329(.A0(men_men_n342_), .A1(x4), .B0(men_men_n345_), .Y(men_men_n346_));
  NOi21      u330(.An(x4), .B(x0), .Y(men_men_n347_));
  XO2        u331(.A(x4), .B(x0), .Y(men_men_n348_));
  OAI210     u332(.A0(men_men_n348_), .A1(men_men_n117_), .B0(men_men_n263_), .Y(men_men_n349_));
  AOI220     u333(.A0(men_men_n349_), .A1(x8), .B0(men_men_n347_), .B1(men_men_n93_), .Y(men_men_n350_));
  NO2        u334(.A(men_men_n350_), .B(x3), .Y(men_men_n351_));
  INV        u335(.A(men_men_n93_), .Y(men_men_n352_));
  NO2        u336(.A(men_men_n92_), .B(x4), .Y(men_men_n353_));
  AOI220     u337(.A0(men_men_n353_), .A1(men_men_n42_), .B0(men_men_n127_), .B1(men_men_n352_), .Y(men_men_n354_));
  NO3        u338(.A(men_men_n348_), .B(men_men_n169_), .C(x2), .Y(men_men_n355_));
  INV        u339(.A(men_men_n355_), .Y(men_men_n356_));
  NA4        u340(.A(men_men_n356_), .B(men_men_n354_), .C(men_men_n223_), .D(x6), .Y(men_men_n357_));
  OAI220     u341(.A0(men_men_n300_), .A1(men_men_n90_), .B0(men_men_n186_), .B1(men_men_n92_), .Y(men_men_n358_));
  NO2        u342(.A(men_men_n41_), .B(x0), .Y(men_men_n359_));
  OR2        u343(.A(men_men_n353_), .B(men_men_n359_), .Y(men_men_n360_));
  NO2        u344(.A(men_men_n155_), .B(men_men_n106_), .Y(men_men_n361_));
  AOI220     u345(.A0(men_men_n361_), .A1(men_men_n360_), .B0(men_men_n358_), .B1(men_men_n58_), .Y(men_men_n362_));
  NO2        u346(.A(men_men_n155_), .B(men_men_n79_), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n35_), .B(x2), .Y(men_men_n364_));
  NOi21      u348(.An(men_men_n123_), .B(men_men_n27_), .Y(men_men_n365_));
  AOI210     u349(.A0(men_men_n364_), .A1(men_men_n363_), .B0(men_men_n365_), .Y(men_men_n366_));
  OAI210     u350(.A0(men_men_n362_), .A1(men_men_n59_), .B0(men_men_n366_), .Y(men_men_n367_));
  OAI220     u351(.A0(men_men_n367_), .A1(x6), .B0(men_men_n357_), .B1(men_men_n351_), .Y(men_men_n368_));
  INV        u352(.A(men_men_n313_), .Y(men_men_n369_));
  AOI210     u353(.A0(men_men_n369_), .A1(men_men_n18_), .B0(men_men_n158_), .Y(men_men_n370_));
  AO220      u354(.A0(men_men_n370_), .A1(men_men_n368_), .B0(men_men_n346_), .B1(men_men_n330_), .Y(men_men_n371_));
  NA2        u355(.A(men_men_n364_), .B(x6), .Y(men_men_n372_));
  AOI210     u356(.A0(x6), .A1(x1), .B0(men_men_n157_), .Y(men_men_n373_));
  NA2        u357(.A(men_men_n353_), .B(x0), .Y(men_men_n374_));
  NA2        u358(.A(men_men_n82_), .B(x6), .Y(men_men_n375_));
  OAI210     u359(.A0(men_men_n374_), .A1(men_men_n373_), .B0(men_men_n375_), .Y(men_men_n376_));
  NA2        u360(.A(men_men_n376_), .B(men_men_n372_), .Y(men_men_n377_));
  NA3        u361(.A(men_men_n377_), .B(men_men_n371_), .C(men_men_n319_), .Y(men_men_n378_));
  AOI210     u362(.A0(men_men_n203_), .A1(x8), .B0(men_men_n111_), .Y(men_men_n379_));
  NA2        u363(.A(men_men_n379_), .B(men_men_n339_), .Y(men_men_n380_));
  NA3        u364(.A(men_men_n380_), .B(men_men_n200_), .C(men_men_n158_), .Y(men_men_n381_));
  OAI210     u365(.A0(men_men_n28_), .A1(x1), .B0(men_men_n231_), .Y(men_men_n382_));
  AO220      u366(.A0(men_men_n382_), .A1(men_men_n154_), .B0(men_men_n110_), .B1(x4), .Y(men_men_n383_));
  NA3        u367(.A(x7), .B(x3), .C(x0), .Y(men_men_n384_));
  NA2        u368(.A(men_men_n222_), .B(x0), .Y(men_men_n385_));
  OAI220     u369(.A0(men_men_n385_), .A1(x2), .B0(men_men_n384_), .B1(men_men_n352_), .Y(men_men_n386_));
  AOI210     u370(.A0(men_men_n383_), .A1(men_men_n119_), .B0(men_men_n386_), .Y(men_men_n387_));
  AOI210     u371(.A0(men_men_n387_), .A1(men_men_n381_), .B0(men_men_n25_), .Y(men_men_n388_));
  NA3        u372(.A(men_men_n121_), .B(men_men_n222_), .C(x0), .Y(men_men_n389_));
  NAi31      u373(.An(men_men_n48_), .B(men_men_n289_), .C(men_men_n182_), .Y(men_men_n390_));
  NA2        u374(.A(men_men_n390_), .B(men_men_n389_), .Y(men_men_n391_));
  OAI210     u375(.A0(men_men_n391_), .A1(men_men_n388_), .B0(x6), .Y(men_men_n392_));
  AOI210     u376(.A0(men_men_n38_), .A1(men_men_n32_), .B0(x0), .Y(men_men_n393_));
  NA2        u377(.A(men_men_n200_), .B(men_men_n158_), .Y(men_men_n394_));
  AOI210     u378(.A0(men_men_n129_), .A1(men_men_n252_), .B0(x1), .Y(men_men_n395_));
  OAI210     u379(.A0(men_men_n394_), .A1(x8), .B0(men_men_n395_), .Y(men_men_n396_));
  INV        u380(.A(men_men_n170_), .Y(men_men_n397_));
  NA3        u381(.A(men_men_n397_), .B(men_men_n152_), .C(x9), .Y(men_men_n398_));
  NO4        u382(.A(men_men_n128_), .B(men_men_n300_), .C(x9), .D(x2), .Y(men_men_n399_));
  NOi21      u383(.An(men_men_n126_), .B(men_men_n186_), .Y(men_men_n400_));
  NO3        u384(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n18_), .Y(men_men_n401_));
  NO3        u385(.A(x9), .B(men_men_n158_), .C(x0), .Y(men_men_n402_));
  AOI220     u386(.A0(men_men_n402_), .A1(men_men_n248_), .B0(men_men_n363_), .B1(men_men_n158_), .Y(men_men_n403_));
  NA4        u387(.A(men_men_n403_), .B(men_men_n401_), .C(men_men_n398_), .D(men_men_n48_), .Y(men_men_n404_));
  OAI210     u388(.A0(men_men_n396_), .A1(men_men_n393_), .B0(men_men_n404_), .Y(men_men_n405_));
  INV        u389(.A(men_men_n136_), .Y(men_men_n406_));
  NO3        u390(.A(men_men_n406_), .B(men_men_n126_), .C(men_men_n41_), .Y(men_men_n407_));
  NOi31      u391(.An(x1), .B(x8), .C(x7), .Y(men_men_n408_));
  AOI210     u392(.A0(men_men_n127_), .A1(x3), .B0(men_men_n408_), .Y(men_men_n409_));
  AOI210     u393(.A0(men_men_n263_), .A1(men_men_n57_), .B0(men_men_n125_), .Y(men_men_n410_));
  OAI210     u394(.A0(men_men_n410_), .A1(x3), .B0(men_men_n409_), .Y(men_men_n411_));
  NO3        u395(.A(men_men_n411_), .B(men_men_n407_), .C(x2), .Y(men_men_n412_));
  OAI220     u396(.A0(men_men_n348_), .A1(men_men_n304_), .B0(men_men_n300_), .B1(men_men_n41_), .Y(men_men_n413_));
  AOI210     u397(.A0(x9), .A1(men_men_n46_), .B0(men_men_n384_), .Y(men_men_n414_));
  AOI220     u398(.A0(men_men_n414_), .A1(men_men_n92_), .B0(men_men_n413_), .B1(men_men_n158_), .Y(men_men_n415_));
  NO2        u399(.A(men_men_n415_), .B(men_men_n51_), .Y(men_men_n416_));
  NO2        u400(.A(men_men_n416_), .B(men_men_n412_), .Y(men_men_n417_));
  AOI210     u401(.A0(men_men_n417_), .A1(men_men_n405_), .B0(men_men_n25_), .Y(men_men_n418_));
  NA4        u402(.A(men_men_n31_), .B(men_men_n92_), .C(x2), .D(men_men_n17_), .Y(men_men_n419_));
  NO3        u403(.A(men_men_n65_), .B(men_men_n18_), .C(x0), .Y(men_men_n420_));
  NA2        u404(.A(men_men_n420_), .B(men_men_n264_), .Y(men_men_n421_));
  NO2        u405(.A(men_men_n421_), .B(men_men_n103_), .Y(men_men_n422_));
  NO3        u406(.A(men_men_n268_), .B(men_men_n181_), .C(men_men_n38_), .Y(men_men_n423_));
  OAI210     u407(.A0(men_men_n423_), .A1(men_men_n422_), .B0(x7), .Y(men_men_n424_));
  NA2        u408(.A(men_men_n227_), .B(x7), .Y(men_men_n425_));
  NA3        u409(.A(men_men_n425_), .B(men_men_n157_), .C(men_men_n137_), .Y(men_men_n426_));
  NA3        u410(.A(men_men_n426_), .B(men_men_n424_), .C(men_men_n419_), .Y(men_men_n427_));
  OAI210     u411(.A0(men_men_n427_), .A1(men_men_n418_), .B0(men_men_n36_), .Y(men_men_n428_));
  NO2        u412(.A(men_men_n402_), .B(men_men_n210_), .Y(men_men_n429_));
  NO4        u413(.A(men_men_n429_), .B(men_men_n76_), .C(x4), .D(men_men_n51_), .Y(men_men_n430_));
  NA2        u414(.A(men_men_n359_), .B(men_men_n182_), .Y(men_men_n431_));
  OAI220     u415(.A0(men_men_n277_), .A1(men_men_n66_), .B0(men_men_n166_), .B1(men_men_n41_), .Y(men_men_n432_));
  NA2        u416(.A(x3), .B(men_men_n51_), .Y(men_men_n433_));
  AOI210     u417(.A0(men_men_n170_), .A1(men_men_n27_), .B0(men_men_n71_), .Y(men_men_n434_));
  OAI210     u418(.A0(men_men_n154_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n435_));
  NO3        u419(.A(men_men_n408_), .B(x3), .C(men_men_n51_), .Y(men_men_n436_));
  AOI210     u420(.A0(men_men_n436_), .A1(men_men_n435_), .B0(men_men_n434_), .Y(men_men_n437_));
  OAI210     u421(.A0(men_men_n159_), .A1(men_men_n433_), .B0(men_men_n437_), .Y(men_men_n438_));
  AOI220     u422(.A0(men_men_n438_), .A1(x0), .B0(men_men_n432_), .B1(men_men_n138_), .Y(men_men_n439_));
  AOI210     u423(.A0(men_men_n439_), .A1(men_men_n431_), .B0(men_men_n235_), .Y(men_men_n440_));
  INV        u424(.A(x5), .Y(men_men_n441_));
  NO4        u425(.A(men_men_n106_), .B(men_men_n441_), .C(men_men_n57_), .D(men_men_n32_), .Y(men_men_n442_));
  NO3        u426(.A(men_men_n442_), .B(men_men_n440_), .C(men_men_n430_), .Y(men_men_n443_));
  NA3        u427(.A(men_men_n443_), .B(men_men_n428_), .C(men_men_n392_), .Y(men_men_n444_));
  AOI210     u428(.A0(men_men_n378_), .A1(men_men_n25_), .B0(men_men_n444_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule