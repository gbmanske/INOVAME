// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n132_, new_new_n133_, new_new_n134_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n996_, new_new_n997_, new_new_n998_, new_new_n999_,
    new_new_n1000_, new_new_n1001_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA3        g031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  OAI210     g034(.A0(new_new_n56_), .A1(new_new_n55_), .B0(new_new_n54_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_12_), .Y(new_new_n58_));
  NAi21      g036(.An(i_2_), .B(i_7_), .Y(new_new_n59_));
  INV        g037(.A(i_1_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_6_), .Y(new_new_n61_));
  NA3        g039(.A(new_new_n61_), .B(new_new_n59_), .C(new_new_n31_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_10_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NAi31      g042(.An(new_new_n64_), .B(new_new_n62_), .C(new_new_n58_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n50_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NA2        g055(.A(i_2_), .B(i_8_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_9_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_7_), .Y(new_new_n80_));
  NO3        g058(.A(new_new_n80_), .B(new_new_n79_), .C(new_new_n60_), .Y(new_new_n81_));
  INV        g059(.A(i_6_), .Y(new_new_n82_));
  NO2        g060(.A(i_2_), .B(i_7_), .Y(new_new_n83_));
  INV        g061(.A(new_new_n83_), .Y(new_new_n84_));
  NA2        g062(.A(new_new_n81_), .B(new_new_n84_), .Y(new_new_n85_));
  NAi21      g063(.An(i_6_), .B(i_10_), .Y(new_new_n86_));
  NA2        g064(.A(i_6_), .B(i_9_), .Y(new_new_n87_));
  AOI210     g065(.A0(new_new_n87_), .A1(new_new_n86_), .B0(new_new_n60_), .Y(new_new_n88_));
  NA2        g066(.A(i_2_), .B(i_6_), .Y(new_new_n89_));
  NO3        g067(.A(new_new_n89_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n90_));
  NO2        g068(.A(new_new_n90_), .B(new_new_n88_), .Y(new_new_n91_));
  AOI210     g069(.A0(new_new_n91_), .A1(new_new_n85_), .B0(new_new_n77_), .Y(new_new_n92_));
  AN3        g070(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n93_));
  NAi21      g071(.An(i_6_), .B(i_11_), .Y(new_new_n94_));
  NO2        g072(.A(i_5_), .B(i_8_), .Y(new_new_n95_));
  NOi21      g073(.An(new_new_n95_), .B(new_new_n94_), .Y(new_new_n96_));
  AOI220     g074(.A0(new_new_n96_), .A1(new_new_n59_), .B0(new_new_n93_), .B1(new_new_n32_), .Y(new_new_n97_));
  INV        g075(.A(i_7_), .Y(new_new_n98_));
  NA2        g076(.A(new_new_n46_), .B(new_new_n98_), .Y(new_new_n99_));
  NO2        g077(.A(i_0_), .B(i_5_), .Y(new_new_n100_));
  NO2        g078(.A(new_new_n100_), .B(new_new_n82_), .Y(new_new_n101_));
  NA2        g079(.A(i_12_), .B(i_3_), .Y(new_new_n102_));
  INV        g080(.A(new_new_n102_), .Y(new_new_n103_));
  NA3        g081(.A(new_new_n103_), .B(new_new_n101_), .C(new_new_n99_), .Y(new_new_n104_));
  NAi21      g082(.An(i_7_), .B(i_11_), .Y(new_new_n105_));
  AN2        g083(.A(i_2_), .B(i_10_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(i_7_), .Y(new_new_n107_));
  OR2        g085(.A(new_new_n77_), .B(new_new_n55_), .Y(new_new_n108_));
  NO2        g086(.A(i_8_), .B(new_new_n98_), .Y(new_new_n109_));
  NO3        g087(.A(new_new_n109_), .B(new_new_n108_), .C(new_new_n107_), .Y(new_new_n110_));
  NA2        g088(.A(i_12_), .B(i_7_), .Y(new_new_n111_));
  NA2        g089(.A(i_11_), .B(i_12_), .Y(new_new_n112_));
  INV        g090(.A(new_new_n112_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n113_), .B(new_new_n110_), .Y(new_new_n114_));
  NA3        g092(.A(new_new_n114_), .B(new_new_n104_), .C(new_new_n97_), .Y(new_new_n115_));
  NOi21      g093(.An(i_1_), .B(i_5_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(i_11_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n98_), .B(new_new_n37_), .Y(new_new_n118_));
  NA2        g096(.A(i_7_), .B(new_new_n25_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(new_new_n118_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(new_new_n46_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n87_), .B(new_new_n86_), .Y(new_new_n122_));
  NAi21      g100(.An(i_3_), .B(i_8_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n59_), .Y(new_new_n124_));
  NOi31      g102(.An(new_new_n124_), .B(new_new_n122_), .C(new_new_n121_), .Y(new_new_n125_));
  NO2        g103(.A(i_1_), .B(new_new_n82_), .Y(new_new_n126_));
  NO2        g104(.A(i_6_), .B(i_5_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(i_3_), .Y(new_new_n128_));
  OAI220     g106(.A0(new_new_n128_), .A1(new_new_n105_), .B0(new_new_n125_), .B1(new_new_n117_), .Y(new_new_n129_));
  NO3        g107(.A(new_new_n129_), .B(new_new_n115_), .C(new_new_n92_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n130_), .B(new_new_n76_), .Y(mai2));
  NO2        g109(.A(new_new_n60_), .B(new_new_n37_), .Y(new_new_n132_));
  NA2        g110(.A(i_6_), .B(new_new_n25_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(new_new_n132_), .Y(new_new_n134_));
  NA4        g112(.A(new_new_n134_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(mai0));
  AN2        g113(.A(i_8_), .B(i_7_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(i_6_), .Y(new_new_n137_));
  NO2        g115(.A(i_12_), .B(i_13_), .Y(new_new_n138_));
  NAi21      g116(.An(i_5_), .B(i_11_), .Y(new_new_n139_));
  NOi21      g117(.An(new_new_n138_), .B(new_new_n139_), .Y(new_new_n140_));
  NO2        g118(.A(i_0_), .B(i_1_), .Y(new_new_n141_));
  NA2        g119(.A(i_2_), .B(i_3_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n142_), .B(i_4_), .Y(new_new_n143_));
  NA3        g121(.A(new_new_n143_), .B(new_new_n141_), .C(new_new_n140_), .Y(new_new_n144_));
  AN2        g122(.A(new_new_n138_), .B(new_new_n79_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(new_new_n27_), .Y(new_new_n146_));
  NA2        g124(.A(i_1_), .B(i_5_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n70_), .B(new_new_n46_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n36_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  OR2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NO3        g129(.A(new_new_n151_), .B(new_new_n77_), .C(i_13_), .Y(new_new_n152_));
  NAi32      g130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n153_));
  NAi21      g131(.An(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  NOi21      g132(.An(i_4_), .B(i_10_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n40_), .Y(new_new_n156_));
  NO2        g134(.A(i_3_), .B(i_5_), .Y(new_new_n157_));
  NO3        g135(.A(new_new_n70_), .B(i_2_), .C(i_1_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n157_), .Y(new_new_n159_));
  OAI210     g137(.A0(new_new_n159_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n160_), .B(new_new_n150_), .Y(new_new_n161_));
  AOI210     g139(.A0(new_new_n161_), .A1(new_new_n144_), .B0(new_new_n137_), .Y(new_new_n162_));
  NA2        g140(.A(i_3_), .B(new_new_n48_), .Y(new_new_n163_));
  NOi21      g141(.An(i_4_), .B(i_9_), .Y(new_new_n164_));
  NOi21      g142(.An(i_11_), .B(i_13_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OR2        g144(.A(new_new_n166_), .B(new_new_n163_), .Y(new_new_n167_));
  NO2        g145(.A(i_4_), .B(i_5_), .Y(new_new_n168_));
  NAi21      g146(.An(i_12_), .B(i_11_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n169_), .B(i_13_), .Y(new_new_n170_));
  NA3        g148(.A(new_new_n170_), .B(new_new_n168_), .C(new_new_n79_), .Y(new_new_n171_));
  AOI210     g149(.A0(new_new_n171_), .A1(new_new_n167_), .B0(new_new_n1001_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n70_), .B(new_new_n60_), .Y(new_new_n173_));
  NA2        g151(.A(new_new_n173_), .B(new_new_n46_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n36_), .B(i_5_), .Y(new_new_n175_));
  NAi31      g153(.An(new_new_n175_), .B(new_new_n145_), .C(i_11_), .Y(new_new_n176_));
  NA2        g154(.A(i_3_), .B(i_5_), .Y(new_new_n177_));
  AOI210     g155(.A0(new_new_n166_), .A1(new_new_n176_), .B0(new_new_n174_), .Y(new_new_n178_));
  NO2        g156(.A(new_new_n70_), .B(i_5_), .Y(new_new_n179_));
  NO2        g157(.A(i_13_), .B(i_10_), .Y(new_new_n180_));
  NA3        g158(.A(new_new_n180_), .B(new_new_n179_), .C(new_new_n44_), .Y(new_new_n181_));
  NO2        g159(.A(i_2_), .B(i_1_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n182_), .B(i_3_), .Y(new_new_n183_));
  NAi21      g161(.An(i_4_), .B(i_12_), .Y(new_new_n184_));
  NO4        g162(.A(new_new_n184_), .B(new_new_n183_), .C(new_new_n181_), .D(new_new_n25_), .Y(new_new_n185_));
  NO3        g163(.A(new_new_n185_), .B(new_new_n178_), .C(new_new_n172_), .Y(new_new_n186_));
  INV        g164(.A(i_8_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n187_), .B(i_7_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n188_), .B(i_6_), .Y(new_new_n189_));
  NO3        g167(.A(i_3_), .B(new_new_n82_), .C(new_new_n48_), .Y(new_new_n190_));
  NA2        g168(.A(new_new_n190_), .B(new_new_n109_), .Y(new_new_n191_));
  NO3        g169(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n192_));
  NA3        g170(.A(new_new_n192_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n193_));
  NO3        g171(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n194_));
  OAI210     g172(.A0(new_new_n93_), .A1(i_12_), .B0(new_new_n194_), .Y(new_new_n195_));
  AOI210     g173(.A0(new_new_n195_), .A1(new_new_n193_), .B0(new_new_n191_), .Y(new_new_n196_));
  NO2        g174(.A(i_3_), .B(i_8_), .Y(new_new_n197_));
  NO3        g175(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n198_));
  NO2        g176(.A(i_13_), .B(i_9_), .Y(new_new_n199_));
  NA3        g177(.A(new_new_n199_), .B(i_6_), .C(new_new_n187_), .Y(new_new_n200_));
  NAi21      g178(.An(i_12_), .B(i_3_), .Y(new_new_n201_));
  NO2        g179(.A(new_new_n44_), .B(i_5_), .Y(new_new_n202_));
  NO3        g180(.A(i_0_), .B(i_2_), .C(new_new_n60_), .Y(new_new_n203_));
  NA3        g181(.A(new_new_n203_), .B(new_new_n202_), .C(i_10_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n204_), .B(new_new_n200_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n205_), .B(new_new_n196_), .Y(new_new_n206_));
  OAI220     g184(.A0(new_new_n206_), .A1(i_4_), .B0(new_new_n189_), .B1(new_new_n186_), .Y(new_new_n207_));
  NAi21      g185(.An(i_12_), .B(i_7_), .Y(new_new_n208_));
  NA3        g186(.A(i_13_), .B(new_new_n187_), .C(i_10_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n209_), .B(new_new_n208_), .Y(new_new_n210_));
  NA2        g188(.A(i_0_), .B(i_5_), .Y(new_new_n211_));
  NA2        g189(.A(new_new_n211_), .B(new_new_n101_), .Y(new_new_n212_));
  OAI220     g190(.A0(new_new_n212_), .A1(new_new_n183_), .B0(new_new_n174_), .B1(new_new_n128_), .Y(new_new_n213_));
  NAi31      g191(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n36_), .B(i_13_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n70_), .B(new_new_n26_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n46_), .B(new_new_n60_), .Y(new_new_n217_));
  NA3        g195(.A(new_new_n217_), .B(new_new_n216_), .C(new_new_n215_), .Y(new_new_n218_));
  INV        g196(.A(i_13_), .Y(new_new_n219_));
  NO2        g197(.A(i_12_), .B(new_new_n219_), .Y(new_new_n220_));
  NA3        g198(.A(new_new_n220_), .B(new_new_n192_), .C(new_new_n190_), .Y(new_new_n221_));
  OAI210     g199(.A0(new_new_n218_), .A1(new_new_n214_), .B0(new_new_n221_), .Y(new_new_n222_));
  AOI220     g200(.A0(new_new_n222_), .A1(new_new_n136_), .B0(new_new_n213_), .B1(new_new_n210_), .Y(new_new_n223_));
  NO2        g201(.A(i_12_), .B(new_new_n37_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n177_), .B(i_4_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n226_));
  OR2        g204(.A(i_8_), .B(i_7_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n82_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n51_), .B(i_1_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n230_));
  INV        g208(.A(i_12_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n44_), .B(new_new_n231_), .Y(new_new_n232_));
  NO3        g210(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n233_));
  NA2        g211(.A(i_2_), .B(i_1_), .Y(new_new_n234_));
  NO2        g212(.A(new_new_n230_), .B(new_new_n226_), .Y(new_new_n235_));
  NO3        g213(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n236_));
  NAi21      g214(.An(i_4_), .B(i_3_), .Y(new_new_n237_));
  NO2        g215(.A(i_0_), .B(i_6_), .Y(new_new_n238_));
  NOi41      g216(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n239_));
  NA2        g217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  NO2        g218(.A(new_new_n234_), .B(new_new_n177_), .Y(new_new_n241_));
  NAi21      g219(.An(new_new_n240_), .B(new_new_n241_), .Y(new_new_n242_));
  INV        g220(.A(new_new_n242_), .Y(new_new_n243_));
  AOI210     g221(.A0(new_new_n243_), .A1(new_new_n40_), .B0(new_new_n235_), .Y(new_new_n244_));
  NO2        g222(.A(i_11_), .B(new_new_n219_), .Y(new_new_n245_));
  NOi21      g223(.An(i_1_), .B(i_6_), .Y(new_new_n246_));
  NAi21      g224(.An(i_3_), .B(i_7_), .Y(new_new_n247_));
  NA2        g225(.A(new_new_n231_), .B(i_9_), .Y(new_new_n248_));
  OR4        g226(.A(new_new_n248_), .B(new_new_n247_), .C(new_new_n246_), .D(new_new_n179_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n250_));
  NO2        g228(.A(i_12_), .B(i_3_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n70_), .B(i_5_), .Y(new_new_n252_));
  NA2        g230(.A(i_3_), .B(i_9_), .Y(new_new_n253_));
  NAi21      g231(.An(i_7_), .B(i_10_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n254_), .B(new_new_n253_), .Y(new_new_n255_));
  NA3        g233(.A(new_new_n255_), .B(new_new_n252_), .C(new_new_n61_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n256_), .B(new_new_n249_), .Y(new_new_n257_));
  NA3        g235(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n258_));
  INV        g236(.A(new_new_n137_), .Y(new_new_n259_));
  NA2        g237(.A(new_new_n231_), .B(i_13_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n260_), .B(new_new_n72_), .Y(new_new_n261_));
  AOI220     g239(.A0(new_new_n261_), .A1(new_new_n259_), .B0(new_new_n257_), .B1(new_new_n245_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n227_), .B(new_new_n37_), .Y(new_new_n263_));
  NA2        g241(.A(i_12_), .B(i_6_), .Y(new_new_n264_));
  OR2        g242(.A(i_13_), .B(i_9_), .Y(new_new_n265_));
  NO3        g243(.A(new_new_n265_), .B(new_new_n264_), .C(new_new_n48_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n237_), .B(i_2_), .Y(new_new_n267_));
  NA2        g245(.A(new_new_n245_), .B(i_9_), .Y(new_new_n268_));
  NA2        g246(.A(new_new_n148_), .B(new_new_n60_), .Y(new_new_n269_));
  NO3        g247(.A(i_11_), .B(new_new_n219_), .C(new_new_n25_), .Y(new_new_n270_));
  NO2        g248(.A(new_new_n247_), .B(i_8_), .Y(new_new_n271_));
  NO2        g249(.A(i_6_), .B(new_new_n48_), .Y(new_new_n272_));
  NA3        g250(.A(new_new_n272_), .B(new_new_n271_), .C(new_new_n270_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n26_), .B(new_new_n82_), .Y(new_new_n274_));
  NA3        g252(.A(new_new_n274_), .B(new_new_n263_), .C(new_new_n220_), .Y(new_new_n275_));
  AOI210     g253(.A0(new_new_n275_), .A1(new_new_n273_), .B0(new_new_n269_), .Y(new_new_n276_));
  INV        g254(.A(new_new_n276_), .Y(new_new_n277_));
  NA4        g255(.A(new_new_n277_), .B(new_new_n262_), .C(new_new_n244_), .D(new_new_n223_), .Y(new_new_n278_));
  NO3        g256(.A(i_12_), .B(new_new_n219_), .C(new_new_n37_), .Y(new_new_n279_));
  INV        g257(.A(new_new_n279_), .Y(new_new_n280_));
  NA2        g258(.A(i_8_), .B(new_new_n98_), .Y(new_new_n281_));
  NOi21      g259(.An(new_new_n157_), .B(new_new_n82_), .Y(new_new_n282_));
  NO3        g260(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n283_));
  AOI220     g261(.A0(new_new_n283_), .A1(new_new_n190_), .B0(new_new_n282_), .B1(new_new_n229_), .Y(new_new_n284_));
  NO2        g262(.A(new_new_n284_), .B(new_new_n281_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n234_), .B(i_0_), .Y(new_new_n286_));
  AOI220     g264(.A0(new_new_n286_), .A1(new_new_n188_), .B0(i_1_), .B1(new_new_n136_), .Y(new_new_n287_));
  NA2        g265(.A(new_new_n272_), .B(new_new_n26_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n288_), .B(new_new_n287_), .Y(new_new_n289_));
  NA2        g267(.A(i_0_), .B(i_1_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n290_), .B(i_2_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n56_), .B(i_6_), .Y(new_new_n292_));
  NA3        g270(.A(new_new_n292_), .B(new_new_n291_), .C(new_new_n157_), .Y(new_new_n293_));
  OAI210     g271(.A0(new_new_n159_), .A1(new_new_n137_), .B0(new_new_n293_), .Y(new_new_n294_));
  NO3        g272(.A(new_new_n294_), .B(new_new_n289_), .C(new_new_n285_), .Y(new_new_n295_));
  NO2        g273(.A(i_3_), .B(i_10_), .Y(new_new_n296_));
  NA3        g274(.A(new_new_n296_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n297_));
  NO2        g275(.A(i_2_), .B(new_new_n98_), .Y(new_new_n298_));
  NA2        g276(.A(i_1_), .B(new_new_n36_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n299_), .B(i_8_), .Y(new_new_n300_));
  NA2        g278(.A(new_new_n300_), .B(new_new_n298_), .Y(new_new_n301_));
  AN2        g279(.A(i_3_), .B(i_10_), .Y(new_new_n302_));
  NA4        g280(.A(new_new_n302_), .B(new_new_n192_), .C(new_new_n170_), .D(new_new_n168_), .Y(new_new_n303_));
  NO2        g281(.A(i_5_), .B(new_new_n37_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n305_));
  OR2        g283(.A(new_new_n301_), .B(new_new_n297_), .Y(new_new_n306_));
  OAI220     g284(.A0(new_new_n306_), .A1(i_6_), .B0(new_new_n295_), .B1(new_new_n280_), .Y(new_new_n307_));
  NO4        g285(.A(new_new_n307_), .B(new_new_n278_), .C(new_new_n207_), .D(new_new_n162_), .Y(new_new_n308_));
  NO3        g286(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n56_), .B(new_new_n82_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n286_), .B(new_new_n310_), .Y(new_new_n311_));
  NO3        g289(.A(i_6_), .B(new_new_n187_), .C(i_7_), .Y(new_new_n312_));
  NA2        g290(.A(new_new_n312_), .B(new_new_n192_), .Y(new_new_n313_));
  AOI210     g291(.A0(new_new_n313_), .A1(new_new_n311_), .B0(new_new_n163_), .Y(new_new_n314_));
  NO2        g292(.A(i_2_), .B(i_3_), .Y(new_new_n315_));
  OR2        g293(.A(i_0_), .B(i_5_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n211_), .B(new_new_n316_), .Y(new_new_n317_));
  NA4        g295(.A(new_new_n317_), .B(new_new_n228_), .C(new_new_n315_), .D(i_1_), .Y(new_new_n318_));
  NA3        g296(.A(new_new_n286_), .B(new_new_n282_), .C(new_new_n109_), .Y(new_new_n319_));
  NAi21      g297(.An(i_8_), .B(i_7_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n320_), .B(i_6_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n151_), .B(new_new_n46_), .Y(new_new_n322_));
  NA3        g300(.A(new_new_n322_), .B(new_new_n321_), .C(new_new_n157_), .Y(new_new_n323_));
  NA3        g301(.A(new_new_n323_), .B(new_new_n319_), .C(new_new_n318_), .Y(new_new_n324_));
  OAI210     g302(.A0(new_new_n324_), .A1(new_new_n314_), .B0(i_4_), .Y(new_new_n325_));
  NO2        g303(.A(i_12_), .B(i_10_), .Y(new_new_n326_));
  NOi21      g304(.An(i_5_), .B(i_0_), .Y(new_new_n327_));
  NA4        g305(.A(new_new_n80_), .B(new_new_n36_), .C(new_new_n82_), .D(i_8_), .Y(new_new_n328_));
  NO2        g306(.A(i_6_), .B(i_8_), .Y(new_new_n329_));
  NOi21      g307(.An(i_0_), .B(i_2_), .Y(new_new_n330_));
  AN2        g308(.A(new_new_n330_), .B(new_new_n329_), .Y(new_new_n331_));
  NO2        g309(.A(i_1_), .B(i_7_), .Y(new_new_n332_));
  AO220      g310(.A0(new_new_n332_), .A1(new_new_n331_), .B0(new_new_n321_), .B1(new_new_n229_), .Y(new_new_n333_));
  NA3        g311(.A(new_new_n333_), .B(i_4_), .C(i_5_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(new_new_n325_), .Y(new_new_n335_));
  NO3        g313(.A(new_new_n227_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n336_));
  NO3        g314(.A(new_new_n320_), .B(i_2_), .C(i_1_), .Y(new_new_n337_));
  OAI210     g315(.A0(new_new_n337_), .A1(new_new_n336_), .B0(i_6_), .Y(new_new_n338_));
  NA3        g316(.A(new_new_n246_), .B(new_new_n298_), .C(new_new_n187_), .Y(new_new_n339_));
  AOI210     g317(.A0(new_new_n339_), .A1(new_new_n338_), .B0(new_new_n317_), .Y(new_new_n340_));
  NOi21      g318(.An(new_new_n147_), .B(new_new_n101_), .Y(new_new_n341_));
  NO2        g319(.A(new_new_n341_), .B(new_new_n119_), .Y(new_new_n342_));
  OAI210     g320(.A0(new_new_n342_), .A1(new_new_n340_), .B0(i_3_), .Y(new_new_n343_));
  INV        g321(.A(new_new_n80_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n290_), .B(new_new_n78_), .Y(new_new_n345_));
  NA2        g323(.A(new_new_n345_), .B(new_new_n127_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n89_), .B(new_new_n187_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n347_), .B(new_new_n60_), .Y(new_new_n348_));
  AOI210     g326(.A0(new_new_n348_), .A1(new_new_n346_), .B0(new_new_n344_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n187_), .B(i_9_), .Y(new_new_n350_));
  NA2        g328(.A(new_new_n350_), .B(i_1_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n351_), .B(new_new_n46_), .Y(new_new_n352_));
  NO3        g330(.A(new_new_n352_), .B(new_new_n349_), .C(new_new_n289_), .Y(new_new_n353_));
  AOI210     g331(.A0(new_new_n353_), .A1(new_new_n343_), .B0(new_new_n156_), .Y(new_new_n354_));
  AOI210     g332(.A0(new_new_n335_), .A1(new_new_n309_), .B0(new_new_n354_), .Y(new_new_n355_));
  NOi32      g333(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n356_));
  INV        g334(.A(new_new_n356_), .Y(new_new_n357_));
  NAi21      g335(.An(i_0_), .B(i_6_), .Y(new_new_n358_));
  NAi21      g336(.An(i_1_), .B(i_5_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n359_), .B(new_new_n358_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n360_), .B(new_new_n25_), .Y(new_new_n361_));
  OAI210     g339(.A0(new_new_n361_), .A1(new_new_n153_), .B0(new_new_n240_), .Y(new_new_n362_));
  NAi41      g340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n153_), .B(new_new_n151_), .Y(new_new_n364_));
  NOi32      g342(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n365_));
  NO2        g343(.A(i_1_), .B(new_new_n98_), .Y(new_new_n366_));
  NAi21      g344(.An(i_3_), .B(i_4_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(i_9_), .Y(new_new_n368_));
  AN2        g346(.A(i_6_), .B(i_7_), .Y(new_new_n369_));
  OAI210     g347(.A0(new_new_n369_), .A1(new_new_n366_), .B0(new_new_n368_), .Y(new_new_n370_));
  NA2        g348(.A(i_2_), .B(i_7_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n367_), .B(i_10_), .Y(new_new_n372_));
  NA3        g350(.A(new_new_n372_), .B(new_new_n371_), .C(new_new_n238_), .Y(new_new_n373_));
  AOI210     g351(.A0(new_new_n373_), .A1(new_new_n370_), .B0(new_new_n179_), .Y(new_new_n374_));
  AOI210     g352(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n375_));
  OAI210     g353(.A0(new_new_n375_), .A1(new_new_n182_), .B0(new_new_n372_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n376_), .B(i_5_), .Y(new_new_n377_));
  NO4        g355(.A(new_new_n377_), .B(new_new_n374_), .C(new_new_n364_), .D(new_new_n362_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n378_), .B(new_new_n357_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n56_), .B(new_new_n25_), .Y(new_new_n380_));
  AN2        g358(.A(i_12_), .B(i_5_), .Y(new_new_n381_));
  NO2        g359(.A(i_4_), .B(new_new_n26_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n382_), .B(new_new_n381_), .Y(new_new_n383_));
  NO2        g361(.A(i_11_), .B(i_6_), .Y(new_new_n384_));
  NA3        g362(.A(new_new_n384_), .B(new_new_n322_), .C(new_new_n219_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n385_), .B(new_new_n383_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n237_), .B(i_5_), .Y(new_new_n387_));
  NO2        g365(.A(i_5_), .B(i_10_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n138_), .B(new_new_n45_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(new_new_n237_), .Y(new_new_n390_));
  OAI210     g368(.A0(new_new_n390_), .A1(new_new_n386_), .B0(new_new_n380_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n386_), .B(new_new_n392_), .Y(new_new_n393_));
  NO3        g371(.A(new_new_n82_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n394_));
  NO2        g372(.A(i_11_), .B(i_12_), .Y(new_new_n395_));
  NA2        g373(.A(new_new_n388_), .B(new_new_n231_), .Y(new_new_n396_));
  NA3        g374(.A(new_new_n109_), .B(i_4_), .C(i_11_), .Y(new_new_n397_));
  NO2        g375(.A(new_new_n397_), .B(new_new_n214_), .Y(new_new_n398_));
  NAi21      g376(.An(i_13_), .B(i_0_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(new_new_n234_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n398_), .B(new_new_n400_), .Y(new_new_n401_));
  NA3        g379(.A(new_new_n401_), .B(new_new_n393_), .C(new_new_n391_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n44_), .B(new_new_n219_), .Y(new_new_n403_));
  NO3        g381(.A(i_1_), .B(i_12_), .C(new_new_n82_), .Y(new_new_n404_));
  NO2        g382(.A(i_0_), .B(i_11_), .Y(new_new_n405_));
  INV        g383(.A(i_5_), .Y(new_new_n406_));
  AN2        g384(.A(i_1_), .B(i_6_), .Y(new_new_n407_));
  NOi21      g385(.An(i_2_), .B(i_12_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n408_), .B(new_new_n407_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n409_), .B(new_new_n406_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n136_), .B(i_9_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n411_), .B(i_4_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n410_), .B(new_new_n412_), .Y(new_new_n413_));
  NAi21      g391(.An(i_9_), .B(i_4_), .Y(new_new_n414_));
  OR2        g392(.A(i_13_), .B(i_10_), .Y(new_new_n415_));
  NO3        g393(.A(new_new_n415_), .B(new_new_n112_), .C(new_new_n414_), .Y(new_new_n416_));
  OR2        g394(.A(new_new_n209_), .B(new_new_n208_), .Y(new_new_n417_));
  NO2        g395(.A(new_new_n98_), .B(new_new_n25_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n279_), .B(new_new_n418_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n272_), .B(new_new_n203_), .Y(new_new_n420_));
  OAI220     g398(.A0(new_new_n420_), .A1(new_new_n417_), .B0(new_new_n419_), .B1(new_new_n341_), .Y(new_new_n421_));
  INV        g399(.A(new_new_n421_), .Y(new_new_n422_));
  AOI210     g400(.A0(new_new_n422_), .A1(new_new_n413_), .B0(new_new_n26_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n319_), .B(new_new_n318_), .Y(new_new_n424_));
  AOI220     g402(.A0(new_new_n292_), .A1(new_new_n283_), .B0(new_new_n286_), .B1(new_new_n310_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n425_), .B(new_new_n163_), .Y(new_new_n426_));
  NO2        g404(.A(new_new_n177_), .B(new_new_n82_), .Y(new_new_n427_));
  AOI220     g405(.A0(new_new_n427_), .A1(new_new_n291_), .B0(new_new_n274_), .B1(new_new_n203_), .Y(new_new_n428_));
  NO2        g406(.A(new_new_n428_), .B(new_new_n281_), .Y(new_new_n429_));
  NO3        g407(.A(new_new_n429_), .B(new_new_n426_), .C(new_new_n424_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n190_), .B(new_new_n93_), .Y(new_new_n431_));
  NA3        g409(.A(new_new_n322_), .B(new_new_n157_), .C(new_new_n82_), .Y(new_new_n432_));
  AOI210     g410(.A0(new_new_n432_), .A1(new_new_n431_), .B0(new_new_n320_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n187_), .B(i_10_), .Y(new_new_n434_));
  NA3        g412(.A(new_new_n252_), .B(new_new_n61_), .C(i_2_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n292_), .B(new_new_n229_), .Y(new_new_n436_));
  OAI220     g414(.A0(new_new_n436_), .A1(new_new_n177_), .B0(new_new_n435_), .B1(new_new_n434_), .Y(new_new_n437_));
  NO2        g415(.A(i_3_), .B(new_new_n48_), .Y(new_new_n438_));
  NA3        g416(.A(new_new_n332_), .B(new_new_n331_), .C(new_new_n438_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n312_), .B(new_new_n317_), .Y(new_new_n440_));
  OAI210     g418(.A0(new_new_n440_), .A1(new_new_n183_), .B0(new_new_n439_), .Y(new_new_n441_));
  NO3        g419(.A(new_new_n441_), .B(new_new_n437_), .C(new_new_n433_), .Y(new_new_n442_));
  AOI210     g420(.A0(new_new_n442_), .A1(new_new_n430_), .B0(new_new_n268_), .Y(new_new_n443_));
  NO4        g421(.A(new_new_n443_), .B(new_new_n423_), .C(new_new_n402_), .D(new_new_n379_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n60_), .B(i_4_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n70_), .B(i_13_), .Y(new_new_n446_));
  NO2        g424(.A(i_10_), .B(i_9_), .Y(new_new_n447_));
  NAi21      g425(.An(i_12_), .B(i_8_), .Y(new_new_n448_));
  NO2        g426(.A(new_new_n448_), .B(i_3_), .Y(new_new_n449_));
  INV        g427(.A(i_0_), .Y(new_new_n450_));
  NO3        g428(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n264_), .B(new_new_n94_), .Y(new_new_n452_));
  NA2        g430(.A(new_new_n452_), .B(new_new_n451_), .Y(new_new_n453_));
  NA2        g431(.A(i_8_), .B(i_9_), .Y(new_new_n454_));
  NO3        g432(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n455_));
  NA3        g433(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n456_));
  OR2        g434(.A(new_new_n290_), .B(new_new_n200_), .Y(new_new_n457_));
  BUFFER     g435(.A(new_new_n293_), .Y(new_new_n458_));
  OA220      g436(.A0(new_new_n458_), .A1(new_new_n156_), .B0(new_new_n457_), .B1(new_new_n226_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n93_), .B(i_13_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n427_), .B(new_new_n380_), .Y(new_new_n461_));
  NO2        g439(.A(i_2_), .B(i_13_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n461_), .B(new_new_n460_), .Y(new_new_n463_));
  NO3        g441(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n464_));
  NO2        g442(.A(i_6_), .B(i_7_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n465_), .B(new_new_n464_), .Y(new_new_n466_));
  NO2        g444(.A(i_11_), .B(i_1_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n70_), .B(i_3_), .Y(new_new_n468_));
  NOi21      g446(.An(i_2_), .B(i_7_), .Y(new_new_n469_));
  NAi31      g447(.An(i_11_), .B(new_new_n469_), .C(new_new_n468_), .Y(new_new_n470_));
  INV        g448(.A(new_new_n415_), .Y(new_new_n471_));
  NA3        g449(.A(new_new_n471_), .B(new_new_n445_), .C(new_new_n72_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n470_), .Y(new_new_n473_));
  NO2        g451(.A(i_6_), .B(i_10_), .Y(new_new_n474_));
  NA4        g452(.A(new_new_n474_), .B(new_new_n309_), .C(i_8_), .D(new_new_n231_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n475_), .B(new_new_n149_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n151_), .B(i_3_), .Y(new_new_n478_));
  NAi31      g456(.An(new_new_n477_), .B(new_new_n478_), .C(new_new_n220_), .Y(new_new_n479_));
  NA3        g457(.A(new_new_n392_), .B(new_new_n173_), .C(new_new_n143_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n480_), .B(new_new_n479_), .Y(new_new_n481_));
  NO4        g459(.A(new_new_n481_), .B(new_new_n476_), .C(new_new_n473_), .D(new_new_n463_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n455_), .B(new_new_n388_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n483_), .B(new_new_n218_), .Y(new_new_n484_));
  NAi21      g462(.An(new_new_n209_), .B(new_new_n395_), .Y(new_new_n485_));
  NO2        g463(.A(new_new_n26_), .B(i_5_), .Y(new_new_n486_));
  NO2        g464(.A(i_0_), .B(new_new_n82_), .Y(new_new_n487_));
  NA3        g465(.A(new_new_n487_), .B(new_new_n486_), .C(new_new_n136_), .Y(new_new_n488_));
  OR3        g466(.A(new_new_n299_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n27_), .B(i_10_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n309_), .B(new_new_n233_), .Y(new_new_n492_));
  OAI220     g470(.A0(new_new_n492_), .A1(new_new_n435_), .B0(new_new_n491_), .B1(new_new_n460_), .Y(new_new_n493_));
  NA3        g471(.A(new_new_n302_), .B(new_new_n217_), .C(new_new_n70_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n494_), .B(new_new_n466_), .Y(new_new_n495_));
  NO4        g473(.A(new_new_n495_), .B(new_new_n493_), .C(new_new_n490_), .D(new_new_n484_), .Y(new_new_n496_));
  NA3        g474(.A(new_new_n496_), .B(new_new_n482_), .C(new_new_n459_), .Y(new_new_n497_));
  NA3        g475(.A(new_new_n302_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n498_));
  INV        g476(.A(new_new_n498_), .Y(new_new_n499_));
  BUFFER     g477(.A(new_new_n283_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n500_), .B(new_new_n499_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n309_), .B(new_new_n158_), .Y(new_new_n502_));
  OAI210     g480(.A0(new_new_n502_), .A1(new_new_n226_), .B0(new_new_n303_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n503_), .B(new_new_n321_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n381_), .B(new_new_n219_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n356_), .B(new_new_n70_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n369_), .B(new_new_n365_), .Y(new_new_n507_));
  OR2        g485(.A(new_new_n505_), .B(new_new_n507_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n36_), .B(i_8_), .Y(new_new_n509_));
  NAi41      g487(.An(new_new_n506_), .B(new_new_n474_), .C(new_new_n509_), .D(new_new_n46_), .Y(new_new_n510_));
  AOI210     g488(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n416_), .Y(new_new_n511_));
  NA3        g489(.A(new_new_n511_), .B(new_new_n510_), .C(new_new_n508_), .Y(new_new_n512_));
  INV        g490(.A(new_new_n512_), .Y(new_new_n513_));
  NO2        g491(.A(i_7_), .B(new_new_n193_), .Y(new_new_n514_));
  OR2        g492(.A(new_new_n177_), .B(i_4_), .Y(new_new_n515_));
  NO2        g493(.A(new_new_n515_), .B(new_new_n82_), .Y(new_new_n516_));
  NA2        g494(.A(new_new_n516_), .B(new_new_n514_), .Y(new_new_n517_));
  NA4        g495(.A(new_new_n517_), .B(new_new_n513_), .C(new_new_n504_), .D(new_new_n501_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n387_), .B(new_new_n291_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n383_), .B(new_new_n519_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n997_), .B(new_new_n219_), .Y(new_new_n521_));
  NA2        g499(.A(new_new_n474_), .B(new_new_n27_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n522_), .B(new_new_n521_), .Y(new_new_n523_));
  NOi31      g501(.An(new_new_n312_), .B(new_new_n415_), .C(new_new_n38_), .Y(new_new_n524_));
  OAI210     g502(.A0(new_new_n524_), .A1(new_new_n523_), .B0(new_new_n520_), .Y(new_new_n525_));
  NO2        g503(.A(i_8_), .B(i_7_), .Y(new_new_n526_));
  OAI210     g504(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n527_), .B(new_new_n217_), .Y(new_new_n528_));
  OAI220     g506(.A0(new_new_n46_), .A1(new_new_n515_), .B0(new_new_n528_), .B1(new_new_n237_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n44_), .B(i_10_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n530_), .B(i_6_), .Y(new_new_n531_));
  NA3        g509(.A(new_new_n531_), .B(new_new_n529_), .C(new_new_n526_), .Y(new_new_n532_));
  AOI220     g510(.A0(new_new_n427_), .A1(new_new_n322_), .B0(new_new_n241_), .B1(new_new_n238_), .Y(new_new_n533_));
  OAI220     g511(.A0(new_new_n533_), .A1(new_new_n260_), .B0(new_new_n460_), .B1(new_new_n128_), .Y(new_new_n534_));
  NA2        g512(.A(new_new_n534_), .B(new_new_n263_), .Y(new_new_n535_));
  NOi31      g513(.An(new_new_n286_), .B(new_new_n297_), .C(new_new_n175_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n215_), .B(new_new_n44_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n151_), .B(i_5_), .Y(new_new_n538_));
  NA3        g516(.A(new_new_n538_), .B(new_new_n403_), .C(new_new_n315_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n539_), .B(new_new_n537_), .Y(new_new_n540_));
  OAI210     g518(.A0(new_new_n540_), .A1(new_new_n536_), .B0(new_new_n455_), .Y(new_new_n541_));
  NA4        g519(.A(new_new_n541_), .B(new_new_n535_), .C(new_new_n532_), .D(new_new_n525_), .Y(new_new_n542_));
  NA3        g520(.A(new_new_n211_), .B(new_new_n68_), .C(new_new_n44_), .Y(new_new_n543_));
  NA2        g521(.A(new_new_n279_), .B(new_new_n80_), .Y(new_new_n544_));
  AOI210     g522(.A0(new_new_n543_), .A1(new_new_n346_), .B0(new_new_n544_), .Y(new_new_n545_));
  NA2        g523(.A(new_new_n292_), .B(new_new_n283_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n546_), .B(new_new_n167_), .Y(new_new_n547_));
  NA2        g525(.A(new_new_n217_), .B(new_new_n216_), .Y(new_new_n548_));
  NA2        g526(.A(new_new_n447_), .B(new_new_n215_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n548_), .B(new_new_n549_), .Y(new_new_n550_));
  NO3        g528(.A(new_new_n550_), .B(new_new_n547_), .C(new_new_n545_), .Y(new_new_n551_));
  NO4        g529(.A(new_new_n246_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n552_));
  NO3        g530(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n227_), .B(new_new_n36_), .Y(new_new_n554_));
  AN2        g532(.A(new_new_n554_), .B(new_new_n553_), .Y(new_new_n555_));
  OA210      g533(.A0(new_new_n555_), .A1(new_new_n552_), .B0(new_new_n356_), .Y(new_new_n556_));
  NO2        g534(.A(new_new_n415_), .B(i_1_), .Y(new_new_n557_));
  NOi31      g535(.An(new_new_n557_), .B(new_new_n452_), .C(new_new_n70_), .Y(new_new_n558_));
  AN4        g536(.A(new_new_n558_), .B(new_new_n412_), .C(new_new_n486_), .D(i_2_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n425_), .B(new_new_n171_), .Y(new_new_n560_));
  NO3        g538(.A(new_new_n560_), .B(new_new_n559_), .C(new_new_n556_), .Y(new_new_n561_));
  NOi21      g539(.An(i_10_), .B(i_6_), .Y(new_new_n562_));
  NO2        g540(.A(new_new_n111_), .B(new_new_n23_), .Y(new_new_n563_));
  NA2        g541(.A(new_new_n312_), .B(new_new_n158_), .Y(new_new_n564_));
  AOI220     g542(.A0(new_new_n564_), .A1(new_new_n436_), .B0(new_new_n166_), .B1(new_new_n176_), .Y(new_new_n565_));
  NOi21      g543(.An(new_new_n140_), .B(new_new_n328_), .Y(new_new_n566_));
  NO2        g544(.A(new_new_n566_), .B(new_new_n565_), .Y(new_new_n567_));
  INV        g545(.A(new_new_n315_), .Y(new_new_n568_));
  NO2        g546(.A(i_12_), .B(new_new_n82_), .Y(new_new_n569_));
  NO3        g547(.A(i_4_), .B(new_new_n338_), .C(new_new_n297_), .Y(new_new_n570_));
  OR2        g548(.A(i_2_), .B(i_5_), .Y(new_new_n571_));
  OR2        g549(.A(new_new_n571_), .B(new_new_n407_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n371_), .B(new_new_n238_), .Y(new_new_n573_));
  AOI210     g551(.A0(new_new_n573_), .A1(new_new_n572_), .B0(new_new_n485_), .Y(new_new_n574_));
  NO2        g552(.A(new_new_n574_), .B(new_new_n570_), .Y(new_new_n575_));
  NA4        g553(.A(new_new_n575_), .B(new_new_n567_), .C(new_new_n561_), .D(new_new_n551_), .Y(new_new_n576_));
  NO4        g554(.A(new_new_n576_), .B(new_new_n542_), .C(new_new_n518_), .D(new_new_n497_), .Y(new_new_n577_));
  NA4        g555(.A(new_new_n577_), .B(new_new_n444_), .C(new_new_n355_), .D(new_new_n308_), .Y(mai7));
  NO2        g556(.A(new_new_n89_), .B(new_new_n52_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n474_), .B(new_new_n80_), .Y(new_new_n580_));
  NA2        g558(.A(i_11_), .B(new_new_n187_), .Y(new_new_n581_));
  NA3        g559(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n231_), .B(i_4_), .Y(new_new_n583_));
  NA2        g561(.A(new_new_n583_), .B(i_8_), .Y(new_new_n584_));
  NO2        g562(.A(new_new_n102_), .B(new_new_n582_), .Y(new_new_n585_));
  NA2        g563(.A(i_2_), .B(new_new_n82_), .Y(new_new_n586_));
  OAI210     g564(.A0(new_new_n83_), .A1(new_new_n197_), .B0(new_new_n198_), .Y(new_new_n587_));
  NO2        g565(.A(i_7_), .B(new_new_n37_), .Y(new_new_n588_));
  NA2        g566(.A(i_4_), .B(i_8_), .Y(new_new_n589_));
  AOI210     g567(.A0(new_new_n589_), .A1(new_new_n302_), .B0(new_new_n588_), .Y(new_new_n590_));
  OAI220     g568(.A0(new_new_n590_), .A1(new_new_n586_), .B0(new_new_n587_), .B1(i_13_), .Y(new_new_n591_));
  NO3        g569(.A(new_new_n591_), .B(new_new_n585_), .C(new_new_n579_), .Y(new_new_n592_));
  AOI210     g570(.A0(new_new_n123_), .A1(new_new_n59_), .B0(i_10_), .Y(new_new_n593_));
  AOI210     g571(.A0(new_new_n593_), .A1(new_new_n231_), .B0(new_new_n155_), .Y(new_new_n594_));
  OR2        g572(.A(i_6_), .B(i_10_), .Y(new_new_n595_));
  NO2        g573(.A(new_new_n595_), .B(new_new_n23_), .Y(new_new_n596_));
  OR3        g574(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n597_));
  NO3        g575(.A(new_new_n597_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n598_));
  INV        g576(.A(new_new_n194_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n598_), .B(new_new_n596_), .Y(new_new_n600_));
  OA220      g578(.A0(new_new_n600_), .A1(new_new_n568_), .B0(new_new_n594_), .B1(new_new_n265_), .Y(new_new_n601_));
  AOI210     g579(.A0(new_new_n601_), .A1(new_new_n592_), .B0(new_new_n60_), .Y(new_new_n602_));
  NOi21      g580(.An(i_11_), .B(i_7_), .Y(new_new_n603_));
  AO210      g581(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n604_));
  NO2        g582(.A(new_new_n604_), .B(new_new_n603_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n605_), .B(new_new_n199_), .Y(new_new_n606_));
  NA3        g584(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n606_), .B(new_new_n60_), .Y(new_new_n608_));
  NO3        g586(.A(new_new_n254_), .B(new_new_n201_), .C(new_new_n581_), .Y(new_new_n609_));
  OAI210     g587(.A0(new_new_n609_), .A1(new_new_n220_), .B0(new_new_n60_), .Y(new_new_n610_));
  OR2        g588(.A(new_new_n201_), .B(new_new_n105_), .Y(new_new_n611_));
  NO2        g589(.A(new_new_n60_), .B(i_9_), .Y(new_new_n612_));
  NO2        g590(.A(i_1_), .B(i_12_), .Y(new_new_n613_));
  INV        g591(.A(new_new_n610_), .Y(new_new_n614_));
  OAI210     g592(.A0(new_new_n614_), .A1(new_new_n608_), .B0(i_6_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n607_), .B(new_new_n105_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n616_), .B(new_new_n569_), .Y(new_new_n617_));
  NO2        g595(.A(i_6_), .B(i_11_), .Y(new_new_n618_));
  NA2        g596(.A(new_new_n617_), .B(new_new_n453_), .Y(new_new_n619_));
  NO4        g597(.A(new_new_n208_), .B(new_new_n123_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n620_), .B(new_new_n612_), .Y(new_new_n621_));
  NA2        g599(.A(new_new_n231_), .B(i_6_), .Y(new_new_n622_));
  NO3        g600(.A(new_new_n595_), .B(new_new_n227_), .C(new_new_n23_), .Y(new_new_n623_));
  AOI210     g601(.A0(i_1_), .A1(new_new_n255_), .B0(new_new_n623_), .Y(new_new_n624_));
  OAI210     g602(.A0(new_new_n624_), .A1(new_new_n44_), .B0(new_new_n621_), .Y(new_new_n625_));
  NA3        g603(.A(new_new_n526_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n132_), .B(i_9_), .Y(new_new_n627_));
  NA3        g605(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n46_), .B(i_1_), .Y(new_new_n629_));
  NA3        g607(.A(new_new_n629_), .B(new_new_n264_), .C(new_new_n44_), .Y(new_new_n630_));
  OAI220     g608(.A0(new_new_n630_), .A1(new_new_n628_), .B0(new_new_n627_), .B1(new_new_n996_), .Y(new_new_n631_));
  NA3        g609(.A(new_new_n612_), .B(new_new_n315_), .C(i_6_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n632_), .B(new_new_n23_), .Y(new_new_n633_));
  AOI210     g611(.A0(new_new_n467_), .A1(new_new_n418_), .B0(new_new_n236_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n634_), .B(new_new_n586_), .Y(new_new_n635_));
  NAi21      g613(.An(new_new_n626_), .B(new_new_n88_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n629_), .B(new_new_n264_), .Y(new_new_n637_));
  NO2        g615(.A(i_11_), .B(new_new_n37_), .Y(new_new_n638_));
  NA2        g616(.A(new_new_n638_), .B(new_new_n24_), .Y(new_new_n639_));
  OAI210     g617(.A0(new_new_n639_), .A1(new_new_n637_), .B0(new_new_n636_), .Y(new_new_n640_));
  OR4        g618(.A(new_new_n640_), .B(new_new_n635_), .C(new_new_n633_), .D(new_new_n631_), .Y(new_new_n641_));
  NO3        g619(.A(new_new_n641_), .B(new_new_n625_), .C(new_new_n619_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n231_), .B(new_new_n98_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n643_), .B(new_new_n603_), .Y(new_new_n644_));
  NA2        g622(.A(new_new_n644_), .B(i_1_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n597_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n414_), .B(new_new_n82_), .Y(new_new_n647_));
  NA2        g625(.A(new_new_n646_), .B(new_new_n46_), .Y(new_new_n648_));
  NA2        g626(.A(i_3_), .B(new_new_n187_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n649_), .B(new_new_n111_), .Y(new_new_n650_));
  AN2        g628(.A(new_new_n650_), .B(new_new_n531_), .Y(new_new_n651_));
  NO2        g629(.A(new_new_n227_), .B(new_new_n44_), .Y(new_new_n652_));
  NO3        g630(.A(new_new_n652_), .B(new_new_n305_), .C(new_new_n232_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n112_), .B(new_new_n37_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n654_), .B(i_6_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n82_), .B(i_9_), .Y(new_new_n656_));
  NO2        g634(.A(new_new_n656_), .B(new_new_n60_), .Y(new_new_n657_));
  NO2        g635(.A(new_new_n657_), .B(new_new_n613_), .Y(new_new_n658_));
  NO4        g636(.A(new_new_n658_), .B(new_new_n655_), .C(new_new_n653_), .D(i_4_), .Y(new_new_n659_));
  NA2        g637(.A(i_1_), .B(i_3_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n454_), .B(new_new_n89_), .Y(new_new_n661_));
  AOI210     g639(.A0(new_new_n652_), .A1(new_new_n562_), .B0(new_new_n661_), .Y(new_new_n662_));
  NO2        g640(.A(new_new_n662_), .B(new_new_n660_), .Y(new_new_n663_));
  NO3        g641(.A(new_new_n663_), .B(new_new_n659_), .C(new_new_n651_), .Y(new_new_n664_));
  NA4        g642(.A(new_new_n664_), .B(new_new_n648_), .C(new_new_n642_), .D(new_new_n615_), .Y(new_new_n665_));
  NO3        g643(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n666_));
  NOi21      g644(.An(new_new_n666_), .B(i_10_), .Y(new_new_n667_));
  OA210      g645(.A0(new_new_n667_), .A1(new_new_n239_), .B0(new_new_n82_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n369_), .B(new_new_n368_), .Y(new_new_n669_));
  NA3        g647(.A(new_new_n474_), .B(new_new_n509_), .C(new_new_n46_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n670_), .B(new_new_n669_), .Y(new_new_n671_));
  OAI210     g649(.A0(new_new_n671_), .A1(new_new_n668_), .B0(i_1_), .Y(new_new_n672_));
  AOI210     g650(.A0(new_new_n264_), .A1(new_new_n94_), .B0(i_1_), .Y(new_new_n673_));
  NO2        g651(.A(new_new_n367_), .B(i_2_), .Y(new_new_n674_));
  NA2        g652(.A(new_new_n674_), .B(new_new_n673_), .Y(new_new_n675_));
  OAI210     g653(.A0(new_new_n632_), .A1(new_new_n448_), .B0(new_new_n675_), .Y(new_new_n676_));
  INV        g654(.A(new_new_n676_), .Y(new_new_n677_));
  AOI210     g655(.A0(new_new_n677_), .A1(new_new_n672_), .B0(i_13_), .Y(new_new_n678_));
  OR2        g656(.A(i_11_), .B(i_7_), .Y(new_new_n679_));
  NO2        g657(.A(new_new_n52_), .B(i_12_), .Y(new_new_n680_));
  INV        g658(.A(new_new_n680_), .Y(new_new_n681_));
  NO2        g659(.A(new_new_n469_), .B(new_new_n24_), .Y(new_new_n682_));
  AOI220     g660(.A0(new_new_n682_), .A1(new_new_n647_), .B0(new_new_n239_), .B1(new_new_n126_), .Y(new_new_n683_));
  OAI220     g661(.A0(new_new_n683_), .A1(new_new_n41_), .B0(new_new_n681_), .B1(new_new_n89_), .Y(new_new_n684_));
  INV        g662(.A(new_new_n684_), .Y(new_new_n685_));
  NA2        g663(.A(new_new_n384_), .B(new_new_n629_), .Y(new_new_n686_));
  NO2        g664(.A(new_new_n686_), .B(new_new_n237_), .Y(new_new_n687_));
  AOI210     g665(.A0(new_new_n448_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n688_));
  NOi31      g666(.An(new_new_n688_), .B(new_new_n580_), .C(new_new_n44_), .Y(new_new_n689_));
  NA2        g667(.A(new_new_n122_), .B(i_13_), .Y(new_new_n690_));
  NO2        g668(.A(new_new_n628_), .B(new_new_n111_), .Y(new_new_n691_));
  INV        g669(.A(new_new_n691_), .Y(new_new_n692_));
  OAI220     g670(.A0(new_new_n692_), .A1(new_new_n68_), .B0(new_new_n690_), .B1(new_new_n673_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n26_), .B(new_new_n187_), .Y(new_new_n694_));
  NA2        g672(.A(new_new_n694_), .B(i_7_), .Y(new_new_n695_));
  NO3        g673(.A(new_new_n469_), .B(new_new_n231_), .C(new_new_n82_), .Y(new_new_n696_));
  NA2        g674(.A(new_new_n696_), .B(new_new_n695_), .Y(new_new_n697_));
  AOI220     g675(.A0(new_new_n384_), .A1(new_new_n629_), .B0(new_new_n88_), .B1(new_new_n99_), .Y(new_new_n698_));
  OAI220     g676(.A0(new_new_n698_), .A1(new_new_n584_), .B0(new_new_n697_), .B1(new_new_n599_), .Y(new_new_n699_));
  NO4        g677(.A(new_new_n699_), .B(new_new_n693_), .C(new_new_n689_), .D(new_new_n687_), .Y(new_new_n700_));
  OR2        g678(.A(i_11_), .B(i_6_), .Y(new_new_n701_));
  NA3        g679(.A(new_new_n583_), .B(new_new_n694_), .C(i_7_), .Y(new_new_n702_));
  AOI210     g680(.A0(new_new_n702_), .A1(new_new_n692_), .B0(new_new_n701_), .Y(new_new_n703_));
  NA3        g681(.A(new_new_n408_), .B(new_new_n588_), .C(new_new_n94_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n618_), .B(i_13_), .Y(new_new_n705_));
  NA2        g683(.A(new_new_n99_), .B(new_new_n694_), .Y(new_new_n706_));
  NAi21      g684(.An(i_11_), .B(i_12_), .Y(new_new_n707_));
  NOi41      g685(.An(new_new_n107_), .B(new_new_n707_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n708_), .B(new_new_n706_), .Y(new_new_n709_));
  NA3        g687(.A(new_new_n709_), .B(new_new_n705_), .C(new_new_n704_), .Y(new_new_n710_));
  OAI210     g688(.A0(new_new_n710_), .A1(new_new_n703_), .B0(new_new_n60_), .Y(new_new_n711_));
  NO2        g689(.A(i_2_), .B(i_12_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n366_), .B(new_new_n712_), .Y(new_new_n713_));
  NA2        g691(.A(i_8_), .B(new_new_n25_), .Y(new_new_n714_));
  NO3        g692(.A(new_new_n714_), .B(new_new_n382_), .C(new_new_n583_), .Y(new_new_n715_));
  OAI210     g693(.A0(new_new_n715_), .A1(new_new_n368_), .B0(new_new_n366_), .Y(new_new_n716_));
  NO2        g694(.A(new_new_n123_), .B(i_2_), .Y(new_new_n717_));
  NA2        g695(.A(new_new_n717_), .B(new_new_n613_), .Y(new_new_n718_));
  NA3        g696(.A(new_new_n718_), .B(new_new_n716_), .C(new_new_n713_), .Y(new_new_n719_));
  NA3        g697(.A(new_new_n719_), .B(new_new_n45_), .C(new_new_n219_), .Y(new_new_n720_));
  NA4        g698(.A(new_new_n720_), .B(new_new_n711_), .C(new_new_n700_), .D(new_new_n685_), .Y(new_new_n721_));
  OR4        g699(.A(new_new_n721_), .B(new_new_n678_), .C(new_new_n665_), .D(new_new_n602_), .Y(mai5));
  NA2        g700(.A(new_new_n644_), .B(new_new_n267_), .Y(new_new_n723_));
  AN2        g701(.A(new_new_n24_), .B(i_10_), .Y(new_new_n724_));
  NA3        g702(.A(new_new_n724_), .B(new_new_n712_), .C(new_new_n105_), .Y(new_new_n725_));
  NO2        g703(.A(new_new_n584_), .B(i_11_), .Y(new_new_n726_));
  NA2        g704(.A(new_new_n83_), .B(new_new_n726_), .Y(new_new_n727_));
  NA3        g705(.A(new_new_n727_), .B(new_new_n725_), .C(new_new_n723_), .Y(new_new_n728_));
  NO3        g706(.A(i_11_), .B(new_new_n231_), .C(i_13_), .Y(new_new_n729_));
  NO2        g707(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n730_));
  NA2        g708(.A(i_12_), .B(i_8_), .Y(new_new_n731_));
  OAI210     g709(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n731_), .Y(new_new_n732_));
  INV        g710(.A(new_new_n447_), .Y(new_new_n733_));
  AOI220     g711(.A0(new_new_n315_), .A1(new_new_n563_), .B0(new_new_n732_), .B1(new_new_n730_), .Y(new_new_n734_));
  INV        g712(.A(new_new_n734_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n735_), .B(new_new_n728_), .Y(new_new_n736_));
  INV        g714(.A(new_new_n165_), .Y(new_new_n737_));
  INV        g715(.A(new_new_n239_), .Y(new_new_n738_));
  OAI210     g716(.A0(new_new_n674_), .A1(new_new_n449_), .B0(new_new_n107_), .Y(new_new_n739_));
  AOI210     g717(.A0(new_new_n739_), .A1(new_new_n738_), .B0(new_new_n737_), .Y(new_new_n740_));
  NO2        g718(.A(new_new_n454_), .B(new_new_n26_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n741_), .B(new_new_n418_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n742_), .B(i_2_), .Y(new_new_n743_));
  INV        g721(.A(new_new_n743_), .Y(new_new_n744_));
  AOI210     g722(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n415_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n745_), .A1(new_new_n744_), .B0(new_new_n740_), .Y(new_new_n746_));
  NO2        g724(.A(new_new_n184_), .B(new_new_n120_), .Y(new_new_n747_));
  OAI210     g725(.A0(new_new_n747_), .A1(new_new_n730_), .B0(i_2_), .Y(new_new_n748_));
  INV        g726(.A(new_new_n166_), .Y(new_new_n749_));
  NO3        g727(.A(new_new_n604_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n750_));
  AOI210     g728(.A0(new_new_n749_), .A1(new_new_n83_), .B0(new_new_n750_), .Y(new_new_n751_));
  AOI210     g729(.A0(new_new_n751_), .A1(new_new_n748_), .B0(new_new_n187_), .Y(new_new_n752_));
  OA210      g730(.A0(new_new_n605_), .A1(new_new_n121_), .B0(i_13_), .Y(new_new_n753_));
  NA2        g731(.A(new_new_n145_), .B(new_new_n581_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n754_), .B(new_new_n371_), .Y(new_new_n755_));
  AOI210     g733(.A0(new_new_n201_), .A1(new_new_n142_), .B0(new_new_n509_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n756_), .B(new_new_n418_), .Y(new_new_n757_));
  NO2        g735(.A(new_new_n99_), .B(new_new_n44_), .Y(new_new_n758_));
  INV        g736(.A(new_new_n298_), .Y(new_new_n759_));
  NA4        g737(.A(new_new_n759_), .B(new_new_n302_), .C(new_new_n119_), .D(new_new_n42_), .Y(new_new_n760_));
  OAI210     g738(.A0(new_new_n760_), .A1(new_new_n758_), .B0(new_new_n757_), .Y(new_new_n761_));
  NO4        g739(.A(new_new_n761_), .B(new_new_n755_), .C(new_new_n753_), .D(new_new_n752_), .Y(new_new_n762_));
  NA2        g740(.A(new_new_n563_), .B(new_new_n28_), .Y(new_new_n763_));
  NA2        g741(.A(new_new_n729_), .B(new_new_n271_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n764_), .B(new_new_n763_), .Y(new_new_n765_));
  NO2        g743(.A(new_new_n59_), .B(i_12_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n766_), .B(new_new_n121_), .Y(new_new_n767_));
  NO2        g745(.A(new_new_n767_), .B(new_new_n581_), .Y(new_new_n768_));
  AOI220     g746(.A0(new_new_n768_), .A1(new_new_n36_), .B0(new_new_n765_), .B1(new_new_n46_), .Y(new_new_n769_));
  NA4        g747(.A(new_new_n769_), .B(new_new_n762_), .C(new_new_n746_), .D(new_new_n736_), .Y(mai6));
  NO3        g748(.A(new_new_n250_), .B(new_new_n304_), .C(i_1_), .Y(new_new_n771_));
  NO2        g749(.A(new_new_n179_), .B(new_new_n133_), .Y(new_new_n772_));
  OAI210     g750(.A0(new_new_n772_), .A1(new_new_n771_), .B0(new_new_n717_), .Y(new_new_n773_));
  NO2        g751(.A(new_new_n214_), .B(new_new_n477_), .Y(new_new_n774_));
  INV        g752(.A(new_new_n327_), .Y(new_new_n775_));
  AO210      g753(.A0(new_new_n775_), .A1(new_new_n773_), .B0(i_12_), .Y(new_new_n776_));
  NA2        g754(.A(new_new_n372_), .B(new_new_n332_), .Y(new_new_n777_));
  NA2        g755(.A(new_new_n569_), .B(new_new_n60_), .Y(new_new_n778_));
  NA2        g756(.A(new_new_n667_), .B(new_new_n68_), .Y(new_new_n779_));
  NA3        g757(.A(new_new_n779_), .B(new_new_n778_), .C(new_new_n777_), .Y(new_new_n780_));
  NA2        g758(.A(new_new_n780_), .B(new_new_n70_), .Y(new_new_n781_));
  INV        g759(.A(new_new_n326_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n72_), .B(new_new_n126_), .Y(new_new_n783_));
  INV        g761(.A(new_new_n119_), .Y(new_new_n784_));
  NA2        g762(.A(new_new_n784_), .B(new_new_n46_), .Y(new_new_n785_));
  AOI210     g763(.A0(new_new_n785_), .A1(new_new_n783_), .B0(new_new_n782_), .Y(new_new_n786_));
  NO2        g764(.A(new_new_n507_), .B(new_new_n179_), .Y(new_new_n787_));
  NO2        g765(.A(new_new_n32_), .B(i_11_), .Y(new_new_n788_));
  NA3        g766(.A(new_new_n788_), .B(new_new_n465_), .C(new_new_n388_), .Y(new_new_n789_));
  NAi32      g767(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n790_));
  NO2        g768(.A(new_new_n701_), .B(new_new_n790_), .Y(new_new_n791_));
  OAI210     g769(.A0(new_new_n666_), .A1(new_new_n554_), .B0(new_new_n553_), .Y(new_new_n792_));
  NAi31      g770(.An(new_new_n791_), .B(new_new_n792_), .C(new_new_n789_), .Y(new_new_n793_));
  OR3        g771(.A(new_new_n793_), .B(new_new_n787_), .C(new_new_n786_), .Y(new_new_n794_));
  NO2        g772(.A(new_new_n679_), .B(i_2_), .Y(new_new_n795_));
  NA2        g773(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n796_));
  NO2        g774(.A(new_new_n796_), .B(new_new_n407_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n797_), .B(new_new_n795_), .Y(new_new_n798_));
  AO210      g776(.A0(new_new_n360_), .A1(new_new_n350_), .B0(new_new_n394_), .Y(new_new_n799_));
  NA3        g777(.A(new_new_n799_), .B(new_new_n251_), .C(i_7_), .Y(new_new_n800_));
  OR2        g778(.A(new_new_n605_), .B(new_new_n449_), .Y(new_new_n801_));
  NA3        g779(.A(new_new_n801_), .B(new_new_n141_), .C(new_new_n66_), .Y(new_new_n802_));
  AO210      g780(.A0(new_new_n483_), .A1(new_new_n733_), .B0(new_new_n36_), .Y(new_new_n803_));
  NA4        g781(.A(new_new_n803_), .B(new_new_n802_), .C(new_new_n800_), .D(new_new_n798_), .Y(new_new_n804_));
  NO2        g782(.A(i_6_), .B(i_11_), .Y(new_new_n805_));
  AOI220     g783(.A0(new_new_n805_), .A1(new_new_n553_), .B0(new_new_n774_), .B1(new_new_n695_), .Y(new_new_n806_));
  NA3        g784(.A(new_new_n371_), .B(new_new_n233_), .C(new_new_n141_), .Y(new_new_n807_));
  NA2        g785(.A(new_new_n394_), .B(new_new_n67_), .Y(new_new_n808_));
  NA4        g786(.A(new_new_n808_), .B(new_new_n807_), .C(new_new_n806_), .D(new_new_n587_), .Y(new_new_n809_));
  AOI210     g787(.A0(new_new_n449_), .A1(new_new_n447_), .B0(new_new_n552_), .Y(new_new_n810_));
  NO2        g788(.A(new_new_n595_), .B(new_new_n99_), .Y(new_new_n811_));
  OAI210     g789(.A0(new_new_n811_), .A1(new_new_n108_), .B0(new_new_n405_), .Y(new_new_n812_));
  INV        g790(.A(new_new_n238_), .Y(new_new_n813_));
  INV        g791(.A(new_new_n572_), .Y(new_new_n814_));
  NA3        g792(.A(new_new_n814_), .B(new_new_n326_), .C(i_7_), .Y(new_new_n815_));
  NA3        g793(.A(new_new_n815_), .B(new_new_n812_), .C(new_new_n810_), .Y(new_new_n816_));
  NO4        g794(.A(new_new_n816_), .B(new_new_n809_), .C(new_new_n804_), .D(new_new_n794_), .Y(new_new_n817_));
  NA4        g795(.A(new_new_n817_), .B(new_new_n781_), .C(new_new_n776_), .D(new_new_n378_), .Y(mai3));
  NA2        g796(.A(i_6_), .B(i_7_), .Y(new_new_n819_));
  NO2        g797(.A(new_new_n819_), .B(i_0_), .Y(new_new_n820_));
  NO2        g798(.A(i_11_), .B(new_new_n231_), .Y(new_new_n821_));
  OAI210     g799(.A0(new_new_n820_), .A1(new_new_n286_), .B0(new_new_n821_), .Y(new_new_n822_));
  NO2        g800(.A(new_new_n822_), .B(new_new_n187_), .Y(new_new_n823_));
  NO3        g801(.A(new_new_n450_), .B(new_new_n86_), .C(new_new_n44_), .Y(new_new_n824_));
  OA210      g802(.A0(new_new_n824_), .A1(new_new_n823_), .B0(new_new_n168_), .Y(new_new_n825_));
  NA2        g803(.A(new_new_n807_), .B(new_new_n370_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n826_), .B(new_new_n40_), .Y(new_new_n827_));
  NO3        g805(.A(new_new_n611_), .B(new_new_n454_), .C(new_new_n126_), .Y(new_new_n828_));
  AN2        g806(.A(new_new_n452_), .B(new_new_n53_), .Y(new_new_n829_));
  NO2        g807(.A(new_new_n829_), .B(new_new_n828_), .Y(new_new_n830_));
  AOI210     g808(.A0(new_new_n830_), .A1(new_new_n827_), .B0(new_new_n48_), .Y(new_new_n831_));
  NO4        g809(.A(new_new_n375_), .B(new_new_n381_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n832_));
  NA2        g810(.A(new_new_n688_), .B(new_new_n656_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n330_), .B(new_new_n438_), .Y(new_new_n834_));
  OAI220     g812(.A0(new_new_n834_), .A1(new_new_n833_), .B0(new_new_n999_), .B1(new_new_n60_), .Y(new_new_n835_));
  NOi21      g813(.An(i_5_), .B(i_9_), .Y(new_new_n836_));
  NA2        g814(.A(new_new_n836_), .B(new_new_n446_), .Y(new_new_n837_));
  BUFFER     g815(.A(new_new_n264_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n838_), .B(new_new_n467_), .Y(new_new_n839_));
  NO3        g817(.A(new_new_n411_), .B(new_new_n264_), .C(new_new_n70_), .Y(new_new_n840_));
  NO2        g818(.A(new_new_n169_), .B(new_new_n142_), .Y(new_new_n841_));
  AOI210     g819(.A0(new_new_n841_), .A1(new_new_n238_), .B0(new_new_n840_), .Y(new_new_n842_));
  OAI220     g820(.A0(new_new_n842_), .A1(new_new_n175_), .B0(new_new_n839_), .B1(new_new_n837_), .Y(new_new_n843_));
  NO4        g821(.A(new_new_n843_), .B(new_new_n835_), .C(new_new_n831_), .D(new_new_n825_), .Y(new_new_n844_));
  NA2        g822(.A(new_new_n179_), .B(new_new_n24_), .Y(new_new_n845_));
  NA2        g823(.A(new_new_n309_), .B(new_new_n124_), .Y(new_new_n846_));
  NAi21      g824(.An(new_new_n156_), .B(new_new_n438_), .Y(new_new_n847_));
  OAI220     g825(.A0(new_new_n847_), .A1(new_new_n813_), .B0(new_new_n846_), .B1(new_new_n396_), .Y(new_new_n848_));
  INV        g826(.A(new_new_n848_), .Y(new_new_n849_));
  NO4        g827(.A(new_new_n571_), .B(new_new_n208_), .C(new_new_n415_), .D(new_new_n407_), .Y(new_new_n850_));
  NA2        g828(.A(new_new_n729_), .B(new_new_n327_), .Y(new_new_n851_));
  AOI210     g829(.A0(new_new_n474_), .A1(new_new_n83_), .B0(new_new_n55_), .Y(new_new_n852_));
  OAI220     g830(.A0(new_new_n852_), .A1(new_new_n851_), .B0(new_new_n639_), .B1(new_new_n528_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n248_), .B(new_new_n147_), .Y(new_new_n854_));
  NA2        g832(.A(i_0_), .B(i_10_), .Y(new_new_n855_));
  AN2        g833(.A(new_new_n854_), .B(i_6_), .Y(new_new_n856_));
  AOI220     g834(.A0(new_new_n330_), .A1(new_new_n95_), .B0(new_new_n179_), .B1(new_new_n80_), .Y(new_new_n857_));
  NA2        g835(.A(new_new_n557_), .B(i_4_), .Y(new_new_n858_));
  NA2        g836(.A(new_new_n182_), .B(new_new_n197_), .Y(new_new_n859_));
  OAI220     g837(.A0(new_new_n859_), .A1(new_new_n851_), .B0(new_new_n858_), .B1(new_new_n857_), .Y(new_new_n860_));
  NO3        g838(.A(new_new_n860_), .B(new_new_n856_), .C(new_new_n853_), .Y(new_new_n861_));
  NA2        g839(.A(new_new_n861_), .B(new_new_n849_), .Y(new_new_n862_));
  NA2        g840(.A(new_new_n392_), .B(new_new_n173_), .Y(new_new_n863_));
  NA2        g841(.A(new_new_n863_), .B(new_new_n154_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n169_), .B(i_0_), .Y(new_new_n865_));
  INV        g843(.A(new_new_n865_), .Y(new_new_n866_));
  NA2        g844(.A(new_new_n465_), .B(new_new_n225_), .Y(new_new_n867_));
  INV        g845(.A(new_new_n404_), .Y(new_new_n868_));
  OAI220     g846(.A0(new_new_n868_), .A1(new_new_n837_), .B0(new_new_n867_), .B1(new_new_n866_), .Y(new_new_n869_));
  NO2        g847(.A(new_new_n869_), .B(new_new_n864_), .Y(new_new_n870_));
  NA2        g848(.A(new_new_n638_), .B(new_new_n116_), .Y(new_new_n871_));
  NO2        g849(.A(i_6_), .B(new_new_n871_), .Y(new_new_n872_));
  AOI210     g850(.A0(new_new_n448_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n873_));
  NA2        g851(.A(new_new_n165_), .B(new_new_n100_), .Y(new_new_n874_));
  NOi32      g852(.An(new_new_n873_), .Bn(new_new_n182_), .C(new_new_n874_), .Y(new_new_n875_));
  NO2        g853(.A(new_new_n875_), .B(new_new_n872_), .Y(new_new_n876_));
  NOi21      g854(.An(i_7_), .B(i_5_), .Y(new_new_n877_));
  NOi31      g855(.An(new_new_n877_), .B(i_0_), .C(new_new_n707_), .Y(new_new_n878_));
  NA3        g856(.A(new_new_n878_), .B(new_new_n382_), .C(i_6_), .Y(new_new_n879_));
  OA210      g857(.A0(new_new_n874_), .A1(new_new_n507_), .B0(new_new_n879_), .Y(new_new_n880_));
  NO3        g858(.A(new_new_n399_), .B(new_new_n363_), .C(new_new_n359_), .Y(new_new_n881_));
  NO2        g859(.A(new_new_n258_), .B(new_new_n316_), .Y(new_new_n882_));
  NO2        g860(.A(new_new_n707_), .B(new_new_n253_), .Y(new_new_n883_));
  AOI210     g861(.A0(new_new_n883_), .A1(new_new_n882_), .B0(new_new_n881_), .Y(new_new_n884_));
  NA4        g862(.A(new_new_n884_), .B(new_new_n880_), .C(new_new_n876_), .D(new_new_n870_), .Y(new_new_n885_));
  NO2        g863(.A(new_new_n845_), .B(new_new_n234_), .Y(new_new_n886_));
  AN2        g864(.A(new_new_n329_), .B(new_new_n327_), .Y(new_new_n887_));
  AN2        g865(.A(new_new_n887_), .B(new_new_n841_), .Y(new_new_n888_));
  OAI210     g866(.A0(new_new_n888_), .A1(new_new_n886_), .B0(i_10_), .Y(new_new_n889_));
  OA210      g867(.A0(new_new_n465_), .A1(new_new_n217_), .B0(new_new_n464_), .Y(new_new_n890_));
  NA3        g868(.A(new_new_n464_), .B(new_new_n408_), .C(new_new_n45_), .Y(new_new_n891_));
  INV        g869(.A(new_new_n891_), .Y(new_new_n892_));
  INV        g870(.A(new_new_n181_), .Y(new_new_n893_));
  AOI220     g871(.A0(new_new_n893_), .A1(new_new_n465_), .B0(new_new_n892_), .B1(new_new_n70_), .Y(new_new_n894_));
  NO2        g872(.A(new_new_n72_), .B(new_new_n731_), .Y(new_new_n895_));
  INV        g873(.A(new_new_n895_), .Y(new_new_n896_));
  NO2        g874(.A(new_new_n896_), .B(new_new_n47_), .Y(new_new_n897_));
  NO2        g875(.A(new_new_n582_), .B(new_new_n102_), .Y(new_new_n898_));
  NA2        g876(.A(new_new_n898_), .B(i_0_), .Y(new_new_n899_));
  NO2        g877(.A(new_new_n899_), .B(new_new_n82_), .Y(new_new_n900_));
  NO3        g878(.A(new_new_n900_), .B(new_new_n897_), .C(new_new_n512_), .Y(new_new_n901_));
  NA3        g879(.A(new_new_n901_), .B(new_new_n894_), .C(new_new_n889_), .Y(new_new_n902_));
  NO3        g880(.A(new_new_n902_), .B(new_new_n885_), .C(new_new_n862_), .Y(new_new_n903_));
  NO2        g881(.A(i_0_), .B(new_new_n707_), .Y(new_new_n904_));
  NA2        g882(.A(new_new_n70_), .B(new_new_n44_), .Y(new_new_n905_));
  NA2        g883(.A(new_new_n855_), .B(new_new_n905_), .Y(new_new_n906_));
  NO3        g884(.A(new_new_n102_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n907_));
  AO220      g885(.A0(new_new_n907_), .A1(new_new_n906_), .B0(new_new_n904_), .B1(new_new_n168_), .Y(new_new_n908_));
  AOI210     g886(.A0(new_new_n778_), .A1(new_new_n669_), .B0(new_new_n874_), .Y(new_new_n909_));
  AOI210     g887(.A0(new_new_n908_), .A1(new_new_n347_), .B0(new_new_n909_), .Y(new_new_n910_));
  NO2        g888(.A(new_new_n792_), .B(new_new_n399_), .Y(new_new_n911_));
  NA3        g889(.A(new_new_n820_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n912_));
  NA2        g890(.A(new_new_n821_), .B(i_9_), .Y(new_new_n913_));
  AOI210     g891(.A0(new_new_n912_), .A1(new_new_n488_), .B0(new_new_n913_), .Y(new_new_n914_));
  NA2        g892(.A(new_new_n238_), .B(new_new_n224_), .Y(new_new_n915_));
  NO2        g893(.A(new_new_n915_), .B(new_new_n147_), .Y(new_new_n916_));
  NO3        g894(.A(new_new_n916_), .B(new_new_n914_), .C(new_new_n911_), .Y(new_new_n917_));
  NA2        g895(.A(new_new_n917_), .B(new_new_n910_), .Y(new_new_n918_));
  NA2        g896(.A(new_new_n887_), .B(new_new_n371_), .Y(new_new_n919_));
  AOI210     g897(.A0(new_new_n297_), .A1(new_new_n156_), .B0(new_new_n919_), .Y(new_new_n920_));
  NA3        g898(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n921_));
  NA2        g899(.A(i_5_), .B(new_new_n478_), .Y(new_new_n922_));
  AOI210     g900(.A0(new_new_n921_), .A1(new_new_n156_), .B0(new_new_n922_), .Y(new_new_n923_));
  NO2        g901(.A(new_new_n923_), .B(new_new_n920_), .Y(new_new_n924_));
  NO3        g902(.A(new_new_n855_), .B(new_new_n836_), .C(new_new_n184_), .Y(new_new_n925_));
  AOI220     g903(.A0(new_new_n925_), .A1(i_11_), .B0(new_new_n558_), .B1(new_new_n72_), .Y(new_new_n926_));
  NO3        g904(.A(new_new_n202_), .B(new_new_n381_), .C(i_0_), .Y(new_new_n927_));
  OAI210     g905(.A0(new_new_n927_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n928_));
  INV        g906(.A(new_new_n211_), .Y(new_new_n929_));
  OAI220     g907(.A0(new_new_n521_), .A1(new_new_n133_), .B0(new_new_n622_), .B1(new_new_n599_), .Y(new_new_n930_));
  NA3        g908(.A(new_new_n930_), .B(i_7_), .C(new_new_n929_), .Y(new_new_n931_));
  NA4        g909(.A(new_new_n931_), .B(new_new_n928_), .C(new_new_n926_), .D(new_new_n924_), .Y(new_new_n932_));
  NA2        g910(.A(new_new_n350_), .B(new_new_n170_), .Y(new_new_n933_));
  OR2        g911(.A(new_new_n933_), .B(new_new_n1000_), .Y(new_new_n934_));
  AOI210     g912(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n169_), .Y(new_new_n935_));
  NA2        g913(.A(new_new_n935_), .B(new_new_n890_), .Y(new_new_n936_));
  NA3        g914(.A(new_new_n388_), .B(new_new_n331_), .C(new_new_n215_), .Y(new_new_n937_));
  INV        g915(.A(new_new_n937_), .Y(new_new_n938_));
  NOi31      g916(.An(new_new_n387_), .B(new_new_n905_), .C(new_new_n234_), .Y(new_new_n939_));
  NO2        g917(.A(new_new_n939_), .B(new_new_n938_), .Y(new_new_n940_));
  NA3        g918(.A(new_new_n940_), .B(new_new_n936_), .C(new_new_n934_), .Y(new_new_n941_));
  NA3        g919(.A(new_new_n302_), .B(i_5_), .C(new_new_n187_), .Y(new_new_n942_));
  NAi31      g920(.An(new_new_n236_), .B(new_new_n942_), .C(new_new_n237_), .Y(new_new_n943_));
  NO4        g921(.A(new_new_n234_), .B(new_new_n202_), .C(i_0_), .D(i_12_), .Y(new_new_n944_));
  NA2        g922(.A(new_new_n944_), .B(new_new_n943_), .Y(new_new_n945_));
  AN2        g923(.A(new_new_n855_), .B(new_new_n147_), .Y(new_new_n946_));
  NO4        g924(.A(new_new_n946_), .B(i_12_), .C(new_new_n626_), .D(new_new_n126_), .Y(new_new_n947_));
  NA2        g925(.A(new_new_n947_), .B(new_new_n211_), .Y(new_new_n948_));
  NA3        g926(.A(new_new_n95_), .B(new_new_n562_), .C(i_11_), .Y(new_new_n949_));
  NA2        g927(.A(new_new_n877_), .B(new_new_n462_), .Y(new_new_n950_));
  NA2        g928(.A(new_new_n61_), .B(new_new_n98_), .Y(new_new_n951_));
  OAI220     g929(.A0(new_new_n951_), .A1(new_new_n942_), .B0(new_new_n950_), .B1(new_new_n657_), .Y(new_new_n952_));
  NA2        g930(.A(new_new_n952_), .B(new_new_n865_), .Y(new_new_n953_));
  NA3        g931(.A(new_new_n953_), .B(new_new_n948_), .C(new_new_n945_), .Y(new_new_n954_));
  NO4        g932(.A(new_new_n954_), .B(new_new_n941_), .C(new_new_n932_), .D(new_new_n918_), .Y(new_new_n955_));
  OAI210     g933(.A0(new_new_n795_), .A1(new_new_n788_), .B0(new_new_n37_), .Y(new_new_n956_));
  NA3        g934(.A(new_new_n873_), .B(new_new_n366_), .C(i_5_), .Y(new_new_n957_));
  NA3        g935(.A(new_new_n957_), .B(new_new_n956_), .C(new_new_n594_), .Y(new_new_n958_));
  NA2        g936(.A(new_new_n958_), .B(new_new_n199_), .Y(new_new_n959_));
  BUFFER     g937(.A(new_new_n367_), .Y(new_new_n960_));
  NA2        g938(.A(new_new_n180_), .B(new_new_n182_), .Y(new_new_n961_));
  AO210      g939(.A0(new_new_n960_), .A1(new_new_n33_), .B0(new_new_n961_), .Y(new_new_n962_));
  OAI210     g940(.A0(new_new_n598_), .A1(new_new_n596_), .B0(new_new_n315_), .Y(new_new_n963_));
  NAi31      g941(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n964_));
  AOI210     g942(.A0(new_new_n112_), .A1(new_new_n67_), .B0(new_new_n964_), .Y(new_new_n965_));
  NO2        g943(.A(new_new_n965_), .B(new_new_n623_), .Y(new_new_n966_));
  NA3        g944(.A(new_new_n966_), .B(new_new_n963_), .C(new_new_n962_), .Y(new_new_n967_));
  NO2        g945(.A(new_new_n456_), .B(new_new_n264_), .Y(new_new_n968_));
  NO4        g946(.A(new_new_n227_), .B(new_new_n139_), .C(new_new_n660_), .D(new_new_n37_), .Y(new_new_n969_));
  NO3        g947(.A(new_new_n969_), .B(new_new_n968_), .C(new_new_n850_), .Y(new_new_n970_));
  OAI210     g948(.A0(new_new_n949_), .A1(new_new_n142_), .B0(new_new_n970_), .Y(new_new_n971_));
  AOI210     g949(.A0(new_new_n967_), .A1(new_new_n48_), .B0(new_new_n971_), .Y(new_new_n972_));
  AOI210     g950(.A0(new_new_n972_), .A1(new_new_n959_), .B0(new_new_n70_), .Y(new_new_n973_));
  NO2        g951(.A(new_new_n555_), .B(new_new_n377_), .Y(new_new_n974_));
  NO2        g952(.A(new_new_n974_), .B(new_new_n737_), .Y(new_new_n975_));
  INV        g953(.A(new_new_n73_), .Y(new_new_n976_));
  AOI210     g954(.A0(new_new_n935_), .A1(i_5_), .B0(new_new_n878_), .Y(new_new_n977_));
  AOI210     g955(.A0(new_new_n977_), .A1(new_new_n976_), .B0(new_new_n660_), .Y(new_new_n978_));
  NA2        g956(.A(new_new_n258_), .B(new_new_n54_), .Y(new_new_n979_));
  AOI220     g957(.A0(new_new_n979_), .A1(new_new_n73_), .B0(new_new_n345_), .B1(new_new_n250_), .Y(new_new_n980_));
  NO2        g958(.A(new_new_n980_), .B(new_new_n231_), .Y(new_new_n981_));
  NA3        g959(.A(new_new_n93_), .B(new_new_n304_), .C(new_new_n31_), .Y(new_new_n982_));
  INV        g960(.A(new_new_n982_), .Y(new_new_n983_));
  NO3        g961(.A(new_new_n983_), .B(new_new_n981_), .C(new_new_n978_), .Y(new_new_n984_));
  OAI210     g962(.A0(new_new_n266_), .A1(new_new_n152_), .B0(new_new_n83_), .Y(new_new_n985_));
  NO2        g963(.A(new_new_n985_), .B(i_11_), .Y(new_new_n986_));
  OAI210     g964(.A0(new_new_n998_), .A1(new_new_n873_), .B0(new_new_n199_), .Y(new_new_n987_));
  NA2        g965(.A(new_new_n158_), .B(i_5_), .Y(new_new_n988_));
  NO2        g966(.A(new_new_n987_), .B(new_new_n988_), .Y(new_new_n989_));
  NO2        g967(.A(new_new_n989_), .B(new_new_n986_), .Y(new_new_n990_));
  OAI210     g968(.A0(new_new_n984_), .A1(i_4_), .B0(new_new_n990_), .Y(new_new_n991_));
  NO3        g969(.A(new_new_n991_), .B(new_new_n975_), .C(new_new_n973_), .Y(new_new_n992_));
  NA4        g970(.A(new_new_n992_), .B(new_new_n955_), .C(new_new_n903_), .D(new_new_n844_), .Y(mai4));
  INV        g971(.A(i_2_), .Y(new_new_n996_));
  INV        g972(.A(i_12_), .Y(new_new_n997_));
  INV        g973(.A(i_12_), .Y(new_new_n998_));
  INV        g974(.A(new_new_n832_), .Y(new_new_n999_));
  INV        g975(.A(new_new_n157_), .Y(new_new_n1000_));
  INV        g976(.A(i_1_), .Y(new_new_n1001_));
endmodule


