//Benchmark atmr_9sym_175_0.25

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, ori00, mai00, men00;
  ONE        o0(.Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  INV        m002(.A(i_5_), .Y(mai_mai_n13_));
  NOi21      m003(.An(i_3_), .B(i_7_), .Y(mai_mai_n14_));
  INV        m004(.A(i_0_), .Y(mai_mai_n15_));
  INV        m005(.A(i_4_), .Y(mai_mai_n16_));
  NA2        m006(.A(i_0_), .B(mai_mai_n16_), .Y(mai_mai_n17_));
  INV        m007(.A(i_7_), .Y(mai_mai_n18_));
  NA3        m008(.A(i_6_), .B(i_5_), .C(mai_mai_n18_), .Y(mai_mai_n19_));
  NO2        m009(.A(mai_mai_n19_), .B(mai_mai_n17_), .Y(mai_mai_n20_));
  NA2        m010(.A(mai_mai_n20_), .B(mai_mai_n11_), .Y(mai_mai_n21_));
  NA2        m011(.A(mai_mai_n15_), .B(i_5_), .Y(mai_mai_n22_));
  NO2        m012(.A(i_2_), .B(i_4_), .Y(mai_mai_n23_));
  INV        m013(.A(i_2_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_5_), .B(i_0_), .Y(mai_mai_n25_));
  NOi21      m015(.An(i_6_), .B(i_8_), .Y(mai_mai_n26_));
  NOi21      m016(.An(i_7_), .B(i_1_), .Y(mai_mai_n27_));
  NOi21      m017(.An(i_5_), .B(i_6_), .Y(mai_mai_n28_));
  AOI220     m018(.A0(mai_mai_n28_), .A1(mai_mai_n27_), .B0(mai_mai_n26_), .B1(mai_mai_n25_), .Y(mai_mai_n29_));
  NO3        m019(.A(mai_mai_n29_), .B(mai_mai_n24_), .C(i_4_), .Y(mai_mai_n30_));
  NOi21      m020(.An(i_0_), .B(i_4_), .Y(mai_mai_n31_));
  XO2        m021(.A(i_1_), .B(i_3_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_7_), .B(i_5_), .Y(mai_mai_n33_));
  AN3        m023(.A(mai_mai_n33_), .B(mai_mai_n32_), .C(mai_mai_n31_), .Y(mai_mai_n34_));
  INV        m024(.A(i_1_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_3_), .B(i_0_), .Y(mai_mai_n36_));
  NA2        m026(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n37_));
  NA3        m027(.A(i_6_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n38_));
  AOI210     m028(.A0(mai_mai_n38_), .A1(mai_mai_n19_), .B0(mai_mai_n37_), .Y(mai_mai_n39_));
  NO3        m029(.A(mai_mai_n39_), .B(mai_mai_n34_), .C(mai_mai_n30_), .Y(mai_mai_n40_));
  INV        m030(.A(i_8_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_4_), .B(i_0_), .Y(mai_mai_n42_));
  INV        m032(.A(mai_mai_n14_), .Y(mai_mai_n43_));
  NA2        m033(.A(i_1_), .B(mai_mai_n13_), .Y(mai_mai_n44_));
  NOi21      m034(.An(i_2_), .B(i_8_), .Y(mai_mai_n45_));
  NO2        m035(.A(mai_mai_n45_), .B(mai_mai_n31_), .Y(mai_mai_n46_));
  NO3        m036(.A(mai_mai_n46_), .B(mai_mai_n44_), .C(mai_mai_n43_), .Y(mai_mai_n47_));
  INV        m037(.A(mai_mai_n47_), .Y(mai_mai_n48_));
  NOi31      m038(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n49_));
  NA2        m039(.A(mai_mai_n49_), .B(i_0_), .Y(mai_mai_n50_));
  NOi21      m040(.An(i_4_), .B(i_3_), .Y(mai_mai_n51_));
  NOi21      m041(.An(i_1_), .B(i_4_), .Y(mai_mai_n52_));
  OAI210     m042(.A0(mai_mai_n52_), .A1(mai_mai_n51_), .B0(mai_mai_n45_), .Y(mai_mai_n53_));
  NA2        m043(.A(mai_mai_n53_), .B(mai_mai_n50_), .Y(mai_mai_n54_));
  AN2        m044(.A(i_8_), .B(i_7_), .Y(mai_mai_n55_));
  NA2        m045(.A(mai_mai_n55_), .B(mai_mai_n12_), .Y(mai_mai_n56_));
  NOi21      m046(.An(i_8_), .B(i_7_), .Y(mai_mai_n57_));
  NA3        m047(.A(mai_mai_n57_), .B(mai_mai_n51_), .C(i_6_), .Y(mai_mai_n58_));
  OAI210     m048(.A0(mai_mai_n56_), .A1(mai_mai_n44_), .B0(mai_mai_n58_), .Y(mai_mai_n59_));
  AOI220     m049(.A0(mai_mai_n59_), .A1(mai_mai_n24_), .B0(mai_mai_n54_), .B1(mai_mai_n28_), .Y(mai_mai_n60_));
  NA4        m050(.A(mai_mai_n60_), .B(mai_mai_n48_), .C(mai_mai_n40_), .D(mai_mai_n21_), .Y(mai_mai_n61_));
  NA2        m051(.A(i_8_), .B(mai_mai_n18_), .Y(mai_mai_n62_));
  AOI220     m052(.A0(mai_mai_n36_), .A1(i_1_), .B0(mai_mai_n32_), .B1(i_2_), .Y(mai_mai_n63_));
  NOi21      m053(.An(i_1_), .B(i_2_), .Y(mai_mai_n64_));
  NO2        m054(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n65_));
  NA2        m055(.A(mai_mai_n65_), .B(mai_mai_n13_), .Y(mai_mai_n66_));
  NA3        m056(.A(mai_mai_n57_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n67_));
  INV        m057(.A(mai_mai_n66_), .Y(mai_mai_n68_));
  NAi21      m058(.An(i_3_), .B(i_6_), .Y(mai_mai_n69_));
  NO3        m059(.A(mai_mai_n69_), .B(i_0_), .C(mai_mai_n41_), .Y(mai_mai_n70_));
  NA2        m060(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n71_));
  NOi21      m061(.An(i_7_), .B(i_8_), .Y(mai_mai_n72_));
  NA2        m062(.A(mai_mai_n72_), .B(mai_mai_n12_), .Y(mai_mai_n73_));
  OAI210     m063(.A0(mai_mai_n73_), .A1(mai_mai_n11_), .B0(mai_mai_n71_), .Y(mai_mai_n74_));
  OAI210     m064(.A0(mai_mai_n74_), .A1(mai_mai_n70_), .B0(mai_mai_n64_), .Y(mai_mai_n75_));
  NA3        m065(.A(mai_mai_n57_), .B(mai_mai_n24_), .C(i_3_), .Y(mai_mai_n76_));
  NA2        m066(.A(mai_mai_n35_), .B(i_6_), .Y(mai_mai_n77_));
  AOI210     m067(.A0(mai_mai_n77_), .A1(mai_mai_n17_), .B0(mai_mai_n76_), .Y(mai_mai_n78_));
  NAi21      m068(.An(i_6_), .B(i_0_), .Y(mai_mai_n79_));
  NOi21      m069(.An(i_4_), .B(i_6_), .Y(mai_mai_n80_));
  NA2        m070(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n81_));
  NOi21      m071(.An(mai_mai_n33_), .B(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m072(.A(mai_mai_n82_), .B(mai_mai_n78_), .Y(mai_mai_n83_));
  NA2        m073(.A(mai_mai_n83_), .B(mai_mai_n75_), .Y(mai_mai_n84_));
  NA2        m074(.A(mai_mai_n45_), .B(mai_mai_n14_), .Y(mai_mai_n85_));
  NOi31      m075(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n86_));
  NOi31      m076(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n87_));
  OAI210     m077(.A0(mai_mai_n87_), .A1(mai_mai_n86_), .B0(i_7_), .Y(mai_mai_n88_));
  NA3        m078(.A(mai_mai_n88_), .B(mai_mai_n85_), .C(mai_mai_n81_), .Y(mai_mai_n89_));
  NA2        m079(.A(mai_mai_n89_), .B(mai_mai_n31_), .Y(mai_mai_n90_));
  NA2        m080(.A(mai_mai_n51_), .B(mai_mai_n27_), .Y(mai_mai_n91_));
  AOI210     m081(.A0(mai_mai_n91_), .A1(mai_mai_n67_), .B0(mai_mai_n22_), .Y(mai_mai_n92_));
  NA3        m082(.A(mai_mai_n57_), .B(mai_mai_n49_), .C(i_6_), .Y(mai_mai_n93_));
  INV        m083(.A(mai_mai_n93_), .Y(mai_mai_n94_));
  NOi21      m084(.An(i_0_), .B(i_2_), .Y(mai_mai_n95_));
  NA3        m085(.A(mai_mai_n95_), .B(mai_mai_n27_), .C(mai_mai_n80_), .Y(mai_mai_n96_));
  NA3        m086(.A(mai_mai_n95_), .B(mai_mai_n51_), .C(mai_mai_n26_), .Y(mai_mai_n97_));
  NA2        m087(.A(mai_mai_n97_), .B(mai_mai_n96_), .Y(mai_mai_n98_));
  NA4        m088(.A(mai_mai_n49_), .B(i_6_), .C(mai_mai_n13_), .D(i_7_), .Y(mai_mai_n99_));
  NA4        m089(.A(mai_mai_n52_), .B(mai_mai_n28_), .C(mai_mai_n15_), .D(i_8_), .Y(mai_mai_n100_));
  NA2        m090(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  NO4        m091(.A(mai_mai_n101_), .B(mai_mai_n98_), .C(mai_mai_n94_), .D(mai_mai_n92_), .Y(mai_mai_n102_));
  NA2        m092(.A(mai_mai_n55_), .B(mai_mai_n23_), .Y(mai_mai_n103_));
  AOI210     m093(.A0(mai_mai_n103_), .A1(mai_mai_n85_), .B0(mai_mai_n77_), .Y(mai_mai_n104_));
  NO4        m094(.A(i_2_), .B(mai_mai_n16_), .C(mai_mai_n11_), .D(mai_mai_n13_), .Y(mai_mai_n105_));
  NA2        m095(.A(i_2_), .B(i_4_), .Y(mai_mai_n106_));
  AOI210     m096(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(mai_mai_n106_), .Y(mai_mai_n107_));
  NO2        m097(.A(i_8_), .B(i_7_), .Y(mai_mai_n108_));
  OA210      m098(.A0(mai_mai_n107_), .A1(mai_mai_n105_), .B0(mai_mai_n108_), .Y(mai_mai_n109_));
  NO2        m099(.A(mai_mai_n109_), .B(mai_mai_n104_), .Y(mai_mai_n110_));
  NA2        m100(.A(mai_mai_n72_), .B(mai_mai_n12_), .Y(mai_mai_n111_));
  NA3        m101(.A(i_2_), .B(i_1_), .C(mai_mai_n13_), .Y(mai_mai_n112_));
  NA2        m102(.A(mai_mai_n42_), .B(i_3_), .Y(mai_mai_n113_));
  AOI210     m103(.A0(mai_mai_n113_), .A1(mai_mai_n112_), .B0(mai_mai_n111_), .Y(mai_mai_n114_));
  NA3        m104(.A(mai_mai_n95_), .B(mai_mai_n57_), .C(mai_mai_n80_), .Y(mai_mai_n115_));
  OAI210     m105(.A0(mai_mai_n76_), .A1(mai_mai_n22_), .B0(mai_mai_n115_), .Y(mai_mai_n116_));
  NO2        m106(.A(mai_mai_n116_), .B(mai_mai_n114_), .Y(mai_mai_n117_));
  NA4        m107(.A(mai_mai_n117_), .B(mai_mai_n110_), .C(mai_mai_n102_), .D(mai_mai_n90_), .Y(mai_mai_n118_));
  OR4        m108(.A(mai_mai_n118_), .B(mai_mai_n84_), .C(mai_mai_n68_), .D(mai_mai_n61_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NA3        u013(.A(i_6_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n24_));
  NOi21      u014(.An(i_8_), .B(i_6_), .Y(men_men_n25_));
  NOi21      u015(.An(i_1_), .B(i_8_), .Y(men_men_n26_));
  AOI220     u016(.A0(men_men_n26_), .A1(i_2_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n22_), .Y(men_men_n28_));
  AOI210     u018(.A0(men_men_n28_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n29_));
  NA2        u019(.A(i_0_), .B(men_men_n14_), .Y(men_men_n30_));
  NA2        u020(.A(men_men_n17_), .B(i_5_), .Y(men_men_n31_));
  NO2        u021(.A(i_2_), .B(i_4_), .Y(men_men_n32_));
  NA3        u022(.A(men_men_n32_), .B(i_6_), .C(i_8_), .Y(men_men_n33_));
  AOI210     u023(.A0(men_men_n31_), .A1(men_men_n30_), .B0(men_men_n33_), .Y(men_men_n34_));
  INV        u024(.A(i_2_), .Y(men_men_n35_));
  NOi21      u025(.An(i_5_), .B(i_0_), .Y(men_men_n36_));
  NOi21      u026(.An(i_6_), .B(i_8_), .Y(men_men_n37_));
  NOi21      u027(.An(i_0_), .B(i_4_), .Y(men_men_n38_));
  NOi21      u028(.An(i_7_), .B(i_5_), .Y(men_men_n39_));
  INV        u029(.A(i_1_), .Y(men_men_n40_));
  NOi21      u030(.An(i_3_), .B(i_0_), .Y(men_men_n41_));
  INV        u031(.A(men_men_n34_), .Y(men_men_n42_));
  INV        u032(.A(i_8_), .Y(men_men_n43_));
  NA2        u033(.A(i_1_), .B(men_men_n11_), .Y(men_men_n44_));
  NO4        u034(.A(men_men_n44_), .B(men_men_n30_), .C(i_2_), .D(men_men_n43_), .Y(men_men_n45_));
  NOi21      u035(.An(i_4_), .B(i_0_), .Y(men_men_n46_));
  AOI210     u036(.A0(men_men_n46_), .A1(men_men_n25_), .B0(men_men_n15_), .Y(men_men_n47_));
  NA2        u037(.A(i_1_), .B(men_men_n14_), .Y(men_men_n48_));
  NOi21      u038(.An(i_2_), .B(i_8_), .Y(men_men_n49_));
  NO3        u039(.A(men_men_n49_), .B(men_men_n46_), .C(men_men_n38_), .Y(men_men_n50_));
  NO3        u040(.A(men_men_n50_), .B(men_men_n48_), .C(men_men_n47_), .Y(men_men_n51_));
  NO2        u041(.A(men_men_n51_), .B(men_men_n45_), .Y(men_men_n52_));
  NOi21      u042(.An(i_4_), .B(i_3_), .Y(men_men_n53_));
  NOi21      u043(.An(i_1_), .B(i_4_), .Y(men_men_n54_));
  AN2        u044(.A(i_8_), .B(i_7_), .Y(men_men_n55_));
  NOi21      u045(.An(i_8_), .B(i_7_), .Y(men_men_n56_));
  NA3        u046(.A(men_men_n52_), .B(men_men_n42_), .C(men_men_n29_), .Y(men_men_n57_));
  NA2        u047(.A(i_8_), .B(i_7_), .Y(men_men_n58_));
  NO3        u048(.A(men_men_n58_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n59_));
  NOi21      u049(.An(i_1_), .B(i_2_), .Y(men_men_n60_));
  NA3        u050(.A(men_men_n60_), .B(men_men_n46_), .C(i_6_), .Y(men_men_n61_));
  INV        u051(.A(men_men_n61_), .Y(men_men_n62_));
  OAI210     u052(.A0(men_men_n62_), .A1(men_men_n59_), .B0(men_men_n14_), .Y(men_men_n63_));
  NA3        u053(.A(men_men_n56_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n64_));
  NA3        u054(.A(men_men_n26_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n65_));
  NA2        u055(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NOi32      u056(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n67_));
  NA2        u057(.A(men_men_n67_), .B(i_3_), .Y(men_men_n68_));
  NA3        u058(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n69_));
  NA2        u059(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NO2        u060(.A(i_0_), .B(i_4_), .Y(men_men_n71_));
  AOI220     u061(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n66_), .B1(men_men_n53_), .Y(men_men_n72_));
  NA2        u062(.A(men_men_n72_), .B(men_men_n63_), .Y(men_men_n73_));
  NOi21      u063(.An(i_7_), .B(i_8_), .Y(men_men_n74_));
  NOi31      u064(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n75_));
  AOI210     u065(.A0(men_men_n74_), .A1(men_men_n12_), .B0(men_men_n75_), .Y(men_men_n76_));
  NO2        u066(.A(men_men_n76_), .B(men_men_n11_), .Y(men_men_n77_));
  NA2        u067(.A(men_men_n77_), .B(men_men_n60_), .Y(men_men_n78_));
  NA3        u068(.A(men_men_n25_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n79_));
  AOI210     u069(.A0(men_men_n22_), .A1(men_men_n44_), .B0(men_men_n79_), .Y(men_men_n80_));
  AOI220     u070(.A0(men_men_n41_), .A1(men_men_n40_), .B0(men_men_n18_), .B1(men_men_n35_), .Y(men_men_n81_));
  NA3        u071(.A(men_men_n21_), .B(i_5_), .C(i_7_), .Y(men_men_n82_));
  OAI210     u072(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n83_));
  NA3        u073(.A(men_men_n58_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n84_));
  OAI220     u074(.A0(men_men_n84_), .A1(men_men_n83_), .B0(men_men_n82_), .B1(men_men_n81_), .Y(men_men_n85_));
  NO2        u075(.A(men_men_n85_), .B(men_men_n80_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n40_), .B(i_6_), .Y(men_men_n87_));
  NOi21      u077(.An(i_2_), .B(i_1_), .Y(men_men_n88_));
  AN3        u078(.A(men_men_n74_), .B(men_men_n88_), .C(men_men_n46_), .Y(men_men_n89_));
  NAi21      u079(.An(i_6_), .B(i_0_), .Y(men_men_n90_));
  NA3        u080(.A(men_men_n54_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n91_));
  NOi21      u081(.An(i_4_), .B(i_6_), .Y(men_men_n92_));
  NOi21      u082(.An(i_5_), .B(i_3_), .Y(men_men_n93_));
  NA3        u083(.A(men_men_n93_), .B(men_men_n60_), .C(men_men_n92_), .Y(men_men_n94_));
  OAI210     u084(.A0(men_men_n91_), .A1(men_men_n90_), .B0(men_men_n94_), .Y(men_men_n95_));
  NO2        u085(.A(men_men_n95_), .B(men_men_n89_), .Y(men_men_n96_));
  NOi21      u086(.An(i_6_), .B(i_1_), .Y(men_men_n97_));
  AOI220     u087(.A0(men_men_n97_), .A1(i_7_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n98_));
  NOi31      u088(.An(men_men_n46_), .B(men_men_n98_), .C(i_2_), .Y(men_men_n99_));
  NA2        u089(.A(men_men_n56_), .B(men_men_n12_), .Y(men_men_n100_));
  NA2        u090(.A(men_men_n37_), .B(men_men_n14_), .Y(men_men_n101_));
  NOi21      u091(.An(i_3_), .B(i_1_), .Y(men_men_n102_));
  NA2        u092(.A(men_men_n102_), .B(i_4_), .Y(men_men_n103_));
  AOI210     u093(.A0(men_men_n101_), .A1(men_men_n100_), .B0(men_men_n103_), .Y(men_men_n104_));
  AOI220     u094(.A0(men_men_n74_), .A1(men_men_n14_), .B0(men_men_n92_), .B1(men_men_n23_), .Y(men_men_n105_));
  NOi31      u095(.An(men_men_n41_), .B(men_men_n105_), .C(men_men_n35_), .Y(men_men_n106_));
  NO3        u096(.A(men_men_n106_), .B(men_men_n104_), .C(men_men_n99_), .Y(men_men_n107_));
  NA4        u097(.A(men_men_n107_), .B(men_men_n96_), .C(men_men_n86_), .D(men_men_n78_), .Y(men_men_n108_));
  NOi31      u098(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n109_));
  NA3        u099(.A(men_men_n37_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n110_));
  INV        u100(.A(men_men_n110_), .Y(men_men_n111_));
  NA2        u101(.A(men_men_n111_), .B(men_men_n38_), .Y(men_men_n112_));
  NA4        u102(.A(men_men_n55_), .B(men_men_n88_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n113_));
  NAi31      u103(.An(men_men_n90_), .B(men_men_n74_), .C(men_men_n88_), .Y(men_men_n114_));
  NA2        u104(.A(men_men_n114_), .B(men_men_n113_), .Y(men_men_n115_));
  NA3        u105(.A(men_men_n46_), .B(men_men_n39_), .C(men_men_n18_), .Y(men_men_n116_));
  NOi32      u106(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n117_));
  NA2        u107(.A(men_men_n117_), .B(men_men_n109_), .Y(men_men_n118_));
  NA2        u108(.A(men_men_n118_), .B(men_men_n116_), .Y(men_men_n119_));
  NA4        u109(.A(men_men_n54_), .B(men_men_n41_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n120_));
  INV        u110(.A(men_men_n120_), .Y(men_men_n121_));
  NO3        u111(.A(men_men_n121_), .B(men_men_n119_), .C(men_men_n115_), .Y(men_men_n122_));
  NOi21      u112(.An(i_5_), .B(i_2_), .Y(men_men_n123_));
  NA2        u113(.A(men_men_n123_), .B(men_men_n74_), .Y(men_men_n124_));
  NO2        u114(.A(men_men_n124_), .B(men_men_n87_), .Y(men_men_n125_));
  NA4        u115(.A(men_men_n102_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n126_));
  NO2        u116(.A(men_men_n126_), .B(i_4_), .Y(men_men_n127_));
  NO2        u117(.A(men_men_n127_), .B(men_men_n125_), .Y(men_men_n128_));
  NA4        u118(.A(men_men_n93_), .B(men_men_n55_), .C(men_men_n40_), .D(men_men_n21_), .Y(men_men_n129_));
  NA3        u119(.A(men_men_n75_), .B(men_men_n102_), .C(i_0_), .Y(men_men_n130_));
  NA3        u120(.A(men_men_n49_), .B(men_men_n36_), .C(men_men_n15_), .Y(men_men_n131_));
  NOi31      u121(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n132_));
  OAI210     u122(.A0(men_men_n117_), .A1(men_men_n67_), .B0(men_men_n132_), .Y(men_men_n133_));
  NA4        u123(.A(men_men_n133_), .B(men_men_n131_), .C(men_men_n130_), .D(men_men_n129_), .Y(men_men_n134_));
  INV        u124(.A(men_men_n134_), .Y(men_men_n135_));
  NA4        u125(.A(men_men_n135_), .B(men_men_n128_), .C(men_men_n122_), .D(men_men_n112_), .Y(men_men_n136_));
  OR4        u126(.A(men_men_n136_), .B(men_men_n108_), .C(men_men_n73_), .D(men_men_n57_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule