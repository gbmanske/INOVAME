// Benchmark "top" written by ABC on Fri Jun 21 17:49:24 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1080_, new_new_n1081_, new_new_n1082_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g0028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g0029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g0032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g0062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g0063(.A(i_6_), .Y(new_new_n86_));
  NO2        g0064(.A(i_2_), .B(i_7_), .Y(new_new_n87_));
  OAI210     g0065(.A0(new_new_n85_), .A1(new_new_n82_), .B0(i_2_), .Y(new_new_n88_));
  NAi21      g0066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g0067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g0068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n63_), .Y(new_new_n91_));
  NA2        g0069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g0070(.A(new_new_n92_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g0071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n88_), .B0(new_new_n80_), .Y(new_new_n95_));
  AN3        g0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g0074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g0075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g0076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g0077(.A0(new_new_n99_), .A1(new_new_n62_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g0078(.A(i_7_), .Y(new_new_n101_));
  NA2        g0079(.A(new_new_n46_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g0080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g0081(.A(new_new_n103_), .B(new_new_n86_), .Y(new_new_n104_));
  NA2        g0082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g0083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g0084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g0085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  AN2        g0086(.A(i_2_), .B(i_10_), .Y(new_new_n109_));
  NO2        g0087(.A(new_new_n109_), .B(i_7_), .Y(new_new_n110_));
  OR2        g0088(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n111_));
  NO2        g0089(.A(i_8_), .B(new_new_n101_), .Y(new_new_n112_));
  NO3        g0090(.A(new_new_n112_), .B(new_new_n111_), .C(new_new_n110_), .Y(new_new_n113_));
  NA2        g0091(.A(i_12_), .B(i_7_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n115_));
  NA2        g0093(.A(new_new_n115_), .B(i_0_), .Y(new_new_n116_));
  NA2        g0094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  OAI210     g0095(.A0(new_new_n116_), .A1(new_new_n114_), .B0(new_new_n117_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n118_), .B(new_new_n113_), .Y(new_new_n119_));
  NA3        g0097(.A(new_new_n119_), .B(new_new_n107_), .C(new_new_n100_), .Y(new_new_n120_));
  NOi21      g0098(.An(i_1_), .B(i_5_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n121_), .B(i_11_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g0101(.A(i_7_), .B(new_new_n25_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(new_new_n123_), .Y(new_new_n125_));
  NO2        g0103(.A(new_new_n125_), .B(new_new_n46_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n127_));
  NAi21      g0105(.An(i_3_), .B(i_8_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n62_), .Y(new_new_n129_));
  NOi31      g0107(.An(new_new_n129_), .B(new_new_n127_), .C(new_new_n126_), .Y(new_new_n130_));
  NO2        g0108(.A(i_1_), .B(new_new_n86_), .Y(new_new_n131_));
  NO2        g0109(.A(i_6_), .B(i_5_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(i_3_), .Y(new_new_n133_));
  AO210      g0111(.A0(new_new_n133_), .A1(new_new_n47_), .B0(new_new_n131_), .Y(new_new_n134_));
  OAI220     g0112(.A0(new_new_n134_), .A1(new_new_n108_), .B0(new_new_n130_), .B1(new_new_n122_), .Y(new_new_n135_));
  NO3        g0113(.A(new_new_n135_), .B(new_new_n120_), .C(new_new_n95_), .Y(new_new_n136_));
  NA3        g0114(.A(new_new_n136_), .B(new_new_n79_), .C(new_new_n56_), .Y(men2));
  NO2        g0115(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n138_));
  NA2        g0116(.A(i_6_), .B(new_new_n25_), .Y(new_new_n139_));
  NA2        g0117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g0118(.A(new_new_n140_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(men0));
  AN2        g0119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g0121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g0122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g0123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g0124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g0125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NO2        g0126(.A(new_new_n148_), .B(i_4_), .Y(new_new_n149_));
  NA3        g0127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  OR2        g0128(.A(new_new_n150_), .B(new_new_n25_), .Y(new_new_n151_));
  AN2        g0129(.A(new_new_n144_), .B(new_new_n83_), .Y(new_new_n152_));
  NO2        g0130(.A(new_new_n152_), .B(new_new_n27_), .Y(new_new_n153_));
  NA2        g0131(.A(i_1_), .B(i_5_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n73_), .B(new_new_n46_), .Y(new_new_n155_));
  NA2        g0133(.A(new_new_n155_), .B(new_new_n36_), .Y(new_new_n156_));
  NO3        g0134(.A(new_new_n156_), .B(new_new_n154_), .C(new_new_n153_), .Y(new_new_n157_));
  OR2        g0135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n159_));
  NAi32      g0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n160_));
  NAi21      g0138(.An(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NOi21      g0139(.An(i_4_), .B(i_10_), .Y(new_new_n162_));
  NA2        g0140(.A(new_new_n162_), .B(new_new_n40_), .Y(new_new_n163_));
  NO2        g0141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  NO3        g0142(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OAI210     g0144(.A0(new_new_n166_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n167_));
  NO2        g0145(.A(new_new_n167_), .B(new_new_n157_), .Y(new_new_n168_));
  AOI210     g0146(.A0(new_new_n168_), .A1(new_new_n151_), .B0(new_new_n143_), .Y(new_new_n169_));
  NA3        g0147(.A(new_new_n73_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n170_));
  NA2        g0148(.A(i_3_), .B(new_new_n48_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_4_), .B(i_9_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_11_), .B(i_13_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n173_), .B(new_new_n172_), .Y(new_new_n174_));
  OR2        g0152(.A(new_new_n174_), .B(new_new_n171_), .Y(new_new_n175_));
  NO2        g0153(.A(i_4_), .B(i_5_), .Y(new_new_n176_));
  NAi21      g0154(.An(i_12_), .B(i_11_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n177_), .B(i_13_), .Y(new_new_n178_));
  NA3        g0156(.A(new_new_n178_), .B(new_new_n176_), .C(new_new_n83_), .Y(new_new_n179_));
  AOI210     g0157(.A0(new_new_n179_), .A1(new_new_n175_), .B0(new_new_n170_), .Y(new_new_n180_));
  NO2        g0158(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n181_), .B(new_new_n46_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n36_), .B(i_5_), .Y(new_new_n183_));
  NAi31      g0161(.An(new_new_n183_), .B(new_new_n152_), .C(i_11_), .Y(new_new_n184_));
  NA2        g0162(.A(i_3_), .B(i_5_), .Y(new_new_n185_));
  OR2        g0163(.A(new_new_n185_), .B(new_new_n174_), .Y(new_new_n186_));
  AOI210     g0164(.A0(new_new_n186_), .A1(new_new_n184_), .B0(new_new_n182_), .Y(new_new_n187_));
  NO2        g0165(.A(new_new_n73_), .B(i_5_), .Y(new_new_n188_));
  NO2        g0166(.A(i_13_), .B(i_10_), .Y(new_new_n189_));
  NA3        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n44_), .Y(new_new_n190_));
  NO2        g0168(.A(i_2_), .B(i_1_), .Y(new_new_n191_));
  NA2        g0169(.A(new_new_n191_), .B(i_3_), .Y(new_new_n192_));
  NAi21      g0170(.An(i_4_), .B(i_12_), .Y(new_new_n193_));
  NO4        g0171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n190_), .D(new_new_n25_), .Y(new_new_n194_));
  NO3        g0172(.A(new_new_n194_), .B(new_new_n187_), .C(new_new_n180_), .Y(new_new_n195_));
  INV        g0173(.A(i_8_), .Y(new_new_n196_));
  NO2        g0174(.A(new_new_n196_), .B(i_7_), .Y(new_new_n197_));
  NA2        g0175(.A(new_new_n197_), .B(i_6_), .Y(new_new_n198_));
  NO3        g0176(.A(i_3_), .B(new_new_n86_), .C(new_new_n48_), .Y(new_new_n199_));
  NA2        g0177(.A(new_new_n199_), .B(new_new_n112_), .Y(new_new_n200_));
  NO3        g0178(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n201_));
  NA3        g0179(.A(new_new_n201_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n202_));
  NO3        g0180(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n203_));
  OAI210     g0181(.A0(new_new_n96_), .A1(i_12_), .B0(new_new_n203_), .Y(new_new_n204_));
  AOI210     g0182(.A0(new_new_n204_), .A1(new_new_n202_), .B0(new_new_n200_), .Y(new_new_n205_));
  NO2        g0183(.A(i_3_), .B(i_8_), .Y(new_new_n206_));
  NO3        g0184(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n207_));
  NA3        g0185(.A(new_new_n207_), .B(new_new_n206_), .C(new_new_n40_), .Y(new_new_n208_));
  NO2        g0186(.A(new_new_n103_), .B(new_new_n58_), .Y(new_new_n209_));
  INV        g0187(.A(new_new_n209_), .Y(new_new_n210_));
  NO2        g0188(.A(i_13_), .B(i_9_), .Y(new_new_n211_));
  NA3        g0189(.A(new_new_n211_), .B(i_6_), .C(new_new_n196_), .Y(new_new_n212_));
  NAi21      g0190(.An(i_12_), .B(i_3_), .Y(new_new_n213_));
  NO2        g0191(.A(new_new_n44_), .B(i_5_), .Y(new_new_n214_));
  NO3        g0192(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n215_));
  NA3        g0193(.A(new_new_n215_), .B(new_new_n214_), .C(i_10_), .Y(new_new_n216_));
  OAI220     g0194(.A0(new_new_n216_), .A1(new_new_n212_), .B0(new_new_n210_), .B1(new_new_n208_), .Y(new_new_n217_));
  AOI210     g0195(.A0(new_new_n217_), .A1(i_7_), .B0(new_new_n205_), .Y(new_new_n218_));
  OAI220     g0196(.A0(new_new_n218_), .A1(i_4_), .B0(new_new_n198_), .B1(new_new_n195_), .Y(new_new_n219_));
  NAi21      g0197(.An(i_12_), .B(i_7_), .Y(new_new_n220_));
  NA3        g0198(.A(i_13_), .B(new_new_n196_), .C(i_10_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n222_));
  NA2        g0200(.A(i_0_), .B(i_5_), .Y(new_new_n223_));
  NA2        g0201(.A(new_new_n223_), .B(new_new_n104_), .Y(new_new_n224_));
  OAI220     g0202(.A0(new_new_n224_), .A1(new_new_n192_), .B0(new_new_n182_), .B1(new_new_n133_), .Y(new_new_n225_));
  NAi31      g0203(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n226_));
  NO2        g0204(.A(new_new_n36_), .B(i_13_), .Y(new_new_n227_));
  NO2        g0205(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n229_));
  NA3        g0207(.A(new_new_n229_), .B(new_new_n228_), .C(new_new_n227_), .Y(new_new_n230_));
  INV        g0208(.A(i_13_), .Y(new_new_n231_));
  NO2        g0209(.A(i_12_), .B(new_new_n231_), .Y(new_new_n232_));
  NA3        g0210(.A(new_new_n232_), .B(new_new_n201_), .C(new_new_n199_), .Y(new_new_n233_));
  OAI210     g0211(.A0(new_new_n230_), .A1(new_new_n226_), .B0(new_new_n233_), .Y(new_new_n234_));
  AOI220     g0212(.A0(new_new_n234_), .A1(new_new_n142_), .B0(new_new_n225_), .B1(new_new_n222_), .Y(new_new_n235_));
  NO2        g0213(.A(i_12_), .B(new_new_n37_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n185_), .B(i_4_), .Y(new_new_n237_));
  NA2        g0215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  OR2        g0216(.A(i_8_), .B(i_7_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n239_), .B(new_new_n86_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n53_), .B(i_1_), .Y(new_new_n241_));
  NA2        g0219(.A(new_new_n241_), .B(new_new_n240_), .Y(new_new_n242_));
  INV        g0220(.A(i_12_), .Y(new_new_n243_));
  NO2        g0221(.A(new_new_n44_), .B(new_new_n243_), .Y(new_new_n244_));
  NO3        g0222(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n245_));
  NA2        g0223(.A(i_2_), .B(i_1_), .Y(new_new_n246_));
  NO2        g0224(.A(new_new_n242_), .B(new_new_n238_), .Y(new_new_n247_));
  NO3        g0225(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n248_));
  NAi21      g0226(.An(i_4_), .B(i_3_), .Y(new_new_n249_));
  NO2        g0227(.A(i_0_), .B(i_6_), .Y(new_new_n250_));
  NOi41      g0228(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n251_));
  NA2        g0229(.A(new_new_n251_), .B(new_new_n250_), .Y(new_new_n252_));
  NO2        g0230(.A(new_new_n246_), .B(new_new_n185_), .Y(new_new_n253_));
  NAi21      g0231(.An(new_new_n252_), .B(new_new_n253_), .Y(new_new_n254_));
  INV        g0232(.A(new_new_n254_), .Y(new_new_n255_));
  AOI220     g0233(.A0(new_new_n255_), .A1(new_new_n40_), .B0(new_new_n247_), .B1(new_new_n211_), .Y(new_new_n256_));
  NO2        g0234(.A(i_11_), .B(new_new_n231_), .Y(new_new_n257_));
  NOi21      g0235(.An(i_1_), .B(i_6_), .Y(new_new_n258_));
  NAi21      g0236(.An(i_3_), .B(i_7_), .Y(new_new_n259_));
  NA2        g0237(.A(new_new_n243_), .B(i_9_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n261_));
  NO2        g0239(.A(i_12_), .B(i_3_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n73_), .B(i_5_), .Y(new_new_n263_));
  NA2        g0241(.A(i_3_), .B(i_9_), .Y(new_new_n264_));
  NAi21      g0242(.An(i_7_), .B(i_10_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n266_));
  NA3        g0244(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n267_));
  INV        g0245(.A(new_new_n143_), .Y(new_new_n268_));
  NA2        g0246(.A(new_new_n243_), .B(i_13_), .Y(new_new_n269_));
  NO2        g0247(.A(new_new_n269_), .B(new_new_n75_), .Y(new_new_n270_));
  NA2        g0248(.A(new_new_n270_), .B(new_new_n268_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n239_), .B(new_new_n37_), .Y(new_new_n272_));
  NA2        g0250(.A(i_12_), .B(i_6_), .Y(new_new_n273_));
  OR2        g0251(.A(i_13_), .B(i_9_), .Y(new_new_n274_));
  NO3        g0252(.A(new_new_n274_), .B(new_new_n273_), .C(new_new_n48_), .Y(new_new_n275_));
  NO2        g0253(.A(new_new_n249_), .B(i_2_), .Y(new_new_n276_));
  NA3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n44_), .Y(new_new_n277_));
  NA2        g0255(.A(new_new_n257_), .B(i_9_), .Y(new_new_n278_));
  NA2        g0256(.A(new_new_n263_), .B(new_new_n64_), .Y(new_new_n279_));
  OAI210     g0257(.A0(new_new_n279_), .A1(new_new_n278_), .B0(new_new_n277_), .Y(new_new_n280_));
  NA2        g0258(.A(new_new_n155_), .B(new_new_n63_), .Y(new_new_n281_));
  NO3        g0259(.A(i_11_), .B(new_new_n231_), .C(new_new_n25_), .Y(new_new_n282_));
  NO2        g0260(.A(new_new_n259_), .B(i_8_), .Y(new_new_n283_));
  NO2        g0261(.A(i_6_), .B(new_new_n48_), .Y(new_new_n284_));
  NA3        g0262(.A(new_new_n284_), .B(new_new_n283_), .C(new_new_n282_), .Y(new_new_n285_));
  NO3        g0263(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n286_));
  NA3        g0264(.A(new_new_n286_), .B(new_new_n272_), .C(new_new_n232_), .Y(new_new_n287_));
  AOI210     g0265(.A0(new_new_n287_), .A1(new_new_n285_), .B0(new_new_n281_), .Y(new_new_n288_));
  AOI210     g0266(.A0(new_new_n280_), .A1(new_new_n272_), .B0(new_new_n288_), .Y(new_new_n289_));
  NA4        g0267(.A(new_new_n289_), .B(new_new_n271_), .C(new_new_n256_), .D(new_new_n235_), .Y(new_new_n290_));
  NO3        g0268(.A(i_12_), .B(new_new_n231_), .C(new_new_n37_), .Y(new_new_n291_));
  INV        g0269(.A(new_new_n291_), .Y(new_new_n292_));
  NA2        g0270(.A(i_8_), .B(new_new_n101_), .Y(new_new_n293_));
  NO3        g0271(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n294_));
  AOI220     g0272(.A0(new_new_n294_), .A1(new_new_n199_), .B0(new_new_n164_), .B1(new_new_n241_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n295_), .B(new_new_n293_), .Y(new_new_n296_));
  NO3        g0274(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n246_), .B(i_0_), .Y(new_new_n298_));
  AOI220     g0276(.A0(new_new_n298_), .A1(new_new_n197_), .B0(new_new_n297_), .B1(new_new_n142_), .Y(new_new_n299_));
  NA2        g0277(.A(new_new_n284_), .B(new_new_n26_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n300_), .B(new_new_n299_), .Y(new_new_n301_));
  NA2        g0279(.A(i_0_), .B(i_1_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n302_), .B(i_2_), .Y(new_new_n303_));
  NO2        g0281(.A(new_new_n59_), .B(i_6_), .Y(new_new_n304_));
  NA3        g0282(.A(new_new_n304_), .B(new_new_n303_), .C(new_new_n164_), .Y(new_new_n305_));
  OAI210     g0283(.A0(new_new_n166_), .A1(new_new_n143_), .B0(new_new_n305_), .Y(new_new_n306_));
  NO3        g0284(.A(new_new_n306_), .B(new_new_n301_), .C(new_new_n296_), .Y(new_new_n307_));
  NO2        g0285(.A(i_3_), .B(i_10_), .Y(new_new_n308_));
  NA3        g0286(.A(new_new_n308_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n309_));
  NO2        g0287(.A(i_2_), .B(new_new_n101_), .Y(new_new_n310_));
  NA2        g0288(.A(i_1_), .B(new_new_n36_), .Y(new_new_n311_));
  NO2        g0289(.A(new_new_n311_), .B(i_8_), .Y(new_new_n312_));
  NA2        g0290(.A(new_new_n312_), .B(new_new_n310_), .Y(new_new_n313_));
  AN2        g0291(.A(i_3_), .B(i_10_), .Y(new_new_n314_));
  NA4        g0292(.A(new_new_n314_), .B(new_new_n201_), .C(new_new_n178_), .D(new_new_n176_), .Y(new_new_n315_));
  NO2        g0293(.A(i_5_), .B(new_new_n37_), .Y(new_new_n316_));
  NO2        g0294(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n317_));
  OR2        g0295(.A(new_new_n313_), .B(new_new_n309_), .Y(new_new_n318_));
  OAI220     g0296(.A0(new_new_n318_), .A1(i_6_), .B0(new_new_n307_), .B1(new_new_n292_), .Y(new_new_n319_));
  NO4        g0297(.A(new_new_n319_), .B(new_new_n290_), .C(new_new_n219_), .D(new_new_n169_), .Y(new_new_n320_));
  NO3        g0298(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n321_));
  NO2        g0299(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n322_));
  NA2        g0300(.A(new_new_n298_), .B(new_new_n322_), .Y(new_new_n323_));
  NO3        g0301(.A(i_6_), .B(new_new_n196_), .C(i_7_), .Y(new_new_n324_));
  NA2        g0302(.A(new_new_n324_), .B(new_new_n201_), .Y(new_new_n325_));
  AOI210     g0303(.A0(new_new_n325_), .A1(new_new_n323_), .B0(new_new_n171_), .Y(new_new_n326_));
  NO2        g0304(.A(i_2_), .B(i_3_), .Y(new_new_n327_));
  OR2        g0305(.A(i_0_), .B(i_5_), .Y(new_new_n328_));
  NA2        g0306(.A(new_new_n223_), .B(new_new_n328_), .Y(new_new_n329_));
  NA4        g0307(.A(new_new_n329_), .B(new_new_n240_), .C(new_new_n327_), .D(i_1_), .Y(new_new_n330_));
  NA3        g0308(.A(new_new_n298_), .B(new_new_n164_), .C(new_new_n112_), .Y(new_new_n331_));
  NAi21      g0309(.An(i_8_), .B(i_7_), .Y(new_new_n332_));
  NO2        g0310(.A(new_new_n332_), .B(i_6_), .Y(new_new_n333_));
  NO2        g0311(.A(new_new_n158_), .B(new_new_n46_), .Y(new_new_n334_));
  NA3        g0312(.A(new_new_n334_), .B(new_new_n333_), .C(new_new_n164_), .Y(new_new_n335_));
  NA3        g0313(.A(new_new_n335_), .B(new_new_n331_), .C(new_new_n330_), .Y(new_new_n336_));
  OAI210     g0314(.A0(new_new_n336_), .A1(new_new_n326_), .B0(i_4_), .Y(new_new_n337_));
  NO2        g0315(.A(i_12_), .B(i_10_), .Y(new_new_n338_));
  NOi21      g0316(.An(i_5_), .B(i_0_), .Y(new_new_n339_));
  NO3        g0317(.A(new_new_n311_), .B(new_new_n339_), .C(new_new_n128_), .Y(new_new_n340_));
  NA4        g0318(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n341_));
  NA2        g0319(.A(new_new_n340_), .B(new_new_n338_), .Y(new_new_n342_));
  NO2        g0320(.A(i_6_), .B(i_8_), .Y(new_new_n343_));
  NOi21      g0321(.An(i_0_), .B(i_2_), .Y(new_new_n344_));
  AN2        g0322(.A(new_new_n344_), .B(new_new_n343_), .Y(new_new_n345_));
  NO2        g0323(.A(i_1_), .B(i_7_), .Y(new_new_n346_));
  AO220      g0324(.A0(new_new_n346_), .A1(new_new_n345_), .B0(new_new_n333_), .B1(new_new_n241_), .Y(new_new_n347_));
  NA3        g0325(.A(new_new_n347_), .B(i_4_), .C(i_5_), .Y(new_new_n348_));
  NA3        g0326(.A(new_new_n348_), .B(new_new_n342_), .C(new_new_n337_), .Y(new_new_n349_));
  NO3        g0327(.A(new_new_n239_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n350_));
  NO3        g0328(.A(new_new_n332_), .B(i_2_), .C(i_1_), .Y(new_new_n351_));
  OAI210     g0329(.A0(new_new_n351_), .A1(new_new_n350_), .B0(i_6_), .Y(new_new_n352_));
  NA2        g0330(.A(new_new_n258_), .B(new_new_n310_), .Y(new_new_n353_));
  AOI210     g0331(.A0(new_new_n353_), .A1(new_new_n352_), .B0(new_new_n329_), .Y(new_new_n354_));
  NOi21      g0332(.An(new_new_n154_), .B(new_new_n104_), .Y(new_new_n355_));
  NO2        g0333(.A(new_new_n355_), .B(new_new_n124_), .Y(new_new_n356_));
  OAI210     g0334(.A0(new_new_n356_), .A1(new_new_n354_), .B0(i_3_), .Y(new_new_n357_));
  INV        g0335(.A(new_new_n84_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n302_), .B(new_new_n81_), .Y(new_new_n359_));
  NA2        g0337(.A(new_new_n359_), .B(new_new_n132_), .Y(new_new_n360_));
  NO2        g0338(.A(new_new_n92_), .B(new_new_n196_), .Y(new_new_n361_));
  NA2        g0339(.A(new_new_n361_), .B(new_new_n63_), .Y(new_new_n362_));
  AOI210     g0340(.A0(new_new_n362_), .A1(new_new_n360_), .B0(new_new_n358_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n196_), .B(i_9_), .Y(new_new_n364_));
  NO2        g0342(.A(new_new_n363_), .B(new_new_n301_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n365_), .A1(new_new_n357_), .B0(new_new_n163_), .Y(new_new_n366_));
  AOI210     g0344(.A0(new_new_n349_), .A1(new_new_n321_), .B0(new_new_n366_), .Y(new_new_n367_));
  NOi32      g0345(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n368_));
  INV        g0346(.A(new_new_n368_), .Y(new_new_n369_));
  NAi21      g0347(.An(i_0_), .B(i_6_), .Y(new_new_n370_));
  NAi21      g0348(.An(i_1_), .B(i_5_), .Y(new_new_n371_));
  NA2        g0349(.A(new_new_n371_), .B(new_new_n370_), .Y(new_new_n372_));
  NA2        g0350(.A(new_new_n372_), .B(new_new_n25_), .Y(new_new_n373_));
  OAI210     g0351(.A0(new_new_n373_), .A1(new_new_n160_), .B0(new_new_n252_), .Y(new_new_n374_));
  NAi41      g0352(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n375_));
  AOI210     g0353(.A0(new_new_n375_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n376_));
  NOi32      g0354(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n377_));
  NO2        g0355(.A(i_1_), .B(new_new_n101_), .Y(new_new_n378_));
  NAi21      g0356(.An(i_3_), .B(i_4_), .Y(new_new_n379_));
  NO2        g0357(.A(new_new_n379_), .B(i_9_), .Y(new_new_n380_));
  AN2        g0358(.A(i_6_), .B(i_7_), .Y(new_new_n381_));
  OAI210     g0359(.A0(new_new_n381_), .A1(new_new_n378_), .B0(new_new_n380_), .Y(new_new_n382_));
  NA2        g0360(.A(i_2_), .B(i_7_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n379_), .B(i_10_), .Y(new_new_n384_));
  NA3        g0362(.A(new_new_n384_), .B(new_new_n383_), .C(new_new_n250_), .Y(new_new_n385_));
  AOI210     g0363(.A0(new_new_n385_), .A1(new_new_n382_), .B0(new_new_n188_), .Y(new_new_n386_));
  AOI210     g0364(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n387_));
  OAI210     g0365(.A0(new_new_n387_), .A1(new_new_n191_), .B0(new_new_n384_), .Y(new_new_n388_));
  AOI220     g0366(.A0(new_new_n384_), .A1(new_new_n346_), .B0(new_new_n245_), .B1(new_new_n191_), .Y(new_new_n389_));
  AOI210     g0367(.A0(new_new_n389_), .A1(new_new_n388_), .B0(i_5_), .Y(new_new_n390_));
  NO4        g0368(.A(new_new_n390_), .B(new_new_n386_), .C(new_new_n376_), .D(new_new_n374_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(new_new_n369_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n393_));
  AN2        g0371(.A(i_12_), .B(i_5_), .Y(new_new_n394_));
  NO2        g0372(.A(i_4_), .B(new_new_n26_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n395_), .B(new_new_n394_), .Y(new_new_n396_));
  NO2        g0374(.A(i_11_), .B(i_6_), .Y(new_new_n397_));
  NA3        g0375(.A(new_new_n397_), .B(new_new_n334_), .C(new_new_n231_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n398_), .B(new_new_n396_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n249_), .B(i_5_), .Y(new_new_n400_));
  NO2        g0378(.A(i_5_), .B(i_10_), .Y(new_new_n401_));
  NA2        g0379(.A(new_new_n400_), .B(new_new_n201_), .Y(new_new_n402_));
  NA2        g0380(.A(new_new_n144_), .B(new_new_n45_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(new_new_n402_), .Y(new_new_n404_));
  OAI210     g0382(.A0(new_new_n404_), .A1(new_new_n399_), .B0(new_new_n393_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n406_));
  NO2        g0384(.A(new_new_n150_), .B(new_new_n86_), .Y(new_new_n407_));
  OAI210     g0385(.A0(new_new_n407_), .A1(new_new_n399_), .B0(new_new_n406_), .Y(new_new_n408_));
  NO3        g0386(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n409_));
  NO2        g0387(.A(i_11_), .B(i_12_), .Y(new_new_n410_));
  NA2        g0388(.A(new_new_n401_), .B(new_new_n243_), .Y(new_new_n411_));
  NA3        g0389(.A(new_new_n112_), .B(i_4_), .C(i_11_), .Y(new_new_n412_));
  OAI220     g0390(.A0(new_new_n412_), .A1(new_new_n226_), .B0(new_new_n411_), .B1(new_new_n341_), .Y(new_new_n413_));
  NAi21      g0391(.An(i_13_), .B(i_0_), .Y(new_new_n414_));
  NO2        g0392(.A(new_new_n414_), .B(new_new_n246_), .Y(new_new_n415_));
  NA2        g0393(.A(new_new_n413_), .B(new_new_n415_), .Y(new_new_n416_));
  NA3        g0394(.A(new_new_n416_), .B(new_new_n408_), .C(new_new_n405_), .Y(new_new_n417_));
  NA2        g0395(.A(new_new_n44_), .B(new_new_n231_), .Y(new_new_n418_));
  NO3        g0396(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n419_));
  NO2        g0397(.A(i_0_), .B(i_11_), .Y(new_new_n420_));
  INV        g0398(.A(i_5_), .Y(new_new_n421_));
  AN2        g0399(.A(i_1_), .B(i_6_), .Y(new_new_n422_));
  NOi21      g0400(.An(i_2_), .B(i_12_), .Y(new_new_n423_));
  NA2        g0401(.A(new_new_n423_), .B(new_new_n422_), .Y(new_new_n424_));
  NO2        g0402(.A(new_new_n424_), .B(new_new_n421_), .Y(new_new_n425_));
  NA2        g0403(.A(new_new_n142_), .B(i_9_), .Y(new_new_n426_));
  NO2        g0404(.A(new_new_n426_), .B(i_4_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n425_), .B(new_new_n427_), .Y(new_new_n428_));
  NAi21      g0406(.An(i_9_), .B(i_4_), .Y(new_new_n429_));
  OR2        g0407(.A(i_13_), .B(i_10_), .Y(new_new_n430_));
  NO3        g0408(.A(new_new_n430_), .B(new_new_n117_), .C(new_new_n429_), .Y(new_new_n431_));
  NO2        g0409(.A(new_new_n174_), .B(new_new_n123_), .Y(new_new_n432_));
  OR2        g0410(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n433_));
  NO2        g0411(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n434_));
  NA2        g0412(.A(new_new_n291_), .B(new_new_n434_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n284_), .B(new_new_n215_), .Y(new_new_n436_));
  OAI220     g0414(.A0(new_new_n436_), .A1(new_new_n433_), .B0(new_new_n435_), .B1(new_new_n355_), .Y(new_new_n437_));
  INV        g0415(.A(new_new_n437_), .Y(new_new_n438_));
  AOI210     g0416(.A0(new_new_n438_), .A1(new_new_n428_), .B0(new_new_n26_), .Y(new_new_n439_));
  NA2        g0417(.A(new_new_n331_), .B(new_new_n330_), .Y(new_new_n440_));
  AOI220     g0418(.A0(new_new_n304_), .A1(new_new_n294_), .B0(new_new_n298_), .B1(new_new_n322_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n441_), .B(new_new_n171_), .Y(new_new_n442_));
  NO2        g0420(.A(new_new_n185_), .B(new_new_n86_), .Y(new_new_n443_));
  AOI220     g0421(.A0(new_new_n443_), .A1(new_new_n303_), .B0(new_new_n286_), .B1(new_new_n215_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n444_), .B(new_new_n293_), .Y(new_new_n445_));
  NO3        g0423(.A(new_new_n445_), .B(new_new_n442_), .C(new_new_n440_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n199_), .B(new_new_n96_), .Y(new_new_n447_));
  NA3        g0425(.A(new_new_n334_), .B(new_new_n164_), .C(new_new_n86_), .Y(new_new_n448_));
  AOI210     g0426(.A0(new_new_n448_), .A1(new_new_n447_), .B0(new_new_n332_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n304_), .B(new_new_n241_), .Y(new_new_n450_));
  NO2        g0428(.A(new_new_n450_), .B(new_new_n185_), .Y(new_new_n451_));
  NO2        g0429(.A(i_3_), .B(new_new_n48_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n451_), .B(new_new_n449_), .Y(new_new_n453_));
  AOI210     g0431(.A0(new_new_n453_), .A1(new_new_n446_), .B0(new_new_n278_), .Y(new_new_n454_));
  NO4        g0432(.A(new_new_n454_), .B(new_new_n439_), .C(new_new_n417_), .D(new_new_n392_), .Y(new_new_n455_));
  NO2        g0433(.A(new_new_n63_), .B(i_4_), .Y(new_new_n456_));
  NO2        g0434(.A(new_new_n73_), .B(i_13_), .Y(new_new_n457_));
  NO2        g0435(.A(i_10_), .B(i_9_), .Y(new_new_n458_));
  NAi21      g0436(.An(i_12_), .B(i_8_), .Y(new_new_n459_));
  NO2        g0437(.A(new_new_n459_), .B(i_3_), .Y(new_new_n460_));
  NO2        g0438(.A(new_new_n46_), .B(i_4_), .Y(new_new_n461_));
  NA2        g0439(.A(new_new_n461_), .B(new_new_n104_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n462_), .B(new_new_n208_), .Y(new_new_n463_));
  NA2        g0441(.A(new_new_n317_), .B(i_0_), .Y(new_new_n464_));
  NO3        g0442(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n273_), .B(new_new_n97_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n466_), .B(new_new_n465_), .Y(new_new_n467_));
  NA2        g0445(.A(i_8_), .B(i_9_), .Y(new_new_n468_));
  AOI210     g0446(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n469_));
  OR2        g0447(.A(new_new_n469_), .B(new_new_n468_), .Y(new_new_n470_));
  NA2        g0448(.A(new_new_n291_), .B(new_new_n209_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n471_), .B(new_new_n470_), .Y(new_new_n472_));
  NA2        g0450(.A(new_new_n257_), .B(new_new_n316_), .Y(new_new_n473_));
  NO3        g0451(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n474_));
  INV        g0452(.A(new_new_n474_), .Y(new_new_n475_));
  NA3        g0453(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n476_));
  NA4        g0454(.A(new_new_n145_), .B(new_new_n115_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n477_));
  OAI220     g0455(.A0(new_new_n477_), .A1(new_new_n476_), .B0(new_new_n475_), .B1(new_new_n473_), .Y(new_new_n478_));
  NO3        g0456(.A(new_new_n478_), .B(new_new_n472_), .C(new_new_n463_), .Y(new_new_n479_));
  OR2        g0457(.A(new_new_n302_), .B(new_new_n212_), .Y(new_new_n480_));
  BUFFER     g0458(.A(new_new_n305_), .Y(new_new_n481_));
  OA220      g0459(.A0(new_new_n481_), .A1(new_new_n163_), .B0(new_new_n480_), .B1(new_new_n238_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n96_), .B(i_13_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n443_), .B(new_new_n393_), .Y(new_new_n484_));
  NO2        g0462(.A(i_2_), .B(i_13_), .Y(new_new_n485_));
  NA3        g0463(.A(new_new_n485_), .B(new_new_n162_), .C(new_new_n99_), .Y(new_new_n486_));
  OAI220     g0464(.A0(new_new_n486_), .A1(new_new_n243_), .B0(new_new_n484_), .B1(new_new_n483_), .Y(new_new_n487_));
  NO3        g0465(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n488_));
  NO2        g0466(.A(i_6_), .B(i_7_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n490_));
  NO2        g0468(.A(i_11_), .B(i_1_), .Y(new_new_n491_));
  NO2        g0469(.A(new_new_n73_), .B(i_3_), .Y(new_new_n492_));
  OR2        g0470(.A(i_11_), .B(i_8_), .Y(new_new_n493_));
  NOi21      g0471(.An(i_2_), .B(i_7_), .Y(new_new_n494_));
  NAi31      g0472(.An(new_new_n493_), .B(new_new_n494_), .C(new_new_n492_), .Y(new_new_n495_));
  INV        g0473(.A(new_new_n430_), .Y(new_new_n496_));
  NA3        g0474(.A(new_new_n496_), .B(new_new_n456_), .C(new_new_n75_), .Y(new_new_n497_));
  NO2        g0475(.A(new_new_n497_), .B(new_new_n495_), .Y(new_new_n498_));
  NO2        g0476(.A(i_3_), .B(new_new_n196_), .Y(new_new_n499_));
  NO2        g0477(.A(i_6_), .B(i_10_), .Y(new_new_n500_));
  NA4        g0478(.A(new_new_n500_), .B(new_new_n321_), .C(new_new_n499_), .D(new_new_n243_), .Y(new_new_n501_));
  NO2        g0479(.A(new_new_n501_), .B(new_new_n156_), .Y(new_new_n502_));
  NA2        g0480(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n503_));
  NO2        g0481(.A(new_new_n158_), .B(i_3_), .Y(new_new_n504_));
  NAi31      g0482(.An(new_new_n503_), .B(new_new_n504_), .C(new_new_n232_), .Y(new_new_n505_));
  NA3        g0483(.A(new_new_n406_), .B(new_new_n181_), .C(new_new_n149_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n506_), .B(new_new_n505_), .Y(new_new_n507_));
  NO4        g0485(.A(new_new_n507_), .B(new_new_n502_), .C(new_new_n498_), .D(new_new_n487_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n474_), .B(new_new_n401_), .Y(new_new_n509_));
  NO2        g0487(.A(new_new_n509_), .B(new_new_n230_), .Y(new_new_n510_));
  NAi21      g0488(.An(new_new_n221_), .B(new_new_n410_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n346_), .B(new_new_n223_), .Y(new_new_n512_));
  NO2        g0490(.A(new_new_n26_), .B(i_5_), .Y(new_new_n513_));
  NO2        g0491(.A(i_0_), .B(new_new_n86_), .Y(new_new_n514_));
  NA3        g0492(.A(new_new_n514_), .B(new_new_n513_), .C(new_new_n142_), .Y(new_new_n515_));
  OR3        g0493(.A(new_new_n311_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n516_));
  OAI220     g0494(.A0(new_new_n516_), .A1(new_new_n515_), .B0(new_new_n512_), .B1(new_new_n511_), .Y(new_new_n517_));
  NA4        g0495(.A(new_new_n314_), .B(new_new_n229_), .C(new_new_n73_), .D(new_new_n243_), .Y(new_new_n518_));
  NO2        g0496(.A(new_new_n518_), .B(new_new_n490_), .Y(new_new_n519_));
  NO3        g0497(.A(new_new_n519_), .B(new_new_n517_), .C(new_new_n510_), .Y(new_new_n520_));
  NA4        g0498(.A(new_new_n520_), .B(new_new_n508_), .C(new_new_n482_), .D(new_new_n479_), .Y(new_new_n521_));
  NA3        g0499(.A(new_new_n314_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n522_));
  INV        g0500(.A(new_new_n522_), .Y(new_new_n523_));
  AN2        g0501(.A(new_new_n294_), .B(new_new_n240_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n524_), .B(new_new_n523_), .Y(new_new_n525_));
  NA2        g0503(.A(new_new_n122_), .B(new_new_n111_), .Y(new_new_n526_));
  AN2        g0504(.A(new_new_n526_), .B(new_new_n465_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n321_), .B(new_new_n165_), .Y(new_new_n528_));
  OAI210     g0506(.A0(new_new_n528_), .A1(new_new_n238_), .B0(new_new_n315_), .Y(new_new_n529_));
  AOI220     g0507(.A0(new_new_n529_), .A1(new_new_n333_), .B0(new_new_n527_), .B1(new_new_n317_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n394_), .B(new_new_n231_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n368_), .B(new_new_n73_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n381_), .B(new_new_n377_), .Y(new_new_n533_));
  AO210      g0511(.A0(new_new_n532_), .A1(new_new_n531_), .B0(new_new_n533_), .Y(new_new_n534_));
  NO2        g0512(.A(new_new_n36_), .B(i_8_), .Y(new_new_n535_));
  AOI210     g0513(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n431_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n536_), .B(new_new_n534_), .Y(new_new_n537_));
  INV        g0515(.A(new_new_n537_), .Y(new_new_n538_));
  NA2        g0516(.A(new_new_n263_), .B(new_new_n64_), .Y(new_new_n539_));
  OAI210     g0517(.A0(i_8_), .A1(new_new_n539_), .B0(new_new_n134_), .Y(new_new_n540_));
  NO2        g0518(.A(i_7_), .B(new_new_n202_), .Y(new_new_n541_));
  OR2        g0519(.A(new_new_n185_), .B(i_4_), .Y(new_new_n542_));
  NO2        g0520(.A(new_new_n542_), .B(new_new_n86_), .Y(new_new_n543_));
  AOI220     g0521(.A0(new_new_n543_), .A1(new_new_n541_), .B0(new_new_n540_), .B1(new_new_n432_), .Y(new_new_n544_));
  NA4        g0522(.A(new_new_n544_), .B(new_new_n538_), .C(new_new_n530_), .D(new_new_n525_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n400_), .B(new_new_n303_), .Y(new_new_n546_));
  OAI210     g0524(.A0(new_new_n396_), .A1(new_new_n170_), .B0(new_new_n546_), .Y(new_new_n547_));
  NA2        g0525(.A(new_new_n1082_), .B(new_new_n231_), .Y(new_new_n548_));
  NA2        g0526(.A(new_new_n500_), .B(new_new_n27_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n549_), .B(new_new_n548_), .Y(new_new_n550_));
  NOi31      g0528(.An(new_new_n324_), .B(new_new_n430_), .C(new_new_n38_), .Y(new_new_n551_));
  OAI210     g0529(.A0(new_new_n551_), .A1(new_new_n550_), .B0(new_new_n547_), .Y(new_new_n552_));
  NO2        g0530(.A(i_8_), .B(i_7_), .Y(new_new_n553_));
  OAI210     g0531(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n554_), .B(new_new_n229_), .Y(new_new_n555_));
  AOI220     g0533(.A0(new_new_n334_), .A1(new_new_n40_), .B0(new_new_n241_), .B1(new_new_n211_), .Y(new_new_n556_));
  OAI220     g0534(.A0(new_new_n556_), .A1(new_new_n542_), .B0(new_new_n555_), .B1(new_new_n249_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n44_), .B(i_10_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n558_), .B(i_6_), .Y(new_new_n559_));
  NA3        g0537(.A(new_new_n559_), .B(new_new_n557_), .C(new_new_n553_), .Y(new_new_n560_));
  AOI220     g0538(.A0(new_new_n443_), .A1(new_new_n334_), .B0(new_new_n253_), .B1(new_new_n250_), .Y(new_new_n561_));
  NO2        g0539(.A(new_new_n561_), .B(new_new_n269_), .Y(new_new_n562_));
  NA2        g0540(.A(new_new_n562_), .B(new_new_n272_), .Y(new_new_n563_));
  NOi31      g0541(.An(new_new_n298_), .B(new_new_n309_), .C(new_new_n183_), .Y(new_new_n564_));
  NA3        g0542(.A(new_new_n314_), .B(new_new_n176_), .C(new_new_n96_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n227_), .B(new_new_n44_), .Y(new_new_n566_));
  NO2        g0544(.A(new_new_n158_), .B(i_5_), .Y(new_new_n567_));
  NA3        g0545(.A(new_new_n567_), .B(new_new_n418_), .C(new_new_n327_), .Y(new_new_n568_));
  OAI210     g0546(.A0(new_new_n568_), .A1(new_new_n566_), .B0(new_new_n565_), .Y(new_new_n569_));
  OAI210     g0547(.A0(new_new_n569_), .A1(new_new_n564_), .B0(new_new_n474_), .Y(new_new_n570_));
  NA4        g0548(.A(new_new_n570_), .B(new_new_n563_), .C(new_new_n560_), .D(new_new_n552_), .Y(new_new_n571_));
  NA3        g0549(.A(new_new_n223_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n572_));
  NA2        g0550(.A(new_new_n291_), .B(new_new_n84_), .Y(new_new_n573_));
  AOI210     g0551(.A0(new_new_n572_), .A1(new_new_n360_), .B0(new_new_n573_), .Y(new_new_n574_));
  NA2        g0552(.A(new_new_n304_), .B(new_new_n294_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n575_), .B(new_new_n175_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n577_));
  NA2        g0555(.A(new_new_n458_), .B(new_new_n227_), .Y(new_new_n578_));
  NO2        g0556(.A(new_new_n577_), .B(new_new_n578_), .Y(new_new_n579_));
  NA2        g0557(.A(i_0_), .B(new_new_n48_), .Y(new_new_n580_));
  NO3        g0558(.A(new_new_n579_), .B(new_new_n576_), .C(new_new_n574_), .Y(new_new_n581_));
  NO4        g0559(.A(new_new_n258_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n582_));
  NO3        g0560(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n239_), .B(new_new_n36_), .Y(new_new_n584_));
  AN2        g0562(.A(new_new_n584_), .B(new_new_n583_), .Y(new_new_n585_));
  OA210      g0563(.A0(new_new_n585_), .A1(new_new_n582_), .B0(new_new_n368_), .Y(new_new_n586_));
  NO2        g0564(.A(new_new_n430_), .B(i_1_), .Y(new_new_n587_));
  NOi31      g0565(.An(new_new_n587_), .B(new_new_n466_), .C(new_new_n73_), .Y(new_new_n588_));
  AN4        g0566(.A(new_new_n588_), .B(new_new_n427_), .C(new_new_n513_), .D(i_2_), .Y(new_new_n589_));
  NO2        g0567(.A(new_new_n441_), .B(new_new_n179_), .Y(new_new_n590_));
  NO3        g0568(.A(new_new_n590_), .B(new_new_n589_), .C(new_new_n586_), .Y(new_new_n591_));
  NOi21      g0569(.An(i_10_), .B(i_6_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n593_));
  AOI220     g0571(.A0(new_new_n291_), .A1(new_new_n593_), .B0(new_new_n282_), .B1(new_new_n592_), .Y(new_new_n594_));
  NO2        g0572(.A(new_new_n594_), .B(new_new_n464_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n114_), .B(new_new_n23_), .Y(new_new_n596_));
  NA2        g0574(.A(new_new_n324_), .B(new_new_n165_), .Y(new_new_n597_));
  AOI220     g0575(.A0(new_new_n597_), .A1(new_new_n450_), .B0(new_new_n186_), .B1(new_new_n184_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n598_), .B(new_new_n595_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n532_), .B(new_new_n389_), .Y(new_new_n600_));
  INV        g0578(.A(new_new_n327_), .Y(new_new_n601_));
  NO2        g0579(.A(i_12_), .B(new_new_n86_), .Y(new_new_n602_));
  NA3        g0580(.A(new_new_n602_), .B(new_new_n282_), .C(new_new_n580_), .Y(new_new_n603_));
  NA3        g0581(.A(new_new_n397_), .B(new_new_n291_), .C(new_new_n223_), .Y(new_new_n604_));
  AOI210     g0582(.A0(new_new_n604_), .A1(new_new_n603_), .B0(new_new_n601_), .Y(new_new_n605_));
  NO3        g0583(.A(i_4_), .B(new_new_n352_), .C(new_new_n309_), .Y(new_new_n606_));
  OR2        g0584(.A(i_2_), .B(i_5_), .Y(new_new_n607_));
  OR2        g0585(.A(new_new_n607_), .B(new_new_n422_), .Y(new_new_n608_));
  NO2        g0586(.A(new_new_n608_), .B(new_new_n511_), .Y(new_new_n609_));
  NO4        g0587(.A(new_new_n609_), .B(new_new_n606_), .C(new_new_n605_), .D(new_new_n600_), .Y(new_new_n610_));
  NA4        g0588(.A(new_new_n610_), .B(new_new_n599_), .C(new_new_n591_), .D(new_new_n581_), .Y(new_new_n611_));
  NO4        g0589(.A(new_new_n611_), .B(new_new_n571_), .C(new_new_n545_), .D(new_new_n521_), .Y(new_new_n612_));
  NA4        g0590(.A(new_new_n612_), .B(new_new_n455_), .C(new_new_n367_), .D(new_new_n320_), .Y(men7));
  NO2        g0591(.A(new_new_n92_), .B(new_new_n54_), .Y(new_new_n614_));
  NO2        g0592(.A(new_new_n108_), .B(new_new_n89_), .Y(new_new_n615_));
  NA2        g0593(.A(new_new_n500_), .B(new_new_n84_), .Y(new_new_n616_));
  NA2        g0594(.A(i_11_), .B(new_new_n196_), .Y(new_new_n617_));
  NA3        g0595(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n618_));
  NO2        g0596(.A(new_new_n243_), .B(i_4_), .Y(new_new_n619_));
  NA2        g0597(.A(new_new_n619_), .B(i_8_), .Y(new_new_n620_));
  NO2        g0598(.A(new_new_n105_), .B(new_new_n618_), .Y(new_new_n621_));
  NA2        g0599(.A(i_2_), .B(new_new_n86_), .Y(new_new_n622_));
  OAI210     g0600(.A0(new_new_n87_), .A1(new_new_n206_), .B0(new_new_n207_), .Y(new_new_n623_));
  NO2        g0601(.A(i_7_), .B(new_new_n37_), .Y(new_new_n624_));
  NA2        g0602(.A(i_4_), .B(i_8_), .Y(new_new_n625_));
  AOI210     g0603(.A0(new_new_n625_), .A1(new_new_n314_), .B0(new_new_n624_), .Y(new_new_n626_));
  OAI220     g0604(.A0(new_new_n626_), .A1(new_new_n622_), .B0(new_new_n623_), .B1(i_13_), .Y(new_new_n627_));
  NO3        g0605(.A(new_new_n627_), .B(new_new_n621_), .C(new_new_n614_), .Y(new_new_n628_));
  AOI210     g0606(.A0(new_new_n128_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n629_));
  AOI210     g0607(.A0(new_new_n629_), .A1(new_new_n243_), .B0(new_new_n162_), .Y(new_new_n630_));
  OR2        g0608(.A(i_6_), .B(i_10_), .Y(new_new_n631_));
  NO2        g0609(.A(new_new_n631_), .B(new_new_n23_), .Y(new_new_n632_));
  OR3        g0610(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n633_));
  NO3        g0611(.A(new_new_n633_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n634_));
  INV        g0612(.A(new_new_n203_), .Y(new_new_n635_));
  NO2        g0613(.A(new_new_n634_), .B(new_new_n632_), .Y(new_new_n636_));
  OA220      g0614(.A0(new_new_n636_), .A1(new_new_n601_), .B0(new_new_n630_), .B1(new_new_n274_), .Y(new_new_n637_));
  AOI210     g0615(.A0(new_new_n637_), .A1(new_new_n628_), .B0(new_new_n63_), .Y(new_new_n638_));
  NOi21      g0616(.An(i_11_), .B(i_7_), .Y(new_new_n639_));
  AO210      g0617(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n640_));
  NO2        g0618(.A(new_new_n640_), .B(new_new_n639_), .Y(new_new_n641_));
  NA2        g0619(.A(new_new_n641_), .B(new_new_n211_), .Y(new_new_n642_));
  NA3        g0620(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n643_));
  NAi31      g0621(.An(new_new_n643_), .B(new_new_n220_), .C(i_11_), .Y(new_new_n644_));
  AOI210     g0622(.A0(new_new_n644_), .A1(new_new_n642_), .B0(new_new_n63_), .Y(new_new_n645_));
  NO3        g0623(.A(new_new_n265_), .B(new_new_n213_), .C(new_new_n617_), .Y(new_new_n646_));
  OAI210     g0624(.A0(new_new_n646_), .A1(new_new_n232_), .B0(new_new_n63_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n423_), .B(new_new_n31_), .Y(new_new_n648_));
  OR2        g0626(.A(new_new_n213_), .B(new_new_n108_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n649_), .B(new_new_n648_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n63_), .B(i_9_), .Y(new_new_n651_));
  NO2        g0629(.A(new_new_n651_), .B(i_4_), .Y(new_new_n652_));
  NA2        g0630(.A(new_new_n652_), .B(new_new_n650_), .Y(new_new_n653_));
  NO2        g0631(.A(i_1_), .B(i_12_), .Y(new_new_n654_));
  NA2        g0632(.A(new_new_n653_), .B(new_new_n647_), .Y(new_new_n655_));
  OAI210     g0633(.A0(new_new_n655_), .A1(new_new_n645_), .B0(i_6_), .Y(new_new_n656_));
  NO2        g0634(.A(new_new_n643_), .B(new_new_n108_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n657_), .B(new_new_n602_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n243_), .B(new_new_n86_), .Y(new_new_n659_));
  NO2        g0637(.A(new_new_n659_), .B(i_11_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n658_), .B(new_new_n467_), .Y(new_new_n661_));
  NO4        g0639(.A(new_new_n220_), .B(new_new_n128_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(new_new_n651_), .Y(new_new_n663_));
  NA2        g0641(.A(new_new_n243_), .B(i_6_), .Y(new_new_n664_));
  NO3        g0642(.A(new_new_n631_), .B(new_new_n239_), .C(new_new_n23_), .Y(new_new_n665_));
  AOI210     g0643(.A0(i_1_), .A1(new_new_n266_), .B0(new_new_n665_), .Y(new_new_n666_));
  OAI210     g0644(.A0(new_new_n666_), .A1(new_new_n44_), .B0(new_new_n663_), .Y(new_new_n667_));
  NA3        g0645(.A(new_new_n553_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n138_), .B(i_9_), .Y(new_new_n669_));
  NA3        g0647(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n670_));
  NO2        g0648(.A(new_new_n46_), .B(i_1_), .Y(new_new_n671_));
  NA3        g0649(.A(new_new_n671_), .B(new_new_n273_), .C(new_new_n44_), .Y(new_new_n672_));
  OAI220     g0650(.A0(new_new_n672_), .A1(new_new_n670_), .B0(new_new_n669_), .B1(new_new_n1080_), .Y(new_new_n673_));
  AOI210     g0651(.A0(new_new_n491_), .A1(new_new_n434_), .B0(new_new_n248_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n622_), .Y(new_new_n675_));
  NAi21      g0653(.An(new_new_n668_), .B(new_new_n91_), .Y(new_new_n676_));
  NA2        g0654(.A(new_new_n671_), .B(new_new_n273_), .Y(new_new_n677_));
  NO2        g0655(.A(i_11_), .B(new_new_n37_), .Y(new_new_n678_));
  NA2        g0656(.A(new_new_n678_), .B(new_new_n24_), .Y(new_new_n679_));
  OAI210     g0657(.A0(new_new_n679_), .A1(new_new_n677_), .B0(new_new_n676_), .Y(new_new_n680_));
  OR3        g0658(.A(new_new_n680_), .B(new_new_n675_), .C(new_new_n673_), .Y(new_new_n681_));
  NO3        g0659(.A(new_new_n681_), .B(new_new_n667_), .C(new_new_n661_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n243_), .B(new_new_n101_), .Y(new_new_n683_));
  NO2        g0661(.A(new_new_n683_), .B(new_new_n639_), .Y(new_new_n684_));
  NA2        g0662(.A(new_new_n684_), .B(i_1_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n685_), .B(new_new_n633_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n429_), .B(new_new_n86_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n686_), .B(new_new_n46_), .Y(new_new_n688_));
  NA2        g0666(.A(i_3_), .B(new_new_n196_), .Y(new_new_n689_));
  NO2        g0667(.A(new_new_n689_), .B(new_new_n114_), .Y(new_new_n690_));
  AN2        g0668(.A(new_new_n690_), .B(new_new_n559_), .Y(new_new_n691_));
  NO2        g0669(.A(new_new_n239_), .B(new_new_n44_), .Y(new_new_n692_));
  NO3        g0670(.A(new_new_n692_), .B(new_new_n317_), .C(new_new_n244_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n694_), .B(i_6_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n86_), .B(i_9_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n696_), .B(new_new_n63_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n697_), .B(new_new_n654_), .Y(new_new_n698_));
  NO4        g0676(.A(new_new_n698_), .B(new_new_n695_), .C(new_new_n693_), .D(i_4_), .Y(new_new_n699_));
  NA2        g0677(.A(i_1_), .B(i_3_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n468_), .B(new_new_n92_), .Y(new_new_n701_));
  AOI210     g0679(.A0(new_new_n692_), .A1(new_new_n592_), .B0(new_new_n701_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n702_), .B(new_new_n700_), .Y(new_new_n703_));
  NO3        g0681(.A(new_new_n703_), .B(new_new_n699_), .C(new_new_n691_), .Y(new_new_n704_));
  NA4        g0682(.A(new_new_n704_), .B(new_new_n688_), .C(new_new_n682_), .D(new_new_n656_), .Y(new_new_n705_));
  NO3        g0683(.A(new_new_n493_), .B(i_3_), .C(i_7_), .Y(new_new_n706_));
  NOi21      g0684(.An(new_new_n706_), .B(i_10_), .Y(new_new_n707_));
  OA210      g0685(.A0(new_new_n707_), .A1(new_new_n251_), .B0(new_new_n86_), .Y(new_new_n708_));
  NA2        g0686(.A(new_new_n381_), .B(new_new_n380_), .Y(new_new_n709_));
  NA3        g0687(.A(new_new_n500_), .B(new_new_n535_), .C(new_new_n46_), .Y(new_new_n710_));
  NO3        g0688(.A(new_new_n494_), .B(new_new_n625_), .C(new_new_n86_), .Y(new_new_n711_));
  NA2        g0689(.A(new_new_n711_), .B(new_new_n25_), .Y(new_new_n712_));
  NA3        g0690(.A(new_new_n162_), .B(new_new_n84_), .C(new_new_n86_), .Y(new_new_n713_));
  NA4        g0691(.A(new_new_n713_), .B(new_new_n712_), .C(new_new_n710_), .D(new_new_n709_), .Y(new_new_n714_));
  OAI210     g0692(.A0(new_new_n714_), .A1(new_new_n708_), .B0(i_1_), .Y(new_new_n715_));
  AOI210     g0693(.A0(new_new_n273_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n716_));
  NO2        g0694(.A(new_new_n379_), .B(i_2_), .Y(new_new_n717_));
  NA2        g0695(.A(new_new_n717_), .B(new_new_n716_), .Y(new_new_n718_));
  AOI210     g0696(.A0(new_new_n718_), .A1(new_new_n715_), .B0(i_13_), .Y(new_new_n719_));
  OR2        g0697(.A(i_11_), .B(i_7_), .Y(new_new_n720_));
  NO2        g0698(.A(new_new_n54_), .B(i_12_), .Y(new_new_n721_));
  INV        g0699(.A(new_new_n721_), .Y(new_new_n722_));
  NO2        g0700(.A(new_new_n494_), .B(new_new_n24_), .Y(new_new_n723_));
  AOI220     g0701(.A0(new_new_n723_), .A1(new_new_n687_), .B0(new_new_n251_), .B1(new_new_n131_), .Y(new_new_n724_));
  OAI220     g0702(.A0(new_new_n724_), .A1(new_new_n41_), .B0(new_new_n722_), .B1(new_new_n92_), .Y(new_new_n725_));
  INV        g0703(.A(new_new_n725_), .Y(new_new_n726_));
  NA2        g0704(.A(new_new_n397_), .B(new_new_n671_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n727_), .B(new_new_n249_), .Y(new_new_n728_));
  AOI210     g0706(.A0(new_new_n459_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n729_));
  NOi31      g0707(.An(new_new_n729_), .B(new_new_n616_), .C(new_new_n44_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n127_), .B(i_13_), .Y(new_new_n731_));
  NO2        g0709(.A(new_new_n670_), .B(new_new_n114_), .Y(new_new_n732_));
  INV        g0710(.A(new_new_n732_), .Y(new_new_n733_));
  NO2        g0711(.A(new_new_n731_), .B(new_new_n716_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n26_), .B(new_new_n196_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n735_), .B(i_7_), .Y(new_new_n736_));
  NO3        g0714(.A(new_new_n494_), .B(new_new_n243_), .C(new_new_n86_), .Y(new_new_n737_));
  NA2        g0715(.A(new_new_n737_), .B(new_new_n736_), .Y(new_new_n738_));
  AOI220     g0716(.A0(new_new_n397_), .A1(new_new_n671_), .B0(new_new_n91_), .B1(new_new_n102_), .Y(new_new_n739_));
  OAI220     g0717(.A0(new_new_n739_), .A1(new_new_n620_), .B0(new_new_n738_), .B1(new_new_n635_), .Y(new_new_n740_));
  NO4        g0718(.A(new_new_n740_), .B(new_new_n734_), .C(new_new_n730_), .D(new_new_n728_), .Y(new_new_n741_));
  OR2        g0719(.A(i_11_), .B(i_6_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n619_), .B(new_new_n735_), .C(i_7_), .Y(new_new_n743_));
  AOI210     g0721(.A0(new_new_n743_), .A1(new_new_n733_), .B0(new_new_n742_), .Y(new_new_n744_));
  NA3        g0722(.A(new_new_n423_), .B(new_new_n624_), .C(new_new_n97_), .Y(new_new_n745_));
  NA2        g0723(.A(new_new_n660_), .B(i_13_), .Y(new_new_n746_));
  NA2        g0724(.A(new_new_n102_), .B(new_new_n735_), .Y(new_new_n747_));
  NAi21      g0725(.An(i_11_), .B(i_12_), .Y(new_new_n748_));
  NOi41      g0726(.An(new_new_n110_), .B(new_new_n748_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n749_));
  NA2        g0727(.A(new_new_n749_), .B(new_new_n747_), .Y(new_new_n750_));
  NA3        g0728(.A(new_new_n750_), .B(new_new_n746_), .C(new_new_n745_), .Y(new_new_n751_));
  OAI210     g0729(.A0(new_new_n751_), .A1(new_new_n744_), .B0(new_new_n63_), .Y(new_new_n752_));
  NO2        g0730(.A(i_2_), .B(i_12_), .Y(new_new_n753_));
  NA2        g0731(.A(new_new_n378_), .B(new_new_n753_), .Y(new_new_n754_));
  NA2        g0732(.A(i_8_), .B(new_new_n25_), .Y(new_new_n755_));
  NO3        g0733(.A(new_new_n755_), .B(new_new_n395_), .C(new_new_n619_), .Y(new_new_n756_));
  OAI210     g0734(.A0(new_new_n756_), .A1(new_new_n380_), .B0(new_new_n378_), .Y(new_new_n757_));
  NO2        g0735(.A(new_new_n128_), .B(i_2_), .Y(new_new_n758_));
  NA2        g0736(.A(new_new_n758_), .B(new_new_n654_), .Y(new_new_n759_));
  NA3        g0737(.A(new_new_n759_), .B(new_new_n757_), .C(new_new_n754_), .Y(new_new_n760_));
  NA3        g0738(.A(new_new_n760_), .B(new_new_n45_), .C(new_new_n231_), .Y(new_new_n761_));
  NA4        g0739(.A(new_new_n761_), .B(new_new_n752_), .C(new_new_n741_), .D(new_new_n726_), .Y(new_new_n762_));
  OR4        g0740(.A(new_new_n762_), .B(new_new_n719_), .C(new_new_n705_), .D(new_new_n638_), .Y(men5));
  AOI210     g0741(.A0(new_new_n684_), .A1(new_new_n276_), .B0(new_new_n432_), .Y(new_new_n764_));
  AN2        g0742(.A(new_new_n24_), .B(i_10_), .Y(new_new_n765_));
  NA3        g0743(.A(new_new_n765_), .B(new_new_n753_), .C(new_new_n108_), .Y(new_new_n766_));
  NO2        g0744(.A(new_new_n620_), .B(i_11_), .Y(new_new_n767_));
  NA2        g0745(.A(new_new_n87_), .B(new_new_n767_), .Y(new_new_n768_));
  NA3        g0746(.A(new_new_n768_), .B(new_new_n766_), .C(new_new_n764_), .Y(new_new_n769_));
  NO3        g0747(.A(i_11_), .B(new_new_n243_), .C(i_13_), .Y(new_new_n770_));
  NO2        g0748(.A(new_new_n124_), .B(new_new_n23_), .Y(new_new_n771_));
  NA2        g0749(.A(i_12_), .B(i_8_), .Y(new_new_n772_));
  OAI210     g0750(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n772_), .Y(new_new_n773_));
  INV        g0751(.A(new_new_n458_), .Y(new_new_n774_));
  AOI220     g0752(.A0(new_new_n327_), .A1(new_new_n596_), .B0(new_new_n773_), .B1(new_new_n771_), .Y(new_new_n775_));
  INV        g0753(.A(new_new_n775_), .Y(new_new_n776_));
  NO2        g0754(.A(new_new_n776_), .B(new_new_n769_), .Y(new_new_n777_));
  INV        g0755(.A(new_new_n173_), .Y(new_new_n778_));
  INV        g0756(.A(new_new_n251_), .Y(new_new_n779_));
  OAI210     g0757(.A0(new_new_n717_), .A1(new_new_n460_), .B0(new_new_n110_), .Y(new_new_n780_));
  AOI210     g0758(.A0(new_new_n780_), .A1(new_new_n779_), .B0(new_new_n778_), .Y(new_new_n781_));
  NO2        g0759(.A(new_new_n468_), .B(new_new_n26_), .Y(new_new_n782_));
  NO2        g0760(.A(new_new_n782_), .B(new_new_n434_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(i_2_), .Y(new_new_n784_));
  INV        g0762(.A(new_new_n784_), .Y(new_new_n785_));
  AOI210     g0763(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n430_), .Y(new_new_n786_));
  AOI210     g0764(.A0(new_new_n786_), .A1(new_new_n785_), .B0(new_new_n781_), .Y(new_new_n787_));
  NO2        g0765(.A(new_new_n193_), .B(new_new_n125_), .Y(new_new_n788_));
  OAI210     g0766(.A0(new_new_n788_), .A1(new_new_n771_), .B0(i_2_), .Y(new_new_n789_));
  INV        g0767(.A(new_new_n174_), .Y(new_new_n790_));
  NO3        g0768(.A(new_new_n640_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n791_));
  AOI210     g0769(.A0(new_new_n790_), .A1(new_new_n87_), .B0(new_new_n791_), .Y(new_new_n792_));
  AOI210     g0770(.A0(new_new_n792_), .A1(new_new_n789_), .B0(new_new_n196_), .Y(new_new_n793_));
  OA210      g0771(.A0(new_new_n641_), .A1(new_new_n126_), .B0(i_13_), .Y(new_new_n794_));
  NA2        g0772(.A(new_new_n203_), .B(new_new_n206_), .Y(new_new_n795_));
  NA2        g0773(.A(new_new_n152_), .B(new_new_n617_), .Y(new_new_n796_));
  AOI210     g0774(.A0(new_new_n796_), .A1(new_new_n795_), .B0(new_new_n383_), .Y(new_new_n797_));
  AOI210     g0775(.A0(new_new_n213_), .A1(new_new_n148_), .B0(new_new_n535_), .Y(new_new_n798_));
  NA2        g0776(.A(new_new_n798_), .B(new_new_n434_), .Y(new_new_n799_));
  NO2        g0777(.A(new_new_n102_), .B(new_new_n44_), .Y(new_new_n800_));
  INV        g0778(.A(new_new_n310_), .Y(new_new_n801_));
  NA4        g0779(.A(new_new_n801_), .B(new_new_n314_), .C(new_new_n124_), .D(new_new_n42_), .Y(new_new_n802_));
  OAI210     g0780(.A0(new_new_n802_), .A1(new_new_n800_), .B0(new_new_n799_), .Y(new_new_n803_));
  NO4        g0781(.A(new_new_n803_), .B(new_new_n797_), .C(new_new_n794_), .D(new_new_n793_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n596_), .B(new_new_n28_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n770_), .B(new_new_n283_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n806_), .B(new_new_n805_), .Y(new_new_n807_));
  NO2        g0785(.A(new_new_n62_), .B(i_12_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n808_), .B(new_new_n126_), .Y(new_new_n809_));
  NO2        g0787(.A(new_new_n809_), .B(new_new_n617_), .Y(new_new_n810_));
  AOI220     g0788(.A0(new_new_n810_), .A1(new_new_n36_), .B0(new_new_n807_), .B1(new_new_n46_), .Y(new_new_n811_));
  NA4        g0789(.A(new_new_n811_), .B(new_new_n804_), .C(new_new_n787_), .D(new_new_n777_), .Y(men6));
  NO3        g0790(.A(new_new_n261_), .B(new_new_n316_), .C(i_1_), .Y(new_new_n813_));
  NO2        g0791(.A(new_new_n188_), .B(new_new_n139_), .Y(new_new_n814_));
  OAI210     g0792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n758_), .Y(new_new_n815_));
  NA4        g0793(.A(new_new_n401_), .B(new_new_n499_), .C(new_new_n71_), .D(new_new_n101_), .Y(new_new_n816_));
  INV        g0794(.A(new_new_n816_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n226_), .B(new_new_n503_), .Y(new_new_n818_));
  NO2        g0796(.A(new_new_n817_), .B(new_new_n339_), .Y(new_new_n819_));
  AO210      g0797(.A0(new_new_n819_), .A1(new_new_n815_), .B0(i_12_), .Y(new_new_n820_));
  NA2        g0798(.A(new_new_n602_), .B(new_new_n63_), .Y(new_new_n821_));
  NA2        g0799(.A(new_new_n707_), .B(new_new_n71_), .Y(new_new_n822_));
  NA2        g0800(.A(new_new_n822_), .B(new_new_n821_), .Y(new_new_n823_));
  NA2        g0801(.A(new_new_n823_), .B(new_new_n73_), .Y(new_new_n824_));
  INV        g0802(.A(new_new_n338_), .Y(new_new_n825_));
  NA2        g0803(.A(new_new_n75_), .B(new_new_n131_), .Y(new_new_n826_));
  INV        g0804(.A(new_new_n124_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n827_), .B(new_new_n46_), .Y(new_new_n828_));
  AOI210     g0806(.A0(new_new_n828_), .A1(new_new_n826_), .B0(new_new_n825_), .Y(new_new_n829_));
  NO2        g0807(.A(new_new_n258_), .B(i_9_), .Y(new_new_n830_));
  NA2        g0808(.A(new_new_n830_), .B(new_new_n808_), .Y(new_new_n831_));
  AOI210     g0809(.A0(new_new_n831_), .A1(new_new_n533_), .B0(new_new_n188_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n32_), .B(i_11_), .Y(new_new_n833_));
  NA3        g0811(.A(new_new_n833_), .B(new_new_n489_), .C(new_new_n401_), .Y(new_new_n834_));
  NAi32      g0812(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n835_));
  NO2        g0813(.A(new_new_n742_), .B(new_new_n835_), .Y(new_new_n836_));
  OAI210     g0814(.A0(new_new_n706_), .A1(new_new_n584_), .B0(new_new_n583_), .Y(new_new_n837_));
  NAi31      g0815(.An(new_new_n836_), .B(new_new_n837_), .C(new_new_n834_), .Y(new_new_n838_));
  OR3        g0816(.A(new_new_n838_), .B(new_new_n832_), .C(new_new_n829_), .Y(new_new_n839_));
  NO2        g0817(.A(new_new_n720_), .B(i_2_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n841_));
  NO2        g0819(.A(new_new_n841_), .B(new_new_n422_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n842_), .B(new_new_n840_), .Y(new_new_n843_));
  AO210      g0821(.A0(new_new_n372_), .A1(new_new_n364_), .B0(new_new_n409_), .Y(new_new_n844_));
  NA3        g0822(.A(new_new_n844_), .B(new_new_n262_), .C(i_7_), .Y(new_new_n845_));
  BUFFER     g0823(.A(new_new_n641_), .Y(new_new_n846_));
  NA3        g0824(.A(new_new_n846_), .B(new_new_n147_), .C(new_new_n69_), .Y(new_new_n847_));
  AO210      g0825(.A0(new_new_n509_), .A1(new_new_n774_), .B0(new_new_n36_), .Y(new_new_n848_));
  NA4        g0826(.A(new_new_n848_), .B(new_new_n847_), .C(new_new_n845_), .D(new_new_n843_), .Y(new_new_n849_));
  NO2        g0827(.A(new_new_n659_), .B(i_11_), .Y(new_new_n850_));
  AOI220     g0828(.A0(new_new_n850_), .A1(new_new_n583_), .B0(new_new_n818_), .B1(new_new_n736_), .Y(new_new_n851_));
  NA3        g0829(.A(new_new_n383_), .B(new_new_n245_), .C(new_new_n147_), .Y(new_new_n852_));
  NA2        g0830(.A(new_new_n409_), .B(new_new_n70_), .Y(new_new_n853_));
  NA4        g0831(.A(new_new_n853_), .B(new_new_n852_), .C(new_new_n851_), .D(new_new_n623_), .Y(new_new_n854_));
  AOI210     g0832(.A0(new_new_n460_), .A1(new_new_n458_), .B0(new_new_n582_), .Y(new_new_n855_));
  NA2        g0833(.A(new_new_n111_), .B(new_new_n420_), .Y(new_new_n856_));
  NA2        g0834(.A(new_new_n250_), .B(new_new_n46_), .Y(new_new_n857_));
  INV        g0835(.A(new_new_n608_), .Y(new_new_n858_));
  NA3        g0836(.A(new_new_n858_), .B(new_new_n338_), .C(i_7_), .Y(new_new_n859_));
  NA3        g0837(.A(new_new_n859_), .B(new_new_n856_), .C(new_new_n855_), .Y(new_new_n860_));
  NO4        g0838(.A(new_new_n860_), .B(new_new_n854_), .C(new_new_n849_), .D(new_new_n839_), .Y(new_new_n861_));
  NA4        g0839(.A(new_new_n861_), .B(new_new_n824_), .C(new_new_n820_), .D(new_new_n391_), .Y(men3));
  NA2        g0840(.A(i_12_), .B(i_10_), .Y(new_new_n863_));
  NA2        g0841(.A(i_6_), .B(i_7_), .Y(new_new_n864_));
  NO2        g0842(.A(new_new_n864_), .B(i_0_), .Y(new_new_n865_));
  NO2        g0843(.A(i_11_), .B(new_new_n243_), .Y(new_new_n866_));
  OAI210     g0844(.A0(new_new_n865_), .A1(new_new_n298_), .B0(new_new_n866_), .Y(new_new_n867_));
  NO2        g0845(.A(new_new_n867_), .B(new_new_n196_), .Y(new_new_n868_));
  NO3        g0846(.A(new_new_n464_), .B(new_new_n89_), .C(new_new_n44_), .Y(new_new_n869_));
  OA210      g0847(.A0(new_new_n869_), .A1(new_new_n868_), .B0(new_new_n176_), .Y(new_new_n870_));
  NA3        g0848(.A(new_new_n852_), .B(new_new_n623_), .C(new_new_n382_), .Y(new_new_n871_));
  NA2        g0849(.A(new_new_n871_), .B(new_new_n40_), .Y(new_new_n872_));
  NO3        g0850(.A(new_new_n649_), .B(new_new_n468_), .C(new_new_n131_), .Y(new_new_n873_));
  AN2        g0851(.A(new_new_n466_), .B(new_new_n55_), .Y(new_new_n874_));
  NO2        g0852(.A(new_new_n874_), .B(new_new_n873_), .Y(new_new_n875_));
  AOI210     g0853(.A0(new_new_n875_), .A1(new_new_n872_), .B0(new_new_n48_), .Y(new_new_n876_));
  NO4        g0854(.A(new_new_n387_), .B(new_new_n394_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n188_), .B(new_new_n592_), .Y(new_new_n878_));
  NOi21      g0856(.An(new_new_n878_), .B(new_new_n877_), .Y(new_new_n879_));
  NA2        g0857(.A(new_new_n729_), .B(new_new_n696_), .Y(new_new_n880_));
  NA2        g0858(.A(new_new_n344_), .B(new_new_n452_), .Y(new_new_n881_));
  OAI220     g0859(.A0(new_new_n881_), .A1(new_new_n880_), .B0(new_new_n879_), .B1(new_new_n63_), .Y(new_new_n882_));
  NOi21      g0860(.An(i_5_), .B(i_9_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n883_), .B(new_new_n457_), .Y(new_new_n884_));
  AOI210     g0862(.A0(new_new_n273_), .A1(new_new_n491_), .B0(new_new_n711_), .Y(new_new_n885_));
  NO3        g0863(.A(new_new_n426_), .B(new_new_n273_), .C(new_new_n73_), .Y(new_new_n886_));
  NO2        g0864(.A(new_new_n177_), .B(new_new_n148_), .Y(new_new_n887_));
  AOI210     g0865(.A0(new_new_n887_), .A1(new_new_n250_), .B0(new_new_n886_), .Y(new_new_n888_));
  OAI220     g0866(.A0(new_new_n888_), .A1(new_new_n183_), .B0(new_new_n885_), .B1(new_new_n884_), .Y(new_new_n889_));
  NO4        g0867(.A(new_new_n889_), .B(new_new_n882_), .C(new_new_n876_), .D(new_new_n870_), .Y(new_new_n890_));
  NA2        g0868(.A(new_new_n188_), .B(new_new_n24_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n321_), .B(new_new_n129_), .Y(new_new_n892_));
  NAi21      g0870(.An(new_new_n163_), .B(new_new_n452_), .Y(new_new_n893_));
  OAI220     g0871(.A0(new_new_n893_), .A1(new_new_n857_), .B0(new_new_n892_), .B1(new_new_n411_), .Y(new_new_n894_));
  INV        g0872(.A(new_new_n894_), .Y(new_new_n895_));
  NO2        g0873(.A(new_new_n401_), .B(new_new_n302_), .Y(new_new_n896_));
  NA2        g0874(.A(new_new_n896_), .B(new_new_n732_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n593_), .B(i_0_), .Y(new_new_n898_));
  NO3        g0876(.A(new_new_n898_), .B(new_new_n396_), .C(new_new_n87_), .Y(new_new_n899_));
  INV        g0877(.A(new_new_n899_), .Y(new_new_n900_));
  INV        g0878(.A(new_new_n489_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n770_), .B(new_new_n339_), .Y(new_new_n902_));
  INV        g0880(.A(new_new_n58_), .Y(new_new_n903_));
  OAI220     g0881(.A0(new_new_n903_), .A1(new_new_n902_), .B0(new_new_n679_), .B1(new_new_n555_), .Y(new_new_n904_));
  NO2        g0882(.A(new_new_n260_), .B(new_new_n154_), .Y(new_new_n905_));
  NA2        g0883(.A(i_0_), .B(i_10_), .Y(new_new_n906_));
  OAI210     g0884(.A0(new_new_n906_), .A1(new_new_n86_), .B0(new_new_n558_), .Y(new_new_n907_));
  NO4        g0885(.A(new_new_n114_), .B(new_new_n58_), .C(new_new_n689_), .D(i_5_), .Y(new_new_n908_));
  AO220      g0886(.A0(new_new_n908_), .A1(new_new_n907_), .B0(new_new_n905_), .B1(i_6_), .Y(new_new_n909_));
  AOI220     g0887(.A0(new_new_n344_), .A1(new_new_n98_), .B0(new_new_n188_), .B1(new_new_n84_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n587_), .B(i_4_), .Y(new_new_n911_));
  NA2        g0889(.A(new_new_n191_), .B(new_new_n206_), .Y(new_new_n912_));
  OAI220     g0890(.A0(new_new_n912_), .A1(new_new_n902_), .B0(new_new_n911_), .B1(new_new_n910_), .Y(new_new_n913_));
  NO3        g0891(.A(new_new_n913_), .B(new_new_n909_), .C(new_new_n904_), .Y(new_new_n914_));
  NA4        g0892(.A(new_new_n914_), .B(new_new_n900_), .C(new_new_n897_), .D(new_new_n895_), .Y(new_new_n915_));
  NO2        g0893(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n916_));
  NA2        g0894(.A(i_11_), .B(i_9_), .Y(new_new_n917_));
  NO3        g0895(.A(i_12_), .B(new_new_n917_), .C(new_new_n622_), .Y(new_new_n918_));
  AN2        g0896(.A(new_new_n918_), .B(new_new_n916_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n48_), .B(i_7_), .Y(new_new_n920_));
  NA2        g0898(.A(new_new_n406_), .B(new_new_n181_), .Y(new_new_n921_));
  NA2        g0899(.A(new_new_n921_), .B(new_new_n161_), .Y(new_new_n922_));
  NO2        g0900(.A(new_new_n917_), .B(new_new_n73_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n177_), .B(i_0_), .Y(new_new_n924_));
  INV        g0902(.A(new_new_n924_), .Y(new_new_n925_));
  NA2        g0903(.A(new_new_n489_), .B(new_new_n237_), .Y(new_new_n926_));
  INV        g0904(.A(new_new_n419_), .Y(new_new_n927_));
  OAI220     g0905(.A0(new_new_n927_), .A1(new_new_n884_), .B0(new_new_n926_), .B1(new_new_n925_), .Y(new_new_n928_));
  NO3        g0906(.A(new_new_n928_), .B(new_new_n922_), .C(new_new_n919_), .Y(new_new_n929_));
  NA2        g0907(.A(new_new_n678_), .B(new_new_n121_), .Y(new_new_n930_));
  NO2        g0908(.A(i_6_), .B(new_new_n930_), .Y(new_new_n931_));
  AOI210     g0909(.A0(new_new_n459_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n173_), .B(new_new_n103_), .Y(new_new_n933_));
  NOi32      g0911(.An(new_new_n932_), .Bn(new_new_n191_), .C(new_new_n933_), .Y(new_new_n934_));
  NO2        g0912(.A(new_new_n934_), .B(new_new_n931_), .Y(new_new_n935_));
  NOi21      g0913(.An(i_7_), .B(i_5_), .Y(new_new_n936_));
  NOi31      g0914(.An(new_new_n936_), .B(i_0_), .C(new_new_n748_), .Y(new_new_n937_));
  NA3        g0915(.A(new_new_n937_), .B(new_new_n395_), .C(i_6_), .Y(new_new_n938_));
  OA210      g0916(.A0(new_new_n933_), .A1(new_new_n533_), .B0(new_new_n938_), .Y(new_new_n939_));
  NO3        g0917(.A(new_new_n414_), .B(new_new_n375_), .C(new_new_n371_), .Y(new_new_n940_));
  NO2        g0918(.A(new_new_n267_), .B(new_new_n328_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n748_), .B(new_new_n264_), .Y(new_new_n942_));
  AOI210     g0920(.A0(new_new_n942_), .A1(new_new_n941_), .B0(new_new_n940_), .Y(new_new_n943_));
  NA4        g0921(.A(new_new_n943_), .B(new_new_n939_), .C(new_new_n935_), .D(new_new_n929_), .Y(new_new_n944_));
  NO2        g0922(.A(new_new_n891_), .B(new_new_n246_), .Y(new_new_n945_));
  AN2        g0923(.A(new_new_n343_), .B(new_new_n339_), .Y(new_new_n946_));
  AN2        g0924(.A(new_new_n946_), .B(new_new_n887_), .Y(new_new_n947_));
  OAI210     g0925(.A0(new_new_n947_), .A1(new_new_n945_), .B0(i_10_), .Y(new_new_n948_));
  NO2        g0926(.A(new_new_n863_), .B(new_new_n327_), .Y(new_new_n949_));
  NA2        g0927(.A(new_new_n949_), .B(new_new_n923_), .Y(new_new_n950_));
  NA3        g0928(.A(new_new_n488_), .B(new_new_n423_), .C(new_new_n45_), .Y(new_new_n951_));
  OAI210     g0929(.A0(new_new_n893_), .A1(new_new_n901_), .B0(new_new_n951_), .Y(new_new_n952_));
  NO2        g0930(.A(new_new_n262_), .B(new_new_n46_), .Y(new_new_n953_));
  NO2        g0931(.A(new_new_n953_), .B(new_new_n190_), .Y(new_new_n954_));
  AOI220     g0932(.A0(new_new_n954_), .A1(new_new_n489_), .B0(new_new_n952_), .B1(new_new_n73_), .Y(new_new_n955_));
  NA3        g0933(.A(new_new_n841_), .B(new_new_n393_), .C(new_new_n659_), .Y(new_new_n956_));
  NA2        g0934(.A(new_new_n92_), .B(new_new_n44_), .Y(new_new_n957_));
  NO2        g0935(.A(new_new_n75_), .B(new_new_n772_), .Y(new_new_n958_));
  AOI220     g0936(.A0(new_new_n958_), .A1(new_new_n957_), .B0(new_new_n176_), .B1(new_new_n615_), .Y(new_new_n959_));
  AOI210     g0937(.A0(new_new_n959_), .A1(new_new_n956_), .B0(new_new_n47_), .Y(new_new_n960_));
  NA2        g0938(.A(new_new_n723_), .B(new_new_n567_), .Y(new_new_n961_));
  NO2        g0939(.A(new_new_n618_), .B(new_new_n105_), .Y(new_new_n962_));
  NA2        g0940(.A(new_new_n962_), .B(i_0_), .Y(new_new_n963_));
  OAI220     g0941(.A0(new_new_n963_), .A1(new_new_n86_), .B0(new_new_n961_), .B1(new_new_n174_), .Y(new_new_n964_));
  NO3        g0942(.A(new_new_n964_), .B(new_new_n960_), .C(new_new_n537_), .Y(new_new_n965_));
  NA4        g0943(.A(new_new_n965_), .B(new_new_n955_), .C(new_new_n950_), .D(new_new_n948_), .Y(new_new_n966_));
  NO3        g0944(.A(new_new_n966_), .B(new_new_n944_), .C(new_new_n915_), .Y(new_new_n967_));
  NO2        g0945(.A(i_0_), .B(new_new_n748_), .Y(new_new_n968_));
  NA2        g0946(.A(new_new_n73_), .B(new_new_n44_), .Y(new_new_n969_));
  NA2        g0947(.A(new_new_n906_), .B(new_new_n969_), .Y(new_new_n970_));
  NO3        g0948(.A(new_new_n105_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n971_));
  AO220      g0949(.A0(new_new_n971_), .A1(new_new_n970_), .B0(new_new_n968_), .B1(new_new_n176_), .Y(new_new_n972_));
  AOI210     g0950(.A0(new_new_n821_), .A1(new_new_n709_), .B0(new_new_n933_), .Y(new_new_n973_));
  AOI210     g0951(.A0(new_new_n972_), .A1(new_new_n361_), .B0(new_new_n973_), .Y(new_new_n974_));
  NA2        g0952(.A(new_new_n758_), .B(new_new_n146_), .Y(new_new_n975_));
  INV        g0953(.A(new_new_n975_), .Y(new_new_n976_));
  NA3        g0954(.A(new_new_n976_), .B(new_new_n696_), .C(new_new_n73_), .Y(new_new_n977_));
  NO2        g0955(.A(new_new_n837_), .B(new_new_n414_), .Y(new_new_n978_));
  NA3        g0956(.A(new_new_n865_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n866_), .B(i_9_), .Y(new_new_n980_));
  AOI210     g0958(.A0(new_new_n979_), .A1(new_new_n515_), .B0(new_new_n980_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n250_), .B(new_new_n236_), .Y(new_new_n982_));
  AOI210     g0960(.A0(new_new_n982_), .A1(new_new_n898_), .B0(new_new_n154_), .Y(new_new_n983_));
  NO3        g0961(.A(new_new_n983_), .B(new_new_n981_), .C(new_new_n978_), .Y(new_new_n984_));
  NA3        g0962(.A(new_new_n984_), .B(new_new_n977_), .C(new_new_n974_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n946_), .B(new_new_n383_), .Y(new_new_n986_));
  AOI210     g0964(.A0(new_new_n309_), .A1(new_new_n163_), .B0(new_new_n986_), .Y(new_new_n987_));
  NA3        g0965(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n920_), .B(new_new_n504_), .Y(new_new_n989_));
  AOI210     g0967(.A0(new_new_n988_), .A1(new_new_n163_), .B0(new_new_n989_), .Y(new_new_n990_));
  NO2        g0968(.A(new_new_n990_), .B(new_new_n987_), .Y(new_new_n991_));
  NO3        g0969(.A(new_new_n906_), .B(new_new_n883_), .C(new_new_n193_), .Y(new_new_n992_));
  AOI220     g0970(.A0(new_new_n992_), .A1(i_11_), .B0(new_new_n588_), .B1(new_new_n75_), .Y(new_new_n993_));
  NO3        g0971(.A(new_new_n214_), .B(new_new_n394_), .C(i_0_), .Y(new_new_n994_));
  OAI210     g0972(.A0(new_new_n994_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n995_));
  INV        g0973(.A(new_new_n223_), .Y(new_new_n996_));
  OAI220     g0974(.A0(new_new_n548_), .A1(new_new_n139_), .B0(new_new_n664_), .B1(new_new_n635_), .Y(new_new_n997_));
  NA3        g0975(.A(new_new_n997_), .B(i_7_), .C(new_new_n996_), .Y(new_new_n998_));
  NA4        g0976(.A(new_new_n998_), .B(new_new_n995_), .C(new_new_n993_), .D(new_new_n991_), .Y(new_new_n999_));
  NO2        g0977(.A(new_new_n249_), .B(new_new_n92_), .Y(new_new_n1000_));
  NA2        g0978(.A(new_new_n1000_), .B(new_new_n968_), .Y(new_new_n1001_));
  AOI220     g0979(.A0(new_new_n936_), .A1(new_new_n504_), .B0(new_new_n865_), .B1(new_new_n164_), .Y(new_new_n1002_));
  NA2        g0980(.A(new_new_n364_), .B(new_new_n178_), .Y(new_new_n1003_));
  OA220      g0981(.A0(new_new_n1003_), .A1(new_new_n1002_), .B0(new_new_n1001_), .B1(i_5_), .Y(new_new_n1004_));
  AOI210     g0982(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n177_), .Y(new_new_n1005_));
  NA3        g0983(.A(new_new_n632_), .B(new_new_n188_), .C(new_new_n84_), .Y(new_new_n1006_));
  NA2        g0984(.A(new_new_n1006_), .B(new_new_n565_), .Y(new_new_n1007_));
  INV        g0985(.A(new_new_n486_), .Y(new_new_n1008_));
  NO2        g0986(.A(new_new_n1008_), .B(new_new_n1007_), .Y(new_new_n1009_));
  NA3        g0987(.A(new_new_n401_), .B(new_new_n173_), .C(new_new_n172_), .Y(new_new_n1010_));
  NA3        g0988(.A(new_new_n401_), .B(new_new_n345_), .C(new_new_n227_), .Y(new_new_n1011_));
  INV        g0989(.A(new_new_n1011_), .Y(new_new_n1012_));
  NOi31      g0990(.An(new_new_n400_), .B(new_new_n969_), .C(new_new_n246_), .Y(new_new_n1013_));
  NO3        g0991(.A(new_new_n917_), .B(new_new_n223_), .C(new_new_n193_), .Y(new_new_n1014_));
  NO4        g0992(.A(new_new_n1014_), .B(new_new_n1013_), .C(new_new_n1012_), .D(new_new_n1081_), .Y(new_new_n1015_));
  NA3        g0993(.A(new_new_n1015_), .B(new_new_n1009_), .C(new_new_n1004_), .Y(new_new_n1016_));
  INV        g0994(.A(new_new_n634_), .Y(new_new_n1017_));
  NO3        g0995(.A(new_new_n1017_), .B(new_new_n580_), .C(new_new_n358_), .Y(new_new_n1018_));
  NO2        g0996(.A(new_new_n86_), .B(i_5_), .Y(new_new_n1019_));
  NA3        g0997(.A(new_new_n866_), .B(new_new_n109_), .C(new_new_n124_), .Y(new_new_n1020_));
  INV        g0998(.A(new_new_n1020_), .Y(new_new_n1021_));
  AOI210     g0999(.A0(new_new_n1021_), .A1(new_new_n1019_), .B0(new_new_n1018_), .Y(new_new_n1022_));
  NA3        g1000(.A(new_new_n314_), .B(i_5_), .C(new_new_n196_), .Y(new_new_n1023_));
  NAi31      g1001(.An(new_new_n248_), .B(new_new_n1023_), .C(new_new_n249_), .Y(new_new_n1024_));
  NO4        g1002(.A(new_new_n246_), .B(new_new_n214_), .C(i_0_), .D(i_12_), .Y(new_new_n1025_));
  AOI220     g1003(.A0(new_new_n1025_), .A1(new_new_n1024_), .B0(new_new_n817_), .B1(new_new_n178_), .Y(new_new_n1026_));
  AN2        g1004(.A(new_new_n906_), .B(new_new_n154_), .Y(new_new_n1027_));
  NO4        g1005(.A(new_new_n1027_), .B(i_12_), .C(new_new_n668_), .D(new_new_n131_), .Y(new_new_n1028_));
  NA2        g1006(.A(new_new_n1028_), .B(new_new_n223_), .Y(new_new_n1029_));
  NA3        g1007(.A(new_new_n98_), .B(new_new_n592_), .C(i_11_), .Y(new_new_n1030_));
  NO2        g1008(.A(new_new_n1030_), .B(new_new_n156_), .Y(new_new_n1031_));
  NA2        g1009(.A(new_new_n936_), .B(new_new_n485_), .Y(new_new_n1032_));
  NA2        g1010(.A(new_new_n64_), .B(new_new_n101_), .Y(new_new_n1033_));
  OAI220     g1011(.A0(new_new_n1033_), .A1(new_new_n1023_), .B0(new_new_n1032_), .B1(new_new_n697_), .Y(new_new_n1034_));
  AOI210     g1012(.A0(new_new_n1034_), .A1(new_new_n924_), .B0(new_new_n1031_), .Y(new_new_n1035_));
  NA4        g1013(.A(new_new_n1035_), .B(new_new_n1029_), .C(new_new_n1026_), .D(new_new_n1022_), .Y(new_new_n1036_));
  NO4        g1014(.A(new_new_n1036_), .B(new_new_n1016_), .C(new_new_n999_), .D(new_new_n985_), .Y(new_new_n1037_));
  OAI210     g1015(.A0(new_new_n840_), .A1(new_new_n833_), .B0(new_new_n37_), .Y(new_new_n1038_));
  NA3        g1016(.A(new_new_n932_), .B(new_new_n378_), .C(i_5_), .Y(new_new_n1039_));
  NA3        g1017(.A(new_new_n1039_), .B(new_new_n1038_), .C(new_new_n630_), .Y(new_new_n1040_));
  NA2        g1018(.A(new_new_n1040_), .B(new_new_n211_), .Y(new_new_n1041_));
  NA2        g1019(.A(new_new_n189_), .B(new_new_n191_), .Y(new_new_n1042_));
  AO210      g1020(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n1042_), .Y(new_new_n1043_));
  OAI210     g1021(.A0(new_new_n634_), .A1(new_new_n632_), .B0(new_new_n327_), .Y(new_new_n1044_));
  INV        g1022(.A(new_new_n665_), .Y(new_new_n1045_));
  NA3        g1023(.A(new_new_n1045_), .B(new_new_n1044_), .C(new_new_n1043_), .Y(new_new_n1046_));
  NO2        g1024(.A(new_new_n476_), .B(new_new_n273_), .Y(new_new_n1047_));
  NO4        g1025(.A(new_new_n239_), .B(new_new_n145_), .C(new_new_n700_), .D(new_new_n37_), .Y(new_new_n1048_));
  NO2        g1026(.A(new_new_n1048_), .B(new_new_n1047_), .Y(new_new_n1049_));
  OAI210     g1027(.A0(new_new_n1030_), .A1(new_new_n148_), .B0(new_new_n1049_), .Y(new_new_n1050_));
  AOI210     g1028(.A0(new_new_n1046_), .A1(new_new_n48_), .B0(new_new_n1050_), .Y(new_new_n1051_));
  AOI210     g1029(.A0(new_new_n1051_), .A1(new_new_n1041_), .B0(new_new_n73_), .Y(new_new_n1052_));
  NO2        g1030(.A(new_new_n585_), .B(new_new_n390_), .Y(new_new_n1053_));
  NO2        g1031(.A(new_new_n1053_), .B(new_new_n778_), .Y(new_new_n1054_));
  INV        g1032(.A(new_new_n76_), .Y(new_new_n1055_));
  AOI210     g1033(.A0(new_new_n1005_), .A1(new_new_n920_), .B0(new_new_n937_), .Y(new_new_n1056_));
  AOI210     g1034(.A0(new_new_n1056_), .A1(new_new_n1055_), .B0(new_new_n700_), .Y(new_new_n1057_));
  NA2        g1035(.A(new_new_n267_), .B(new_new_n57_), .Y(new_new_n1058_));
  AOI220     g1036(.A0(new_new_n1058_), .A1(new_new_n76_), .B0(new_new_n359_), .B1(new_new_n261_), .Y(new_new_n1059_));
  NO2        g1037(.A(new_new_n1059_), .B(new_new_n243_), .Y(new_new_n1060_));
  NA3        g1038(.A(new_new_n96_), .B(new_new_n316_), .C(new_new_n31_), .Y(new_new_n1061_));
  INV        g1039(.A(new_new_n1061_), .Y(new_new_n1062_));
  NO3        g1040(.A(new_new_n1062_), .B(new_new_n1060_), .C(new_new_n1057_), .Y(new_new_n1063_));
  OAI210     g1041(.A0(new_new_n275_), .A1(new_new_n159_), .B0(new_new_n87_), .Y(new_new_n1064_));
  NA3        g1042(.A(new_new_n782_), .B(new_new_n298_), .C(new_new_n80_), .Y(new_new_n1065_));
  AOI210     g1043(.A0(new_new_n1065_), .A1(new_new_n1064_), .B0(i_11_), .Y(new_new_n1066_));
  NA2        g1044(.A(new_new_n625_), .B(new_new_n220_), .Y(new_new_n1067_));
  OAI210     g1045(.A0(new_new_n1067_), .A1(new_new_n932_), .B0(new_new_n211_), .Y(new_new_n1068_));
  NA2        g1046(.A(new_new_n165_), .B(i_5_), .Y(new_new_n1069_));
  NO2        g1047(.A(new_new_n1068_), .B(new_new_n1069_), .Y(new_new_n1070_));
  NO3        g1048(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1071_));
  OAI210     g1049(.A0(new_new_n941_), .A1(new_new_n316_), .B0(new_new_n1071_), .Y(new_new_n1072_));
  NO2        g1050(.A(new_new_n1072_), .B(new_new_n748_), .Y(new_new_n1073_));
  NO3        g1051(.A(new_new_n1073_), .B(new_new_n1070_), .C(new_new_n1066_), .Y(new_new_n1074_));
  OAI210     g1052(.A0(new_new_n1063_), .A1(i_4_), .B0(new_new_n1074_), .Y(new_new_n1075_));
  NO3        g1053(.A(new_new_n1075_), .B(new_new_n1054_), .C(new_new_n1052_), .Y(new_new_n1076_));
  NA4        g1054(.A(new_new_n1076_), .B(new_new_n1037_), .C(new_new_n967_), .D(new_new_n890_), .Y(men4));
  INV        g1055(.A(i_2_), .Y(new_new_n1080_));
  INV        g1056(.A(new_new_n1010_), .Y(new_new_n1081_));
  INV        g1057(.A(i_12_), .Y(new_new_n1082_));
endmodule


