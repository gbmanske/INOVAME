//Benchmark atmr_misex3_1774_0.0156

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1533_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1540_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1543_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1549_, mai_mai_n1550_, mai_mai_n1551_, mai_mai_n1552_, mai_mai_n1556_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1609_, men_men_n1610_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(g), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(g), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o0010(.A(ori_ori_n38_), .B(n), .Y(ori_ori_n39_));
  INV        o0011(.A(h), .Y(ori_ori_n40_));
  NAi21      o0012(.An(j), .B(l), .Y(ori_ori_n41_));
  NAi32      o0013(.An(n), .Bn(g), .C(m), .Y(ori_ori_n42_));
  NO3        o0014(.A(ori_ori_n42_), .B(ori_ori_n41_), .C(ori_ori_n40_), .Y(ori_ori_n43_));
  NAi31      o0015(.An(n), .B(m), .C(l), .Y(ori_ori_n44_));
  INV        o0016(.A(i), .Y(ori_ori_n45_));
  AN2        o0017(.A(h), .B(g), .Y(ori_ori_n46_));
  NA2        o0018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NAi21      o0020(.An(n), .B(m), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(l), .Y(ori_ori_n50_));
  NOi32      o0022(.An(k), .Bn(h), .C(g), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NO2        o0024(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  NO3        o0025(.A(ori_ori_n53_), .B(ori_ori_n48_), .C(ori_ori_n43_), .Y(ori_ori_n54_));
  AOI210     o0026(.A0(ori_ori_n54_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n55_));
  INV        o0027(.A(c), .Y(ori_ori_n56_));
  NA2        o0028(.A(e), .B(b), .Y(ori_ori_n57_));
  NO2        o0029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0030(.A(d), .Y(ori_ori_n59_));
  NAi21      o0031(.An(i), .B(h), .Y(ori_ori_n60_));
  NAi31      o0032(.An(i), .B(l), .C(j), .Y(ori_ori_n61_));
  NAi41      o0033(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n62_));
  NA2        o0034(.A(g), .B(f), .Y(ori_ori_n63_));
  NAi21      o0035(.An(i), .B(j), .Y(ori_ori_n64_));
  NAi32      o0036(.An(n), .Bn(k), .C(m), .Y(ori_ori_n65_));
  NAi31      o0037(.An(l), .B(m), .C(k), .Y(ori_ori_n66_));
  NAi21      o0038(.An(e), .B(h), .Y(ori_ori_n67_));
  NAi41      o0039(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n68_));
  INV        o0040(.A(m), .Y(ori_ori_n69_));
  NOi21      o0041(.An(k), .B(l), .Y(ori_ori_n70_));
  NA2        o0042(.A(ori_ori_n70_), .B(ori_ori_n69_), .Y(ori_ori_n71_));
  AN4        o0043(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n72_));
  NOi31      o0044(.An(h), .B(g), .C(f), .Y(ori_ori_n73_));
  NA2        o0045(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NAi32      o0046(.An(m), .Bn(k), .C(j), .Y(ori_ori_n75_));
  NOi32      o0047(.An(h), .Bn(g), .C(f), .Y(ori_ori_n76_));
  NA2        o0048(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  OA220      o0049(.A0(ori_ori_n77_), .A1(ori_ori_n75_), .B0(ori_ori_n74_), .B1(ori_ori_n71_), .Y(ori_ori_n78_));
  INV        o0050(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  INV        o0051(.A(n), .Y(ori_ori_n80_));
  NOi32      o0052(.An(e), .Bn(b), .C(d), .Y(ori_ori_n81_));
  NA2        o0053(.A(ori_ori_n81_), .B(ori_ori_n80_), .Y(ori_ori_n82_));
  INV        o0054(.A(j), .Y(ori_ori_n83_));
  AN3        o0055(.A(m), .B(k), .C(i), .Y(ori_ori_n84_));
  NA3        o0056(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(g), .Y(ori_ori_n85_));
  NO2        o0057(.A(ori_ori_n85_), .B(f), .Y(ori_ori_n86_));
  NAi32      o0058(.An(g), .Bn(f), .C(h), .Y(ori_ori_n87_));
  NAi31      o0059(.An(j), .B(m), .C(l), .Y(ori_ori_n88_));
  NO2        o0060(.A(ori_ori_n88_), .B(ori_ori_n87_), .Y(ori_ori_n89_));
  NA2        o0061(.A(m), .B(l), .Y(ori_ori_n90_));
  NAi31      o0062(.An(k), .B(j), .C(g), .Y(ori_ori_n91_));
  NO3        o0063(.A(ori_ori_n91_), .B(ori_ori_n90_), .C(f), .Y(ori_ori_n92_));
  AN2        o0064(.A(j), .B(g), .Y(ori_ori_n93_));
  NOi32      o0065(.An(m), .Bn(l), .C(i), .Y(ori_ori_n94_));
  NOi21      o0066(.An(g), .B(i), .Y(ori_ori_n95_));
  NOi32      o0067(.An(m), .Bn(j), .C(k), .Y(ori_ori_n96_));
  AOI220     o0068(.A0(ori_ori_n96_), .A1(ori_ori_n95_), .B0(ori_ori_n94_), .B1(ori_ori_n93_), .Y(ori_ori_n97_));
  NO2        o0069(.A(ori_ori_n97_), .B(f), .Y(ori_ori_n98_));
  NO4        o0070(.A(ori_ori_n98_), .B(ori_ori_n92_), .C(ori_ori_n89_), .D(ori_ori_n86_), .Y(ori_ori_n99_));
  NAi41      o0071(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n100_));
  AN2        o0072(.A(e), .B(b), .Y(ori_ori_n101_));
  NOi31      o0073(.An(c), .B(h), .C(f), .Y(ori_ori_n102_));
  NA2        o0074(.A(ori_ori_n102_), .B(ori_ori_n101_), .Y(ori_ori_n103_));
  NO2        o0075(.A(ori_ori_n103_), .B(ori_ori_n100_), .Y(ori_ori_n104_));
  NOi21      o0076(.An(g), .B(f), .Y(ori_ori_n105_));
  NOi21      o0077(.An(i), .B(h), .Y(ori_ori_n106_));
  NA3        o0078(.A(ori_ori_n106_), .B(ori_ori_n105_), .C(ori_ori_n36_), .Y(ori_ori_n107_));
  INV        o0079(.A(a), .Y(ori_ori_n108_));
  NA2        o0080(.A(ori_ori_n101_), .B(ori_ori_n108_), .Y(ori_ori_n109_));
  INV        o0081(.A(l), .Y(ori_ori_n110_));
  NOi21      o0082(.An(m), .B(n), .Y(ori_ori_n111_));
  AN2        o0083(.A(k), .B(h), .Y(ori_ori_n112_));
  NO2        o0084(.A(ori_ori_n107_), .B(ori_ori_n82_), .Y(ori_ori_n113_));
  INV        o0085(.A(b), .Y(ori_ori_n114_));
  NA2        o0086(.A(l), .B(j), .Y(ori_ori_n115_));
  AN2        o0087(.A(k), .B(i), .Y(ori_ori_n116_));
  NA2        o0088(.A(ori_ori_n116_), .B(ori_ori_n115_), .Y(ori_ori_n117_));
  NA2        o0089(.A(g), .B(e), .Y(ori_ori_n118_));
  NOi32      o0090(.An(c), .Bn(a), .C(d), .Y(ori_ori_n119_));
  NA2        o0091(.A(ori_ori_n119_), .B(ori_ori_n111_), .Y(ori_ori_n120_));
  NO2        o0092(.A(ori_ori_n113_), .B(ori_ori_n104_), .Y(ori_ori_n121_));
  OAI210     o0093(.A0(ori_ori_n99_), .A1(ori_ori_n82_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  NOi31      o0094(.An(k), .B(m), .C(j), .Y(ori_ori_n123_));
  NA3        o0095(.A(ori_ori_n123_), .B(ori_ori_n73_), .C(ori_ori_n72_), .Y(ori_ori_n124_));
  NOi31      o0096(.An(k), .B(m), .C(i), .Y(ori_ori_n125_));
  INV        o0097(.A(ori_ori_n124_), .Y(ori_ori_n126_));
  NOi32      o0098(.An(f), .Bn(b), .C(e), .Y(ori_ori_n127_));
  NAi21      o0099(.An(g), .B(h), .Y(ori_ori_n128_));
  NAi21      o0100(.An(m), .B(n), .Y(ori_ori_n129_));
  NAi21      o0101(.An(j), .B(k), .Y(ori_ori_n130_));
  NO3        o0102(.A(ori_ori_n130_), .B(ori_ori_n129_), .C(ori_ori_n128_), .Y(ori_ori_n131_));
  NAi41      o0103(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n132_));
  NAi31      o0104(.An(j), .B(k), .C(h), .Y(ori_ori_n133_));
  NA2        o0105(.A(ori_ori_n131_), .B(ori_ori_n127_), .Y(ori_ori_n134_));
  NO2        o0106(.A(k), .B(j), .Y(ori_ori_n135_));
  NO2        o0107(.A(ori_ori_n135_), .B(ori_ori_n129_), .Y(ori_ori_n136_));
  AN2        o0108(.A(k), .B(j), .Y(ori_ori_n137_));
  NAi21      o0109(.An(c), .B(b), .Y(ori_ori_n138_));
  NA2        o0110(.A(f), .B(d), .Y(ori_ori_n139_));
  NO4        o0111(.A(ori_ori_n139_), .B(ori_ori_n138_), .C(ori_ori_n137_), .D(ori_ori_n128_), .Y(ori_ori_n140_));
  NA2        o0112(.A(h), .B(c), .Y(ori_ori_n141_));
  NAi31      o0113(.An(f), .B(e), .C(b), .Y(ori_ori_n142_));
  NA2        o0114(.A(ori_ori_n140_), .B(ori_ori_n136_), .Y(ori_ori_n143_));
  NA2        o0115(.A(d), .B(b), .Y(ori_ori_n144_));
  NAi21      o0116(.An(e), .B(f), .Y(ori_ori_n145_));
  NO2        o0117(.A(ori_ori_n145_), .B(ori_ori_n144_), .Y(ori_ori_n146_));
  NA2        o0118(.A(b), .B(a), .Y(ori_ori_n147_));
  NAi21      o0119(.An(e), .B(g), .Y(ori_ori_n148_));
  NAi21      o0120(.An(c), .B(d), .Y(ori_ori_n149_));
  NAi31      o0121(.An(l), .B(k), .C(h), .Y(ori_ori_n150_));
  NO2        o0122(.A(ori_ori_n129_), .B(ori_ori_n150_), .Y(ori_ori_n151_));
  NA2        o0123(.A(ori_ori_n151_), .B(ori_ori_n146_), .Y(ori_ori_n152_));
  NAi41      o0124(.An(ori_ori_n126_), .B(ori_ori_n152_), .C(ori_ori_n143_), .D(ori_ori_n134_), .Y(ori_ori_n153_));
  NAi31      o0125(.An(e), .B(f), .C(b), .Y(ori_ori_n154_));
  NOi21      o0126(.An(g), .B(d), .Y(ori_ori_n155_));
  NO2        o0127(.A(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NOi21      o0128(.An(h), .B(i), .Y(ori_ori_n157_));
  NOi21      o0129(.An(k), .B(m), .Y(ori_ori_n158_));
  NA3        o0130(.A(ori_ori_n158_), .B(ori_ori_n157_), .C(n), .Y(ori_ori_n159_));
  NOi21      o0131(.An(ori_ori_n156_), .B(ori_ori_n159_), .Y(ori_ori_n160_));
  NOi21      o0132(.An(h), .B(g), .Y(ori_ori_n161_));
  NAi31      o0133(.An(l), .B(j), .C(h), .Y(ori_ori_n162_));
  NOi32      o0134(.An(n), .Bn(k), .C(m), .Y(ori_ori_n163_));
  NA2        o0135(.A(l), .B(i), .Y(ori_ori_n164_));
  NAi31      o0136(.An(d), .B(f), .C(c), .Y(ori_ori_n165_));
  NAi31      o0137(.An(e), .B(f), .C(c), .Y(ori_ori_n166_));
  NA2        o0138(.A(ori_ori_n166_), .B(ori_ori_n165_), .Y(ori_ori_n167_));
  NA2        o0139(.A(j), .B(h), .Y(ori_ori_n168_));
  OR3        o0140(.A(n), .B(m), .C(k), .Y(ori_ori_n169_));
  NO2        o0141(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  NAi32      o0142(.An(m), .Bn(k), .C(n), .Y(ori_ori_n171_));
  NO2        o0143(.A(ori_ori_n171_), .B(ori_ori_n168_), .Y(ori_ori_n172_));
  AOI220     o0144(.A0(ori_ori_n172_), .A1(ori_ori_n156_), .B0(ori_ori_n170_), .B1(ori_ori_n167_), .Y(ori_ori_n173_));
  NO2        o0145(.A(n), .B(m), .Y(ori_ori_n174_));
  NA2        o0146(.A(ori_ori_n174_), .B(ori_ori_n50_), .Y(ori_ori_n175_));
  NAi21      o0147(.An(f), .B(e), .Y(ori_ori_n176_));
  NA2        o0148(.A(d), .B(c), .Y(ori_ori_n177_));
  NO2        o0149(.A(ori_ori_n177_), .B(ori_ori_n176_), .Y(ori_ori_n178_));
  NOi21      o0150(.An(ori_ori_n178_), .B(ori_ori_n175_), .Y(ori_ori_n179_));
  NAi31      o0151(.An(m), .B(n), .C(b), .Y(ori_ori_n180_));
  NA2        o0152(.A(k), .B(i), .Y(ori_ori_n181_));
  NAi21      o0153(.An(h), .B(f), .Y(ori_ori_n182_));
  NO2        o0154(.A(ori_ori_n182_), .B(ori_ori_n181_), .Y(ori_ori_n183_));
  NO2        o0155(.A(ori_ori_n180_), .B(ori_ori_n149_), .Y(ori_ori_n184_));
  NA2        o0156(.A(ori_ori_n184_), .B(ori_ori_n183_), .Y(ori_ori_n185_));
  NOi32      o0157(.An(f), .Bn(c), .C(d), .Y(ori_ori_n186_));
  NOi32      o0158(.An(f), .Bn(c), .C(e), .Y(ori_ori_n187_));
  NO2        o0159(.A(ori_ori_n187_), .B(ori_ori_n186_), .Y(ori_ori_n188_));
  NO3        o0160(.A(n), .B(m), .C(j), .Y(ori_ori_n189_));
  NA2        o0161(.A(ori_ori_n189_), .B(ori_ori_n112_), .Y(ori_ori_n190_));
  AO210      o0162(.A0(ori_ori_n190_), .A1(ori_ori_n175_), .B0(ori_ori_n188_), .Y(ori_ori_n191_));
  NAi41      o0163(.An(ori_ori_n179_), .B(ori_ori_n191_), .C(ori_ori_n185_), .D(ori_ori_n173_), .Y(ori_ori_n192_));
  OR3        o0164(.A(ori_ori_n192_), .B(ori_ori_n160_), .C(ori_ori_n153_), .Y(ori_ori_n193_));
  NO4        o0165(.A(ori_ori_n193_), .B(ori_ori_n122_), .C(ori_ori_n79_), .D(ori_ori_n55_), .Y(ori_ori_n194_));
  NA3        o0166(.A(m), .B(ori_ori_n110_), .C(j), .Y(ori_ori_n195_));
  NAi31      o0167(.An(n), .B(h), .C(g), .Y(ori_ori_n196_));
  NO2        o0168(.A(ori_ori_n196_), .B(ori_ori_n195_), .Y(ori_ori_n197_));
  NOi32      o0169(.An(m), .Bn(k), .C(l), .Y(ori_ori_n198_));
  NA3        o0170(.A(ori_ori_n198_), .B(ori_ori_n83_), .C(g), .Y(ori_ori_n199_));
  NO2        o0171(.A(ori_ori_n199_), .B(n), .Y(ori_ori_n200_));
  NOi21      o0172(.An(k), .B(j), .Y(ori_ori_n201_));
  NA4        o0173(.A(ori_ori_n201_), .B(ori_ori_n111_), .C(i), .D(g), .Y(ori_ori_n202_));
  AN2        o0174(.A(i), .B(g), .Y(ori_ori_n203_));
  NA3        o0175(.A(ori_ori_n70_), .B(ori_ori_n203_), .C(ori_ori_n111_), .Y(ori_ori_n204_));
  NA2        o0176(.A(ori_ori_n204_), .B(ori_ori_n202_), .Y(ori_ori_n205_));
  NO3        o0177(.A(ori_ori_n205_), .B(ori_ori_n200_), .C(ori_ori_n197_), .Y(ori_ori_n206_));
  NAi41      o0178(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n207_));
  INV        o0179(.A(ori_ori_n207_), .Y(ori_ori_n208_));
  INV        o0180(.A(f), .Y(ori_ori_n209_));
  INV        o0181(.A(g), .Y(ori_ori_n210_));
  NOi31      o0182(.An(i), .B(j), .C(h), .Y(ori_ori_n211_));
  NOi21      o0183(.An(l), .B(m), .Y(ori_ori_n212_));
  NA2        o0184(.A(ori_ori_n212_), .B(ori_ori_n211_), .Y(ori_ori_n213_));
  NO3        o0185(.A(ori_ori_n213_), .B(ori_ori_n210_), .C(ori_ori_n209_), .Y(ori_ori_n214_));
  NA2        o0186(.A(ori_ori_n214_), .B(ori_ori_n208_), .Y(ori_ori_n215_));
  OAI210     o0187(.A0(ori_ori_n206_), .A1(ori_ori_n32_), .B0(ori_ori_n215_), .Y(ori_ori_n216_));
  NOi21      o0188(.An(n), .B(m), .Y(ori_ori_n217_));
  NOi32      o0189(.An(l), .Bn(i), .C(j), .Y(ori_ori_n218_));
  NA2        o0190(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n219_));
  OA220      o0191(.A0(ori_ori_n219_), .A1(ori_ori_n103_), .B0(ori_ori_n75_), .B1(ori_ori_n74_), .Y(ori_ori_n220_));
  NAi21      o0192(.An(j), .B(h), .Y(ori_ori_n221_));
  XN2        o0193(.A(i), .B(h), .Y(ori_ori_n222_));
  NA2        o0194(.A(ori_ori_n222_), .B(ori_ori_n221_), .Y(ori_ori_n223_));
  NOi31      o0195(.An(k), .B(n), .C(m), .Y(ori_ori_n224_));
  NOi31      o0196(.An(ori_ori_n224_), .B(ori_ori_n177_), .C(ori_ori_n176_), .Y(ori_ori_n225_));
  NA2        o0197(.A(ori_ori_n225_), .B(ori_ori_n223_), .Y(ori_ori_n226_));
  NAi31      o0198(.An(f), .B(e), .C(c), .Y(ori_ori_n227_));
  NO4        o0199(.A(ori_ori_n227_), .B(ori_ori_n169_), .C(ori_ori_n168_), .D(ori_ori_n59_), .Y(ori_ori_n228_));
  NA3        o0200(.A(e), .B(c), .C(b), .Y(ori_ori_n229_));
  NAi32      o0201(.An(m), .Bn(i), .C(k), .Y(ori_ori_n230_));
  INV        o0202(.A(k), .Y(ori_ori_n231_));
  INV        o0203(.A(ori_ori_n228_), .Y(ori_ori_n232_));
  NAi21      o0204(.An(n), .B(a), .Y(ori_ori_n233_));
  NO2        o0205(.A(ori_ori_n233_), .B(ori_ori_n144_), .Y(ori_ori_n234_));
  NAi41      o0206(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n235_));
  NO2        o0207(.A(ori_ori_n235_), .B(e), .Y(ori_ori_n236_));
  NA2        o0208(.A(ori_ori_n236_), .B(ori_ori_n234_), .Y(ori_ori_n237_));
  AN4        o0209(.A(ori_ori_n237_), .B(ori_ori_n232_), .C(ori_ori_n226_), .D(ori_ori_n220_), .Y(ori_ori_n238_));
  OR2        o0210(.A(h), .B(g), .Y(ori_ori_n239_));
  NO2        o0211(.A(ori_ori_n239_), .B(ori_ori_n100_), .Y(ori_ori_n240_));
  NA2        o0212(.A(ori_ori_n240_), .B(ori_ori_n127_), .Y(ori_ori_n241_));
  NAi41      o0213(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n242_));
  NO2        o0214(.A(ori_ori_n242_), .B(ori_ori_n209_), .Y(ori_ori_n243_));
  NA2        o0215(.A(ori_ori_n158_), .B(ori_ori_n106_), .Y(ori_ori_n244_));
  NAi21      o0216(.An(ori_ori_n244_), .B(ori_ori_n243_), .Y(ori_ori_n245_));
  NO2        o0217(.A(n), .B(a), .Y(ori_ori_n246_));
  NAi31      o0218(.An(ori_ori_n235_), .B(ori_ori_n246_), .C(ori_ori_n101_), .Y(ori_ori_n247_));
  AN2        o0219(.A(ori_ori_n247_), .B(ori_ori_n245_), .Y(ori_ori_n248_));
  NAi21      o0220(.An(h), .B(i), .Y(ori_ori_n249_));
  NA2        o0221(.A(ori_ori_n174_), .B(k), .Y(ori_ori_n250_));
  NO2        o0222(.A(ori_ori_n250_), .B(ori_ori_n249_), .Y(ori_ori_n251_));
  NA2        o0223(.A(ori_ori_n251_), .B(ori_ori_n186_), .Y(ori_ori_n252_));
  NA3        o0224(.A(ori_ori_n252_), .B(ori_ori_n248_), .C(ori_ori_n241_), .Y(ori_ori_n253_));
  NOi21      o0225(.An(g), .B(e), .Y(ori_ori_n254_));
  NO2        o0226(.A(ori_ori_n68_), .B(ori_ori_n69_), .Y(ori_ori_n255_));
  NA2        o0227(.A(ori_ori_n255_), .B(ori_ori_n254_), .Y(ori_ori_n256_));
  NOi32      o0228(.An(l), .Bn(j), .C(i), .Y(ori_ori_n257_));
  AOI210     o0229(.A0(ori_ori_n70_), .A1(ori_ori_n83_), .B0(ori_ori_n257_), .Y(ori_ori_n258_));
  NAi21      o0230(.An(f), .B(g), .Y(ori_ori_n259_));
  NO2        o0231(.A(ori_ori_n259_), .B(ori_ori_n62_), .Y(ori_ori_n260_));
  NO2        o0232(.A(ori_ori_n65_), .B(ori_ori_n115_), .Y(ori_ori_n261_));
  NO2        o0233(.A(ori_ori_n258_), .B(ori_ori_n256_), .Y(ori_ori_n262_));
  NOi41      o0234(.An(ori_ori_n238_), .B(ori_ori_n262_), .C(ori_ori_n253_), .D(ori_ori_n216_), .Y(ori_ori_n263_));
  NO4        o0235(.A(ori_ori_n197_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n264_));
  NO2        o0236(.A(ori_ori_n264_), .B(ori_ori_n109_), .Y(ori_ori_n265_));
  NA3        o0237(.A(ori_ori_n59_), .B(c), .C(b), .Y(ori_ori_n266_));
  NAi21      o0238(.An(h), .B(g), .Y(ori_ori_n267_));
  NO2        o0239(.A(ori_ori_n244_), .B(ori_ori_n259_), .Y(ori_ori_n268_));
  NAi31      o0240(.An(g), .B(k), .C(h), .Y(ori_ori_n269_));
  NA4        o0241(.A(ori_ori_n158_), .B(ori_ori_n76_), .C(ori_ori_n72_), .D(ori_ori_n115_), .Y(ori_ori_n270_));
  NA3        o0242(.A(ori_ori_n158_), .B(ori_ori_n157_), .C(ori_ori_n80_), .Y(ori_ori_n271_));
  NO2        o0243(.A(ori_ori_n271_), .B(ori_ori_n188_), .Y(ori_ori_n272_));
  NOi21      o0244(.An(ori_ori_n270_), .B(ori_ori_n272_), .Y(ori_ori_n273_));
  NA3        o0245(.A(e), .B(c), .C(b), .Y(ori_ori_n274_));
  NAi32      o0246(.An(k), .Bn(i), .C(j), .Y(ori_ori_n275_));
  NAi31      o0247(.An(h), .B(l), .C(i), .Y(ori_ori_n276_));
  NA3        o0248(.A(ori_ori_n276_), .B(ori_ori_n275_), .C(ori_ori_n162_), .Y(ori_ori_n277_));
  NOi21      o0249(.An(ori_ori_n277_), .B(ori_ori_n49_), .Y(ori_ori_n278_));
  NA2        o0250(.A(ori_ori_n260_), .B(ori_ori_n278_), .Y(ori_ori_n279_));
  NAi21      o0251(.An(l), .B(k), .Y(ori_ori_n280_));
  NO2        o0252(.A(ori_ori_n280_), .B(ori_ori_n49_), .Y(ori_ori_n281_));
  NOi21      o0253(.An(l), .B(j), .Y(ori_ori_n282_));
  NA2        o0254(.A(ori_ori_n161_), .B(ori_ori_n282_), .Y(ori_ori_n283_));
  NA3        o0255(.A(ori_ori_n116_), .B(ori_ori_n115_), .C(g), .Y(ori_ori_n284_));
  OR3        o0256(.A(ori_ori_n68_), .B(ori_ori_n69_), .C(e), .Y(ori_ori_n285_));
  AOI210     o0257(.A0(ori_ori_n284_), .A1(ori_ori_n283_), .B0(ori_ori_n285_), .Y(ori_ori_n286_));
  INV        o0258(.A(ori_ori_n286_), .Y(ori_ori_n287_));
  NAi32      o0259(.An(j), .Bn(h), .C(i), .Y(ori_ori_n288_));
  NAi21      o0260(.An(m), .B(l), .Y(ori_ori_n289_));
  NO3        o0261(.A(ori_ori_n289_), .B(ori_ori_n288_), .C(ori_ori_n80_), .Y(ori_ori_n290_));
  NA2        o0262(.A(h), .B(g), .Y(ori_ori_n291_));
  NA3        o0263(.A(ori_ori_n287_), .B(ori_ori_n279_), .C(ori_ori_n273_), .Y(ori_ori_n292_));
  NO2        o0264(.A(ori_ori_n142_), .B(d), .Y(ori_ori_n293_));
  NA2        o0265(.A(ori_ori_n293_), .B(ori_ori_n53_), .Y(ori_ori_n294_));
  NO2        o0266(.A(ori_ori_n103_), .B(ori_ori_n100_), .Y(ori_ori_n295_));
  NAi32      o0267(.An(n), .Bn(m), .C(l), .Y(ori_ori_n296_));
  NO2        o0268(.A(ori_ori_n296_), .B(ori_ori_n288_), .Y(ori_ori_n297_));
  NA2        o0269(.A(ori_ori_n297_), .B(ori_ori_n178_), .Y(ori_ori_n298_));
  NAi31      o0270(.An(k), .B(l), .C(j), .Y(ori_ori_n299_));
  OAI210     o0271(.A0(ori_ori_n280_), .A1(j), .B0(ori_ori_n299_), .Y(ori_ori_n300_));
  NOi21      o0272(.An(ori_ori_n300_), .B(ori_ori_n118_), .Y(ori_ori_n301_));
  NA2        o0273(.A(ori_ori_n298_), .B(ori_ori_n294_), .Y(ori_ori_n302_));
  NO3        o0274(.A(ori_ori_n302_), .B(ori_ori_n292_), .C(ori_ori_n265_), .Y(ori_ori_n303_));
  NA2        o0275(.A(ori_ori_n251_), .B(ori_ori_n187_), .Y(ori_ori_n304_));
  NAi21      o0276(.An(m), .B(k), .Y(ori_ori_n305_));
  NO2        o0277(.A(ori_ori_n222_), .B(ori_ori_n305_), .Y(ori_ori_n306_));
  NAi41      o0278(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n307_));
  NO2        o0279(.A(ori_ori_n307_), .B(ori_ori_n148_), .Y(ori_ori_n308_));
  NA2        o0280(.A(ori_ori_n308_), .B(ori_ori_n306_), .Y(ori_ori_n309_));
  NAi31      o0281(.An(i), .B(l), .C(h), .Y(ori_ori_n310_));
  NA2        o0282(.A(e), .B(c), .Y(ori_ori_n311_));
  NO3        o0283(.A(ori_ori_n311_), .B(n), .C(d), .Y(ori_ori_n312_));
  NOi21      o0284(.An(f), .B(h), .Y(ori_ori_n313_));
  NA2        o0285(.A(ori_ori_n313_), .B(ori_ori_n116_), .Y(ori_ori_n314_));
  NO2        o0286(.A(ori_ori_n314_), .B(ori_ori_n210_), .Y(ori_ori_n315_));
  NAi31      o0287(.An(d), .B(e), .C(b), .Y(ori_ori_n316_));
  NO2        o0288(.A(ori_ori_n129_), .B(ori_ori_n316_), .Y(ori_ori_n317_));
  NA2        o0289(.A(ori_ori_n317_), .B(ori_ori_n315_), .Y(ori_ori_n318_));
  NA3        o0290(.A(ori_ori_n318_), .B(ori_ori_n309_), .C(ori_ori_n304_), .Y(ori_ori_n319_));
  NO4        o0291(.A(ori_ori_n307_), .B(ori_ori_n75_), .C(ori_ori_n67_), .D(ori_ori_n210_), .Y(ori_ori_n320_));
  NA2        o0292(.A(ori_ori_n246_), .B(ori_ori_n101_), .Y(ori_ori_n321_));
  OR2        o0293(.A(ori_ori_n321_), .B(ori_ori_n199_), .Y(ori_ori_n322_));
  NOi31      o0294(.An(l), .B(n), .C(m), .Y(ori_ori_n323_));
  NA2        o0295(.A(ori_ori_n323_), .B(ori_ori_n211_), .Y(ori_ori_n324_));
  NO2        o0296(.A(ori_ori_n324_), .B(ori_ori_n188_), .Y(ori_ori_n325_));
  NAi32      o0297(.An(ori_ori_n325_), .Bn(ori_ori_n320_), .C(ori_ori_n322_), .Y(ori_ori_n326_));
  NAi32      o0298(.An(m), .Bn(j), .C(k), .Y(ori_ori_n327_));
  NAi41      o0299(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n328_));
  OAI210     o0300(.A0(ori_ori_n207_), .A1(ori_ori_n327_), .B0(ori_ori_n328_), .Y(ori_ori_n329_));
  NOi31      o0301(.An(j), .B(m), .C(k), .Y(ori_ori_n330_));
  NO2        o0302(.A(ori_ori_n123_), .B(ori_ori_n330_), .Y(ori_ori_n331_));
  AN3        o0303(.A(h), .B(g), .C(f), .Y(ori_ori_n332_));
  NAi31      o0304(.An(ori_ori_n331_), .B(ori_ori_n332_), .C(ori_ori_n329_), .Y(ori_ori_n333_));
  NOi32      o0305(.An(m), .Bn(j), .C(l), .Y(ori_ori_n334_));
  NO2        o0306(.A(ori_ori_n334_), .B(ori_ori_n94_), .Y(ori_ori_n335_));
  NAi32      o0307(.An(ori_ori_n335_), .Bn(ori_ori_n196_), .C(ori_ori_n293_), .Y(ori_ori_n336_));
  NO2        o0308(.A(ori_ori_n289_), .B(ori_ori_n288_), .Y(ori_ori_n337_));
  NO2        o0309(.A(ori_ori_n213_), .B(g), .Y(ori_ori_n338_));
  NO2        o0310(.A(ori_ori_n154_), .B(ori_ori_n80_), .Y(ori_ori_n339_));
  AOI220     o0311(.A0(ori_ori_n339_), .A1(ori_ori_n338_), .B0(ori_ori_n243_), .B1(ori_ori_n337_), .Y(ori_ori_n340_));
  NA2        o0312(.A(ori_ori_n230_), .B(ori_ori_n75_), .Y(ori_ori_n341_));
  NA3        o0313(.A(ori_ori_n341_), .B(ori_ori_n332_), .C(ori_ori_n208_), .Y(ori_ori_n342_));
  NA4        o0314(.A(ori_ori_n342_), .B(ori_ori_n340_), .C(ori_ori_n336_), .D(ori_ori_n333_), .Y(ori_ori_n343_));
  NA3        o0315(.A(h), .B(g), .C(f), .Y(ori_ori_n344_));
  NO2        o0316(.A(ori_ori_n344_), .B(ori_ori_n71_), .Y(ori_ori_n345_));
  NA2        o0317(.A(ori_ori_n328_), .B(ori_ori_n207_), .Y(ori_ori_n346_));
  NA2        o0318(.A(ori_ori_n161_), .B(e), .Y(ori_ori_n347_));
  NO2        o0319(.A(ori_ori_n347_), .B(ori_ori_n41_), .Y(ori_ori_n348_));
  NA2        o0320(.A(ori_ori_n346_), .B(ori_ori_n345_), .Y(ori_ori_n349_));
  NOi32      o0321(.An(j), .Bn(g), .C(i), .Y(ori_ori_n350_));
  NA3        o0322(.A(ori_ori_n350_), .B(ori_ori_n280_), .C(ori_ori_n111_), .Y(ori_ori_n351_));
  AO210      o0323(.A0(ori_ori_n109_), .A1(ori_ori_n32_), .B0(ori_ori_n351_), .Y(ori_ori_n352_));
  NOi32      o0324(.An(e), .Bn(b), .C(a), .Y(ori_ori_n353_));
  AN2        o0325(.A(l), .B(j), .Y(ori_ori_n354_));
  NO2        o0326(.A(ori_ori_n305_), .B(ori_ori_n354_), .Y(ori_ori_n355_));
  NO3        o0327(.A(ori_ori_n307_), .B(ori_ori_n67_), .C(ori_ori_n210_), .Y(ori_ori_n356_));
  NA3        o0328(.A(ori_ori_n204_), .B(ori_ori_n202_), .C(ori_ori_n35_), .Y(ori_ori_n357_));
  AOI220     o0329(.A0(ori_ori_n357_), .A1(ori_ori_n353_), .B0(ori_ori_n356_), .B1(ori_ori_n355_), .Y(ori_ori_n358_));
  NO2        o0330(.A(ori_ori_n316_), .B(n), .Y(ori_ori_n359_));
  NA2        o0331(.A(ori_ori_n203_), .B(k), .Y(ori_ori_n360_));
  NA3        o0332(.A(m), .B(ori_ori_n110_), .C(ori_ori_n209_), .Y(ori_ori_n361_));
  NA4        o0333(.A(ori_ori_n198_), .B(ori_ori_n83_), .C(g), .D(ori_ori_n209_), .Y(ori_ori_n362_));
  OAI210     o0334(.A0(ori_ori_n361_), .A1(ori_ori_n360_), .B0(ori_ori_n362_), .Y(ori_ori_n363_));
  NA2        o0335(.A(ori_ori_n51_), .B(ori_ori_n111_), .Y(ori_ori_n364_));
  NA2        o0336(.A(ori_ori_n363_), .B(ori_ori_n359_), .Y(ori_ori_n365_));
  NA4        o0337(.A(ori_ori_n365_), .B(ori_ori_n358_), .C(ori_ori_n352_), .D(ori_ori_n349_), .Y(ori_ori_n366_));
  NO4        o0338(.A(ori_ori_n366_), .B(ori_ori_n343_), .C(ori_ori_n326_), .D(ori_ori_n319_), .Y(ori_ori_n367_));
  NA4        o0339(.A(ori_ori_n367_), .B(ori_ori_n303_), .C(ori_ori_n263_), .D(ori_ori_n194_), .Y(ori10));
  NA3        o0340(.A(m), .B(k), .C(i), .Y(ori_ori_n369_));
  NO3        o0341(.A(ori_ori_n369_), .B(j), .C(ori_ori_n210_), .Y(ori_ori_n370_));
  NOi21      o0342(.An(e), .B(f), .Y(ori_ori_n371_));
  NO4        o0343(.A(ori_ori_n149_), .B(ori_ori_n371_), .C(n), .D(ori_ori_n108_), .Y(ori_ori_n372_));
  NAi31      o0344(.An(b), .B(f), .C(c), .Y(ori_ori_n373_));
  INV        o0345(.A(ori_ori_n373_), .Y(ori_ori_n374_));
  NOi32      o0346(.An(k), .Bn(h), .C(j), .Y(ori_ori_n375_));
  NA2        o0347(.A(ori_ori_n375_), .B(ori_ori_n217_), .Y(ori_ori_n376_));
  NA2        o0348(.A(ori_ori_n159_), .B(ori_ori_n376_), .Y(ori_ori_n377_));
  AOI220     o0349(.A0(ori_ori_n377_), .A1(ori_ori_n374_), .B0(ori_ori_n372_), .B1(ori_ori_n370_), .Y(ori_ori_n378_));
  AN2        o0350(.A(j), .B(h), .Y(ori_ori_n379_));
  NO3        o0351(.A(n), .B(m), .C(k), .Y(ori_ori_n380_));
  NA2        o0352(.A(ori_ori_n380_), .B(ori_ori_n379_), .Y(ori_ori_n381_));
  NO3        o0353(.A(ori_ori_n381_), .B(ori_ori_n149_), .C(ori_ori_n209_), .Y(ori_ori_n382_));
  OR2        o0354(.A(m), .B(k), .Y(ori_ori_n383_));
  NO2        o0355(.A(ori_ori_n168_), .B(ori_ori_n383_), .Y(ori_ori_n384_));
  NA4        o0356(.A(n), .B(f), .C(c), .D(ori_ori_n114_), .Y(ori_ori_n385_));
  NOi21      o0357(.An(ori_ori_n384_), .B(ori_ori_n385_), .Y(ori_ori_n386_));
  NOi32      o0358(.An(d), .Bn(a), .C(c), .Y(ori_ori_n387_));
  NA2        o0359(.A(ori_ori_n387_), .B(ori_ori_n176_), .Y(ori_ori_n388_));
  NAi21      o0360(.An(i), .B(g), .Y(ori_ori_n389_));
  NAi31      o0361(.An(k), .B(m), .C(j), .Y(ori_ori_n390_));
  NO3        o0362(.A(ori_ori_n390_), .B(ori_ori_n389_), .C(n), .Y(ori_ori_n391_));
  NOi21      o0363(.An(ori_ori_n391_), .B(ori_ori_n388_), .Y(ori_ori_n392_));
  NO3        o0364(.A(ori_ori_n392_), .B(ori_ori_n386_), .C(ori_ori_n382_), .Y(ori_ori_n393_));
  NO2        o0365(.A(ori_ori_n385_), .B(ori_ori_n289_), .Y(ori_ori_n394_));
  NOi32      o0366(.An(f), .Bn(d), .C(c), .Y(ori_ori_n395_));
  AOI220     o0367(.A0(ori_ori_n395_), .A1(ori_ori_n297_), .B0(ori_ori_n394_), .B1(ori_ori_n211_), .Y(ori_ori_n396_));
  NA3        o0368(.A(ori_ori_n396_), .B(ori_ori_n393_), .C(ori_ori_n378_), .Y(ori_ori_n397_));
  NO2        o0369(.A(ori_ori_n59_), .B(ori_ori_n114_), .Y(ori_ori_n398_));
  NA2        o0370(.A(ori_ori_n246_), .B(ori_ori_n398_), .Y(ori_ori_n399_));
  INV        o0371(.A(e), .Y(ori_ori_n400_));
  NA2        o0372(.A(ori_ori_n46_), .B(e), .Y(ori_ori_n401_));
  OAI220     o0373(.A0(ori_ori_n401_), .A1(ori_ori_n195_), .B0(ori_ori_n199_), .B1(ori_ori_n400_), .Y(ori_ori_n402_));
  AN2        o0374(.A(g), .B(e), .Y(ori_ori_n403_));
  NA3        o0375(.A(ori_ori_n403_), .B(ori_ori_n198_), .C(i), .Y(ori_ori_n404_));
  OAI210     o0376(.A0(ori_ori_n85_), .A1(ori_ori_n400_), .B0(ori_ori_n404_), .Y(ori_ori_n405_));
  NO2        o0377(.A(ori_ori_n97_), .B(ori_ori_n400_), .Y(ori_ori_n406_));
  NO3        o0378(.A(ori_ori_n406_), .B(ori_ori_n405_), .C(ori_ori_n402_), .Y(ori_ori_n407_));
  NOi32      o0379(.An(h), .Bn(e), .C(g), .Y(ori_ori_n408_));
  NA3        o0380(.A(ori_ori_n408_), .B(ori_ori_n282_), .C(m), .Y(ori_ori_n409_));
  NOi21      o0381(.An(g), .B(h), .Y(ori_ori_n410_));
  AN3        o0382(.A(m), .B(l), .C(i), .Y(ori_ori_n411_));
  NA3        o0383(.A(ori_ori_n411_), .B(ori_ori_n410_), .C(e), .Y(ori_ori_n412_));
  AN3        o0384(.A(h), .B(g), .C(e), .Y(ori_ori_n413_));
  NA2        o0385(.A(ori_ori_n413_), .B(ori_ori_n94_), .Y(ori_ori_n414_));
  AN3        o0386(.A(ori_ori_n414_), .B(ori_ori_n412_), .C(ori_ori_n409_), .Y(ori_ori_n415_));
  AOI210     o0387(.A0(ori_ori_n415_), .A1(ori_ori_n407_), .B0(ori_ori_n399_), .Y(ori_ori_n416_));
  NA3        o0388(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(e), .Y(ori_ori_n417_));
  NO2        o0389(.A(ori_ori_n417_), .B(ori_ori_n399_), .Y(ori_ori_n418_));
  NA3        o0390(.A(ori_ori_n387_), .B(ori_ori_n176_), .C(ori_ori_n80_), .Y(ori_ori_n419_));
  NAi31      o0391(.An(b), .B(c), .C(a), .Y(ori_ori_n420_));
  NO2        o0392(.A(ori_ori_n420_), .B(n), .Y(ori_ori_n421_));
  NA2        o0393(.A(ori_ori_n51_), .B(m), .Y(ori_ori_n422_));
  NO2        o0394(.A(ori_ori_n422_), .B(ori_ori_n145_), .Y(ori_ori_n423_));
  NA2        o0395(.A(ori_ori_n423_), .B(ori_ori_n421_), .Y(ori_ori_n424_));
  INV        o0396(.A(ori_ori_n424_), .Y(ori_ori_n425_));
  NO4        o0397(.A(ori_ori_n425_), .B(ori_ori_n418_), .C(ori_ori_n416_), .D(ori_ori_n397_), .Y(ori_ori_n426_));
  NA2        o0398(.A(i), .B(g), .Y(ori_ori_n427_));
  NOi21      o0399(.An(a), .B(n), .Y(ori_ori_n428_));
  NOi21      o0400(.An(d), .B(c), .Y(ori_ori_n429_));
  NA2        o0401(.A(ori_ori_n429_), .B(ori_ori_n428_), .Y(ori_ori_n430_));
  NA3        o0402(.A(i), .B(g), .C(f), .Y(ori_ori_n431_));
  OR2        o0403(.A(ori_ori_n431_), .B(ori_ori_n66_), .Y(ori_ori_n432_));
  NA3        o0404(.A(ori_ori_n411_), .B(ori_ori_n410_), .C(ori_ori_n176_), .Y(ori_ori_n433_));
  AOI210     o0405(.A0(ori_ori_n433_), .A1(ori_ori_n432_), .B0(ori_ori_n430_), .Y(ori_ori_n434_));
  INV        o0406(.A(ori_ori_n434_), .Y(ori_ori_n435_));
  OR2        o0407(.A(n), .B(m), .Y(ori_ori_n436_));
  NO2        o0408(.A(ori_ori_n436_), .B(ori_ori_n150_), .Y(ori_ori_n437_));
  NO2        o0409(.A(ori_ori_n177_), .B(ori_ori_n145_), .Y(ori_ori_n438_));
  OAI210     o0410(.A0(ori_ori_n437_), .A1(ori_ori_n170_), .B0(ori_ori_n438_), .Y(ori_ori_n439_));
  INV        o0411(.A(ori_ori_n364_), .Y(ori_ori_n440_));
  NA3        o0412(.A(ori_ori_n440_), .B(ori_ori_n353_), .C(d), .Y(ori_ori_n441_));
  NO2        o0413(.A(ori_ori_n420_), .B(ori_ori_n49_), .Y(ori_ori_n442_));
  NO3        o0414(.A(ori_ori_n63_), .B(ori_ori_n110_), .C(e), .Y(ori_ori_n443_));
  NAi21      o0415(.An(k), .B(j), .Y(ori_ori_n444_));
  NA2        o0416(.A(ori_ori_n249_), .B(ori_ori_n444_), .Y(ori_ori_n445_));
  NA3        o0417(.A(ori_ori_n445_), .B(ori_ori_n443_), .C(ori_ori_n442_), .Y(ori_ori_n446_));
  NAi21      o0418(.An(e), .B(d), .Y(ori_ori_n447_));
  INV        o0419(.A(ori_ori_n447_), .Y(ori_ori_n448_));
  NO2        o0420(.A(ori_ori_n250_), .B(ori_ori_n209_), .Y(ori_ori_n449_));
  NA3        o0421(.A(ori_ori_n449_), .B(ori_ori_n448_), .C(ori_ori_n223_), .Y(ori_ori_n450_));
  NA4        o0422(.A(ori_ori_n450_), .B(ori_ori_n446_), .C(ori_ori_n441_), .D(ori_ori_n439_), .Y(ori_ori_n451_));
  NO2        o0423(.A(ori_ori_n324_), .B(ori_ori_n209_), .Y(ori_ori_n452_));
  NA2        o0424(.A(ori_ori_n452_), .B(ori_ori_n448_), .Y(ori_ori_n453_));
  NOi31      o0425(.An(n), .B(m), .C(k), .Y(ori_ori_n454_));
  AOI220     o0426(.A0(ori_ori_n454_), .A1(ori_ori_n379_), .B0(ori_ori_n217_), .B1(ori_ori_n50_), .Y(ori_ori_n455_));
  NAi31      o0427(.An(g), .B(f), .C(c), .Y(ori_ori_n456_));
  OR3        o0428(.A(ori_ori_n456_), .B(ori_ori_n455_), .C(e), .Y(ori_ori_n457_));
  NA3        o0429(.A(ori_ori_n457_), .B(ori_ori_n453_), .C(ori_ori_n298_), .Y(ori_ori_n458_));
  NOi41      o0430(.An(ori_ori_n435_), .B(ori_ori_n458_), .C(ori_ori_n451_), .D(ori_ori_n262_), .Y(ori_ori_n459_));
  NOi32      o0431(.An(c), .Bn(a), .C(b), .Y(ori_ori_n460_));
  NA2        o0432(.A(ori_ori_n460_), .B(ori_ori_n111_), .Y(ori_ori_n461_));
  INV        o0433(.A(ori_ori_n269_), .Y(ori_ori_n462_));
  AN2        o0434(.A(e), .B(d), .Y(ori_ori_n463_));
  NA2        o0435(.A(ori_ori_n463_), .B(ori_ori_n462_), .Y(ori_ori_n464_));
  INV        o0436(.A(ori_ori_n145_), .Y(ori_ori_n465_));
  NO2        o0437(.A(ori_ori_n128_), .B(ori_ori_n41_), .Y(ori_ori_n466_));
  NO2        o0438(.A(ori_ori_n63_), .B(e), .Y(ori_ori_n467_));
  NOi31      o0439(.An(j), .B(k), .C(i), .Y(ori_ori_n468_));
  NOi21      o0440(.An(ori_ori_n162_), .B(ori_ori_n468_), .Y(ori_ori_n469_));
  NA4        o0441(.A(ori_ori_n310_), .B(ori_ori_n469_), .C(ori_ori_n258_), .D(ori_ori_n117_), .Y(ori_ori_n470_));
  AOI220     o0442(.A0(ori_ori_n470_), .A1(ori_ori_n467_), .B0(ori_ori_n466_), .B1(ori_ori_n465_), .Y(ori_ori_n471_));
  AOI210     o0443(.A0(ori_ori_n471_), .A1(ori_ori_n464_), .B0(ori_ori_n461_), .Y(ori_ori_n472_));
  NO2        o0444(.A(ori_ori_n205_), .B(ori_ori_n200_), .Y(ori_ori_n473_));
  NOi21      o0445(.An(a), .B(b), .Y(ori_ori_n474_));
  NA3        o0446(.A(e), .B(d), .C(c), .Y(ori_ori_n475_));
  NAi21      o0447(.An(ori_ori_n475_), .B(ori_ori_n474_), .Y(ori_ori_n476_));
  NO2        o0448(.A(ori_ori_n419_), .B(ori_ori_n199_), .Y(ori_ori_n477_));
  NOi21      o0449(.An(ori_ori_n476_), .B(ori_ori_n477_), .Y(ori_ori_n478_));
  AOI210     o0450(.A0(ori_ori_n264_), .A1(ori_ori_n473_), .B0(ori_ori_n478_), .Y(ori_ori_n479_));
  NO4        o0451(.A(ori_ori_n182_), .B(ori_ori_n100_), .C(ori_ori_n56_), .D(b), .Y(ori_ori_n480_));
  NA2        o0452(.A(ori_ori_n374_), .B(ori_ori_n151_), .Y(ori_ori_n481_));
  OR2        o0453(.A(k), .B(j), .Y(ori_ori_n482_));
  NA2        o0454(.A(l), .B(k), .Y(ori_ori_n483_));
  NA3        o0455(.A(ori_ori_n483_), .B(ori_ori_n482_), .C(ori_ori_n217_), .Y(ori_ori_n484_));
  AOI210     o0456(.A0(ori_ori_n230_), .A1(ori_ori_n327_), .B0(ori_ori_n80_), .Y(ori_ori_n485_));
  NOi21      o0457(.An(ori_ori_n484_), .B(ori_ori_n485_), .Y(ori_ori_n486_));
  OR3        o0458(.A(ori_ori_n486_), .B(ori_ori_n141_), .C(ori_ori_n132_), .Y(ori_ori_n487_));
  NA2        o0459(.A(ori_ori_n270_), .B(ori_ori_n124_), .Y(ori_ori_n488_));
  NO3        o0460(.A(ori_ori_n419_), .B(ori_ori_n88_), .C(ori_ori_n128_), .Y(ori_ori_n489_));
  NO2        o0461(.A(ori_ori_n489_), .B(ori_ori_n488_), .Y(ori_ori_n490_));
  NA3        o0462(.A(ori_ori_n490_), .B(ori_ori_n487_), .C(ori_ori_n481_), .Y(ori_ori_n491_));
  NO4        o0463(.A(ori_ori_n491_), .B(ori_ori_n480_), .C(ori_ori_n479_), .D(ori_ori_n472_), .Y(ori_ori_n492_));
  INV        o0464(.A(e), .Y(ori_ori_n493_));
  NO2        o0465(.A(ori_ori_n182_), .B(ori_ori_n56_), .Y(ori_ori_n494_));
  NAi31      o0466(.An(j), .B(l), .C(i), .Y(ori_ori_n495_));
  OAI210     o0467(.A0(ori_ori_n495_), .A1(ori_ori_n129_), .B0(ori_ori_n100_), .Y(ori_ori_n496_));
  NA3        o0468(.A(ori_ori_n496_), .B(ori_ori_n494_), .C(ori_ori_n493_), .Y(ori_ori_n497_));
  NO3        o0469(.A(ori_ori_n388_), .B(ori_ori_n335_), .C(ori_ori_n196_), .Y(ori_ori_n498_));
  NO2        o0470(.A(ori_ori_n388_), .B(ori_ori_n364_), .Y(ori_ori_n499_));
  NO4        o0471(.A(ori_ori_n499_), .B(ori_ori_n498_), .C(ori_ori_n179_), .D(ori_ori_n295_), .Y(ori_ori_n500_));
  NA3        o0472(.A(ori_ori_n500_), .B(ori_ori_n497_), .C(ori_ori_n238_), .Y(ori_ori_n501_));
  OAI210     o0473(.A0(ori_ori_n125_), .A1(ori_ori_n123_), .B0(n), .Y(ori_ori_n502_));
  NO2        o0474(.A(ori_ori_n502_), .B(ori_ori_n128_), .Y(ori_ori_n503_));
  AN2        o0475(.A(ori_ori_n503_), .B(ori_ori_n187_), .Y(ori_ori_n504_));
  XO2        o0476(.A(i), .B(h), .Y(ori_ori_n505_));
  NA3        o0477(.A(ori_ori_n505_), .B(ori_ori_n158_), .C(n), .Y(ori_ori_n506_));
  NAi41      o0478(.An(ori_ori_n290_), .B(ori_ori_n506_), .C(ori_ori_n455_), .D(ori_ori_n376_), .Y(ori_ori_n507_));
  NOi32      o0479(.An(ori_ori_n507_), .Bn(ori_ori_n467_), .C(ori_ori_n266_), .Y(ori_ori_n508_));
  NAi31      o0480(.An(c), .B(f), .C(d), .Y(ori_ori_n509_));
  AOI210     o0481(.A0(ori_ori_n271_), .A1(ori_ori_n190_), .B0(ori_ori_n509_), .Y(ori_ori_n510_));
  NOi21      o0482(.An(ori_ori_n78_), .B(ori_ori_n510_), .Y(ori_ori_n511_));
  NA3        o0483(.A(ori_ori_n372_), .B(ori_ori_n94_), .C(ori_ori_n93_), .Y(ori_ori_n512_));
  NA2        o0484(.A(ori_ori_n224_), .B(ori_ori_n106_), .Y(ori_ori_n513_));
  AOI210     o0485(.A0(ori_ori_n513_), .A1(ori_ori_n175_), .B0(ori_ori_n509_), .Y(ori_ori_n514_));
  AOI210     o0486(.A0(ori_ori_n351_), .A1(ori_ori_n35_), .B0(ori_ori_n476_), .Y(ori_ori_n515_));
  NOi31      o0487(.An(ori_ori_n512_), .B(ori_ori_n515_), .C(ori_ori_n514_), .Y(ori_ori_n516_));
  AN2        o0488(.A(ori_ori_n278_), .B(ori_ori_n260_), .Y(ori_ori_n517_));
  NA3        o0489(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n518_));
  NO2        o0490(.A(ori_ori_n518_), .B(ori_ori_n430_), .Y(ori_ori_n519_));
  NO2        o0491(.A(ori_ori_n519_), .B(ori_ori_n286_), .Y(ori_ori_n520_));
  NAi41      o0492(.An(ori_ori_n517_), .B(ori_ori_n520_), .C(ori_ori_n516_), .D(ori_ori_n511_), .Y(ori_ori_n521_));
  NO4        o0493(.A(ori_ori_n521_), .B(ori_ori_n508_), .C(ori_ori_n504_), .D(ori_ori_n501_), .Y(ori_ori_n522_));
  NA4        o0494(.A(ori_ori_n522_), .B(ori_ori_n492_), .C(ori_ori_n459_), .D(ori_ori_n426_), .Y(ori11));
  NO2        o0495(.A(ori_ori_n68_), .B(f), .Y(ori_ori_n524_));
  NA2        o0496(.A(j), .B(g), .Y(ori_ori_n525_));
  NAi31      o0497(.An(i), .B(m), .C(l), .Y(ori_ori_n526_));
  NA3        o0498(.A(m), .B(k), .C(j), .Y(ori_ori_n527_));
  OAI220     o0499(.A0(ori_ori_n527_), .A1(ori_ori_n128_), .B0(ori_ori_n526_), .B1(ori_ori_n525_), .Y(ori_ori_n528_));
  NA2        o0500(.A(ori_ori_n528_), .B(ori_ori_n524_), .Y(ori_ori_n529_));
  NOi32      o0501(.An(e), .Bn(b), .C(f), .Y(ori_ori_n530_));
  NA2        o0502(.A(ori_ori_n46_), .B(j), .Y(ori_ori_n531_));
  NAi31      o0503(.An(d), .B(e), .C(a), .Y(ori_ori_n532_));
  NO2        o0504(.A(ori_ori_n532_), .B(n), .Y(ori_ori_n533_));
  NA2        o0505(.A(ori_ori_n533_), .B(ori_ori_n98_), .Y(ori_ori_n534_));
  NAi41      o0506(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n535_));
  NA2        o0507(.A(j), .B(i), .Y(ori_ori_n536_));
  NAi31      o0508(.An(n), .B(m), .C(k), .Y(ori_ori_n537_));
  NO3        o0509(.A(ori_ori_n537_), .B(ori_ori_n536_), .C(ori_ori_n110_), .Y(ori_ori_n538_));
  NO4        o0510(.A(n), .B(d), .C(ori_ori_n114_), .D(a), .Y(ori_ori_n539_));
  OR2        o0511(.A(n), .B(c), .Y(ori_ori_n540_));
  NO2        o0512(.A(ori_ori_n540_), .B(ori_ori_n147_), .Y(ori_ori_n541_));
  NO2        o0513(.A(ori_ori_n541_), .B(ori_ori_n539_), .Y(ori_ori_n542_));
  NOi32      o0514(.An(g), .Bn(f), .C(i), .Y(ori_ori_n543_));
  AOI220     o0515(.A0(ori_ori_n543_), .A1(ori_ori_n96_), .B0(ori_ori_n528_), .B1(f), .Y(ori_ori_n544_));
  NO2        o0516(.A(ori_ori_n269_), .B(ori_ori_n49_), .Y(ori_ori_n545_));
  NO2        o0517(.A(ori_ori_n544_), .B(ori_ori_n542_), .Y(ori_ori_n546_));
  INV        o0518(.A(ori_ori_n546_), .Y(ori_ori_n547_));
  NA2        o0519(.A(ori_ori_n137_), .B(ori_ori_n34_), .Y(ori_ori_n548_));
  OAI220     o0520(.A0(ori_ori_n548_), .A1(m), .B0(ori_ori_n531_), .B1(ori_ori_n230_), .Y(ori_ori_n549_));
  NOi41      o0521(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n550_));
  NAi32      o0522(.An(e), .Bn(b), .C(c), .Y(ori_ori_n551_));
  OR2        o0523(.A(ori_ori_n551_), .B(ori_ori_n80_), .Y(ori_ori_n552_));
  AN2        o0524(.A(ori_ori_n328_), .B(ori_ori_n307_), .Y(ori_ori_n553_));
  NA2        o0525(.A(ori_ori_n553_), .B(ori_ori_n552_), .Y(ori_ori_n554_));
  OA210      o0526(.A0(ori_ori_n554_), .A1(ori_ori_n550_), .B0(ori_ori_n549_), .Y(ori_ori_n555_));
  OAI220     o0527(.A0(ori_ori_n390_), .A1(ori_ori_n389_), .B0(ori_ori_n526_), .B1(ori_ori_n525_), .Y(ori_ori_n556_));
  NAi31      o0528(.An(d), .B(c), .C(a), .Y(ori_ori_n557_));
  NO2        o0529(.A(ori_ori_n557_), .B(n), .Y(ori_ori_n558_));
  NO3        o0530(.A(ori_ori_n61_), .B(ori_ori_n49_), .C(ori_ori_n210_), .Y(ori_ori_n559_));
  NO2        o0531(.A(ori_ori_n227_), .B(ori_ori_n108_), .Y(ori_ori_n560_));
  OAI210     o0532(.A0(ori_ori_n559_), .A1(ori_ori_n391_), .B0(ori_ori_n560_), .Y(ori_ori_n561_));
  INV        o0533(.A(ori_ori_n561_), .Y(ori_ori_n562_));
  INV        o0534(.A(ori_ori_n421_), .Y(ori_ori_n563_));
  NA2        o0535(.A(ori_ori_n556_), .B(f), .Y(ori_ori_n564_));
  NAi32      o0536(.An(d), .Bn(a), .C(b), .Y(ori_ori_n565_));
  NO2        o0537(.A(ori_ori_n565_), .B(ori_ori_n49_), .Y(ori_ori_n566_));
  NA2        o0538(.A(h), .B(f), .Y(ori_ori_n567_));
  NO2        o0539(.A(ori_ori_n567_), .B(ori_ori_n91_), .Y(ori_ori_n568_));
  NO3        o0540(.A(ori_ori_n171_), .B(ori_ori_n168_), .C(g), .Y(ori_ori_n569_));
  AOI220     o0541(.A0(ori_ori_n569_), .A1(ori_ori_n58_), .B0(ori_ori_n568_), .B1(ori_ori_n566_), .Y(ori_ori_n570_));
  OAI210     o0542(.A0(ori_ori_n564_), .A1(ori_ori_n563_), .B0(ori_ori_n570_), .Y(ori_ori_n571_));
  AN3        o0543(.A(j), .B(h), .C(g), .Y(ori_ori_n572_));
  NO2        o0544(.A(ori_ori_n144_), .B(c), .Y(ori_ori_n573_));
  NA3        o0545(.A(ori_ori_n573_), .B(ori_ori_n572_), .C(ori_ori_n454_), .Y(ori_ori_n574_));
  NA3        o0546(.A(f), .B(d), .C(b), .Y(ori_ori_n575_));
  NO4        o0547(.A(ori_ori_n575_), .B(ori_ori_n171_), .C(ori_ori_n168_), .D(g), .Y(ori_ori_n576_));
  NAi21      o0548(.An(ori_ori_n576_), .B(ori_ori_n574_), .Y(ori_ori_n577_));
  NO4        o0549(.A(ori_ori_n577_), .B(ori_ori_n571_), .C(ori_ori_n562_), .D(ori_ori_n555_), .Y(ori_ori_n578_));
  AN4        o0550(.A(ori_ori_n578_), .B(ori_ori_n547_), .C(ori_ori_n534_), .D(ori_ori_n529_), .Y(ori_ori_n579_));
  INV        o0551(.A(k), .Y(ori_ori_n580_));
  NA3        o0552(.A(l), .B(ori_ori_n580_), .C(i), .Y(ori_ori_n581_));
  INV        o0553(.A(ori_ori_n581_), .Y(ori_ori_n582_));
  NA4        o0554(.A(ori_ori_n387_), .B(ori_ori_n410_), .C(ori_ori_n176_), .D(ori_ori_n111_), .Y(ori_ori_n583_));
  NAi32      o0555(.An(h), .Bn(f), .C(g), .Y(ori_ori_n584_));
  NAi41      o0556(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n585_));
  OAI210     o0557(.A0(ori_ori_n532_), .A1(n), .B0(ori_ori_n585_), .Y(ori_ori_n586_));
  NA2        o0558(.A(ori_ori_n586_), .B(m), .Y(ori_ori_n587_));
  NAi31      o0559(.An(h), .B(g), .C(f), .Y(ori_ori_n588_));
  OR2        o0560(.A(ori_ori_n587_), .B(ori_ori_n584_), .Y(ori_ori_n589_));
  NO3        o0561(.A(ori_ori_n584_), .B(ori_ori_n68_), .C(ori_ori_n69_), .Y(ori_ori_n590_));
  NO4        o0562(.A(ori_ori_n588_), .B(ori_ori_n540_), .C(ori_ori_n147_), .D(ori_ori_n69_), .Y(ori_ori_n591_));
  OR2        o0563(.A(ori_ori_n591_), .B(ori_ori_n590_), .Y(ori_ori_n592_));
  NAi31      o0564(.An(ori_ori_n592_), .B(ori_ori_n589_), .C(ori_ori_n583_), .Y(ori_ori_n593_));
  NAi31      o0565(.An(f), .B(h), .C(g), .Y(ori_ori_n594_));
  NOi32      o0566(.An(b), .Bn(a), .C(c), .Y(ori_ori_n595_));
  NOi32      o0567(.An(d), .Bn(a), .C(e), .Y(ori_ori_n596_));
  NA2        o0568(.A(ori_ori_n596_), .B(ori_ori_n111_), .Y(ori_ori_n597_));
  NO2        o0569(.A(n), .B(c), .Y(ori_ori_n598_));
  NA3        o0570(.A(ori_ori_n598_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n599_));
  NAi32      o0571(.An(n), .Bn(f), .C(m), .Y(ori_ori_n600_));
  NA3        o0572(.A(ori_ori_n600_), .B(ori_ori_n599_), .C(ori_ori_n597_), .Y(ori_ori_n601_));
  NOi32      o0573(.An(e), .Bn(a), .C(d), .Y(ori_ori_n602_));
  AOI210     o0574(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n602_), .Y(ori_ori_n603_));
  AOI210     o0575(.A0(ori_ori_n603_), .A1(ori_ori_n209_), .B0(ori_ori_n548_), .Y(ori_ori_n604_));
  NA2        o0576(.A(ori_ori_n604_), .B(ori_ori_n601_), .Y(ori_ori_n605_));
  OAI210     o0577(.A0(ori_ori_n245_), .A1(ori_ori_n83_), .B0(ori_ori_n605_), .Y(ori_ori_n606_));
  AOI210     o0578(.A0(ori_ori_n593_), .A1(ori_ori_n582_), .B0(ori_ori_n606_), .Y(ori_ori_n607_));
  NO3        o0579(.A(ori_ori_n305_), .B(ori_ori_n60_), .C(n), .Y(ori_ori_n608_));
  NA3        o0580(.A(ori_ori_n509_), .B(ori_ori_n166_), .C(ori_ori_n165_), .Y(ori_ori_n609_));
  NA2        o0581(.A(ori_ori_n456_), .B(ori_ori_n227_), .Y(ori_ori_n610_));
  OR2        o0582(.A(ori_ori_n610_), .B(ori_ori_n609_), .Y(ori_ori_n611_));
  NA2        o0583(.A(ori_ori_n611_), .B(ori_ori_n608_), .Y(ori_ori_n612_));
  NO2        o0584(.A(ori_ori_n612_), .B(ori_ori_n83_), .Y(ori_ori_n613_));
  NA3        o0585(.A(ori_ori_n550_), .B(ori_ori_n330_), .C(ori_ori_n46_), .Y(ori_ori_n614_));
  NOi32      o0586(.An(e), .Bn(c), .C(f), .Y(ori_ori_n615_));
  NOi21      o0587(.An(f), .B(g), .Y(ori_ori_n616_));
  NO2        o0588(.A(ori_ori_n616_), .B(ori_ori_n207_), .Y(ori_ori_n617_));
  AOI220     o0589(.A0(ori_ori_n617_), .A1(ori_ori_n384_), .B0(ori_ori_n615_), .B1(ori_ori_n170_), .Y(ori_ori_n618_));
  NA3        o0590(.A(ori_ori_n618_), .B(ori_ori_n614_), .C(ori_ori_n173_), .Y(ori_ori_n619_));
  AOI210     o0591(.A0(ori_ori_n535_), .A1(ori_ori_n388_), .B0(ori_ori_n291_), .Y(ori_ori_n620_));
  NA2        o0592(.A(ori_ori_n620_), .B(ori_ori_n261_), .Y(ori_ori_n621_));
  NOi21      o0593(.An(j), .B(l), .Y(ori_ori_n622_));
  NAi21      o0594(.An(k), .B(h), .Y(ori_ori_n623_));
  NO2        o0595(.A(ori_ori_n623_), .B(ori_ori_n259_), .Y(ori_ori_n624_));
  NA2        o0596(.A(ori_ori_n624_), .B(ori_ori_n622_), .Y(ori_ori_n625_));
  OR2        o0597(.A(ori_ori_n625_), .B(ori_ori_n587_), .Y(ori_ori_n626_));
  NOi31      o0598(.An(m), .B(n), .C(k), .Y(ori_ori_n627_));
  NA2        o0599(.A(ori_ori_n622_), .B(ori_ori_n627_), .Y(ori_ori_n628_));
  NO2        o0600(.A(ori_ori_n388_), .B(ori_ori_n291_), .Y(ori_ori_n629_));
  NAi21      o0601(.An(ori_ori_n628_), .B(ori_ori_n629_), .Y(ori_ori_n630_));
  NO2        o0602(.A(ori_ori_n299_), .B(ori_ori_n594_), .Y(ori_ori_n631_));
  NO2        o0603(.A(ori_ori_n532_), .B(ori_ori_n49_), .Y(ori_ori_n632_));
  NA2        o0604(.A(ori_ori_n632_), .B(ori_ori_n631_), .Y(ori_ori_n633_));
  NA4        o0605(.A(ori_ori_n633_), .B(ori_ori_n630_), .C(ori_ori_n626_), .D(ori_ori_n621_), .Y(ori_ori_n634_));
  NA2        o0606(.A(ori_ori_n106_), .B(ori_ori_n36_), .Y(ori_ori_n635_));
  NO2        o0607(.A(k), .B(ori_ori_n210_), .Y(ori_ori_n636_));
  INV        o0608(.A(ori_ori_n353_), .Y(ori_ori_n637_));
  NO2        o0609(.A(ori_ori_n637_), .B(n), .Y(ori_ori_n638_));
  NAi31      o0610(.An(ori_ori_n635_), .B(ori_ori_n638_), .C(ori_ori_n636_), .Y(ori_ori_n639_));
  NO2        o0611(.A(ori_ori_n531_), .B(ori_ori_n171_), .Y(ori_ori_n640_));
  NA3        o0612(.A(ori_ori_n551_), .B(ori_ori_n266_), .C(ori_ori_n142_), .Y(ori_ori_n641_));
  NA2        o0613(.A(ori_ori_n505_), .B(ori_ori_n158_), .Y(ori_ori_n642_));
  NO3        o0614(.A(ori_ori_n385_), .B(ori_ori_n642_), .C(ori_ori_n83_), .Y(ori_ori_n643_));
  AOI210     o0615(.A0(ori_ori_n641_), .A1(ori_ori_n640_), .B0(ori_ori_n643_), .Y(ori_ori_n644_));
  AN3        o0616(.A(f), .B(d), .C(b), .Y(ori_ori_n645_));
  OAI210     o0617(.A0(ori_ori_n645_), .A1(ori_ori_n127_), .B0(n), .Y(ori_ori_n646_));
  NA3        o0618(.A(ori_ori_n505_), .B(ori_ori_n158_), .C(ori_ori_n210_), .Y(ori_ori_n647_));
  AOI210     o0619(.A0(ori_ori_n646_), .A1(ori_ori_n229_), .B0(ori_ori_n647_), .Y(ori_ori_n648_));
  NAi31      o0620(.An(m), .B(n), .C(k), .Y(ori_ori_n649_));
  OR2        o0621(.A(ori_ori_n132_), .B(ori_ori_n60_), .Y(ori_ori_n650_));
  OAI210     o0622(.A0(ori_ori_n650_), .A1(ori_ori_n649_), .B0(ori_ori_n247_), .Y(ori_ori_n651_));
  OAI210     o0623(.A0(ori_ori_n651_), .A1(ori_ori_n648_), .B0(j), .Y(ori_ori_n652_));
  NA3        o0624(.A(ori_ori_n652_), .B(ori_ori_n644_), .C(ori_ori_n639_), .Y(ori_ori_n653_));
  NO4        o0625(.A(ori_ori_n653_), .B(ori_ori_n634_), .C(ori_ori_n619_), .D(ori_ori_n613_), .Y(ori_ori_n654_));
  NA2        o0626(.A(ori_ori_n372_), .B(ori_ori_n161_), .Y(ori_ori_n655_));
  NAi31      o0627(.An(g), .B(h), .C(f), .Y(ori_ori_n656_));
  OA210      o0628(.A0(ori_ori_n532_), .A1(n), .B0(ori_ori_n585_), .Y(ori_ori_n657_));
  NO2        o0629(.A(ori_ori_n657_), .B(ori_ori_n87_), .Y(ori_ori_n658_));
  INV        o0630(.A(ori_ori_n658_), .Y(ori_ori_n659_));
  AOI210     o0631(.A0(ori_ori_n659_), .A1(ori_ori_n655_), .B0(ori_ori_n527_), .Y(ori_ori_n660_));
  NO3        o0632(.A(g), .B(ori_ori_n209_), .C(ori_ori_n56_), .Y(ori_ori_n661_));
  NAi21      o0633(.An(h), .B(j), .Y(ori_ori_n662_));
  NO2        o0634(.A(ori_ori_n513_), .B(ori_ori_n83_), .Y(ori_ori_n663_));
  OAI210     o0635(.A0(ori_ori_n663_), .A1(ori_ori_n384_), .B0(ori_ori_n661_), .Y(ori_ori_n664_));
  OR2        o0636(.A(ori_ori_n68_), .B(ori_ori_n69_), .Y(ori_ori_n665_));
  NA2        o0637(.A(ori_ori_n595_), .B(ori_ori_n332_), .Y(ori_ori_n666_));
  OA220      o0638(.A0(ori_ori_n628_), .A1(ori_ori_n666_), .B0(ori_ori_n625_), .B1(ori_ori_n665_), .Y(ori_ori_n667_));
  AN2        o0639(.A(h), .B(f), .Y(ori_ori_n668_));
  NA2        o0640(.A(ori_ori_n668_), .B(ori_ori_n37_), .Y(ori_ori_n669_));
  NA2        o0641(.A(ori_ori_n96_), .B(ori_ori_n46_), .Y(ori_ori_n670_));
  OAI220     o0642(.A0(ori_ori_n670_), .A1(ori_ori_n321_), .B0(ori_ori_n669_), .B1(ori_ori_n461_), .Y(ori_ori_n671_));
  AOI210     o0643(.A0(ori_ori_n565_), .A1(ori_ori_n420_), .B0(ori_ori_n49_), .Y(ori_ori_n672_));
  OAI220     o0644(.A0(ori_ori_n588_), .A1(ori_ori_n581_), .B0(ori_ori_n314_), .B1(ori_ori_n525_), .Y(ori_ori_n673_));
  AOI210     o0645(.A0(ori_ori_n673_), .A1(ori_ori_n672_), .B0(ori_ori_n671_), .Y(ori_ori_n674_));
  NA3        o0646(.A(ori_ori_n674_), .B(ori_ori_n667_), .C(ori_ori_n664_), .Y(ori_ori_n675_));
  NO2        o0647(.A(ori_ori_n249_), .B(f), .Y(ori_ori_n676_));
  NO2        o0648(.A(ori_ori_n616_), .B(ori_ori_n60_), .Y(ori_ori_n677_));
  NO3        o0649(.A(ori_ori_n677_), .B(ori_ori_n676_), .C(ori_ori_n34_), .Y(ori_ori_n678_));
  NA2        o0650(.A(ori_ori_n317_), .B(ori_ori_n137_), .Y(ori_ori_n679_));
  NA2        o0651(.A(ori_ori_n129_), .B(ori_ori_n49_), .Y(ori_ori_n680_));
  AOI220     o0652(.A0(ori_ori_n680_), .A1(ori_ori_n530_), .B0(ori_ori_n353_), .B1(ori_ori_n111_), .Y(ori_ori_n681_));
  OA220      o0653(.A0(ori_ori_n681_), .A1(ori_ori_n548_), .B0(ori_ori_n351_), .B1(ori_ori_n109_), .Y(ori_ori_n682_));
  OAI210     o0654(.A0(ori_ori_n679_), .A1(ori_ori_n678_), .B0(ori_ori_n682_), .Y(ori_ori_n683_));
  NO3        o0655(.A(ori_ori_n395_), .B(ori_ori_n187_), .C(ori_ori_n186_), .Y(ori_ori_n684_));
  NA2        o0656(.A(ori_ori_n684_), .B(ori_ori_n227_), .Y(ori_ori_n685_));
  NA3        o0657(.A(ori_ori_n685_), .B(ori_ori_n251_), .C(j), .Y(ori_ori_n686_));
  NO3        o0658(.A(ori_ori_n456_), .B(ori_ori_n168_), .C(i), .Y(ori_ori_n687_));
  NA2        o0659(.A(ori_ori_n460_), .B(ori_ori_n80_), .Y(ori_ori_n688_));
  NO4        o0660(.A(ori_ori_n527_), .B(ori_ori_n688_), .C(ori_ori_n128_), .D(ori_ori_n209_), .Y(ori_ori_n689_));
  INV        o0661(.A(ori_ori_n689_), .Y(ori_ori_n690_));
  NA4        o0662(.A(ori_ori_n690_), .B(ori_ori_n686_), .C(ori_ori_n512_), .D(ori_ori_n393_), .Y(ori_ori_n691_));
  NO4        o0663(.A(ori_ori_n691_), .B(ori_ori_n683_), .C(ori_ori_n675_), .D(ori_ori_n660_), .Y(ori_ori_n692_));
  NA4        o0664(.A(ori_ori_n692_), .B(ori_ori_n654_), .C(ori_ori_n607_), .D(ori_ori_n579_), .Y(ori08));
  NO2        o0665(.A(k), .B(h), .Y(ori_ori_n694_));
  AO210      o0666(.A0(ori_ori_n249_), .A1(ori_ori_n444_), .B0(ori_ori_n694_), .Y(ori_ori_n695_));
  NO2        o0667(.A(ori_ori_n695_), .B(ori_ori_n289_), .Y(ori_ori_n696_));
  NA2        o0668(.A(ori_ori_n615_), .B(ori_ori_n80_), .Y(ori_ori_n697_));
  NA2        o0669(.A(ori_ori_n697_), .B(ori_ori_n456_), .Y(ori_ori_n698_));
  AOI210     o0670(.A0(ori_ori_n698_), .A1(ori_ori_n696_), .B0(ori_ori_n489_), .Y(ori_ori_n699_));
  NA2        o0671(.A(ori_ori_n80_), .B(ori_ori_n108_), .Y(ori_ori_n700_));
  NO2        o0672(.A(ori_ori_n700_), .B(ori_ori_n57_), .Y(ori_ori_n701_));
  NO4        o0673(.A(ori_ori_n369_), .B(ori_ori_n110_), .C(j), .D(ori_ori_n210_), .Y(ori_ori_n702_));
  NA2        o0674(.A(ori_ori_n575_), .B(ori_ori_n229_), .Y(ori_ori_n703_));
  AOI220     o0675(.A0(ori_ori_n703_), .A1(ori_ori_n338_), .B0(ori_ori_n702_), .B1(ori_ori_n701_), .Y(ori_ori_n704_));
  AOI210     o0676(.A0(ori_ori_n575_), .A1(ori_ori_n154_), .B0(ori_ori_n80_), .Y(ori_ori_n705_));
  NA4        o0677(.A(ori_ori_n212_), .B(ori_ori_n137_), .C(ori_ori_n45_), .D(h), .Y(ori_ori_n706_));
  AN2        o0678(.A(l), .B(k), .Y(ori_ori_n707_));
  NA4        o0679(.A(ori_ori_n707_), .B(ori_ori_n106_), .C(ori_ori_n69_), .D(ori_ori_n210_), .Y(ori_ori_n708_));
  OAI210     o0680(.A0(ori_ori_n706_), .A1(g), .B0(ori_ori_n708_), .Y(ori_ori_n709_));
  NA2        o0681(.A(ori_ori_n709_), .B(ori_ori_n705_), .Y(ori_ori_n710_));
  NA4        o0682(.A(ori_ori_n710_), .B(ori_ori_n704_), .C(ori_ori_n699_), .D(ori_ori_n340_), .Y(ori_ori_n711_));
  AN2        o0683(.A(ori_ori_n533_), .B(ori_ori_n92_), .Y(ori_ori_n712_));
  NO4        o0684(.A(ori_ori_n168_), .B(ori_ori_n383_), .C(ori_ori_n110_), .D(g), .Y(ori_ori_n713_));
  AOI210     o0685(.A0(ori_ori_n713_), .A1(ori_ori_n703_), .B0(ori_ori_n519_), .Y(ori_ori_n714_));
  NO2        o0686(.A(ori_ori_n38_), .B(ori_ori_n209_), .Y(ori_ori_n715_));
  NA2        o0687(.A(ori_ori_n617_), .B(ori_ori_n337_), .Y(ori_ori_n716_));
  NAi31      o0688(.An(ori_ori_n712_), .B(ori_ori_n716_), .C(ori_ori_n714_), .Y(ori_ori_n717_));
  OAI210     o0689(.A0(ori_ori_n551_), .A1(ori_ori_n47_), .B0(ori_ori_n650_), .Y(ori_ori_n718_));
  NO2        o0690(.A(ori_ori_n483_), .B(ori_ori_n129_), .Y(ori_ori_n719_));
  NA2        o0691(.A(ori_ori_n719_), .B(ori_ori_n718_), .Y(ori_ori_n720_));
  NO3        o0692(.A(ori_ori_n305_), .B(ori_ori_n128_), .C(ori_ori_n41_), .Y(ori_ori_n721_));
  NAi21      o0693(.An(ori_ori_n721_), .B(ori_ori_n708_), .Y(ori_ori_n722_));
  NA2        o0694(.A(ori_ori_n695_), .B(ori_ori_n133_), .Y(ori_ori_n723_));
  AOI220     o0695(.A0(ori_ori_n723_), .A1(ori_ori_n394_), .B0(ori_ori_n722_), .B1(ori_ori_n72_), .Y(ori_ori_n724_));
  NA2        o0696(.A(ori_ori_n720_), .B(ori_ori_n724_), .Y(ori_ori_n725_));
  NA2        o0697(.A(ori_ori_n353_), .B(ori_ori_n43_), .Y(ori_ori_n726_));
  NA3        o0698(.A(ori_ori_n685_), .B(ori_ori_n323_), .C(ori_ori_n375_), .Y(ori_ori_n727_));
  NA3        o0699(.A(m), .B(l), .C(k), .Y(ori_ori_n728_));
  NA3        o0700(.A(ori_ori_n111_), .B(k), .C(ori_ori_n83_), .Y(ori_ori_n729_));
  NA2        o0701(.A(ori_ori_n727_), .B(ori_ori_n726_), .Y(ori_ori_n730_));
  NO4        o0702(.A(ori_ori_n730_), .B(ori_ori_n725_), .C(ori_ori_n717_), .D(ori_ori_n711_), .Y(ori_ori_n731_));
  NA2        o0703(.A(ori_ori_n617_), .B(ori_ori_n384_), .Y(ori_ori_n732_));
  NOi31      o0704(.An(g), .B(h), .C(f), .Y(ori_ori_n733_));
  NA2        o0705(.A(ori_ori_n632_), .B(ori_ori_n733_), .Y(ori_ori_n734_));
  OR2        o0706(.A(ori_ori_n734_), .B(ori_ori_n536_), .Y(ori_ori_n735_));
  NO3        o0707(.A(ori_ori_n388_), .B(ori_ori_n525_), .C(h), .Y(ori_ori_n736_));
  AOI210     o0708(.A0(ori_ori_n736_), .A1(ori_ori_n111_), .B0(ori_ori_n499_), .Y(ori_ori_n737_));
  NA4        o0709(.A(ori_ori_n737_), .B(ori_ori_n735_), .C(ori_ori_n732_), .D(ori_ori_n248_), .Y(ori_ori_n738_));
  NA2        o0710(.A(ori_ori_n707_), .B(ori_ori_n69_), .Y(ori_ori_n739_));
  NO4        o0711(.A(ori_ori_n684_), .B(ori_ori_n168_), .C(n), .D(i), .Y(ori_ori_n740_));
  NOi21      o0712(.An(h), .B(j), .Y(ori_ori_n741_));
  NA2        o0713(.A(ori_ori_n741_), .B(f), .Y(ori_ori_n742_));
  NO2        o0714(.A(ori_ori_n740_), .B(ori_ori_n687_), .Y(ori_ori_n743_));
  NO2        o0715(.A(ori_ori_n743_), .B(ori_ori_n739_), .Y(ori_ori_n744_));
  AOI210     o0716(.A0(ori_ori_n738_), .A1(l), .B0(ori_ori_n744_), .Y(ori_ori_n745_));
  NO2        o0717(.A(j), .B(i), .Y(ori_ori_n746_));
  NA3        o0718(.A(ori_ori_n746_), .B(ori_ori_n76_), .C(l), .Y(ori_ori_n747_));
  NA2        o0719(.A(ori_ori_n746_), .B(ori_ori_n33_), .Y(ori_ori_n748_));
  OR2        o0720(.A(ori_ori_n747_), .B(ori_ori_n587_), .Y(ori_ori_n749_));
  NO3        o0721(.A(ori_ori_n149_), .B(ori_ori_n49_), .C(ori_ori_n108_), .Y(ori_ori_n750_));
  NO3        o0722(.A(ori_ori_n540_), .B(ori_ori_n147_), .C(ori_ori_n69_), .Y(ori_ori_n751_));
  NO3        o0723(.A(ori_ori_n483_), .B(ori_ori_n431_), .C(j), .Y(ori_ori_n752_));
  OAI210     o0724(.A0(ori_ori_n751_), .A1(ori_ori_n750_), .B0(ori_ori_n752_), .Y(ori_ori_n753_));
  OAI210     o0725(.A0(ori_ori_n734_), .A1(ori_ori_n61_), .B0(ori_ori_n753_), .Y(ori_ori_n754_));
  INV        o0726(.A(j), .Y(ori_ori_n755_));
  NO3        o0727(.A(ori_ori_n289_), .B(ori_ori_n755_), .C(ori_ori_n40_), .Y(ori_ori_n756_));
  AOI210     o0728(.A0(ori_ori_n530_), .A1(n), .B0(ori_ori_n550_), .Y(ori_ori_n757_));
  NA2        o0729(.A(ori_ori_n757_), .B(ori_ori_n553_), .Y(ori_ori_n758_));
  AN3        o0730(.A(ori_ori_n758_), .B(ori_ori_n756_), .C(ori_ori_n95_), .Y(ori_ori_n759_));
  NO3        o0731(.A(ori_ori_n168_), .B(ori_ori_n383_), .C(ori_ori_n110_), .Y(ori_ori_n760_));
  AOI220     o0732(.A0(ori_ori_n760_), .A1(ori_ori_n243_), .B0(ori_ori_n610_), .B1(ori_ori_n297_), .Y(ori_ori_n761_));
  NAi31      o0733(.An(ori_ori_n603_), .B(ori_ori_n89_), .C(ori_ori_n80_), .Y(ori_ori_n762_));
  NA2        o0734(.A(ori_ori_n762_), .B(ori_ori_n761_), .Y(ori_ori_n763_));
  NO2        o0735(.A(ori_ori_n289_), .B(ori_ori_n133_), .Y(ori_ori_n764_));
  AOI220     o0736(.A0(ori_ori_n764_), .A1(ori_ori_n617_), .B0(ori_ori_n721_), .B1(ori_ori_n705_), .Y(ori_ori_n765_));
  NO2        o0737(.A(ori_ori_n728_), .B(ori_ori_n87_), .Y(ori_ori_n766_));
  NA2        o0738(.A(ori_ori_n766_), .B(ori_ori_n586_), .Y(ori_ori_n767_));
  NO2        o0739(.A(ori_ori_n588_), .B(ori_ori_n115_), .Y(ori_ori_n768_));
  OAI210     o0740(.A0(ori_ori_n768_), .A1(ori_ori_n752_), .B0(ori_ori_n672_), .Y(ori_ori_n769_));
  NA3        o0741(.A(ori_ori_n769_), .B(ori_ori_n767_), .C(ori_ori_n765_), .Y(ori_ori_n770_));
  OR4        o0742(.A(ori_ori_n770_), .B(ori_ori_n763_), .C(ori_ori_n759_), .D(ori_ori_n754_), .Y(ori_ori_n771_));
  NA3        o0743(.A(ori_ori_n757_), .B(ori_ori_n553_), .C(ori_ori_n552_), .Y(ori_ori_n772_));
  NA4        o0744(.A(ori_ori_n772_), .B(ori_ori_n212_), .C(ori_ori_n444_), .D(ori_ori_n34_), .Y(ori_ori_n773_));
  NO4        o0745(.A(ori_ori_n483_), .B(ori_ori_n427_), .C(j), .D(f), .Y(ori_ori_n774_));
  OAI220     o0746(.A0(ori_ori_n706_), .A1(ori_ori_n697_), .B0(ori_ori_n321_), .B1(ori_ori_n38_), .Y(ori_ori_n775_));
  AOI210     o0747(.A0(ori_ori_n774_), .A1(ori_ori_n255_), .B0(ori_ori_n775_), .Y(ori_ori_n776_));
  NA3        o0748(.A(ori_ori_n543_), .B(ori_ori_n282_), .C(h), .Y(ori_ori_n777_));
  NOi21      o0749(.An(ori_ori_n672_), .B(ori_ori_n777_), .Y(ori_ori_n778_));
  NO2        o0750(.A(ori_ori_n88_), .B(ori_ori_n47_), .Y(ori_ori_n779_));
  NO2        o0751(.A(ori_ori_n777_), .B(ori_ori_n599_), .Y(ori_ori_n780_));
  AOI210     o0752(.A0(ori_ori_n779_), .A1(ori_ori_n638_), .B0(ori_ori_n780_), .Y(ori_ori_n781_));
  NAi41      o0753(.An(ori_ori_n778_), .B(ori_ori_n781_), .C(ori_ori_n776_), .D(ori_ori_n773_), .Y(ori_ori_n782_));
  NA2        o0754(.A(ori_ori_n766_), .B(ori_ori_n234_), .Y(ori_ori_n783_));
  NO2        o0755(.A(ori_ori_n657_), .B(ori_ori_n69_), .Y(ori_ori_n784_));
  AOI210     o0756(.A0(ori_ori_n774_), .A1(ori_ori_n784_), .B0(ori_ori_n325_), .Y(ori_ori_n785_));
  OAI210     o0757(.A0(ori_ori_n728_), .A1(ori_ori_n656_), .B0(ori_ori_n518_), .Y(ori_ori_n786_));
  NA3        o0758(.A(ori_ori_n246_), .B(ori_ori_n59_), .C(b), .Y(ori_ori_n787_));
  AOI220     o0759(.A0(ori_ori_n598_), .A1(ori_ori_n29_), .B0(ori_ori_n460_), .B1(ori_ori_n80_), .Y(ori_ori_n788_));
  NA2        o0760(.A(ori_ori_n788_), .B(ori_ori_n787_), .Y(ori_ori_n789_));
  NA2        o0761(.A(ori_ori_n789_), .B(ori_ori_n786_), .Y(ori_ori_n790_));
  NA3        o0762(.A(ori_ori_n790_), .B(ori_ori_n785_), .C(ori_ori_n783_), .Y(ori_ori_n791_));
  NOi41      o0763(.An(ori_ori_n749_), .B(ori_ori_n791_), .C(ori_ori_n782_), .D(ori_ori_n771_), .Y(ori_ori_n792_));
  NO3        o0764(.A(ori_ori_n331_), .B(ori_ori_n291_), .C(ori_ori_n110_), .Y(ori_ori_n793_));
  NA2        o0765(.A(ori_ori_n793_), .B(ori_ori_n758_), .Y(ori_ori_n794_));
  NO3        o0766(.A(ori_ori_n525_), .B(ori_ori_n90_), .C(h), .Y(ori_ori_n795_));
  NA2        o0767(.A(ori_ori_n795_), .B(ori_ori_n701_), .Y(ori_ori_n796_));
  NA3        o0768(.A(ori_ori_n796_), .B(ori_ori_n794_), .C(ori_ori_n396_), .Y(ori_ori_n797_));
  OR2        o0769(.A(ori_ori_n656_), .B(ori_ori_n88_), .Y(ori_ori_n798_));
  NOi31      o0770(.An(b), .B(d), .C(a), .Y(ori_ori_n799_));
  NO2        o0771(.A(ori_ori_n799_), .B(ori_ori_n596_), .Y(ori_ori_n800_));
  NO2        o0772(.A(ori_ori_n800_), .B(n), .Y(ori_ori_n801_));
  NOi21      o0773(.An(ori_ori_n788_), .B(ori_ori_n801_), .Y(ori_ori_n802_));
  NO2        o0774(.A(ori_ori_n802_), .B(ori_ori_n798_), .Y(ori_ori_n803_));
  NO2        o0775(.A(ori_ori_n551_), .B(ori_ori_n80_), .Y(ori_ori_n804_));
  NA2        o0776(.A(ori_ori_n793_), .B(ori_ori_n804_), .Y(ori_ori_n805_));
  OAI210     o0777(.A0(ori_ori_n706_), .A1(ori_ori_n385_), .B0(ori_ori_n805_), .Y(ori_ori_n806_));
  NO2        o0778(.A(ori_ori_n684_), .B(n), .Y(ori_ori_n807_));
  AOI220     o0779(.A0(ori_ori_n764_), .A1(ori_ori_n661_), .B0(ori_ori_n807_), .B1(ori_ori_n696_), .Y(ori_ori_n808_));
  NO2        o0780(.A(ori_ori_n311_), .B(ori_ori_n233_), .Y(ori_ori_n809_));
  OAI210     o0781(.A0(ori_ori_n92_), .A1(ori_ori_n89_), .B0(ori_ori_n809_), .Y(ori_ori_n810_));
  INV        o0782(.A(ori_ori_n810_), .Y(ori_ori_n811_));
  NA2        o0783(.A(ori_ori_n713_), .B(ori_ori_n339_), .Y(ori_ori_n812_));
  OAI210     o0784(.A0(ori_ori_n591_), .A1(ori_ori_n590_), .B0(ori_ori_n354_), .Y(ori_ori_n813_));
  AN2        o0785(.A(ori_ori_n813_), .B(ori_ori_n812_), .Y(ori_ori_n814_));
  NAi31      o0786(.An(ori_ori_n811_), .B(ori_ori_n814_), .C(ori_ori_n808_), .Y(ori_ori_n815_));
  NO4        o0787(.A(ori_ori_n815_), .B(ori_ori_n806_), .C(ori_ori_n803_), .D(ori_ori_n797_), .Y(ori_ori_n816_));
  NA4        o0788(.A(ori_ori_n816_), .B(ori_ori_n792_), .C(ori_ori_n745_), .D(ori_ori_n731_), .Y(ori09));
  INV        o0789(.A(ori_ori_n120_), .Y(ori_ori_n818_));
  NA2        o0790(.A(f), .B(e), .Y(ori_ori_n819_));
  NO2        o0791(.A(ori_ori_n222_), .B(ori_ori_n110_), .Y(ori_ori_n820_));
  NA2        o0792(.A(ori_ori_n820_), .B(g), .Y(ori_ori_n821_));
  NA4        o0793(.A(ori_ori_n299_), .B(ori_ori_n469_), .C(ori_ori_n258_), .D(ori_ori_n117_), .Y(ori_ori_n822_));
  AOI210     o0794(.A0(ori_ori_n822_), .A1(g), .B0(ori_ori_n466_), .Y(ori_ori_n823_));
  AOI210     o0795(.A0(ori_ori_n823_), .A1(ori_ori_n821_), .B0(ori_ori_n819_), .Y(ori_ori_n824_));
  NA2        o0796(.A(ori_ori_n437_), .B(e), .Y(ori_ori_n825_));
  NO2        o0797(.A(ori_ori_n825_), .B(ori_ori_n509_), .Y(ori_ori_n826_));
  AOI210     o0798(.A0(ori_ori_n824_), .A1(ori_ori_n818_), .B0(ori_ori_n826_), .Y(ori_ori_n827_));
  NA3        o0799(.A(m), .B(l), .C(i), .Y(ori_ori_n828_));
  OAI220     o0800(.A0(ori_ori_n588_), .A1(ori_ori_n828_), .B0(ori_ori_n344_), .B1(ori_ori_n526_), .Y(ori_ori_n829_));
  NA4        o0801(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(g), .D(f), .Y(ori_ori_n830_));
  NAi31      o0802(.An(ori_ori_n829_), .B(ori_ori_n830_), .C(ori_ori_n432_), .Y(ori_ori_n831_));
  NA3        o0803(.A(ori_ori_n798_), .B(ori_ori_n564_), .C(ori_ori_n518_), .Y(ori_ori_n832_));
  OA210      o0804(.A0(ori_ori_n832_), .A1(ori_ori_n831_), .B0(ori_ori_n801_), .Y(ori_ori_n833_));
  INV        o0805(.A(ori_ori_n328_), .Y(ori_ori_n834_));
  NO2        o0806(.A(ori_ori_n125_), .B(ori_ori_n123_), .Y(ori_ori_n835_));
  NOi31      o0807(.An(k), .B(m), .C(l), .Y(ori_ori_n836_));
  NO2        o0808(.A(ori_ori_n330_), .B(ori_ori_n836_), .Y(ori_ori_n837_));
  AOI210     o0809(.A0(ori_ori_n837_), .A1(ori_ori_n835_), .B0(ori_ori_n594_), .Y(ori_ori_n838_));
  NA2        o0810(.A(ori_ori_n787_), .B(ori_ori_n321_), .Y(ori_ori_n839_));
  NA2        o0811(.A(ori_ori_n332_), .B(ori_ori_n334_), .Y(ori_ori_n840_));
  OAI210     o0812(.A0(ori_ori_n199_), .A1(ori_ori_n209_), .B0(ori_ori_n840_), .Y(ori_ori_n841_));
  AOI220     o0813(.A0(ori_ori_n841_), .A1(ori_ori_n839_), .B0(ori_ori_n838_), .B1(ori_ori_n834_), .Y(ori_ori_n842_));
  NA2        o0814(.A(ori_ori_n164_), .B(ori_ori_n112_), .Y(ori_ori_n843_));
  NA3        o0815(.A(ori_ori_n843_), .B(ori_ori_n695_), .C(ori_ori_n133_), .Y(ori_ori_n844_));
  NA3        o0816(.A(ori_ori_n844_), .B(ori_ori_n184_), .C(ori_ori_n31_), .Y(ori_ori_n845_));
  NA4        o0817(.A(ori_ori_n845_), .B(ori_ori_n842_), .C(ori_ori_n618_), .D(ori_ori_n78_), .Y(ori_ori_n846_));
  NO2        o0818(.A(ori_ori_n584_), .B(ori_ori_n495_), .Y(ori_ori_n847_));
  NA2        o0819(.A(ori_ori_n847_), .B(ori_ori_n184_), .Y(ori_ori_n848_));
  NOi21      o0820(.An(f), .B(d), .Y(ori_ori_n849_));
  NA2        o0821(.A(ori_ori_n849_), .B(m), .Y(ori_ori_n850_));
  NO2        o0822(.A(ori_ori_n850_), .B(ori_ori_n52_), .Y(ori_ori_n851_));
  NOi32      o0823(.An(g), .Bn(f), .C(d), .Y(ori_ori_n852_));
  NA4        o0824(.A(ori_ori_n852_), .B(ori_ori_n598_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n853_));
  NOi21      o0825(.An(ori_ori_n300_), .B(ori_ori_n853_), .Y(ori_ori_n854_));
  AOI210     o0826(.A0(ori_ori_n851_), .A1(ori_ori_n541_), .B0(ori_ori_n854_), .Y(ori_ori_n855_));
  NA3        o0827(.A(ori_ori_n299_), .B(ori_ori_n258_), .C(ori_ori_n117_), .Y(ori_ori_n856_));
  AN2        o0828(.A(f), .B(d), .Y(ori_ori_n857_));
  NA3        o0829(.A(ori_ori_n474_), .B(ori_ori_n857_), .C(ori_ori_n80_), .Y(ori_ori_n858_));
  NO3        o0830(.A(ori_ori_n858_), .B(ori_ori_n69_), .C(ori_ori_n210_), .Y(ori_ori_n859_));
  NA2        o0831(.A(ori_ori_n856_), .B(ori_ori_n859_), .Y(ori_ori_n860_));
  NAi41      o0832(.An(ori_ori_n488_), .B(ori_ori_n860_), .C(ori_ori_n855_), .D(ori_ori_n848_), .Y(ori_ori_n861_));
  NO4        o0833(.A(ori_ori_n616_), .B(ori_ori_n129_), .C(ori_ori_n316_), .D(ori_ori_n150_), .Y(ori_ori_n862_));
  NO2        o0834(.A(ori_ori_n649_), .B(ori_ori_n316_), .Y(ori_ori_n863_));
  AN2        o0835(.A(ori_ori_n863_), .B(ori_ori_n676_), .Y(ori_ori_n864_));
  NO2        o0836(.A(ori_ori_n864_), .B(ori_ori_n862_), .Y(ori_ori_n865_));
  NA3        o0837(.A(ori_ori_n158_), .B(ori_ori_n106_), .C(ori_ori_n105_), .Y(ori_ori_n866_));
  OAI220     o0838(.A0(ori_ori_n858_), .A1(ori_ori_n422_), .B0(ori_ori_n328_), .B1(ori_ori_n866_), .Y(ori_ori_n867_));
  NOi31      o0839(.An(ori_ori_n220_), .B(ori_ori_n867_), .C(ori_ori_n295_), .Y(ori_ori_n868_));
  NA2        o0840(.A(c), .B(ori_ori_n114_), .Y(ori_ori_n869_));
  NO2        o0841(.A(ori_ori_n869_), .B(ori_ori_n400_), .Y(ori_ori_n870_));
  NA3        o0842(.A(ori_ori_n870_), .B(ori_ori_n507_), .C(f), .Y(ori_ori_n871_));
  OR2        o0843(.A(ori_ori_n656_), .B(ori_ori_n537_), .Y(ori_ori_n872_));
  INV        o0844(.A(ori_ori_n872_), .Y(ori_ori_n873_));
  NA2        o0845(.A(ori_ori_n800_), .B(ori_ori_n109_), .Y(ori_ori_n874_));
  NA2        o0846(.A(ori_ori_n874_), .B(ori_ori_n873_), .Y(ori_ori_n875_));
  NA4        o0847(.A(ori_ori_n875_), .B(ori_ori_n871_), .C(ori_ori_n868_), .D(ori_ori_n865_), .Y(ori_ori_n876_));
  NO4        o0848(.A(ori_ori_n876_), .B(ori_ori_n861_), .C(ori_ori_n846_), .D(ori_ori_n833_), .Y(ori_ori_n877_));
  OR2        o0849(.A(ori_ori_n858_), .B(ori_ori_n69_), .Y(ori_ori_n878_));
  NA2        o0850(.A(ori_ori_n110_), .B(j), .Y(ori_ori_n879_));
  NA2        o0851(.A(ori_ori_n820_), .B(g), .Y(ori_ori_n880_));
  AOI210     o0852(.A0(ori_ori_n880_), .A1(ori_ori_n283_), .B0(ori_ori_n878_), .Y(ori_ori_n881_));
  NO2        o0853(.A(ori_ori_n321_), .B(ori_ori_n830_), .Y(ori_ori_n882_));
  NO2        o0854(.A(ori_ori_n133_), .B(ori_ori_n129_), .Y(ori_ori_n883_));
  NO2        o0855(.A(ori_ori_n227_), .B(ori_ori_n221_), .Y(ori_ori_n884_));
  AOI220     o0856(.A0(ori_ori_n884_), .A1(ori_ori_n224_), .B0(ori_ori_n293_), .B1(ori_ori_n883_), .Y(ori_ori_n885_));
  NO2        o0857(.A(ori_ori_n422_), .B(ori_ori_n819_), .Y(ori_ori_n886_));
  NA2        o0858(.A(ori_ori_n886_), .B(ori_ori_n558_), .Y(ori_ori_n887_));
  NA2        o0859(.A(ori_ori_n887_), .B(ori_ori_n885_), .Y(ori_ori_n888_));
  NA2        o0860(.A(e), .B(d), .Y(ori_ori_n889_));
  OAI220     o0861(.A0(ori_ori_n889_), .A1(c), .B0(ori_ori_n311_), .B1(d), .Y(ori_ori_n890_));
  NA3        o0862(.A(ori_ori_n890_), .B(ori_ori_n449_), .C(ori_ori_n505_), .Y(ori_ori_n891_));
  AOI210     o0863(.A0(ori_ori_n513_), .A1(ori_ori_n175_), .B0(ori_ori_n227_), .Y(ori_ori_n892_));
  AOI210     o0864(.A0(ori_ori_n617_), .A1(ori_ori_n337_), .B0(ori_ori_n892_), .Y(ori_ori_n893_));
  NA2        o0865(.A(ori_ori_n275_), .B(ori_ori_n162_), .Y(ori_ori_n894_));
  NA2        o0866(.A(ori_ori_n859_), .B(ori_ori_n894_), .Y(ori_ori_n895_));
  NA3        o0867(.A(ori_ori_n163_), .B(ori_ori_n81_), .C(ori_ori_n34_), .Y(ori_ori_n896_));
  NA4        o0868(.A(ori_ori_n896_), .B(ori_ori_n895_), .C(ori_ori_n893_), .D(ori_ori_n891_), .Y(ori_ori_n897_));
  NO4        o0869(.A(ori_ori_n897_), .B(ori_ori_n888_), .C(ori_ori_n882_), .D(ori_ori_n881_), .Y(ori_ori_n898_));
  OR2        o0870(.A(ori_ori_n697_), .B(ori_ori_n213_), .Y(ori_ori_n899_));
  OAI220     o0871(.A0(ori_ori_n616_), .A1(ori_ori_n60_), .B0(ori_ori_n291_), .B1(j), .Y(ori_ori_n900_));
  AOI220     o0872(.A0(ori_ori_n900_), .A1(ori_ori_n863_), .B0(ori_ori_n608_), .B1(ori_ori_n615_), .Y(ori_ori_n901_));
  OAI210     o0873(.A0(ori_ori_n825_), .A1(ori_ori_n165_), .B0(ori_ori_n901_), .Y(ori_ori_n902_));
  OAI210     o0874(.A0(ori_ori_n820_), .A1(ori_ori_n894_), .B0(ori_ori_n852_), .Y(ori_ori_n903_));
  NO2        o0875(.A(ori_ori_n903_), .B(ori_ori_n599_), .Y(ori_ori_n904_));
  AOI210     o0876(.A0(ori_ori_n116_), .A1(ori_ori_n115_), .B0(ori_ori_n257_), .Y(ori_ori_n905_));
  NO2        o0877(.A(ori_ori_n905_), .B(ori_ori_n853_), .Y(ori_ori_n906_));
  AO210      o0878(.A0(ori_ori_n839_), .A1(ori_ori_n829_), .B0(ori_ori_n906_), .Y(ori_ori_n907_));
  NOi31      o0879(.An(ori_ori_n541_), .B(ori_ori_n850_), .C(ori_ori_n283_), .Y(ori_ori_n908_));
  NO4        o0880(.A(ori_ori_n908_), .B(ori_ori_n907_), .C(ori_ori_n904_), .D(ori_ori_n902_), .Y(ori_ori_n909_));
  AO220      o0881(.A0(ori_ori_n449_), .A1(ori_ori_n741_), .B0(ori_ori_n170_), .B1(f), .Y(ori_ori_n910_));
  OAI210     o0882(.A0(ori_ori_n910_), .A1(ori_ori_n452_), .B0(ori_ori_n890_), .Y(ori_ori_n911_));
  NO2        o0883(.A(ori_ori_n431_), .B(ori_ori_n66_), .Y(ori_ori_n912_));
  OAI210     o0884(.A0(ori_ori_n832_), .A1(ori_ori_n912_), .B0(ori_ori_n701_), .Y(ori_ori_n913_));
  AN4        o0885(.A(ori_ori_n913_), .B(ori_ori_n911_), .C(ori_ori_n909_), .D(ori_ori_n899_), .Y(ori_ori_n914_));
  NA4        o0886(.A(ori_ori_n914_), .B(ori_ori_n898_), .C(ori_ori_n877_), .D(ori_ori_n827_), .Y(ori12));
  NO2        o0887(.A(ori_ori_n447_), .B(c), .Y(ori_ori_n916_));
  NO4        o0888(.A(ori_ori_n436_), .B(ori_ori_n249_), .C(ori_ori_n580_), .D(ori_ori_n210_), .Y(ori_ori_n917_));
  NA2        o0889(.A(ori_ori_n917_), .B(ori_ori_n916_), .Y(ori_ori_n918_));
  NA2        o0890(.A(ori_ori_n541_), .B(ori_ori_n912_), .Y(ori_ori_n919_));
  NO2        o0891(.A(ori_ori_n447_), .B(ori_ori_n114_), .Y(ori_ori_n920_));
  NO2        o0892(.A(ori_ori_n835_), .B(ori_ori_n344_), .Y(ori_ori_n921_));
  NO2        o0893(.A(ori_ori_n656_), .B(ori_ori_n369_), .Y(ori_ori_n922_));
  AOI220     o0894(.A0(ori_ori_n922_), .A1(ori_ori_n539_), .B0(ori_ori_n921_), .B1(ori_ori_n920_), .Y(ori_ori_n923_));
  NA4        o0895(.A(ori_ori_n923_), .B(ori_ori_n919_), .C(ori_ori_n918_), .D(ori_ori_n435_), .Y(ori_ori_n924_));
  AOI210     o0896(.A0(ori_ori_n230_), .A1(ori_ori_n327_), .B0(ori_ori_n196_), .Y(ori_ori_n925_));
  OR2        o0897(.A(ori_ori_n925_), .B(ori_ori_n917_), .Y(ori_ori_n926_));
  AOI210     o0898(.A0(ori_ori_n324_), .A1(ori_ori_n381_), .B0(ori_ori_n210_), .Y(ori_ori_n927_));
  OAI210     o0899(.A0(ori_ori_n927_), .A1(ori_ori_n926_), .B0(ori_ori_n395_), .Y(ori_ori_n928_));
  NO2        o0900(.A(ori_ori_n635_), .B(ori_ori_n259_), .Y(ori_ori_n929_));
  NO2        o0901(.A(ori_ori_n588_), .B(ori_ori_n828_), .Y(ori_ori_n930_));
  NO2        o0902(.A(ori_ori_n149_), .B(ori_ori_n233_), .Y(ori_ori_n931_));
  NA3        o0903(.A(ori_ori_n931_), .B(ori_ori_n236_), .C(i), .Y(ori_ori_n932_));
  NA2        o0904(.A(ori_ori_n932_), .B(ori_ori_n928_), .Y(ori_ori_n933_));
  OR2        o0905(.A(ori_ori_n312_), .B(ori_ori_n920_), .Y(ori_ori_n934_));
  NA2        o0906(.A(ori_ori_n934_), .B(ori_ori_n345_), .Y(ori_ori_n935_));
  NO3        o0907(.A(ori_ori_n129_), .B(ori_ori_n150_), .C(ori_ori_n210_), .Y(ori_ori_n936_));
  NA2        o0908(.A(ori_ori_n936_), .B(ori_ori_n530_), .Y(ori_ori_n937_));
  NA4        o0909(.A(ori_ori_n437_), .B(ori_ori_n429_), .C(ori_ori_n176_), .D(g), .Y(ori_ori_n938_));
  NA3        o0910(.A(ori_ori_n938_), .B(ori_ori_n937_), .C(ori_ori_n935_), .Y(ori_ori_n939_));
  NO3        o0911(.A(ori_ori_n659_), .B(ori_ori_n88_), .C(ori_ori_n45_), .Y(ori_ori_n940_));
  NO4        o0912(.A(ori_ori_n940_), .B(ori_ori_n939_), .C(ori_ori_n933_), .D(ori_ori_n924_), .Y(ori_ori_n941_));
  NO2        o0913(.A(ori_ori_n361_), .B(ori_ori_n360_), .Y(ori_ori_n942_));
  INV        o0914(.A(ori_ori_n68_), .Y(ori_ori_n943_));
  NA2        o0915(.A(ori_ori_n551_), .B(ori_ori_n142_), .Y(ori_ori_n944_));
  NOi21      o0916(.An(ori_ori_n34_), .B(ori_ori_n649_), .Y(ori_ori_n945_));
  AOI220     o0917(.A0(ori_ori_n945_), .A1(ori_ori_n944_), .B0(ori_ori_n943_), .B1(ori_ori_n942_), .Y(ori_ori_n946_));
  OAI210     o0918(.A0(ori_ori_n247_), .A1(ori_ori_n45_), .B0(ori_ori_n946_), .Y(ori_ori_n947_));
  INV        o0919(.A(ori_ori_n309_), .Y(ori_ori_n948_));
  NO2        o0920(.A(ori_ori_n49_), .B(ori_ori_n45_), .Y(ori_ori_n949_));
  NO2        o0921(.A(ori_ori_n502_), .B(ori_ori_n291_), .Y(ori_ori_n950_));
  INV        o0922(.A(ori_ori_n950_), .Y(ori_ori_n951_));
  NO2        o0923(.A(ori_ori_n951_), .B(ori_ori_n142_), .Y(ori_ori_n952_));
  INV        o0924(.A(ori_ori_n358_), .Y(ori_ori_n953_));
  NO4        o0925(.A(ori_ori_n953_), .B(ori_ori_n952_), .C(ori_ori_n948_), .D(ori_ori_n947_), .Y(ori_ori_n954_));
  NA2        o0926(.A(ori_ori_n337_), .B(g), .Y(ori_ori_n955_));
  NA2        o0927(.A(ori_ori_n161_), .B(i), .Y(ori_ori_n956_));
  NA2        o0928(.A(ori_ori_n46_), .B(i), .Y(ori_ori_n957_));
  OAI220     o0929(.A0(ori_ori_n957_), .A1(ori_ori_n195_), .B0(ori_ori_n956_), .B1(ori_ori_n88_), .Y(ori_ori_n958_));
  AOI210     o0930(.A0(ori_ori_n411_), .A1(ori_ori_n37_), .B0(ori_ori_n958_), .Y(ori_ori_n959_));
  NO2        o0931(.A(ori_ori_n142_), .B(ori_ori_n80_), .Y(ori_ori_n960_));
  OR2        o0932(.A(ori_ori_n960_), .B(ori_ori_n550_), .Y(ori_ori_n961_));
  NA2        o0933(.A(ori_ori_n551_), .B(ori_ori_n373_), .Y(ori_ori_n962_));
  AOI210     o0934(.A0(ori_ori_n962_), .A1(n), .B0(ori_ori_n961_), .Y(ori_ori_n963_));
  OAI220     o0935(.A0(ori_ori_n963_), .A1(ori_ori_n955_), .B0(ori_ori_n959_), .B1(ori_ori_n321_), .Y(ori_ori_n964_));
  NO2        o0936(.A(ori_ori_n656_), .B(ori_ori_n495_), .Y(ori_ori_n965_));
  NA3        o0937(.A(ori_ori_n332_), .B(ori_ori_n622_), .C(i), .Y(ori_ori_n966_));
  OAI210     o0938(.A0(ori_ori_n431_), .A1(ori_ori_n299_), .B0(ori_ori_n966_), .Y(ori_ori_n967_));
  OAI220     o0939(.A0(ori_ori_n967_), .A1(ori_ori_n965_), .B0(ori_ori_n672_), .B1(ori_ori_n751_), .Y(ori_ori_n968_));
  NA2        o0940(.A(ori_ori_n602_), .B(ori_ori_n111_), .Y(ori_ori_n969_));
  OR3        o0941(.A(ori_ori_n299_), .B(ori_ori_n427_), .C(f), .Y(ori_ori_n970_));
  NA3        o0942(.A(ori_ori_n622_), .B(ori_ori_n76_), .C(i), .Y(ori_ori_n971_));
  OA220      o0943(.A0(ori_ori_n971_), .A1(ori_ori_n969_), .B0(ori_ori_n970_), .B1(ori_ori_n587_), .Y(ori_ori_n972_));
  NA3        o0944(.A(ori_ori_n313_), .B(ori_ori_n116_), .C(g), .Y(ori_ori_n973_));
  AOI210     o0945(.A0(ori_ori_n669_), .A1(ori_ori_n973_), .B0(m), .Y(ori_ori_n974_));
  OAI210     o0946(.A0(ori_ori_n974_), .A1(ori_ori_n921_), .B0(ori_ori_n312_), .Y(ori_ori_n975_));
  INV        o0947(.A(ori_ori_n688_), .Y(ori_ori_n976_));
  NA2        o0948(.A(ori_ori_n830_), .B(ori_ori_n432_), .Y(ori_ori_n977_));
  NA2        o0949(.A(ori_ori_n218_), .B(ori_ori_n73_), .Y(ori_ori_n978_));
  NA2        o0950(.A(ori_ori_n978_), .B(ori_ori_n971_), .Y(ori_ori_n979_));
  AOI220     o0951(.A0(ori_ori_n979_), .A1(ori_ori_n255_), .B0(ori_ori_n977_), .B1(ori_ori_n976_), .Y(ori_ori_n980_));
  NA4        o0952(.A(ori_ori_n980_), .B(ori_ori_n975_), .C(ori_ori_n972_), .D(ori_ori_n968_), .Y(ori_ori_n981_));
  NO2        o0953(.A(ori_ori_n369_), .B(ori_ori_n87_), .Y(ori_ori_n982_));
  OAI210     o0954(.A0(ori_ori_n982_), .A1(ori_ori_n929_), .B0(ori_ori_n234_), .Y(ori_ori_n983_));
  NA2        o0955(.A(ori_ori_n658_), .B(ori_ori_n84_), .Y(ori_ori_n984_));
  NO2        o0956(.A(ori_ori_n455_), .B(ori_ori_n210_), .Y(ori_ori_n985_));
  AOI220     o0957(.A0(ori_ori_n985_), .A1(ori_ori_n374_), .B0(ori_ori_n934_), .B1(ori_ori_n214_), .Y(ori_ori_n986_));
  AOI220     o0958(.A0(ori_ori_n922_), .A1(ori_ori_n931_), .B0(ori_ori_n586_), .B1(ori_ori_n86_), .Y(ori_ori_n987_));
  NA4        o0959(.A(ori_ori_n987_), .B(ori_ori_n986_), .C(ori_ori_n984_), .D(ori_ori_n983_), .Y(ori_ori_n988_));
  OAI210     o0960(.A0(ori_ori_n977_), .A1(ori_ori_n930_), .B0(ori_ori_n539_), .Y(ori_ori_n989_));
  OAI210     o0961(.A0(ori_ori_n361_), .A1(ori_ori_n360_), .B0(ori_ori_n107_), .Y(ori_ori_n990_));
  NA2        o0962(.A(ori_ori_n990_), .B(ori_ori_n533_), .Y(ori_ori_n991_));
  NA2        o0963(.A(ori_ori_n974_), .B(ori_ori_n920_), .Y(ori_ori_n992_));
  NO3        o0964(.A(ori_ori_n879_), .B(ori_ori_n49_), .C(ori_ori_n45_), .Y(ori_ori_n993_));
  AOI220     o0965(.A0(ori_ori_n993_), .A1(ori_ori_n620_), .B0(ori_ori_n640_), .B1(ori_ori_n530_), .Y(ori_ori_n994_));
  NA4        o0966(.A(ori_ori_n994_), .B(ori_ori_n992_), .C(ori_ori_n991_), .D(ori_ori_n989_), .Y(ori_ori_n995_));
  NO4        o0967(.A(ori_ori_n995_), .B(ori_ori_n988_), .C(ori_ori_n981_), .D(ori_ori_n964_), .Y(ori_ori_n996_));
  NAi31      o0968(.An(ori_ori_n138_), .B(ori_ori_n413_), .C(n), .Y(ori_ori_n997_));
  NO3        o0969(.A(ori_ori_n123_), .B(ori_ori_n330_), .C(ori_ori_n836_), .Y(ori_ori_n998_));
  NO2        o0970(.A(ori_ori_n998_), .B(ori_ori_n997_), .Y(ori_ori_n999_));
  NO3        o0971(.A(ori_ori_n267_), .B(ori_ori_n138_), .C(ori_ori_n400_), .Y(ori_ori_n1000_));
  AOI210     o0972(.A0(ori_ori_n1000_), .A1(ori_ori_n496_), .B0(ori_ori_n999_), .Y(ori_ori_n1001_));
  NA2        o0973(.A(ori_ori_n489_), .B(i), .Y(ori_ori_n1002_));
  NA2        o0974(.A(ori_ori_n1002_), .B(ori_ori_n1001_), .Y(ori_ori_n1003_));
  NA2        o0975(.A(ori_ori_n227_), .B(ori_ori_n166_), .Y(ori_ori_n1004_));
  NO3        o0976(.A(ori_ori_n297_), .B(ori_ori_n437_), .C(ori_ori_n170_), .Y(ori_ori_n1005_));
  NOi31      o0977(.An(ori_ori_n1004_), .B(ori_ori_n1005_), .C(ori_ori_n210_), .Y(ori_ori_n1006_));
  NAi21      o0978(.An(ori_ori_n551_), .B(ori_ori_n985_), .Y(ori_ori_n1007_));
  NA2        o0979(.A(ori_ori_n480_), .B(g), .Y(ori_ori_n1008_));
  NA2        o0980(.A(ori_ori_n1008_), .B(ori_ori_n1007_), .Y(ori_ori_n1009_));
  NA2        o0981(.A(ori_ori_n925_), .B(ori_ori_n916_), .Y(ori_ori_n1010_));
  OAI220     o0982(.A0(ori_ori_n922_), .A1(ori_ori_n930_), .B0(ori_ori_n541_), .B1(ori_ori_n421_), .Y(ori_ori_n1011_));
  NA3        o0983(.A(ori_ori_n1011_), .B(ori_ori_n1010_), .C(ori_ori_n614_), .Y(ori_ori_n1012_));
  OAI210     o0984(.A0(ori_ori_n925_), .A1(ori_ori_n917_), .B0(ori_ori_n1004_), .Y(ori_ori_n1013_));
  NA3        o0985(.A(ori_ori_n962_), .B(ori_ori_n485_), .C(ori_ori_n46_), .Y(ori_ori_n1014_));
  AOI210     o0986(.A0(ori_ori_n372_), .A1(ori_ori_n370_), .B0(ori_ori_n320_), .Y(ori_ori_n1015_));
  NA3        o0987(.A(ori_ori_n1015_), .B(ori_ori_n1014_), .C(ori_ori_n1013_), .Y(ori_ori_n1016_));
  OR2        o0988(.A(ori_ori_n1016_), .B(ori_ori_n1012_), .Y(ori_ori_n1017_));
  NO4        o0989(.A(ori_ori_n1017_), .B(ori_ori_n1009_), .C(ori_ori_n1006_), .D(ori_ori_n1003_), .Y(ori_ori_n1018_));
  NA4        o0990(.A(ori_ori_n1018_), .B(ori_ori_n996_), .C(ori_ori_n954_), .D(ori_ori_n941_), .Y(ori13));
  AN2        o0991(.A(c), .B(b), .Y(ori_ori_n1020_));
  NAi32      o0992(.An(d), .Bn(c), .C(e), .Y(ori_ori_n1021_));
  AN2        o0993(.A(d), .B(c), .Y(ori_ori_n1022_));
  NA2        o0994(.A(ori_ori_n1022_), .B(ori_ori_n114_), .Y(ori_ori_n1023_));
  NO3        o0995(.A(m), .B(i), .C(h), .Y(ori_ori_n1024_));
  NA3        o0996(.A(k), .B(j), .C(i), .Y(ori_ori_n1025_));
  AN3        o0997(.A(g), .B(f), .C(c), .Y(ori_ori_n1026_));
  NA3        o0998(.A(l), .B(k), .C(j), .Y(ori_ori_n1027_));
  NA2        o0999(.A(i), .B(h), .Y(ori_ori_n1028_));
  NO3        o1000(.A(ori_ori_n1028_), .B(ori_ori_n1027_), .C(ori_ori_n129_), .Y(ori_ori_n1029_));
  NO3        o1001(.A(ori_ori_n139_), .B(ori_ori_n274_), .C(ori_ori_n210_), .Y(ori_ori_n1030_));
  NA3        o1002(.A(c), .B(b), .C(a), .Y(ori_ori_n1031_));
  NO2        o1003(.A(ori_ori_n526_), .B(ori_ori_n594_), .Y(ori_ori_n1032_));
  NA4        o1004(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(g), .D(ori_ori_n209_), .Y(ori_ori_n1033_));
  NA4        o1005(.A(ori_ori_n572_), .B(m), .C(ori_ori_n110_), .D(ori_ori_n209_), .Y(ori_ori_n1034_));
  NA3        o1006(.A(ori_ori_n1034_), .B(ori_ori_n362_), .C(ori_ori_n1033_), .Y(ori_ori_n1035_));
  NO3        o1007(.A(ori_ori_n1035_), .B(ori_ori_n1032_), .C(ori_ori_n990_), .Y(ori_ori_n1036_));
  NOi41      o1008(.An(ori_ori_n798_), .B(ori_ori_n841_), .C(ori_ori_n831_), .D(ori_ori_n715_), .Y(ori_ori_n1037_));
  OAI220     o1009(.A0(ori_ori_n1037_), .A1(ori_ori_n688_), .B0(ori_ori_n1036_), .B1(ori_ori_n585_), .Y(ori_ori_n1038_));
  NOi31      o1010(.An(m), .B(n), .C(f), .Y(ori_ori_n1039_));
  NA2        o1011(.A(ori_ori_n1039_), .B(ori_ori_n51_), .Y(ori_ori_n1040_));
  AN2        o1012(.A(e), .B(c), .Y(ori_ori_n1041_));
  NA2        o1013(.A(ori_ori_n1041_), .B(a), .Y(ori_ori_n1042_));
  OAI220     o1014(.A0(ori_ori_n1042_), .A1(ori_ori_n1040_), .B0(ori_ori_n872_), .B1(ori_ori_n420_), .Y(ori_ori_n1043_));
  NA2        o1015(.A(ori_ori_n505_), .B(l), .Y(ori_ori_n1044_));
  NO2        o1016(.A(ori_ori_n274_), .B(a), .Y(ori_ori_n1045_));
  NO2        o1017(.A(ori_ori_n83_), .B(g), .Y(ori_ori_n1046_));
  NO4        o1018(.A(ori_ori_n1043_), .B(ori_ori_n1038_), .C(ori_ori_n811_), .D(ori_ori_n562_), .Y(ori_ori_n1047_));
  NA2        o1019(.A(c), .B(b), .Y(ori_ori_n1048_));
  NO2        o1020(.A(ori_ori_n700_), .B(ori_ori_n1048_), .Y(ori_ori_n1049_));
  OAI210     o1021(.A0(ori_ori_n850_), .A1(ori_ori_n823_), .B0(ori_ori_n407_), .Y(ori_ori_n1050_));
  OAI210     o1022(.A0(ori_ori_n1050_), .A1(ori_ori_n851_), .B0(ori_ori_n1049_), .Y(ori_ori_n1051_));
  NAi21      o1023(.An(ori_ori_n415_), .B(ori_ori_n1049_), .Y(ori_ori_n1052_));
  NA3        o1024(.A(ori_ori_n421_), .B(ori_ori_n556_), .C(f), .Y(ori_ori_n1053_));
  OAI210     o1025(.A0(ori_ori_n545_), .A1(ori_ori_n39_), .B0(ori_ori_n1045_), .Y(ori_ori_n1054_));
  NA3        o1026(.A(ori_ori_n1054_), .B(ori_ori_n1053_), .C(ori_ori_n1052_), .Y(ori_ori_n1055_));
  NA2        o1027(.A(ori_ori_n258_), .B(ori_ori_n117_), .Y(ori_ori_n1056_));
  OAI210     o1028(.A0(ori_ori_n1056_), .A1(ori_ori_n277_), .B0(g), .Y(ori_ori_n1057_));
  NAi21      o1029(.An(f), .B(d), .Y(ori_ori_n1058_));
  NO2        o1030(.A(ori_ori_n1058_), .B(ori_ori_n1031_), .Y(ori_ori_n1059_));
  INV        o1031(.A(ori_ori_n1059_), .Y(ori_ori_n1060_));
  AOI210     o1032(.A0(ori_ori_n1057_), .A1(ori_ori_n283_), .B0(ori_ori_n1060_), .Y(ori_ori_n1061_));
  AOI210     o1033(.A0(ori_ori_n1061_), .A1(ori_ori_n111_), .B0(ori_ori_n1055_), .Y(ori_ori_n1062_));
  NA3        o1034(.A(ori_ori_n905_), .B(ori_ori_n1044_), .C(ori_ori_n469_), .Y(ori_ori_n1063_));
  NA2        o1035(.A(ori_ori_n440_), .B(ori_ori_n1059_), .Y(ori_ori_n1064_));
  NA4        o1036(.A(ori_ori_n1064_), .B(ori_ori_n1062_), .C(ori_ori_n1051_), .D(ori_ori_n1047_), .Y(ori00));
  NA2        o1037(.A(ori_ori_n886_), .B(ori_ori_n931_), .Y(ori_ori_n1066_));
  INV        o1038(.A(ori_ori_n712_), .Y(ori_ori_n1067_));
  NA3        o1039(.A(ori_ori_n1067_), .B(ori_ori_n1066_), .C(ori_ori_n991_), .Y(ori_ori_n1068_));
  NA2        o1040(.A(ori_ori_n507_), .B(f), .Y(ori_ori_n1069_));
  OAI210     o1041(.A0(ori_ori_n998_), .A1(ori_ori_n40_), .B0(ori_ori_n642_), .Y(ori_ori_n1070_));
  NA3        o1042(.A(ori_ori_n1070_), .B(ori_ori_n254_), .C(n), .Y(ori_ori_n1071_));
  AOI210     o1043(.A0(ori_ori_n1071_), .A1(ori_ori_n1069_), .B0(ori_ori_n1023_), .Y(ori_ori_n1072_));
  NO2        o1044(.A(ori_ori_n1072_), .B(ori_ori_n1068_), .Y(ori_ori_n1073_));
  NA3        o1045(.A(ori_ori_n163_), .B(ori_ori_n46_), .C(ori_ori_n45_), .Y(ori_ori_n1074_));
  NA3        o1046(.A(d), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n1075_));
  NO2        o1047(.A(ori_ori_n1075_), .B(ori_ori_n1074_), .Y(ori_ori_n1076_));
  INV        o1048(.A(ori_ori_n574_), .Y(ori_ori_n1077_));
  NO3        o1049(.A(ori_ori_n1077_), .B(ori_ori_n1076_), .C(ori_ori_n908_), .Y(ori_ori_n1078_));
  NO4        o1050(.A(ori_ori_n486_), .B(ori_ori_n347_), .C(ori_ori_n1048_), .D(ori_ori_n59_), .Y(ori_ori_n1079_));
  NA3        o1051(.A(ori_ori_n375_), .B(ori_ori_n217_), .C(g), .Y(ori_ori_n1080_));
  OR2        o1052(.A(ori_ori_n1080_), .B(ori_ori_n1075_), .Y(ori_ori_n1081_));
  NO2        o1053(.A(h), .B(g), .Y(ori_ori_n1082_));
  NA4        o1054(.A(ori_ori_n496_), .B(ori_ori_n463_), .C(ori_ori_n1082_), .D(ori_ori_n1020_), .Y(ori_ori_n1083_));
  OAI220     o1055(.A0(ori_ori_n526_), .A1(ori_ori_n594_), .B0(ori_ori_n88_), .B1(ori_ori_n87_), .Y(ori_ori_n1084_));
  AOI220     o1056(.A0(ori_ori_n1084_), .A1(ori_ori_n533_), .B0(ori_ori_n936_), .B1(ori_ori_n573_), .Y(ori_ori_n1085_));
  AOI220     o1057(.A0(ori_ori_n306_), .A1(ori_ori_n243_), .B0(ori_ori_n172_), .B1(ori_ori_n146_), .Y(ori_ori_n1086_));
  NA4        o1058(.A(ori_ori_n1086_), .B(ori_ori_n1085_), .C(ori_ori_n1083_), .D(ori_ori_n1081_), .Y(ori_ori_n1087_));
  NO3        o1059(.A(ori_ori_n1087_), .B(ori_ori_n1079_), .C(ori_ori_n262_), .Y(ori_ori_n1088_));
  AOI210     o1060(.A0(ori_ori_n243_), .A1(ori_ori_n337_), .B0(ori_ori_n576_), .Y(ori_ori_n1089_));
  NA2        o1061(.A(ori_ori_n1089_), .B(ori_ori_n152_), .Y(ori_ori_n1090_));
  NO2        o1062(.A(ori_ori_n235_), .B(ori_ori_n176_), .Y(ori_ori_n1091_));
  NA2        o1063(.A(ori_ori_n1091_), .B(ori_ori_n421_), .Y(ori_ori_n1092_));
  INV        o1064(.A(ori_ori_n1092_), .Y(ori_ori_n1093_));
  NO2        o1065(.A(ori_ori_n269_), .B(ori_ori_n69_), .Y(ori_ori_n1094_));
  NO3        o1066(.A(ori_ori_n420_), .B(ori_ori_n819_), .C(n), .Y(ori_ori_n1095_));
  NA2        o1067(.A(ori_ori_n1095_), .B(ori_ori_n1094_), .Y(ori_ori_n1096_));
  INV        o1068(.A(ori_ori_n1096_), .Y(ori_ori_n1097_));
  NO4        o1069(.A(ori_ori_n1097_), .B(ori_ori_n1093_), .C(ori_ori_n1090_), .D(ori_ori_n517_), .Y(ori_ori_n1098_));
  AN3        o1070(.A(ori_ori_n1098_), .B(ori_ori_n1088_), .C(ori_ori_n1078_), .Y(ori_ori_n1099_));
  NA2        o1071(.A(ori_ori_n533_), .B(ori_ori_n98_), .Y(ori_ori_n1100_));
  NA3        o1072(.A(ori_ori_n1039_), .B(ori_ori_n602_), .C(ori_ori_n462_), .Y(ori_ori_n1101_));
  NA3        o1073(.A(ori_ori_n1101_), .B(ori_ori_n1100_), .C(ori_ori_n237_), .Y(ori_ori_n1102_));
  NA2        o1074(.A(ori_ori_n1035_), .B(ori_ori_n533_), .Y(ori_ori_n1103_));
  NA4        o1075(.A(ori_ori_n645_), .B(ori_ori_n201_), .C(ori_ori_n217_), .D(ori_ori_n161_), .Y(ori_ori_n1104_));
  NA3        o1076(.A(ori_ori_n1104_), .B(ori_ori_n1103_), .C(ori_ori_n287_), .Y(ori_ori_n1105_));
  OAI210     o1077(.A0(ori_ori_n461_), .A1(ori_ori_n118_), .B0(ori_ori_n853_), .Y(ori_ori_n1106_));
  NA2        o1078(.A(ori_ori_n1106_), .B(ori_ori_n1063_), .Y(ori_ori_n1107_));
  NO2        o1079(.A(ori_ori_n213_), .B(ori_ori_n210_), .Y(ori_ori_n1108_));
  NA2        o1080(.A(n), .B(e), .Y(ori_ori_n1109_));
  NO2        o1081(.A(ori_ori_n1109_), .B(ori_ori_n144_), .Y(ori_ori_n1110_));
  AOI220     o1082(.A0(ori_ori_n1110_), .A1(ori_ori_n268_), .B0(ori_ori_n834_), .B1(ori_ori_n1108_), .Y(ori_ori_n1111_));
  OAI210     o1083(.A0(ori_ori_n348_), .A1(ori_ori_n301_), .B0(ori_ori_n442_), .Y(ori_ori_n1112_));
  NA3        o1084(.A(ori_ori_n1112_), .B(ori_ori_n1111_), .C(ori_ori_n1107_), .Y(ori_ori_n1113_));
  NA2        o1085(.A(ori_ori_n1110_), .B(ori_ori_n838_), .Y(ori_ori_n1114_));
  AOI220     o1086(.A0(ori_ori_n945_), .A1(ori_ori_n573_), .B0(ori_ori_n645_), .B1(ori_ori_n240_), .Y(ori_ori_n1115_));
  NO2        o1087(.A(ori_ori_n64_), .B(h), .Y(ori_ori_n1116_));
  NA3        o1088(.A(ori_ori_n1115_), .B(ori_ori_n1114_), .C(ori_ori_n855_), .Y(ori_ori_n1117_));
  NO4        o1089(.A(ori_ori_n1117_), .B(ori_ori_n1113_), .C(ori_ori_n1105_), .D(ori_ori_n1102_), .Y(ori_ori_n1118_));
  NA2        o1090(.A(ori_ori_n824_), .B(ori_ori_n750_), .Y(ori_ori_n1119_));
  NA4        o1091(.A(ori_ori_n1119_), .B(ori_ori_n1118_), .C(ori_ori_n1099_), .D(ori_ori_n1073_), .Y(ori01));
  NO2        o1092(.A(ori_ori_n477_), .B(ori_ori_n272_), .Y(ori_ori_n1121_));
  NA2        o1093(.A(ori_ori_n386_), .B(i), .Y(ori_ori_n1122_));
  NA3        o1094(.A(ori_ori_n1122_), .B(ori_ori_n1121_), .C(ori_ori_n1010_), .Y(ori_ori_n1123_));
  NA2        o1095(.A(ori_ori_n586_), .B(ori_ori_n86_), .Y(ori_ori_n1124_));
  NA2        o1096(.A(ori_ori_n551_), .B(ori_ori_n266_), .Y(ori_ori_n1125_));
  NA2        o1097(.A(ori_ori_n950_), .B(ori_ori_n1125_), .Y(ori_ori_n1126_));
  NA4        o1098(.A(ori_ori_n1126_), .B(ori_ori_n1124_), .C(ori_ori_n901_), .D(ori_ori_n322_), .Y(ori_ori_n1127_));
  NA2        o1099(.A(ori_ori_n45_), .B(f), .Y(ori_ori_n1128_));
  NA2        o1100(.A(ori_ori_n707_), .B(ori_ori_n93_), .Y(ori_ori_n1129_));
  NO2        o1101(.A(ori_ori_n1129_), .B(ori_ori_n1128_), .Y(ori_ori_n1130_));
  INV        o1102(.A(ori_ori_n116_), .Y(ori_ori_n1131_));
  OA220      o1103(.A0(ori_ori_n1131_), .A1(ori_ori_n583_), .B0(ori_ori_n657_), .B1(ori_ori_n362_), .Y(ori_ori_n1132_));
  NAi41      o1104(.An(ori_ori_n160_), .B(ori_ori_n1132_), .C(ori_ori_n1104_), .D(ori_ori_n885_), .Y(ori_ori_n1133_));
  NO3        o1105(.A(ori_ori_n778_), .B(ori_ori_n671_), .C(ori_ori_n510_), .Y(ori_ori_n1134_));
  NA4        o1106(.A(ori_ori_n707_), .B(ori_ori_n93_), .C(ori_ori_n45_), .D(ori_ori_n209_), .Y(ori_ori_n1135_));
  OA220      o1107(.A0(ori_ori_n1135_), .A1(ori_ori_n665_), .B0(ori_ori_n190_), .B1(ori_ori_n188_), .Y(ori_ori_n1136_));
  NA3        o1108(.A(ori_ori_n1136_), .B(ori_ori_n1134_), .C(ori_ori_n134_), .Y(ori_ori_n1137_));
  NO4        o1109(.A(ori_ori_n1137_), .B(ori_ori_n1133_), .C(ori_ori_n1127_), .D(ori_ori_n1123_), .Y(ori_ori_n1138_));
  INV        o1110(.A(ori_ori_n1080_), .Y(ori_ori_n1139_));
  NA2        o1111(.A(ori_ori_n1139_), .B(ori_ori_n530_), .Y(ori_ori_n1140_));
  NA2        o1112(.A(ori_ori_n535_), .B(ori_ori_n388_), .Y(ori_ori_n1141_));
  NOi21      o1113(.An(ori_ori_n559_), .B(ori_ori_n580_), .Y(ori_ori_n1142_));
  NA2        o1114(.A(ori_ori_n1142_), .B(ori_ori_n1141_), .Y(ori_ori_n1143_));
  AOI210     o1115(.A0(ori_ori_n199_), .A1(ori_ori_n85_), .B0(ori_ori_n209_), .Y(ori_ori_n1144_));
  OAI210     o1116(.A0(ori_ori_n801_), .A1(ori_ori_n421_), .B0(ori_ori_n1144_), .Y(ori_ori_n1145_));
  AN3        o1117(.A(m), .B(l), .C(k), .Y(ori_ori_n1146_));
  OAI210     o1118(.A0(ori_ori_n350_), .A1(ori_ori_n34_), .B0(ori_ori_n1146_), .Y(ori_ori_n1147_));
  NA2        o1119(.A(ori_ori_n198_), .B(ori_ori_n34_), .Y(ori_ori_n1148_));
  AO210      o1120(.A0(ori_ori_n1148_), .A1(ori_ori_n1147_), .B0(ori_ori_n321_), .Y(ori_ori_n1149_));
  NA4        o1121(.A(ori_ori_n1149_), .B(ori_ori_n1145_), .C(ori_ori_n1143_), .D(ori_ori_n1140_), .Y(ori_ori_n1150_));
  NA2        o1122(.A(ori_ori_n592_), .B(ori_ori_n116_), .Y(ori_ori_n1151_));
  OAI210     o1123(.A0(ori_ori_n1131_), .A1(ori_ori_n589_), .B0(ori_ori_n1151_), .Y(ori_ori_n1152_));
  NA2        o1124(.A(ori_ori_n271_), .B(ori_ori_n190_), .Y(ori_ori_n1153_));
  NA2        o1125(.A(ori_ori_n1153_), .B(ori_ori_n661_), .Y(ori_ori_n1154_));
  OAI210     o1126(.A0(ori_ori_n1130_), .A1(ori_ori_n315_), .B0(ori_ori_n672_), .Y(ori_ori_n1155_));
  NA3        o1127(.A(ori_ori_n1155_), .B(ori_ori_n1154_), .C(ori_ori_n781_), .Y(ori_ori_n1156_));
  NO3        o1128(.A(ori_ori_n1156_), .B(ori_ori_n1152_), .C(ori_ori_n1150_), .Y(ori_ori_n1157_));
  NA3        o1129(.A(ori_ori_n598_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1158_));
  NO2        o1130(.A(ori_ori_n1158_), .B(ori_ori_n199_), .Y(ori_ori_n1159_));
  AOI210     o1131(.A0(ori_ori_n503_), .A1(ori_ori_n58_), .B0(ori_ori_n1159_), .Y(ori_ori_n1160_));
  OR3        o1132(.A(ori_ori_n1129_), .B(ori_ori_n599_), .C(ori_ori_n1128_), .Y(ori_ori_n1161_));
  NO2        o1133(.A(ori_ori_n1135_), .B(ori_ori_n969_), .Y(ori_ori_n1162_));
  NO2        o1134(.A(ori_ori_n202_), .B(ori_ori_n109_), .Y(ori_ori_n1163_));
  NO3        o1135(.A(ori_ori_n1163_), .B(ori_ori_n1162_), .C(ori_ori_n1076_), .Y(ori_ori_n1164_));
  NA4        o1136(.A(ori_ori_n1164_), .B(ori_ori_n1161_), .C(ori_ori_n1160_), .D(ori_ori_n749_), .Y(ori_ori_n1165_));
  NO2        o1137(.A(ori_ori_n956_), .B(ori_ori_n229_), .Y(ori_ori_n1166_));
  NO2        o1138(.A(ori_ori_n957_), .B(ori_ori_n553_), .Y(ori_ori_n1167_));
  OAI210     o1139(.A0(ori_ori_n1167_), .A1(ori_ori_n1166_), .B0(ori_ori_n330_), .Y(ori_ori_n1168_));
  NA2        o1140(.A(ori_ori_n568_), .B(ori_ori_n566_), .Y(ori_ori_n1169_));
  NO3        o1141(.A(ori_ori_n75_), .B(ori_ori_n291_), .C(ori_ori_n45_), .Y(ori_ori_n1170_));
  NA2        o1142(.A(ori_ori_n1170_), .B(ori_ori_n550_), .Y(ori_ori_n1171_));
  NA3        o1143(.A(ori_ori_n1171_), .B(ori_ori_n1169_), .C(ori_ori_n667_), .Y(ori_ori_n1172_));
  OR2        o1144(.A(ori_ori_n1080_), .B(ori_ori_n1075_), .Y(ori_ori_n1173_));
  NO2        o1145(.A(ori_ori_n362_), .B(ori_ori_n68_), .Y(ori_ori_n1174_));
  INV        o1146(.A(ori_ori_n1174_), .Y(ori_ori_n1175_));
  NA2        o1147(.A(ori_ori_n1170_), .B(ori_ori_n804_), .Y(ori_ori_n1176_));
  NA4        o1148(.A(ori_ori_n1176_), .B(ori_ori_n1175_), .C(ori_ori_n1173_), .D(ori_ori_n378_), .Y(ori_ori_n1177_));
  NOi41      o1149(.An(ori_ori_n1168_), .B(ori_ori_n1177_), .C(ori_ori_n1172_), .D(ori_ori_n1165_), .Y(ori_ori_n1178_));
  NO2        o1150(.A(ori_ori_n128_), .B(ori_ori_n45_), .Y(ori_ori_n1179_));
  NO2        o1151(.A(ori_ori_n45_), .B(ori_ori_n40_), .Y(ori_ori_n1180_));
  AO220      o1152(.A0(ori_ori_n1180_), .A1(ori_ori_n617_), .B0(ori_ori_n1179_), .B1(ori_ori_n705_), .Y(ori_ori_n1181_));
  NA2        o1153(.A(ori_ori_n1181_), .B(ori_ori_n330_), .Y(ori_ori_n1182_));
  INV        o1154(.A(ori_ori_n132_), .Y(ori_ori_n1183_));
  NO3        o1155(.A(ori_ori_n1028_), .B(ori_ori_n171_), .C(ori_ori_n83_), .Y(ori_ori_n1184_));
  AOI220     o1156(.A0(ori_ori_n1184_), .A1(ori_ori_n1183_), .B0(ori_ori_n1170_), .B1(ori_ori_n960_), .Y(ori_ori_n1185_));
  NA2        o1157(.A(ori_ori_n1185_), .B(ori_ori_n1182_), .Y(ori_ori_n1186_));
  NO2        o1158(.A(ori_ori_n610_), .B(ori_ori_n609_), .Y(ori_ori_n1187_));
  NO4        o1159(.A(ori_ori_n1028_), .B(ori_ori_n1187_), .C(ori_ori_n169_), .D(ori_ori_n83_), .Y(ori_ori_n1188_));
  NO3        o1160(.A(ori_ori_n1188_), .B(ori_ori_n1186_), .C(ori_ori_n634_), .Y(ori_ori_n1189_));
  NA4        o1161(.A(ori_ori_n1189_), .B(ori_ori_n1178_), .C(ori_ori_n1157_), .D(ori_ori_n1138_), .Y(ori06));
  NO2        o1162(.A(ori_ori_n221_), .B(ori_ori_n100_), .Y(ori_ori_n1191_));
  OAI210     o1163(.A0(ori_ori_n1191_), .A1(ori_ori_n1184_), .B0(ori_ori_n374_), .Y(ori_ori_n1192_));
  NO3        o1164(.A(ori_ori_n595_), .B(ori_ori_n799_), .C(ori_ori_n596_), .Y(ori_ori_n1193_));
  OR2        o1165(.A(ori_ori_n1193_), .B(ori_ori_n872_), .Y(ori_ori_n1194_));
  NA3        o1166(.A(ori_ori_n1194_), .B(ori_ori_n1192_), .C(ori_ori_n1168_), .Y(ori_ori_n1195_));
  NO3        o1167(.A(ori_ori_n1195_), .B(ori_ori_n1172_), .C(ori_ori_n253_), .Y(ori_ori_n1196_));
  NO2        o1168(.A(ori_ori_n291_), .B(ori_ori_n45_), .Y(ori_ori_n1197_));
  AOI210     o1169(.A0(ori_ori_n1197_), .A1(ori_ori_n961_), .B0(ori_ori_n1166_), .Y(ori_ori_n1198_));
  AOI210     o1170(.A0(ori_ori_n1197_), .A1(ori_ori_n554_), .B0(ori_ori_n1181_), .Y(ori_ori_n1199_));
  AOI210     o1171(.A0(ori_ori_n1199_), .A1(ori_ori_n1198_), .B0(ori_ori_n327_), .Y(ori_ori_n1200_));
  OAI210     o1172(.A0(ori_ori_n85_), .A1(ori_ori_n40_), .B0(ori_ori_n670_), .Y(ori_ori_n1201_));
  NA2        o1173(.A(ori_ori_n1201_), .B(ori_ori_n638_), .Y(ori_ori_n1202_));
  NO2        o1174(.A(ori_ori_n513_), .B(ori_ori_n166_), .Y(ori_ori_n1203_));
  NO2        o1175(.A(ori_ori_n603_), .B(ori_ori_n1040_), .Y(ori_ori_n1204_));
  OAI210     o1176(.A0(ori_ori_n456_), .A1(ori_ori_n244_), .B0(ori_ori_n896_), .Y(ori_ori_n1205_));
  NO3        o1177(.A(ori_ori_n1205_), .B(ori_ori_n1204_), .C(ori_ori_n1203_), .Y(ori_ori_n1206_));
  NO2        o1178(.A(ori_ori_n361_), .B(ori_ori_n133_), .Y(ori_ori_n1207_));
  NA2        o1179(.A(ori_ori_n1207_), .B(ori_ori_n586_), .Y(ori_ori_n1208_));
  NA3        o1180(.A(ori_ori_n1208_), .B(ori_ori_n1206_), .C(ori_ori_n1202_), .Y(ori_ori_n1209_));
  NO2        o1181(.A(ori_ori_n742_), .B(ori_ori_n360_), .Y(ori_ori_n1210_));
  INV        o1182(.A(ori_ori_n672_), .Y(ori_ori_n1211_));
  NOi21      o1183(.An(ori_ori_n1210_), .B(ori_ori_n1211_), .Y(ori_ori_n1212_));
  AN2        o1184(.A(ori_ori_n945_), .B(ori_ori_n641_), .Y(ori_ori_n1213_));
  NO4        o1185(.A(ori_ori_n1213_), .B(ori_ori_n1212_), .C(ori_ori_n1209_), .D(ori_ori_n1200_), .Y(ori_ori_n1214_));
  NO2        o1186(.A(ori_ori_n729_), .B(ori_ori_n47_), .Y(ori_ori_n1215_));
  NA2        o1187(.A(ori_ori_n353_), .B(ori_ori_n1215_), .Y(ori_ori_n1216_));
  NO3        o1188(.A(ori_ori_n239_), .B(ori_ori_n100_), .C(ori_ori_n274_), .Y(ori_ori_n1217_));
  OAI220     o1189(.A0(ori_ori_n697_), .A1(ori_ori_n244_), .B0(ori_ori_n509_), .B1(ori_ori_n513_), .Y(ori_ori_n1218_));
  OAI210     o1190(.A0(l), .A1(i), .B0(k), .Y(ori_ori_n1219_));
  NO3        o1191(.A(ori_ori_n1219_), .B(ori_ori_n594_), .C(j), .Y(ori_ori_n1220_));
  NO3        o1192(.A(ori_ori_n1218_), .B(ori_ori_n1217_), .C(ori_ori_n1043_), .Y(ori_ori_n1221_));
  NA3        o1193(.A(ori_ori_n788_), .B(ori_ori_n787_), .C(ori_ori_n430_), .Y(ori_ori_n1222_));
  NAi31      o1194(.An(ori_ori_n742_), .B(ori_ori_n1222_), .C(ori_ori_n198_), .Y(ori_ori_n1223_));
  NA4        o1195(.A(ori_ori_n1223_), .B(ori_ori_n1221_), .C(ori_ori_n1216_), .D(ori_ori_n1115_), .Y(ori_ori_n1224_));
  NOi21      o1196(.An(ori_ori_n1193_), .B(ori_ori_n460_), .Y(ori_ori_n1225_));
  OR3        o1197(.A(ori_ori_n1225_), .B(ori_ori_n777_), .C(ori_ori_n537_), .Y(ori_ori_n1226_));
  NA2        o1198(.A(ori_ori_n568_), .B(ori_ori_n442_), .Y(ori_ori_n1227_));
  NA2        o1199(.A(ori_ori_n1220_), .B(ori_ori_n784_), .Y(ori_ori_n1228_));
  NA3        o1200(.A(ori_ori_n1228_), .B(ori_ori_n1227_), .C(ori_ori_n1226_), .Y(ori_ori_n1229_));
  AOI220     o1201(.A0(ori_ori_n1210_), .A1(ori_ori_n750_), .B0(ori_ori_n1207_), .B1(ori_ori_n234_), .Y(ori_ori_n1230_));
  AN2        o1202(.A(ori_ori_n917_), .B(ori_ori_n916_), .Y(ori_ori_n1231_));
  NO4        o1203(.A(ori_ori_n1231_), .B(ori_ori_n864_), .C(ori_ori_n499_), .D(ori_ori_n480_), .Y(ori_ori_n1232_));
  NA3        o1204(.A(ori_ori_n1232_), .B(ori_ori_n1230_), .C(ori_ori_n1176_), .Y(ori_ori_n1233_));
  NAi21      o1205(.An(j), .B(i), .Y(ori_ori_n1234_));
  NO4        o1206(.A(ori_ori_n1187_), .B(ori_ori_n1234_), .C(ori_ori_n436_), .D(ori_ori_n231_), .Y(ori_ori_n1235_));
  NO4        o1207(.A(ori_ori_n1235_), .B(ori_ori_n1233_), .C(ori_ori_n1229_), .D(ori_ori_n1224_), .Y(ori_ori_n1236_));
  NA4        o1208(.A(ori_ori_n1236_), .B(ori_ori_n1214_), .C(ori_ori_n1196_), .D(ori_ori_n1189_), .Y(ori07));
  NAi32      o1209(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1238_));
  NO3        o1210(.A(ori_ori_n1238_), .B(g), .C(f), .Y(ori_ori_n1239_));
  NAi21      o1211(.An(f), .B(c), .Y(ori_ori_n1240_));
  OR2        o1212(.A(e), .B(d), .Y(ori_ori_n1241_));
  NOi31      o1213(.An(n), .B(m), .C(b), .Y(ori_ori_n1242_));
  NOi41      o1214(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1243_));
  NO2        o1215(.A(ori_ori_n1025_), .B(ori_ori_n296_), .Y(ori_ori_n1244_));
  NA2        o1216(.A(ori_ori_n538_), .B(ori_ori_n76_), .Y(ori_ori_n1245_));
  NA2        o1217(.A(ori_ori_n1116_), .B(ori_ori_n281_), .Y(ori_ori_n1246_));
  NA2        o1218(.A(ori_ori_n1246_), .B(ori_ori_n1245_), .Y(ori_ori_n1247_));
  NO2        o1219(.A(ori_ori_n1247_), .B(ori_ori_n1239_), .Y(ori_ori_n1248_));
  NO3        o1220(.A(e), .B(d), .C(c), .Y(ori_ori_n1249_));
  NO2        o1221(.A(ori_ori_n129_), .B(ori_ori_n210_), .Y(ori_ori_n1250_));
  NA2        o1222(.A(ori_ori_n1250_), .B(ori_ori_n1249_), .Y(ori_ori_n1251_));
  INV        o1223(.A(ori_ori_n1251_), .Y(ori_ori_n1252_));
  NA3        o1224(.A(ori_ori_n694_), .B(ori_ori_n680_), .C(ori_ori_n110_), .Y(ori_ori_n1253_));
  NO2        o1225(.A(ori_ori_n1253_), .B(ori_ori_n45_), .Y(ori_ori_n1254_));
  NO2        o1226(.A(l), .B(k), .Y(ori_ori_n1255_));
  NO3        o1227(.A(ori_ori_n436_), .B(d), .C(c), .Y(ori_ori_n1256_));
  NO2        o1228(.A(ori_ori_n1254_), .B(ori_ori_n1252_), .Y(ori_ori_n1257_));
  NO2        o1229(.A(g), .B(c), .Y(ori_ori_n1258_));
  NO2        o1230(.A(ori_ori_n447_), .B(a), .Y(ori_ori_n1259_));
  NA2        o1231(.A(ori_ori_n1259_), .B(ori_ori_n111_), .Y(ori_ori_n1260_));
  NA2        o1232(.A(ori_ori_n135_), .B(ori_ori_n217_), .Y(ori_ori_n1261_));
  NO2        o1233(.A(ori_ori_n1261_), .B(ori_ori_n1354_), .Y(ori_ori_n1262_));
  NO2        o1234(.A(ori_ori_n748_), .B(ori_ori_n182_), .Y(ori_ori_n1263_));
  NOi31      o1235(.An(m), .B(n), .C(b), .Y(ori_ori_n1264_));
  NOi31      o1236(.An(f), .B(d), .C(c), .Y(ori_ori_n1265_));
  NA2        o1237(.A(ori_ori_n1265_), .B(ori_ori_n1264_), .Y(ori_ori_n1266_));
  INV        o1238(.A(ori_ori_n1266_), .Y(ori_ori_n1267_));
  NO3        o1239(.A(ori_ori_n1267_), .B(ori_ori_n1263_), .C(ori_ori_n1262_), .Y(ori_ori_n1268_));
  NA2        o1240(.A(ori_ori_n1026_), .B(ori_ori_n463_), .Y(ori_ori_n1269_));
  NO2        o1241(.A(ori_ori_n1269_), .B(ori_ori_n436_), .Y(ori_ori_n1270_));
  NO3        o1242(.A(ori_ori_n41_), .B(i), .C(h), .Y(ori_ori_n1271_));
  NO2        o1243(.A(ori_ori_n1024_), .B(ori_ori_n1270_), .Y(ori_ori_n1272_));
  AN3        o1244(.A(ori_ori_n1272_), .B(ori_ori_n1268_), .C(ori_ori_n1260_), .Y(ori_ori_n1273_));
  NA2        o1245(.A(ori_ori_n1242_), .B(ori_ori_n371_), .Y(ori_ori_n1274_));
  INV        o1246(.A(ori_ori_n1274_), .Y(ori_ori_n1275_));
  INV        o1247(.A(ori_ori_n1029_), .Y(ori_ori_n1276_));
  NAi21      o1248(.An(ori_ori_n1275_), .B(ori_ori_n1276_), .Y(ori_ori_n1277_));
  NO4        o1249(.A(ori_ori_n129_), .B(g), .C(f), .D(e), .Y(ori_ori_n1278_));
  NA2        o1250(.A(ori_ori_n1243_), .B(ori_ori_n1255_), .Y(ori_ori_n1279_));
  INV        o1251(.A(ori_ori_n1279_), .Y(ori_ori_n1280_));
  OR3        o1252(.A(ori_ori_n537_), .B(ori_ori_n536_), .C(ori_ori_n110_), .Y(ori_ori_n1281_));
  NA2        o1253(.A(ori_ori_n1039_), .B(ori_ori_n400_), .Y(ori_ori_n1282_));
  NO2        o1254(.A(ori_ori_n1282_), .B(ori_ori_n429_), .Y(ori_ori_n1283_));
  AO210      o1255(.A0(ori_ori_n1283_), .A1(ori_ori_n114_), .B0(ori_ori_n1280_), .Y(ori_ori_n1284_));
  NO2        o1256(.A(ori_ori_n1284_), .B(ori_ori_n1277_), .Y(ori_ori_n1285_));
  NA4        o1257(.A(ori_ori_n1285_), .B(ori_ori_n1273_), .C(ori_ori_n1257_), .D(ori_ori_n1248_), .Y(ori_ori_n1286_));
  NO2        o1258(.A(ori_ori_n1048_), .B(ori_ori_n108_), .Y(ori_ori_n1287_));
  NO2        o1259(.A(ori_ori_n383_), .B(j), .Y(ori_ori_n1288_));
  NA2        o1260(.A(ori_ori_n1271_), .B(ori_ori_n1039_), .Y(ori_ori_n1289_));
  INV        o1261(.A(ori_ori_n1289_), .Y(ori_ori_n1290_));
  NA2        o1262(.A(ori_ori_n1288_), .B(ori_ori_n157_), .Y(ori_ori_n1291_));
  INV        o1263(.A(ori_ori_n1291_), .Y(ori_ori_n1292_));
  NO2        o1264(.A(ori_ori_n1292_), .B(ori_ori_n1290_), .Y(ori_ori_n1293_));
  INV        o1265(.A(ori_ori_n49_), .Y(ori_ori_n1294_));
  NA2        o1266(.A(ori_ori_n1294_), .B(ori_ori_n1082_), .Y(ori_ori_n1295_));
  INV        o1267(.A(ori_ori_n1295_), .Y(ori_ori_n1296_));
  NO2        o1268(.A(ori_ori_n662_), .B(ori_ori_n171_), .Y(ori_ori_n1297_));
  NO2        o1269(.A(ori_ori_n1297_), .B(ori_ori_n1296_), .Y(ori_ori_n1298_));
  NO3        o1270(.A(ori_ori_n1031_), .B(ori_ori_n1241_), .C(ori_ori_n49_), .Y(ori_ori_n1299_));
  NA3        o1271(.A(ori_ori_n1287_), .B(ori_ori_n463_), .C(f), .Y(ori_ori_n1300_));
  INV        o1272(.A(ori_ori_n174_), .Y(ori_ori_n1301_));
  NO2        o1273(.A(ori_ori_n1352_), .B(ori_ori_n1300_), .Y(ori_ori_n1302_));
  NO2        o1274(.A(ori_ori_n1234_), .B(ori_ori_n169_), .Y(ori_ori_n1303_));
  NOi21      o1275(.An(d), .B(f), .Y(ori_ori_n1304_));
  INV        o1276(.A(ori_ori_n1302_), .Y(ori_ori_n1305_));
  NA3        o1277(.A(ori_ori_n1305_), .B(ori_ori_n1298_), .C(ori_ori_n1293_), .Y(ori_ori_n1306_));
  NA2        o1278(.A(h), .B(ori_ori_n1244_), .Y(ori_ori_n1307_));
  OAI210     o1279(.A0(ori_ori_n1278_), .A1(ori_ori_n1242_), .B0(ori_ori_n869_), .Y(ori_ori_n1308_));
  NO2        o1280(.A(ori_ori_n1021_), .B(ori_ori_n129_), .Y(ori_ori_n1309_));
  NA2        o1281(.A(ori_ori_n1309_), .B(ori_ori_n616_), .Y(ori_ori_n1310_));
  NA3        o1282(.A(ori_ori_n1310_), .B(ori_ori_n1308_), .C(ori_ori_n1307_), .Y(ori_ori_n1311_));
  NA2        o1283(.A(ori_ori_n1258_), .B(ori_ori_n1304_), .Y(ori_ori_n1312_));
  NO2        o1284(.A(ori_ori_n1312_), .B(m), .Y(ori_ori_n1313_));
  NO2        o1285(.A(ori_ori_n149_), .B(ori_ori_n176_), .Y(ori_ori_n1314_));
  OAI210     o1286(.A0(ori_ori_n1314_), .A1(ori_ori_n108_), .B0(ori_ori_n1264_), .Y(ori_ori_n1315_));
  INV        o1287(.A(ori_ori_n1315_), .Y(ori_ori_n1316_));
  NO3        o1288(.A(ori_ori_n1316_), .B(ori_ori_n1313_), .C(ori_ori_n1311_), .Y(ori_ori_n1317_));
  NO2        o1289(.A(ori_ori_n1240_), .B(e), .Y(ori_ori_n1318_));
  NA2        o1290(.A(ori_ori_n1318_), .B(ori_ori_n398_), .Y(ori_ori_n1319_));
  BUFFER     o1291(.A(ori_ori_n129_), .Y(ori_ori_n1320_));
  NO2        o1292(.A(ori_ori_n1320_), .B(ori_ori_n1319_), .Y(ori_ori_n1321_));
  NO2        o1293(.A(ori_ori_n1281_), .B(ori_ori_n344_), .Y(ori_ori_n1322_));
  NO2        o1294(.A(ori_ori_n1322_), .B(ori_ori_n1321_), .Y(ori_ori_n1323_));
  NO2        o1295(.A(ori_ori_n176_), .B(c), .Y(ori_ori_n1324_));
  NA2        o1296(.A(ori_ori_n1324_), .B(ori_ori_n174_), .Y(ori_ori_n1325_));
  INV        o1297(.A(ori_ori_n1325_), .Y(ori_ori_n1326_));
  NO2        o1298(.A(ori_ori_n1256_), .B(ori_ori_n1299_), .Y(ori_ori_n1327_));
  INV        o1299(.A(ori_ori_n1046_), .Y(ori_ori_n1328_));
  OAI210     o1300(.A0(ori_ori_n1328_), .A1(ori_ori_n65_), .B0(ori_ori_n1327_), .Y(ori_ori_n1329_));
  OR2        o1301(.A(h), .B(ori_ori_n536_), .Y(ori_ori_n1330_));
  NO2        o1302(.A(ori_ori_n1330_), .B(ori_ori_n169_), .Y(ori_ori_n1331_));
  NA2        o1303(.A(ori_ori_n1030_), .B(ori_ori_n217_), .Y(ori_ori_n1332_));
  NO2        o1304(.A(ori_ori_n49_), .B(l), .Y(ori_ori_n1333_));
  INV        o1305(.A(ori_ori_n482_), .Y(ori_ori_n1334_));
  NA2        o1306(.A(ori_ori_n1334_), .B(ori_ori_n1333_), .Y(ori_ori_n1335_));
  NA2        o1307(.A(ori_ori_n1335_), .B(ori_ori_n1332_), .Y(ori_ori_n1336_));
  NO4        o1308(.A(ori_ori_n1336_), .B(ori_ori_n1331_), .C(ori_ori_n1329_), .D(ori_ori_n1326_), .Y(ori_ori_n1337_));
  NA3        o1309(.A(ori_ori_n1337_), .B(ori_ori_n1323_), .C(ori_ori_n1317_), .Y(ori_ori_n1338_));
  NA3        o1310(.A(ori_ori_n949_), .B(ori_ori_n135_), .C(ori_ori_n46_), .Y(ori_ori_n1339_));
  INV        o1311(.A(ori_ori_n1339_), .Y(ori_ori_n1340_));
  NA2        o1312(.A(ori_ori_n1303_), .B(h), .Y(ori_ori_n1341_));
  INV        o1313(.A(ori_ori_n1341_), .Y(ori_ori_n1342_));
  NO2        o1314(.A(ori_ori_n1342_), .B(ori_ori_n1340_), .Y(ori_ori_n1343_));
  INV        o1315(.A(ori_ori_n1318_), .Y(ori_ori_n1344_));
  NO2        o1316(.A(ori_ori_n1344_), .B(ori_ori_n1301_), .Y(ori_ori_n1345_));
  INV        o1317(.A(ori_ori_n1345_), .Y(ori_ori_n1346_));
  NO2        o1318(.A(ori_ori_n1282_), .B(d), .Y(ori_ori_n1347_));
  NA3        o1319(.A(ori_ori_n1353_), .B(ori_ori_n1346_), .C(ori_ori_n1343_), .Y(ori_ori_n1348_));
  OR4        o1320(.A(ori_ori_n1348_), .B(ori_ori_n1338_), .C(ori_ori_n1306_), .D(ori_ori_n1286_), .Y(ori04));
  INV        o1321(.A(ori_ori_n111_), .Y(ori_ori_n1352_));
  INV        o1322(.A(ori_ori_n1347_), .Y(ori_ori_n1353_));
  INV        o1323(.A(h), .Y(ori_ori_n1354_));
  ZERO       o1324(.Y(ori02));
  ZERO       o1325(.Y(ori03));
  ZERO       o1326(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO2        m0025(.A(mai_mai_n53_), .B(mai_mai_n39_), .Y(mai_mai_n54_));
  NO2        m0026(.A(mai_mai_n54_), .B(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NA3        m0031(.A(g), .B(mai_mai_n59_), .C(a), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(h), .Y(mai_mai_n61_));
  NAi31      m0033(.An(i), .B(l), .C(j), .Y(mai_mai_n62_));
  OAI220     m0034(.A0(mai_mai_n62_), .A1(mai_mai_n49_), .B0(mai_mai_n61_), .B1(mai_mai_n44_), .Y(mai_mai_n63_));
  NAi31      m0035(.An(mai_mai_n60_), .B(mai_mai_n63_), .C(mai_mai_n58_), .Y(mai_mai_n64_));
  NAi41      m0036(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(g), .B(f), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi21      m0039(.An(i), .B(j), .Y(mai_mai_n68_));
  NAi32      m0040(.An(n), .Bn(k), .C(m), .Y(mai_mai_n69_));
  NO2        m0041(.A(mai_mai_n69_), .B(mai_mai_n68_), .Y(mai_mai_n70_));
  NAi31      m0042(.An(l), .B(m), .C(k), .Y(mai_mai_n71_));
  NAi21      m0043(.An(e), .B(h), .Y(mai_mai_n72_));
  NAi41      m0044(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n74_));
  INV        m0046(.A(m), .Y(mai_mai_n75_));
  NOi21      m0047(.An(k), .B(l), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  AN4        m0049(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n78_));
  NOi31      m0050(.An(h), .B(g), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  NAi32      m0052(.An(m), .Bn(k), .C(j), .Y(mai_mai_n81_));
  NOi32      m0053(.An(h), .Bn(g), .C(f), .Y(mai_mai_n82_));
  NA2        m0054(.A(mai_mai_n82_), .B(mai_mai_n78_), .Y(mai_mai_n83_));
  OA220      m0055(.A0(mai_mai_n83_), .A1(mai_mai_n81_), .B0(mai_mai_n80_), .B1(mai_mai_n77_), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(mai_mai_n74_), .C(mai_mai_n64_), .Y(mai_mai_n85_));
  INV        m0057(.A(n), .Y(mai_mai_n86_));
  NOi32      m0058(.An(e), .Bn(b), .C(d), .Y(mai_mai_n87_));
  NA2        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .Y(mai_mai_n88_));
  INV        m0060(.A(j), .Y(mai_mai_n89_));
  AN3        m0061(.A(m), .B(k), .C(i), .Y(mai_mai_n90_));
  NA3        m0062(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(g), .Y(mai_mai_n91_));
  NAi32      m0063(.An(g), .Bn(f), .C(h), .Y(mai_mai_n92_));
  NAi31      m0064(.An(j), .B(m), .C(l), .Y(mai_mai_n93_));
  NA2        m0065(.A(m), .B(l), .Y(mai_mai_n94_));
  NAi31      m0066(.An(k), .B(j), .C(g), .Y(mai_mai_n95_));
  NO3        m0067(.A(mai_mai_n95_), .B(mai_mai_n94_), .C(f), .Y(mai_mai_n96_));
  AN2        m0068(.A(j), .B(g), .Y(mai_mai_n97_));
  NOi32      m0069(.An(m), .Bn(l), .C(i), .Y(mai_mai_n98_));
  NOi21      m0070(.An(g), .B(i), .Y(mai_mai_n99_));
  NOi32      m0071(.An(m), .Bn(j), .C(k), .Y(mai_mai_n100_));
  AOI220     m0072(.A0(mai_mai_n100_), .A1(mai_mai_n99_), .B0(mai_mai_n98_), .B1(mai_mai_n97_), .Y(mai_mai_n101_));
  NAi41      m0073(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n102_));
  AN2        m0074(.A(e), .B(b), .Y(mai_mai_n103_));
  NOi31      m0075(.An(c), .B(h), .C(f), .Y(mai_mai_n104_));
  NA2        m0076(.A(mai_mai_n104_), .B(mai_mai_n103_), .Y(mai_mai_n105_));
  NO2        m0077(.A(mai_mai_n105_), .B(mai_mai_n102_), .Y(mai_mai_n106_));
  NOi21      m0078(.An(g), .B(f), .Y(mai_mai_n107_));
  NOi21      m0079(.An(i), .B(h), .Y(mai_mai_n108_));
  INV        m0080(.A(a), .Y(mai_mai_n109_));
  NA2        m0081(.A(mai_mai_n103_), .B(mai_mai_n109_), .Y(mai_mai_n110_));
  INV        m0082(.A(l), .Y(mai_mai_n111_));
  NOi21      m0083(.An(m), .B(n), .Y(mai_mai_n112_));
  AN2        m0084(.A(k), .B(h), .Y(mai_mai_n113_));
  INV        m0085(.A(b), .Y(mai_mai_n114_));
  NA2        m0086(.A(l), .B(j), .Y(mai_mai_n115_));
  AN2        m0087(.A(k), .B(i), .Y(mai_mai_n116_));
  NA2        m0088(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NA2        m0089(.A(g), .B(e), .Y(mai_mai_n118_));
  NOi32      m0090(.An(c), .Bn(a), .C(d), .Y(mai_mai_n119_));
  NA2        m0091(.A(mai_mai_n119_), .B(mai_mai_n112_), .Y(mai_mai_n120_));
  NO4        m0092(.A(mai_mai_n120_), .B(mai_mai_n118_), .C(mai_mai_n117_), .D(mai_mai_n114_), .Y(mai_mai_n121_));
  NO2        m0093(.A(mai_mai_n121_), .B(mai_mai_n106_), .Y(mai_mai_n122_));
  OAI210     m0094(.A0(mai_mai_n91_), .A1(mai_mai_n88_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  NOi31      m0095(.An(k), .B(m), .C(j), .Y(mai_mai_n124_));
  NOi31      m0096(.An(k), .B(m), .C(i), .Y(mai_mai_n125_));
  NA3        m0097(.A(mai_mai_n125_), .B(mai_mai_n82_), .C(mai_mai_n78_), .Y(mai_mai_n126_));
  INV        m0098(.A(mai_mai_n126_), .Y(mai_mai_n127_));
  NOi32      m0099(.An(f), .Bn(b), .C(e), .Y(mai_mai_n128_));
  NAi21      m0100(.An(g), .B(h), .Y(mai_mai_n129_));
  NAi21      m0101(.An(m), .B(n), .Y(mai_mai_n130_));
  NAi21      m0102(.An(j), .B(k), .Y(mai_mai_n131_));
  NO3        m0103(.A(mai_mai_n131_), .B(mai_mai_n130_), .C(mai_mai_n129_), .Y(mai_mai_n132_));
  NAi41      m0104(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n133_));
  NAi31      m0105(.An(j), .B(k), .C(h), .Y(mai_mai_n134_));
  NO3        m0106(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n130_), .Y(mai_mai_n135_));
  AOI210     m0107(.A0(mai_mai_n132_), .A1(mai_mai_n128_), .B0(mai_mai_n135_), .Y(mai_mai_n136_));
  NO2        m0108(.A(k), .B(j), .Y(mai_mai_n137_));
  NO2        m0109(.A(mai_mai_n137_), .B(mai_mai_n130_), .Y(mai_mai_n138_));
  AN2        m0110(.A(k), .B(j), .Y(mai_mai_n139_));
  NAi21      m0111(.An(c), .B(b), .Y(mai_mai_n140_));
  NA2        m0112(.A(f), .B(d), .Y(mai_mai_n141_));
  NO4        m0113(.A(mai_mai_n141_), .B(mai_mai_n140_), .C(mai_mai_n139_), .D(mai_mai_n129_), .Y(mai_mai_n142_));
  NA2        m0114(.A(h), .B(c), .Y(mai_mai_n143_));
  NAi31      m0115(.An(f), .B(e), .C(b), .Y(mai_mai_n144_));
  NA2        m0116(.A(mai_mai_n142_), .B(mai_mai_n138_), .Y(mai_mai_n145_));
  NA2        m0117(.A(d), .B(b), .Y(mai_mai_n146_));
  NAi21      m0118(.An(e), .B(f), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n147_), .B(mai_mai_n146_), .Y(mai_mai_n148_));
  NA2        m0120(.A(b), .B(a), .Y(mai_mai_n149_));
  NAi21      m0121(.An(e), .B(g), .Y(mai_mai_n150_));
  NAi21      m0122(.An(c), .B(d), .Y(mai_mai_n151_));
  NAi31      m0123(.An(l), .B(k), .C(h), .Y(mai_mai_n152_));
  NO2        m0124(.A(mai_mai_n130_), .B(mai_mai_n152_), .Y(mai_mai_n153_));
  NAi31      m0125(.An(mai_mai_n127_), .B(mai_mai_n145_), .C(mai_mai_n136_), .Y(mai_mai_n154_));
  NAi31      m0126(.An(e), .B(f), .C(b), .Y(mai_mai_n155_));
  NOi21      m0127(.An(g), .B(d), .Y(mai_mai_n156_));
  NO2        m0128(.A(mai_mai_n156_), .B(mai_mai_n155_), .Y(mai_mai_n157_));
  NOi21      m0129(.An(h), .B(i), .Y(mai_mai_n158_));
  NOi21      m0130(.An(k), .B(m), .Y(mai_mai_n159_));
  NA3        m0131(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(n), .Y(mai_mai_n160_));
  NOi21      m0132(.An(mai_mai_n157_), .B(mai_mai_n160_), .Y(mai_mai_n161_));
  NOi21      m0133(.An(h), .B(g), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n141_), .B(mai_mai_n140_), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  NAi31      m0136(.An(l), .B(j), .C(h), .Y(mai_mai_n165_));
  NO2        m0137(.A(mai_mai_n165_), .B(mai_mai_n49_), .Y(mai_mai_n166_));
  NA2        m0138(.A(mai_mai_n166_), .B(mai_mai_n67_), .Y(mai_mai_n167_));
  NOi32      m0139(.An(n), .Bn(k), .C(m), .Y(mai_mai_n168_));
  NA2        m0140(.A(l), .B(i), .Y(mai_mai_n169_));
  NA2        m0141(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  OAI210     m0142(.A0(mai_mai_n170_), .A1(mai_mai_n164_), .B0(mai_mai_n167_), .Y(mai_mai_n171_));
  NAi31      m0143(.An(d), .B(f), .C(c), .Y(mai_mai_n172_));
  NAi31      m0144(.An(e), .B(f), .C(c), .Y(mai_mai_n173_));
  NA2        m0145(.A(mai_mai_n173_), .B(mai_mai_n172_), .Y(mai_mai_n174_));
  NA2        m0146(.A(j), .B(h), .Y(mai_mai_n175_));
  OR3        m0147(.A(n), .B(m), .C(k), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n176_), .B(mai_mai_n175_), .Y(mai_mai_n177_));
  NAi32      m0149(.An(m), .Bn(k), .C(n), .Y(mai_mai_n178_));
  NO2        m0150(.A(mai_mai_n178_), .B(mai_mai_n175_), .Y(mai_mai_n179_));
  AOI220     m0151(.A0(mai_mai_n179_), .A1(mai_mai_n157_), .B0(mai_mai_n177_), .B1(mai_mai_n174_), .Y(mai_mai_n180_));
  NO2        m0152(.A(n), .B(m), .Y(mai_mai_n181_));
  NA2        m0153(.A(mai_mai_n181_), .B(mai_mai_n50_), .Y(mai_mai_n182_));
  NAi21      m0154(.An(f), .B(e), .Y(mai_mai_n183_));
  NA2        m0155(.A(d), .B(c), .Y(mai_mai_n184_));
  NO2        m0156(.A(mai_mai_n184_), .B(mai_mai_n183_), .Y(mai_mai_n185_));
  NOi21      m0157(.An(mai_mai_n185_), .B(mai_mai_n182_), .Y(mai_mai_n186_));
  NAi21      m0158(.An(d), .B(c), .Y(mai_mai_n187_));
  NAi31      m0159(.An(m), .B(n), .C(b), .Y(mai_mai_n188_));
  NA2        m0160(.A(k), .B(i), .Y(mai_mai_n189_));
  NAi21      m0161(.An(h), .B(f), .Y(mai_mai_n190_));
  NO2        m0162(.A(mai_mai_n190_), .B(mai_mai_n189_), .Y(mai_mai_n191_));
  NO2        m0163(.A(mai_mai_n188_), .B(mai_mai_n151_), .Y(mai_mai_n192_));
  NA2        m0164(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  NOi32      m0165(.An(f), .Bn(c), .C(d), .Y(mai_mai_n194_));
  NOi32      m0166(.An(f), .Bn(c), .C(e), .Y(mai_mai_n195_));
  NO2        m0167(.A(mai_mai_n195_), .B(mai_mai_n194_), .Y(mai_mai_n196_));
  NO3        m0168(.A(n), .B(m), .C(j), .Y(mai_mai_n197_));
  NA2        m0169(.A(mai_mai_n197_), .B(mai_mai_n113_), .Y(mai_mai_n198_));
  AO210      m0170(.A0(mai_mai_n198_), .A1(mai_mai_n182_), .B0(mai_mai_n196_), .Y(mai_mai_n199_));
  NAi41      m0171(.An(mai_mai_n186_), .B(mai_mai_n199_), .C(mai_mai_n193_), .D(mai_mai_n180_), .Y(mai_mai_n200_));
  OR4        m0172(.A(mai_mai_n200_), .B(mai_mai_n171_), .C(mai_mai_n161_), .D(mai_mai_n154_), .Y(mai_mai_n201_));
  NO4        m0173(.A(mai_mai_n201_), .B(mai_mai_n123_), .C(mai_mai_n85_), .D(mai_mai_n55_), .Y(mai_mai_n202_));
  NA3        m0174(.A(m), .B(mai_mai_n111_), .C(j), .Y(mai_mai_n203_));
  NAi31      m0175(.An(n), .B(h), .C(g), .Y(mai_mai_n204_));
  NO2        m0176(.A(mai_mai_n204_), .B(mai_mai_n203_), .Y(mai_mai_n205_));
  NOi32      m0177(.An(m), .Bn(k), .C(l), .Y(mai_mai_n206_));
  NA3        m0178(.A(mai_mai_n206_), .B(mai_mai_n89_), .C(g), .Y(mai_mai_n207_));
  NO2        m0179(.A(mai_mai_n207_), .B(n), .Y(mai_mai_n208_));
  AN2        m0180(.A(i), .B(g), .Y(mai_mai_n209_));
  NA3        m0181(.A(mai_mai_n76_), .B(mai_mai_n209_), .C(mai_mai_n112_), .Y(mai_mai_n210_));
  NAi41      m0182(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n211_));
  INV        m0183(.A(mai_mai_n211_), .Y(mai_mai_n212_));
  INV        m0184(.A(f), .Y(mai_mai_n213_));
  INV        m0185(.A(g), .Y(mai_mai_n214_));
  NOi31      m0186(.An(i), .B(j), .C(h), .Y(mai_mai_n215_));
  NOi21      m0187(.An(l), .B(m), .Y(mai_mai_n216_));
  NA2        m0188(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n217_));
  NO3        m0189(.A(mai_mai_n217_), .B(mai_mai_n214_), .C(mai_mai_n213_), .Y(mai_mai_n218_));
  NA2        m0190(.A(mai_mai_n218_), .B(mai_mai_n212_), .Y(mai_mai_n219_));
  INV        m0191(.A(mai_mai_n219_), .Y(mai_mai_n220_));
  NOi21      m0192(.An(n), .B(m), .Y(mai_mai_n221_));
  NOi32      m0193(.An(l), .Bn(i), .C(j), .Y(mai_mai_n222_));
  NA2        m0194(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n223_));
  OA220      m0195(.A0(mai_mai_n223_), .A1(mai_mai_n105_), .B0(mai_mai_n81_), .B1(mai_mai_n80_), .Y(mai_mai_n224_));
  NAi21      m0196(.An(j), .B(h), .Y(mai_mai_n225_));
  XN2        m0197(.A(i), .B(h), .Y(mai_mai_n226_));
  NA2        m0198(.A(mai_mai_n226_), .B(mai_mai_n225_), .Y(mai_mai_n227_));
  NOi31      m0199(.An(k), .B(n), .C(m), .Y(mai_mai_n228_));
  NOi31      m0200(.An(mai_mai_n228_), .B(mai_mai_n184_), .C(mai_mai_n183_), .Y(mai_mai_n229_));
  NA2        m0201(.A(mai_mai_n229_), .B(mai_mai_n227_), .Y(mai_mai_n230_));
  NAi31      m0202(.An(f), .B(e), .C(c), .Y(mai_mai_n231_));
  NO4        m0203(.A(mai_mai_n231_), .B(mai_mai_n176_), .C(mai_mai_n175_), .D(mai_mai_n59_), .Y(mai_mai_n232_));
  NA4        m0204(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n233_));
  NAi32      m0205(.An(m), .Bn(i), .C(k), .Y(mai_mai_n234_));
  NO3        m0206(.A(mai_mai_n234_), .B(mai_mai_n92_), .C(mai_mai_n233_), .Y(mai_mai_n235_));
  INV        m0207(.A(k), .Y(mai_mai_n236_));
  NO2        m0208(.A(mai_mai_n235_), .B(mai_mai_n232_), .Y(mai_mai_n237_));
  NAi21      m0209(.An(n), .B(a), .Y(mai_mai_n238_));
  NO2        m0210(.A(mai_mai_n238_), .B(mai_mai_n146_), .Y(mai_mai_n239_));
  NAi41      m0211(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n240_));
  NO2        m0212(.A(mai_mai_n240_), .B(e), .Y(mai_mai_n241_));
  NO3        m0213(.A(mai_mai_n147_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n242_));
  OAI210     m0214(.A0(mai_mai_n242_), .A1(mai_mai_n241_), .B0(mai_mai_n239_), .Y(mai_mai_n243_));
  AN4        m0215(.A(mai_mai_n243_), .B(mai_mai_n237_), .C(mai_mai_n230_), .D(mai_mai_n224_), .Y(mai_mai_n244_));
  OR2        m0216(.A(h), .B(g), .Y(mai_mai_n245_));
  NO2        m0217(.A(mai_mai_n245_), .B(mai_mai_n102_), .Y(mai_mai_n246_));
  NA2        m0218(.A(mai_mai_n246_), .B(mai_mai_n128_), .Y(mai_mai_n247_));
  NAi31      m0219(.An(e), .B(d), .C(b), .Y(mai_mai_n248_));
  NA2        m0220(.A(mai_mai_n159_), .B(mai_mai_n108_), .Y(mai_mai_n249_));
  NO2        m0221(.A(n), .B(a), .Y(mai_mai_n250_));
  NAi31      m0222(.An(mai_mai_n240_), .B(mai_mai_n250_), .C(mai_mai_n103_), .Y(mai_mai_n251_));
  NAi21      m0223(.An(h), .B(i), .Y(mai_mai_n252_));
  NA2        m0224(.A(mai_mai_n181_), .B(k), .Y(mai_mai_n253_));
  NO2        m0225(.A(mai_mai_n253_), .B(mai_mai_n252_), .Y(mai_mai_n254_));
  NA2        m0226(.A(mai_mai_n254_), .B(mai_mai_n194_), .Y(mai_mai_n255_));
  NA3        m0227(.A(mai_mai_n255_), .B(mai_mai_n251_), .C(mai_mai_n247_), .Y(mai_mai_n256_));
  NOi21      m0228(.An(g), .B(e), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n258_), .B(mai_mai_n257_), .Y(mai_mai_n259_));
  NOi32      m0231(.An(l), .Bn(j), .C(i), .Y(mai_mai_n260_));
  AOI210     m0232(.A0(mai_mai_n76_), .A1(mai_mai_n89_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  NO2        m0233(.A(mai_mai_n252_), .B(mai_mai_n44_), .Y(mai_mai_n262_));
  NAi21      m0234(.An(f), .B(g), .Y(mai_mai_n263_));
  NO2        m0235(.A(mai_mai_n263_), .B(mai_mai_n65_), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n69_), .B(mai_mai_n115_), .Y(mai_mai_n265_));
  AOI220     m0237(.A0(mai_mai_n265_), .A1(mai_mai_n264_), .B0(mai_mai_n262_), .B1(mai_mai_n67_), .Y(mai_mai_n266_));
  OAI210     m0238(.A0(mai_mai_n261_), .A1(mai_mai_n259_), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  NO3        m0239(.A(mai_mai_n131_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n268_));
  NOi41      m0240(.An(mai_mai_n244_), .B(mai_mai_n267_), .C(mai_mai_n256_), .D(mai_mai_n220_), .Y(mai_mai_n269_));
  NO4        m0241(.A(mai_mai_n205_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n270_));
  NO2        m0242(.A(mai_mai_n270_), .B(mai_mai_n110_), .Y(mai_mai_n271_));
  NA3        m0243(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n272_));
  NAi21      m0244(.An(h), .B(g), .Y(mai_mai_n273_));
  OR4        m0245(.A(mai_mai_n273_), .B(mai_mai_n272_), .C(mai_mai_n223_), .D(e), .Y(mai_mai_n274_));
  NO2        m0246(.A(mai_mai_n249_), .B(mai_mai_n263_), .Y(mai_mai_n275_));
  NAi31      m0247(.An(g), .B(k), .C(h), .Y(mai_mai_n276_));
  NO3        m0248(.A(mai_mai_n130_), .B(mai_mai_n276_), .C(l), .Y(mai_mai_n277_));
  NAi31      m0249(.An(e), .B(d), .C(a), .Y(mai_mai_n278_));
  NA2        m0250(.A(mai_mai_n277_), .B(mai_mai_n128_), .Y(mai_mai_n279_));
  NA2        m0251(.A(mai_mai_n279_), .B(mai_mai_n274_), .Y(mai_mai_n280_));
  NA4        m0252(.A(mai_mai_n159_), .B(mai_mai_n82_), .C(mai_mai_n78_), .D(mai_mai_n115_), .Y(mai_mai_n281_));
  NA3        m0253(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(mai_mai_n86_), .Y(mai_mai_n282_));
  NO2        m0254(.A(mai_mai_n282_), .B(mai_mai_n196_), .Y(mai_mai_n283_));
  NOi21      m0255(.An(mai_mai_n281_), .B(mai_mai_n283_), .Y(mai_mai_n284_));
  NA3        m0256(.A(e), .B(c), .C(b), .Y(mai_mai_n285_));
  NO2        m0257(.A(mai_mai_n60_), .B(mai_mai_n285_), .Y(mai_mai_n286_));
  NAi32      m0258(.An(k), .Bn(i), .C(j), .Y(mai_mai_n287_));
  NAi31      m0259(.An(h), .B(l), .C(i), .Y(mai_mai_n288_));
  NA3        m0260(.A(mai_mai_n288_), .B(mai_mai_n287_), .C(mai_mai_n165_), .Y(mai_mai_n289_));
  NOi21      m0261(.An(mai_mai_n289_), .B(mai_mai_n49_), .Y(mai_mai_n290_));
  OAI210     m0262(.A0(mai_mai_n264_), .A1(mai_mai_n286_), .B0(mai_mai_n290_), .Y(mai_mai_n291_));
  NAi21      m0263(.An(l), .B(k), .Y(mai_mai_n292_));
  NO2        m0264(.A(mai_mai_n292_), .B(mai_mai_n49_), .Y(mai_mai_n293_));
  NOi21      m0265(.An(l), .B(j), .Y(mai_mai_n294_));
  NA2        m0266(.A(mai_mai_n162_), .B(mai_mai_n294_), .Y(mai_mai_n295_));
  NAi32      m0267(.An(j), .Bn(h), .C(i), .Y(mai_mai_n296_));
  NAi21      m0268(.An(m), .B(l), .Y(mai_mai_n297_));
  NO3        m0269(.A(mai_mai_n297_), .B(mai_mai_n296_), .C(mai_mai_n86_), .Y(mai_mai_n298_));
  NA2        m0270(.A(h), .B(g), .Y(mai_mai_n299_));
  NA2        m0271(.A(mai_mai_n168_), .B(mai_mai_n45_), .Y(mai_mai_n300_));
  NO2        m0272(.A(mai_mai_n300_), .B(mai_mai_n299_), .Y(mai_mai_n301_));
  OAI210     m0273(.A0(mai_mai_n301_), .A1(mai_mai_n298_), .B0(mai_mai_n163_), .Y(mai_mai_n302_));
  NA3        m0274(.A(mai_mai_n302_), .B(mai_mai_n291_), .C(mai_mai_n284_), .Y(mai_mai_n303_));
  NO2        m0275(.A(mai_mai_n144_), .B(d), .Y(mai_mai_n304_));
  NA2        m0276(.A(mai_mai_n304_), .B(mai_mai_n53_), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n105_), .B(mai_mai_n102_), .Y(mai_mai_n306_));
  NAi32      m0278(.An(n), .Bn(m), .C(l), .Y(mai_mai_n307_));
  NO2        m0279(.A(mai_mai_n307_), .B(mai_mai_n296_), .Y(mai_mai_n308_));
  NA2        m0280(.A(mai_mai_n308_), .B(mai_mai_n185_), .Y(mai_mai_n309_));
  NO2        m0281(.A(mai_mai_n120_), .B(mai_mai_n114_), .Y(mai_mai_n310_));
  NAi31      m0282(.An(k), .B(l), .C(j), .Y(mai_mai_n311_));
  OAI210     m0283(.A0(mai_mai_n292_), .A1(j), .B0(mai_mai_n311_), .Y(mai_mai_n312_));
  NOi21      m0284(.An(mai_mai_n312_), .B(mai_mai_n118_), .Y(mai_mai_n313_));
  NA2        m0285(.A(mai_mai_n313_), .B(mai_mai_n310_), .Y(mai_mai_n314_));
  NA3        m0286(.A(mai_mai_n314_), .B(mai_mai_n309_), .C(mai_mai_n305_), .Y(mai_mai_n315_));
  NO4        m0287(.A(mai_mai_n315_), .B(mai_mai_n303_), .C(mai_mai_n280_), .D(mai_mai_n271_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n254_), .B(mai_mai_n195_), .Y(mai_mai_n317_));
  NAi21      m0289(.An(m), .B(k), .Y(mai_mai_n318_));
  NO2        m0290(.A(mai_mai_n226_), .B(mai_mai_n318_), .Y(mai_mai_n319_));
  NAi41      m0291(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n320_));
  NO2        m0292(.A(mai_mai_n320_), .B(mai_mai_n150_), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n321_), .B(mai_mai_n319_), .Y(mai_mai_n322_));
  NAi31      m0294(.An(i), .B(l), .C(h), .Y(mai_mai_n323_));
  NO4        m0295(.A(mai_mai_n323_), .B(mai_mai_n150_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n324_));
  NA2        m0296(.A(e), .B(c), .Y(mai_mai_n325_));
  NO3        m0297(.A(mai_mai_n325_), .B(n), .C(d), .Y(mai_mai_n326_));
  NOi21      m0298(.An(f), .B(h), .Y(mai_mai_n327_));
  NA2        m0299(.A(mai_mai_n327_), .B(mai_mai_n116_), .Y(mai_mai_n328_));
  NO2        m0300(.A(mai_mai_n328_), .B(mai_mai_n214_), .Y(mai_mai_n329_));
  NAi31      m0301(.An(d), .B(e), .C(b), .Y(mai_mai_n330_));
  NO2        m0302(.A(mai_mai_n130_), .B(mai_mai_n330_), .Y(mai_mai_n331_));
  NA2        m0303(.A(mai_mai_n331_), .B(mai_mai_n329_), .Y(mai_mai_n332_));
  NAi41      m0304(.An(mai_mai_n324_), .B(mai_mai_n332_), .C(mai_mai_n322_), .D(mai_mai_n317_), .Y(mai_mai_n333_));
  NO4        m0305(.A(mai_mai_n320_), .B(mai_mai_n81_), .C(mai_mai_n72_), .D(mai_mai_n214_), .Y(mai_mai_n334_));
  NA2        m0306(.A(mai_mai_n250_), .B(mai_mai_n103_), .Y(mai_mai_n335_));
  OR2        m0307(.A(mai_mai_n335_), .B(mai_mai_n207_), .Y(mai_mai_n336_));
  NOi31      m0308(.An(l), .B(n), .C(m), .Y(mai_mai_n337_));
  NA2        m0309(.A(mai_mai_n337_), .B(mai_mai_n215_), .Y(mai_mai_n338_));
  NO2        m0310(.A(mai_mai_n338_), .B(mai_mai_n196_), .Y(mai_mai_n339_));
  NAi32      m0311(.An(mai_mai_n339_), .Bn(mai_mai_n334_), .C(mai_mai_n336_), .Y(mai_mai_n340_));
  NAi32      m0312(.An(m), .Bn(j), .C(k), .Y(mai_mai_n341_));
  NAi41      m0313(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n342_));
  OAI210     m0314(.A0(mai_mai_n211_), .A1(mai_mai_n341_), .B0(mai_mai_n342_), .Y(mai_mai_n343_));
  NOi31      m0315(.An(j), .B(m), .C(k), .Y(mai_mai_n344_));
  NO2        m0316(.A(mai_mai_n124_), .B(mai_mai_n344_), .Y(mai_mai_n345_));
  AN3        m0317(.A(h), .B(g), .C(f), .Y(mai_mai_n346_));
  NAi31      m0318(.An(mai_mai_n345_), .B(mai_mai_n346_), .C(mai_mai_n343_), .Y(mai_mai_n347_));
  NOi32      m0319(.An(m), .Bn(j), .C(l), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n348_), .B(mai_mai_n98_), .Y(mai_mai_n349_));
  NO2        m0321(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n350_));
  NO2        m0322(.A(mai_mai_n217_), .B(g), .Y(mai_mai_n351_));
  NA2        m0323(.A(mai_mai_n234_), .B(mai_mai_n81_), .Y(mai_mai_n352_));
  NA3        m0324(.A(mai_mai_n352_), .B(mai_mai_n346_), .C(mai_mai_n212_), .Y(mai_mai_n353_));
  NA2        m0325(.A(mai_mai_n353_), .B(mai_mai_n347_), .Y(mai_mai_n354_));
  NA3        m0326(.A(h), .B(g), .C(f), .Y(mai_mai_n355_));
  NO2        m0327(.A(mai_mai_n355_), .B(mai_mai_n77_), .Y(mai_mai_n356_));
  NA2        m0328(.A(mai_mai_n342_), .B(mai_mai_n211_), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n162_), .B(e), .Y(mai_mai_n358_));
  NO2        m0330(.A(mai_mai_n358_), .B(mai_mai_n41_), .Y(mai_mai_n359_));
  AOI220     m0331(.A0(mai_mai_n359_), .A1(mai_mai_n310_), .B0(mai_mai_n357_), .B1(mai_mai_n356_), .Y(mai_mai_n360_));
  NOi32      m0332(.An(j), .Bn(g), .C(i), .Y(mai_mai_n361_));
  NA3        m0333(.A(mai_mai_n361_), .B(mai_mai_n292_), .C(mai_mai_n112_), .Y(mai_mai_n362_));
  OR2        m0334(.A(mai_mai_n110_), .B(mai_mai_n362_), .Y(mai_mai_n363_));
  NOi32      m0335(.An(e), .Bn(b), .C(a), .Y(mai_mai_n364_));
  AN2        m0336(.A(l), .B(j), .Y(mai_mai_n365_));
  NO2        m0337(.A(mai_mai_n318_), .B(mai_mai_n365_), .Y(mai_mai_n366_));
  NO3        m0338(.A(mai_mai_n320_), .B(mai_mai_n72_), .C(mai_mai_n214_), .Y(mai_mai_n367_));
  NA2        m0339(.A(mai_mai_n210_), .B(mai_mai_n35_), .Y(mai_mai_n368_));
  AOI220     m0340(.A0(mai_mai_n368_), .A1(mai_mai_n364_), .B0(mai_mai_n367_), .B1(mai_mai_n366_), .Y(mai_mai_n369_));
  NA2        m0341(.A(mai_mai_n209_), .B(k), .Y(mai_mai_n370_));
  NA3        m0342(.A(m), .B(mai_mai_n111_), .C(mai_mai_n213_), .Y(mai_mai_n371_));
  NAi41      m0343(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n372_));
  NA2        m0344(.A(mai_mai_n51_), .B(mai_mai_n112_), .Y(mai_mai_n373_));
  NO2        m0345(.A(mai_mai_n373_), .B(mai_mai_n372_), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n374_), .B(b), .Y(mai_mai_n375_));
  NA4        m0347(.A(mai_mai_n375_), .B(mai_mai_n369_), .C(mai_mai_n363_), .D(mai_mai_n360_), .Y(mai_mai_n376_));
  NO4        m0348(.A(mai_mai_n376_), .B(mai_mai_n354_), .C(mai_mai_n340_), .D(mai_mai_n333_), .Y(mai_mai_n377_));
  NA4        m0349(.A(mai_mai_n377_), .B(mai_mai_n316_), .C(mai_mai_n269_), .D(mai_mai_n202_), .Y(mai10));
  NA3        m0350(.A(m), .B(k), .C(i), .Y(mai_mai_n379_));
  NO3        m0351(.A(mai_mai_n379_), .B(j), .C(mai_mai_n214_), .Y(mai_mai_n380_));
  NOi21      m0352(.An(e), .B(f), .Y(mai_mai_n381_));
  NO4        m0353(.A(mai_mai_n151_), .B(mai_mai_n381_), .C(n), .D(mai_mai_n109_), .Y(mai_mai_n382_));
  NAi31      m0354(.An(b), .B(f), .C(c), .Y(mai_mai_n383_));
  INV        m0355(.A(mai_mai_n383_), .Y(mai_mai_n384_));
  NOi32      m0356(.An(k), .Bn(h), .C(j), .Y(mai_mai_n385_));
  NA2        m0357(.A(mai_mai_n385_), .B(mai_mai_n221_), .Y(mai_mai_n386_));
  NA2        m0358(.A(mai_mai_n160_), .B(mai_mai_n386_), .Y(mai_mai_n387_));
  AOI220     m0359(.A0(mai_mai_n387_), .A1(mai_mai_n384_), .B0(mai_mai_n382_), .B1(mai_mai_n380_), .Y(mai_mai_n388_));
  AN2        m0360(.A(j), .B(h), .Y(mai_mai_n389_));
  NO3        m0361(.A(n), .B(m), .C(k), .Y(mai_mai_n390_));
  NA2        m0362(.A(mai_mai_n390_), .B(mai_mai_n389_), .Y(mai_mai_n391_));
  NO3        m0363(.A(mai_mai_n391_), .B(mai_mai_n151_), .C(mai_mai_n213_), .Y(mai_mai_n392_));
  OR2        m0364(.A(m), .B(k), .Y(mai_mai_n393_));
  NO2        m0365(.A(mai_mai_n175_), .B(mai_mai_n393_), .Y(mai_mai_n394_));
  NA4        m0366(.A(n), .B(f), .C(c), .D(mai_mai_n114_), .Y(mai_mai_n395_));
  NOi21      m0367(.An(mai_mai_n394_), .B(mai_mai_n395_), .Y(mai_mai_n396_));
  NOi32      m0368(.An(d), .Bn(a), .C(c), .Y(mai_mai_n397_));
  NA2        m0369(.A(mai_mai_n397_), .B(mai_mai_n183_), .Y(mai_mai_n398_));
  NAi21      m0370(.An(i), .B(g), .Y(mai_mai_n399_));
  NAi31      m0371(.An(k), .B(m), .C(j), .Y(mai_mai_n400_));
  NO2        m0372(.A(mai_mai_n396_), .B(mai_mai_n392_), .Y(mai_mai_n401_));
  NO2        m0373(.A(mai_mai_n395_), .B(mai_mai_n297_), .Y(mai_mai_n402_));
  NOi32      m0374(.An(f), .Bn(d), .C(c), .Y(mai_mai_n403_));
  AOI220     m0375(.A0(mai_mai_n403_), .A1(mai_mai_n308_), .B0(mai_mai_n402_), .B1(mai_mai_n215_), .Y(mai_mai_n404_));
  NA3        m0376(.A(mai_mai_n404_), .B(mai_mai_n401_), .C(mai_mai_n388_), .Y(mai_mai_n405_));
  NO2        m0377(.A(mai_mai_n59_), .B(mai_mai_n114_), .Y(mai_mai_n406_));
  NA2        m0378(.A(mai_mai_n250_), .B(mai_mai_n406_), .Y(mai_mai_n407_));
  INV        m0379(.A(e), .Y(mai_mai_n408_));
  NA2        m0380(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n409_));
  OAI220     m0381(.A0(mai_mai_n409_), .A1(mai_mai_n203_), .B0(mai_mai_n207_), .B1(mai_mai_n408_), .Y(mai_mai_n410_));
  AN2        m0382(.A(g), .B(e), .Y(mai_mai_n411_));
  NA3        m0383(.A(mai_mai_n411_), .B(mai_mai_n206_), .C(i), .Y(mai_mai_n412_));
  INV        m0384(.A(mai_mai_n412_), .Y(mai_mai_n413_));
  NO2        m0385(.A(mai_mai_n101_), .B(mai_mai_n408_), .Y(mai_mai_n414_));
  NO3        m0386(.A(mai_mai_n414_), .B(mai_mai_n413_), .C(mai_mai_n410_), .Y(mai_mai_n415_));
  NOi32      m0387(.An(h), .Bn(e), .C(g), .Y(mai_mai_n416_));
  NA3        m0388(.A(mai_mai_n416_), .B(mai_mai_n294_), .C(m), .Y(mai_mai_n417_));
  NOi21      m0389(.An(g), .B(h), .Y(mai_mai_n418_));
  AN3        m0390(.A(m), .B(l), .C(i), .Y(mai_mai_n419_));
  NA3        m0391(.A(mai_mai_n419_), .B(mai_mai_n418_), .C(e), .Y(mai_mai_n420_));
  AN3        m0392(.A(h), .B(g), .C(e), .Y(mai_mai_n421_));
  NA2        m0393(.A(mai_mai_n421_), .B(mai_mai_n98_), .Y(mai_mai_n422_));
  AN3        m0394(.A(mai_mai_n422_), .B(mai_mai_n420_), .C(mai_mai_n417_), .Y(mai_mai_n423_));
  AOI210     m0395(.A0(mai_mai_n423_), .A1(mai_mai_n415_), .B0(mai_mai_n407_), .Y(mai_mai_n424_));
  NA3        m0396(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n425_));
  NO2        m0397(.A(mai_mai_n425_), .B(mai_mai_n407_), .Y(mai_mai_n426_));
  NA3        m0398(.A(mai_mai_n397_), .B(mai_mai_n183_), .C(mai_mai_n86_), .Y(mai_mai_n427_));
  NAi31      m0399(.An(b), .B(c), .C(a), .Y(mai_mai_n428_));
  NO2        m0400(.A(mai_mai_n428_), .B(n), .Y(mai_mai_n429_));
  OAI210     m0401(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n430_));
  NO2        m0402(.A(mai_mai_n430_), .B(mai_mai_n147_), .Y(mai_mai_n431_));
  NA2        m0403(.A(mai_mai_n431_), .B(mai_mai_n429_), .Y(mai_mai_n432_));
  INV        m0404(.A(mai_mai_n432_), .Y(mai_mai_n433_));
  NO4        m0405(.A(mai_mai_n433_), .B(mai_mai_n426_), .C(mai_mai_n424_), .D(mai_mai_n405_), .Y(mai_mai_n434_));
  NA2        m0406(.A(i), .B(g), .Y(mai_mai_n435_));
  NO3        m0407(.A(mai_mai_n278_), .B(mai_mai_n435_), .C(c), .Y(mai_mai_n436_));
  NOi21      m0408(.An(a), .B(n), .Y(mai_mai_n437_));
  NOi21      m0409(.An(d), .B(c), .Y(mai_mai_n438_));
  NA2        m0410(.A(mai_mai_n438_), .B(mai_mai_n437_), .Y(mai_mai_n439_));
  NA3        m0411(.A(i), .B(g), .C(f), .Y(mai_mai_n440_));
  OR2        m0412(.A(mai_mai_n440_), .B(mai_mai_n71_), .Y(mai_mai_n441_));
  NA3        m0413(.A(mai_mai_n419_), .B(mai_mai_n418_), .C(mai_mai_n183_), .Y(mai_mai_n442_));
  AOI210     m0414(.A0(mai_mai_n442_), .A1(mai_mai_n441_), .B0(mai_mai_n439_), .Y(mai_mai_n443_));
  AOI210     m0415(.A0(mai_mai_n436_), .A1(mai_mai_n293_), .B0(mai_mai_n443_), .Y(mai_mai_n444_));
  OR2        m0416(.A(n), .B(m), .Y(mai_mai_n445_));
  NO2        m0417(.A(mai_mai_n445_), .B(mai_mai_n152_), .Y(mai_mai_n446_));
  NO2        m0418(.A(mai_mai_n184_), .B(mai_mai_n147_), .Y(mai_mai_n447_));
  OAI210     m0419(.A0(mai_mai_n446_), .A1(mai_mai_n177_), .B0(mai_mai_n447_), .Y(mai_mai_n448_));
  INV        m0420(.A(mai_mai_n373_), .Y(mai_mai_n449_));
  NA3        m0421(.A(mai_mai_n449_), .B(mai_mai_n364_), .C(d), .Y(mai_mai_n450_));
  NO2        m0422(.A(mai_mai_n428_), .B(mai_mai_n49_), .Y(mai_mai_n451_));
  NO3        m0423(.A(mai_mai_n66_), .B(mai_mai_n111_), .C(e), .Y(mai_mai_n452_));
  NAi21      m0424(.An(k), .B(j), .Y(mai_mai_n453_));
  NA2        m0425(.A(mai_mai_n252_), .B(mai_mai_n453_), .Y(mai_mai_n454_));
  NA3        m0426(.A(mai_mai_n454_), .B(mai_mai_n452_), .C(mai_mai_n451_), .Y(mai_mai_n455_));
  NAi21      m0427(.An(e), .B(d), .Y(mai_mai_n456_));
  INV        m0428(.A(mai_mai_n456_), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n253_), .B(mai_mai_n213_), .Y(mai_mai_n458_));
  NA3        m0430(.A(mai_mai_n458_), .B(mai_mai_n457_), .C(mai_mai_n227_), .Y(mai_mai_n459_));
  NA4        m0431(.A(mai_mai_n459_), .B(mai_mai_n455_), .C(mai_mai_n450_), .D(mai_mai_n448_), .Y(mai_mai_n460_));
  NO2        m0432(.A(mai_mai_n338_), .B(mai_mai_n213_), .Y(mai_mai_n461_));
  NA2        m0433(.A(mai_mai_n461_), .B(mai_mai_n457_), .Y(mai_mai_n462_));
  NOi31      m0434(.An(n), .B(m), .C(k), .Y(mai_mai_n463_));
  AOI220     m0435(.A0(mai_mai_n463_), .A1(mai_mai_n389_), .B0(mai_mai_n221_), .B1(mai_mai_n50_), .Y(mai_mai_n464_));
  NAi31      m0436(.An(g), .B(f), .C(c), .Y(mai_mai_n465_));
  OR3        m0437(.A(mai_mai_n465_), .B(mai_mai_n464_), .C(e), .Y(mai_mai_n466_));
  NA3        m0438(.A(mai_mai_n466_), .B(mai_mai_n462_), .C(mai_mai_n309_), .Y(mai_mai_n467_));
  NOi41      m0439(.An(mai_mai_n444_), .B(mai_mai_n467_), .C(mai_mai_n460_), .D(mai_mai_n267_), .Y(mai_mai_n468_));
  NOi32      m0440(.An(c), .Bn(a), .C(b), .Y(mai_mai_n469_));
  NA2        m0441(.A(mai_mai_n469_), .B(mai_mai_n112_), .Y(mai_mai_n470_));
  INV        m0442(.A(mai_mai_n276_), .Y(mai_mai_n471_));
  AN2        m0443(.A(e), .B(d), .Y(mai_mai_n472_));
  NA2        m0444(.A(mai_mai_n472_), .B(mai_mai_n471_), .Y(mai_mai_n473_));
  INV        m0445(.A(mai_mai_n147_), .Y(mai_mai_n474_));
  NO2        m0446(.A(mai_mai_n129_), .B(mai_mai_n41_), .Y(mai_mai_n475_));
  NO2        m0447(.A(mai_mai_n66_), .B(e), .Y(mai_mai_n476_));
  NOi31      m0448(.An(j), .B(k), .C(i), .Y(mai_mai_n477_));
  NOi21      m0449(.An(mai_mai_n165_), .B(mai_mai_n477_), .Y(mai_mai_n478_));
  NA4        m0450(.A(mai_mai_n323_), .B(mai_mai_n478_), .C(mai_mai_n261_), .D(mai_mai_n117_), .Y(mai_mai_n479_));
  AOI220     m0451(.A0(mai_mai_n479_), .A1(mai_mai_n476_), .B0(mai_mai_n475_), .B1(mai_mai_n474_), .Y(mai_mai_n480_));
  AOI210     m0452(.A0(mai_mai_n480_), .A1(mai_mai_n473_), .B0(mai_mai_n470_), .Y(mai_mai_n481_));
  INV        m0453(.A(mai_mai_n208_), .Y(mai_mai_n482_));
  NOi21      m0454(.An(a), .B(b), .Y(mai_mai_n483_));
  NA3        m0455(.A(e), .B(d), .C(c), .Y(mai_mai_n484_));
  NAi21      m0456(.An(mai_mai_n484_), .B(mai_mai_n483_), .Y(mai_mai_n485_));
  NO2        m0457(.A(mai_mai_n427_), .B(mai_mai_n207_), .Y(mai_mai_n486_));
  NOi21      m0458(.An(mai_mai_n485_), .B(mai_mai_n486_), .Y(mai_mai_n487_));
  AOI210     m0459(.A0(mai_mai_n270_), .A1(mai_mai_n482_), .B0(mai_mai_n487_), .Y(mai_mai_n488_));
  NO4        m0460(.A(mai_mai_n190_), .B(mai_mai_n102_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n489_));
  NA2        m0461(.A(mai_mai_n384_), .B(mai_mai_n153_), .Y(mai_mai_n490_));
  OR2        m0462(.A(k), .B(j), .Y(mai_mai_n491_));
  NA2        m0463(.A(l), .B(k), .Y(mai_mai_n492_));
  NA3        m0464(.A(mai_mai_n492_), .B(mai_mai_n491_), .C(mai_mai_n221_), .Y(mai_mai_n493_));
  AOI210     m0465(.A0(mai_mai_n234_), .A1(mai_mai_n341_), .B0(mai_mai_n86_), .Y(mai_mai_n494_));
  NOi21      m0466(.An(mai_mai_n493_), .B(mai_mai_n494_), .Y(mai_mai_n495_));
  OR3        m0467(.A(mai_mai_n495_), .B(mai_mai_n143_), .C(mai_mai_n133_), .Y(mai_mai_n496_));
  NA2        m0468(.A(mai_mai_n281_), .B(mai_mai_n126_), .Y(mai_mai_n497_));
  NA2        m0469(.A(mai_mai_n397_), .B(mai_mai_n112_), .Y(mai_mai_n498_));
  NO4        m0470(.A(mai_mai_n498_), .B(mai_mai_n95_), .C(mai_mai_n111_), .D(e), .Y(mai_mai_n499_));
  NO3        m0471(.A(mai_mai_n427_), .B(mai_mai_n93_), .C(mai_mai_n129_), .Y(mai_mai_n500_));
  NO4        m0472(.A(mai_mai_n500_), .B(mai_mai_n499_), .C(mai_mai_n497_), .D(mai_mai_n324_), .Y(mai_mai_n501_));
  NA3        m0473(.A(mai_mai_n501_), .B(mai_mai_n496_), .C(mai_mai_n490_), .Y(mai_mai_n502_));
  NO4        m0474(.A(mai_mai_n502_), .B(mai_mai_n489_), .C(mai_mai_n488_), .D(mai_mai_n481_), .Y(mai_mai_n503_));
  NA2        m0475(.A(mai_mai_n70_), .B(mai_mai_n67_), .Y(mai_mai_n504_));
  NOi21      m0476(.An(d), .B(e), .Y(mai_mai_n505_));
  NAi31      m0477(.An(j), .B(l), .C(i), .Y(mai_mai_n506_));
  OAI210     m0478(.A0(mai_mai_n506_), .A1(mai_mai_n130_), .B0(mai_mai_n102_), .Y(mai_mai_n507_));
  NO3        m0479(.A(mai_mai_n398_), .B(mai_mai_n349_), .C(mai_mai_n204_), .Y(mai_mai_n508_));
  NO2        m0480(.A(mai_mai_n398_), .B(mai_mai_n373_), .Y(mai_mai_n509_));
  NO4        m0481(.A(mai_mai_n509_), .B(mai_mai_n508_), .C(mai_mai_n186_), .D(mai_mai_n306_), .Y(mai_mai_n510_));
  NA3        m0482(.A(mai_mai_n510_), .B(mai_mai_n504_), .C(mai_mai_n244_), .Y(mai_mai_n511_));
  OAI210     m0483(.A0(mai_mai_n125_), .A1(mai_mai_n124_), .B0(n), .Y(mai_mai_n512_));
  NO2        m0484(.A(mai_mai_n512_), .B(mai_mai_n129_), .Y(mai_mai_n513_));
  OA210      m0485(.A0(mai_mai_n246_), .A1(mai_mai_n513_), .B0(mai_mai_n195_), .Y(mai_mai_n514_));
  XO2        m0486(.A(i), .B(h), .Y(mai_mai_n515_));
  NA3        m0487(.A(mai_mai_n515_), .B(mai_mai_n159_), .C(n), .Y(mai_mai_n516_));
  NAi41      m0488(.An(mai_mai_n298_), .B(mai_mai_n516_), .C(mai_mai_n464_), .D(mai_mai_n386_), .Y(mai_mai_n517_));
  NOi32      m0489(.An(mai_mai_n517_), .Bn(mai_mai_n476_), .C(mai_mai_n272_), .Y(mai_mai_n518_));
  NAi31      m0490(.An(c), .B(f), .C(d), .Y(mai_mai_n519_));
  AOI210     m0491(.A0(mai_mai_n282_), .A1(mai_mai_n198_), .B0(mai_mai_n519_), .Y(mai_mai_n520_));
  NOi21      m0492(.An(mai_mai_n84_), .B(mai_mai_n520_), .Y(mai_mai_n521_));
  NA3        m0493(.A(mai_mai_n382_), .B(mai_mai_n98_), .C(mai_mai_n97_), .Y(mai_mai_n522_));
  NA2        m0494(.A(mai_mai_n228_), .B(mai_mai_n108_), .Y(mai_mai_n523_));
  AOI210     m0495(.A0(mai_mai_n523_), .A1(mai_mai_n182_), .B0(mai_mai_n519_), .Y(mai_mai_n524_));
  AOI210     m0496(.A0(mai_mai_n362_), .A1(mai_mai_n35_), .B0(mai_mai_n485_), .Y(mai_mai_n525_));
  NOi31      m0497(.An(mai_mai_n522_), .B(mai_mai_n525_), .C(mai_mai_n524_), .Y(mai_mai_n526_));
  AO220      m0498(.A0(mai_mai_n290_), .A1(mai_mai_n264_), .B0(mai_mai_n166_), .B1(mai_mai_n67_), .Y(mai_mai_n527_));
  NA3        m0499(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n528_));
  NAi31      m0500(.An(mai_mai_n527_), .B(mai_mai_n526_), .C(mai_mai_n521_), .Y(mai_mai_n529_));
  NO4        m0501(.A(mai_mai_n529_), .B(mai_mai_n518_), .C(mai_mai_n514_), .D(mai_mai_n511_), .Y(mai_mai_n530_));
  NA4        m0502(.A(mai_mai_n530_), .B(mai_mai_n503_), .C(mai_mai_n468_), .D(mai_mai_n434_), .Y(mai11));
  NO2        m0503(.A(mai_mai_n73_), .B(f), .Y(mai_mai_n532_));
  NA2        m0504(.A(j), .B(g), .Y(mai_mai_n533_));
  NAi31      m0505(.An(i), .B(m), .C(l), .Y(mai_mai_n534_));
  NA3        m0506(.A(m), .B(k), .C(j), .Y(mai_mai_n535_));
  OAI220     m0507(.A0(mai_mai_n535_), .A1(mai_mai_n129_), .B0(mai_mai_n534_), .B1(mai_mai_n533_), .Y(mai_mai_n536_));
  NA2        m0508(.A(mai_mai_n536_), .B(mai_mai_n532_), .Y(mai_mai_n537_));
  NOi32      m0509(.An(e), .Bn(b), .C(f), .Y(mai_mai_n538_));
  NA2        m0510(.A(mai_mai_n260_), .B(mai_mai_n112_), .Y(mai_mai_n539_));
  NA2        m0511(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n540_));
  NO2        m0512(.A(mai_mai_n540_), .B(mai_mai_n300_), .Y(mai_mai_n541_));
  NAi31      m0513(.An(d), .B(e), .C(a), .Y(mai_mai_n542_));
  NA2        m0514(.A(mai_mai_n541_), .B(mai_mai_n538_), .Y(mai_mai_n543_));
  NAi41      m0515(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n544_));
  AN2        m0516(.A(mai_mai_n544_), .B(mai_mai_n372_), .Y(mai_mai_n545_));
  AOI210     m0517(.A0(mai_mai_n545_), .A1(mai_mai_n398_), .B0(mai_mai_n273_), .Y(mai_mai_n546_));
  NA2        m0518(.A(j), .B(i), .Y(mai_mai_n547_));
  NAi31      m0519(.An(n), .B(m), .C(k), .Y(mai_mai_n548_));
  NO3        m0520(.A(mai_mai_n548_), .B(mai_mai_n547_), .C(mai_mai_n111_), .Y(mai_mai_n549_));
  NO4        m0521(.A(n), .B(d), .C(mai_mai_n114_), .D(a), .Y(mai_mai_n550_));
  OR2        m0522(.A(n), .B(c), .Y(mai_mai_n551_));
  NO2        m0523(.A(mai_mai_n551_), .B(mai_mai_n149_), .Y(mai_mai_n552_));
  NO2        m0524(.A(mai_mai_n552_), .B(mai_mai_n550_), .Y(mai_mai_n553_));
  NOi32      m0525(.An(g), .Bn(f), .C(i), .Y(mai_mai_n554_));
  AOI220     m0526(.A0(mai_mai_n554_), .A1(mai_mai_n100_), .B0(mai_mai_n536_), .B1(f), .Y(mai_mai_n555_));
  NO2        m0527(.A(mai_mai_n276_), .B(mai_mai_n49_), .Y(mai_mai_n556_));
  NO2        m0528(.A(mai_mai_n555_), .B(mai_mai_n553_), .Y(mai_mai_n557_));
  AOI210     m0529(.A0(mai_mai_n549_), .A1(mai_mai_n546_), .B0(mai_mai_n557_), .Y(mai_mai_n558_));
  NA2        m0530(.A(mai_mai_n139_), .B(mai_mai_n34_), .Y(mai_mai_n559_));
  OAI220     m0531(.A0(mai_mai_n559_), .A1(m), .B0(mai_mai_n540_), .B1(mai_mai_n234_), .Y(mai_mai_n560_));
  NOi41      m0532(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n561_));
  NAi32      m0533(.An(e), .Bn(b), .C(c), .Y(mai_mai_n562_));
  OR2        m0534(.A(mai_mai_n562_), .B(mai_mai_n86_), .Y(mai_mai_n563_));
  AN2        m0535(.A(mai_mai_n342_), .B(mai_mai_n320_), .Y(mai_mai_n564_));
  NA2        m0536(.A(mai_mai_n564_), .B(mai_mai_n563_), .Y(mai_mai_n565_));
  OA210      m0537(.A0(mai_mai_n565_), .A1(mai_mai_n561_), .B0(mai_mai_n560_), .Y(mai_mai_n566_));
  OAI220     m0538(.A0(mai_mai_n400_), .A1(mai_mai_n399_), .B0(mai_mai_n534_), .B1(mai_mai_n533_), .Y(mai_mai_n567_));
  NAi31      m0539(.An(d), .B(c), .C(a), .Y(mai_mai_n568_));
  NO2        m0540(.A(mai_mai_n568_), .B(n), .Y(mai_mai_n569_));
  NA3        m0541(.A(mai_mai_n569_), .B(mai_mai_n567_), .C(e), .Y(mai_mai_n570_));
  NO3        m0542(.A(mai_mai_n62_), .B(mai_mai_n49_), .C(mai_mai_n214_), .Y(mai_mai_n571_));
  INV        m0543(.A(mai_mai_n570_), .Y(mai_mai_n572_));
  NO2        m0544(.A(mai_mai_n278_), .B(n), .Y(mai_mai_n573_));
  NO2        m0545(.A(mai_mai_n429_), .B(mai_mai_n573_), .Y(mai_mai_n574_));
  NA2        m0546(.A(mai_mai_n567_), .B(f), .Y(mai_mai_n575_));
  NAi32      m0547(.An(d), .Bn(a), .C(b), .Y(mai_mai_n576_));
  NO2        m0548(.A(mai_mai_n576_), .B(mai_mai_n49_), .Y(mai_mai_n577_));
  NA2        m0549(.A(h), .B(f), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n578_), .B(mai_mai_n95_), .Y(mai_mai_n579_));
  NO3        m0551(.A(mai_mai_n178_), .B(mai_mai_n175_), .C(g), .Y(mai_mai_n580_));
  AOI220     m0552(.A0(mai_mai_n580_), .A1(mai_mai_n58_), .B0(mai_mai_n579_), .B1(mai_mai_n577_), .Y(mai_mai_n581_));
  OAI210     m0553(.A0(mai_mai_n575_), .A1(mai_mai_n574_), .B0(mai_mai_n581_), .Y(mai_mai_n582_));
  AN3        m0554(.A(j), .B(h), .C(g), .Y(mai_mai_n583_));
  NO2        m0555(.A(mai_mai_n146_), .B(c), .Y(mai_mai_n584_));
  NA3        m0556(.A(mai_mai_n584_), .B(mai_mai_n583_), .C(mai_mai_n463_), .Y(mai_mai_n585_));
  NA3        m0557(.A(f), .B(d), .C(b), .Y(mai_mai_n586_));
  NO4        m0558(.A(mai_mai_n586_), .B(mai_mai_n178_), .C(mai_mai_n175_), .D(g), .Y(mai_mai_n587_));
  NAi21      m0559(.An(mai_mai_n587_), .B(mai_mai_n585_), .Y(mai_mai_n588_));
  NO4        m0560(.A(mai_mai_n588_), .B(mai_mai_n582_), .C(mai_mai_n572_), .D(mai_mai_n566_), .Y(mai_mai_n589_));
  AN4        m0561(.A(mai_mai_n589_), .B(mai_mai_n558_), .C(mai_mai_n543_), .D(mai_mai_n537_), .Y(mai_mai_n590_));
  INV        m0562(.A(k), .Y(mai_mai_n591_));
  NA3        m0563(.A(l), .B(mai_mai_n591_), .C(i), .Y(mai_mai_n592_));
  INV        m0564(.A(mai_mai_n592_), .Y(mai_mai_n593_));
  NA4        m0565(.A(mai_mai_n397_), .B(mai_mai_n418_), .C(mai_mai_n183_), .D(mai_mai_n112_), .Y(mai_mai_n594_));
  NAi32      m0566(.An(h), .Bn(f), .C(g), .Y(mai_mai_n595_));
  NAi41      m0567(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n596_));
  OAI210     m0568(.A0(mai_mai_n542_), .A1(n), .B0(mai_mai_n596_), .Y(mai_mai_n597_));
  NAi31      m0569(.An(h), .B(g), .C(f), .Y(mai_mai_n598_));
  OR3        m0570(.A(mai_mai_n598_), .B(mai_mai_n278_), .C(mai_mai_n49_), .Y(mai_mai_n599_));
  NA4        m0571(.A(mai_mai_n418_), .B(mai_mai_n119_), .C(mai_mai_n112_), .D(e), .Y(mai_mai_n600_));
  AN2        m0572(.A(mai_mai_n600_), .B(mai_mai_n599_), .Y(mai_mai_n601_));
  BUFFER     m0573(.A(mai_mai_n601_), .Y(mai_mai_n602_));
  NO3        m0574(.A(mai_mai_n595_), .B(mai_mai_n73_), .C(mai_mai_n75_), .Y(mai_mai_n603_));
  NAi31      m0575(.An(mai_mai_n603_), .B(mai_mai_n602_), .C(mai_mai_n594_), .Y(mai_mai_n604_));
  NAi31      m0576(.An(f), .B(h), .C(g), .Y(mai_mai_n605_));
  NO4        m0577(.A(mai_mai_n311_), .B(mai_mai_n605_), .C(mai_mai_n73_), .D(mai_mai_n75_), .Y(mai_mai_n606_));
  NOi32      m0578(.An(b), .Bn(a), .C(c), .Y(mai_mai_n607_));
  NOi41      m0579(.An(mai_mai_n607_), .B(mai_mai_n355_), .C(mai_mai_n69_), .D(mai_mai_n115_), .Y(mai_mai_n608_));
  OR2        m0580(.A(mai_mai_n608_), .B(mai_mai_n606_), .Y(mai_mai_n609_));
  NOi32      m0581(.An(d), .Bn(a), .C(e), .Y(mai_mai_n610_));
  NA2        m0582(.A(mai_mai_n610_), .B(mai_mai_n112_), .Y(mai_mai_n611_));
  NO2        m0583(.A(n), .B(c), .Y(mai_mai_n612_));
  NOi32      m0584(.An(e), .Bn(a), .C(d), .Y(mai_mai_n613_));
  AOI210     m0585(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n613_), .Y(mai_mai_n614_));
  AOI210     m0586(.A0(mai_mai_n604_), .A1(mai_mai_n593_), .B0(mai_mai_n609_), .Y(mai_mai_n615_));
  NO3        m0587(.A(mai_mai_n318_), .B(mai_mai_n61_), .C(n), .Y(mai_mai_n616_));
  NA3        m0588(.A(mai_mai_n519_), .B(mai_mai_n173_), .C(mai_mai_n172_), .Y(mai_mai_n617_));
  NA2        m0589(.A(mai_mai_n465_), .B(mai_mai_n231_), .Y(mai_mai_n618_));
  OR2        m0590(.A(mai_mai_n618_), .B(mai_mai_n617_), .Y(mai_mai_n619_));
  NA2        m0591(.A(mai_mai_n76_), .B(mai_mai_n112_), .Y(mai_mai_n620_));
  NO2        m0592(.A(mai_mai_n620_), .B(mai_mai_n45_), .Y(mai_mai_n621_));
  AOI220     m0593(.A0(mai_mai_n621_), .A1(mai_mai_n546_), .B0(mai_mai_n619_), .B1(mai_mai_n616_), .Y(mai_mai_n622_));
  NO2        m0594(.A(mai_mai_n622_), .B(mai_mai_n89_), .Y(mai_mai_n623_));
  NA3        m0595(.A(mai_mai_n561_), .B(mai_mai_n344_), .C(mai_mai_n46_), .Y(mai_mai_n624_));
  NOi32      m0596(.An(e), .Bn(c), .C(f), .Y(mai_mai_n625_));
  NOi21      m0597(.An(f), .B(g), .Y(mai_mai_n626_));
  NO2        m0598(.A(mai_mai_n626_), .B(mai_mai_n211_), .Y(mai_mai_n627_));
  AOI220     m0599(.A0(mai_mai_n627_), .A1(mai_mai_n394_), .B0(mai_mai_n625_), .B1(mai_mai_n177_), .Y(mai_mai_n628_));
  NA3        m0600(.A(mai_mai_n628_), .B(mai_mai_n624_), .C(mai_mai_n180_), .Y(mai_mai_n629_));
  AOI210     m0601(.A0(mai_mai_n545_), .A1(mai_mai_n398_), .B0(mai_mai_n299_), .Y(mai_mai_n630_));
  NA2        m0602(.A(mai_mai_n630_), .B(mai_mai_n265_), .Y(mai_mai_n631_));
  NOi21      m0603(.An(j), .B(l), .Y(mai_mai_n632_));
  NAi21      m0604(.An(k), .B(h), .Y(mai_mai_n633_));
  NO2        m0605(.A(mai_mai_n633_), .B(mai_mai_n263_), .Y(mai_mai_n634_));
  NOi31      m0606(.An(m), .B(n), .C(k), .Y(mai_mai_n635_));
  NA2        m0607(.A(mai_mai_n632_), .B(mai_mai_n635_), .Y(mai_mai_n636_));
  AOI210     m0608(.A0(mai_mai_n398_), .A1(mai_mai_n372_), .B0(mai_mai_n299_), .Y(mai_mai_n637_));
  NAi21      m0609(.An(mai_mai_n636_), .B(mai_mai_n637_), .Y(mai_mai_n638_));
  NO2        m0610(.A(mai_mai_n278_), .B(mai_mai_n49_), .Y(mai_mai_n639_));
  NA2        m0611(.A(mai_mai_n639_), .B(mai_mai_n579_), .Y(mai_mai_n640_));
  NA3        m0612(.A(mai_mai_n640_), .B(mai_mai_n638_), .C(mai_mai_n631_), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n108_), .B(mai_mai_n36_), .Y(mai_mai_n642_));
  NO2        m0614(.A(k), .B(mai_mai_n214_), .Y(mai_mai_n643_));
  INV        m0615(.A(mai_mai_n364_), .Y(mai_mai_n644_));
  NO2        m0616(.A(mai_mai_n644_), .B(n), .Y(mai_mai_n645_));
  NAi31      m0617(.An(mai_mai_n642_), .B(mai_mai_n645_), .C(mai_mai_n643_), .Y(mai_mai_n646_));
  NO2        m0618(.A(mai_mai_n540_), .B(mai_mai_n178_), .Y(mai_mai_n647_));
  NA3        m0619(.A(mai_mai_n562_), .B(mai_mai_n272_), .C(mai_mai_n144_), .Y(mai_mai_n648_));
  NA2        m0620(.A(mai_mai_n515_), .B(mai_mai_n159_), .Y(mai_mai_n649_));
  NO3        m0621(.A(mai_mai_n395_), .B(mai_mai_n649_), .C(mai_mai_n89_), .Y(mai_mai_n650_));
  AOI210     m0622(.A0(mai_mai_n648_), .A1(mai_mai_n647_), .B0(mai_mai_n650_), .Y(mai_mai_n651_));
  AN3        m0623(.A(f), .B(d), .C(b), .Y(mai_mai_n652_));
  OAI210     m0624(.A0(mai_mai_n652_), .A1(mai_mai_n128_), .B0(n), .Y(mai_mai_n653_));
  NA3        m0625(.A(mai_mai_n515_), .B(mai_mai_n159_), .C(mai_mai_n214_), .Y(mai_mai_n654_));
  AOI210     m0626(.A0(mai_mai_n653_), .A1(mai_mai_n233_), .B0(mai_mai_n654_), .Y(mai_mai_n655_));
  NAi31      m0627(.An(m), .B(n), .C(k), .Y(mai_mai_n656_));
  INV        m0628(.A(mai_mai_n251_), .Y(mai_mai_n657_));
  OAI210     m0629(.A0(mai_mai_n657_), .A1(mai_mai_n655_), .B0(j), .Y(mai_mai_n658_));
  NA3        m0630(.A(mai_mai_n658_), .B(mai_mai_n651_), .C(mai_mai_n646_), .Y(mai_mai_n659_));
  NO4        m0631(.A(mai_mai_n659_), .B(mai_mai_n641_), .C(mai_mai_n629_), .D(mai_mai_n623_), .Y(mai_mai_n660_));
  NA2        m0632(.A(mai_mai_n382_), .B(mai_mai_n162_), .Y(mai_mai_n661_));
  NAi31      m0633(.An(g), .B(h), .C(f), .Y(mai_mai_n662_));
  OR3        m0634(.A(mai_mai_n662_), .B(mai_mai_n278_), .C(n), .Y(mai_mai_n663_));
  OA210      m0635(.A0(mai_mai_n542_), .A1(n), .B0(mai_mai_n596_), .Y(mai_mai_n664_));
  NA3        m0636(.A(mai_mai_n416_), .B(mai_mai_n119_), .C(mai_mai_n86_), .Y(mai_mai_n665_));
  OAI210     m0637(.A0(mai_mai_n664_), .A1(mai_mai_n92_), .B0(mai_mai_n665_), .Y(mai_mai_n666_));
  NOi21      m0638(.An(mai_mai_n663_), .B(mai_mai_n666_), .Y(mai_mai_n667_));
  AOI210     m0639(.A0(mai_mai_n667_), .A1(mai_mai_n661_), .B0(mai_mai_n535_), .Y(mai_mai_n668_));
  NO3        m0640(.A(g), .B(mai_mai_n213_), .C(mai_mai_n56_), .Y(mai_mai_n669_));
  NAi21      m0641(.An(h), .B(j), .Y(mai_mai_n670_));
  NO2        m0642(.A(mai_mai_n523_), .B(mai_mai_n89_), .Y(mai_mai_n671_));
  OAI210     m0643(.A0(mai_mai_n671_), .A1(mai_mai_n394_), .B0(mai_mai_n669_), .Y(mai_mai_n672_));
  OR2        m0644(.A(mai_mai_n73_), .B(mai_mai_n75_), .Y(mai_mai_n673_));
  NA3        m0645(.A(mai_mai_n532_), .B(mai_mai_n100_), .C(mai_mai_n99_), .Y(mai_mai_n674_));
  AN2        m0646(.A(h), .B(f), .Y(mai_mai_n675_));
  NA2        m0647(.A(mai_mai_n675_), .B(mai_mai_n37_), .Y(mai_mai_n676_));
  NA2        m0648(.A(mai_mai_n100_), .B(mai_mai_n46_), .Y(mai_mai_n677_));
  OAI220     m0649(.A0(mai_mai_n677_), .A1(mai_mai_n335_), .B0(mai_mai_n676_), .B1(mai_mai_n470_), .Y(mai_mai_n678_));
  AOI210     m0650(.A0(mai_mai_n576_), .A1(mai_mai_n428_), .B0(mai_mai_n49_), .Y(mai_mai_n679_));
  OAI220     m0651(.A0(mai_mai_n598_), .A1(mai_mai_n592_), .B0(mai_mai_n328_), .B1(mai_mai_n533_), .Y(mai_mai_n680_));
  AOI210     m0652(.A0(mai_mai_n680_), .A1(mai_mai_n679_), .B0(mai_mai_n678_), .Y(mai_mai_n681_));
  NA3        m0653(.A(mai_mai_n681_), .B(mai_mai_n674_), .C(mai_mai_n672_), .Y(mai_mai_n682_));
  NO2        m0654(.A(mai_mai_n252_), .B(f), .Y(mai_mai_n683_));
  NO2        m0655(.A(mai_mai_n626_), .B(mai_mai_n61_), .Y(mai_mai_n684_));
  NO3        m0656(.A(mai_mai_n684_), .B(mai_mai_n683_), .C(mai_mai_n34_), .Y(mai_mai_n685_));
  NA2        m0657(.A(mai_mai_n331_), .B(mai_mai_n139_), .Y(mai_mai_n686_));
  NA2        m0658(.A(mai_mai_n130_), .B(mai_mai_n49_), .Y(mai_mai_n687_));
  AOI220     m0659(.A0(mai_mai_n687_), .A1(mai_mai_n538_), .B0(mai_mai_n364_), .B1(mai_mai_n112_), .Y(mai_mai_n688_));
  OA220      m0660(.A0(mai_mai_n688_), .A1(mai_mai_n559_), .B0(mai_mai_n362_), .B1(mai_mai_n110_), .Y(mai_mai_n689_));
  OAI210     m0661(.A0(mai_mai_n686_), .A1(mai_mai_n685_), .B0(mai_mai_n689_), .Y(mai_mai_n690_));
  NO3        m0662(.A(mai_mai_n403_), .B(mai_mai_n195_), .C(mai_mai_n194_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n691_), .B(mai_mai_n231_), .Y(mai_mai_n692_));
  NA3        m0664(.A(mai_mai_n692_), .B(mai_mai_n254_), .C(j), .Y(mai_mai_n693_));
  NO3        m0665(.A(mai_mai_n465_), .B(mai_mai_n175_), .C(i), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n469_), .B(mai_mai_n86_), .Y(mai_mai_n695_));
  NO4        m0667(.A(mai_mai_n535_), .B(mai_mai_n695_), .C(mai_mai_n129_), .D(mai_mai_n213_), .Y(mai_mai_n696_));
  INV        m0668(.A(mai_mai_n696_), .Y(mai_mai_n697_));
  NA4        m0669(.A(mai_mai_n697_), .B(mai_mai_n693_), .C(mai_mai_n522_), .D(mai_mai_n401_), .Y(mai_mai_n698_));
  NO4        m0670(.A(mai_mai_n698_), .B(mai_mai_n690_), .C(mai_mai_n682_), .D(mai_mai_n668_), .Y(mai_mai_n699_));
  NA4        m0671(.A(mai_mai_n699_), .B(mai_mai_n660_), .C(mai_mai_n615_), .D(mai_mai_n590_), .Y(mai08));
  NO2        m0672(.A(k), .B(h), .Y(mai_mai_n701_));
  AO210      m0673(.A0(mai_mai_n252_), .A1(mai_mai_n453_), .B0(mai_mai_n701_), .Y(mai_mai_n702_));
  NO2        m0674(.A(mai_mai_n702_), .B(mai_mai_n297_), .Y(mai_mai_n703_));
  NA2        m0675(.A(mai_mai_n625_), .B(mai_mai_n86_), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n704_), .B(mai_mai_n465_), .Y(mai_mai_n705_));
  AOI210     m0677(.A0(mai_mai_n705_), .A1(mai_mai_n703_), .B0(mai_mai_n500_), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n86_), .B(mai_mai_n109_), .Y(mai_mai_n707_));
  NO2        m0679(.A(mai_mai_n707_), .B(mai_mai_n57_), .Y(mai_mai_n708_));
  NO4        m0680(.A(mai_mai_n379_), .B(mai_mai_n111_), .C(j), .D(mai_mai_n214_), .Y(mai_mai_n709_));
  NA2        m0681(.A(mai_mai_n586_), .B(mai_mai_n233_), .Y(mai_mai_n710_));
  AOI220     m0682(.A0(mai_mai_n710_), .A1(mai_mai_n351_), .B0(mai_mai_n709_), .B1(mai_mai_n708_), .Y(mai_mai_n711_));
  AOI210     m0683(.A0(mai_mai_n586_), .A1(mai_mai_n155_), .B0(mai_mai_n86_), .Y(mai_mai_n712_));
  NA4        m0684(.A(mai_mai_n216_), .B(mai_mai_n139_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n713_));
  AN2        m0685(.A(l), .B(k), .Y(mai_mai_n714_));
  NA4        m0686(.A(mai_mai_n714_), .B(mai_mai_n108_), .C(mai_mai_n75_), .D(mai_mai_n214_), .Y(mai_mai_n715_));
  OAI210     m0687(.A0(mai_mai_n713_), .A1(g), .B0(mai_mai_n715_), .Y(mai_mai_n716_));
  NA2        m0688(.A(mai_mai_n716_), .B(mai_mai_n712_), .Y(mai_mai_n717_));
  NA3        m0689(.A(mai_mai_n717_), .B(mai_mai_n711_), .C(mai_mai_n706_), .Y(mai_mai_n718_));
  NO4        m0690(.A(mai_mai_n175_), .B(mai_mai_n393_), .C(mai_mai_n111_), .D(g), .Y(mai_mai_n719_));
  NA2        m0691(.A(mai_mai_n719_), .B(mai_mai_n710_), .Y(mai_mai_n720_));
  NO2        m0692(.A(mai_mai_n38_), .B(mai_mai_n213_), .Y(mai_mai_n721_));
  AOI220     m0693(.A0(mai_mai_n627_), .A1(mai_mai_n350_), .B0(mai_mai_n721_), .B1(mai_mai_n573_), .Y(mai_mai_n722_));
  NA2        m0694(.A(mai_mai_n722_), .B(mai_mai_n720_), .Y(mai_mai_n723_));
  NO2        m0695(.A(mai_mai_n545_), .B(mai_mai_n35_), .Y(mai_mai_n724_));
  INV        m0696(.A(mai_mai_n724_), .Y(mai_mai_n725_));
  NO3        m0697(.A(mai_mai_n318_), .B(mai_mai_n129_), .C(mai_mai_n41_), .Y(mai_mai_n726_));
  NA2        m0698(.A(mai_mai_n702_), .B(mai_mai_n134_), .Y(mai_mai_n727_));
  AOI220     m0699(.A0(mai_mai_n727_), .A1(mai_mai_n402_), .B0(mai_mai_n726_), .B1(mai_mai_n78_), .Y(mai_mai_n728_));
  OAI210     m0700(.A0(mai_mai_n725_), .A1(mai_mai_n89_), .B0(mai_mai_n728_), .Y(mai_mai_n729_));
  NA2        m0701(.A(mai_mai_n364_), .B(mai_mai_n43_), .Y(mai_mai_n730_));
  NA3        m0702(.A(mai_mai_n692_), .B(mai_mai_n337_), .C(mai_mai_n385_), .Y(mai_mai_n731_));
  NA2        m0703(.A(mai_mai_n714_), .B(mai_mai_n221_), .Y(mai_mai_n732_));
  NO2        m0704(.A(mai_mai_n732_), .B(mai_mai_n330_), .Y(mai_mai_n733_));
  AOI210     m0705(.A0(mai_mai_n733_), .A1(mai_mai_n683_), .B0(mai_mai_n499_), .Y(mai_mai_n734_));
  NA3        m0706(.A(m), .B(l), .C(k), .Y(mai_mai_n735_));
  AOI210     m0707(.A0(mai_mai_n665_), .A1(mai_mai_n663_), .B0(mai_mai_n735_), .Y(mai_mai_n736_));
  NO2        m0708(.A(mai_mai_n544_), .B(mai_mai_n273_), .Y(mai_mai_n737_));
  NOi21      m0709(.An(mai_mai_n737_), .B(mai_mai_n539_), .Y(mai_mai_n738_));
  NA4        m0710(.A(mai_mai_n112_), .B(l), .C(k), .D(mai_mai_n89_), .Y(mai_mai_n739_));
  NA3        m0711(.A(mai_mai_n119_), .B(mai_mai_n411_), .C(i), .Y(mai_mai_n740_));
  NO2        m0712(.A(mai_mai_n740_), .B(mai_mai_n739_), .Y(mai_mai_n741_));
  NO3        m0713(.A(mai_mai_n741_), .B(mai_mai_n738_), .C(mai_mai_n736_), .Y(mai_mai_n742_));
  NA4        m0714(.A(mai_mai_n742_), .B(mai_mai_n734_), .C(mai_mai_n731_), .D(mai_mai_n730_), .Y(mai_mai_n743_));
  NO4        m0715(.A(mai_mai_n743_), .B(mai_mai_n729_), .C(mai_mai_n723_), .D(mai_mai_n718_), .Y(mai_mai_n744_));
  NA2        m0716(.A(mai_mai_n627_), .B(mai_mai_n394_), .Y(mai_mai_n745_));
  OR2        m0717(.A(mai_mai_n599_), .B(mai_mai_n547_), .Y(mai_mai_n746_));
  NO3        m0718(.A(mai_mai_n398_), .B(mai_mai_n533_), .C(h), .Y(mai_mai_n747_));
  AOI210     m0719(.A0(mai_mai_n747_), .A1(mai_mai_n112_), .B0(mai_mai_n509_), .Y(mai_mai_n748_));
  NA4        m0720(.A(mai_mai_n748_), .B(mai_mai_n746_), .C(mai_mai_n745_), .D(mai_mai_n251_), .Y(mai_mai_n749_));
  NA2        m0721(.A(mai_mai_n714_), .B(mai_mai_n75_), .Y(mai_mai_n750_));
  NO4        m0722(.A(mai_mai_n691_), .B(mai_mai_n175_), .C(n), .D(i), .Y(mai_mai_n751_));
  NOi21      m0723(.An(h), .B(j), .Y(mai_mai_n752_));
  NA2        m0724(.A(mai_mai_n752_), .B(f), .Y(mai_mai_n753_));
  NO2        m0725(.A(mai_mai_n753_), .B(mai_mai_n248_), .Y(mai_mai_n754_));
  NO3        m0726(.A(mai_mai_n754_), .B(mai_mai_n751_), .C(mai_mai_n694_), .Y(mai_mai_n755_));
  OAI220     m0727(.A0(mai_mai_n755_), .A1(mai_mai_n750_), .B0(mai_mai_n601_), .B1(mai_mai_n62_), .Y(mai_mai_n756_));
  AOI210     m0728(.A0(mai_mai_n749_), .A1(l), .B0(mai_mai_n756_), .Y(mai_mai_n757_));
  NO2        m0729(.A(j), .B(i), .Y(mai_mai_n758_));
  NA3        m0730(.A(mai_mai_n758_), .B(mai_mai_n82_), .C(l), .Y(mai_mai_n759_));
  NA2        m0731(.A(mai_mai_n758_), .B(mai_mai_n33_), .Y(mai_mai_n760_));
  NA2        m0732(.A(mai_mai_n421_), .B(mai_mai_n119_), .Y(mai_mai_n761_));
  OR2        m0733(.A(mai_mai_n761_), .B(mai_mai_n760_), .Y(mai_mai_n762_));
  NO3        m0734(.A(mai_mai_n151_), .B(mai_mai_n49_), .C(mai_mai_n109_), .Y(mai_mai_n763_));
  NO3        m0735(.A(mai_mai_n551_), .B(mai_mai_n149_), .C(mai_mai_n75_), .Y(mai_mai_n764_));
  NO3        m0736(.A(mai_mai_n492_), .B(mai_mai_n440_), .C(j), .Y(mai_mai_n765_));
  OAI210     m0737(.A0(mai_mai_n764_), .A1(mai_mai_n763_), .B0(mai_mai_n765_), .Y(mai_mai_n766_));
  INV        m0738(.A(mai_mai_n766_), .Y(mai_mai_n767_));
  NA2        m0739(.A(k), .B(j), .Y(mai_mai_n768_));
  NO3        m0740(.A(mai_mai_n297_), .B(mai_mai_n768_), .C(mai_mai_n40_), .Y(mai_mai_n769_));
  AOI210     m0741(.A0(mai_mai_n538_), .A1(n), .B0(mai_mai_n561_), .Y(mai_mai_n770_));
  NA2        m0742(.A(mai_mai_n770_), .B(mai_mai_n564_), .Y(mai_mai_n771_));
  AN3        m0743(.A(mai_mai_n771_), .B(mai_mai_n769_), .C(mai_mai_n99_), .Y(mai_mai_n772_));
  NA2        m0744(.A(mai_mai_n618_), .B(mai_mai_n308_), .Y(mai_mai_n773_));
  INV        m0745(.A(mai_mai_n773_), .Y(mai_mai_n774_));
  NO2        m0746(.A(mai_mai_n297_), .B(mai_mai_n134_), .Y(mai_mai_n775_));
  AOI220     m0747(.A0(mai_mai_n775_), .A1(mai_mai_n627_), .B0(mai_mai_n726_), .B1(mai_mai_n712_), .Y(mai_mai_n776_));
  NO2        m0748(.A(mai_mai_n735_), .B(mai_mai_n92_), .Y(mai_mai_n777_));
  NA2        m0749(.A(mai_mai_n777_), .B(mai_mai_n597_), .Y(mai_mai_n778_));
  NO2        m0750(.A(mai_mai_n598_), .B(mai_mai_n115_), .Y(mai_mai_n779_));
  OAI210     m0751(.A0(mai_mai_n779_), .A1(mai_mai_n765_), .B0(mai_mai_n679_), .Y(mai_mai_n780_));
  NA3        m0752(.A(mai_mai_n780_), .B(mai_mai_n778_), .C(mai_mai_n776_), .Y(mai_mai_n781_));
  OR4        m0753(.A(mai_mai_n781_), .B(mai_mai_n774_), .C(mai_mai_n772_), .D(mai_mai_n767_), .Y(mai_mai_n782_));
  NA3        m0754(.A(mai_mai_n770_), .B(mai_mai_n564_), .C(mai_mai_n563_), .Y(mai_mai_n783_));
  NA4        m0755(.A(mai_mai_n783_), .B(mai_mai_n216_), .C(mai_mai_n453_), .D(mai_mai_n34_), .Y(mai_mai_n784_));
  OAI220     m0756(.A0(mai_mai_n713_), .A1(mai_mai_n704_), .B0(mai_mai_n335_), .B1(mai_mai_n38_), .Y(mai_mai_n785_));
  INV        m0757(.A(mai_mai_n785_), .Y(mai_mai_n786_));
  NA3        m0758(.A(mai_mai_n554_), .B(mai_mai_n294_), .C(h), .Y(mai_mai_n787_));
  NOi21      m0759(.An(mai_mai_n679_), .B(mai_mai_n787_), .Y(mai_mai_n788_));
  NO2        m0760(.A(mai_mai_n93_), .B(mai_mai_n47_), .Y(mai_mai_n789_));
  NO2        m0761(.A(mai_mai_n759_), .B(mai_mai_n673_), .Y(mai_mai_n790_));
  AOI210     m0762(.A0(mai_mai_n789_), .A1(mai_mai_n645_), .B0(mai_mai_n790_), .Y(mai_mai_n791_));
  NAi41      m0763(.An(mai_mai_n788_), .B(mai_mai_n791_), .C(mai_mai_n786_), .D(mai_mai_n784_), .Y(mai_mai_n792_));
  OR2        m0764(.A(mai_mai_n777_), .B(mai_mai_n96_), .Y(mai_mai_n793_));
  AOI220     m0765(.A0(mai_mai_n793_), .A1(mai_mai_n239_), .B0(mai_mai_n765_), .B1(mai_mai_n639_), .Y(mai_mai_n794_));
  INV        m0766(.A(mai_mai_n339_), .Y(mai_mai_n795_));
  OAI210     m0767(.A0(mai_mai_n735_), .A1(mai_mai_n662_), .B0(mai_mai_n528_), .Y(mai_mai_n796_));
  NA3        m0768(.A(mai_mai_n250_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n797_));
  AOI220     m0769(.A0(mai_mai_n612_), .A1(mai_mai_n29_), .B0(mai_mai_n469_), .B1(mai_mai_n86_), .Y(mai_mai_n798_));
  NA2        m0770(.A(mai_mai_n798_), .B(mai_mai_n797_), .Y(mai_mai_n799_));
  NO2        m0771(.A(mai_mai_n787_), .B(mai_mai_n498_), .Y(mai_mai_n800_));
  AOI210     m0772(.A0(mai_mai_n799_), .A1(mai_mai_n796_), .B0(mai_mai_n800_), .Y(mai_mai_n801_));
  NA3        m0773(.A(mai_mai_n801_), .B(mai_mai_n795_), .C(mai_mai_n794_), .Y(mai_mai_n802_));
  NOi41      m0774(.An(mai_mai_n762_), .B(mai_mai_n802_), .C(mai_mai_n792_), .D(mai_mai_n782_), .Y(mai_mai_n803_));
  OR3        m0775(.A(mai_mai_n713_), .B(mai_mai_n233_), .C(g), .Y(mai_mai_n804_));
  NO3        m0776(.A(mai_mai_n345_), .B(mai_mai_n299_), .C(mai_mai_n111_), .Y(mai_mai_n805_));
  NA2        m0777(.A(mai_mai_n805_), .B(mai_mai_n771_), .Y(mai_mai_n806_));
  NA2        m0778(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n807_));
  NO3        m0779(.A(mai_mai_n807_), .B(mai_mai_n760_), .C(mai_mai_n278_), .Y(mai_mai_n808_));
  NO3        m0780(.A(mai_mai_n533_), .B(mai_mai_n94_), .C(h), .Y(mai_mai_n809_));
  AOI210     m0781(.A0(mai_mai_n809_), .A1(mai_mai_n708_), .B0(mai_mai_n808_), .Y(mai_mai_n810_));
  NA4        m0782(.A(mai_mai_n810_), .B(mai_mai_n806_), .C(mai_mai_n804_), .D(mai_mai_n404_), .Y(mai_mai_n811_));
  OR2        m0783(.A(mai_mai_n662_), .B(mai_mai_n93_), .Y(mai_mai_n812_));
  NOi31      m0784(.An(b), .B(d), .C(a), .Y(mai_mai_n813_));
  NO2        m0785(.A(mai_mai_n813_), .B(mai_mai_n610_), .Y(mai_mai_n814_));
  NO2        m0786(.A(mai_mai_n814_), .B(n), .Y(mai_mai_n815_));
  NOi21      m0787(.An(mai_mai_n798_), .B(mai_mai_n815_), .Y(mai_mai_n816_));
  OAI220     m0788(.A0(mai_mai_n816_), .A1(mai_mai_n812_), .B0(mai_mai_n787_), .B1(mai_mai_n611_), .Y(mai_mai_n817_));
  NO2        m0789(.A(mai_mai_n562_), .B(mai_mai_n86_), .Y(mai_mai_n818_));
  NO3        m0790(.A(mai_mai_n626_), .B(mai_mai_n330_), .C(mai_mai_n115_), .Y(mai_mai_n819_));
  NOi21      m0791(.An(mai_mai_n819_), .B(mai_mai_n160_), .Y(mai_mai_n820_));
  AOI210     m0792(.A0(mai_mai_n805_), .A1(mai_mai_n818_), .B0(mai_mai_n820_), .Y(mai_mai_n821_));
  OAI210     m0793(.A0(mai_mai_n713_), .A1(mai_mai_n395_), .B0(mai_mai_n821_), .Y(mai_mai_n822_));
  NO2        m0794(.A(mai_mai_n691_), .B(n), .Y(mai_mai_n823_));
  AOI220     m0795(.A0(mai_mai_n775_), .A1(mai_mai_n669_), .B0(mai_mai_n823_), .B1(mai_mai_n703_), .Y(mai_mai_n824_));
  NO2        m0796(.A(mai_mai_n325_), .B(mai_mai_n238_), .Y(mai_mai_n825_));
  NA2        m0797(.A(mai_mai_n119_), .B(mai_mai_n86_), .Y(mai_mai_n826_));
  AOI210     m0798(.A0(mai_mai_n425_), .A1(mai_mai_n417_), .B0(mai_mai_n826_), .Y(mai_mai_n827_));
  NA2        m0799(.A(mai_mai_n733_), .B(mai_mai_n34_), .Y(mai_mai_n828_));
  NAi21      m0800(.An(mai_mai_n739_), .B(mai_mai_n436_), .Y(mai_mai_n829_));
  NO2        m0801(.A(mai_mai_n273_), .B(i), .Y(mai_mai_n830_));
  NAi41      m0802(.An(mai_mai_n827_), .B(mai_mai_n829_), .C(mai_mai_n828_), .D(mai_mai_n824_), .Y(mai_mai_n831_));
  NO4        m0803(.A(mai_mai_n831_), .B(mai_mai_n822_), .C(mai_mai_n817_), .D(mai_mai_n811_), .Y(mai_mai_n832_));
  NA4        m0804(.A(mai_mai_n832_), .B(mai_mai_n803_), .C(mai_mai_n757_), .D(mai_mai_n744_), .Y(mai09));
  INV        m0805(.A(mai_mai_n120_), .Y(mai_mai_n834_));
  NA2        m0806(.A(f), .B(e), .Y(mai_mai_n835_));
  NO2        m0807(.A(mai_mai_n226_), .B(mai_mai_n111_), .Y(mai_mai_n836_));
  NA2        m0808(.A(mai_mai_n836_), .B(g), .Y(mai_mai_n837_));
  NA4        m0809(.A(mai_mai_n311_), .B(mai_mai_n478_), .C(mai_mai_n261_), .D(mai_mai_n117_), .Y(mai_mai_n838_));
  AOI210     m0810(.A0(mai_mai_n838_), .A1(g), .B0(mai_mai_n475_), .Y(mai_mai_n839_));
  AOI210     m0811(.A0(mai_mai_n839_), .A1(mai_mai_n837_), .B0(mai_mai_n835_), .Y(mai_mai_n840_));
  NA2        m0812(.A(mai_mai_n446_), .B(e), .Y(mai_mai_n841_));
  NO2        m0813(.A(mai_mai_n841_), .B(mai_mai_n519_), .Y(mai_mai_n842_));
  AOI210     m0814(.A0(mai_mai_n840_), .A1(mai_mai_n834_), .B0(mai_mai_n842_), .Y(mai_mai_n843_));
  NO2        m0815(.A(mai_mai_n207_), .B(mai_mai_n213_), .Y(mai_mai_n844_));
  NA3        m0816(.A(m), .B(l), .C(i), .Y(mai_mai_n845_));
  OAI220     m0817(.A0(mai_mai_n598_), .A1(mai_mai_n845_), .B0(mai_mai_n355_), .B1(mai_mai_n534_), .Y(mai_mai_n846_));
  NA4        m0818(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(g), .D(f), .Y(mai_mai_n847_));
  NAi31      m0819(.An(mai_mai_n846_), .B(mai_mai_n847_), .C(mai_mai_n441_), .Y(mai_mai_n848_));
  OR2        m0820(.A(mai_mai_n848_), .B(mai_mai_n844_), .Y(mai_mai_n849_));
  NA3        m0821(.A(mai_mai_n812_), .B(mai_mai_n575_), .C(mai_mai_n528_), .Y(mai_mai_n850_));
  OA210      m0822(.A0(mai_mai_n850_), .A1(mai_mai_n849_), .B0(mai_mai_n815_), .Y(mai_mai_n851_));
  INV        m0823(.A(mai_mai_n342_), .Y(mai_mai_n852_));
  NO2        m0824(.A(mai_mai_n125_), .B(mai_mai_n124_), .Y(mai_mai_n853_));
  NOi31      m0825(.An(k), .B(m), .C(l), .Y(mai_mai_n854_));
  NO2        m0826(.A(mai_mai_n344_), .B(mai_mai_n854_), .Y(mai_mai_n855_));
  AOI210     m0827(.A0(mai_mai_n855_), .A1(mai_mai_n853_), .B0(mai_mai_n605_), .Y(mai_mai_n856_));
  NA2        m0828(.A(mai_mai_n797_), .B(mai_mai_n335_), .Y(mai_mai_n857_));
  NA2        m0829(.A(mai_mai_n346_), .B(mai_mai_n348_), .Y(mai_mai_n858_));
  OAI210     m0830(.A0(mai_mai_n207_), .A1(mai_mai_n213_), .B0(mai_mai_n858_), .Y(mai_mai_n859_));
  AOI220     m0831(.A0(mai_mai_n859_), .A1(mai_mai_n857_), .B0(mai_mai_n856_), .B1(mai_mai_n852_), .Y(mai_mai_n860_));
  NA2        m0832(.A(mai_mai_n169_), .B(mai_mai_n113_), .Y(mai_mai_n861_));
  NA3        m0833(.A(mai_mai_n861_), .B(mai_mai_n702_), .C(mai_mai_n134_), .Y(mai_mai_n862_));
  NA3        m0834(.A(mai_mai_n862_), .B(mai_mai_n192_), .C(mai_mai_n31_), .Y(mai_mai_n863_));
  NA4        m0835(.A(mai_mai_n863_), .B(mai_mai_n860_), .C(mai_mai_n628_), .D(mai_mai_n84_), .Y(mai_mai_n864_));
  NO2        m0836(.A(mai_mai_n595_), .B(mai_mai_n506_), .Y(mai_mai_n865_));
  NA2        m0837(.A(mai_mai_n865_), .B(mai_mai_n192_), .Y(mai_mai_n866_));
  NOi21      m0838(.An(f), .B(d), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n867_), .B(m), .Y(mai_mai_n868_));
  NO2        m0840(.A(mai_mai_n868_), .B(mai_mai_n52_), .Y(mai_mai_n869_));
  NOi32      m0841(.An(g), .Bn(f), .C(d), .Y(mai_mai_n870_));
  NA4        m0842(.A(mai_mai_n870_), .B(mai_mai_n612_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n871_));
  NA2        m0843(.A(mai_mai_n869_), .B(mai_mai_n552_), .Y(mai_mai_n872_));
  NA3        m0844(.A(mai_mai_n311_), .B(mai_mai_n261_), .C(mai_mai_n117_), .Y(mai_mai_n873_));
  AN2        m0845(.A(f), .B(d), .Y(mai_mai_n874_));
  NA3        m0846(.A(mai_mai_n483_), .B(mai_mai_n874_), .C(mai_mai_n86_), .Y(mai_mai_n875_));
  NO3        m0847(.A(mai_mai_n875_), .B(mai_mai_n75_), .C(mai_mai_n214_), .Y(mai_mai_n876_));
  NO2        m0848(.A(mai_mai_n287_), .B(mai_mai_n56_), .Y(mai_mai_n877_));
  NA2        m0849(.A(mai_mai_n873_), .B(mai_mai_n876_), .Y(mai_mai_n878_));
  NAi41      m0850(.An(mai_mai_n497_), .B(mai_mai_n878_), .C(mai_mai_n872_), .D(mai_mai_n866_), .Y(mai_mai_n879_));
  NO4        m0851(.A(mai_mai_n626_), .B(mai_mai_n130_), .C(mai_mai_n330_), .D(mai_mai_n152_), .Y(mai_mai_n880_));
  NO2        m0852(.A(mai_mai_n656_), .B(mai_mai_n330_), .Y(mai_mai_n881_));
  AN2        m0853(.A(mai_mai_n881_), .B(mai_mai_n683_), .Y(mai_mai_n882_));
  NO3        m0854(.A(mai_mai_n882_), .B(mai_mai_n880_), .C(mai_mai_n235_), .Y(mai_mai_n883_));
  NA2        m0855(.A(mai_mai_n610_), .B(mai_mai_n86_), .Y(mai_mai_n884_));
  NO2        m0856(.A(mai_mai_n858_), .B(mai_mai_n884_), .Y(mai_mai_n885_));
  NA3        m0857(.A(mai_mai_n159_), .B(mai_mai_n108_), .C(mai_mai_n107_), .Y(mai_mai_n886_));
  OAI220     m0858(.A0(mai_mai_n875_), .A1(mai_mai_n430_), .B0(mai_mai_n342_), .B1(mai_mai_n886_), .Y(mai_mai_n887_));
  NOi41      m0859(.An(mai_mai_n224_), .B(mai_mai_n887_), .C(mai_mai_n885_), .D(mai_mai_n306_), .Y(mai_mai_n888_));
  NA2        m0860(.A(c), .B(mai_mai_n114_), .Y(mai_mai_n889_));
  NO2        m0861(.A(mai_mai_n889_), .B(mai_mai_n408_), .Y(mai_mai_n890_));
  NA3        m0862(.A(mai_mai_n890_), .B(mai_mai_n517_), .C(f), .Y(mai_mai_n891_));
  OR2        m0863(.A(mai_mai_n662_), .B(mai_mai_n548_), .Y(mai_mai_n892_));
  INV        m0864(.A(mai_mai_n892_), .Y(mai_mai_n893_));
  NA2        m0865(.A(mai_mai_n814_), .B(mai_mai_n110_), .Y(mai_mai_n894_));
  NA2        m0866(.A(mai_mai_n894_), .B(mai_mai_n893_), .Y(mai_mai_n895_));
  NA4        m0867(.A(mai_mai_n895_), .B(mai_mai_n891_), .C(mai_mai_n888_), .D(mai_mai_n883_), .Y(mai_mai_n896_));
  NO4        m0868(.A(mai_mai_n896_), .B(mai_mai_n879_), .C(mai_mai_n864_), .D(mai_mai_n851_), .Y(mai_mai_n897_));
  OR2        m0869(.A(mai_mai_n875_), .B(mai_mai_n75_), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n111_), .B(j), .Y(mai_mai_n899_));
  NA2        m0871(.A(mai_mai_n836_), .B(g), .Y(mai_mai_n900_));
  AOI210     m0872(.A0(mai_mai_n900_), .A1(mai_mai_n295_), .B0(mai_mai_n898_), .Y(mai_mai_n901_));
  NO2        m0873(.A(mai_mai_n134_), .B(mai_mai_n130_), .Y(mai_mai_n902_));
  NO2        m0874(.A(mai_mai_n231_), .B(mai_mai_n225_), .Y(mai_mai_n903_));
  AOI220     m0875(.A0(mai_mai_n903_), .A1(mai_mai_n228_), .B0(mai_mai_n304_), .B1(mai_mai_n902_), .Y(mai_mai_n904_));
  NO2        m0876(.A(mai_mai_n430_), .B(mai_mai_n835_), .Y(mai_mai_n905_));
  NA2        m0877(.A(mai_mai_n905_), .B(mai_mai_n569_), .Y(mai_mai_n906_));
  NA2        m0878(.A(mai_mai_n906_), .B(mai_mai_n904_), .Y(mai_mai_n907_));
  NA2        m0879(.A(e), .B(d), .Y(mai_mai_n908_));
  OAI220     m0880(.A0(mai_mai_n908_), .A1(c), .B0(mai_mai_n325_), .B1(d), .Y(mai_mai_n909_));
  NA3        m0881(.A(mai_mai_n909_), .B(mai_mai_n458_), .C(mai_mai_n515_), .Y(mai_mai_n910_));
  AOI210     m0882(.A0(mai_mai_n523_), .A1(mai_mai_n182_), .B0(mai_mai_n231_), .Y(mai_mai_n911_));
  AOI210     m0883(.A0(mai_mai_n627_), .A1(mai_mai_n350_), .B0(mai_mai_n911_), .Y(mai_mai_n912_));
  NA2        m0884(.A(mai_mai_n287_), .B(mai_mai_n165_), .Y(mai_mai_n913_));
  NA2        m0885(.A(mai_mai_n876_), .B(mai_mai_n913_), .Y(mai_mai_n914_));
  NA3        m0886(.A(mai_mai_n168_), .B(mai_mai_n87_), .C(mai_mai_n34_), .Y(mai_mai_n915_));
  NA4        m0887(.A(mai_mai_n915_), .B(mai_mai_n914_), .C(mai_mai_n912_), .D(mai_mai_n910_), .Y(mai_mai_n916_));
  NO3        m0888(.A(mai_mai_n916_), .B(mai_mai_n907_), .C(mai_mai_n901_), .Y(mai_mai_n917_));
  NA2        m0889(.A(mai_mai_n852_), .B(mai_mai_n31_), .Y(mai_mai_n918_));
  AO210      m0890(.A0(mai_mai_n918_), .A1(mai_mai_n704_), .B0(mai_mai_n217_), .Y(mai_mai_n919_));
  OAI220     m0891(.A0(mai_mai_n626_), .A1(mai_mai_n61_), .B0(mai_mai_n299_), .B1(j), .Y(mai_mai_n920_));
  AOI220     m0892(.A0(mai_mai_n920_), .A1(mai_mai_n881_), .B0(mai_mai_n616_), .B1(mai_mai_n625_), .Y(mai_mai_n921_));
  OAI210     m0893(.A0(mai_mai_n841_), .A1(mai_mai_n172_), .B0(mai_mai_n921_), .Y(mai_mai_n922_));
  AOI210     m0894(.A0(mai_mai_n116_), .A1(mai_mai_n115_), .B0(mai_mai_n260_), .Y(mai_mai_n923_));
  NO2        m0895(.A(mai_mai_n923_), .B(mai_mai_n871_), .Y(mai_mai_n924_));
  AO210      m0896(.A0(mai_mai_n857_), .A1(mai_mai_n846_), .B0(mai_mai_n924_), .Y(mai_mai_n925_));
  NO2        m0897(.A(mai_mai_n925_), .B(mai_mai_n922_), .Y(mai_mai_n926_));
  AO220      m0898(.A0(mai_mai_n458_), .A1(mai_mai_n752_), .B0(mai_mai_n177_), .B1(f), .Y(mai_mai_n927_));
  OAI210     m0899(.A0(mai_mai_n927_), .A1(mai_mai_n461_), .B0(mai_mai_n909_), .Y(mai_mai_n928_));
  NA2        m0900(.A(mai_mai_n850_), .B(mai_mai_n708_), .Y(mai_mai_n929_));
  AN4        m0901(.A(mai_mai_n929_), .B(mai_mai_n928_), .C(mai_mai_n926_), .D(mai_mai_n919_), .Y(mai_mai_n930_));
  NA4        m0902(.A(mai_mai_n930_), .B(mai_mai_n917_), .C(mai_mai_n897_), .D(mai_mai_n843_), .Y(mai12));
  NO2        m0903(.A(mai_mai_n456_), .B(c), .Y(mai_mai_n932_));
  NO4        m0904(.A(mai_mai_n445_), .B(mai_mai_n252_), .C(mai_mai_n591_), .D(mai_mai_n214_), .Y(mai_mai_n933_));
  NA2        m0905(.A(mai_mai_n933_), .B(mai_mai_n932_), .Y(mai_mai_n934_));
  NO2        m0906(.A(mai_mai_n456_), .B(mai_mai_n114_), .Y(mai_mai_n935_));
  NO2        m0907(.A(mai_mai_n853_), .B(mai_mai_n355_), .Y(mai_mai_n936_));
  NO2        m0908(.A(mai_mai_n662_), .B(mai_mai_n379_), .Y(mai_mai_n937_));
  AOI220     m0909(.A0(mai_mai_n937_), .A1(mai_mai_n550_), .B0(mai_mai_n936_), .B1(mai_mai_n935_), .Y(mai_mai_n938_));
  NA3        m0910(.A(mai_mai_n938_), .B(mai_mai_n934_), .C(mai_mai_n444_), .Y(mai_mai_n939_));
  AOI210     m0911(.A0(mai_mai_n234_), .A1(mai_mai_n341_), .B0(mai_mai_n204_), .Y(mai_mai_n940_));
  OR2        m0912(.A(mai_mai_n940_), .B(mai_mai_n933_), .Y(mai_mai_n941_));
  AOI210     m0913(.A0(mai_mai_n338_), .A1(mai_mai_n391_), .B0(mai_mai_n214_), .Y(mai_mai_n942_));
  OAI210     m0914(.A0(mai_mai_n942_), .A1(mai_mai_n941_), .B0(mai_mai_n403_), .Y(mai_mai_n943_));
  NO2        m0915(.A(mai_mai_n642_), .B(mai_mai_n263_), .Y(mai_mai_n944_));
  NO2        m0916(.A(mai_mai_n598_), .B(mai_mai_n845_), .Y(mai_mai_n945_));
  AOI220     m0917(.A0(mai_mai_n945_), .A1(mai_mai_n573_), .B0(mai_mai_n825_), .B1(mai_mai_n944_), .Y(mai_mai_n946_));
  NO2        m0918(.A(mai_mai_n151_), .B(mai_mai_n238_), .Y(mai_mai_n947_));
  NA2        m0919(.A(mai_mai_n946_), .B(mai_mai_n943_), .Y(mai_mai_n948_));
  OR2        m0920(.A(mai_mai_n326_), .B(mai_mai_n935_), .Y(mai_mai_n949_));
  NA2        m0921(.A(mai_mai_n949_), .B(mai_mai_n356_), .Y(mai_mai_n950_));
  NO3        m0922(.A(mai_mai_n130_), .B(mai_mai_n152_), .C(mai_mai_n214_), .Y(mai_mai_n951_));
  NA2        m0923(.A(mai_mai_n951_), .B(mai_mai_n538_), .Y(mai_mai_n952_));
  NA4        m0924(.A(mai_mai_n446_), .B(mai_mai_n438_), .C(mai_mai_n183_), .D(g), .Y(mai_mai_n953_));
  NA3        m0925(.A(mai_mai_n953_), .B(mai_mai_n952_), .C(mai_mai_n950_), .Y(mai_mai_n954_));
  NO3        m0926(.A(mai_mai_n667_), .B(mai_mai_n93_), .C(mai_mai_n45_), .Y(mai_mai_n955_));
  NO4        m0927(.A(mai_mai_n955_), .B(mai_mai_n954_), .C(mai_mai_n948_), .D(mai_mai_n939_), .Y(mai_mai_n956_));
  NO2        m0928(.A(mai_mai_n371_), .B(mai_mai_n370_), .Y(mai_mai_n957_));
  NA2        m0929(.A(mai_mai_n596_), .B(mai_mai_n73_), .Y(mai_mai_n958_));
  NA2        m0930(.A(mai_mai_n562_), .B(mai_mai_n144_), .Y(mai_mai_n959_));
  NOi21      m0931(.An(mai_mai_n34_), .B(mai_mai_n656_), .Y(mai_mai_n960_));
  AOI220     m0932(.A0(mai_mai_n960_), .A1(mai_mai_n959_), .B0(mai_mai_n958_), .B1(mai_mai_n957_), .Y(mai_mai_n961_));
  OAI210     m0933(.A0(mai_mai_n251_), .A1(mai_mai_n45_), .B0(mai_mai_n961_), .Y(mai_mai_n962_));
  NA2        m0934(.A(mai_mai_n436_), .B(mai_mai_n265_), .Y(mai_mai_n963_));
  NO3        m0935(.A(mai_mai_n826_), .B(mai_mai_n91_), .C(mai_mai_n408_), .Y(mai_mai_n964_));
  NAi31      m0936(.An(mai_mai_n964_), .B(mai_mai_n963_), .C(mai_mai_n322_), .Y(mai_mai_n965_));
  NO2        m0937(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n966_));
  NO2        m0938(.A(mai_mai_n512_), .B(mai_mai_n299_), .Y(mai_mai_n967_));
  INV        m0939(.A(mai_mai_n967_), .Y(mai_mai_n968_));
  NO2        m0940(.A(mai_mai_n968_), .B(mai_mai_n144_), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n635_), .B(mai_mai_n365_), .Y(mai_mai_n970_));
  OAI210     m0942(.A0(mai_mai_n740_), .A1(mai_mai_n970_), .B0(mai_mai_n369_), .Y(mai_mai_n971_));
  NO4        m0943(.A(mai_mai_n971_), .B(mai_mai_n969_), .C(mai_mai_n965_), .D(mai_mai_n962_), .Y(mai_mai_n972_));
  NA2        m0944(.A(mai_mai_n350_), .B(g), .Y(mai_mai_n973_));
  NA2        m0945(.A(mai_mai_n162_), .B(i), .Y(mai_mai_n974_));
  NA2        m0946(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n975_));
  OAI220     m0947(.A0(mai_mai_n975_), .A1(mai_mai_n203_), .B0(mai_mai_n974_), .B1(mai_mai_n93_), .Y(mai_mai_n976_));
  AOI210     m0948(.A0(mai_mai_n419_), .A1(mai_mai_n37_), .B0(mai_mai_n976_), .Y(mai_mai_n977_));
  NO2        m0949(.A(mai_mai_n144_), .B(mai_mai_n86_), .Y(mai_mai_n978_));
  OR2        m0950(.A(mai_mai_n978_), .B(mai_mai_n561_), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n562_), .B(mai_mai_n383_), .Y(mai_mai_n980_));
  AOI210     m0952(.A0(mai_mai_n980_), .A1(n), .B0(mai_mai_n979_), .Y(mai_mai_n981_));
  OAI220     m0953(.A0(mai_mai_n981_), .A1(mai_mai_n973_), .B0(mai_mai_n977_), .B1(mai_mai_n335_), .Y(mai_mai_n982_));
  NO2        m0954(.A(mai_mai_n662_), .B(mai_mai_n506_), .Y(mai_mai_n983_));
  NA3        m0955(.A(mai_mai_n346_), .B(mai_mai_n632_), .C(i), .Y(mai_mai_n984_));
  OAI210     m0956(.A0(mai_mai_n440_), .A1(mai_mai_n311_), .B0(mai_mai_n984_), .Y(mai_mai_n985_));
  OAI210     m0957(.A0(mai_mai_n985_), .A1(mai_mai_n983_), .B0(mai_mai_n679_), .Y(mai_mai_n986_));
  OR3        m0958(.A(mai_mai_n311_), .B(mai_mai_n435_), .C(f), .Y(mai_mai_n987_));
  NA3        m0959(.A(mai_mai_n327_), .B(mai_mai_n116_), .C(g), .Y(mai_mai_n988_));
  AOI210     m0960(.A0(mai_mai_n676_), .A1(mai_mai_n988_), .B0(m), .Y(mai_mai_n989_));
  OAI210     m0961(.A0(mai_mai_n989_), .A1(mai_mai_n936_), .B0(mai_mai_n326_), .Y(mai_mai_n990_));
  NA2        m0962(.A(mai_mai_n695_), .B(mai_mai_n884_), .Y(mai_mai_n991_));
  NA2        m0963(.A(mai_mai_n847_), .B(mai_mai_n441_), .Y(mai_mai_n992_));
  INV        m0964(.A(mai_mai_n987_), .Y(mai_mai_n993_));
  AOI220     m0965(.A0(mai_mai_n993_), .A1(mai_mai_n258_), .B0(mai_mai_n992_), .B1(mai_mai_n991_), .Y(mai_mai_n994_));
  NA3        m0966(.A(mai_mai_n994_), .B(mai_mai_n990_), .C(mai_mai_n986_), .Y(mai_mai_n995_));
  NO2        m0967(.A(mai_mai_n379_), .B(mai_mai_n92_), .Y(mai_mai_n996_));
  OAI210     m0968(.A0(mai_mai_n996_), .A1(mai_mai_n944_), .B0(mai_mai_n239_), .Y(mai_mai_n997_));
  NA2        m0969(.A(mai_mai_n666_), .B(mai_mai_n90_), .Y(mai_mai_n998_));
  NO2        m0970(.A(mai_mai_n464_), .B(mai_mai_n214_), .Y(mai_mai_n999_));
  AOI220     m0971(.A0(mai_mai_n999_), .A1(mai_mai_n384_), .B0(mai_mai_n949_), .B1(mai_mai_n218_), .Y(mai_mai_n1000_));
  NA2        m0972(.A(mai_mai_n937_), .B(mai_mai_n947_), .Y(mai_mai_n1001_));
  NA4        m0973(.A(mai_mai_n1001_), .B(mai_mai_n1000_), .C(mai_mai_n998_), .D(mai_mai_n997_), .Y(mai_mai_n1002_));
  OAI210     m0974(.A0(mai_mai_n992_), .A1(mai_mai_n945_), .B0(mai_mai_n550_), .Y(mai_mai_n1003_));
  AOI210     m0975(.A0(mai_mai_n420_), .A1(mai_mai_n412_), .B0(mai_mai_n826_), .Y(mai_mai_n1004_));
  INV        m0976(.A(mai_mai_n1004_), .Y(mai_mai_n1005_));
  NA2        m0977(.A(mai_mai_n989_), .B(mai_mai_n935_), .Y(mai_mai_n1006_));
  NO3        m0978(.A(mai_mai_n899_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n1007_));
  AOI220     m0979(.A0(mai_mai_n1007_), .A1(mai_mai_n630_), .B0(mai_mai_n647_), .B1(mai_mai_n538_), .Y(mai_mai_n1008_));
  NA4        m0980(.A(mai_mai_n1008_), .B(mai_mai_n1006_), .C(mai_mai_n1005_), .D(mai_mai_n1003_), .Y(mai_mai_n1009_));
  NO4        m0981(.A(mai_mai_n1009_), .B(mai_mai_n1002_), .C(mai_mai_n995_), .D(mai_mai_n982_), .Y(mai_mai_n1010_));
  NAi31      m0982(.An(mai_mai_n140_), .B(mai_mai_n421_), .C(n), .Y(mai_mai_n1011_));
  NO3        m0983(.A(mai_mai_n124_), .B(mai_mai_n344_), .C(mai_mai_n854_), .Y(mai_mai_n1012_));
  NO2        m0984(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .Y(mai_mai_n1013_));
  NO3        m0985(.A(mai_mai_n273_), .B(mai_mai_n140_), .C(mai_mai_n408_), .Y(mai_mai_n1014_));
  AOI210     m0986(.A0(mai_mai_n1014_), .A1(mai_mai_n507_), .B0(mai_mai_n1013_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(mai_mai_n500_), .B(i), .Y(mai_mai_n1016_));
  NA2        m0988(.A(mai_mai_n1016_), .B(mai_mai_n1015_), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n231_), .B(mai_mai_n173_), .Y(mai_mai_n1018_));
  NO3        m0990(.A(mai_mai_n308_), .B(mai_mai_n446_), .C(mai_mai_n177_), .Y(mai_mai_n1019_));
  NOi31      m0991(.An(mai_mai_n1018_), .B(mai_mai_n1019_), .C(mai_mai_n214_), .Y(mai_mai_n1020_));
  NAi21      m0992(.An(mai_mai_n562_), .B(mai_mai_n999_), .Y(mai_mai_n1021_));
  NA2        m0993(.A(mai_mai_n439_), .B(mai_mai_n884_), .Y(mai_mai_n1022_));
  NO3        m0994(.A(mai_mai_n440_), .B(mai_mai_n311_), .C(mai_mai_n75_), .Y(mai_mai_n1023_));
  AOI220     m0995(.A0(mai_mai_n1023_), .A1(mai_mai_n1022_), .B0(mai_mai_n489_), .B1(g), .Y(mai_mai_n1024_));
  NA2        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1021_), .Y(mai_mai_n1025_));
  OAI220     m0997(.A0(mai_mai_n1011_), .A1(mai_mai_n234_), .B0(mai_mai_n984_), .B1(mai_mai_n611_), .Y(mai_mai_n1026_));
  NO2        m0998(.A(mai_mai_n663_), .B(mai_mai_n379_), .Y(mai_mai_n1027_));
  NA2        m0999(.A(mai_mai_n940_), .B(mai_mai_n932_), .Y(mai_mai_n1028_));
  NO3        m1000(.A(mai_mai_n551_), .B(mai_mai_n149_), .C(mai_mai_n213_), .Y(mai_mai_n1029_));
  OAI210     m1001(.A0(mai_mai_n1029_), .A1(mai_mai_n532_), .B0(mai_mai_n380_), .Y(mai_mai_n1030_));
  OAI220     m1002(.A0(mai_mai_n937_), .A1(mai_mai_n945_), .B0(mai_mai_n552_), .B1(mai_mai_n429_), .Y(mai_mai_n1031_));
  NA4        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1030_), .C(mai_mai_n1028_), .D(mai_mai_n624_), .Y(mai_mai_n1032_));
  OAI210     m1004(.A0(mai_mai_n940_), .A1(mai_mai_n933_), .B0(mai_mai_n1018_), .Y(mai_mai_n1033_));
  NA3        m1005(.A(mai_mai_n980_), .B(mai_mai_n494_), .C(mai_mai_n46_), .Y(mai_mai_n1034_));
  INV        m1006(.A(mai_mai_n334_), .Y(mai_mai_n1035_));
  NA4        m1007(.A(mai_mai_n1035_), .B(mai_mai_n1034_), .C(mai_mai_n1033_), .D(mai_mai_n274_), .Y(mai_mai_n1036_));
  OR4        m1008(.A(mai_mai_n1036_), .B(mai_mai_n1032_), .C(mai_mai_n1027_), .D(mai_mai_n1026_), .Y(mai_mai_n1037_));
  NO4        m1009(.A(mai_mai_n1037_), .B(mai_mai_n1025_), .C(mai_mai_n1020_), .D(mai_mai_n1017_), .Y(mai_mai_n1038_));
  NA4        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1010_), .C(mai_mai_n972_), .D(mai_mai_n956_), .Y(mai13));
  NA2        m1011(.A(mai_mai_n46_), .B(mai_mai_n89_), .Y(mai_mai_n1040_));
  AN2        m1012(.A(c), .B(b), .Y(mai_mai_n1041_));
  NA3        m1013(.A(mai_mai_n250_), .B(mai_mai_n1041_), .C(m), .Y(mai_mai_n1042_));
  NA2        m1014(.A(mai_mai_n505_), .B(f), .Y(mai_mai_n1043_));
  NO4        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1042_), .C(mai_mai_n1040_), .D(mai_mai_n592_), .Y(mai_mai_n1044_));
  NA2        m1016(.A(mai_mai_n265_), .B(mai_mai_n1041_), .Y(mai_mai_n1045_));
  NO4        m1017(.A(mai_mai_n1045_), .B(mai_mai_n1043_), .C(mai_mai_n974_), .D(a), .Y(mai_mai_n1046_));
  NAi32      m1018(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1047_));
  NA2        m1019(.A(mai_mai_n139_), .B(mai_mai_n45_), .Y(mai_mai_n1048_));
  NO4        m1020(.A(mai_mai_n1048_), .B(mai_mai_n1047_), .C(mai_mai_n598_), .D(mai_mai_n307_), .Y(mai_mai_n1049_));
  NA2        m1021(.A(mai_mai_n670_), .B(mai_mai_n225_), .Y(mai_mai_n1050_));
  NA2        m1022(.A(mai_mai_n411_), .B(mai_mai_n213_), .Y(mai_mai_n1051_));
  AN2        m1023(.A(d), .B(c), .Y(mai_mai_n1052_));
  NA2        m1024(.A(mai_mai_n1052_), .B(mai_mai_n114_), .Y(mai_mai_n1053_));
  NO4        m1025(.A(mai_mai_n1053_), .B(mai_mai_n1051_), .C(mai_mai_n178_), .D(mai_mai_n169_), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n505_), .B(c), .Y(mai_mai_n1055_));
  NO4        m1027(.A(mai_mai_n1048_), .B(mai_mai_n595_), .C(mai_mai_n1055_), .D(mai_mai_n307_), .Y(mai_mai_n1056_));
  AO210      m1028(.A0(mai_mai_n1054_), .A1(mai_mai_n1050_), .B0(mai_mai_n1056_), .Y(mai_mai_n1057_));
  OR4        m1029(.A(mai_mai_n1057_), .B(mai_mai_n1049_), .C(mai_mai_n1046_), .D(mai_mai_n1044_), .Y(mai_mai_n1058_));
  NAi32      m1030(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1059_));
  NO2        m1031(.A(mai_mai_n1059_), .B(mai_mai_n146_), .Y(mai_mai_n1060_));
  NA2        m1032(.A(mai_mai_n1060_), .B(g), .Y(mai_mai_n1061_));
  OR3        m1033(.A(mai_mai_n225_), .B(mai_mai_n178_), .C(mai_mai_n169_), .Y(mai_mai_n1062_));
  NO2        m1034(.A(mai_mai_n1062_), .B(mai_mai_n1061_), .Y(mai_mai_n1063_));
  NO2        m1035(.A(mai_mai_n1055_), .B(mai_mai_n307_), .Y(mai_mai_n1064_));
  NO2        m1036(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1065_));
  NA2        m1037(.A(mai_mai_n634_), .B(mai_mai_n1065_), .Y(mai_mai_n1066_));
  NOi21      m1038(.An(mai_mai_n1064_), .B(mai_mai_n1066_), .Y(mai_mai_n1067_));
  NO2        m1039(.A(mai_mai_n768_), .B(mai_mai_n111_), .Y(mai_mai_n1068_));
  NOi41      m1040(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1069_));
  NA2        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1068_), .Y(mai_mai_n1070_));
  NO2        m1042(.A(mai_mai_n1070_), .B(mai_mai_n1061_), .Y(mai_mai_n1071_));
  OR3        m1043(.A(e), .B(d), .C(c), .Y(mai_mai_n1072_));
  NA3        m1044(.A(k), .B(j), .C(i), .Y(mai_mai_n1073_));
  NO3        m1045(.A(mai_mai_n1073_), .B(mai_mai_n307_), .C(mai_mai_n92_), .Y(mai_mai_n1074_));
  NOi21      m1046(.An(mai_mai_n1074_), .B(mai_mai_n1072_), .Y(mai_mai_n1075_));
  OR4        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1071_), .C(mai_mai_n1067_), .D(mai_mai_n1063_), .Y(mai_mai_n1076_));
  NA3        m1048(.A(mai_mai_n472_), .B(mai_mai_n337_), .C(mai_mai_n56_), .Y(mai_mai_n1077_));
  NO2        m1049(.A(mai_mai_n1077_), .B(mai_mai_n1066_), .Y(mai_mai_n1078_));
  NO4        m1050(.A(mai_mai_n1077_), .B(mai_mai_n595_), .C(mai_mai_n453_), .D(mai_mai_n45_), .Y(mai_mai_n1079_));
  NO2        m1051(.A(f), .B(c), .Y(mai_mai_n1080_));
  NOi21      m1052(.An(mai_mai_n1080_), .B(mai_mai_n445_), .Y(mai_mai_n1081_));
  NA2        m1053(.A(mai_mai_n1081_), .B(mai_mai_n59_), .Y(mai_mai_n1082_));
  OR2        m1054(.A(k), .B(i), .Y(mai_mai_n1083_));
  NO3        m1055(.A(mai_mai_n1083_), .B(mai_mai_n245_), .C(l), .Y(mai_mai_n1084_));
  NOi31      m1056(.An(mai_mai_n1084_), .B(mai_mai_n1082_), .C(j), .Y(mai_mai_n1085_));
  OR3        m1057(.A(mai_mai_n1085_), .B(mai_mai_n1079_), .C(mai_mai_n1078_), .Y(mai_mai_n1086_));
  OR3        m1058(.A(mai_mai_n1086_), .B(mai_mai_n1076_), .C(mai_mai_n1058_), .Y(mai02));
  OR2        m1059(.A(l), .B(k), .Y(mai_mai_n1088_));
  OR3        m1060(.A(h), .B(g), .C(f), .Y(mai_mai_n1089_));
  OR3        m1061(.A(n), .B(m), .C(i), .Y(mai_mai_n1090_));
  NO4        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1089_), .C(mai_mai_n1088_), .D(mai_mai_n1072_), .Y(mai_mai_n1091_));
  NOi31      m1063(.An(e), .B(d), .C(c), .Y(mai_mai_n1092_));
  AOI210     m1064(.A0(mai_mai_n1074_), .A1(mai_mai_n1092_), .B0(mai_mai_n1049_), .Y(mai_mai_n1093_));
  AN3        m1065(.A(g), .B(f), .C(c), .Y(mai_mai_n1094_));
  NA3        m1066(.A(mai_mai_n1094_), .B(mai_mai_n472_), .C(h), .Y(mai_mai_n1095_));
  OR2        m1067(.A(mai_mai_n1073_), .B(mai_mai_n307_), .Y(mai_mai_n1096_));
  OR2        m1068(.A(mai_mai_n1096_), .B(mai_mai_n1095_), .Y(mai_mai_n1097_));
  NO3        m1069(.A(mai_mai_n1077_), .B(mai_mai_n1048_), .C(mai_mai_n595_), .Y(mai_mai_n1098_));
  NO2        m1070(.A(mai_mai_n1098_), .B(mai_mai_n1063_), .Y(mai_mai_n1099_));
  NA3        m1071(.A(l), .B(k), .C(j), .Y(mai_mai_n1100_));
  NA2        m1072(.A(i), .B(h), .Y(mai_mai_n1101_));
  NO3        m1073(.A(mai_mai_n1101_), .B(mai_mai_n1100_), .C(mai_mai_n130_), .Y(mai_mai_n1102_));
  NO3        m1074(.A(mai_mai_n141_), .B(mai_mai_n285_), .C(mai_mai_n214_), .Y(mai_mai_n1103_));
  AOI210     m1075(.A0(mai_mai_n1103_), .A1(mai_mai_n1102_), .B0(mai_mai_n1067_), .Y(mai_mai_n1104_));
  NA3        m1076(.A(c), .B(b), .C(a), .Y(mai_mai_n1105_));
  NO3        m1077(.A(mai_mai_n1105_), .B(mai_mai_n908_), .C(mai_mai_n213_), .Y(mai_mai_n1106_));
  NO4        m1078(.A(mai_mai_n1073_), .B(mai_mai_n299_), .C(mai_mai_n49_), .D(mai_mai_n111_), .Y(mai_mai_n1107_));
  AOI210     m1079(.A0(mai_mai_n1107_), .A1(mai_mai_n1106_), .B0(mai_mai_n1078_), .Y(mai_mai_n1108_));
  AN4        m1080(.A(mai_mai_n1108_), .B(mai_mai_n1104_), .C(mai_mai_n1099_), .D(mai_mai_n1097_), .Y(mai_mai_n1109_));
  NO2        m1081(.A(mai_mai_n1053_), .B(mai_mai_n1051_), .Y(mai_mai_n1110_));
  NA2        m1082(.A(mai_mai_n1070_), .B(mai_mai_n1062_), .Y(mai_mai_n1111_));
  AOI210     m1083(.A0(mai_mai_n1111_), .A1(mai_mai_n1110_), .B0(mai_mai_n1044_), .Y(mai_mai_n1112_));
  NAi41      m1084(.An(mai_mai_n1091_), .B(mai_mai_n1112_), .C(mai_mai_n1109_), .D(mai_mai_n1093_), .Y(mai03));
  NOi41      m1085(.An(mai_mai_n812_), .B(mai_mai_n859_), .C(mai_mai_n848_), .D(mai_mai_n721_), .Y(mai_mai_n1114_));
  NO2        m1086(.A(mai_mai_n1114_), .B(mai_mai_n695_), .Y(mai_mai_n1115_));
  NOi31      m1087(.An(i), .B(k), .C(j), .Y(mai_mai_n1116_));
  NA4        m1088(.A(mai_mai_n1116_), .B(mai_mai_n1092_), .C(mai_mai_n346_), .D(mai_mai_n337_), .Y(mai_mai_n1117_));
  OAI210     m1089(.A0(mai_mai_n826_), .A1(mai_mai_n422_), .B0(mai_mai_n1117_), .Y(mai_mai_n1118_));
  NOi31      m1090(.An(m), .B(n), .C(f), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n1119_), .B(mai_mai_n51_), .Y(mai_mai_n1120_));
  AN2        m1092(.A(e), .B(c), .Y(mai_mai_n1121_));
  NA2        m1093(.A(mai_mai_n1121_), .B(a), .Y(mai_mai_n1122_));
  OAI220     m1094(.A0(mai_mai_n1122_), .A1(mai_mai_n1120_), .B0(mai_mai_n892_), .B1(mai_mai_n428_), .Y(mai_mai_n1123_));
  NA2        m1095(.A(mai_mai_n515_), .B(l), .Y(mai_mai_n1124_));
  NOi31      m1096(.An(mai_mai_n870_), .B(mai_mai_n1042_), .C(mai_mai_n1124_), .Y(mai_mai_n1125_));
  NO4        m1097(.A(mai_mai_n1125_), .B(mai_mai_n1123_), .C(mai_mai_n1118_), .D(mai_mai_n1004_), .Y(mai_mai_n1126_));
  NO2        m1098(.A(mai_mai_n285_), .B(a), .Y(mai_mai_n1127_));
  INV        m1099(.A(mai_mai_n1049_), .Y(mai_mai_n1128_));
  NO2        m1100(.A(mai_mai_n1101_), .B(mai_mai_n492_), .Y(mai_mai_n1129_));
  NO2        m1101(.A(mai_mai_n89_), .B(g), .Y(mai_mai_n1130_));
  AOI210     m1102(.A0(mai_mai_n1130_), .A1(mai_mai_n1129_), .B0(mai_mai_n1084_), .Y(mai_mai_n1131_));
  OR2        m1103(.A(mai_mai_n1131_), .B(mai_mai_n1082_), .Y(mai_mai_n1132_));
  NA3        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1128_), .C(mai_mai_n1126_), .Y(mai_mai_n1133_));
  NO4        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1115_), .C(mai_mai_n827_), .D(mai_mai_n572_), .Y(mai_mai_n1134_));
  NA2        m1106(.A(c), .B(b), .Y(mai_mai_n1135_));
  NO2        m1107(.A(mai_mai_n707_), .B(mai_mai_n1135_), .Y(mai_mai_n1136_));
  OAI210     m1108(.A0(mai_mai_n868_), .A1(mai_mai_n839_), .B0(mai_mai_n415_), .Y(mai_mai_n1137_));
  OAI210     m1109(.A0(mai_mai_n1137_), .A1(mai_mai_n869_), .B0(mai_mai_n1136_), .Y(mai_mai_n1138_));
  NAi21      m1110(.An(mai_mai_n423_), .B(mai_mai_n1136_), .Y(mai_mai_n1139_));
  NA3        m1111(.A(mai_mai_n429_), .B(mai_mai_n567_), .C(f), .Y(mai_mai_n1140_));
  OAI210     m1112(.A0(mai_mai_n556_), .A1(mai_mai_n39_), .B0(mai_mai_n1127_), .Y(mai_mai_n1141_));
  NA3        m1113(.A(mai_mai_n1141_), .B(mai_mai_n1140_), .C(mai_mai_n1139_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n261_), .B(mai_mai_n117_), .Y(mai_mai_n1143_));
  OAI210     m1115(.A0(mai_mai_n1143_), .A1(mai_mai_n289_), .B0(g), .Y(mai_mai_n1144_));
  NAi21      m1116(.An(f), .B(d), .Y(mai_mai_n1145_));
  NO2        m1117(.A(mai_mai_n1145_), .B(mai_mai_n1105_), .Y(mai_mai_n1146_));
  INV        m1118(.A(mai_mai_n1146_), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n1144_), .B(mai_mai_n1147_), .Y(mai_mai_n1148_));
  AOI210     m1120(.A0(mai_mai_n1148_), .A1(mai_mai_n112_), .B0(mai_mai_n1142_), .Y(mai_mai_n1149_));
  NA2        m1121(.A(mai_mai_n475_), .B(mai_mai_n474_), .Y(mai_mai_n1150_));
  NO2        m1122(.A(mai_mai_n184_), .B(mai_mai_n238_), .Y(mai_mai_n1151_));
  NA2        m1123(.A(mai_mai_n1151_), .B(m), .Y(mai_mai_n1152_));
  NA3        m1124(.A(mai_mai_n923_), .B(mai_mai_n1124_), .C(mai_mai_n478_), .Y(mai_mai_n1153_));
  OAI210     m1125(.A0(mai_mai_n1153_), .A1(mai_mai_n312_), .B0(mai_mai_n476_), .Y(mai_mai_n1154_));
  AOI210     m1126(.A0(mai_mai_n1154_), .A1(mai_mai_n1150_), .B0(mai_mai_n1152_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n569_), .B(mai_mai_n410_), .Y(mai_mai_n1156_));
  NA2        m1128(.A(mai_mai_n158_), .B(mai_mai_n33_), .Y(mai_mai_n1157_));
  AOI210     m1129(.A0(mai_mai_n970_), .A1(mai_mai_n1157_), .B0(mai_mai_n214_), .Y(mai_mai_n1158_));
  OAI210     m1130(.A0(mai_mai_n1158_), .A1(mai_mai_n449_), .B0(mai_mai_n1146_), .Y(mai_mai_n1159_));
  NO2        m1131(.A(mai_mai_n373_), .B(mai_mai_n372_), .Y(mai_mai_n1160_));
  AOI210     m1132(.A0(mai_mai_n1151_), .A1(mai_mai_n431_), .B0(mai_mai_n964_), .Y(mai_mai_n1161_));
  NAi41      m1133(.An(mai_mai_n1160_), .B(mai_mai_n1161_), .C(mai_mai_n1159_), .D(mai_mai_n1156_), .Y(mai_mai_n1162_));
  NO2        m1134(.A(mai_mai_n1162_), .B(mai_mai_n1155_), .Y(mai_mai_n1163_));
  NA4        m1135(.A(mai_mai_n1163_), .B(mai_mai_n1149_), .C(mai_mai_n1138_), .D(mai_mai_n1134_), .Y(mai00));
  AOI210     m1136(.A0(mai_mai_n298_), .A1(mai_mai_n214_), .B0(mai_mai_n277_), .Y(mai_mai_n1165_));
  NO2        m1137(.A(mai_mai_n1165_), .B(mai_mai_n586_), .Y(mai_mai_n1166_));
  AOI210     m1138(.A0(mai_mai_n905_), .A1(mai_mai_n947_), .B0(mai_mai_n1118_), .Y(mai_mai_n1167_));
  NO2        m1139(.A(mai_mai_n1098_), .B(mai_mai_n964_), .Y(mai_mai_n1168_));
  NA3        m1140(.A(mai_mai_n1168_), .B(mai_mai_n1167_), .C(mai_mai_n1005_), .Y(mai_mai_n1169_));
  NA2        m1141(.A(mai_mai_n517_), .B(f), .Y(mai_mai_n1170_));
  OAI210     m1142(.A0(mai_mai_n1012_), .A1(mai_mai_n40_), .B0(mai_mai_n649_), .Y(mai_mai_n1171_));
  NA3        m1143(.A(mai_mai_n1171_), .B(mai_mai_n257_), .C(n), .Y(mai_mai_n1172_));
  AOI210     m1144(.A0(mai_mai_n1172_), .A1(mai_mai_n1170_), .B0(mai_mai_n1053_), .Y(mai_mai_n1173_));
  NO4        m1145(.A(mai_mai_n1173_), .B(mai_mai_n1169_), .C(mai_mai_n1166_), .D(mai_mai_n1076_), .Y(mai_mai_n1174_));
  NA3        m1146(.A(mai_mai_n168_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1175_));
  NA3        m1147(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1176_));
  NOi31      m1148(.An(n), .B(m), .C(i), .Y(mai_mai_n1177_));
  NA3        m1149(.A(mai_mai_n1177_), .B(mai_mai_n652_), .C(mai_mai_n51_), .Y(mai_mai_n1178_));
  OAI210     m1150(.A0(mai_mai_n1176_), .A1(mai_mai_n1175_), .B0(mai_mai_n1178_), .Y(mai_mai_n1179_));
  INV        m1151(.A(mai_mai_n585_), .Y(mai_mai_n1180_));
  NO3        m1152(.A(mai_mai_n1180_), .B(mai_mai_n1179_), .C(mai_mai_n1160_), .Y(mai_mai_n1181_));
  NO4        m1153(.A(mai_mai_n495_), .B(mai_mai_n358_), .C(mai_mai_n1135_), .D(mai_mai_n59_), .Y(mai_mai_n1182_));
  NA3        m1154(.A(mai_mai_n385_), .B(mai_mai_n221_), .C(g), .Y(mai_mai_n1183_));
  OA220      m1155(.A0(mai_mai_n1183_), .A1(mai_mai_n1176_), .B0(mai_mai_n386_), .B1(mai_mai_n133_), .Y(mai_mai_n1184_));
  NO2        m1156(.A(h), .B(g), .Y(mai_mai_n1185_));
  NA4        m1157(.A(mai_mai_n507_), .B(mai_mai_n472_), .C(mai_mai_n1185_), .D(mai_mai_n1041_), .Y(mai_mai_n1186_));
  NA2        m1158(.A(mai_mai_n951_), .B(mai_mai_n584_), .Y(mai_mai_n1187_));
  NA3        m1159(.A(mai_mai_n1187_), .B(mai_mai_n1186_), .C(mai_mai_n1184_), .Y(mai_mai_n1188_));
  NO3        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1182_), .C(mai_mai_n267_), .Y(mai_mai_n1189_));
  INV        m1161(.A(mai_mai_n324_), .Y(mai_mai_n1190_));
  INV        m1162(.A(mai_mai_n587_), .Y(mai_mai_n1191_));
  NA2        m1163(.A(mai_mai_n1191_), .B(mai_mai_n1190_), .Y(mai_mai_n1192_));
  NO2        m1164(.A(mai_mai_n240_), .B(mai_mai_n183_), .Y(mai_mai_n1193_));
  NA2        m1165(.A(mai_mai_n1193_), .B(mai_mai_n429_), .Y(mai_mai_n1194_));
  NA3        m1166(.A(mai_mai_n181_), .B(mai_mai_n111_), .C(g), .Y(mai_mai_n1195_));
  NA3        m1167(.A(mai_mai_n472_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1196_));
  NOi31      m1168(.An(mai_mai_n877_), .B(mai_mai_n1196_), .C(mai_mai_n1195_), .Y(mai_mai_n1197_));
  NAi31      m1169(.An(mai_mai_n188_), .B(mai_mai_n865_), .C(mai_mai_n472_), .Y(mai_mai_n1198_));
  NAi31      m1170(.An(mai_mai_n1197_), .B(mai_mai_n1198_), .C(mai_mai_n1194_), .Y(mai_mai_n1199_));
  NO2        m1171(.A(mai_mai_n276_), .B(mai_mai_n75_), .Y(mai_mai_n1200_));
  NO3        m1172(.A(mai_mai_n428_), .B(mai_mai_n835_), .C(n), .Y(mai_mai_n1201_));
  AOI210     m1173(.A0(mai_mai_n1201_), .A1(mai_mai_n1200_), .B0(mai_mai_n1091_), .Y(mai_mai_n1202_));
  NAi31      m1174(.An(mai_mai_n1056_), .B(mai_mai_n1202_), .C(mai_mai_n74_), .Y(mai_mai_n1203_));
  NO4        m1175(.A(mai_mai_n1203_), .B(mai_mai_n1199_), .C(mai_mai_n1192_), .D(mai_mai_n527_), .Y(mai_mai_n1204_));
  AN3        m1176(.A(mai_mai_n1204_), .B(mai_mai_n1189_), .C(mai_mai_n1181_), .Y(mai_mai_n1205_));
  NA3        m1177(.A(mai_mai_n1119_), .B(mai_mai_n613_), .C(mai_mai_n471_), .Y(mai_mai_n1206_));
  NA3        m1178(.A(mai_mai_n1206_), .B(mai_mai_n570_), .C(mai_mai_n243_), .Y(mai_mai_n1207_));
  OAI210     m1179(.A0(mai_mai_n470_), .A1(mai_mai_n118_), .B0(mai_mai_n871_), .Y(mai_mai_n1208_));
  AOI220     m1180(.A0(mai_mai_n1208_), .A1(mai_mai_n1153_), .B0(mai_mai_n569_), .B1(mai_mai_n410_), .Y(mai_mai_n1209_));
  OR4        m1181(.A(mai_mai_n1053_), .B(mai_mai_n273_), .C(mai_mai_n223_), .D(e), .Y(mai_mai_n1210_));
  NO2        m1182(.A(mai_mai_n217_), .B(mai_mai_n214_), .Y(mai_mai_n1211_));
  NA2        m1183(.A(n), .B(e), .Y(mai_mai_n1212_));
  NO2        m1184(.A(mai_mai_n1212_), .B(mai_mai_n146_), .Y(mai_mai_n1213_));
  AOI220     m1185(.A0(mai_mai_n1213_), .A1(mai_mai_n275_), .B0(mai_mai_n852_), .B1(mai_mai_n1211_), .Y(mai_mai_n1214_));
  OAI210     m1186(.A0(mai_mai_n359_), .A1(mai_mai_n313_), .B0(mai_mai_n451_), .Y(mai_mai_n1215_));
  NA4        m1187(.A(mai_mai_n1215_), .B(mai_mai_n1214_), .C(mai_mai_n1210_), .D(mai_mai_n1209_), .Y(mai_mai_n1216_));
  AOI210     m1188(.A0(mai_mai_n1213_), .A1(mai_mai_n856_), .B0(mai_mai_n827_), .Y(mai_mai_n1217_));
  AOI220     m1189(.A0(mai_mai_n960_), .A1(mai_mai_n584_), .B0(mai_mai_n652_), .B1(mai_mai_n246_), .Y(mai_mai_n1218_));
  NO2        m1190(.A(mai_mai_n68_), .B(h), .Y(mai_mai_n1219_));
  NO3        m1191(.A(mai_mai_n1053_), .B(mai_mai_n1051_), .C(mai_mai_n732_), .Y(mai_mai_n1220_));
  NO2        m1192(.A(mai_mai_n1088_), .B(mai_mai_n130_), .Y(mai_mai_n1221_));
  AN2        m1193(.A(mai_mai_n1221_), .B(mai_mai_n1103_), .Y(mai_mai_n1222_));
  OAI210     m1194(.A0(mai_mai_n1222_), .A1(mai_mai_n1220_), .B0(mai_mai_n1219_), .Y(mai_mai_n1223_));
  NA4        m1195(.A(mai_mai_n1223_), .B(mai_mai_n1218_), .C(mai_mai_n1217_), .D(mai_mai_n872_), .Y(mai_mai_n1224_));
  NO3        m1196(.A(mai_mai_n1224_), .B(mai_mai_n1216_), .C(mai_mai_n1207_), .Y(mai_mai_n1225_));
  NA2        m1197(.A(mai_mai_n840_), .B(mai_mai_n763_), .Y(mai_mai_n1226_));
  NA4        m1198(.A(mai_mai_n1226_), .B(mai_mai_n1225_), .C(mai_mai_n1205_), .D(mai_mai_n1174_), .Y(mai01));
  AN2        m1199(.A(mai_mai_n1030_), .B(mai_mai_n1028_), .Y(mai_mai_n1228_));
  NO4        m1200(.A(mai_mai_n808_), .B(mai_mai_n800_), .C(mai_mai_n486_), .D(mai_mai_n283_), .Y(mai_mai_n1229_));
  NA2        m1201(.A(mai_mai_n396_), .B(i), .Y(mai_mai_n1230_));
  NA3        m1202(.A(mai_mai_n1230_), .B(mai_mai_n1229_), .C(mai_mai_n1228_), .Y(mai_mai_n1231_));
  NA2        m1203(.A(mai_mai_n562_), .B(mai_mai_n272_), .Y(mai_mai_n1232_));
  NA2        m1204(.A(mai_mai_n967_), .B(mai_mai_n1232_), .Y(mai_mai_n1233_));
  NA3        m1205(.A(mai_mai_n1233_), .B(mai_mai_n921_), .C(mai_mai_n336_), .Y(mai_mai_n1234_));
  NA2        m1206(.A(mai_mai_n45_), .B(f), .Y(mai_mai_n1235_));
  NA2        m1207(.A(mai_mai_n714_), .B(mai_mai_n97_), .Y(mai_mai_n1236_));
  NO2        m1208(.A(mai_mai_n1236_), .B(mai_mai_n1235_), .Y(mai_mai_n1237_));
  NO2        m1209(.A(mai_mai_n787_), .B(mai_mai_n611_), .Y(mai_mai_n1238_));
  AOI210     m1210(.A0(mai_mai_n1237_), .A1(mai_mai_n639_), .B0(mai_mai_n1238_), .Y(mai_mai_n1239_));
  INV        m1211(.A(mai_mai_n116_), .Y(mai_mai_n1240_));
  OR2        m1212(.A(mai_mai_n1240_), .B(mai_mai_n594_), .Y(mai_mai_n1241_));
  NAi41      m1213(.An(mai_mai_n161_), .B(mai_mai_n1241_), .C(mai_mai_n1239_), .D(mai_mai_n904_), .Y(mai_mai_n1242_));
  NO3        m1214(.A(mai_mai_n788_), .B(mai_mai_n678_), .C(mai_mai_n520_), .Y(mai_mai_n1243_));
  OR2        m1215(.A(mai_mai_n198_), .B(mai_mai_n196_), .Y(mai_mai_n1244_));
  NA3        m1216(.A(mai_mai_n1244_), .B(mai_mai_n1243_), .C(mai_mai_n136_), .Y(mai_mai_n1245_));
  NO4        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1242_), .C(mai_mai_n1234_), .D(mai_mai_n1231_), .Y(mai_mai_n1246_));
  INV        m1218(.A(mai_mai_n1183_), .Y(mai_mai_n1247_));
  OAI210     m1219(.A0(mai_mai_n1247_), .A1(mai_mai_n301_), .B0(mai_mai_n538_), .Y(mai_mai_n1248_));
  NA2        m1220(.A(mai_mai_n545_), .B(mai_mai_n398_), .Y(mai_mai_n1249_));
  NOi21      m1221(.An(mai_mai_n571_), .B(mai_mai_n591_), .Y(mai_mai_n1250_));
  NA2        m1222(.A(mai_mai_n1250_), .B(mai_mai_n1249_), .Y(mai_mai_n1251_));
  AOI210     m1223(.A0(mai_mai_n207_), .A1(mai_mai_n91_), .B0(mai_mai_n213_), .Y(mai_mai_n1252_));
  OAI210     m1224(.A0(mai_mai_n815_), .A1(mai_mai_n429_), .B0(mai_mai_n1252_), .Y(mai_mai_n1253_));
  AN3        m1225(.A(m), .B(l), .C(k), .Y(mai_mai_n1254_));
  OAI210     m1226(.A0(mai_mai_n361_), .A1(mai_mai_n34_), .B0(mai_mai_n1254_), .Y(mai_mai_n1255_));
  NA2        m1227(.A(mai_mai_n206_), .B(mai_mai_n34_), .Y(mai_mai_n1256_));
  AO210      m1228(.A0(mai_mai_n1256_), .A1(mai_mai_n1255_), .B0(mai_mai_n335_), .Y(mai_mai_n1257_));
  NA4        m1229(.A(mai_mai_n1257_), .B(mai_mai_n1253_), .C(mai_mai_n1251_), .D(mai_mai_n1248_), .Y(mai_mai_n1258_));
  AOI210     m1230(.A0(mai_mai_n603_), .A1(mai_mai_n116_), .B0(mai_mai_n609_), .Y(mai_mai_n1259_));
  OAI210     m1231(.A0(mai_mai_n1240_), .A1(mai_mai_n602_), .B0(mai_mai_n1259_), .Y(mai_mai_n1260_));
  NA2        m1232(.A(mai_mai_n282_), .B(mai_mai_n198_), .Y(mai_mai_n1261_));
  NA2        m1233(.A(mai_mai_n1261_), .B(mai_mai_n669_), .Y(mai_mai_n1262_));
  NO3        m1234(.A(mai_mai_n826_), .B(mai_mai_n207_), .C(mai_mai_n408_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n1263_), .B(mai_mai_n964_), .Y(mai_mai_n1264_));
  OAI210     m1236(.A0(mai_mai_n1237_), .A1(mai_mai_n329_), .B0(mai_mai_n679_), .Y(mai_mai_n1265_));
  NA4        m1237(.A(mai_mai_n1265_), .B(mai_mai_n1264_), .C(mai_mai_n1262_), .D(mai_mai_n791_), .Y(mai_mai_n1266_));
  NO3        m1238(.A(mai_mai_n1266_), .B(mai_mai_n1260_), .C(mai_mai_n1258_), .Y(mai_mai_n1267_));
  NA2        m1239(.A(mai_mai_n513_), .B(mai_mai_n58_), .Y(mai_mai_n1268_));
  INV        m1240(.A(mai_mai_n1179_), .Y(mai_mai_n1269_));
  NA3        m1241(.A(mai_mai_n1269_), .B(mai_mai_n1268_), .C(mai_mai_n762_), .Y(mai_mai_n1270_));
  NO2        m1242(.A(mai_mai_n974_), .B(mai_mai_n233_), .Y(mai_mai_n1271_));
  NO2        m1243(.A(mai_mai_n975_), .B(mai_mai_n564_), .Y(mai_mai_n1272_));
  OAI210     m1244(.A0(mai_mai_n1272_), .A1(mai_mai_n1271_), .B0(mai_mai_n344_), .Y(mai_mai_n1273_));
  NA2        m1245(.A(mai_mai_n579_), .B(mai_mai_n577_), .Y(mai_mai_n1274_));
  NO3        m1246(.A(mai_mai_n81_), .B(mai_mai_n299_), .C(mai_mai_n45_), .Y(mai_mai_n1275_));
  NA2        m1247(.A(mai_mai_n1275_), .B(mai_mai_n561_), .Y(mai_mai_n1276_));
  NA2        m1248(.A(mai_mai_n1276_), .B(mai_mai_n1274_), .Y(mai_mai_n1277_));
  OR2        m1249(.A(mai_mai_n1183_), .B(mai_mai_n1176_), .Y(mai_mai_n1278_));
  NA2        m1250(.A(mai_mai_n1275_), .B(mai_mai_n818_), .Y(mai_mai_n1279_));
  NA3        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1278_), .C(mai_mai_n388_), .Y(mai_mai_n1280_));
  NOi41      m1252(.An(mai_mai_n1273_), .B(mai_mai_n1280_), .C(mai_mai_n1277_), .D(mai_mai_n1270_), .Y(mai_mai_n1281_));
  NO2        m1253(.A(mai_mai_n129_), .B(mai_mai_n45_), .Y(mai_mai_n1282_));
  NO2        m1254(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1283_));
  AO220      m1255(.A0(mai_mai_n1283_), .A1(mai_mai_n627_), .B0(mai_mai_n1282_), .B1(mai_mai_n712_), .Y(mai_mai_n1284_));
  NA2        m1256(.A(mai_mai_n1284_), .B(mai_mai_n344_), .Y(mai_mai_n1285_));
  NO3        m1257(.A(mai_mai_n1101_), .B(mai_mai_n178_), .C(mai_mai_n89_), .Y(mai_mai_n1286_));
  NA2        m1258(.A(mai_mai_n1275_), .B(mai_mai_n978_), .Y(mai_mai_n1287_));
  NA2        m1259(.A(mai_mai_n1287_), .B(mai_mai_n1285_), .Y(mai_mai_n1288_));
  NO2        m1260(.A(mai_mai_n618_), .B(mai_mai_n617_), .Y(mai_mai_n1289_));
  NO4        m1261(.A(mai_mai_n1101_), .B(mai_mai_n1289_), .C(mai_mai_n176_), .D(mai_mai_n89_), .Y(mai_mai_n1290_));
  NO3        m1262(.A(mai_mai_n1290_), .B(mai_mai_n1288_), .C(mai_mai_n641_), .Y(mai_mai_n1291_));
  NA4        m1263(.A(mai_mai_n1291_), .B(mai_mai_n1281_), .C(mai_mai_n1267_), .D(mai_mai_n1246_), .Y(mai06));
  NO2        m1264(.A(mai_mai_n409_), .B(mai_mai_n568_), .Y(mai_mai_n1293_));
  INV        m1265(.A(mai_mai_n739_), .Y(mai_mai_n1294_));
  NA2        m1266(.A(mai_mai_n1294_), .B(mai_mai_n1293_), .Y(mai_mai_n1295_));
  NO2        m1267(.A(mai_mai_n225_), .B(mai_mai_n102_), .Y(mai_mai_n1296_));
  OAI210     m1268(.A0(mai_mai_n1296_), .A1(mai_mai_n1286_), .B0(mai_mai_n384_), .Y(mai_mai_n1297_));
  NO3        m1269(.A(mai_mai_n607_), .B(mai_mai_n813_), .C(mai_mai_n610_), .Y(mai_mai_n1298_));
  OR2        m1270(.A(mai_mai_n1298_), .B(mai_mai_n892_), .Y(mai_mai_n1299_));
  NA4        m1271(.A(mai_mai_n1299_), .B(mai_mai_n1297_), .C(mai_mai_n1295_), .D(mai_mai_n1273_), .Y(mai_mai_n1300_));
  NO3        m1272(.A(mai_mai_n1300_), .B(mai_mai_n1277_), .C(mai_mai_n256_), .Y(mai_mai_n1301_));
  NO2        m1273(.A(mai_mai_n299_), .B(mai_mai_n45_), .Y(mai_mai_n1302_));
  AOI210     m1274(.A0(mai_mai_n1302_), .A1(mai_mai_n979_), .B0(mai_mai_n1271_), .Y(mai_mai_n1303_));
  AOI210     m1275(.A0(mai_mai_n1302_), .A1(mai_mai_n565_), .B0(mai_mai_n1284_), .Y(mai_mai_n1304_));
  AOI210     m1276(.A0(mai_mai_n1304_), .A1(mai_mai_n1303_), .B0(mai_mai_n341_), .Y(mai_mai_n1305_));
  INV        m1277(.A(mai_mai_n677_), .Y(mai_mai_n1306_));
  NA2        m1278(.A(mai_mai_n1306_), .B(mai_mai_n645_), .Y(mai_mai_n1307_));
  NO2        m1279(.A(mai_mai_n523_), .B(mai_mai_n173_), .Y(mai_mai_n1308_));
  NOi21      m1280(.An(mai_mai_n135_), .B(mai_mai_n45_), .Y(mai_mai_n1309_));
  NO2        m1281(.A(mai_mai_n614_), .B(mai_mai_n1120_), .Y(mai_mai_n1310_));
  OAI210     m1282(.A0(mai_mai_n465_), .A1(mai_mai_n249_), .B0(mai_mai_n915_), .Y(mai_mai_n1311_));
  NO4        m1283(.A(mai_mai_n1311_), .B(mai_mai_n1310_), .C(mai_mai_n1309_), .D(mai_mai_n1308_), .Y(mai_mai_n1312_));
  OR2        m1284(.A(mai_mai_n608_), .B(mai_mai_n606_), .Y(mai_mai_n1313_));
  INV        m1285(.A(mai_mai_n1313_), .Y(mai_mai_n1314_));
  NA3        m1286(.A(mai_mai_n1314_), .B(mai_mai_n1312_), .C(mai_mai_n1307_), .Y(mai_mai_n1315_));
  NO2        m1287(.A(mai_mai_n753_), .B(mai_mai_n370_), .Y(mai_mai_n1316_));
  NO3        m1288(.A(mai_mai_n679_), .B(mai_mai_n764_), .C(mai_mai_n639_), .Y(mai_mai_n1317_));
  NOi21      m1289(.An(mai_mai_n1316_), .B(mai_mai_n1317_), .Y(mai_mai_n1318_));
  AN2        m1290(.A(mai_mai_n960_), .B(mai_mai_n648_), .Y(mai_mai_n1319_));
  NO4        m1291(.A(mai_mai_n1319_), .B(mai_mai_n1318_), .C(mai_mai_n1315_), .D(mai_mai_n1305_), .Y(mai_mai_n1320_));
  NO2        m1292(.A(mai_mai_n807_), .B(mai_mai_n278_), .Y(mai_mai_n1321_));
  OAI220     m1293(.A0(mai_mai_n739_), .A1(mai_mai_n47_), .B0(mai_mai_n225_), .B1(mai_mai_n620_), .Y(mai_mai_n1322_));
  OAI210     m1294(.A0(mai_mai_n278_), .A1(c), .B0(mai_mai_n644_), .Y(mai_mai_n1323_));
  AOI220     m1295(.A0(mai_mai_n1323_), .A1(mai_mai_n1322_), .B0(mai_mai_n1321_), .B1(mai_mai_n268_), .Y(mai_mai_n1324_));
  NO3        m1296(.A(mai_mai_n245_), .B(mai_mai_n102_), .C(mai_mai_n285_), .Y(mai_mai_n1325_));
  OAI220     m1297(.A0(mai_mai_n704_), .A1(mai_mai_n249_), .B0(mai_mai_n519_), .B1(mai_mai_n523_), .Y(mai_mai_n1326_));
  OAI210     m1298(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1327_));
  NO3        m1299(.A(mai_mai_n1327_), .B(mai_mai_n605_), .C(j), .Y(mai_mai_n1328_));
  NOi21      m1300(.An(mai_mai_n1328_), .B(mai_mai_n673_), .Y(mai_mai_n1329_));
  NO4        m1301(.A(mai_mai_n1329_), .B(mai_mai_n1326_), .C(mai_mai_n1325_), .D(mai_mai_n1123_), .Y(mai_mai_n1330_));
  NA4        m1302(.A(mai_mai_n798_), .B(mai_mai_n797_), .C(mai_mai_n439_), .D(mai_mai_n884_), .Y(mai_mai_n1331_));
  NAi31      m1303(.An(mai_mai_n753_), .B(mai_mai_n1331_), .C(mai_mai_n206_), .Y(mai_mai_n1332_));
  NA4        m1304(.A(mai_mai_n1332_), .B(mai_mai_n1330_), .C(mai_mai_n1324_), .D(mai_mai_n1218_), .Y(mai_mai_n1333_));
  NOi31      m1305(.An(mai_mai_n1298_), .B(mai_mai_n469_), .C(mai_mai_n397_), .Y(mai_mai_n1334_));
  OR3        m1306(.A(mai_mai_n1334_), .B(mai_mai_n787_), .C(mai_mai_n548_), .Y(mai_mai_n1335_));
  OR3        m1307(.A(mai_mai_n372_), .B(mai_mai_n225_), .C(mai_mai_n620_), .Y(mai_mai_n1336_));
  AOI210     m1308(.A0(mai_mai_n579_), .A1(mai_mai_n451_), .B0(mai_mai_n374_), .Y(mai_mai_n1337_));
  NA3        m1309(.A(mai_mai_n1337_), .B(mai_mai_n1336_), .C(mai_mai_n1335_), .Y(mai_mai_n1338_));
  AN2        m1310(.A(mai_mai_n933_), .B(mai_mai_n932_), .Y(mai_mai_n1339_));
  NO4        m1311(.A(mai_mai_n1339_), .B(mai_mai_n882_), .C(mai_mai_n509_), .D(mai_mai_n489_), .Y(mai_mai_n1340_));
  NA2        m1312(.A(mai_mai_n1340_), .B(mai_mai_n1279_), .Y(mai_mai_n1341_));
  NAi21      m1313(.An(j), .B(i), .Y(mai_mai_n1342_));
  NO4        m1314(.A(mai_mai_n1289_), .B(mai_mai_n1342_), .C(mai_mai_n445_), .D(mai_mai_n236_), .Y(mai_mai_n1343_));
  NO4        m1315(.A(mai_mai_n1343_), .B(mai_mai_n1341_), .C(mai_mai_n1338_), .D(mai_mai_n1333_), .Y(mai_mai_n1344_));
  NA4        m1316(.A(mai_mai_n1344_), .B(mai_mai_n1320_), .C(mai_mai_n1301_), .D(mai_mai_n1291_), .Y(mai07));
  NOi21      m1317(.An(j), .B(k), .Y(mai_mai_n1346_));
  NA4        m1318(.A(mai_mai_n181_), .B(mai_mai_n108_), .C(mai_mai_n1346_), .D(f), .Y(mai_mai_n1347_));
  NAi32      m1319(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1348_));
  NO3        m1320(.A(mai_mai_n1348_), .B(g), .C(f), .Y(mai_mai_n1349_));
  OAI210     m1321(.A0(mai_mai_n323_), .A1(mai_mai_n491_), .B0(mai_mai_n1349_), .Y(mai_mai_n1350_));
  NAi21      m1322(.An(f), .B(c), .Y(mai_mai_n1351_));
  OR2        m1323(.A(e), .B(d), .Y(mai_mai_n1352_));
  OAI220     m1324(.A0(mai_mai_n1352_), .A1(mai_mai_n1351_), .B0(mai_mai_n633_), .B1(mai_mai_n325_), .Y(mai_mai_n1353_));
  NA3        m1325(.A(mai_mai_n1353_), .B(mai_mai_n1065_), .C(mai_mai_n181_), .Y(mai_mai_n1354_));
  NOi31      m1326(.An(n), .B(m), .C(b), .Y(mai_mai_n1355_));
  NO3        m1327(.A(mai_mai_n130_), .B(mai_mai_n453_), .C(h), .Y(mai_mai_n1356_));
  NA3        m1328(.A(mai_mai_n1354_), .B(mai_mai_n1350_), .C(mai_mai_n1347_), .Y(mai_mai_n1357_));
  NOi41      m1329(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1358_));
  NOi21      m1330(.An(h), .B(k), .Y(mai_mai_n1359_));
  NO2        m1331(.A(k), .B(i), .Y(mai_mai_n1360_));
  NA3        m1332(.A(mai_mai_n1360_), .B(mai_mai_n903_), .C(mai_mai_n181_), .Y(mai_mai_n1361_));
  NA2        m1333(.A(mai_mai_n89_), .B(mai_mai_n45_), .Y(mai_mai_n1362_));
  NO2        m1334(.A(mai_mai_n1059_), .B(mai_mai_n445_), .Y(mai_mai_n1363_));
  NA3        m1335(.A(mai_mai_n1363_), .B(mai_mai_n1362_), .C(mai_mai_n214_), .Y(mai_mai_n1364_));
  NO2        m1336(.A(mai_mai_n1073_), .B(mai_mai_n307_), .Y(mai_mai_n1365_));
  NA2        m1337(.A(mai_mai_n549_), .B(mai_mai_n82_), .Y(mai_mai_n1366_));
  NA2        m1338(.A(mai_mai_n1219_), .B(mai_mai_n293_), .Y(mai_mai_n1367_));
  NA4        m1339(.A(mai_mai_n1367_), .B(mai_mai_n1366_), .C(mai_mai_n1364_), .D(mai_mai_n1361_), .Y(mai_mai_n1368_));
  NO2        m1340(.A(mai_mai_n1368_), .B(mai_mai_n1357_), .Y(mai_mai_n1369_));
  NO3        m1341(.A(e), .B(d), .C(c), .Y(mai_mai_n1370_));
  NA2        m1342(.A(mai_mai_n1556_), .B(mai_mai_n1370_), .Y(mai_mai_n1371_));
  NO2        m1343(.A(mai_mai_n1371_), .B(mai_mai_n214_), .Y(mai_mai_n1372_));
  OR2        m1344(.A(h), .B(f), .Y(mai_mai_n1373_));
  NO3        m1345(.A(n), .B(m), .C(i), .Y(mai_mai_n1374_));
  OAI210     m1346(.A0(mai_mai_n1121_), .A1(mai_mai_n156_), .B0(mai_mai_n1374_), .Y(mai_mai_n1375_));
  NO2        m1347(.A(mai_mai_n1375_), .B(mai_mai_n1373_), .Y(mai_mai_n1376_));
  NA3        m1348(.A(mai_mai_n701_), .B(mai_mai_n687_), .C(mai_mai_n111_), .Y(mai_mai_n1377_));
  NO2        m1349(.A(mai_mai_n1377_), .B(mai_mai_n45_), .Y(mai_mai_n1378_));
  NA2        m1350(.A(mai_mai_n1374_), .B(mai_mai_n643_), .Y(mai_mai_n1379_));
  NO2        m1351(.A(l), .B(k), .Y(mai_mai_n1380_));
  NOi41      m1352(.An(mai_mai_n554_), .B(mai_mai_n1380_), .C(mai_mai_n484_), .D(mai_mai_n445_), .Y(mai_mai_n1381_));
  NO3        m1353(.A(mai_mai_n445_), .B(d), .C(c), .Y(mai_mai_n1382_));
  NO4        m1354(.A(mai_mai_n1381_), .B(mai_mai_n1378_), .C(mai_mai_n1376_), .D(mai_mai_n1372_), .Y(mai_mai_n1383_));
  NO2        m1355(.A(mai_mai_n147_), .B(h), .Y(mai_mai_n1384_));
  NO2        m1356(.A(mai_mai_n1083_), .B(l), .Y(mai_mai_n1385_));
  NO2        m1357(.A(g), .B(c), .Y(mai_mai_n1386_));
  NA3        m1358(.A(mai_mai_n1386_), .B(mai_mai_n141_), .C(mai_mai_n189_), .Y(mai_mai_n1387_));
  NO2        m1359(.A(mai_mai_n1387_), .B(mai_mai_n1385_), .Y(mai_mai_n1388_));
  NA2        m1360(.A(mai_mai_n1388_), .B(mai_mai_n181_), .Y(mai_mai_n1389_));
  OAI210     m1361(.A0(mai_mai_n1359_), .A1(mai_mai_n213_), .B0(mai_mai_n1083_), .Y(mai_mai_n1390_));
  NO2        m1362(.A(mai_mai_n456_), .B(a), .Y(mai_mai_n1391_));
  NA3        m1363(.A(mai_mai_n1391_), .B(mai_mai_n1390_), .C(mai_mai_n112_), .Y(mai_mai_n1392_));
  NO2        m1364(.A(i), .B(h), .Y(mai_mai_n1393_));
  NA2        m1365(.A(mai_mai_n1393_), .B(mai_mai_n221_), .Y(mai_mai_n1394_));
  AOI210     m1366(.A0(mai_mai_n1145_), .A1(h), .B0(mai_mai_n416_), .Y(mai_mai_n1395_));
  NA2        m1367(.A(mai_mai_n137_), .B(mai_mai_n221_), .Y(mai_mai_n1396_));
  AOI210     m1368(.A0(mai_mai_n257_), .A1(mai_mai_n114_), .B0(mai_mai_n538_), .Y(mai_mai_n1397_));
  OAI220     m1369(.A0(mai_mai_n1397_), .A1(mai_mai_n1394_), .B0(mai_mai_n1396_), .B1(mai_mai_n1395_), .Y(mai_mai_n1398_));
  NO2        m1370(.A(mai_mai_n760_), .B(mai_mai_n190_), .Y(mai_mai_n1399_));
  NOi31      m1371(.An(m), .B(n), .C(b), .Y(mai_mai_n1400_));
  NOi31      m1372(.An(f), .B(d), .C(c), .Y(mai_mai_n1401_));
  NA2        m1373(.A(mai_mai_n1401_), .B(mai_mai_n1400_), .Y(mai_mai_n1402_));
  INV        m1374(.A(mai_mai_n1402_), .Y(mai_mai_n1403_));
  NO3        m1375(.A(mai_mai_n1403_), .B(mai_mai_n1399_), .C(mai_mai_n1398_), .Y(mai_mai_n1404_));
  NA2        m1376(.A(mai_mai_n1094_), .B(mai_mai_n472_), .Y(mai_mai_n1405_));
  NO4        m1377(.A(mai_mai_n1405_), .B(mai_mai_n1068_), .C(mai_mai_n445_), .D(mai_mai_n45_), .Y(mai_mai_n1406_));
  OAI210     m1378(.A0(mai_mai_n184_), .A1(mai_mai_n533_), .B0(mai_mai_n1069_), .Y(mai_mai_n1407_));
  NO3        m1379(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1408_));
  INV        m1380(.A(mai_mai_n1407_), .Y(mai_mai_n1409_));
  NO2        m1381(.A(mai_mai_n1409_), .B(mai_mai_n1406_), .Y(mai_mai_n1410_));
  AN4        m1382(.A(mai_mai_n1410_), .B(mai_mai_n1404_), .C(mai_mai_n1392_), .D(mai_mai_n1389_), .Y(mai_mai_n1411_));
  NA2        m1383(.A(mai_mai_n1355_), .B(mai_mai_n381_), .Y(mai_mai_n1412_));
  NO2        m1384(.A(mai_mai_n1412_), .B(mai_mai_n1050_), .Y(mai_mai_n1413_));
  NA2        m1385(.A(mai_mai_n1382_), .B(mai_mai_n215_), .Y(mai_mai_n1414_));
  NO2        m1386(.A(mai_mai_n190_), .B(b), .Y(mai_mai_n1415_));
  AOI220     m1387(.A0(mai_mai_n1177_), .A1(mai_mai_n1415_), .B0(mai_mai_n1102_), .B1(mai_mai_n1405_), .Y(mai_mai_n1416_));
  NAi31      m1388(.An(mai_mai_n1413_), .B(mai_mai_n1416_), .C(mai_mai_n1414_), .Y(mai_mai_n1417_));
  NO4        m1389(.A(mai_mai_n130_), .B(g), .C(f), .D(e), .Y(mai_mai_n1418_));
  NA3        m1390(.A(mai_mai_n1360_), .B(mai_mai_n294_), .C(h), .Y(mai_mai_n1419_));
  NA2        m1391(.A(mai_mai_n197_), .B(mai_mai_n99_), .Y(mai_mai_n1420_));
  OR2        m1392(.A(e), .B(a), .Y(mai_mai_n1421_));
  NO2        m1393(.A(mai_mai_n1352_), .B(mai_mai_n1351_), .Y(mai_mai_n1422_));
  AOI210     m1394(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1422_), .Y(mai_mai_n1423_));
  NO2        m1395(.A(mai_mai_n1423_), .B(mai_mai_n1090_), .Y(mai_mai_n1424_));
  NOi41      m1396(.An(h), .B(f), .C(e), .D(a), .Y(mai_mai_n1425_));
  NA2        m1397(.A(mai_mai_n1425_), .B(mai_mai_n112_), .Y(mai_mai_n1426_));
  NA2        m1398(.A(mai_mai_n1358_), .B(mai_mai_n1380_), .Y(mai_mai_n1427_));
  NA2        m1399(.A(mai_mai_n1427_), .B(mai_mai_n1426_), .Y(mai_mai_n1428_));
  OR3        m1400(.A(mai_mai_n548_), .B(mai_mai_n547_), .C(mai_mai_n111_), .Y(mai_mai_n1429_));
  NA2        m1401(.A(mai_mai_n1119_), .B(mai_mai_n408_), .Y(mai_mai_n1430_));
  OAI220     m1402(.A0(mai_mai_n1430_), .A1(mai_mai_n438_), .B0(mai_mai_n1429_), .B1(mai_mai_n299_), .Y(mai_mai_n1431_));
  AO210      m1403(.A0(mai_mai_n1431_), .A1(mai_mai_n114_), .B0(mai_mai_n1428_), .Y(mai_mai_n1432_));
  NO3        m1404(.A(mai_mai_n1432_), .B(mai_mai_n1424_), .C(mai_mai_n1417_), .Y(mai_mai_n1433_));
  NA4        m1405(.A(mai_mai_n1433_), .B(mai_mai_n1411_), .C(mai_mai_n1383_), .D(mai_mai_n1369_), .Y(mai_mai_n1434_));
  NO2        m1406(.A(mai_mai_n1135_), .B(mai_mai_n109_), .Y(mai_mai_n1435_));
  NA2        m1407(.A(mai_mai_n381_), .B(mai_mai_n56_), .Y(mai_mai_n1436_));
  AOI210     m1408(.A0(mai_mai_n1436_), .A1(mai_mai_n1059_), .B0(mai_mai_n1379_), .Y(mai_mai_n1437_));
  NA2        m1409(.A(mai_mai_n215_), .B(mai_mai_n181_), .Y(mai_mai_n1438_));
  AOI210     m1410(.A0(mai_mai_n1438_), .A1(mai_mai_n1195_), .B0(mai_mai_n1436_), .Y(mai_mai_n1439_));
  NO2        m1411(.A(mai_mai_n1095_), .B(mai_mai_n1090_), .Y(mai_mai_n1440_));
  NO3        m1412(.A(mai_mai_n1440_), .B(mai_mai_n1439_), .C(mai_mai_n1437_), .Y(mai_mai_n1441_));
  NO2        m1413(.A(mai_mai_n393_), .B(j), .Y(mai_mai_n1442_));
  NA3        m1414(.A(mai_mai_n1408_), .B(mai_mai_n1352_), .C(mai_mai_n1119_), .Y(mai_mai_n1443_));
  NAi41      m1415(.An(mai_mai_n1393_), .B(mai_mai_n1081_), .C(mai_mai_n169_), .D(mai_mai_n150_), .Y(mai_mai_n1444_));
  NA2        m1416(.A(mai_mai_n1444_), .B(mai_mai_n1443_), .Y(mai_mai_n1445_));
  NA3        m1417(.A(g), .B(mai_mai_n1442_), .C(mai_mai_n158_), .Y(mai_mai_n1446_));
  INV        m1418(.A(mai_mai_n1446_), .Y(mai_mai_n1447_));
  NO3        m1419(.A(mai_mai_n753_), .B(mai_mai_n176_), .C(mai_mai_n411_), .Y(mai_mai_n1448_));
  NO3        m1420(.A(mai_mai_n1448_), .B(mai_mai_n1447_), .C(mai_mai_n1445_), .Y(mai_mai_n1449_));
  AOI210     m1421(.A0(mai_mai_n1438_), .A1(mai_mai_n1420_), .B0(mai_mai_n1059_), .Y(mai_mai_n1450_));
  OR2        m1422(.A(n), .B(i), .Y(mai_mai_n1451_));
  OAI210     m1423(.A0(mai_mai_n1451_), .A1(mai_mai_n1080_), .B0(mai_mai_n49_), .Y(mai_mai_n1452_));
  AOI220     m1424(.A0(mai_mai_n1452_), .A1(mai_mai_n1185_), .B0(mai_mai_n830_), .B1(mai_mai_n197_), .Y(mai_mai_n1453_));
  INV        m1425(.A(mai_mai_n1453_), .Y(mai_mai_n1454_));
  OAI220     m1426(.A0(mai_mai_n670_), .A1(g), .B0(mai_mai_n225_), .B1(c), .Y(mai_mai_n1455_));
  AOI210     m1427(.A0(mai_mai_n1415_), .A1(mai_mai_n41_), .B0(mai_mai_n1455_), .Y(mai_mai_n1456_));
  NO2        m1428(.A(mai_mai_n130_), .B(l), .Y(mai_mai_n1457_));
  NO2        m1429(.A(mai_mai_n225_), .B(k), .Y(mai_mai_n1458_));
  OAI210     m1430(.A0(mai_mai_n1458_), .A1(mai_mai_n1393_), .B0(mai_mai_n1457_), .Y(mai_mai_n1459_));
  OAI220     m1431(.A0(mai_mai_n1459_), .A1(mai_mai_n31_), .B0(mai_mai_n1456_), .B1(mai_mai_n178_), .Y(mai_mai_n1460_));
  NO3        m1432(.A(mai_mai_n1429_), .B(mai_mai_n472_), .C(mai_mai_n355_), .Y(mai_mai_n1461_));
  NO4        m1433(.A(mai_mai_n1461_), .B(mai_mai_n1460_), .C(mai_mai_n1454_), .D(mai_mai_n1450_), .Y(mai_mai_n1462_));
  NO3        m1434(.A(mai_mai_n1105_), .B(mai_mai_n1352_), .C(mai_mai_n49_), .Y(mai_mai_n1463_));
  NO2        m1435(.A(mai_mai_n1090_), .B(h), .Y(mai_mai_n1464_));
  NA3        m1436(.A(mai_mai_n1464_), .B(d), .C(mai_mai_n1051_), .Y(mai_mai_n1465_));
  NO2        m1437(.A(mai_mai_n1465_), .B(c), .Y(mai_mai_n1466_));
  NA3        m1438(.A(mai_mai_n1435_), .B(mai_mai_n472_), .C(f), .Y(mai_mai_n1467_));
  NA2        m1439(.A(mai_mai_n181_), .B(mai_mai_n111_), .Y(mai_mai_n1468_));
  NO2        m1440(.A(mai_mai_n42_), .B(mai_mai_n1467_), .Y(mai_mai_n1469_));
  NO2        m1441(.A(mai_mai_n1342_), .B(mai_mai_n176_), .Y(mai_mai_n1470_));
  NOi21      m1442(.An(d), .B(f), .Y(mai_mai_n1471_));
  NO3        m1443(.A(mai_mai_n1401_), .B(mai_mai_n1471_), .C(mai_mai_n40_), .Y(mai_mai_n1472_));
  NA2        m1444(.A(mai_mai_n1472_), .B(mai_mai_n1470_), .Y(mai_mai_n1473_));
  NO2        m1445(.A(mai_mai_n1352_), .B(f), .Y(mai_mai_n1474_));
  INV        m1446(.A(mai_mai_n1473_), .Y(mai_mai_n1475_));
  NO3        m1447(.A(mai_mai_n1475_), .B(mai_mai_n1469_), .C(mai_mai_n1466_), .Y(mai_mai_n1476_));
  NA4        m1448(.A(mai_mai_n1476_), .B(mai_mai_n1462_), .C(mai_mai_n1449_), .D(mai_mai_n1441_), .Y(mai_mai_n1477_));
  NO3        m1449(.A(mai_mai_n1094_), .B(mai_mai_n1080_), .C(mai_mai_n40_), .Y(mai_mai_n1478_));
  NO2        m1450(.A(mai_mai_n472_), .B(mai_mai_n299_), .Y(mai_mai_n1479_));
  OAI210     m1451(.A0(mai_mai_n1479_), .A1(mai_mai_n1478_), .B0(mai_mai_n1365_), .Y(mai_mai_n1480_));
  OAI210     m1452(.A0(mai_mai_n1418_), .A1(mai_mai_n1355_), .B0(mai_mai_n889_), .Y(mai_mai_n1481_));
  NO2        m1453(.A(mai_mai_n1047_), .B(mai_mai_n130_), .Y(mai_mai_n1482_));
  NA2        m1454(.A(mai_mai_n1482_), .B(mai_mai_n626_), .Y(mai_mai_n1483_));
  NA3        m1455(.A(mai_mai_n1483_), .B(mai_mai_n1481_), .C(mai_mai_n1480_), .Y(mai_mai_n1484_));
  NA2        m1456(.A(mai_mai_n1386_), .B(mai_mai_n1471_), .Y(mai_mai_n1485_));
  NO2        m1457(.A(mai_mai_n1485_), .B(m), .Y(mai_mai_n1486_));
  NO2        m1458(.A(mai_mai_n151_), .B(mai_mai_n183_), .Y(mai_mai_n1487_));
  OAI210     m1459(.A0(mai_mai_n1487_), .A1(mai_mai_n109_), .B0(mai_mai_n1400_), .Y(mai_mai_n1488_));
  INV        m1460(.A(mai_mai_n1488_), .Y(mai_mai_n1489_));
  NO3        m1461(.A(mai_mai_n1489_), .B(mai_mai_n1486_), .C(mai_mai_n1484_), .Y(mai_mai_n1490_));
  NO2        m1462(.A(mai_mai_n1351_), .B(e), .Y(mai_mai_n1491_));
  NA2        m1463(.A(mai_mai_n1491_), .B(mai_mai_n406_), .Y(mai_mai_n1492_));
  OAI210     m1464(.A0(mai_mai_n1474_), .A1(mai_mai_n1130_), .B0(mai_mai_n635_), .Y(mai_mai_n1493_));
  OR3        m1465(.A(mai_mai_n1458_), .B(mai_mai_n1219_), .C(mai_mai_n130_), .Y(mai_mai_n1494_));
  OAI220     m1466(.A0(mai_mai_n1494_), .A1(mai_mai_n1492_), .B0(mai_mai_n1493_), .B1(mai_mai_n447_), .Y(mai_mai_n1495_));
  INV        m1467(.A(mai_mai_n1495_), .Y(mai_mai_n1496_));
  NO2        m1468(.A(mai_mai_n183_), .B(c), .Y(mai_mai_n1497_));
  OAI210     m1469(.A0(mai_mai_n1497_), .A1(mai_mai_n1491_), .B0(mai_mai_n181_), .Y(mai_mai_n1498_));
  AOI220     m1470(.A0(mai_mai_n1498_), .A1(mai_mai_n1082_), .B0(mai_mai_n540_), .B1(mai_mai_n370_), .Y(mai_mai_n1499_));
  NA2        m1471(.A(mai_mai_n547_), .B(g), .Y(mai_mai_n1500_));
  AOI210     m1472(.A0(mai_mai_n1500_), .A1(mai_mai_n1382_), .B0(mai_mai_n1463_), .Y(mai_mai_n1501_));
  NO2        m1473(.A(mai_mai_n1421_), .B(f), .Y(mai_mai_n1502_));
  NA2        m1474(.A(mai_mai_n1130_), .B(a), .Y(mai_mai_n1503_));
  OAI220     m1475(.A0(mai_mai_n1503_), .A1(mai_mai_n69_), .B0(mai_mai_n1501_), .B1(mai_mai_n213_), .Y(mai_mai_n1504_));
  AOI210     m1476(.A0(mai_mai_n908_), .A1(mai_mai_n418_), .B0(mai_mai_n104_), .Y(mai_mai_n1505_));
  OR2        m1477(.A(mai_mai_n1505_), .B(mai_mai_n547_), .Y(mai_mai_n1506_));
  NA2        m1478(.A(mai_mai_n1502_), .B(mai_mai_n1362_), .Y(mai_mai_n1507_));
  OAI220     m1479(.A0(mai_mai_n1507_), .A1(mai_mai_n49_), .B0(mai_mai_n1506_), .B1(mai_mai_n176_), .Y(mai_mai_n1508_));
  NA4        m1480(.A(mai_mai_n1103_), .B(mai_mai_n1100_), .C(mai_mai_n221_), .D(mai_mai_n68_), .Y(mai_mai_n1509_));
  NA2        m1481(.A(mai_mai_n1356_), .B(mai_mai_n184_), .Y(mai_mai_n1510_));
  NO2        m1482(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1511_));
  OAI210     m1483(.A0(mai_mai_n1421_), .A1(mai_mai_n867_), .B0(mai_mai_n491_), .Y(mai_mai_n1512_));
  OAI210     m1484(.A0(mai_mai_n1512_), .A1(mai_mai_n1106_), .B0(mai_mai_n1511_), .Y(mai_mai_n1513_));
  NO2        m1485(.A(mai_mai_n252_), .B(g), .Y(mai_mai_n1514_));
  NO2        m1486(.A(m), .B(i), .Y(mai_mai_n1515_));
  BUFFER     m1487(.A(mai_mai_n1515_), .Y(mai_mai_n1516_));
  AOI220     m1488(.A0(mai_mai_n1516_), .A1(mai_mai_n1384_), .B0(mai_mai_n1081_), .B1(mai_mai_n1514_), .Y(mai_mai_n1517_));
  NA4        m1489(.A(mai_mai_n1517_), .B(mai_mai_n1513_), .C(mai_mai_n1510_), .D(mai_mai_n1509_), .Y(mai_mai_n1518_));
  NO4        m1490(.A(mai_mai_n1518_), .B(mai_mai_n1508_), .C(mai_mai_n1504_), .D(mai_mai_n1499_), .Y(mai_mai_n1519_));
  NA3        m1491(.A(mai_mai_n1519_), .B(mai_mai_n1496_), .C(mai_mai_n1490_), .Y(mai_mai_n1520_));
  NA3        m1492(.A(mai_mai_n966_), .B(mai_mai_n137_), .C(mai_mai_n46_), .Y(mai_mai_n1521_));
  AOI210     m1493(.A0(mai_mai_n148_), .A1(c), .B0(mai_mai_n1521_), .Y(mai_mai_n1522_));
  INV        m1494(.A(mai_mai_n187_), .Y(mai_mai_n1523_));
  NA2        m1495(.A(mai_mai_n1523_), .B(mai_mai_n1464_), .Y(mai_mai_n1524_));
  OR2        m1496(.A(mai_mai_n131_), .B(mai_mai_n1412_), .Y(mai_mai_n1525_));
  NO2        m1497(.A(mai_mai_n72_), .B(c), .Y(mai_mai_n1526_));
  NA2        m1498(.A(mai_mai_n1470_), .B(mai_mai_n1526_), .Y(mai_mai_n1527_));
  NA3        m1499(.A(mai_mai_n1527_), .B(mai_mai_n1525_), .C(mai_mai_n1524_), .Y(mai_mai_n1528_));
  NO2        m1500(.A(mai_mai_n1528_), .B(mai_mai_n1522_), .Y(mai_mai_n1529_));
  AOI210     m1501(.A0(mai_mai_n156_), .A1(mai_mai_n56_), .B0(mai_mai_n1491_), .Y(mai_mai_n1530_));
  NO2        m1502(.A(mai_mai_n1530_), .B(mai_mai_n1468_), .Y(mai_mai_n1531_));
  NOi21      m1503(.An(mai_mai_n1356_), .B(e), .Y(mai_mai_n1532_));
  NO2        m1504(.A(mai_mai_n1532_), .B(mai_mai_n1531_), .Y(mai_mai_n1533_));
  AN2        m1505(.A(mai_mai_n1103_), .B(mai_mai_n1088_), .Y(mai_mai_n1534_));
  AOI220     m1506(.A0(mai_mai_n1515_), .A1(mai_mai_n643_), .B0(mai_mai_n1065_), .B1(mai_mai_n159_), .Y(mai_mai_n1535_));
  NOi31      m1507(.An(mai_mai_n30_), .B(mai_mai_n1535_), .C(n), .Y(mai_mai_n1536_));
  AOI210     m1508(.A0(mai_mai_n1534_), .A1(mai_mai_n1177_), .B0(mai_mai_n1536_), .Y(mai_mai_n1537_));
  NO2        m1509(.A(mai_mai_n1467_), .B(mai_mai_n69_), .Y(mai_mai_n1538_));
  NA2        m1510(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1539_));
  NO2        m1511(.A(mai_mai_n1360_), .B(mai_mai_n116_), .Y(mai_mai_n1540_));
  OAI220     m1512(.A0(mai_mai_n1540_), .A1(mai_mai_n1412_), .B0(mai_mai_n1430_), .B1(mai_mai_n1539_), .Y(mai_mai_n1541_));
  NO2        m1513(.A(mai_mai_n1541_), .B(mai_mai_n1538_), .Y(mai_mai_n1542_));
  NA4        m1514(.A(mai_mai_n1542_), .B(mai_mai_n1537_), .C(mai_mai_n1533_), .D(mai_mai_n1529_), .Y(mai_mai_n1543_));
  OR4        m1515(.A(mai_mai_n1543_), .B(mai_mai_n1520_), .C(mai_mai_n1477_), .D(mai_mai_n1434_), .Y(mai04));
  NOi31      m1516(.An(mai_mai_n1418_), .B(mai_mai_n1419_), .C(mai_mai_n1053_), .Y(mai_mai_n1545_));
  NA2        m1517(.A(mai_mai_n1474_), .B(mai_mai_n830_), .Y(mai_mai_n1546_));
  NO4        m1518(.A(mai_mai_n1546_), .B(mai_mai_n1042_), .C(mai_mai_n492_), .D(j), .Y(mai_mai_n1547_));
  OR3        m1519(.A(mai_mai_n1547_), .B(mai_mai_n1545_), .C(mai_mai_n1071_), .Y(mai_mai_n1548_));
  NO2        m1520(.A(mai_mai_n1362_), .B(mai_mai_n92_), .Y(mai_mai_n1549_));
  AOI210     m1521(.A0(mai_mai_n1549_), .A1(mai_mai_n1064_), .B0(mai_mai_n1197_), .Y(mai_mai_n1550_));
  NA2        m1522(.A(mai_mai_n1550_), .B(mai_mai_n1223_), .Y(mai_mai_n1551_));
  NO4        m1523(.A(mai_mai_n1551_), .B(mai_mai_n1548_), .C(mai_mai_n1079_), .D(mai_mai_n1058_), .Y(mai_mai_n1552_));
  NA4        m1524(.A(mai_mai_n1552_), .B(mai_mai_n1132_), .C(mai_mai_n1117_), .D(mai_mai_n1109_), .Y(mai05));
  INV        m1525(.A(m), .Y(mai_mai_n1556_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  INV        u0023(.A(men_men_n51_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(g), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(g), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(g), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(g), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(g), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n96_), .C(f), .Y(men_men_n98_));
  AN2        u0070(.A(j), .B(g), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(l), .C(i), .Y(men_men_n100_));
  NOi21      u0072(.An(g), .B(i), .Y(men_men_n101_));
  NOi32      u0073(.An(m), .Bn(j), .C(k), .Y(men_men_n102_));
  AOI220     u0074(.A0(men_men_n102_), .A1(men_men_n101_), .B0(men_men_n100_), .B1(men_men_n99_), .Y(men_men_n103_));
  NO2        u0075(.A(men_men_n103_), .B(f), .Y(men_men_n104_));
  NO3        u0076(.A(men_men_n104_), .B(men_men_n98_), .C(men_men_n95_), .Y(men_men_n105_));
  NAi41      u0077(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n106_));
  AN2        u0078(.A(e), .B(b), .Y(men_men_n107_));
  NOi31      u0079(.An(c), .B(h), .C(f), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NO2        u0081(.A(men_men_n109_), .B(men_men_n106_), .Y(men_men_n110_));
  NOi21      u0082(.An(g), .B(f), .Y(men_men_n111_));
  NOi21      u0083(.An(i), .B(h), .Y(men_men_n112_));
  NA3        u0084(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n36_), .Y(men_men_n113_));
  INV        u0085(.A(a), .Y(men_men_n114_));
  NA2        u0086(.A(men_men_n107_), .B(men_men_n114_), .Y(men_men_n115_));
  INV        u0087(.A(l), .Y(men_men_n116_));
  NOi21      u0088(.An(m), .B(n), .Y(men_men_n117_));
  AN2        u0089(.A(k), .B(h), .Y(men_men_n118_));
  NO2        u0090(.A(men_men_n113_), .B(men_men_n88_), .Y(men_men_n119_));
  INV        u0091(.A(b), .Y(men_men_n120_));
  NA2        u0092(.A(l), .B(j), .Y(men_men_n121_));
  AN2        u0093(.A(k), .B(i), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n121_), .Y(men_men_n123_));
  NA2        u0095(.A(g), .B(e), .Y(men_men_n124_));
  NOi32      u0096(.An(c), .Bn(a), .C(d), .Y(men_men_n125_));
  NA2        u0097(.A(men_men_n125_), .B(men_men_n117_), .Y(men_men_n126_));
  NO4        u0098(.A(men_men_n126_), .B(men_men_n124_), .C(men_men_n123_), .D(men_men_n120_), .Y(men_men_n127_));
  NO3        u0099(.A(men_men_n127_), .B(men_men_n119_), .C(men_men_n110_), .Y(men_men_n128_));
  OAI210     u0100(.A0(men_men_n105_), .A1(men_men_n88_), .B0(men_men_n128_), .Y(men_men_n129_));
  NOi31      u0101(.An(k), .B(m), .C(j), .Y(men_men_n130_));
  NA3        u0102(.A(men_men_n130_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n131_));
  NOi31      u0103(.An(k), .B(m), .C(i), .Y(men_men_n132_));
  NA3        u0104(.A(men_men_n132_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n133_));
  NA2        u0105(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n134_));
  NOi32      u0106(.An(f), .Bn(b), .C(e), .Y(men_men_n135_));
  NAi21      u0107(.An(g), .B(h), .Y(men_men_n136_));
  NAi21      u0108(.An(m), .B(n), .Y(men_men_n137_));
  NAi21      u0109(.An(j), .B(k), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n139_));
  NAi41      u0111(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n140_));
  NAi31      u0112(.An(j), .B(k), .C(h), .Y(men_men_n141_));
  NO3        u0113(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n137_), .Y(men_men_n142_));
  AOI210     u0114(.A0(men_men_n139_), .A1(men_men_n135_), .B0(men_men_n142_), .Y(men_men_n143_));
  NO2        u0115(.A(k), .B(j), .Y(men_men_n144_));
  AN2        u0116(.A(k), .B(j), .Y(men_men_n145_));
  NAi21      u0117(.An(c), .B(b), .Y(men_men_n146_));
  NA2        u0118(.A(f), .B(d), .Y(men_men_n147_));
  NA2        u0119(.A(h), .B(c), .Y(men_men_n148_));
  NAi31      u0120(.An(f), .B(e), .C(b), .Y(men_men_n149_));
  NA2        u0121(.A(d), .B(b), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(f), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n151_), .B(men_men_n150_), .Y(men_men_n152_));
  NA2        u0124(.A(b), .B(a), .Y(men_men_n153_));
  NAi21      u0125(.An(e), .B(g), .Y(men_men_n154_));
  NAi21      u0126(.An(c), .B(d), .Y(men_men_n155_));
  NAi31      u0127(.An(l), .B(k), .C(h), .Y(men_men_n156_));
  NO2        u0128(.A(men_men_n137_), .B(men_men_n156_), .Y(men_men_n157_));
  NA2        u0129(.A(men_men_n157_), .B(men_men_n152_), .Y(men_men_n158_));
  NAi31      u0130(.An(men_men_n134_), .B(men_men_n158_), .C(men_men_n143_), .Y(men_men_n159_));
  NAi31      u0131(.An(e), .B(f), .C(b), .Y(men_men_n160_));
  NOi21      u0132(.An(g), .B(d), .Y(men_men_n161_));
  NO2        u0133(.A(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  NOi21      u0134(.An(h), .B(i), .Y(men_men_n163_));
  NOi21      u0135(.An(k), .B(m), .Y(men_men_n164_));
  NA3        u0136(.A(men_men_n164_), .B(men_men_n163_), .C(n), .Y(men_men_n165_));
  NOi21      u0137(.An(men_men_n162_), .B(men_men_n165_), .Y(men_men_n166_));
  NOi21      u0138(.An(h), .B(g), .Y(men_men_n167_));
  NO2        u0139(.A(men_men_n147_), .B(men_men_n146_), .Y(men_men_n168_));
  NA2        u0140(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  NAi31      u0141(.An(l), .B(j), .C(h), .Y(men_men_n170_));
  NO2        u0142(.A(men_men_n170_), .B(men_men_n49_), .Y(men_men_n171_));
  NA2        u0143(.A(men_men_n171_), .B(men_men_n67_), .Y(men_men_n172_));
  NOi32      u0144(.An(n), .Bn(k), .C(m), .Y(men_men_n173_));
  NA2        u0145(.A(l), .B(i), .Y(men_men_n174_));
  INV        u0146(.A(men_men_n173_), .Y(men_men_n175_));
  OAI210     u0147(.A0(men_men_n175_), .A1(men_men_n169_), .B0(men_men_n172_), .Y(men_men_n176_));
  NAi31      u0148(.An(d), .B(f), .C(c), .Y(men_men_n177_));
  NAi31      u0149(.An(e), .B(f), .C(c), .Y(men_men_n178_));
  NA2        u0150(.A(men_men_n178_), .B(men_men_n177_), .Y(men_men_n179_));
  NA2        u0151(.A(j), .B(h), .Y(men_men_n180_));
  OR3        u0152(.A(n), .B(m), .C(k), .Y(men_men_n181_));
  NO2        u0153(.A(men_men_n181_), .B(men_men_n180_), .Y(men_men_n182_));
  NAi32      u0154(.An(m), .Bn(k), .C(n), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n183_), .B(men_men_n180_), .Y(men_men_n184_));
  AOI220     u0156(.A0(men_men_n184_), .A1(men_men_n162_), .B0(men_men_n182_), .B1(men_men_n179_), .Y(men_men_n185_));
  NO2        u0157(.A(n), .B(m), .Y(men_men_n186_));
  NA2        u0158(.A(men_men_n186_), .B(men_men_n50_), .Y(men_men_n187_));
  NAi21      u0159(.An(f), .B(e), .Y(men_men_n188_));
  NA2        u0160(.A(d), .B(c), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NOi21      u0162(.An(men_men_n190_), .B(men_men_n187_), .Y(men_men_n191_));
  NAi21      u0163(.An(d), .B(c), .Y(men_men_n192_));
  NAi31      u0164(.An(m), .B(n), .C(b), .Y(men_men_n193_));
  NA2        u0165(.A(k), .B(i), .Y(men_men_n194_));
  NAi21      u0166(.An(h), .B(f), .Y(men_men_n195_));
  NO2        u0167(.A(men_men_n195_), .B(men_men_n194_), .Y(men_men_n196_));
  NO2        u0168(.A(men_men_n193_), .B(men_men_n155_), .Y(men_men_n197_));
  NA2        u0169(.A(men_men_n197_), .B(men_men_n196_), .Y(men_men_n198_));
  NOi32      u0170(.An(f), .Bn(c), .C(d), .Y(men_men_n199_));
  NOi32      u0171(.An(f), .Bn(c), .C(e), .Y(men_men_n200_));
  NO2        u0172(.A(men_men_n200_), .B(men_men_n199_), .Y(men_men_n201_));
  NO3        u0173(.A(n), .B(m), .C(j), .Y(men_men_n202_));
  NA2        u0174(.A(men_men_n202_), .B(men_men_n118_), .Y(men_men_n203_));
  AO210      u0175(.A0(men_men_n203_), .A1(men_men_n187_), .B0(men_men_n201_), .Y(men_men_n204_));
  NAi41      u0176(.An(men_men_n191_), .B(men_men_n204_), .C(men_men_n198_), .D(men_men_n185_), .Y(men_men_n205_));
  OR4        u0177(.A(men_men_n205_), .B(men_men_n176_), .C(men_men_n166_), .D(men_men_n159_), .Y(men_men_n206_));
  NO4        u0178(.A(men_men_n206_), .B(men_men_n129_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n207_));
  NA3        u0179(.A(m), .B(men_men_n116_), .C(j), .Y(men_men_n208_));
  NAi31      u0180(.An(n), .B(h), .C(g), .Y(men_men_n209_));
  NO2        u0181(.A(men_men_n209_), .B(men_men_n208_), .Y(men_men_n210_));
  NOi32      u0182(.An(m), .Bn(k), .C(l), .Y(men_men_n211_));
  NA3        u0183(.A(men_men_n211_), .B(men_men_n89_), .C(g), .Y(men_men_n212_));
  NO2        u0184(.A(men_men_n212_), .B(n), .Y(men_men_n213_));
  NOi21      u0185(.An(k), .B(j), .Y(men_men_n214_));
  NA4        u0186(.A(men_men_n214_), .B(men_men_n117_), .C(i), .D(g), .Y(men_men_n215_));
  AN2        u0187(.A(i), .B(g), .Y(men_men_n216_));
  NA3        u0188(.A(men_men_n76_), .B(men_men_n216_), .C(men_men_n117_), .Y(men_men_n217_));
  NA2        u0189(.A(men_men_n217_), .B(men_men_n215_), .Y(men_men_n218_));
  NO3        u0190(.A(men_men_n218_), .B(men_men_n213_), .C(men_men_n210_), .Y(men_men_n219_));
  NAi41      u0191(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n220_));
  INV        u0192(.A(men_men_n220_), .Y(men_men_n221_));
  INV        u0193(.A(f), .Y(men_men_n222_));
  INV        u0194(.A(g), .Y(men_men_n223_));
  NOi31      u0195(.An(i), .B(j), .C(h), .Y(men_men_n224_));
  NOi21      u0196(.An(l), .B(m), .Y(men_men_n225_));
  NA2        u0197(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  NO3        u0198(.A(men_men_n226_), .B(men_men_n223_), .C(men_men_n222_), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n227_), .B(men_men_n221_), .Y(men_men_n228_));
  OAI210     u0200(.A0(men_men_n219_), .A1(men_men_n32_), .B0(men_men_n228_), .Y(men_men_n229_));
  NOi21      u0201(.An(n), .B(m), .Y(men_men_n230_));
  NOi32      u0202(.An(l), .Bn(i), .C(j), .Y(men_men_n231_));
  NA2        u0203(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  OA220      u0204(.A0(men_men_n232_), .A1(men_men_n109_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n233_));
  NAi21      u0205(.An(j), .B(h), .Y(men_men_n234_));
  XN2        u0206(.A(i), .B(h), .Y(men_men_n235_));
  NA2        u0207(.A(men_men_n235_), .B(men_men_n234_), .Y(men_men_n236_));
  NOi31      u0208(.An(k), .B(n), .C(m), .Y(men_men_n237_));
  NOi31      u0209(.An(men_men_n237_), .B(men_men_n189_), .C(men_men_n188_), .Y(men_men_n238_));
  NA2        u0210(.A(men_men_n238_), .B(men_men_n236_), .Y(men_men_n239_));
  NAi31      u0211(.An(f), .B(e), .C(c), .Y(men_men_n240_));
  NO4        u0212(.A(men_men_n240_), .B(men_men_n181_), .C(men_men_n180_), .D(men_men_n59_), .Y(men_men_n241_));
  NA4        u0213(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n242_));
  NAi32      u0214(.An(m), .Bn(i), .C(k), .Y(men_men_n243_));
  NO3        u0215(.A(men_men_n243_), .B(men_men_n93_), .C(men_men_n242_), .Y(men_men_n244_));
  INV        u0216(.A(k), .Y(men_men_n245_));
  NO2        u0217(.A(men_men_n244_), .B(men_men_n241_), .Y(men_men_n246_));
  NAi21      u0218(.An(n), .B(a), .Y(men_men_n247_));
  NO2        u0219(.A(men_men_n247_), .B(men_men_n150_), .Y(men_men_n248_));
  NAi41      u0220(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(e), .Y(men_men_n250_));
  NO3        u0222(.A(men_men_n151_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n251_));
  OAI210     u0223(.A0(men_men_n251_), .A1(men_men_n250_), .B0(men_men_n248_), .Y(men_men_n252_));
  AN4        u0224(.A(men_men_n252_), .B(men_men_n246_), .C(men_men_n239_), .D(men_men_n233_), .Y(men_men_n253_));
  OR2        u0225(.A(h), .B(g), .Y(men_men_n254_));
  NO2        u0226(.A(men_men_n254_), .B(men_men_n106_), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n255_), .B(men_men_n135_), .Y(men_men_n256_));
  NAi41      u0228(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n257_), .B(men_men_n222_), .Y(men_men_n258_));
  NA2        u0230(.A(men_men_n164_), .B(men_men_n112_), .Y(men_men_n259_));
  NAi21      u0231(.An(men_men_n259_), .B(men_men_n258_), .Y(men_men_n260_));
  NO2        u0232(.A(n), .B(a), .Y(men_men_n261_));
  NAi31      u0233(.An(men_men_n249_), .B(men_men_n261_), .C(men_men_n107_), .Y(men_men_n262_));
  AN2        u0234(.A(men_men_n262_), .B(men_men_n260_), .Y(men_men_n263_));
  NAi21      u0235(.An(h), .B(i), .Y(men_men_n264_));
  NA2        u0236(.A(men_men_n186_), .B(k), .Y(men_men_n265_));
  NO2        u0237(.A(men_men_n265_), .B(men_men_n264_), .Y(men_men_n266_));
  NA2        u0238(.A(men_men_n266_), .B(men_men_n199_), .Y(men_men_n267_));
  NA3        u0239(.A(men_men_n267_), .B(men_men_n263_), .C(men_men_n256_), .Y(men_men_n268_));
  NOi21      u0240(.An(g), .B(e), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n270_));
  NA2        u0242(.A(men_men_n270_), .B(men_men_n269_), .Y(men_men_n271_));
  NOi32      u0243(.An(l), .Bn(j), .C(i), .Y(men_men_n272_));
  AOI210     u0244(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n272_), .Y(men_men_n273_));
  NO2        u0245(.A(men_men_n264_), .B(men_men_n44_), .Y(men_men_n274_));
  NAi21      u0246(.An(f), .B(g), .Y(men_men_n275_));
  NO2        u0247(.A(men_men_n275_), .B(men_men_n65_), .Y(men_men_n276_));
  NO2        u0248(.A(men_men_n69_), .B(men_men_n121_), .Y(men_men_n277_));
  AOI220     u0249(.A0(men_men_n277_), .A1(men_men_n276_), .B0(men_men_n274_), .B1(men_men_n67_), .Y(men_men_n278_));
  OAI210     u0250(.A0(men_men_n273_), .A1(men_men_n271_), .B0(men_men_n278_), .Y(men_men_n279_));
  NO3        u0251(.A(men_men_n138_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n280_));
  NOi41      u0252(.An(men_men_n253_), .B(men_men_n279_), .C(men_men_n268_), .D(men_men_n229_), .Y(men_men_n281_));
  NO4        u0253(.A(men_men_n210_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n282_));
  NO2        u0254(.A(men_men_n282_), .B(men_men_n115_), .Y(men_men_n283_));
  NA3        u0255(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n284_));
  NAi21      u0256(.An(h), .B(g), .Y(men_men_n285_));
  OR4        u0257(.A(men_men_n285_), .B(men_men_n284_), .C(men_men_n232_), .D(e), .Y(men_men_n286_));
  NAi31      u0258(.An(g), .B(k), .C(h), .Y(men_men_n287_));
  NO3        u0259(.A(men_men_n137_), .B(men_men_n287_), .C(l), .Y(men_men_n288_));
  NAi31      u0260(.An(e), .B(d), .C(a), .Y(men_men_n289_));
  NA2        u0261(.A(men_men_n288_), .B(men_men_n135_), .Y(men_men_n290_));
  NA2        u0262(.A(men_men_n290_), .B(men_men_n286_), .Y(men_men_n291_));
  NA3        u0263(.A(men_men_n164_), .B(men_men_n163_), .C(men_men_n86_), .Y(men_men_n292_));
  NO2        u0264(.A(men_men_n292_), .B(men_men_n201_), .Y(men_men_n293_));
  INV        u0265(.A(men_men_n293_), .Y(men_men_n294_));
  NA3        u0266(.A(e), .B(c), .C(b), .Y(men_men_n295_));
  NO2        u0267(.A(men_men_n60_), .B(men_men_n295_), .Y(men_men_n296_));
  NAi32      u0268(.An(k), .Bn(i), .C(j), .Y(men_men_n297_));
  NAi31      u0269(.An(h), .B(l), .C(i), .Y(men_men_n298_));
  NA3        u0270(.A(men_men_n298_), .B(men_men_n297_), .C(men_men_n170_), .Y(men_men_n299_));
  NOi21      u0271(.An(men_men_n299_), .B(men_men_n49_), .Y(men_men_n300_));
  OAI210     u0272(.A0(men_men_n276_), .A1(men_men_n296_), .B0(men_men_n300_), .Y(men_men_n301_));
  NAi21      u0273(.An(l), .B(k), .Y(men_men_n302_));
  NO2        u0274(.A(men_men_n302_), .B(men_men_n49_), .Y(men_men_n303_));
  NOi21      u0275(.An(l), .B(j), .Y(men_men_n304_));
  NA2        u0276(.A(men_men_n167_), .B(men_men_n304_), .Y(men_men_n305_));
  NA3        u0277(.A(men_men_n122_), .B(men_men_n121_), .C(g), .Y(men_men_n306_));
  OR3        u0278(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n307_));
  AOI210     u0279(.A0(men_men_n306_), .A1(men_men_n305_), .B0(men_men_n307_), .Y(men_men_n308_));
  INV        u0280(.A(men_men_n308_), .Y(men_men_n309_));
  NAi32      u0281(.An(j), .Bn(h), .C(i), .Y(men_men_n310_));
  NAi21      u0282(.An(m), .B(l), .Y(men_men_n311_));
  NO3        u0283(.A(men_men_n311_), .B(men_men_n310_), .C(men_men_n86_), .Y(men_men_n312_));
  NA2        u0284(.A(h), .B(g), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n173_), .B(men_men_n45_), .Y(men_men_n314_));
  NO2        u0286(.A(men_men_n314_), .B(men_men_n313_), .Y(men_men_n315_));
  OAI210     u0287(.A0(men_men_n315_), .A1(men_men_n312_), .B0(men_men_n168_), .Y(men_men_n316_));
  NA4        u0288(.A(men_men_n316_), .B(men_men_n309_), .C(men_men_n301_), .D(men_men_n294_), .Y(men_men_n317_));
  NO2        u0289(.A(men_men_n149_), .B(d), .Y(men_men_n318_));
  NA2        u0290(.A(men_men_n318_), .B(men_men_n53_), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n109_), .B(men_men_n106_), .Y(men_men_n320_));
  NAi32      u0292(.An(n), .Bn(m), .C(l), .Y(men_men_n321_));
  NO2        u0293(.A(men_men_n321_), .B(men_men_n310_), .Y(men_men_n322_));
  NA2        u0294(.A(men_men_n322_), .B(men_men_n190_), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n126_), .B(men_men_n120_), .Y(men_men_n324_));
  NAi31      u0296(.An(k), .B(l), .C(j), .Y(men_men_n325_));
  OAI210     u0297(.A0(men_men_n302_), .A1(j), .B0(men_men_n325_), .Y(men_men_n326_));
  NOi21      u0298(.An(men_men_n326_), .B(men_men_n124_), .Y(men_men_n327_));
  NA2        u0299(.A(men_men_n327_), .B(men_men_n324_), .Y(men_men_n328_));
  NA3        u0300(.A(men_men_n328_), .B(men_men_n323_), .C(men_men_n319_), .Y(men_men_n329_));
  NO4        u0301(.A(men_men_n329_), .B(men_men_n317_), .C(men_men_n291_), .D(men_men_n283_), .Y(men_men_n330_));
  NA2        u0302(.A(men_men_n266_), .B(men_men_n200_), .Y(men_men_n331_));
  NAi21      u0303(.An(m), .B(k), .Y(men_men_n332_));
  NO2        u0304(.A(men_men_n235_), .B(men_men_n332_), .Y(men_men_n333_));
  NAi41      u0305(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n334_));
  NO2        u0306(.A(men_men_n334_), .B(men_men_n154_), .Y(men_men_n335_));
  NA2        u0307(.A(men_men_n335_), .B(men_men_n333_), .Y(men_men_n336_));
  NAi31      u0308(.An(i), .B(l), .C(h), .Y(men_men_n337_));
  NO4        u0309(.A(men_men_n337_), .B(men_men_n154_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n338_));
  NA2        u0310(.A(e), .B(c), .Y(men_men_n339_));
  NO3        u0311(.A(men_men_n339_), .B(n), .C(d), .Y(men_men_n340_));
  NOi21      u0312(.An(f), .B(h), .Y(men_men_n341_));
  NA2        u0313(.A(men_men_n341_), .B(men_men_n122_), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n342_), .B(men_men_n223_), .Y(men_men_n343_));
  NAi31      u0315(.An(d), .B(e), .C(b), .Y(men_men_n344_));
  NO2        u0316(.A(men_men_n137_), .B(men_men_n344_), .Y(men_men_n345_));
  NA2        u0317(.A(men_men_n345_), .B(men_men_n343_), .Y(men_men_n346_));
  NAi41      u0318(.An(men_men_n338_), .B(men_men_n346_), .C(men_men_n336_), .D(men_men_n331_), .Y(men_men_n347_));
  NO4        u0319(.A(men_men_n334_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n223_), .Y(men_men_n348_));
  NA2        u0320(.A(men_men_n261_), .B(men_men_n107_), .Y(men_men_n349_));
  OR2        u0321(.A(men_men_n349_), .B(men_men_n212_), .Y(men_men_n350_));
  NOi31      u0322(.An(l), .B(n), .C(m), .Y(men_men_n351_));
  NA2        u0323(.A(men_men_n351_), .B(men_men_n224_), .Y(men_men_n352_));
  NO2        u0324(.A(men_men_n352_), .B(men_men_n201_), .Y(men_men_n353_));
  NAi32      u0325(.An(men_men_n353_), .Bn(men_men_n348_), .C(men_men_n350_), .Y(men_men_n354_));
  NAi32      u0326(.An(m), .Bn(j), .C(k), .Y(men_men_n355_));
  NAi41      u0327(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n356_));
  OAI210     u0328(.A0(men_men_n220_), .A1(men_men_n355_), .B0(men_men_n356_), .Y(men_men_n357_));
  NOi31      u0329(.An(j), .B(m), .C(k), .Y(men_men_n358_));
  NO2        u0330(.A(men_men_n130_), .B(men_men_n358_), .Y(men_men_n359_));
  AN3        u0331(.A(h), .B(g), .C(f), .Y(men_men_n360_));
  NAi31      u0332(.An(men_men_n359_), .B(men_men_n360_), .C(men_men_n357_), .Y(men_men_n361_));
  NOi32      u0333(.An(m), .Bn(j), .C(l), .Y(men_men_n362_));
  NO2        u0334(.A(men_men_n362_), .B(men_men_n100_), .Y(men_men_n363_));
  NAi32      u0335(.An(men_men_n363_), .Bn(men_men_n209_), .C(men_men_n318_), .Y(men_men_n364_));
  NO2        u0336(.A(men_men_n311_), .B(men_men_n310_), .Y(men_men_n365_));
  NO2        u0337(.A(men_men_n226_), .B(g), .Y(men_men_n366_));
  NO2        u0338(.A(men_men_n160_), .B(men_men_n86_), .Y(men_men_n367_));
  AOI220     u0339(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n258_), .B1(men_men_n365_), .Y(men_men_n368_));
  NA2        u0340(.A(men_men_n243_), .B(men_men_n81_), .Y(men_men_n369_));
  NA3        u0341(.A(men_men_n369_), .B(men_men_n360_), .C(men_men_n221_), .Y(men_men_n370_));
  NA4        u0342(.A(men_men_n370_), .B(men_men_n368_), .C(men_men_n364_), .D(men_men_n361_), .Y(men_men_n371_));
  NA3        u0343(.A(h), .B(g), .C(f), .Y(men_men_n372_));
  NO2        u0344(.A(men_men_n372_), .B(men_men_n77_), .Y(men_men_n373_));
  INV        u0345(.A(men_men_n220_), .Y(men_men_n374_));
  NA2        u0346(.A(men_men_n167_), .B(e), .Y(men_men_n375_));
  NO2        u0347(.A(men_men_n375_), .B(men_men_n41_), .Y(men_men_n376_));
  AOI220     u0348(.A0(men_men_n376_), .A1(men_men_n324_), .B0(men_men_n374_), .B1(men_men_n373_), .Y(men_men_n377_));
  NOi32      u0349(.An(j), .Bn(g), .C(i), .Y(men_men_n378_));
  NA3        u0350(.A(men_men_n378_), .B(men_men_n302_), .C(men_men_n117_), .Y(men_men_n379_));
  AO210      u0351(.A0(men_men_n115_), .A1(men_men_n32_), .B0(men_men_n379_), .Y(men_men_n380_));
  NOi32      u0352(.An(e), .Bn(b), .C(a), .Y(men_men_n381_));
  AN2        u0353(.A(l), .B(j), .Y(men_men_n382_));
  NO2        u0354(.A(men_men_n332_), .B(men_men_n382_), .Y(men_men_n383_));
  NO3        u0355(.A(men_men_n334_), .B(men_men_n72_), .C(men_men_n223_), .Y(men_men_n384_));
  NA3        u0356(.A(men_men_n217_), .B(men_men_n215_), .C(men_men_n35_), .Y(men_men_n385_));
  AOI220     u0357(.A0(men_men_n385_), .A1(men_men_n381_), .B0(men_men_n384_), .B1(men_men_n383_), .Y(men_men_n386_));
  NO2        u0358(.A(men_men_n344_), .B(n), .Y(men_men_n387_));
  NA2        u0359(.A(men_men_n216_), .B(k), .Y(men_men_n388_));
  NA3        u0360(.A(m), .B(men_men_n116_), .C(men_men_n222_), .Y(men_men_n389_));
  NA4        u0361(.A(men_men_n211_), .B(men_men_n89_), .C(g), .D(men_men_n222_), .Y(men_men_n390_));
  OAI210     u0362(.A0(men_men_n389_), .A1(men_men_n388_), .B0(men_men_n390_), .Y(men_men_n391_));
  NAi41      u0363(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n392_));
  NA2        u0364(.A(men_men_n51_), .B(men_men_n117_), .Y(men_men_n393_));
  NO2        u0365(.A(men_men_n393_), .B(men_men_n392_), .Y(men_men_n394_));
  AOI220     u0366(.A0(men_men_n394_), .A1(b), .B0(men_men_n391_), .B1(men_men_n387_), .Y(men_men_n395_));
  NA4        u0367(.A(men_men_n395_), .B(men_men_n386_), .C(men_men_n380_), .D(men_men_n377_), .Y(men_men_n396_));
  NO4        u0368(.A(men_men_n396_), .B(men_men_n371_), .C(men_men_n354_), .D(men_men_n347_), .Y(men_men_n397_));
  NA4        u0369(.A(men_men_n397_), .B(men_men_n330_), .C(men_men_n281_), .D(men_men_n207_), .Y(men10));
  NA3        u0370(.A(m), .B(k), .C(i), .Y(men_men_n399_));
  NO3        u0371(.A(men_men_n399_), .B(j), .C(men_men_n223_), .Y(men_men_n400_));
  NOi21      u0372(.An(e), .B(f), .Y(men_men_n401_));
  NO4        u0373(.A(men_men_n155_), .B(men_men_n401_), .C(n), .D(men_men_n114_), .Y(men_men_n402_));
  NAi31      u0374(.An(b), .B(f), .C(c), .Y(men_men_n403_));
  INV        u0375(.A(men_men_n403_), .Y(men_men_n404_));
  NOi32      u0376(.An(k), .Bn(h), .C(j), .Y(men_men_n405_));
  NA2        u0377(.A(men_men_n405_), .B(men_men_n230_), .Y(men_men_n406_));
  NA2        u0378(.A(men_men_n165_), .B(men_men_n406_), .Y(men_men_n407_));
  AOI220     u0379(.A0(men_men_n407_), .A1(men_men_n404_), .B0(men_men_n402_), .B1(men_men_n400_), .Y(men_men_n408_));
  AN2        u0380(.A(j), .B(h), .Y(men_men_n409_));
  NO3        u0381(.A(n), .B(m), .C(k), .Y(men_men_n410_));
  NA2        u0382(.A(men_men_n410_), .B(men_men_n409_), .Y(men_men_n411_));
  NO3        u0383(.A(men_men_n411_), .B(men_men_n155_), .C(men_men_n222_), .Y(men_men_n412_));
  OR2        u0384(.A(m), .B(k), .Y(men_men_n413_));
  NO2        u0385(.A(men_men_n180_), .B(men_men_n413_), .Y(men_men_n414_));
  NA4        u0386(.A(n), .B(f), .C(c), .D(men_men_n120_), .Y(men_men_n415_));
  NOi21      u0387(.An(men_men_n414_), .B(men_men_n415_), .Y(men_men_n416_));
  NOi32      u0388(.An(d), .Bn(a), .C(c), .Y(men_men_n417_));
  NA2        u0389(.A(men_men_n417_), .B(men_men_n188_), .Y(men_men_n418_));
  NAi21      u0390(.An(i), .B(g), .Y(men_men_n419_));
  NAi31      u0391(.An(k), .B(m), .C(j), .Y(men_men_n420_));
  NO3        u0392(.A(men_men_n420_), .B(men_men_n419_), .C(n), .Y(men_men_n421_));
  NOi21      u0393(.An(men_men_n421_), .B(men_men_n418_), .Y(men_men_n422_));
  NO3        u0394(.A(men_men_n422_), .B(men_men_n416_), .C(men_men_n412_), .Y(men_men_n423_));
  NO2        u0395(.A(men_men_n415_), .B(men_men_n311_), .Y(men_men_n424_));
  NOi32      u0396(.An(f), .Bn(d), .C(c), .Y(men_men_n425_));
  AOI220     u0397(.A0(men_men_n425_), .A1(men_men_n322_), .B0(men_men_n424_), .B1(men_men_n224_), .Y(men_men_n426_));
  NA3        u0398(.A(men_men_n426_), .B(men_men_n423_), .C(men_men_n408_), .Y(men_men_n427_));
  NO2        u0399(.A(men_men_n59_), .B(men_men_n120_), .Y(men_men_n428_));
  NA2        u0400(.A(men_men_n261_), .B(men_men_n428_), .Y(men_men_n429_));
  INV        u0401(.A(e), .Y(men_men_n430_));
  NA2        u0402(.A(men_men_n46_), .B(e), .Y(men_men_n431_));
  OAI220     u0403(.A0(men_men_n431_), .A1(men_men_n208_), .B0(men_men_n212_), .B1(men_men_n430_), .Y(men_men_n432_));
  AN2        u0404(.A(g), .B(e), .Y(men_men_n433_));
  NA3        u0405(.A(men_men_n433_), .B(men_men_n211_), .C(i), .Y(men_men_n434_));
  OAI210     u0406(.A0(men_men_n91_), .A1(men_men_n430_), .B0(men_men_n434_), .Y(men_men_n435_));
  NO2        u0407(.A(men_men_n103_), .B(men_men_n430_), .Y(men_men_n436_));
  NO3        u0408(.A(men_men_n436_), .B(men_men_n435_), .C(men_men_n432_), .Y(men_men_n437_));
  NOi32      u0409(.An(h), .Bn(e), .C(g), .Y(men_men_n438_));
  NA3        u0410(.A(men_men_n438_), .B(men_men_n304_), .C(m), .Y(men_men_n439_));
  NOi21      u0411(.An(g), .B(h), .Y(men_men_n440_));
  AN3        u0412(.A(m), .B(l), .C(i), .Y(men_men_n441_));
  NA3        u0413(.A(men_men_n441_), .B(men_men_n440_), .C(e), .Y(men_men_n442_));
  AN3        u0414(.A(h), .B(g), .C(e), .Y(men_men_n443_));
  NA2        u0415(.A(men_men_n443_), .B(men_men_n100_), .Y(men_men_n444_));
  AN3        u0416(.A(men_men_n444_), .B(men_men_n442_), .C(men_men_n439_), .Y(men_men_n445_));
  AOI210     u0417(.A0(men_men_n445_), .A1(men_men_n437_), .B0(men_men_n429_), .Y(men_men_n446_));
  NA3        u0418(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n447_));
  NO2        u0419(.A(men_men_n447_), .B(men_men_n429_), .Y(men_men_n448_));
  NAi31      u0420(.An(b), .B(c), .C(a), .Y(men_men_n449_));
  NO2        u0421(.A(men_men_n449_), .B(n), .Y(men_men_n450_));
  OAI210     u0422(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n451_));
  NO2        u0423(.A(men_men_n451_), .B(men_men_n151_), .Y(men_men_n452_));
  NA2        u0424(.A(men_men_n452_), .B(men_men_n450_), .Y(men_men_n453_));
  INV        u0425(.A(men_men_n453_), .Y(men_men_n454_));
  NO4        u0426(.A(men_men_n454_), .B(men_men_n448_), .C(men_men_n446_), .D(men_men_n427_), .Y(men_men_n455_));
  NA2        u0427(.A(i), .B(g), .Y(men_men_n456_));
  NO3        u0428(.A(men_men_n289_), .B(men_men_n456_), .C(c), .Y(men_men_n457_));
  NOi21      u0429(.An(a), .B(n), .Y(men_men_n458_));
  NOi21      u0430(.An(d), .B(c), .Y(men_men_n459_));
  NA2        u0431(.A(men_men_n459_), .B(men_men_n458_), .Y(men_men_n460_));
  NA3        u0432(.A(i), .B(g), .C(f), .Y(men_men_n461_));
  OR2        u0433(.A(men_men_n461_), .B(men_men_n71_), .Y(men_men_n462_));
  NA2        u0434(.A(men_men_n457_), .B(men_men_n303_), .Y(men_men_n463_));
  OR2        u0435(.A(n), .B(m), .Y(men_men_n464_));
  NO2        u0436(.A(men_men_n464_), .B(men_men_n156_), .Y(men_men_n465_));
  NO2        u0437(.A(men_men_n189_), .B(men_men_n151_), .Y(men_men_n466_));
  OAI210     u0438(.A0(men_men_n465_), .A1(men_men_n182_), .B0(men_men_n466_), .Y(men_men_n467_));
  INV        u0439(.A(men_men_n393_), .Y(men_men_n468_));
  NA3        u0440(.A(men_men_n468_), .B(men_men_n381_), .C(d), .Y(men_men_n469_));
  NO2        u0441(.A(men_men_n449_), .B(men_men_n49_), .Y(men_men_n470_));
  NAi21      u0442(.An(k), .B(j), .Y(men_men_n471_));
  NAi21      u0443(.An(e), .B(d), .Y(men_men_n472_));
  INV        u0444(.A(men_men_n472_), .Y(men_men_n473_));
  NO2        u0445(.A(men_men_n265_), .B(men_men_n222_), .Y(men_men_n474_));
  NA3        u0446(.A(men_men_n474_), .B(men_men_n473_), .C(men_men_n236_), .Y(men_men_n475_));
  NA3        u0447(.A(men_men_n475_), .B(men_men_n469_), .C(men_men_n467_), .Y(men_men_n476_));
  NO2        u0448(.A(men_men_n352_), .B(men_men_n222_), .Y(men_men_n477_));
  NA2        u0449(.A(men_men_n477_), .B(men_men_n473_), .Y(men_men_n478_));
  NOi31      u0450(.An(n), .B(m), .C(k), .Y(men_men_n479_));
  AOI220     u0451(.A0(men_men_n479_), .A1(men_men_n409_), .B0(men_men_n230_), .B1(men_men_n50_), .Y(men_men_n480_));
  NAi31      u0452(.An(g), .B(f), .C(c), .Y(men_men_n481_));
  OR3        u0453(.A(men_men_n481_), .B(men_men_n480_), .C(e), .Y(men_men_n482_));
  NA3        u0454(.A(men_men_n482_), .B(men_men_n478_), .C(men_men_n323_), .Y(men_men_n483_));
  NOi41      u0455(.An(men_men_n463_), .B(men_men_n483_), .C(men_men_n476_), .D(men_men_n279_), .Y(men_men_n484_));
  NOi32      u0456(.An(c), .Bn(a), .C(b), .Y(men_men_n485_));
  NA2        u0457(.A(men_men_n485_), .B(men_men_n117_), .Y(men_men_n486_));
  INV        u0458(.A(men_men_n287_), .Y(men_men_n487_));
  AN2        u0459(.A(e), .B(d), .Y(men_men_n488_));
  INV        u0460(.A(men_men_n151_), .Y(men_men_n489_));
  NO2        u0461(.A(men_men_n136_), .B(men_men_n41_), .Y(men_men_n490_));
  NO2        u0462(.A(men_men_n66_), .B(e), .Y(men_men_n491_));
  NOi31      u0463(.An(j), .B(k), .C(i), .Y(men_men_n492_));
  NOi21      u0464(.An(men_men_n170_), .B(men_men_n492_), .Y(men_men_n493_));
  NA4        u0465(.A(men_men_n337_), .B(men_men_n493_), .C(men_men_n273_), .D(men_men_n123_), .Y(men_men_n494_));
  NA2        u0466(.A(men_men_n494_), .B(men_men_n491_), .Y(men_men_n495_));
  NO2        u0467(.A(men_men_n495_), .B(men_men_n486_), .Y(men_men_n496_));
  NO2        u0468(.A(men_men_n218_), .B(men_men_n213_), .Y(men_men_n497_));
  NOi21      u0469(.An(a), .B(b), .Y(men_men_n498_));
  NA3        u0470(.A(e), .B(d), .C(c), .Y(men_men_n499_));
  NAi21      u0471(.An(men_men_n499_), .B(men_men_n498_), .Y(men_men_n500_));
  AOI210     u0472(.A0(men_men_n282_), .A1(men_men_n497_), .B0(men_men_n500_), .Y(men_men_n501_));
  NO4        u0473(.A(men_men_n195_), .B(men_men_n106_), .C(men_men_n56_), .D(b), .Y(men_men_n502_));
  NA2        u0474(.A(men_men_n404_), .B(men_men_n157_), .Y(men_men_n503_));
  OR2        u0475(.A(k), .B(j), .Y(men_men_n504_));
  NA2        u0476(.A(l), .B(k), .Y(men_men_n505_));
  NA3        u0477(.A(men_men_n505_), .B(men_men_n504_), .C(men_men_n230_), .Y(men_men_n506_));
  AOI210     u0478(.A0(men_men_n243_), .A1(men_men_n355_), .B0(men_men_n86_), .Y(men_men_n507_));
  NOi21      u0479(.An(men_men_n506_), .B(men_men_n507_), .Y(men_men_n508_));
  OR3        u0480(.A(men_men_n508_), .B(men_men_n148_), .C(men_men_n140_), .Y(men_men_n509_));
  NA2        u0481(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n510_));
  NA2        u0482(.A(men_men_n417_), .B(men_men_n117_), .Y(men_men_n511_));
  NO4        u0483(.A(men_men_n511_), .B(men_men_n97_), .C(men_men_n116_), .D(e), .Y(men_men_n512_));
  NO3        u0484(.A(men_men_n512_), .B(men_men_n510_), .C(men_men_n338_), .Y(men_men_n513_));
  NA3        u0485(.A(men_men_n513_), .B(men_men_n509_), .C(men_men_n503_), .Y(men_men_n514_));
  NO4        u0486(.A(men_men_n514_), .B(men_men_n502_), .C(men_men_n501_), .D(men_men_n496_), .Y(men_men_n515_));
  NA2        u0487(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n516_));
  NOi21      u0488(.An(d), .B(e), .Y(men_men_n517_));
  NO2        u0489(.A(men_men_n195_), .B(men_men_n56_), .Y(men_men_n518_));
  NAi31      u0490(.An(j), .B(l), .C(i), .Y(men_men_n519_));
  OAI210     u0491(.A0(men_men_n519_), .A1(men_men_n137_), .B0(men_men_n106_), .Y(men_men_n520_));
  NA4        u0492(.A(men_men_n520_), .B(men_men_n518_), .C(men_men_n517_), .D(b), .Y(men_men_n521_));
  NO3        u0493(.A(men_men_n418_), .B(men_men_n363_), .C(men_men_n209_), .Y(men_men_n522_));
  NO2        u0494(.A(men_men_n418_), .B(men_men_n393_), .Y(men_men_n523_));
  NO4        u0495(.A(men_men_n523_), .B(men_men_n522_), .C(men_men_n191_), .D(men_men_n320_), .Y(men_men_n524_));
  NA4        u0496(.A(men_men_n524_), .B(men_men_n521_), .C(men_men_n516_), .D(men_men_n253_), .Y(men_men_n525_));
  OAI210     u0497(.A0(men_men_n132_), .A1(men_men_n130_), .B0(n), .Y(men_men_n526_));
  NO2        u0498(.A(men_men_n526_), .B(men_men_n136_), .Y(men_men_n527_));
  OR2        u0499(.A(men_men_n312_), .B(men_men_n255_), .Y(men_men_n528_));
  OA210      u0500(.A0(men_men_n528_), .A1(men_men_n527_), .B0(men_men_n200_), .Y(men_men_n529_));
  XO2        u0501(.A(i), .B(h), .Y(men_men_n530_));
  NA3        u0502(.A(men_men_n530_), .B(men_men_n164_), .C(n), .Y(men_men_n531_));
  NAi41      u0503(.An(men_men_n312_), .B(men_men_n531_), .C(men_men_n480_), .D(men_men_n406_), .Y(men_men_n532_));
  NOi32      u0504(.An(men_men_n532_), .Bn(men_men_n491_), .C(men_men_n284_), .Y(men_men_n533_));
  NAi31      u0505(.An(c), .B(f), .C(d), .Y(men_men_n534_));
  AOI210     u0506(.A0(men_men_n292_), .A1(men_men_n203_), .B0(men_men_n534_), .Y(men_men_n535_));
  NOi21      u0507(.An(men_men_n84_), .B(men_men_n535_), .Y(men_men_n536_));
  NA2        u0508(.A(men_men_n237_), .B(men_men_n112_), .Y(men_men_n537_));
  AOI210     u0509(.A0(men_men_n537_), .A1(men_men_n187_), .B0(men_men_n534_), .Y(men_men_n538_));
  INV        u0510(.A(men_men_n538_), .Y(men_men_n539_));
  AO220      u0511(.A0(men_men_n300_), .A1(men_men_n276_), .B0(men_men_n171_), .B1(men_men_n67_), .Y(men_men_n540_));
  NA3        u0512(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n541_), .B(men_men_n460_), .Y(men_men_n542_));
  NO2        u0514(.A(men_men_n542_), .B(men_men_n308_), .Y(men_men_n543_));
  NAi41      u0515(.An(men_men_n540_), .B(men_men_n543_), .C(men_men_n539_), .D(men_men_n536_), .Y(men_men_n544_));
  NO4        u0516(.A(men_men_n544_), .B(men_men_n533_), .C(men_men_n529_), .D(men_men_n525_), .Y(men_men_n545_));
  NA4        u0517(.A(men_men_n545_), .B(men_men_n515_), .C(men_men_n484_), .D(men_men_n455_), .Y(men11));
  NO2        u0518(.A(men_men_n73_), .B(f), .Y(men_men_n547_));
  NA2        u0519(.A(j), .B(g), .Y(men_men_n548_));
  NAi31      u0520(.An(i), .B(m), .C(l), .Y(men_men_n549_));
  NA3        u0521(.A(m), .B(k), .C(j), .Y(men_men_n550_));
  OAI220     u0522(.A0(men_men_n550_), .A1(men_men_n136_), .B0(men_men_n549_), .B1(men_men_n548_), .Y(men_men_n551_));
  NA2        u0523(.A(men_men_n551_), .B(men_men_n547_), .Y(men_men_n552_));
  NOi32      u0524(.An(e), .Bn(b), .C(f), .Y(men_men_n553_));
  NA2        u0525(.A(men_men_n272_), .B(men_men_n117_), .Y(men_men_n554_));
  NA2        u0526(.A(men_men_n46_), .B(j), .Y(men_men_n555_));
  NO2        u0527(.A(men_men_n555_), .B(men_men_n314_), .Y(men_men_n556_));
  NAi31      u0528(.An(d), .B(e), .C(a), .Y(men_men_n557_));
  NO2        u0529(.A(men_men_n557_), .B(n), .Y(men_men_n558_));
  AOI220     u0530(.A0(men_men_n558_), .A1(men_men_n104_), .B0(men_men_n556_), .B1(men_men_n553_), .Y(men_men_n559_));
  NAi41      u0531(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n560_));
  AN2        u0532(.A(men_men_n560_), .B(men_men_n392_), .Y(men_men_n561_));
  AOI210     u0533(.A0(men_men_n561_), .A1(men_men_n418_), .B0(men_men_n285_), .Y(men_men_n562_));
  NA2        u0534(.A(j), .B(i), .Y(men_men_n563_));
  NAi31      u0535(.An(n), .B(m), .C(k), .Y(men_men_n564_));
  NO3        u0536(.A(men_men_n564_), .B(men_men_n563_), .C(men_men_n116_), .Y(men_men_n565_));
  NO4        u0537(.A(n), .B(d), .C(men_men_n120_), .D(a), .Y(men_men_n566_));
  OR2        u0538(.A(n), .B(c), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n567_), .B(men_men_n153_), .Y(men_men_n568_));
  NO2        u0540(.A(men_men_n568_), .B(men_men_n566_), .Y(men_men_n569_));
  NOi32      u0541(.An(g), .Bn(f), .C(i), .Y(men_men_n570_));
  AOI220     u0542(.A0(men_men_n570_), .A1(men_men_n102_), .B0(men_men_n551_), .B1(f), .Y(men_men_n571_));
  NO2        u0543(.A(men_men_n287_), .B(men_men_n49_), .Y(men_men_n572_));
  NO2        u0544(.A(men_men_n571_), .B(men_men_n569_), .Y(men_men_n573_));
  AOI210     u0545(.A0(men_men_n565_), .A1(men_men_n562_), .B0(men_men_n573_), .Y(men_men_n574_));
  NA2        u0546(.A(men_men_n145_), .B(men_men_n34_), .Y(men_men_n575_));
  OAI220     u0547(.A0(men_men_n575_), .A1(m), .B0(men_men_n555_), .B1(men_men_n243_), .Y(men_men_n576_));
  NOi41      u0548(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n577_));
  NAi32      u0549(.An(e), .Bn(b), .C(c), .Y(men_men_n578_));
  OR2        u0550(.A(men_men_n578_), .B(men_men_n86_), .Y(men_men_n579_));
  AN2        u0551(.A(men_men_n356_), .B(men_men_n334_), .Y(men_men_n580_));
  NA2        u0552(.A(men_men_n580_), .B(men_men_n579_), .Y(men_men_n581_));
  OA210      u0553(.A0(men_men_n581_), .A1(men_men_n577_), .B0(men_men_n576_), .Y(men_men_n582_));
  OAI220     u0554(.A0(men_men_n420_), .A1(men_men_n419_), .B0(men_men_n549_), .B1(men_men_n548_), .Y(men_men_n583_));
  NAi31      u0555(.An(d), .B(c), .C(a), .Y(men_men_n584_));
  NO2        u0556(.A(men_men_n584_), .B(n), .Y(men_men_n585_));
  NA3        u0557(.A(men_men_n585_), .B(men_men_n583_), .C(e), .Y(men_men_n586_));
  NO3        u0558(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n223_), .Y(men_men_n587_));
  NO2        u0559(.A(men_men_n240_), .B(men_men_n114_), .Y(men_men_n588_));
  OAI210     u0560(.A0(men_men_n587_), .A1(men_men_n421_), .B0(men_men_n588_), .Y(men_men_n589_));
  NA2        u0561(.A(men_men_n589_), .B(men_men_n586_), .Y(men_men_n590_));
  NO2        u0562(.A(men_men_n289_), .B(n), .Y(men_men_n591_));
  NO2        u0563(.A(men_men_n450_), .B(men_men_n591_), .Y(men_men_n592_));
  NA2        u0564(.A(men_men_n583_), .B(f), .Y(men_men_n593_));
  NA2        u0565(.A(h), .B(f), .Y(men_men_n594_));
  NO2        u0566(.A(men_men_n594_), .B(men_men_n97_), .Y(men_men_n595_));
  NO3        u0567(.A(men_men_n183_), .B(men_men_n180_), .C(g), .Y(men_men_n596_));
  NA2        u0568(.A(men_men_n596_), .B(men_men_n58_), .Y(men_men_n597_));
  OAI210     u0569(.A0(men_men_n593_), .A1(men_men_n592_), .B0(men_men_n597_), .Y(men_men_n598_));
  AN3        u0570(.A(j), .B(h), .C(g), .Y(men_men_n599_));
  NO2        u0571(.A(men_men_n150_), .B(c), .Y(men_men_n600_));
  NA3        u0572(.A(men_men_n600_), .B(men_men_n599_), .C(men_men_n479_), .Y(men_men_n601_));
  NA3        u0573(.A(f), .B(d), .C(b), .Y(men_men_n602_));
  INV        u0574(.A(men_men_n601_), .Y(men_men_n603_));
  NO4        u0575(.A(men_men_n603_), .B(men_men_n598_), .C(men_men_n590_), .D(men_men_n582_), .Y(men_men_n604_));
  AN4        u0576(.A(men_men_n604_), .B(men_men_n574_), .C(men_men_n559_), .D(men_men_n552_), .Y(men_men_n605_));
  INV        u0577(.A(k), .Y(men_men_n606_));
  NA3        u0578(.A(l), .B(men_men_n606_), .C(i), .Y(men_men_n607_));
  INV        u0579(.A(men_men_n607_), .Y(men_men_n608_));
  NAi32      u0580(.An(h), .Bn(f), .C(g), .Y(men_men_n609_));
  NAi41      u0581(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n610_));
  OAI210     u0582(.A0(men_men_n557_), .A1(n), .B0(men_men_n610_), .Y(men_men_n611_));
  NA2        u0583(.A(men_men_n611_), .B(m), .Y(men_men_n612_));
  NAi31      u0584(.An(h), .B(g), .C(f), .Y(men_men_n613_));
  OR3        u0585(.A(men_men_n613_), .B(men_men_n289_), .C(men_men_n49_), .Y(men_men_n614_));
  NA4        u0586(.A(men_men_n440_), .B(men_men_n125_), .C(men_men_n117_), .D(e), .Y(men_men_n615_));
  AN2        u0587(.A(men_men_n615_), .B(men_men_n614_), .Y(men_men_n616_));
  OA210      u0588(.A0(men_men_n612_), .A1(men_men_n609_), .B0(men_men_n616_), .Y(men_men_n617_));
  NO3        u0589(.A(men_men_n609_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n618_));
  NO4        u0590(.A(men_men_n613_), .B(men_men_n567_), .C(men_men_n153_), .D(men_men_n75_), .Y(men_men_n619_));
  OR2        u0591(.A(men_men_n619_), .B(men_men_n618_), .Y(men_men_n620_));
  NAi21      u0592(.An(men_men_n620_), .B(men_men_n617_), .Y(men_men_n621_));
  NAi31      u0593(.An(f), .B(h), .C(g), .Y(men_men_n622_));
  NO4        u0594(.A(men_men_n325_), .B(men_men_n622_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n623_));
  NOi32      u0595(.An(b), .Bn(a), .C(c), .Y(men_men_n624_));
  NOi41      u0596(.An(men_men_n624_), .B(men_men_n372_), .C(men_men_n69_), .D(men_men_n121_), .Y(men_men_n625_));
  OR2        u0597(.A(men_men_n625_), .B(men_men_n623_), .Y(men_men_n626_));
  NOi32      u0598(.An(d), .Bn(a), .C(e), .Y(men_men_n627_));
  NA2        u0599(.A(men_men_n627_), .B(men_men_n117_), .Y(men_men_n628_));
  NO2        u0600(.A(n), .B(c), .Y(men_men_n629_));
  NA3        u0601(.A(men_men_n629_), .B(men_men_n29_), .C(m), .Y(men_men_n630_));
  NAi32      u0602(.An(n), .Bn(f), .C(m), .Y(men_men_n631_));
  NA3        u0603(.A(men_men_n631_), .B(men_men_n630_), .C(men_men_n628_), .Y(men_men_n632_));
  NOi32      u0604(.An(e), .Bn(a), .C(d), .Y(men_men_n633_));
  AOI210     u0605(.A0(men_men_n29_), .A1(d), .B0(men_men_n633_), .Y(men_men_n634_));
  AOI210     u0606(.A0(men_men_n634_), .A1(men_men_n222_), .B0(men_men_n575_), .Y(men_men_n635_));
  AOI210     u0607(.A0(men_men_n635_), .A1(men_men_n632_), .B0(men_men_n626_), .Y(men_men_n636_));
  OAI210     u0608(.A0(men_men_n260_), .A1(men_men_n89_), .B0(men_men_n636_), .Y(men_men_n637_));
  AOI210     u0609(.A0(men_men_n621_), .A1(men_men_n608_), .B0(men_men_n637_), .Y(men_men_n638_));
  NO3        u0610(.A(men_men_n332_), .B(men_men_n61_), .C(n), .Y(men_men_n639_));
  NA3        u0611(.A(men_men_n534_), .B(men_men_n178_), .C(men_men_n177_), .Y(men_men_n640_));
  NA2        u0612(.A(men_men_n481_), .B(men_men_n240_), .Y(men_men_n641_));
  OR2        u0613(.A(men_men_n641_), .B(men_men_n640_), .Y(men_men_n642_));
  NA2        u0614(.A(men_men_n76_), .B(men_men_n117_), .Y(men_men_n643_));
  NO2        u0615(.A(men_men_n643_), .B(men_men_n45_), .Y(men_men_n644_));
  AOI220     u0616(.A0(men_men_n644_), .A1(men_men_n562_), .B0(men_men_n642_), .B1(men_men_n639_), .Y(men_men_n645_));
  NO2        u0617(.A(men_men_n645_), .B(men_men_n89_), .Y(men_men_n646_));
  NA3        u0618(.A(men_men_n577_), .B(men_men_n358_), .C(men_men_n46_), .Y(men_men_n647_));
  NOi32      u0619(.An(e), .Bn(c), .C(f), .Y(men_men_n648_));
  NOi21      u0620(.An(f), .B(g), .Y(men_men_n649_));
  NO2        u0621(.A(men_men_n649_), .B(men_men_n220_), .Y(men_men_n650_));
  AOI220     u0622(.A0(men_men_n650_), .A1(men_men_n414_), .B0(men_men_n648_), .B1(men_men_n182_), .Y(men_men_n651_));
  NA3        u0623(.A(men_men_n651_), .B(men_men_n647_), .C(men_men_n185_), .Y(men_men_n652_));
  AOI210     u0624(.A0(men_men_n561_), .A1(men_men_n418_), .B0(men_men_n313_), .Y(men_men_n653_));
  NA2        u0625(.A(men_men_n653_), .B(men_men_n277_), .Y(men_men_n654_));
  NOi21      u0626(.An(j), .B(l), .Y(men_men_n655_));
  NAi21      u0627(.An(k), .B(h), .Y(men_men_n656_));
  NO2        u0628(.A(men_men_n656_), .B(men_men_n275_), .Y(men_men_n657_));
  NA2        u0629(.A(men_men_n657_), .B(men_men_n655_), .Y(men_men_n658_));
  OR2        u0630(.A(men_men_n658_), .B(men_men_n612_), .Y(men_men_n659_));
  NOi31      u0631(.An(m), .B(n), .C(k), .Y(men_men_n660_));
  NA2        u0632(.A(men_men_n655_), .B(men_men_n660_), .Y(men_men_n661_));
  AOI210     u0633(.A0(men_men_n418_), .A1(men_men_n392_), .B0(men_men_n313_), .Y(men_men_n662_));
  NAi21      u0634(.An(men_men_n661_), .B(men_men_n662_), .Y(men_men_n663_));
  NO2        u0635(.A(men_men_n289_), .B(men_men_n49_), .Y(men_men_n664_));
  NO2        u0636(.A(men_men_n325_), .B(men_men_n622_), .Y(men_men_n665_));
  NO2        u0637(.A(men_men_n557_), .B(men_men_n49_), .Y(men_men_n666_));
  AOI220     u0638(.A0(men_men_n666_), .A1(men_men_n665_), .B0(men_men_n664_), .B1(men_men_n595_), .Y(men_men_n667_));
  NA4        u0639(.A(men_men_n667_), .B(men_men_n663_), .C(men_men_n659_), .D(men_men_n654_), .Y(men_men_n668_));
  NA2        u0640(.A(men_men_n112_), .B(men_men_n36_), .Y(men_men_n669_));
  NO2        u0641(.A(k), .B(men_men_n223_), .Y(men_men_n670_));
  NO2        u0642(.A(men_men_n553_), .B(men_men_n381_), .Y(men_men_n671_));
  NO2        u0643(.A(men_men_n671_), .B(n), .Y(men_men_n672_));
  NAi31      u0644(.An(men_men_n669_), .B(men_men_n672_), .C(men_men_n670_), .Y(men_men_n673_));
  NO2        u0645(.A(men_men_n555_), .B(men_men_n183_), .Y(men_men_n674_));
  NA3        u0646(.A(men_men_n578_), .B(men_men_n284_), .C(men_men_n149_), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n530_), .B(men_men_n164_), .Y(men_men_n676_));
  NO3        u0648(.A(men_men_n415_), .B(men_men_n676_), .C(men_men_n89_), .Y(men_men_n677_));
  AOI210     u0649(.A0(men_men_n675_), .A1(men_men_n674_), .B0(men_men_n677_), .Y(men_men_n678_));
  AN3        u0650(.A(f), .B(d), .C(b), .Y(men_men_n679_));
  OAI210     u0651(.A0(men_men_n679_), .A1(men_men_n135_), .B0(n), .Y(men_men_n680_));
  NA3        u0652(.A(men_men_n530_), .B(men_men_n164_), .C(men_men_n223_), .Y(men_men_n681_));
  AOI210     u0653(.A0(men_men_n680_), .A1(men_men_n242_), .B0(men_men_n681_), .Y(men_men_n682_));
  NAi31      u0654(.An(m), .B(n), .C(k), .Y(men_men_n683_));
  OR2        u0655(.A(men_men_n140_), .B(men_men_n61_), .Y(men_men_n684_));
  OAI210     u0656(.A0(men_men_n684_), .A1(men_men_n683_), .B0(men_men_n262_), .Y(men_men_n685_));
  OAI210     u0657(.A0(men_men_n685_), .A1(men_men_n682_), .B0(j), .Y(men_men_n686_));
  NA3        u0658(.A(men_men_n686_), .B(men_men_n678_), .C(men_men_n673_), .Y(men_men_n687_));
  NO4        u0659(.A(men_men_n687_), .B(men_men_n668_), .C(men_men_n652_), .D(men_men_n646_), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n402_), .B(men_men_n167_), .Y(men_men_n689_));
  NAi31      u0661(.An(g), .B(h), .C(f), .Y(men_men_n690_));
  OR3        u0662(.A(men_men_n690_), .B(men_men_n289_), .C(n), .Y(men_men_n691_));
  OA210      u0663(.A0(men_men_n557_), .A1(n), .B0(men_men_n610_), .Y(men_men_n692_));
  NA3        u0664(.A(men_men_n438_), .B(men_men_n125_), .C(men_men_n86_), .Y(men_men_n693_));
  OAI210     u0665(.A0(men_men_n692_), .A1(men_men_n93_), .B0(men_men_n693_), .Y(men_men_n694_));
  NOi21      u0666(.An(men_men_n691_), .B(men_men_n694_), .Y(men_men_n695_));
  AOI210     u0667(.A0(men_men_n695_), .A1(men_men_n689_), .B0(men_men_n550_), .Y(men_men_n696_));
  NO3        u0668(.A(g), .B(men_men_n222_), .C(men_men_n56_), .Y(men_men_n697_));
  NO2        u0669(.A(men_men_n537_), .B(men_men_n89_), .Y(men_men_n698_));
  OAI210     u0670(.A0(men_men_n698_), .A1(men_men_n414_), .B0(men_men_n697_), .Y(men_men_n699_));
  OR2        u0671(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n700_));
  NA2        u0672(.A(men_men_n624_), .B(men_men_n360_), .Y(men_men_n701_));
  OA220      u0673(.A0(men_men_n661_), .A1(men_men_n701_), .B0(men_men_n658_), .B1(men_men_n700_), .Y(men_men_n702_));
  NA3        u0674(.A(men_men_n547_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n703_));
  AN2        u0675(.A(h), .B(f), .Y(men_men_n704_));
  NA2        u0676(.A(men_men_n704_), .B(men_men_n37_), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n102_), .B(men_men_n46_), .Y(men_men_n706_));
  OAI220     u0678(.A0(men_men_n706_), .A1(men_men_n349_), .B0(men_men_n705_), .B1(men_men_n486_), .Y(men_men_n707_));
  INV        u0679(.A(men_men_n707_), .Y(men_men_n708_));
  NA4        u0680(.A(men_men_n708_), .B(men_men_n703_), .C(men_men_n702_), .D(men_men_n699_), .Y(men_men_n709_));
  NO2        u0681(.A(men_men_n264_), .B(f), .Y(men_men_n710_));
  NO2        u0682(.A(men_men_n649_), .B(men_men_n61_), .Y(men_men_n711_));
  NO3        u0683(.A(men_men_n711_), .B(men_men_n710_), .C(men_men_n34_), .Y(men_men_n712_));
  NA2        u0684(.A(men_men_n345_), .B(men_men_n145_), .Y(men_men_n713_));
  NA2        u0685(.A(men_men_n137_), .B(men_men_n49_), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n381_), .B(men_men_n117_), .Y(men_men_n715_));
  OA220      u0687(.A0(men_men_n715_), .A1(men_men_n575_), .B0(men_men_n379_), .B1(men_men_n115_), .Y(men_men_n716_));
  OAI210     u0688(.A0(men_men_n713_), .A1(men_men_n712_), .B0(men_men_n716_), .Y(men_men_n717_));
  NO3        u0689(.A(men_men_n425_), .B(men_men_n200_), .C(men_men_n199_), .Y(men_men_n718_));
  NA2        u0690(.A(men_men_n718_), .B(men_men_n240_), .Y(men_men_n719_));
  NA3        u0691(.A(men_men_n719_), .B(men_men_n266_), .C(j), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n485_), .B(men_men_n86_), .Y(men_men_n721_));
  NA2        u0693(.A(men_men_n720_), .B(men_men_n423_), .Y(men_men_n722_));
  NO4        u0694(.A(men_men_n722_), .B(men_men_n717_), .C(men_men_n709_), .D(men_men_n696_), .Y(men_men_n723_));
  NA4        u0695(.A(men_men_n723_), .B(men_men_n688_), .C(men_men_n638_), .D(men_men_n605_), .Y(men08));
  NO2        u0696(.A(k), .B(h), .Y(men_men_n725_));
  AO210      u0697(.A0(men_men_n264_), .A1(men_men_n471_), .B0(men_men_n725_), .Y(men_men_n726_));
  NO2        u0698(.A(men_men_n726_), .B(men_men_n311_), .Y(men_men_n727_));
  NA2        u0699(.A(men_men_n648_), .B(men_men_n86_), .Y(men_men_n728_));
  NA2        u0700(.A(men_men_n728_), .B(men_men_n481_), .Y(men_men_n729_));
  NA2        u0701(.A(men_men_n729_), .B(men_men_n727_), .Y(men_men_n730_));
  NA2        u0702(.A(men_men_n86_), .B(men_men_n114_), .Y(men_men_n731_));
  NO2        u0703(.A(men_men_n731_), .B(men_men_n57_), .Y(men_men_n732_));
  NO4        u0704(.A(men_men_n399_), .B(men_men_n116_), .C(j), .D(men_men_n223_), .Y(men_men_n733_));
  NA2        u0705(.A(men_men_n602_), .B(men_men_n242_), .Y(men_men_n734_));
  AOI220     u0706(.A0(men_men_n734_), .A1(men_men_n366_), .B0(men_men_n733_), .B1(men_men_n732_), .Y(men_men_n735_));
  AOI210     u0707(.A0(men_men_n602_), .A1(men_men_n160_), .B0(men_men_n86_), .Y(men_men_n736_));
  NA4        u0708(.A(men_men_n225_), .B(men_men_n145_), .C(men_men_n45_), .D(h), .Y(men_men_n737_));
  AN2        u0709(.A(l), .B(k), .Y(men_men_n738_));
  NA4        u0710(.A(men_men_n738_), .B(men_men_n112_), .C(men_men_n75_), .D(men_men_n223_), .Y(men_men_n739_));
  OAI210     u0711(.A0(men_men_n737_), .A1(g), .B0(men_men_n739_), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n740_), .B(men_men_n736_), .Y(men_men_n741_));
  NA4        u0713(.A(men_men_n741_), .B(men_men_n735_), .C(men_men_n730_), .D(men_men_n368_), .Y(men_men_n742_));
  AN2        u0714(.A(men_men_n558_), .B(men_men_n98_), .Y(men_men_n743_));
  NO4        u0715(.A(men_men_n180_), .B(men_men_n413_), .C(men_men_n116_), .D(g), .Y(men_men_n744_));
  AOI210     u0716(.A0(men_men_n744_), .A1(men_men_n734_), .B0(men_men_n542_), .Y(men_men_n745_));
  NO2        u0717(.A(men_men_n38_), .B(men_men_n222_), .Y(men_men_n746_));
  AOI220     u0718(.A0(men_men_n650_), .A1(men_men_n365_), .B0(men_men_n746_), .B1(men_men_n591_), .Y(men_men_n747_));
  NAi31      u0719(.An(men_men_n743_), .B(men_men_n747_), .C(men_men_n745_), .Y(men_men_n748_));
  NO2        u0720(.A(men_men_n561_), .B(men_men_n35_), .Y(men_men_n749_));
  OAI210     u0721(.A0(men_men_n578_), .A1(men_men_n47_), .B0(men_men_n684_), .Y(men_men_n750_));
  NO2        u0722(.A(men_men_n505_), .B(men_men_n137_), .Y(men_men_n751_));
  AOI210     u0723(.A0(men_men_n751_), .A1(men_men_n750_), .B0(men_men_n749_), .Y(men_men_n752_));
  NO3        u0724(.A(men_men_n332_), .B(men_men_n136_), .C(men_men_n41_), .Y(men_men_n753_));
  NAi21      u0725(.An(men_men_n753_), .B(men_men_n739_), .Y(men_men_n754_));
  NA2        u0726(.A(men_men_n726_), .B(men_men_n141_), .Y(men_men_n755_));
  AOI220     u0727(.A0(men_men_n755_), .A1(men_men_n424_), .B0(men_men_n754_), .B1(men_men_n78_), .Y(men_men_n756_));
  OAI210     u0728(.A0(men_men_n752_), .A1(men_men_n89_), .B0(men_men_n756_), .Y(men_men_n757_));
  NA2        u0729(.A(men_men_n381_), .B(men_men_n43_), .Y(men_men_n758_));
  NA3        u0730(.A(men_men_n719_), .B(men_men_n351_), .C(men_men_n405_), .Y(men_men_n759_));
  NA2        u0731(.A(men_men_n738_), .B(men_men_n230_), .Y(men_men_n760_));
  NO2        u0732(.A(men_men_n760_), .B(men_men_n344_), .Y(men_men_n761_));
  AOI210     u0733(.A0(men_men_n761_), .A1(men_men_n710_), .B0(men_men_n512_), .Y(men_men_n762_));
  NA3        u0734(.A(m), .B(l), .C(k), .Y(men_men_n763_));
  AOI210     u0735(.A0(men_men_n693_), .A1(men_men_n691_), .B0(men_men_n763_), .Y(men_men_n764_));
  NO2        u0736(.A(men_men_n560_), .B(men_men_n285_), .Y(men_men_n765_));
  NOi21      u0737(.An(men_men_n765_), .B(men_men_n554_), .Y(men_men_n766_));
  NA4        u0738(.A(men_men_n117_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n767_));
  NA3        u0739(.A(men_men_n125_), .B(men_men_n433_), .C(i), .Y(men_men_n768_));
  NO2        u0740(.A(men_men_n768_), .B(men_men_n767_), .Y(men_men_n769_));
  NO3        u0741(.A(men_men_n769_), .B(men_men_n766_), .C(men_men_n764_), .Y(men_men_n770_));
  NA4        u0742(.A(men_men_n770_), .B(men_men_n762_), .C(men_men_n759_), .D(men_men_n758_), .Y(men_men_n771_));
  NO4        u0743(.A(men_men_n771_), .B(men_men_n757_), .C(men_men_n748_), .D(men_men_n742_), .Y(men_men_n772_));
  NA2        u0744(.A(men_men_n650_), .B(men_men_n414_), .Y(men_men_n773_));
  NOi31      u0745(.An(g), .B(h), .C(f), .Y(men_men_n774_));
  NA2        u0746(.A(men_men_n666_), .B(men_men_n774_), .Y(men_men_n775_));
  AO210      u0747(.A0(men_men_n775_), .A1(men_men_n614_), .B0(men_men_n563_), .Y(men_men_n776_));
  INV        u0748(.A(men_men_n523_), .Y(men_men_n777_));
  NA4        u0749(.A(men_men_n777_), .B(men_men_n776_), .C(men_men_n773_), .D(men_men_n263_), .Y(men_men_n778_));
  NA2        u0750(.A(men_men_n738_), .B(men_men_n75_), .Y(men_men_n779_));
  NO4        u0751(.A(men_men_n718_), .B(men_men_n180_), .C(n), .D(i), .Y(men_men_n780_));
  NOi21      u0752(.An(h), .B(j), .Y(men_men_n781_));
  NA2        u0753(.A(men_men_n781_), .B(f), .Y(men_men_n782_));
  NO2        u0754(.A(men_men_n782_), .B(men_men_n257_), .Y(men_men_n783_));
  NO2        u0755(.A(men_men_n783_), .B(men_men_n780_), .Y(men_men_n784_));
  OAI220     u0756(.A0(men_men_n784_), .A1(men_men_n779_), .B0(men_men_n616_), .B1(men_men_n62_), .Y(men_men_n785_));
  AOI210     u0757(.A0(men_men_n778_), .A1(l), .B0(men_men_n785_), .Y(men_men_n786_));
  NO2        u0758(.A(j), .B(i), .Y(men_men_n787_));
  NA3        u0759(.A(men_men_n787_), .B(men_men_n82_), .C(l), .Y(men_men_n788_));
  NA2        u0760(.A(men_men_n787_), .B(men_men_n33_), .Y(men_men_n789_));
  NA2        u0761(.A(men_men_n443_), .B(men_men_n125_), .Y(men_men_n790_));
  OA220      u0762(.A0(men_men_n790_), .A1(men_men_n789_), .B0(men_men_n788_), .B1(men_men_n612_), .Y(men_men_n791_));
  NO3        u0763(.A(men_men_n155_), .B(men_men_n49_), .C(men_men_n114_), .Y(men_men_n792_));
  NO3        u0764(.A(men_men_n567_), .B(men_men_n153_), .C(men_men_n75_), .Y(men_men_n793_));
  NO3        u0765(.A(men_men_n505_), .B(men_men_n461_), .C(j), .Y(men_men_n794_));
  OAI210     u0766(.A0(men_men_n793_), .A1(men_men_n792_), .B0(men_men_n794_), .Y(men_men_n795_));
  OAI210     u0767(.A0(men_men_n775_), .A1(men_men_n62_), .B0(men_men_n795_), .Y(men_men_n796_));
  NA2        u0768(.A(k), .B(j), .Y(men_men_n797_));
  NO3        u0769(.A(men_men_n311_), .B(men_men_n797_), .C(men_men_n40_), .Y(men_men_n798_));
  AOI210     u0770(.A0(men_men_n553_), .A1(n), .B0(men_men_n577_), .Y(men_men_n799_));
  NA2        u0771(.A(men_men_n799_), .B(men_men_n580_), .Y(men_men_n800_));
  AN3        u0772(.A(men_men_n800_), .B(men_men_n798_), .C(men_men_n101_), .Y(men_men_n801_));
  NO3        u0773(.A(men_men_n180_), .B(men_men_n413_), .C(men_men_n116_), .Y(men_men_n802_));
  AOI220     u0774(.A0(men_men_n802_), .A1(men_men_n258_), .B0(men_men_n641_), .B1(men_men_n322_), .Y(men_men_n803_));
  NAi31      u0775(.An(men_men_n634_), .B(men_men_n95_), .C(men_men_n86_), .Y(men_men_n804_));
  NA2        u0776(.A(men_men_n804_), .B(men_men_n803_), .Y(men_men_n805_));
  NO2        u0777(.A(men_men_n311_), .B(men_men_n141_), .Y(men_men_n806_));
  AOI220     u0778(.A0(men_men_n806_), .A1(men_men_n650_), .B0(men_men_n753_), .B1(men_men_n736_), .Y(men_men_n807_));
  INV        u0779(.A(men_men_n807_), .Y(men_men_n808_));
  OR4        u0780(.A(men_men_n808_), .B(men_men_n805_), .C(men_men_n801_), .D(men_men_n796_), .Y(men_men_n809_));
  NA3        u0781(.A(men_men_n799_), .B(men_men_n580_), .C(men_men_n579_), .Y(men_men_n810_));
  NA4        u0782(.A(men_men_n810_), .B(men_men_n225_), .C(men_men_n471_), .D(men_men_n34_), .Y(men_men_n811_));
  NO4        u0783(.A(men_men_n505_), .B(men_men_n456_), .C(j), .D(f), .Y(men_men_n812_));
  OAI220     u0784(.A0(men_men_n737_), .A1(men_men_n728_), .B0(men_men_n349_), .B1(men_men_n38_), .Y(men_men_n813_));
  AOI210     u0785(.A0(men_men_n812_), .A1(men_men_n270_), .B0(men_men_n813_), .Y(men_men_n814_));
  NA3        u0786(.A(men_men_n570_), .B(men_men_n304_), .C(h), .Y(men_men_n815_));
  NO2        u0787(.A(men_men_n94_), .B(men_men_n47_), .Y(men_men_n816_));
  OAI220     u0788(.A0(men_men_n815_), .A1(men_men_n630_), .B0(men_men_n788_), .B1(men_men_n700_), .Y(men_men_n817_));
  AOI210     u0789(.A0(men_men_n816_), .A1(men_men_n672_), .B0(men_men_n817_), .Y(men_men_n818_));
  NA3        u0790(.A(men_men_n818_), .B(men_men_n814_), .C(men_men_n811_), .Y(men_men_n819_));
  AOI220     u0791(.A0(men_men_n98_), .A1(men_men_n248_), .B0(men_men_n794_), .B1(men_men_n664_), .Y(men_men_n820_));
  NO2        u0792(.A(men_men_n692_), .B(men_men_n75_), .Y(men_men_n821_));
  AOI210     u0793(.A0(men_men_n812_), .A1(men_men_n821_), .B0(men_men_n353_), .Y(men_men_n822_));
  OAI210     u0794(.A0(men_men_n763_), .A1(men_men_n690_), .B0(men_men_n541_), .Y(men_men_n823_));
  NA3        u0795(.A(men_men_n261_), .B(men_men_n59_), .C(b), .Y(men_men_n824_));
  AOI220     u0796(.A0(men_men_n629_), .A1(men_men_n29_), .B0(men_men_n485_), .B1(men_men_n86_), .Y(men_men_n825_));
  NA2        u0797(.A(men_men_n825_), .B(men_men_n824_), .Y(men_men_n826_));
  NO2        u0798(.A(men_men_n815_), .B(men_men_n511_), .Y(men_men_n827_));
  AOI210     u0799(.A0(men_men_n826_), .A1(men_men_n823_), .B0(men_men_n827_), .Y(men_men_n828_));
  NA3        u0800(.A(men_men_n828_), .B(men_men_n822_), .C(men_men_n820_), .Y(men_men_n829_));
  NOi41      u0801(.An(men_men_n791_), .B(men_men_n829_), .C(men_men_n819_), .D(men_men_n809_), .Y(men_men_n830_));
  OR3        u0802(.A(men_men_n737_), .B(men_men_n242_), .C(g), .Y(men_men_n831_));
  NO3        u0803(.A(men_men_n359_), .B(men_men_n313_), .C(men_men_n116_), .Y(men_men_n832_));
  NA2        u0804(.A(men_men_n832_), .B(men_men_n800_), .Y(men_men_n833_));
  NA2        u0805(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n834_));
  NO3        u0806(.A(men_men_n834_), .B(men_men_n789_), .C(men_men_n289_), .Y(men_men_n835_));
  NO3        u0807(.A(men_men_n548_), .B(men_men_n96_), .C(h), .Y(men_men_n836_));
  AOI210     u0808(.A0(men_men_n836_), .A1(men_men_n732_), .B0(men_men_n835_), .Y(men_men_n837_));
  NA4        u0809(.A(men_men_n837_), .B(men_men_n833_), .C(men_men_n831_), .D(men_men_n426_), .Y(men_men_n838_));
  OR2        u0810(.A(men_men_n690_), .B(men_men_n94_), .Y(men_men_n839_));
  NOi31      u0811(.An(b), .B(d), .C(a), .Y(men_men_n840_));
  NO2        u0812(.A(men_men_n840_), .B(men_men_n627_), .Y(men_men_n841_));
  NO2        u0813(.A(men_men_n841_), .B(n), .Y(men_men_n842_));
  NOi21      u0814(.An(men_men_n825_), .B(men_men_n842_), .Y(men_men_n843_));
  OAI220     u0815(.A0(men_men_n843_), .A1(men_men_n839_), .B0(men_men_n815_), .B1(men_men_n628_), .Y(men_men_n844_));
  NO2        u0816(.A(men_men_n578_), .B(men_men_n86_), .Y(men_men_n845_));
  NO3        u0817(.A(men_men_n649_), .B(men_men_n344_), .C(men_men_n121_), .Y(men_men_n846_));
  NOi21      u0818(.An(men_men_n846_), .B(men_men_n165_), .Y(men_men_n847_));
  AOI210     u0819(.A0(men_men_n832_), .A1(men_men_n845_), .B0(men_men_n847_), .Y(men_men_n848_));
  OAI210     u0820(.A0(men_men_n737_), .A1(men_men_n415_), .B0(men_men_n848_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n718_), .B(n), .Y(men_men_n850_));
  AOI220     u0822(.A0(men_men_n806_), .A1(men_men_n697_), .B0(men_men_n850_), .B1(men_men_n727_), .Y(men_men_n851_));
  NO2        u0823(.A(men_men_n339_), .B(men_men_n247_), .Y(men_men_n852_));
  OAI210     u0824(.A0(men_men_n98_), .A1(men_men_n95_), .B0(men_men_n852_), .Y(men_men_n853_));
  NA2        u0825(.A(men_men_n125_), .B(men_men_n86_), .Y(men_men_n854_));
  AOI210     u0826(.A0(men_men_n447_), .A1(men_men_n439_), .B0(men_men_n854_), .Y(men_men_n855_));
  NAi21      u0827(.An(men_men_n855_), .B(men_men_n853_), .Y(men_men_n856_));
  NA2        u0828(.A(men_men_n761_), .B(men_men_n34_), .Y(men_men_n857_));
  NAi21      u0829(.An(men_men_n767_), .B(men_men_n457_), .Y(men_men_n858_));
  NO2        u0830(.A(men_men_n285_), .B(i), .Y(men_men_n859_));
  NA2        u0831(.A(men_men_n744_), .B(men_men_n367_), .Y(men_men_n860_));
  OAI210     u0832(.A0(men_men_n619_), .A1(men_men_n618_), .B0(men_men_n382_), .Y(men_men_n861_));
  AN3        u0833(.A(men_men_n861_), .B(men_men_n860_), .C(men_men_n858_), .Y(men_men_n862_));
  NAi41      u0834(.An(men_men_n856_), .B(men_men_n862_), .C(men_men_n857_), .D(men_men_n851_), .Y(men_men_n863_));
  NO4        u0835(.A(men_men_n863_), .B(men_men_n849_), .C(men_men_n844_), .D(men_men_n838_), .Y(men_men_n864_));
  NA4        u0836(.A(men_men_n864_), .B(men_men_n830_), .C(men_men_n786_), .D(men_men_n772_), .Y(men09));
  INV        u0837(.A(men_men_n126_), .Y(men_men_n866_));
  NA2        u0838(.A(f), .B(e), .Y(men_men_n867_));
  NO2        u0839(.A(men_men_n235_), .B(men_men_n116_), .Y(men_men_n868_));
  NA2        u0840(.A(men_men_n868_), .B(g), .Y(men_men_n869_));
  NA4        u0841(.A(men_men_n325_), .B(men_men_n493_), .C(men_men_n273_), .D(men_men_n123_), .Y(men_men_n870_));
  AOI210     u0842(.A0(men_men_n870_), .A1(g), .B0(men_men_n490_), .Y(men_men_n871_));
  AOI210     u0843(.A0(men_men_n871_), .A1(men_men_n869_), .B0(men_men_n867_), .Y(men_men_n872_));
  NA2        u0844(.A(men_men_n465_), .B(e), .Y(men_men_n873_));
  NO2        u0845(.A(men_men_n873_), .B(men_men_n534_), .Y(men_men_n874_));
  AOI210     u0846(.A0(men_men_n872_), .A1(men_men_n866_), .B0(men_men_n874_), .Y(men_men_n875_));
  NO2        u0847(.A(men_men_n212_), .B(men_men_n222_), .Y(men_men_n876_));
  NA3        u0848(.A(m), .B(l), .C(i), .Y(men_men_n877_));
  OAI220     u0849(.A0(men_men_n613_), .A1(men_men_n877_), .B0(men_men_n372_), .B1(men_men_n549_), .Y(men_men_n878_));
  NA4        u0850(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(f), .Y(men_men_n879_));
  NAi31      u0851(.An(men_men_n878_), .B(men_men_n879_), .C(men_men_n462_), .Y(men_men_n880_));
  OR2        u0852(.A(men_men_n880_), .B(men_men_n876_), .Y(men_men_n881_));
  NA3        u0853(.A(men_men_n839_), .B(men_men_n593_), .C(men_men_n541_), .Y(men_men_n882_));
  OA210      u0854(.A0(men_men_n882_), .A1(men_men_n881_), .B0(men_men_n842_), .Y(men_men_n883_));
  INV        u0855(.A(men_men_n356_), .Y(men_men_n884_));
  NO2        u0856(.A(men_men_n132_), .B(men_men_n130_), .Y(men_men_n885_));
  NOi31      u0857(.An(k), .B(m), .C(l), .Y(men_men_n886_));
  NO2        u0858(.A(men_men_n358_), .B(men_men_n886_), .Y(men_men_n887_));
  AOI210     u0859(.A0(men_men_n887_), .A1(men_men_n885_), .B0(men_men_n622_), .Y(men_men_n888_));
  NA2        u0860(.A(men_men_n824_), .B(men_men_n349_), .Y(men_men_n889_));
  NA2        u0861(.A(men_men_n360_), .B(men_men_n362_), .Y(men_men_n890_));
  OAI210     u0862(.A0(men_men_n212_), .A1(men_men_n222_), .B0(men_men_n890_), .Y(men_men_n891_));
  AOI220     u0863(.A0(men_men_n891_), .A1(men_men_n889_), .B0(men_men_n888_), .B1(men_men_n884_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n174_), .B(men_men_n118_), .Y(men_men_n893_));
  NA3        u0865(.A(men_men_n893_), .B(men_men_n726_), .C(men_men_n141_), .Y(men_men_n894_));
  NA3        u0866(.A(men_men_n894_), .B(men_men_n197_), .C(men_men_n31_), .Y(men_men_n895_));
  NA4        u0867(.A(men_men_n895_), .B(men_men_n892_), .C(men_men_n651_), .D(men_men_n84_), .Y(men_men_n896_));
  NO2        u0868(.A(men_men_n609_), .B(men_men_n519_), .Y(men_men_n897_));
  NOi21      u0869(.An(f), .B(d), .Y(men_men_n898_));
  NA2        u0870(.A(men_men_n898_), .B(m), .Y(men_men_n899_));
  NO2        u0871(.A(men_men_n899_), .B(men_men_n52_), .Y(men_men_n900_));
  NOi32      u0872(.An(g), .Bn(f), .C(d), .Y(men_men_n901_));
  NA4        u0873(.A(men_men_n901_), .B(men_men_n629_), .C(men_men_n29_), .D(m), .Y(men_men_n902_));
  NOi21      u0874(.An(men_men_n326_), .B(men_men_n902_), .Y(men_men_n903_));
  AOI210     u0875(.A0(men_men_n900_), .A1(men_men_n568_), .B0(men_men_n903_), .Y(men_men_n904_));
  AN2        u0876(.A(f), .B(d), .Y(men_men_n905_));
  NA3        u0877(.A(men_men_n498_), .B(men_men_n905_), .C(men_men_n86_), .Y(men_men_n906_));
  NO3        u0878(.A(men_men_n906_), .B(men_men_n75_), .C(men_men_n223_), .Y(men_men_n907_));
  NO2        u0879(.A(men_men_n297_), .B(men_men_n56_), .Y(men_men_n908_));
  NAi21      u0880(.An(men_men_n510_), .B(men_men_n904_), .Y(men_men_n909_));
  NO4        u0881(.A(men_men_n649_), .B(men_men_n137_), .C(men_men_n344_), .D(men_men_n156_), .Y(men_men_n910_));
  NO2        u0882(.A(men_men_n683_), .B(men_men_n344_), .Y(men_men_n911_));
  AN2        u0883(.A(men_men_n911_), .B(men_men_n710_), .Y(men_men_n912_));
  NO3        u0884(.A(men_men_n912_), .B(men_men_n910_), .C(men_men_n244_), .Y(men_men_n913_));
  NA2        u0885(.A(men_men_n627_), .B(men_men_n86_), .Y(men_men_n914_));
  NO2        u0886(.A(men_men_n890_), .B(men_men_n914_), .Y(men_men_n915_));
  NA3        u0887(.A(men_men_n164_), .B(men_men_n112_), .C(men_men_n111_), .Y(men_men_n916_));
  OAI220     u0888(.A0(men_men_n906_), .A1(men_men_n451_), .B0(men_men_n356_), .B1(men_men_n916_), .Y(men_men_n917_));
  NOi41      u0889(.An(men_men_n233_), .B(men_men_n917_), .C(men_men_n915_), .D(men_men_n320_), .Y(men_men_n918_));
  NA2        u0890(.A(c), .B(men_men_n120_), .Y(men_men_n919_));
  NO2        u0891(.A(men_men_n919_), .B(men_men_n430_), .Y(men_men_n920_));
  NA3        u0892(.A(men_men_n920_), .B(men_men_n532_), .C(f), .Y(men_men_n921_));
  OR2        u0893(.A(men_men_n690_), .B(men_men_n564_), .Y(men_men_n922_));
  INV        u0894(.A(men_men_n922_), .Y(men_men_n923_));
  NA2        u0895(.A(men_men_n841_), .B(men_men_n115_), .Y(men_men_n924_));
  NA2        u0896(.A(men_men_n924_), .B(men_men_n923_), .Y(men_men_n925_));
  NA4        u0897(.A(men_men_n925_), .B(men_men_n921_), .C(men_men_n918_), .D(men_men_n913_), .Y(men_men_n926_));
  NO4        u0898(.A(men_men_n926_), .B(men_men_n909_), .C(men_men_n896_), .D(men_men_n883_), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n116_), .B(j), .Y(men_men_n928_));
  NO2        u0900(.A(men_men_n349_), .B(men_men_n879_), .Y(men_men_n929_));
  NO2        u0901(.A(men_men_n240_), .B(men_men_n234_), .Y(men_men_n930_));
  NA2        u0902(.A(men_men_n930_), .B(men_men_n237_), .Y(men_men_n931_));
  NO2        u0903(.A(men_men_n451_), .B(men_men_n867_), .Y(men_men_n932_));
  NA2        u0904(.A(men_men_n932_), .B(men_men_n585_), .Y(men_men_n933_));
  NA2        u0905(.A(men_men_n933_), .B(men_men_n931_), .Y(men_men_n934_));
  NA2        u0906(.A(e), .B(d), .Y(men_men_n935_));
  OAI220     u0907(.A0(men_men_n935_), .A1(c), .B0(men_men_n339_), .B1(d), .Y(men_men_n936_));
  NA3        u0908(.A(men_men_n936_), .B(men_men_n474_), .C(men_men_n530_), .Y(men_men_n937_));
  AOI210     u0909(.A0(men_men_n537_), .A1(men_men_n187_), .B0(men_men_n240_), .Y(men_men_n938_));
  AOI210     u0910(.A0(men_men_n650_), .A1(men_men_n365_), .B0(men_men_n938_), .Y(men_men_n939_));
  NA2        u0911(.A(men_men_n297_), .B(men_men_n170_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n907_), .B(men_men_n940_), .Y(men_men_n941_));
  NA3        u0913(.A(men_men_n173_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n942_));
  NA4        u0914(.A(men_men_n942_), .B(men_men_n941_), .C(men_men_n939_), .D(men_men_n937_), .Y(men_men_n943_));
  NO3        u0915(.A(men_men_n943_), .B(men_men_n934_), .C(men_men_n929_), .Y(men_men_n944_));
  NA2        u0916(.A(men_men_n884_), .B(men_men_n31_), .Y(men_men_n945_));
  AO210      u0917(.A0(men_men_n945_), .A1(men_men_n728_), .B0(men_men_n226_), .Y(men_men_n946_));
  OAI220     u0918(.A0(men_men_n649_), .A1(men_men_n61_), .B0(men_men_n313_), .B1(j), .Y(men_men_n947_));
  AOI220     u0919(.A0(men_men_n947_), .A1(men_men_n911_), .B0(men_men_n639_), .B1(men_men_n648_), .Y(men_men_n948_));
  OAI210     u0920(.A0(men_men_n873_), .A1(men_men_n177_), .B0(men_men_n948_), .Y(men_men_n949_));
  OAI210     u0921(.A0(men_men_n868_), .A1(men_men_n940_), .B0(men_men_n901_), .Y(men_men_n950_));
  NO2        u0922(.A(men_men_n950_), .B(men_men_n630_), .Y(men_men_n951_));
  AOI210     u0923(.A0(men_men_n122_), .A1(men_men_n121_), .B0(men_men_n272_), .Y(men_men_n952_));
  NO2        u0924(.A(men_men_n952_), .B(men_men_n902_), .Y(men_men_n953_));
  AO210      u0925(.A0(men_men_n889_), .A1(men_men_n878_), .B0(men_men_n953_), .Y(men_men_n954_));
  NOi31      u0926(.An(men_men_n568_), .B(men_men_n899_), .C(men_men_n305_), .Y(men_men_n955_));
  NO4        u0927(.A(men_men_n955_), .B(men_men_n954_), .C(men_men_n951_), .D(men_men_n949_), .Y(men_men_n956_));
  AO220      u0928(.A0(men_men_n474_), .A1(men_men_n781_), .B0(men_men_n182_), .B1(f), .Y(men_men_n957_));
  OAI210     u0929(.A0(men_men_n957_), .A1(men_men_n477_), .B0(men_men_n936_), .Y(men_men_n958_));
  NO2        u0930(.A(men_men_n461_), .B(men_men_n71_), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n882_), .A1(men_men_n959_), .B0(men_men_n732_), .Y(men_men_n960_));
  AN4        u0932(.A(men_men_n960_), .B(men_men_n958_), .C(men_men_n956_), .D(men_men_n946_), .Y(men_men_n961_));
  NA4        u0933(.A(men_men_n961_), .B(men_men_n944_), .C(men_men_n927_), .D(men_men_n875_), .Y(men12));
  NO2        u0934(.A(men_men_n472_), .B(c), .Y(men_men_n963_));
  NO4        u0935(.A(men_men_n464_), .B(men_men_n264_), .C(men_men_n606_), .D(men_men_n223_), .Y(men_men_n964_));
  NA2        u0936(.A(men_men_n964_), .B(men_men_n963_), .Y(men_men_n965_));
  NA2        u0937(.A(men_men_n568_), .B(men_men_n959_), .Y(men_men_n966_));
  NO2        u0938(.A(men_men_n472_), .B(men_men_n120_), .Y(men_men_n967_));
  NO2        u0939(.A(men_men_n885_), .B(men_men_n372_), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n690_), .B(men_men_n399_), .Y(men_men_n969_));
  AOI220     u0941(.A0(men_men_n969_), .A1(men_men_n566_), .B0(men_men_n968_), .B1(men_men_n967_), .Y(men_men_n970_));
  NA4        u0942(.A(men_men_n970_), .B(men_men_n966_), .C(men_men_n965_), .D(men_men_n463_), .Y(men_men_n971_));
  AOI210     u0943(.A0(men_men_n243_), .A1(men_men_n355_), .B0(men_men_n209_), .Y(men_men_n972_));
  OR2        u0944(.A(men_men_n972_), .B(men_men_n964_), .Y(men_men_n973_));
  AOI210     u0945(.A0(men_men_n352_), .A1(men_men_n411_), .B0(men_men_n223_), .Y(men_men_n974_));
  OAI210     u0946(.A0(men_men_n974_), .A1(men_men_n973_), .B0(men_men_n425_), .Y(men_men_n975_));
  NO2        u0947(.A(men_men_n669_), .B(men_men_n275_), .Y(men_men_n976_));
  NO2        u0948(.A(men_men_n613_), .B(men_men_n877_), .Y(men_men_n977_));
  AOI220     u0949(.A0(men_men_n977_), .A1(men_men_n591_), .B0(men_men_n852_), .B1(men_men_n976_), .Y(men_men_n978_));
  NO2        u0950(.A(men_men_n155_), .B(men_men_n247_), .Y(men_men_n979_));
  NA3        u0951(.A(men_men_n979_), .B(men_men_n250_), .C(i), .Y(men_men_n980_));
  NA3        u0952(.A(men_men_n980_), .B(men_men_n978_), .C(men_men_n975_), .Y(men_men_n981_));
  OR2        u0953(.A(men_men_n340_), .B(men_men_n967_), .Y(men_men_n982_));
  NA2        u0954(.A(men_men_n982_), .B(men_men_n373_), .Y(men_men_n983_));
  NA4        u0955(.A(men_men_n465_), .B(men_men_n459_), .C(men_men_n188_), .D(g), .Y(men_men_n984_));
  NA2        u0956(.A(men_men_n984_), .B(men_men_n983_), .Y(men_men_n985_));
  NO3        u0957(.A(men_men_n695_), .B(men_men_n94_), .C(men_men_n45_), .Y(men_men_n986_));
  NO4        u0958(.A(men_men_n986_), .B(men_men_n985_), .C(men_men_n981_), .D(men_men_n971_), .Y(men_men_n987_));
  NO2        u0959(.A(men_men_n389_), .B(men_men_n388_), .Y(men_men_n988_));
  INV        u0960(.A(men_men_n610_), .Y(men_men_n989_));
  NA2        u0961(.A(men_men_n578_), .B(men_men_n149_), .Y(men_men_n990_));
  NOi21      u0962(.An(men_men_n34_), .B(men_men_n683_), .Y(men_men_n991_));
  AOI220     u0963(.A0(men_men_n991_), .A1(men_men_n990_), .B0(men_men_n989_), .B1(men_men_n988_), .Y(men_men_n992_));
  OAI210     u0964(.A0(men_men_n262_), .A1(men_men_n45_), .B0(men_men_n992_), .Y(men_men_n993_));
  NA2        u0965(.A(men_men_n457_), .B(men_men_n277_), .Y(men_men_n994_));
  NO3        u0966(.A(men_men_n854_), .B(men_men_n91_), .C(men_men_n430_), .Y(men_men_n995_));
  NAi31      u0967(.An(men_men_n995_), .B(men_men_n994_), .C(men_men_n336_), .Y(men_men_n996_));
  NO2        u0968(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n997_));
  NO2        u0969(.A(men_men_n526_), .B(men_men_n313_), .Y(men_men_n998_));
  NO2        u0970(.A(men_men_n998_), .B(men_men_n385_), .Y(men_men_n999_));
  NO2        u0971(.A(men_men_n999_), .B(men_men_n149_), .Y(men_men_n1000_));
  NA2        u0972(.A(men_men_n660_), .B(men_men_n382_), .Y(men_men_n1001_));
  OAI210     u0973(.A0(men_men_n768_), .A1(men_men_n1001_), .B0(men_men_n386_), .Y(men_men_n1002_));
  NO4        u0974(.A(men_men_n1002_), .B(men_men_n1000_), .C(men_men_n996_), .D(men_men_n993_), .Y(men_men_n1003_));
  NA2        u0975(.A(men_men_n365_), .B(g), .Y(men_men_n1004_));
  NA2        u0976(.A(men_men_n167_), .B(i), .Y(men_men_n1005_));
  NA2        u0977(.A(men_men_n46_), .B(i), .Y(men_men_n1006_));
  OAI220     u0978(.A0(men_men_n1006_), .A1(men_men_n208_), .B0(men_men_n1005_), .B1(men_men_n94_), .Y(men_men_n1007_));
  AOI210     u0979(.A0(men_men_n441_), .A1(men_men_n37_), .B0(men_men_n1007_), .Y(men_men_n1008_));
  NA2        u0980(.A(men_men_n578_), .B(men_men_n403_), .Y(men_men_n1009_));
  AOI210     u0981(.A0(men_men_n1009_), .A1(n), .B0(men_men_n577_), .Y(men_men_n1010_));
  OAI220     u0982(.A0(men_men_n1010_), .A1(men_men_n1004_), .B0(men_men_n1008_), .B1(men_men_n349_), .Y(men_men_n1011_));
  NO2        u0983(.A(men_men_n690_), .B(men_men_n519_), .Y(men_men_n1012_));
  NA3        u0984(.A(men_men_n360_), .B(men_men_n655_), .C(i), .Y(men_men_n1013_));
  OAI210     u0985(.A0(men_men_n461_), .A1(men_men_n325_), .B0(men_men_n1013_), .Y(men_men_n1014_));
  OAI210     u0986(.A0(men_men_n1014_), .A1(men_men_n1012_), .B0(men_men_n793_), .Y(men_men_n1015_));
  NA2        u0987(.A(men_men_n633_), .B(men_men_n117_), .Y(men_men_n1016_));
  OR3        u0988(.A(men_men_n325_), .B(men_men_n456_), .C(f), .Y(men_men_n1017_));
  NA3        u0989(.A(men_men_n655_), .B(men_men_n82_), .C(i), .Y(men_men_n1018_));
  OA220      u0990(.A0(men_men_n1018_), .A1(men_men_n1016_), .B0(men_men_n1017_), .B1(men_men_n612_), .Y(men_men_n1019_));
  NA3        u0991(.A(men_men_n341_), .B(men_men_n122_), .C(g), .Y(men_men_n1020_));
  AOI210     u0992(.A0(men_men_n705_), .A1(men_men_n1020_), .B0(m), .Y(men_men_n1021_));
  OAI210     u0993(.A0(men_men_n1021_), .A1(men_men_n968_), .B0(men_men_n340_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n721_), .B(men_men_n914_), .Y(men_men_n1023_));
  NA2        u0995(.A(men_men_n879_), .B(men_men_n462_), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n231_), .B(men_men_n79_), .Y(men_men_n1025_));
  NA3        u0997(.A(men_men_n1025_), .B(men_men_n1018_), .C(men_men_n1017_), .Y(men_men_n1026_));
  AOI220     u0998(.A0(men_men_n1026_), .A1(men_men_n270_), .B0(men_men_n1024_), .B1(men_men_n1023_), .Y(men_men_n1027_));
  NA4        u0999(.A(men_men_n1027_), .B(men_men_n1022_), .C(men_men_n1019_), .D(men_men_n1015_), .Y(men_men_n1028_));
  NO2        u1000(.A(men_men_n399_), .B(men_men_n93_), .Y(men_men_n1029_));
  OAI210     u1001(.A0(men_men_n1029_), .A1(men_men_n976_), .B0(men_men_n248_), .Y(men_men_n1030_));
  NA2        u1002(.A(men_men_n694_), .B(men_men_n90_), .Y(men_men_n1031_));
  NO2        u1003(.A(men_men_n480_), .B(men_men_n223_), .Y(men_men_n1032_));
  AOI220     u1004(.A0(men_men_n1032_), .A1(men_men_n404_), .B0(men_men_n982_), .B1(men_men_n227_), .Y(men_men_n1033_));
  AOI220     u1005(.A0(men_men_n969_), .A1(men_men_n979_), .B0(men_men_n611_), .B1(men_men_n92_), .Y(men_men_n1034_));
  NA4        u1006(.A(men_men_n1034_), .B(men_men_n1033_), .C(men_men_n1031_), .D(men_men_n1030_), .Y(men_men_n1035_));
  NA2        u1007(.A(men_men_n1024_), .B(men_men_n566_), .Y(men_men_n1036_));
  AOI210     u1008(.A0(men_men_n442_), .A1(men_men_n434_), .B0(men_men_n854_), .Y(men_men_n1037_));
  OAI210     u1009(.A0(men_men_n389_), .A1(men_men_n388_), .B0(men_men_n113_), .Y(men_men_n1038_));
  AOI210     u1010(.A0(men_men_n1038_), .A1(men_men_n558_), .B0(men_men_n1037_), .Y(men_men_n1039_));
  NA2        u1011(.A(men_men_n1021_), .B(men_men_n967_), .Y(men_men_n1040_));
  NO3        u1012(.A(men_men_n928_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1041_));
  AOI220     u1013(.A0(men_men_n1041_), .A1(men_men_n653_), .B0(men_men_n674_), .B1(men_men_n553_), .Y(men_men_n1042_));
  NA4        u1014(.A(men_men_n1042_), .B(men_men_n1040_), .C(men_men_n1039_), .D(men_men_n1036_), .Y(men_men_n1043_));
  NO4        u1015(.A(men_men_n1043_), .B(men_men_n1035_), .C(men_men_n1028_), .D(men_men_n1011_), .Y(men_men_n1044_));
  NAi31      u1016(.An(men_men_n146_), .B(men_men_n443_), .C(n), .Y(men_men_n1045_));
  NO3        u1017(.A(men_men_n130_), .B(men_men_n358_), .C(men_men_n886_), .Y(men_men_n1046_));
  NO2        u1018(.A(men_men_n1046_), .B(men_men_n1045_), .Y(men_men_n1047_));
  NO3        u1019(.A(men_men_n285_), .B(men_men_n146_), .C(men_men_n430_), .Y(men_men_n1048_));
  AOI210     u1020(.A0(men_men_n1048_), .A1(men_men_n520_), .B0(men_men_n1047_), .Y(men_men_n1049_));
  INV        u1021(.A(men_men_n1049_), .Y(men_men_n1050_));
  NA2        u1022(.A(men_men_n240_), .B(men_men_n178_), .Y(men_men_n1051_));
  NO3        u1023(.A(men_men_n322_), .B(men_men_n465_), .C(men_men_n182_), .Y(men_men_n1052_));
  NOi31      u1024(.An(men_men_n1051_), .B(men_men_n1052_), .C(men_men_n223_), .Y(men_men_n1053_));
  NAi21      u1025(.An(men_men_n578_), .B(men_men_n1032_), .Y(men_men_n1054_));
  NA2        u1026(.A(men_men_n460_), .B(men_men_n914_), .Y(men_men_n1055_));
  NO3        u1027(.A(men_men_n461_), .B(men_men_n325_), .C(men_men_n75_), .Y(men_men_n1056_));
  AOI220     u1028(.A0(men_men_n1056_), .A1(men_men_n1055_), .B0(men_men_n502_), .B1(g), .Y(men_men_n1057_));
  NA2        u1029(.A(men_men_n1057_), .B(men_men_n1054_), .Y(men_men_n1058_));
  OAI220     u1030(.A0(men_men_n1045_), .A1(men_men_n243_), .B0(men_men_n1013_), .B1(men_men_n628_), .Y(men_men_n1059_));
  NO2        u1031(.A(men_men_n691_), .B(men_men_n399_), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n972_), .B(men_men_n963_), .Y(men_men_n1061_));
  NO3        u1033(.A(men_men_n567_), .B(men_men_n153_), .C(men_men_n222_), .Y(men_men_n1062_));
  OAI210     u1034(.A0(men_men_n1062_), .A1(men_men_n547_), .B0(men_men_n400_), .Y(men_men_n1063_));
  OAI220     u1035(.A0(men_men_n969_), .A1(men_men_n977_), .B0(men_men_n568_), .B1(men_men_n450_), .Y(men_men_n1064_));
  NA4        u1036(.A(men_men_n1064_), .B(men_men_n1063_), .C(men_men_n1061_), .D(men_men_n647_), .Y(men_men_n1065_));
  OAI210     u1037(.A0(men_men_n972_), .A1(men_men_n964_), .B0(men_men_n1051_), .Y(men_men_n1066_));
  NA3        u1038(.A(men_men_n1009_), .B(men_men_n507_), .C(men_men_n46_), .Y(men_men_n1067_));
  AOI210     u1039(.A0(men_men_n402_), .A1(men_men_n400_), .B0(men_men_n348_), .Y(men_men_n1068_));
  NA4        u1040(.A(men_men_n1068_), .B(men_men_n1067_), .C(men_men_n1066_), .D(men_men_n286_), .Y(men_men_n1069_));
  OR4        u1041(.A(men_men_n1069_), .B(men_men_n1065_), .C(men_men_n1060_), .D(men_men_n1059_), .Y(men_men_n1070_));
  NO4        u1042(.A(men_men_n1070_), .B(men_men_n1058_), .C(men_men_n1053_), .D(men_men_n1050_), .Y(men_men_n1071_));
  NA4        u1043(.A(men_men_n1071_), .B(men_men_n1044_), .C(men_men_n1003_), .D(men_men_n987_), .Y(men13));
  NA2        u1044(.A(men_men_n46_), .B(men_men_n89_), .Y(men_men_n1073_));
  AN2        u1045(.A(c), .B(b), .Y(men_men_n1074_));
  NA3        u1046(.A(men_men_n261_), .B(men_men_n1074_), .C(m), .Y(men_men_n1075_));
  NA2        u1047(.A(men_men_n517_), .B(f), .Y(men_men_n1076_));
  NO4        u1048(.A(men_men_n1076_), .B(men_men_n1075_), .C(men_men_n1073_), .D(men_men_n607_), .Y(men_men_n1077_));
  NA2        u1049(.A(men_men_n277_), .B(men_men_n1074_), .Y(men_men_n1078_));
  NO4        u1050(.A(men_men_n1078_), .B(men_men_n1076_), .C(men_men_n1005_), .D(a), .Y(men_men_n1079_));
  NAi32      u1051(.An(d), .Bn(c), .C(e), .Y(men_men_n1080_));
  NA2        u1052(.A(men_men_n145_), .B(men_men_n45_), .Y(men_men_n1081_));
  NO4        u1053(.A(men_men_n1081_), .B(men_men_n1080_), .C(men_men_n613_), .D(men_men_n321_), .Y(men_men_n1082_));
  NA2        u1054(.A(men_men_n433_), .B(men_men_n222_), .Y(men_men_n1083_));
  AN2        u1055(.A(d), .B(c), .Y(men_men_n1084_));
  NA2        u1056(.A(men_men_n1084_), .B(men_men_n120_), .Y(men_men_n1085_));
  NO4        u1057(.A(men_men_n1085_), .B(men_men_n1083_), .C(men_men_n183_), .D(men_men_n174_), .Y(men_men_n1086_));
  NA2        u1058(.A(men_men_n517_), .B(c), .Y(men_men_n1087_));
  NO4        u1059(.A(men_men_n1081_), .B(men_men_n609_), .C(men_men_n1087_), .D(men_men_n321_), .Y(men_men_n1088_));
  OR2        u1060(.A(men_men_n1086_), .B(men_men_n1088_), .Y(men_men_n1089_));
  OR4        u1061(.A(men_men_n1089_), .B(men_men_n1082_), .C(men_men_n1079_), .D(men_men_n1077_), .Y(men_men_n1090_));
  NAi32      u1062(.An(f), .Bn(e), .C(c), .Y(men_men_n1091_));
  NO2        u1063(.A(men_men_n1091_), .B(men_men_n150_), .Y(men_men_n1092_));
  NA2        u1064(.A(men_men_n1092_), .B(g), .Y(men_men_n1093_));
  OR3        u1065(.A(men_men_n234_), .B(men_men_n183_), .C(men_men_n174_), .Y(men_men_n1094_));
  NO2        u1066(.A(men_men_n1094_), .B(men_men_n1093_), .Y(men_men_n1095_));
  NO2        u1067(.A(men_men_n1087_), .B(men_men_n321_), .Y(men_men_n1096_));
  NO2        u1068(.A(j), .B(men_men_n45_), .Y(men_men_n1097_));
  NA2        u1069(.A(men_men_n657_), .B(men_men_n1097_), .Y(men_men_n1098_));
  NOi21      u1070(.An(men_men_n1096_), .B(men_men_n1098_), .Y(men_men_n1099_));
  NO2        u1071(.A(men_men_n797_), .B(men_men_n116_), .Y(men_men_n1100_));
  NOi41      u1072(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1101_));
  NA2        u1073(.A(men_men_n1101_), .B(men_men_n1100_), .Y(men_men_n1102_));
  NO2        u1074(.A(men_men_n1102_), .B(men_men_n1093_), .Y(men_men_n1103_));
  OR3        u1075(.A(e), .B(d), .C(c), .Y(men_men_n1104_));
  NA3        u1076(.A(k), .B(j), .C(i), .Y(men_men_n1105_));
  NO3        u1077(.A(men_men_n1105_), .B(men_men_n321_), .C(men_men_n93_), .Y(men_men_n1106_));
  NOi21      u1078(.An(men_men_n1106_), .B(men_men_n1104_), .Y(men_men_n1107_));
  OR4        u1079(.A(men_men_n1107_), .B(men_men_n1103_), .C(men_men_n1099_), .D(men_men_n1095_), .Y(men_men_n1108_));
  NA3        u1080(.A(men_men_n488_), .B(men_men_n351_), .C(men_men_n56_), .Y(men_men_n1109_));
  NO2        u1081(.A(men_men_n1109_), .B(men_men_n1098_), .Y(men_men_n1110_));
  NO3        u1082(.A(men_men_n1109_), .B(men_men_n609_), .C(men_men_n471_), .Y(men_men_n1111_));
  NO2        u1083(.A(f), .B(c), .Y(men_men_n1112_));
  NOi21      u1084(.An(men_men_n1112_), .B(men_men_n464_), .Y(men_men_n1113_));
  NA2        u1085(.A(men_men_n1113_), .B(men_men_n59_), .Y(men_men_n1114_));
  OR2        u1086(.A(k), .B(i), .Y(men_men_n1115_));
  NO3        u1087(.A(men_men_n1115_), .B(men_men_n254_), .C(l), .Y(men_men_n1116_));
  NOi31      u1088(.An(men_men_n1116_), .B(men_men_n1114_), .C(j), .Y(men_men_n1117_));
  OR3        u1089(.A(men_men_n1117_), .B(men_men_n1111_), .C(men_men_n1110_), .Y(men_men_n1118_));
  OR3        u1090(.A(men_men_n1118_), .B(men_men_n1108_), .C(men_men_n1090_), .Y(men02));
  OR2        u1091(.A(l), .B(k), .Y(men_men_n1120_));
  OR3        u1092(.A(h), .B(g), .C(f), .Y(men_men_n1121_));
  OR3        u1093(.A(n), .B(m), .C(i), .Y(men_men_n1122_));
  NO4        u1094(.A(men_men_n1122_), .B(men_men_n1121_), .C(men_men_n1120_), .D(men_men_n1104_), .Y(men_men_n1123_));
  NOi31      u1095(.An(e), .B(d), .C(c), .Y(men_men_n1124_));
  AOI210     u1096(.A0(men_men_n1106_), .A1(men_men_n1124_), .B0(men_men_n1082_), .Y(men_men_n1125_));
  AN3        u1097(.A(g), .B(f), .C(c), .Y(men_men_n1126_));
  NA3        u1098(.A(men_men_n1126_), .B(men_men_n488_), .C(h), .Y(men_men_n1127_));
  OR2        u1099(.A(men_men_n1105_), .B(men_men_n321_), .Y(men_men_n1128_));
  OR2        u1100(.A(men_men_n1128_), .B(men_men_n1127_), .Y(men_men_n1129_));
  NO3        u1101(.A(men_men_n1109_), .B(men_men_n1081_), .C(men_men_n609_), .Y(men_men_n1130_));
  NO2        u1102(.A(men_men_n1130_), .B(men_men_n1095_), .Y(men_men_n1131_));
  NA3        u1103(.A(l), .B(k), .C(j), .Y(men_men_n1132_));
  NA2        u1104(.A(i), .B(h), .Y(men_men_n1133_));
  NO3        u1105(.A(men_men_n1133_), .B(men_men_n1132_), .C(men_men_n137_), .Y(men_men_n1134_));
  NO3        u1106(.A(men_men_n147_), .B(men_men_n295_), .C(men_men_n223_), .Y(men_men_n1135_));
  AOI210     u1107(.A0(men_men_n1135_), .A1(men_men_n1134_), .B0(men_men_n1099_), .Y(men_men_n1136_));
  NA3        u1108(.A(c), .B(b), .C(a), .Y(men_men_n1137_));
  NO3        u1109(.A(men_men_n1137_), .B(men_men_n935_), .C(men_men_n222_), .Y(men_men_n1138_));
  NO4        u1110(.A(men_men_n1105_), .B(men_men_n313_), .C(men_men_n49_), .D(men_men_n116_), .Y(men_men_n1139_));
  AOI210     u1111(.A0(men_men_n1139_), .A1(men_men_n1138_), .B0(men_men_n1110_), .Y(men_men_n1140_));
  AN4        u1112(.A(men_men_n1140_), .B(men_men_n1136_), .C(men_men_n1131_), .D(men_men_n1129_), .Y(men_men_n1141_));
  NO2        u1113(.A(men_men_n1085_), .B(men_men_n1083_), .Y(men_men_n1142_));
  NA2        u1114(.A(men_men_n1102_), .B(men_men_n1094_), .Y(men_men_n1143_));
  AOI210     u1115(.A0(men_men_n1143_), .A1(men_men_n1142_), .B0(men_men_n1077_), .Y(men_men_n1144_));
  NAi41      u1116(.An(men_men_n1123_), .B(men_men_n1144_), .C(men_men_n1141_), .D(men_men_n1125_), .Y(men03));
  NO2        u1117(.A(men_men_n549_), .B(men_men_n622_), .Y(men_men_n1146_));
  NA4        u1118(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(men_men_n222_), .Y(men_men_n1147_));
  NA4        u1119(.A(men_men_n599_), .B(m), .C(men_men_n116_), .D(men_men_n222_), .Y(men_men_n1148_));
  NA3        u1120(.A(men_men_n1148_), .B(men_men_n390_), .C(men_men_n1147_), .Y(men_men_n1149_));
  NO3        u1121(.A(men_men_n1149_), .B(men_men_n1146_), .C(men_men_n1038_), .Y(men_men_n1150_));
  NO3        u1122(.A(men_men_n891_), .B(men_men_n880_), .C(men_men_n746_), .Y(men_men_n1151_));
  OAI220     u1123(.A0(men_men_n1151_), .A1(men_men_n721_), .B0(men_men_n1150_), .B1(men_men_n610_), .Y(men_men_n1152_));
  NOi31      u1124(.An(i), .B(k), .C(j), .Y(men_men_n1153_));
  NA4        u1125(.A(men_men_n1153_), .B(men_men_n1124_), .C(men_men_n360_), .D(men_men_n351_), .Y(men_men_n1154_));
  OAI210     u1126(.A0(men_men_n854_), .A1(men_men_n444_), .B0(men_men_n1154_), .Y(men_men_n1155_));
  NOi31      u1127(.An(m), .B(n), .C(f), .Y(men_men_n1156_));
  NA2        u1128(.A(men_men_n1156_), .B(men_men_n51_), .Y(men_men_n1157_));
  AN2        u1129(.A(e), .B(c), .Y(men_men_n1158_));
  NO2        u1130(.A(men_men_n922_), .B(men_men_n449_), .Y(men_men_n1159_));
  NA2        u1131(.A(men_men_n530_), .B(l), .Y(men_men_n1160_));
  NOi31      u1132(.An(men_men_n901_), .B(men_men_n1075_), .C(men_men_n1160_), .Y(men_men_n1161_));
  NO4        u1133(.A(men_men_n1161_), .B(men_men_n1159_), .C(men_men_n1155_), .D(men_men_n1037_), .Y(men_men_n1162_));
  NO2        u1134(.A(men_men_n295_), .B(a), .Y(men_men_n1163_));
  INV        u1135(.A(men_men_n1082_), .Y(men_men_n1164_));
  NO2        u1136(.A(men_men_n1133_), .B(men_men_n505_), .Y(men_men_n1165_));
  NO2        u1137(.A(men_men_n89_), .B(g), .Y(men_men_n1166_));
  AOI210     u1138(.A0(men_men_n1166_), .A1(men_men_n1165_), .B0(men_men_n1116_), .Y(men_men_n1167_));
  OR2        u1139(.A(men_men_n1167_), .B(men_men_n1114_), .Y(men_men_n1168_));
  NA3        u1140(.A(men_men_n1168_), .B(men_men_n1164_), .C(men_men_n1162_), .Y(men_men_n1169_));
  NO4        u1141(.A(men_men_n1169_), .B(men_men_n1152_), .C(men_men_n856_), .D(men_men_n590_), .Y(men_men_n1170_));
  NA2        u1142(.A(c), .B(b), .Y(men_men_n1171_));
  NO2        u1143(.A(men_men_n731_), .B(men_men_n1171_), .Y(men_men_n1172_));
  OAI210     u1144(.A0(men_men_n899_), .A1(men_men_n871_), .B0(men_men_n437_), .Y(men_men_n1173_));
  OAI210     u1145(.A0(men_men_n1173_), .A1(men_men_n900_), .B0(men_men_n1172_), .Y(men_men_n1174_));
  NAi21      u1146(.An(men_men_n445_), .B(men_men_n1172_), .Y(men_men_n1175_));
  OAI210     u1147(.A0(men_men_n572_), .A1(men_men_n39_), .B0(men_men_n1163_), .Y(men_men_n1176_));
  NA2        u1148(.A(men_men_n1176_), .B(men_men_n1175_), .Y(men_men_n1177_));
  INV        u1149(.A(men_men_n273_), .Y(men_men_n1178_));
  OAI210     u1150(.A0(men_men_n1178_), .A1(men_men_n299_), .B0(g), .Y(men_men_n1179_));
  NAi21      u1151(.An(f), .B(d), .Y(men_men_n1180_));
  NO2        u1152(.A(men_men_n1180_), .B(men_men_n1137_), .Y(men_men_n1181_));
  INV        u1153(.A(men_men_n1181_), .Y(men_men_n1182_));
  AOI210     u1154(.A0(men_men_n1179_), .A1(men_men_n305_), .B0(men_men_n1182_), .Y(men_men_n1183_));
  AOI210     u1155(.A0(men_men_n1183_), .A1(men_men_n117_), .B0(men_men_n1177_), .Y(men_men_n1184_));
  NA2        u1156(.A(men_men_n490_), .B(men_men_n489_), .Y(men_men_n1185_));
  NO2        u1157(.A(men_men_n189_), .B(men_men_n247_), .Y(men_men_n1186_));
  NA2        u1158(.A(men_men_n1186_), .B(m), .Y(men_men_n1187_));
  NA3        u1159(.A(men_men_n952_), .B(men_men_n1160_), .C(men_men_n493_), .Y(men_men_n1188_));
  OAI210     u1160(.A0(men_men_n1188_), .A1(men_men_n326_), .B0(men_men_n491_), .Y(men_men_n1189_));
  AOI210     u1161(.A0(men_men_n1189_), .A1(men_men_n1185_), .B0(men_men_n1187_), .Y(men_men_n1190_));
  NA2        u1162(.A(men_men_n585_), .B(men_men_n432_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n163_), .B(men_men_n33_), .Y(men_men_n1192_));
  AOI210     u1164(.A0(men_men_n1001_), .A1(men_men_n1192_), .B0(men_men_n223_), .Y(men_men_n1193_));
  OAI210     u1165(.A0(men_men_n1193_), .A1(men_men_n468_), .B0(men_men_n1181_), .Y(men_men_n1194_));
  NO2        u1166(.A(men_men_n393_), .B(men_men_n392_), .Y(men_men_n1195_));
  AOI210     u1167(.A0(men_men_n1186_), .A1(men_men_n452_), .B0(men_men_n995_), .Y(men_men_n1196_));
  NAi41      u1168(.An(men_men_n1195_), .B(men_men_n1196_), .C(men_men_n1194_), .D(men_men_n1191_), .Y(men_men_n1197_));
  NO2        u1169(.A(men_men_n1197_), .B(men_men_n1190_), .Y(men_men_n1198_));
  NA4        u1170(.A(men_men_n1198_), .B(men_men_n1184_), .C(men_men_n1174_), .D(men_men_n1170_), .Y(men00));
  AOI210     u1171(.A0(men_men_n312_), .A1(men_men_n223_), .B0(men_men_n288_), .Y(men_men_n1200_));
  NO2        u1172(.A(men_men_n1200_), .B(men_men_n602_), .Y(men_men_n1201_));
  AOI210     u1173(.A0(men_men_n932_), .A1(men_men_n979_), .B0(men_men_n1155_), .Y(men_men_n1202_));
  NO3        u1174(.A(men_men_n1130_), .B(men_men_n995_), .C(men_men_n743_), .Y(men_men_n1203_));
  NA3        u1175(.A(men_men_n1203_), .B(men_men_n1202_), .C(men_men_n1039_), .Y(men_men_n1204_));
  NA2        u1176(.A(men_men_n532_), .B(f), .Y(men_men_n1205_));
  OAI210     u1177(.A0(men_men_n1046_), .A1(men_men_n40_), .B0(men_men_n676_), .Y(men_men_n1206_));
  NA3        u1178(.A(men_men_n1206_), .B(men_men_n269_), .C(n), .Y(men_men_n1207_));
  AOI210     u1179(.A0(men_men_n1207_), .A1(men_men_n1205_), .B0(men_men_n1085_), .Y(men_men_n1208_));
  NO4        u1180(.A(men_men_n1208_), .B(men_men_n1204_), .C(men_men_n1201_), .D(men_men_n1108_), .Y(men_men_n1209_));
  NA3        u1181(.A(men_men_n173_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1210_));
  NA3        u1182(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1211_));
  NOi31      u1183(.An(n), .B(m), .C(i), .Y(men_men_n1212_));
  NA3        u1184(.A(men_men_n1212_), .B(men_men_n679_), .C(men_men_n51_), .Y(men_men_n1213_));
  OAI210     u1185(.A0(men_men_n1211_), .A1(men_men_n1210_), .B0(men_men_n1213_), .Y(men_men_n1214_));
  INV        u1186(.A(men_men_n601_), .Y(men_men_n1215_));
  NO4        u1187(.A(men_men_n1215_), .B(men_men_n1214_), .C(men_men_n1195_), .D(men_men_n955_), .Y(men_men_n1216_));
  NO4        u1188(.A(men_men_n508_), .B(men_men_n375_), .C(men_men_n1171_), .D(men_men_n59_), .Y(men_men_n1217_));
  NA3        u1189(.A(men_men_n405_), .B(men_men_n230_), .C(g), .Y(men_men_n1218_));
  OA220      u1190(.A0(men_men_n1218_), .A1(men_men_n1211_), .B0(men_men_n406_), .B1(men_men_n140_), .Y(men_men_n1219_));
  NO2        u1191(.A(h), .B(g), .Y(men_men_n1220_));
  NA4        u1192(.A(men_men_n520_), .B(men_men_n488_), .C(men_men_n1220_), .D(men_men_n1074_), .Y(men_men_n1221_));
  OAI220     u1193(.A0(men_men_n549_), .A1(men_men_n622_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n1222_), .B(men_men_n558_), .Y(men_men_n1223_));
  AOI220     u1195(.A0(men_men_n333_), .A1(men_men_n258_), .B0(men_men_n184_), .B1(men_men_n152_), .Y(men_men_n1224_));
  NA4        u1196(.A(men_men_n1224_), .B(men_men_n1223_), .C(men_men_n1221_), .D(men_men_n1219_), .Y(men_men_n1225_));
  NO3        u1197(.A(men_men_n1225_), .B(men_men_n1217_), .C(men_men_n279_), .Y(men_men_n1226_));
  INV        u1198(.A(men_men_n338_), .Y(men_men_n1227_));
  NA2        u1199(.A(men_men_n258_), .B(men_men_n365_), .Y(men_men_n1228_));
  NA3        u1200(.A(men_men_n1228_), .B(men_men_n1227_), .C(men_men_n158_), .Y(men_men_n1229_));
  NA3        u1201(.A(men_men_n186_), .B(men_men_n116_), .C(g), .Y(men_men_n1230_));
  NA3        u1202(.A(men_men_n488_), .B(men_men_n40_), .C(f), .Y(men_men_n1231_));
  NOi31      u1203(.An(men_men_n908_), .B(men_men_n1231_), .C(men_men_n1230_), .Y(men_men_n1232_));
  NAi31      u1204(.An(men_men_n193_), .B(men_men_n897_), .C(men_men_n488_), .Y(men_men_n1233_));
  NAi21      u1205(.An(men_men_n1232_), .B(men_men_n1233_), .Y(men_men_n1234_));
  INV        u1206(.A(men_men_n1123_), .Y(men_men_n1235_));
  NAi31      u1207(.An(men_men_n1088_), .B(men_men_n1235_), .C(men_men_n74_), .Y(men_men_n1236_));
  NO4        u1208(.A(men_men_n1236_), .B(men_men_n1234_), .C(men_men_n1229_), .D(men_men_n540_), .Y(men_men_n1237_));
  AN3        u1209(.A(men_men_n1237_), .B(men_men_n1226_), .C(men_men_n1216_), .Y(men_men_n1238_));
  NA2        u1210(.A(men_men_n558_), .B(men_men_n104_), .Y(men_men_n1239_));
  NA3        u1211(.A(men_men_n1156_), .B(men_men_n633_), .C(men_men_n487_), .Y(men_men_n1240_));
  NA4        u1212(.A(men_men_n1240_), .B(men_men_n586_), .C(men_men_n1239_), .D(men_men_n252_), .Y(men_men_n1241_));
  NA2        u1213(.A(men_men_n1149_), .B(men_men_n558_), .Y(men_men_n1242_));
  NA4        u1214(.A(men_men_n679_), .B(men_men_n214_), .C(men_men_n230_), .D(men_men_n167_), .Y(men_men_n1243_));
  NA3        u1215(.A(men_men_n1243_), .B(men_men_n1242_), .C(men_men_n309_), .Y(men_men_n1244_));
  OAI210     u1216(.A0(men_men_n486_), .A1(men_men_n124_), .B0(men_men_n902_), .Y(men_men_n1245_));
  AOI220     u1217(.A0(men_men_n1245_), .A1(men_men_n1188_), .B0(men_men_n585_), .B1(men_men_n432_), .Y(men_men_n1246_));
  OR4        u1218(.A(men_men_n1085_), .B(men_men_n285_), .C(men_men_n232_), .D(e), .Y(men_men_n1247_));
  NA2        u1219(.A(n), .B(e), .Y(men_men_n1248_));
  NO2        u1220(.A(men_men_n1248_), .B(men_men_n150_), .Y(men_men_n1249_));
  OAI210     u1221(.A0(men_men_n376_), .A1(men_men_n327_), .B0(men_men_n470_), .Y(men_men_n1250_));
  NA3        u1222(.A(men_men_n1250_), .B(men_men_n1247_), .C(men_men_n1246_), .Y(men_men_n1251_));
  AOI210     u1223(.A0(men_men_n1249_), .A1(men_men_n888_), .B0(men_men_n855_), .Y(men_men_n1252_));
  AOI220     u1224(.A0(men_men_n991_), .A1(men_men_n600_), .B0(men_men_n679_), .B1(men_men_n255_), .Y(men_men_n1253_));
  NO2        u1225(.A(men_men_n68_), .B(h), .Y(men_men_n1254_));
  NO3        u1226(.A(men_men_n1085_), .B(men_men_n1083_), .C(men_men_n760_), .Y(men_men_n1255_));
  INV        u1227(.A(men_men_n137_), .Y(men_men_n1256_));
  AN2        u1228(.A(men_men_n1256_), .B(men_men_n1135_), .Y(men_men_n1257_));
  OAI210     u1229(.A0(men_men_n1257_), .A1(men_men_n1255_), .B0(men_men_n1254_), .Y(men_men_n1258_));
  NA4        u1230(.A(men_men_n1258_), .B(men_men_n1253_), .C(men_men_n1252_), .D(men_men_n904_), .Y(men_men_n1259_));
  NO4        u1231(.A(men_men_n1259_), .B(men_men_n1251_), .C(men_men_n1244_), .D(men_men_n1241_), .Y(men_men_n1260_));
  NA2        u1232(.A(men_men_n872_), .B(men_men_n792_), .Y(men_men_n1261_));
  NA4        u1233(.A(men_men_n1261_), .B(men_men_n1260_), .C(men_men_n1238_), .D(men_men_n1209_), .Y(men01));
  AN2        u1234(.A(men_men_n1063_), .B(men_men_n1061_), .Y(men_men_n1263_));
  NO3        u1235(.A(men_men_n835_), .B(men_men_n827_), .C(men_men_n293_), .Y(men_men_n1264_));
  NA2        u1236(.A(men_men_n416_), .B(i), .Y(men_men_n1265_));
  NA3        u1237(.A(men_men_n1265_), .B(men_men_n1264_), .C(men_men_n1263_), .Y(men_men_n1266_));
  NA2        u1238(.A(men_men_n611_), .B(men_men_n92_), .Y(men_men_n1267_));
  NA2        u1239(.A(men_men_n578_), .B(men_men_n284_), .Y(men_men_n1268_));
  NA2        u1240(.A(men_men_n998_), .B(men_men_n1268_), .Y(men_men_n1269_));
  NA4        u1241(.A(men_men_n1269_), .B(men_men_n1267_), .C(men_men_n948_), .D(men_men_n350_), .Y(men_men_n1270_));
  NA2        u1242(.A(men_men_n45_), .B(f), .Y(men_men_n1271_));
  NA2        u1243(.A(men_men_n738_), .B(men_men_n99_), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n1272_), .B(men_men_n1271_), .Y(men_men_n1273_));
  OAI210     u1245(.A0(men_men_n815_), .A1(men_men_n628_), .B0(men_men_n1243_), .Y(men_men_n1274_));
  AOI210     u1246(.A0(men_men_n1273_), .A1(men_men_n664_), .B0(men_men_n1274_), .Y(men_men_n1275_));
  INV        u1247(.A(men_men_n122_), .Y(men_men_n1276_));
  OR2        u1248(.A(men_men_n692_), .B(men_men_n390_), .Y(men_men_n1277_));
  NAi41      u1249(.An(men_men_n166_), .B(men_men_n1277_), .C(men_men_n1275_), .D(men_men_n931_), .Y(men_men_n1278_));
  NO2        u1250(.A(men_men_n707_), .B(men_men_n535_), .Y(men_men_n1279_));
  NA4        u1251(.A(men_men_n738_), .B(men_men_n99_), .C(men_men_n45_), .D(men_men_n222_), .Y(men_men_n1280_));
  OA220      u1252(.A0(men_men_n1280_), .A1(men_men_n700_), .B0(men_men_n203_), .B1(men_men_n201_), .Y(men_men_n1281_));
  NA3        u1253(.A(men_men_n1281_), .B(men_men_n1279_), .C(men_men_n143_), .Y(men_men_n1282_));
  NO4        u1254(.A(men_men_n1282_), .B(men_men_n1278_), .C(men_men_n1270_), .D(men_men_n1266_), .Y(men_men_n1283_));
  NA2        u1255(.A(men_men_n315_), .B(men_men_n553_), .Y(men_men_n1284_));
  INV        u1256(.A(men_men_n561_), .Y(men_men_n1285_));
  NOi21      u1257(.An(men_men_n587_), .B(men_men_n606_), .Y(men_men_n1286_));
  NA2        u1258(.A(men_men_n1286_), .B(men_men_n1285_), .Y(men_men_n1287_));
  AOI210     u1259(.A0(men_men_n212_), .A1(men_men_n91_), .B0(men_men_n222_), .Y(men_men_n1288_));
  OAI210     u1260(.A0(men_men_n842_), .A1(men_men_n450_), .B0(men_men_n1288_), .Y(men_men_n1289_));
  AN3        u1261(.A(m), .B(l), .C(k), .Y(men_men_n1290_));
  OAI210     u1262(.A0(men_men_n378_), .A1(men_men_n34_), .B0(men_men_n1290_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n211_), .B(men_men_n34_), .Y(men_men_n1292_));
  AO210      u1264(.A0(men_men_n1292_), .A1(men_men_n1291_), .B0(men_men_n349_), .Y(men_men_n1293_));
  NA4        u1265(.A(men_men_n1293_), .B(men_men_n1289_), .C(men_men_n1287_), .D(men_men_n1284_), .Y(men_men_n1294_));
  AOI210     u1266(.A0(men_men_n620_), .A1(men_men_n122_), .B0(men_men_n626_), .Y(men_men_n1295_));
  OAI210     u1267(.A0(men_men_n1276_), .A1(men_men_n617_), .B0(men_men_n1295_), .Y(men_men_n1296_));
  NA2        u1268(.A(men_men_n292_), .B(men_men_n203_), .Y(men_men_n1297_));
  NA2        u1269(.A(men_men_n1297_), .B(men_men_n697_), .Y(men_men_n1298_));
  NO3        u1270(.A(men_men_n854_), .B(men_men_n212_), .C(men_men_n430_), .Y(men_men_n1299_));
  NO2        u1271(.A(men_men_n1299_), .B(men_men_n995_), .Y(men_men_n1300_));
  NA3        u1272(.A(men_men_n1300_), .B(men_men_n1298_), .C(men_men_n818_), .Y(men_men_n1301_));
  NO3        u1273(.A(men_men_n1301_), .B(men_men_n1296_), .C(men_men_n1294_), .Y(men_men_n1302_));
  NA3        u1274(.A(men_men_n629_), .B(men_men_n29_), .C(f), .Y(men_men_n1303_));
  NO2        u1275(.A(men_men_n1303_), .B(men_men_n212_), .Y(men_men_n1304_));
  AOI210     u1276(.A0(men_men_n527_), .A1(men_men_n58_), .B0(men_men_n1304_), .Y(men_men_n1305_));
  OR3        u1277(.A(men_men_n1272_), .B(men_men_n630_), .C(men_men_n1271_), .Y(men_men_n1306_));
  NO2        u1278(.A(men_men_n1280_), .B(men_men_n1016_), .Y(men_men_n1307_));
  NO2        u1279(.A(men_men_n215_), .B(men_men_n115_), .Y(men_men_n1308_));
  NO3        u1280(.A(men_men_n1308_), .B(men_men_n1307_), .C(men_men_n1214_), .Y(men_men_n1309_));
  NA4        u1281(.A(men_men_n1309_), .B(men_men_n1306_), .C(men_men_n1305_), .D(men_men_n791_), .Y(men_men_n1310_));
  NO2        u1282(.A(men_men_n1005_), .B(men_men_n242_), .Y(men_men_n1311_));
  NO2        u1283(.A(men_men_n1006_), .B(men_men_n580_), .Y(men_men_n1312_));
  OAI210     u1284(.A0(men_men_n1312_), .A1(men_men_n1311_), .B0(men_men_n358_), .Y(men_men_n1313_));
  NO3        u1285(.A(men_men_n81_), .B(men_men_n313_), .C(men_men_n45_), .Y(men_men_n1314_));
  NA2        u1286(.A(men_men_n1314_), .B(men_men_n577_), .Y(men_men_n1315_));
  NA2        u1287(.A(men_men_n1315_), .B(men_men_n702_), .Y(men_men_n1316_));
  OR2        u1288(.A(men_men_n1218_), .B(men_men_n1211_), .Y(men_men_n1317_));
  NO2        u1289(.A(men_men_n390_), .B(men_men_n73_), .Y(men_men_n1318_));
  INV        u1290(.A(men_men_n1318_), .Y(men_men_n1319_));
  NA2        u1291(.A(men_men_n1314_), .B(men_men_n845_), .Y(men_men_n1320_));
  NA4        u1292(.A(men_men_n1320_), .B(men_men_n1319_), .C(men_men_n1317_), .D(men_men_n408_), .Y(men_men_n1321_));
  NOi41      u1293(.An(men_men_n1313_), .B(men_men_n1321_), .C(men_men_n1316_), .D(men_men_n1310_), .Y(men_men_n1322_));
  NO2        u1294(.A(men_men_n136_), .B(men_men_n45_), .Y(men_men_n1323_));
  NO2        u1295(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1324_));
  AO220      u1296(.A0(men_men_n1324_), .A1(men_men_n650_), .B0(men_men_n1323_), .B1(men_men_n736_), .Y(men_men_n1325_));
  NA2        u1297(.A(men_men_n1325_), .B(men_men_n358_), .Y(men_men_n1326_));
  INV        u1298(.A(men_men_n140_), .Y(men_men_n1327_));
  NO3        u1299(.A(men_men_n1133_), .B(men_men_n183_), .C(men_men_n89_), .Y(men_men_n1328_));
  NA2        u1300(.A(men_men_n1328_), .B(men_men_n1327_), .Y(men_men_n1329_));
  NA2        u1301(.A(men_men_n1329_), .B(men_men_n1326_), .Y(men_men_n1330_));
  NO2        u1302(.A(men_men_n641_), .B(men_men_n640_), .Y(men_men_n1331_));
  NO4        u1303(.A(men_men_n1133_), .B(men_men_n1331_), .C(men_men_n181_), .D(men_men_n89_), .Y(men_men_n1332_));
  NO3        u1304(.A(men_men_n1332_), .B(men_men_n1330_), .C(men_men_n668_), .Y(men_men_n1333_));
  NA4        u1305(.A(men_men_n1333_), .B(men_men_n1322_), .C(men_men_n1302_), .D(men_men_n1283_), .Y(men06));
  NO2        u1306(.A(men_men_n431_), .B(men_men_n584_), .Y(men_men_n1335_));
  INV        u1307(.A(men_men_n767_), .Y(men_men_n1336_));
  OAI210     u1308(.A0(men_men_n1336_), .A1(men_men_n280_), .B0(men_men_n1335_), .Y(men_men_n1337_));
  NO2        u1309(.A(men_men_n234_), .B(men_men_n106_), .Y(men_men_n1338_));
  OAI210     u1310(.A0(men_men_n1338_), .A1(men_men_n1328_), .B0(men_men_n404_), .Y(men_men_n1339_));
  NO3        u1311(.A(men_men_n624_), .B(men_men_n840_), .C(men_men_n627_), .Y(men_men_n1340_));
  OR2        u1312(.A(men_men_n1340_), .B(men_men_n922_), .Y(men_men_n1341_));
  NA4        u1313(.A(men_men_n1341_), .B(men_men_n1339_), .C(men_men_n1337_), .D(men_men_n1313_), .Y(men_men_n1342_));
  NO3        u1314(.A(men_men_n1342_), .B(men_men_n1316_), .C(men_men_n268_), .Y(men_men_n1343_));
  NO2        u1315(.A(men_men_n313_), .B(men_men_n45_), .Y(men_men_n1344_));
  AOI210     u1316(.A0(men_men_n1344_), .A1(men_men_n577_), .B0(men_men_n1311_), .Y(men_men_n1345_));
  AOI210     u1317(.A0(men_men_n1344_), .A1(men_men_n581_), .B0(men_men_n1325_), .Y(men_men_n1346_));
  AOI210     u1318(.A0(men_men_n1346_), .A1(men_men_n1345_), .B0(men_men_n355_), .Y(men_men_n1347_));
  OAI210     u1319(.A0(men_men_n91_), .A1(men_men_n40_), .B0(men_men_n706_), .Y(men_men_n1348_));
  NA2        u1320(.A(men_men_n1348_), .B(men_men_n672_), .Y(men_men_n1349_));
  NO2        u1321(.A(men_men_n537_), .B(men_men_n178_), .Y(men_men_n1350_));
  NOi21      u1322(.An(men_men_n142_), .B(men_men_n45_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n634_), .B(men_men_n1157_), .Y(men_men_n1352_));
  OAI210     u1324(.A0(men_men_n481_), .A1(men_men_n259_), .B0(men_men_n942_), .Y(men_men_n1353_));
  NO4        u1325(.A(men_men_n1353_), .B(men_men_n1352_), .C(men_men_n1351_), .D(men_men_n1350_), .Y(men_men_n1354_));
  OR2        u1326(.A(men_men_n625_), .B(men_men_n623_), .Y(men_men_n1355_));
  NO2        u1327(.A(men_men_n389_), .B(men_men_n141_), .Y(men_men_n1356_));
  AOI210     u1328(.A0(men_men_n1356_), .A1(men_men_n611_), .B0(men_men_n1355_), .Y(men_men_n1357_));
  NA3        u1329(.A(men_men_n1357_), .B(men_men_n1354_), .C(men_men_n1349_), .Y(men_men_n1358_));
  NO2        u1330(.A(men_men_n782_), .B(men_men_n388_), .Y(men_men_n1359_));
  NO2        u1331(.A(men_men_n793_), .B(men_men_n664_), .Y(men_men_n1360_));
  NOi21      u1332(.An(men_men_n1359_), .B(men_men_n1360_), .Y(men_men_n1361_));
  AN2        u1333(.A(men_men_n991_), .B(men_men_n675_), .Y(men_men_n1362_));
  NO4        u1334(.A(men_men_n1362_), .B(men_men_n1361_), .C(men_men_n1358_), .D(men_men_n1347_), .Y(men_men_n1363_));
  NO2        u1335(.A(men_men_n834_), .B(men_men_n289_), .Y(men_men_n1364_));
  OAI220     u1336(.A0(men_men_n767_), .A1(men_men_n47_), .B0(men_men_n234_), .B1(men_men_n643_), .Y(men_men_n1365_));
  OAI210     u1337(.A0(men_men_n289_), .A1(c), .B0(men_men_n671_), .Y(men_men_n1366_));
  AOI220     u1338(.A0(men_men_n1366_), .A1(men_men_n1365_), .B0(men_men_n1364_), .B1(men_men_n280_), .Y(men_men_n1367_));
  NO3        u1339(.A(men_men_n254_), .B(men_men_n106_), .C(men_men_n295_), .Y(men_men_n1368_));
  OAI220     u1340(.A0(men_men_n728_), .A1(men_men_n259_), .B0(men_men_n534_), .B1(men_men_n537_), .Y(men_men_n1369_));
  OAI210     u1341(.A0(l), .A1(i), .B0(k), .Y(men_men_n1370_));
  NO3        u1342(.A(men_men_n1370_), .B(men_men_n622_), .C(j), .Y(men_men_n1371_));
  NOi21      u1343(.An(men_men_n1371_), .B(men_men_n700_), .Y(men_men_n1372_));
  NO4        u1344(.A(men_men_n1372_), .B(men_men_n1369_), .C(men_men_n1368_), .D(men_men_n1159_), .Y(men_men_n1373_));
  NA4        u1345(.A(men_men_n825_), .B(men_men_n824_), .C(men_men_n460_), .D(men_men_n914_), .Y(men_men_n1374_));
  NAi31      u1346(.An(men_men_n782_), .B(men_men_n1374_), .C(men_men_n211_), .Y(men_men_n1375_));
  NA4        u1347(.A(men_men_n1375_), .B(men_men_n1373_), .C(men_men_n1367_), .D(men_men_n1253_), .Y(men_men_n1376_));
  NOi31      u1348(.An(men_men_n1340_), .B(men_men_n485_), .C(men_men_n417_), .Y(men_men_n1377_));
  OR3        u1349(.A(men_men_n1377_), .B(men_men_n815_), .C(men_men_n564_), .Y(men_men_n1378_));
  OR3        u1350(.A(men_men_n392_), .B(men_men_n234_), .C(men_men_n643_), .Y(men_men_n1379_));
  AOI210     u1351(.A0(men_men_n595_), .A1(men_men_n470_), .B0(men_men_n394_), .Y(men_men_n1380_));
  NA2        u1352(.A(men_men_n1371_), .B(men_men_n821_), .Y(men_men_n1381_));
  NA4        u1353(.A(men_men_n1381_), .B(men_men_n1380_), .C(men_men_n1379_), .D(men_men_n1378_), .Y(men_men_n1382_));
  AOI220     u1354(.A0(men_men_n1359_), .A1(men_men_n792_), .B0(men_men_n1356_), .B1(men_men_n248_), .Y(men_men_n1383_));
  AN2        u1355(.A(men_men_n964_), .B(men_men_n963_), .Y(men_men_n1384_));
  NO4        u1356(.A(men_men_n1384_), .B(men_men_n912_), .C(men_men_n523_), .D(men_men_n502_), .Y(men_men_n1385_));
  NA3        u1357(.A(men_men_n1385_), .B(men_men_n1383_), .C(men_men_n1320_), .Y(men_men_n1386_));
  NAi21      u1358(.An(j), .B(i), .Y(men_men_n1387_));
  NO4        u1359(.A(men_men_n1331_), .B(men_men_n1387_), .C(men_men_n464_), .D(men_men_n245_), .Y(men_men_n1388_));
  NO4        u1360(.A(men_men_n1388_), .B(men_men_n1386_), .C(men_men_n1382_), .D(men_men_n1376_), .Y(men_men_n1389_));
  NA4        u1361(.A(men_men_n1389_), .B(men_men_n1363_), .C(men_men_n1343_), .D(men_men_n1333_), .Y(men07));
  NOi21      u1362(.An(j), .B(k), .Y(men_men_n1391_));
  NA4        u1363(.A(men_men_n186_), .B(men_men_n112_), .C(men_men_n1391_), .D(f), .Y(men_men_n1392_));
  NAi32      u1364(.An(m), .Bn(b), .C(n), .Y(men_men_n1393_));
  NO3        u1365(.A(men_men_n1393_), .B(g), .C(f), .Y(men_men_n1394_));
  OAI210     u1366(.A0(men_men_n337_), .A1(men_men_n504_), .B0(men_men_n1394_), .Y(men_men_n1395_));
  NAi21      u1367(.An(f), .B(c), .Y(men_men_n1396_));
  OR2        u1368(.A(e), .B(d), .Y(men_men_n1397_));
  OAI220     u1369(.A0(men_men_n1397_), .A1(men_men_n1396_), .B0(men_men_n656_), .B1(men_men_n339_), .Y(men_men_n1398_));
  NA3        u1370(.A(men_men_n1398_), .B(men_men_n1097_), .C(men_men_n186_), .Y(men_men_n1399_));
  NOi31      u1371(.An(n), .B(m), .C(b), .Y(men_men_n1400_));
  NO3        u1372(.A(men_men_n137_), .B(men_men_n471_), .C(h), .Y(men_men_n1401_));
  NA3        u1373(.A(men_men_n1399_), .B(men_men_n1395_), .C(men_men_n1392_), .Y(men_men_n1402_));
  NOi41      u1374(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1403_));
  NA3        u1375(.A(men_men_n1403_), .B(men_men_n905_), .C(men_men_n433_), .Y(men_men_n1404_));
  NO2        u1376(.A(men_men_n1404_), .B(men_men_n56_), .Y(men_men_n1405_));
  NA2        u1377(.A(men_men_n1135_), .B(men_men_n230_), .Y(men_men_n1406_));
  NO2        u1378(.A(men_men_n1406_), .B(men_men_n61_), .Y(men_men_n1407_));
  NO2        u1379(.A(k), .B(i), .Y(men_men_n1408_));
  NA3        u1380(.A(men_men_n1408_), .B(men_men_n930_), .C(men_men_n186_), .Y(men_men_n1409_));
  NA2        u1381(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1410_));
  NO2        u1382(.A(men_men_n1091_), .B(men_men_n464_), .Y(men_men_n1411_));
  NA3        u1383(.A(men_men_n1411_), .B(men_men_n1410_), .C(men_men_n223_), .Y(men_men_n1412_));
  NO2        u1384(.A(men_men_n1105_), .B(men_men_n321_), .Y(men_men_n1413_));
  NA2        u1385(.A(men_men_n565_), .B(men_men_n82_), .Y(men_men_n1414_));
  NA2        u1386(.A(men_men_n1254_), .B(men_men_n303_), .Y(men_men_n1415_));
  NA4        u1387(.A(men_men_n1415_), .B(men_men_n1414_), .C(men_men_n1412_), .D(men_men_n1409_), .Y(men_men_n1416_));
  NO4        u1388(.A(men_men_n1416_), .B(men_men_n1407_), .C(men_men_n1405_), .D(men_men_n1402_), .Y(men_men_n1417_));
  NO3        u1389(.A(e), .B(d), .C(c), .Y(men_men_n1418_));
  OAI210     u1390(.A0(men_men_n137_), .A1(men_men_n223_), .B0(men_men_n631_), .Y(men_men_n1419_));
  NA2        u1391(.A(men_men_n1419_), .B(men_men_n1418_), .Y(men_men_n1420_));
  INV        u1392(.A(men_men_n1420_), .Y(men_men_n1421_));
  OR2        u1393(.A(h), .B(f), .Y(men_men_n1422_));
  NO3        u1394(.A(n), .B(m), .C(i), .Y(men_men_n1423_));
  OAI210     u1395(.A0(men_men_n1158_), .A1(men_men_n161_), .B0(men_men_n1423_), .Y(men_men_n1424_));
  NO2        u1396(.A(i), .B(g), .Y(men_men_n1425_));
  OR3        u1397(.A(men_men_n1425_), .B(men_men_n1393_), .C(men_men_n72_), .Y(men_men_n1426_));
  OAI220     u1398(.A0(men_men_n1426_), .A1(men_men_n504_), .B0(men_men_n1424_), .B1(men_men_n1422_), .Y(men_men_n1427_));
  NA3        u1399(.A(men_men_n725_), .B(men_men_n714_), .C(men_men_n116_), .Y(men_men_n1428_));
  NA3        u1400(.A(men_men_n1400_), .B(men_men_n1100_), .C(men_men_n704_), .Y(men_men_n1429_));
  AOI210     u1401(.A0(men_men_n1429_), .A1(men_men_n1428_), .B0(men_men_n45_), .Y(men_men_n1430_));
  NO2        u1402(.A(l), .B(k), .Y(men_men_n1431_));
  NOi41      u1403(.An(men_men_n570_), .B(men_men_n1431_), .C(men_men_n499_), .D(men_men_n464_), .Y(men_men_n1432_));
  NO3        u1404(.A(men_men_n464_), .B(d), .C(c), .Y(men_men_n1433_));
  NO4        u1405(.A(men_men_n1432_), .B(men_men_n1430_), .C(men_men_n1427_), .D(men_men_n1421_), .Y(men_men_n1434_));
  NO2        u1406(.A(men_men_n151_), .B(h), .Y(men_men_n1435_));
  NO2        u1407(.A(men_men_n1115_), .B(l), .Y(men_men_n1436_));
  NO2        u1408(.A(g), .B(c), .Y(men_men_n1437_));
  NA3        u1409(.A(men_men_n1437_), .B(men_men_n147_), .C(men_men_n194_), .Y(men_men_n1438_));
  NO2        u1410(.A(men_men_n1438_), .B(men_men_n1436_), .Y(men_men_n1439_));
  NA2        u1411(.A(men_men_n1439_), .B(men_men_n186_), .Y(men_men_n1440_));
  NO2        u1412(.A(men_men_n472_), .B(a), .Y(men_men_n1441_));
  NA3        u1413(.A(men_men_n1441_), .B(k), .C(men_men_n117_), .Y(men_men_n1442_));
  NO2        u1414(.A(i), .B(h), .Y(men_men_n1443_));
  NA2        u1415(.A(men_men_n1443_), .B(men_men_n230_), .Y(men_men_n1444_));
  AOI210     u1416(.A0(men_men_n1180_), .A1(h), .B0(men_men_n438_), .Y(men_men_n1445_));
  NA2        u1417(.A(men_men_n144_), .B(men_men_n230_), .Y(men_men_n1446_));
  AOI210     u1418(.A0(men_men_n269_), .A1(men_men_n120_), .B0(men_men_n553_), .Y(men_men_n1447_));
  OAI220     u1419(.A0(men_men_n1447_), .A1(men_men_n1444_), .B0(men_men_n1446_), .B1(men_men_n1445_), .Y(men_men_n1448_));
  NO2        u1420(.A(men_men_n789_), .B(men_men_n195_), .Y(men_men_n1449_));
  NOi31      u1421(.An(m), .B(n), .C(b), .Y(men_men_n1450_));
  NOi31      u1422(.An(f), .B(d), .C(c), .Y(men_men_n1451_));
  NA2        u1423(.A(men_men_n1451_), .B(men_men_n1450_), .Y(men_men_n1452_));
  INV        u1424(.A(men_men_n1452_), .Y(men_men_n1453_));
  NO3        u1425(.A(men_men_n1453_), .B(men_men_n1449_), .C(men_men_n1448_), .Y(men_men_n1454_));
  NA2        u1426(.A(men_men_n1126_), .B(men_men_n488_), .Y(men_men_n1455_));
  NO4        u1427(.A(men_men_n1455_), .B(men_men_n1100_), .C(men_men_n464_), .D(men_men_n45_), .Y(men_men_n1456_));
  OAI210     u1428(.A0(men_men_n189_), .A1(men_men_n548_), .B0(men_men_n1101_), .Y(men_men_n1457_));
  NO3        u1429(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1458_));
  INV        u1430(.A(men_men_n1457_), .Y(men_men_n1459_));
  NO2        u1431(.A(men_men_n1459_), .B(men_men_n1456_), .Y(men_men_n1460_));
  AN4        u1432(.A(men_men_n1460_), .B(men_men_n1454_), .C(men_men_n1442_), .D(men_men_n1440_), .Y(men_men_n1461_));
  NA2        u1433(.A(men_men_n1400_), .B(men_men_n401_), .Y(men_men_n1462_));
  NA2        u1434(.A(men_men_n1433_), .B(men_men_n224_), .Y(men_men_n1463_));
  NO2        u1435(.A(men_men_n195_), .B(b), .Y(men_men_n1464_));
  AOI220     u1436(.A0(men_men_n1212_), .A1(men_men_n1464_), .B0(men_men_n1134_), .B1(men_men_n1455_), .Y(men_men_n1465_));
  NO2        u1437(.A(i), .B(men_men_n222_), .Y(men_men_n1466_));
  NA4        u1438(.A(men_men_n1186_), .B(men_men_n1466_), .C(men_men_n107_), .D(m), .Y(men_men_n1467_));
  NA3        u1439(.A(men_men_n1467_), .B(men_men_n1465_), .C(men_men_n1463_), .Y(men_men_n1468_));
  NO4        u1440(.A(men_men_n137_), .B(g), .C(f), .D(e), .Y(men_men_n1469_));
  NA3        u1441(.A(men_men_n1408_), .B(men_men_n304_), .C(h), .Y(men_men_n1470_));
  NA2        u1442(.A(men_men_n202_), .B(men_men_n101_), .Y(men_men_n1471_));
  OR2        u1443(.A(e), .B(a), .Y(men_men_n1472_));
  NO2        u1444(.A(men_men_n1397_), .B(men_men_n1396_), .Y(men_men_n1473_));
  AOI210     u1445(.A0(men_men_n30_), .A1(h), .B0(men_men_n1473_), .Y(men_men_n1474_));
  NO2        u1446(.A(men_men_n1474_), .B(men_men_n1122_), .Y(men_men_n1475_));
  NA2        u1447(.A(men_men_n1403_), .B(men_men_n1431_), .Y(men_men_n1476_));
  INV        u1448(.A(men_men_n1476_), .Y(men_men_n1477_));
  OR3        u1449(.A(men_men_n564_), .B(men_men_n563_), .C(men_men_n116_), .Y(men_men_n1478_));
  NA2        u1450(.A(men_men_n1156_), .B(men_men_n430_), .Y(men_men_n1479_));
  OAI220     u1451(.A0(men_men_n1479_), .A1(men_men_n459_), .B0(men_men_n1478_), .B1(men_men_n313_), .Y(men_men_n1480_));
  AO210      u1452(.A0(men_men_n1480_), .A1(men_men_n120_), .B0(men_men_n1477_), .Y(men_men_n1481_));
  NO3        u1453(.A(men_men_n1481_), .B(men_men_n1475_), .C(men_men_n1468_), .Y(men_men_n1482_));
  NA4        u1454(.A(men_men_n1482_), .B(men_men_n1461_), .C(men_men_n1434_), .D(men_men_n1417_), .Y(men_men_n1483_));
  NO2        u1455(.A(men_men_n1171_), .B(men_men_n114_), .Y(men_men_n1484_));
  NA2        u1456(.A(men_men_n401_), .B(men_men_n56_), .Y(men_men_n1485_));
  NA2        u1457(.A(men_men_n224_), .B(men_men_n186_), .Y(men_men_n1486_));
  AOI210     u1458(.A0(men_men_n1486_), .A1(men_men_n1230_), .B0(men_men_n1485_), .Y(men_men_n1487_));
  NO2        u1459(.A(men_men_n413_), .B(j), .Y(men_men_n1488_));
  NA3        u1460(.A(men_men_n1458_), .B(men_men_n1397_), .C(men_men_n1156_), .Y(men_men_n1489_));
  NAi41      u1461(.An(men_men_n1443_), .B(men_men_n1113_), .C(men_men_n174_), .D(men_men_n154_), .Y(men_men_n1490_));
  NA2        u1462(.A(men_men_n1490_), .B(men_men_n1489_), .Y(men_men_n1491_));
  NA3        u1463(.A(g), .B(men_men_n1488_), .C(men_men_n163_), .Y(men_men_n1492_));
  INV        u1464(.A(men_men_n1492_), .Y(men_men_n1493_));
  NO3        u1465(.A(men_men_n782_), .B(men_men_n181_), .C(men_men_n433_), .Y(men_men_n1494_));
  NO3        u1466(.A(men_men_n1494_), .B(men_men_n1493_), .C(men_men_n1491_), .Y(men_men_n1495_));
  NO3        u1467(.A(men_men_n1122_), .B(men_men_n606_), .C(g), .Y(men_men_n1496_));
  NOi21      u1468(.An(men_men_n1486_), .B(men_men_n1496_), .Y(men_men_n1497_));
  AOI210     u1469(.A0(men_men_n1497_), .A1(men_men_n1471_), .B0(men_men_n1091_), .Y(men_men_n1498_));
  OR2        u1470(.A(n), .B(i), .Y(men_men_n1499_));
  OAI210     u1471(.A0(men_men_n1499_), .A1(men_men_n1112_), .B0(men_men_n49_), .Y(men_men_n1500_));
  AOI220     u1472(.A0(men_men_n1500_), .A1(men_men_n1220_), .B0(men_men_n859_), .B1(men_men_n202_), .Y(men_men_n1501_));
  INV        u1473(.A(men_men_n1501_), .Y(men_men_n1502_));
  NO2        u1474(.A(men_men_n234_), .B(k), .Y(men_men_n1503_));
  NO2        u1475(.A(men_men_n1502_), .B(men_men_n1498_), .Y(men_men_n1504_));
  INV        u1476(.A(men_men_n49_), .Y(men_men_n1505_));
  NO3        u1477(.A(men_men_n1137_), .B(men_men_n1397_), .C(men_men_n49_), .Y(men_men_n1506_));
  NA2        u1478(.A(men_men_n1138_), .B(men_men_n1505_), .Y(men_men_n1507_));
  NO2        u1479(.A(men_men_n1122_), .B(h), .Y(men_men_n1508_));
  NA3        u1480(.A(men_men_n1508_), .B(d), .C(men_men_n1083_), .Y(men_men_n1509_));
  OAI220     u1481(.A0(men_men_n1509_), .A1(c), .B0(men_men_n1507_), .B1(j), .Y(men_men_n1510_));
  NA3        u1482(.A(men_men_n1484_), .B(men_men_n488_), .C(f), .Y(men_men_n1511_));
  NA2        u1483(.A(men_men_n186_), .B(men_men_n116_), .Y(men_men_n1512_));
  NO2        u1484(.A(men_men_n1391_), .B(men_men_n42_), .Y(men_men_n1513_));
  NA2        u1485(.A(men_men_n117_), .B(men_men_n40_), .Y(men_men_n1514_));
  NO2        u1486(.A(men_men_n1514_), .B(men_men_n1511_), .Y(men_men_n1515_));
  AOI210     u1487(.A0(men_men_n548_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1516_));
  NA2        u1488(.A(men_men_n1516_), .B(men_men_n1441_), .Y(men_men_n1517_));
  NO2        u1489(.A(men_men_n1387_), .B(men_men_n181_), .Y(men_men_n1518_));
  NOi21      u1490(.An(d), .B(f), .Y(men_men_n1519_));
  NO3        u1491(.A(men_men_n1451_), .B(men_men_n1519_), .C(men_men_n40_), .Y(men_men_n1520_));
  NA2        u1492(.A(men_men_n1520_), .B(men_men_n1518_), .Y(men_men_n1521_));
  NO2        u1493(.A(men_men_n1397_), .B(f), .Y(men_men_n1522_));
  NA2        u1494(.A(men_men_n1441_), .B(men_men_n1513_), .Y(men_men_n1523_));
  NO2        u1495(.A(men_men_n313_), .B(c), .Y(men_men_n1524_));
  NA2        u1496(.A(men_men_n1524_), .B(men_men_n565_), .Y(men_men_n1525_));
  NA4        u1497(.A(men_men_n1525_), .B(men_men_n1523_), .C(men_men_n1521_), .D(men_men_n1517_), .Y(men_men_n1526_));
  NO3        u1498(.A(men_men_n1526_), .B(men_men_n1515_), .C(men_men_n1510_), .Y(men_men_n1527_));
  NA4        u1499(.A(men_men_n1527_), .B(men_men_n1504_), .C(men_men_n1495_), .D(men_men_n1610_), .Y(men_men_n1528_));
  NO3        u1500(.A(men_men_n1126_), .B(men_men_n1112_), .C(men_men_n40_), .Y(men_men_n1529_));
  NO2        u1501(.A(men_men_n488_), .B(men_men_n313_), .Y(men_men_n1530_));
  OAI210     u1502(.A0(men_men_n1530_), .A1(men_men_n1529_), .B0(men_men_n1413_), .Y(men_men_n1531_));
  OAI210     u1503(.A0(men_men_n1469_), .A1(men_men_n1400_), .B0(men_men_n919_), .Y(men_men_n1532_));
  NO2        u1504(.A(men_men_n1080_), .B(men_men_n137_), .Y(men_men_n1533_));
  NA2        u1505(.A(men_men_n1533_), .B(men_men_n649_), .Y(men_men_n1534_));
  NA3        u1506(.A(men_men_n1534_), .B(men_men_n1532_), .C(men_men_n1531_), .Y(men_men_n1535_));
  NA2        u1507(.A(men_men_n1437_), .B(men_men_n1519_), .Y(men_men_n1536_));
  NO2        u1508(.A(men_men_n1536_), .B(m), .Y(men_men_n1537_));
  NA3        u1509(.A(men_men_n1135_), .B(men_men_n112_), .C(men_men_n230_), .Y(men_men_n1538_));
  NO2        u1510(.A(men_men_n155_), .B(men_men_n188_), .Y(men_men_n1539_));
  OAI210     u1511(.A0(men_men_n1539_), .A1(men_men_n114_), .B0(men_men_n1450_), .Y(men_men_n1540_));
  NA2        u1512(.A(men_men_n1540_), .B(men_men_n1538_), .Y(men_men_n1541_));
  NO3        u1513(.A(men_men_n1541_), .B(men_men_n1537_), .C(men_men_n1535_), .Y(men_men_n1542_));
  NO2        u1514(.A(men_men_n1396_), .B(e), .Y(men_men_n1543_));
  NA2        u1515(.A(men_men_n1543_), .B(men_men_n428_), .Y(men_men_n1544_));
  OAI210     u1516(.A0(men_men_n1522_), .A1(men_men_n1166_), .B0(men_men_n660_), .Y(men_men_n1545_));
  OR3        u1517(.A(men_men_n1503_), .B(men_men_n1254_), .C(men_men_n137_), .Y(men_men_n1546_));
  OAI220     u1518(.A0(men_men_n1546_), .A1(men_men_n1544_), .B0(men_men_n1545_), .B1(men_men_n466_), .Y(men_men_n1547_));
  NO3        u1519(.A(men_men_n1478_), .B(men_men_n372_), .C(a), .Y(men_men_n1548_));
  NO2        u1520(.A(men_men_n1548_), .B(men_men_n1547_), .Y(men_men_n1549_));
  NO2        u1521(.A(men_men_n188_), .B(c), .Y(men_men_n1550_));
  OAI210     u1522(.A0(men_men_n1550_), .A1(men_men_n1543_), .B0(men_men_n186_), .Y(men_men_n1551_));
  AOI220     u1523(.A0(men_men_n1551_), .A1(men_men_n1114_), .B0(men_men_n555_), .B1(men_men_n388_), .Y(men_men_n1552_));
  NA2        u1524(.A(men_men_n563_), .B(g), .Y(men_men_n1553_));
  AOI210     u1525(.A0(men_men_n1553_), .A1(men_men_n1433_), .B0(men_men_n1506_), .Y(men_men_n1554_));
  NO2        u1526(.A(men_men_n1472_), .B(f), .Y(men_men_n1555_));
  NA2        u1527(.A(men_men_n1166_), .B(a), .Y(men_men_n1556_));
  OAI220     u1528(.A0(men_men_n1556_), .A1(men_men_n69_), .B0(men_men_n1554_), .B1(men_men_n222_), .Y(men_men_n1557_));
  AOI210     u1529(.A0(men_men_n935_), .A1(men_men_n440_), .B0(men_men_n108_), .Y(men_men_n1558_));
  OR2        u1530(.A(men_men_n1558_), .B(men_men_n563_), .Y(men_men_n1559_));
  NA2        u1531(.A(men_men_n1555_), .B(men_men_n1410_), .Y(men_men_n1560_));
  OAI220     u1532(.A0(men_men_n1560_), .A1(men_men_n49_), .B0(men_men_n1559_), .B1(men_men_n181_), .Y(men_men_n1561_));
  NA4        u1533(.A(men_men_n1135_), .B(men_men_n1132_), .C(men_men_n230_), .D(men_men_n68_), .Y(men_men_n1562_));
  NA2        u1534(.A(men_men_n1401_), .B(men_men_n189_), .Y(men_men_n1563_));
  NO2        u1535(.A(men_men_n49_), .B(l), .Y(men_men_n1564_));
  OAI210     u1536(.A0(men_men_n1472_), .A1(men_men_n898_), .B0(men_men_n504_), .Y(men_men_n1565_));
  OAI210     u1537(.A0(men_men_n1565_), .A1(men_men_n1138_), .B0(men_men_n1564_), .Y(men_men_n1566_));
  NO2        u1538(.A(men_men_n264_), .B(g), .Y(men_men_n1567_));
  NO2        u1539(.A(m), .B(i), .Y(men_men_n1568_));
  BUFFER     u1540(.A(men_men_n1568_), .Y(men_men_n1569_));
  AOI220     u1541(.A0(men_men_n1569_), .A1(men_men_n1435_), .B0(men_men_n1113_), .B1(men_men_n1567_), .Y(men_men_n1570_));
  NA4        u1542(.A(men_men_n1570_), .B(men_men_n1566_), .C(men_men_n1563_), .D(men_men_n1562_), .Y(men_men_n1571_));
  NO4        u1543(.A(men_men_n1571_), .B(men_men_n1561_), .C(men_men_n1557_), .D(men_men_n1552_), .Y(men_men_n1572_));
  NA3        u1544(.A(men_men_n1572_), .B(men_men_n1549_), .C(men_men_n1542_), .Y(men_men_n1573_));
  NA3        u1545(.A(men_men_n997_), .B(men_men_n144_), .C(men_men_n46_), .Y(men_men_n1574_));
  AOI210     u1546(.A0(men_men_n152_), .A1(c), .B0(men_men_n1574_), .Y(men_men_n1575_));
  INV        u1547(.A(men_men_n192_), .Y(men_men_n1576_));
  NA2        u1548(.A(men_men_n1576_), .B(men_men_n1508_), .Y(men_men_n1577_));
  AO210      u1549(.A0(men_men_n138_), .A1(l), .B0(men_men_n1462_), .Y(men_men_n1578_));
  NO2        u1550(.A(men_men_n72_), .B(c), .Y(men_men_n1579_));
  NO4        u1551(.A(men_men_n1422_), .B(men_men_n193_), .C(men_men_n471_), .D(men_men_n45_), .Y(men_men_n1580_));
  AOI210     u1552(.A0(men_men_n1518_), .A1(men_men_n1579_), .B0(men_men_n1580_), .Y(men_men_n1581_));
  NA3        u1553(.A(men_men_n1581_), .B(men_men_n1578_), .C(men_men_n1577_), .Y(men_men_n1582_));
  NO2        u1554(.A(men_men_n1582_), .B(men_men_n1575_), .Y(men_men_n1583_));
  NO4        u1555(.A(men_men_n234_), .B(men_men_n193_), .C(men_men_n269_), .D(k), .Y(men_men_n1584_));
  AOI210     u1556(.A0(men_men_n161_), .A1(men_men_n56_), .B0(men_men_n1543_), .Y(men_men_n1585_));
  NO2        u1557(.A(men_men_n1585_), .B(men_men_n1512_), .Y(men_men_n1586_));
  NO2        u1558(.A(men_men_n1574_), .B(men_men_n114_), .Y(men_men_n1587_));
  NOi21      u1559(.An(men_men_n1401_), .B(e), .Y(men_men_n1588_));
  NO4        u1560(.A(men_men_n1588_), .B(men_men_n1587_), .C(men_men_n1586_), .D(men_men_n1584_), .Y(men_men_n1589_));
  AOI220     u1561(.A0(men_men_n1568_), .A1(men_men_n670_), .B0(men_men_n1097_), .B1(men_men_n164_), .Y(men_men_n1590_));
  NOi31      u1562(.An(men_men_n30_), .B(men_men_n1590_), .C(n), .Y(men_men_n1591_));
  INV        u1563(.A(men_men_n1591_), .Y(men_men_n1592_));
  NA2        u1564(.A(men_men_n59_), .B(a), .Y(men_men_n1593_));
  NO2        u1565(.A(men_men_n1408_), .B(men_men_n122_), .Y(men_men_n1594_));
  OAI220     u1566(.A0(men_men_n1594_), .A1(men_men_n1462_), .B0(men_men_n1479_), .B1(men_men_n1593_), .Y(men_men_n1595_));
  NA4        u1567(.A(men_men_n1609_), .B(men_men_n1592_), .C(men_men_n1589_), .D(men_men_n1583_), .Y(men_men_n1596_));
  OR4        u1568(.A(men_men_n1596_), .B(men_men_n1573_), .C(men_men_n1528_), .D(men_men_n1483_), .Y(men04));
  NOi31      u1569(.An(men_men_n1469_), .B(men_men_n1470_), .C(men_men_n1085_), .Y(men_men_n1598_));
  NA2        u1570(.A(men_men_n1522_), .B(men_men_n859_), .Y(men_men_n1599_));
  NO4        u1571(.A(men_men_n1599_), .B(men_men_n1075_), .C(men_men_n505_), .D(j), .Y(men_men_n1600_));
  OR3        u1572(.A(men_men_n1600_), .B(men_men_n1598_), .C(men_men_n1103_), .Y(men_men_n1601_));
  NO3        u1573(.A(men_men_n1410_), .B(men_men_n93_), .C(k), .Y(men_men_n1602_));
  AOI210     u1574(.A0(men_men_n1602_), .A1(men_men_n1096_), .B0(men_men_n1232_), .Y(men_men_n1603_));
  NA2        u1575(.A(men_men_n1603_), .B(men_men_n1258_), .Y(men_men_n1604_));
  NO4        u1576(.A(men_men_n1604_), .B(men_men_n1601_), .C(men_men_n1111_), .D(men_men_n1090_), .Y(men_men_n1605_));
  NA4        u1577(.A(men_men_n1605_), .B(men_men_n1168_), .C(men_men_n1154_), .D(men_men_n1141_), .Y(men05));
  INV        u1578(.A(men_men_n1595_), .Y(men_men_n1609_));
  INV        u1579(.A(men_men_n1487_), .Y(men_men_n1610_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule