//Benchmark atmr_misex3_1774_0.5

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1584_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1592_, men_men_n1593_, men_men_n1594_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, men_men_n1602_, men_men_n1603_, men_men_n1604_, men_men_n1605_, men_men_n1606_, men_men_n1607_, men_men_n1608_, men_men_n1609_, men_men_n1610_, men_men_n1611_, men_men_n1612_, men_men_n1613_, men_men_n1614_, men_men_n1615_, men_men_n1616_, men_men_n1617_, men_men_n1618_, men_men_n1619_, men_men_n1620_, men_men_n1621_, men_men_n1622_, men_men_n1623_, men_men_n1624_, men_men_n1625_, men_men_n1626_, men_men_n1627_, men_men_n1628_, men_men_n1629_, men_men_n1630_, men_men_n1631_, men_men_n1632_, men_men_n1633_, men_men_n1634_, men_men_n1635_, men_men_n1636_, men_men_n1637_, men_men_n1638_, men_men_n1639_, men_men_n1640_, men_men_n1641_, men_men_n1642_, men_men_n1643_, men_men_n1644_, men_men_n1645_, men_men_n1646_, men_men_n1647_, men_men_n1648_, men_men_n1649_, men_men_n1650_, men_men_n1651_, men_men_n1652_, men_men_n1654_, men_men_n1655_, men_men_n1656_, men_men_n1657_, men_men_n1658_, men_men_n1659_, men_men_n1660_, men_men_n1661_, men_men_n1665_, men_men_n1666_, men_men_n1667_, men_men_n1668_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  ZERO       o00(.Y(ori10));
  ZERO       o01(.Y(ori11));
  ZERO       o02(.Y(ori08));
  ZERO       o03(.Y(ori09));
  ZERO       o04(.Y(ori12));
  ZERO       o05(.Y(ori13));
  ZERO       o06(.Y(ori02));
  ZERO       o07(.Y(ori03));
  ZERO       o08(.Y(ori00));
  ZERO       o09(.Y(ori01));
  ZERO       o10(.Y(ori06));
  ZERO       o11(.Y(ori07));
  ONE        o12(.Y(ori04));
  ZERO       o13(.Y(ori05));
  NOi32      m000(.An(m), .Bn(l), .C(n), .Y(mai_mai_n29_));
  NOi32      m001(.An(i), .Bn(m), .C(h), .Y(mai_mai_n30_));
  NA2        m002(.A(mai_mai_n30_), .B(mai_mai_n29_), .Y(mai_mai_n31_));
  INV        m003(.A(h), .Y(mai_mai_n32_));
  NAi21      m004(.An(j), .B(l), .Y(mai_mai_n33_));
  NAi32      m005(.An(n), .Bn(m), .C(m), .Y(mai_mai_n34_));
  NO3        m006(.A(mai_mai_n34_), .B(mai_mai_n33_), .C(mai_mai_n32_), .Y(mai_mai_n35_));
  INV        m007(.A(i), .Y(mai_mai_n36_));
  AN2        m008(.A(h), .B(m), .Y(mai_mai_n37_));
  NAi21      m009(.An(n), .B(m), .Y(mai_mai_n38_));
  INV        m010(.A(c), .Y(mai_mai_n39_));
  NAi21      m011(.An(i), .B(h), .Y(mai_mai_n40_));
  INV        m012(.A(h), .Y(mai_mai_n41_));
  NAi31      m013(.An(n), .B(d), .C(b), .Y(mai_mai_n42_));
  INV        m014(.A(m), .Y(mai_mai_n43_));
  AN4        m015(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n44_));
  NA2        m016(.A(h), .B(mai_mai_n44_), .Y(mai_mai_n45_));
  INV        m017(.A(n), .Y(mai_mai_n46_));
  INV        m018(.A(j), .Y(mai_mai_n47_));
  AN3        m019(.A(m), .B(k), .C(i), .Y(mai_mai_n48_));
  NAi32      m020(.An(m), .Bn(f), .C(h), .Y(mai_mai_n49_));
  NAi31      m021(.An(j), .B(m), .C(l), .Y(mai_mai_n50_));
  NO2        m022(.A(mai_mai_n50_), .B(mai_mai_n49_), .Y(mai_mai_n51_));
  NAi41      m023(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n52_));
  AN2        m024(.A(e), .B(b), .Y(mai_mai_n53_));
  NA2        m025(.A(c), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  INV        m026(.A(a), .Y(mai_mai_n55_));
  INV        m027(.A(l), .Y(mai_mai_n56_));
  NOi21      m028(.An(m), .B(n), .Y(mai_mai_n57_));
  INV        m029(.A(b), .Y(mai_mai_n58_));
  NA2        m030(.A(l), .B(j), .Y(mai_mai_n59_));
  NAi21      m031(.An(m), .B(h), .Y(mai_mai_n60_));
  NAi21      m032(.An(m), .B(n), .Y(mai_mai_n61_));
  NAi21      m033(.An(j), .B(h), .Y(mai_mai_n62_));
  INV        m034(.A(mai_mai_n61_), .Y(mai_mai_n63_));
  NAi21      m035(.An(c), .B(b), .Y(mai_mai_n64_));
  NA2        m036(.A(f), .B(d), .Y(mai_mai_n65_));
  NO3        m037(.A(mai_mai_n65_), .B(mai_mai_n64_), .C(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m038(.A(mai_mai_n66_), .B(mai_mai_n63_), .Y(mai_mai_n67_));
  NA2        m039(.A(d), .B(b), .Y(mai_mai_n68_));
  INV        m040(.A(mai_mai_n68_), .Y(mai_mai_n69_));
  BUFFER     m041(.A(c), .Y(mai_mai_n70_));
  NAi31      m042(.An(l), .B(k), .C(h), .Y(mai_mai_n71_));
  INV        m043(.A(mai_mai_n67_), .Y(mai_mai_n72_));
  NAi31      m044(.An(e), .B(f), .C(b), .Y(mai_mai_n73_));
  INV        m045(.A(mai_mai_n73_), .Y(mai_mai_n74_));
  NOi21      m046(.An(k), .B(m), .Y(mai_mai_n75_));
  NA3        m047(.A(mai_mai_n75_), .B(h), .C(n), .Y(mai_mai_n76_));
  NOi21      m048(.An(mai_mai_n74_), .B(mai_mai_n76_), .Y(mai_mai_n77_));
  NA2        m049(.A(j), .B(h), .Y(mai_mai_n78_));
  OR3        m050(.A(n), .B(m), .C(k), .Y(mai_mai_n79_));
  NO2        m051(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  NAi32      m052(.An(m), .Bn(k), .C(n), .Y(mai_mai_n81_));
  NO2        m053(.A(mai_mai_n81_), .B(mai_mai_n78_), .Y(mai_mai_n82_));
  AOI220     m054(.A0(mai_mai_n82_), .A1(mai_mai_n74_), .B0(mai_mai_n80_), .B1(c), .Y(mai_mai_n83_));
  NO2        m055(.A(n), .B(m), .Y(mai_mai_n84_));
  NA2        m056(.A(d), .B(c), .Y(mai_mai_n85_));
  NAi31      m057(.An(m), .B(n), .C(b), .Y(mai_mai_n86_));
  NO2        m058(.A(mai_mai_n86_), .B(mai_mai_n70_), .Y(mai_mai_n87_));
  INV        m059(.A(mai_mai_n83_), .Y(mai_mai_n88_));
  OR3        m060(.A(mai_mai_n88_), .B(mai_mai_n77_), .C(mai_mai_n72_), .Y(mai_mai_n89_));
  INV        m061(.A(mai_mai_n89_), .Y(mai_mai_n90_));
  NAi31      m062(.An(n), .B(h), .C(m), .Y(mai_mai_n91_));
  NA3        m063(.A(mai_mai_n57_), .B(i), .C(m), .Y(mai_mai_n92_));
  AN2        m064(.A(i), .B(m), .Y(mai_mai_n93_));
  INV        m065(.A(m), .Y(mai_mai_n94_));
  NOi21      m066(.An(l), .B(m), .Y(mai_mai_n95_));
  NOi21      m067(.An(n), .B(m), .Y(mai_mai_n96_));
  NA2        m068(.A(i), .B(mai_mai_n96_), .Y(mai_mai_n97_));
  OA220      m069(.A0(mai_mai_n97_), .A1(mai_mai_n54_), .B0(m), .B1(mai_mai_n45_), .Y(mai_mai_n98_));
  INV        m070(.A(h), .Y(mai_mai_n99_));
  NOi31      m071(.An(k), .B(n), .C(m), .Y(mai_mai_n100_));
  NOi21      m072(.An(mai_mai_n100_), .B(mai_mai_n85_), .Y(mai_mai_n101_));
  INV        m073(.A(mai_mai_n101_), .Y(mai_mai_n102_));
  NAi21      m074(.An(n), .B(a), .Y(mai_mai_n103_));
  NAi41      m075(.An(m), .B(m), .C(k), .D(h), .Y(mai_mai_n104_));
  AN2        m076(.A(mai_mai_n102_), .B(mai_mai_n98_), .Y(mai_mai_n105_));
  NO2        m077(.A(h), .B(mai_mai_n52_), .Y(mai_mai_n106_));
  NA2        m078(.A(mai_mai_n106_), .B(b), .Y(mai_mai_n107_));
  NO2        m079(.A(n), .B(a), .Y(mai_mai_n108_));
  NAi31      m080(.An(mai_mai_n104_), .B(mai_mai_n108_), .C(mai_mai_n53_), .Y(mai_mai_n109_));
  NAi21      m081(.An(h), .B(i), .Y(mai_mai_n110_));
  NA2        m082(.A(mai_mai_n84_), .B(k), .Y(mai_mai_n111_));
  NO2        m083(.A(mai_mai_n111_), .B(mai_mai_n110_), .Y(mai_mai_n112_));
  NA2        m084(.A(mai_mai_n109_), .B(mai_mai_n107_), .Y(mai_mai_n113_));
  NAi21      m085(.An(f), .B(m), .Y(mai_mai_n114_));
  NOi21      m086(.An(mai_mai_n105_), .B(mai_mai_n113_), .Y(mai_mai_n115_));
  NAi21      m087(.An(h), .B(m), .Y(mai_mai_n116_));
  NA2        m088(.A(k), .B(h), .Y(mai_mai_n117_));
  INV        m089(.A(a), .Y(mai_mai_n118_));
  NA3        m090(.A(mai_mai_n75_), .B(h), .C(mai_mai_n46_), .Y(mai_mai_n119_));
  NO2        m091(.A(mai_mai_n119_), .B(mai_mai_n581_), .Y(mai_mai_n120_));
  INV        m092(.A(mai_mai_n120_), .Y(mai_mai_n121_));
  NA3        m093(.A(e), .B(c), .C(b), .Y(mai_mai_n122_));
  NO2        m094(.A(mai_mai_n569_), .B(mai_mai_n42_), .Y(mai_mai_n123_));
  INV        m095(.A(mai_mai_n123_), .Y(mai_mai_n124_));
  NAi32      m096(.An(j), .Bn(h), .C(i), .Y(mai_mai_n125_));
  NAi21      m097(.An(m), .B(l), .Y(mai_mai_n126_));
  NO3        m098(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(mai_mai_n46_), .Y(mai_mai_n127_));
  NA2        m099(.A(h), .B(m), .Y(mai_mai_n128_));
  NA2        m100(.A(mai_mai_n127_), .B(b), .Y(mai_mai_n129_));
  NA3        m101(.A(mai_mai_n129_), .B(mai_mai_n124_), .C(mai_mai_n121_), .Y(mai_mai_n130_));
  NAi32      m102(.An(n), .Bn(m), .C(l), .Y(mai_mai_n131_));
  NO2        m103(.A(mai_mai_n131_), .B(mai_mai_n125_), .Y(mai_mai_n132_));
  INV        m104(.A(mai_mai_n130_), .Y(mai_mai_n133_));
  NAi31      m105(.An(d), .B(c), .C(b), .Y(mai_mai_n134_));
  NAi31      m106(.An(d), .B(e), .C(b), .Y(mai_mai_n135_));
  NO3        m107(.A(mai_mai_n134_), .B(m), .C(mai_mai_n41_), .Y(mai_mai_n136_));
  NA2        m108(.A(mai_mai_n108_), .B(mai_mai_n53_), .Y(mai_mai_n137_));
  NOi31      m109(.An(l), .B(n), .C(m), .Y(mai_mai_n138_));
  NA2        m110(.A(mai_mai_n138_), .B(i), .Y(mai_mai_n139_));
  NO2        m111(.A(mai_mai_n139_), .B(mai_mai_n581_), .Y(mai_mai_n140_));
  OR2        m112(.A(mai_mai_n140_), .B(mai_mai_n136_), .Y(mai_mai_n141_));
  NAi32      m113(.An(m), .Bn(j), .C(k), .Y(mai_mai_n142_));
  NAi41      m114(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n143_));
  AN3        m115(.A(h), .B(m), .C(f), .Y(mai_mai_n144_));
  NAi31      m116(.An(m), .B(mai_mai_n144_), .C(b), .Y(mai_mai_n145_));
  NO2        m117(.A(mai_mai_n126_), .B(mai_mai_n125_), .Y(mai_mai_n146_));
  INV        m118(.A(mai_mai_n145_), .Y(mai_mai_n147_));
  NA2        m119(.A(mai_mai_n92_), .B(mai_mai_n31_), .Y(mai_mai_n148_));
  NA2        m120(.A(mai_mai_n148_), .B(b), .Y(mai_mai_n149_));
  NO2        m121(.A(mai_mai_n135_), .B(n), .Y(mai_mai_n150_));
  NA2        m122(.A(h), .B(mai_mai_n57_), .Y(mai_mai_n151_));
  INV        m123(.A(mai_mai_n151_), .Y(mai_mai_n152_));
  AOI220     m124(.A0(mai_mai_n152_), .A1(b), .B0(m), .B1(mai_mai_n150_), .Y(mai_mai_n153_));
  INV        m125(.A(mai_mai_n153_), .Y(mai_mai_n154_));
  NO4        m126(.A(mai_mai_n154_), .B(mai_mai_n147_), .C(mai_mai_n141_), .D(mai_mai_n112_), .Y(mai_mai_n155_));
  NA4        m127(.A(mai_mai_n155_), .B(mai_mai_n133_), .C(mai_mai_n115_), .D(mai_mai_n90_), .Y(mai10));
  NA2        m128(.A(h), .B(mai_mai_n96_), .Y(mai_mai_n157_));
  INV        m129(.A(mai_mai_n76_), .Y(mai_mai_n158_));
  NA2        m130(.A(mai_mai_n158_), .B(c), .Y(mai_mai_n159_));
  NO2        m131(.A(mai_mai_n78_), .B(m), .Y(mai_mai_n160_));
  NA3        m132(.A(n), .B(f), .C(c), .Y(mai_mai_n161_));
  NOi21      m133(.An(mai_mai_n160_), .B(mai_mai_n161_), .Y(mai_mai_n162_));
  INV        m134(.A(mai_mai_n162_), .Y(mai_mai_n163_));
  NO2        m135(.A(mai_mai_n161_), .B(mai_mai_n126_), .Y(mai_mai_n164_));
  AOI220     m136(.A0(d), .A1(mai_mai_n132_), .B0(mai_mai_n164_), .B1(i), .Y(mai_mai_n165_));
  NA3        m137(.A(mai_mai_n165_), .B(mai_mai_n163_), .C(mai_mai_n159_), .Y(mai_mai_n166_));
  NA2        m138(.A(mai_mai_n108_), .B(b), .Y(mai_mai_n167_));
  INV        m139(.A(e), .Y(mai_mai_n168_));
  NA2        m140(.A(m), .B(m), .Y(mai_mai_n169_));
  NO2        m141(.A(mai_mai_n169_), .B(mai_mai_n167_), .Y(mai_mai_n170_));
  NAi31      m142(.An(b), .B(c), .C(a), .Y(mai_mai_n171_));
  NO2        m143(.A(mai_mai_n171_), .B(n), .Y(mai_mai_n172_));
  NA2        m144(.A(h), .B(m), .Y(mai_mai_n173_));
  NO2        m145(.A(mai_mai_n170_), .B(mai_mai_n166_), .Y(mai_mai_n174_));
  NOi21      m146(.An(a), .B(n), .Y(mai_mai_n175_));
  NA2        m147(.A(d), .B(mai_mai_n175_), .Y(mai_mai_n176_));
  NA2        m148(.A(m), .B(m), .Y(mai_mai_n177_));
  NO2        m149(.A(mai_mai_n177_), .B(mai_mai_n176_), .Y(mai_mai_n178_));
  INV        m150(.A(mai_mai_n178_), .Y(mai_mai_n179_));
  OR2        m151(.A(n), .B(m), .Y(mai_mai_n180_));
  NO2        m152(.A(mai_mai_n180_), .B(mai_mai_n71_), .Y(mai_mai_n181_));
  INV        m153(.A(mai_mai_n80_), .Y(mai_mai_n182_));
  INV        m154(.A(mai_mai_n151_), .Y(mai_mai_n183_));
  NA3        m155(.A(mai_mai_n183_), .B(b), .C(d), .Y(mai_mai_n184_));
  NAi21      m156(.An(k), .B(j), .Y(mai_mai_n185_));
  INV        m157(.A(mai_mai_n111_), .Y(mai_mai_n186_));
  NA2        m158(.A(mai_mai_n186_), .B(d), .Y(mai_mai_n187_));
  NA3        m159(.A(mai_mai_n187_), .B(mai_mai_n184_), .C(mai_mai_n182_), .Y(mai_mai_n188_));
  INV        m160(.A(mai_mai_n139_), .Y(mai_mai_n189_));
  NOi21      m161(.An(mai_mai_n179_), .B(mai_mai_n188_), .Y(mai_mai_n190_));
  NOi32      m162(.An(c), .Bn(a), .C(b), .Y(mai_mai_n191_));
  NA2        m163(.A(mai_mai_n191_), .B(mai_mai_n57_), .Y(mai_mai_n192_));
  INV        m164(.A(m), .Y(mai_mai_n193_));
  AOI210     m165(.A0(mai_mai_n193_), .A1(mai_mai_n117_), .B0(mai_mai_n192_), .Y(mai_mai_n194_));
  NO4        m166(.A(h), .B(mai_mai_n52_), .C(mai_mai_n39_), .D(b), .Y(mai_mai_n195_));
  NO3        m167(.A(n), .B(mai_mai_n50_), .C(mai_mai_n60_), .Y(mai_mai_n196_));
  NO3        m168(.A(mai_mai_n196_), .B(mai_mai_n195_), .C(mai_mai_n194_), .Y(mai_mai_n197_));
  NOi21      m169(.An(d), .B(e), .Y(mai_mai_n198_));
  INV        m170(.A(mai_mai_n52_), .Y(mai_mai_n199_));
  NA3        m171(.A(mai_mai_n199_), .B(c), .C(b), .Y(mai_mai_n200_));
  NO2        m172(.A(mai_mai_n583_), .B(mai_mai_n151_), .Y(mai_mai_n201_));
  INV        m173(.A(mai_mai_n201_), .Y(mai_mai_n202_));
  NA3        m174(.A(mai_mai_n202_), .B(mai_mai_n200_), .C(mai_mai_n105_), .Y(mai_mai_n203_));
  NO2        m175(.A(m), .B(mai_mai_n60_), .Y(mai_mai_n204_));
  XO2        m176(.A(i), .B(h), .Y(mai_mai_n205_));
  NA3        m177(.A(mai_mai_n205_), .B(mai_mai_n75_), .C(n), .Y(mai_mai_n206_));
  NAi31      m178(.An(mai_mai_n127_), .B(mai_mai_n206_), .C(mai_mai_n157_), .Y(mai_mai_n207_));
  NA2        m179(.A(mai_mai_n100_), .B(i), .Y(mai_mai_n208_));
  NA2        m180(.A(m), .B(l), .Y(mai_mai_n209_));
  INV        m181(.A(mai_mai_n203_), .Y(mai_mai_n210_));
  NA4        m182(.A(mai_mai_n210_), .B(mai_mai_n197_), .C(mai_mai_n190_), .D(mai_mai_n174_), .Y(mai11));
  NO2        m183(.A(mai_mai_n42_), .B(f), .Y(mai_mai_n212_));
  NA2        m184(.A(j), .B(m), .Y(mai_mai_n213_));
  NA2        m185(.A(k), .B(j), .Y(mai_mai_n214_));
  NA2        m186(.A(m), .B(mai_mai_n212_), .Y(mai_mai_n215_));
  NA2        m187(.A(mai_mai_n37_), .B(j), .Y(mai_mai_n216_));
  NO2        m188(.A(mai_mai_n216_), .B(m), .Y(mai_mai_n217_));
  NAi31      m189(.An(d), .B(e), .C(a), .Y(mai_mai_n218_));
  NO2        m190(.A(mai_mai_n218_), .B(n), .Y(mai_mai_n219_));
  NA2        m191(.A(mai_mai_n217_), .B(b), .Y(mai_mai_n220_));
  NAi31      m192(.An(n), .B(m), .C(k), .Y(mai_mai_n221_));
  NO4        m193(.A(n), .B(d), .C(mai_mai_n58_), .D(a), .Y(mai_mai_n222_));
  INV        m194(.A(mai_mai_n222_), .Y(mai_mai_n223_));
  NO2        m195(.A(mai_mai_n60_), .B(mai_mai_n223_), .Y(mai_mai_n224_));
  INV        m196(.A(mai_mai_n224_), .Y(mai_mai_n225_));
  NA2        m197(.A(k), .B(mai_mai_n30_), .Y(mai_mai_n226_));
  NO2        m198(.A(mai_mai_n216_), .B(m), .Y(mai_mai_n227_));
  NAi21      m199(.An(b), .B(c), .Y(mai_mai_n228_));
  BUFFER     m200(.A(mai_mai_n143_), .Y(mai_mai_n229_));
  NA2        m201(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n230_));
  OA210      m202(.A0(mai_mai_n230_), .A1(c), .B0(mai_mai_n227_), .Y(mai_mai_n231_));
  NO3        m203(.A(i), .B(mai_mai_n38_), .C(mai_mai_n94_), .Y(mai_mai_n232_));
  NA2        m204(.A(mai_mai_n232_), .B(a), .Y(mai_mai_n233_));
  INV        m205(.A(mai_mai_n233_), .Y(mai_mai_n234_));
  NAi32      m206(.An(d), .Bn(a), .C(b), .Y(mai_mai_n235_));
  NO3        m207(.A(mai_mai_n81_), .B(mai_mai_n78_), .C(m), .Y(mai_mai_n236_));
  NA3        m208(.A(f), .B(d), .C(b), .Y(mai_mai_n237_));
  NO3        m209(.A(mai_mai_n236_), .B(mai_mai_n234_), .C(mai_mai_n231_), .Y(mai_mai_n238_));
  AN4        m210(.A(mai_mai_n238_), .B(mai_mai_n225_), .C(mai_mai_n220_), .D(mai_mai_n215_), .Y(mai_mai_n239_));
  NA3        m211(.A(a), .B(m), .C(mai_mai_n57_), .Y(mai_mai_n240_));
  NAi32      m212(.An(h), .Bn(f), .C(m), .Y(mai_mai_n241_));
  NAi41      m213(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n242_));
  OAI210     m214(.A0(mai_mai_n218_), .A1(n), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  NA2        m215(.A(mai_mai_n243_), .B(m), .Y(mai_mai_n244_));
  NAi21      m216(.An(h), .B(m), .Y(mai_mai_n245_));
  OR2        m217(.A(mai_mai_n244_), .B(mai_mai_n241_), .Y(mai_mai_n246_));
  NO2        m218(.A(mai_mai_n241_), .B(mai_mai_n42_), .Y(mai_mai_n247_));
  NAi31      m219(.An(mai_mai_n247_), .B(mai_mai_n246_), .C(mai_mai_n240_), .Y(mai_mai_n248_));
  NAi21      m220(.An(f), .B(h), .Y(mai_mai_n249_));
  NO2        m221(.A(n), .B(c), .Y(mai_mai_n250_));
  INV        m222(.A(mai_mai_n248_), .Y(mai_mai_n251_));
  NO3        m223(.A(m), .B(mai_mai_n40_), .C(n), .Y(mai_mai_n252_));
  NA2        m224(.A(k), .B(mai_mai_n57_), .Y(mai_mai_n253_));
  INV        m225(.A(mai_mai_n252_), .Y(mai_mai_n254_));
  NO2        m226(.A(mai_mai_n254_), .B(mai_mai_n47_), .Y(mai_mai_n255_));
  OR2        m227(.A(mai_mai_n114_), .B(mai_mai_n244_), .Y(mai_mai_n256_));
  NO2        m228(.A(mai_mai_n583_), .B(mai_mai_n128_), .Y(mai_mai_n257_));
  NAi21      m229(.An(n), .B(mai_mai_n257_), .Y(mai_mai_n258_));
  NA2        m230(.A(mai_mai_n258_), .B(mai_mai_n256_), .Y(mai_mai_n259_));
  NO2        m231(.A(mai_mai_n573_), .B(n), .Y(mai_mai_n260_));
  NA2        m232(.A(mai_mai_n260_), .B(m), .Y(mai_mai_n261_));
  NA2        m233(.A(mai_mai_n205_), .B(mai_mai_n75_), .Y(mai_mai_n262_));
  NO3        m234(.A(mai_mai_n161_), .B(mai_mai_n262_), .C(mai_mai_n47_), .Y(mai_mai_n263_));
  INV        m235(.A(mai_mai_n263_), .Y(mai_mai_n264_));
  AN2        m236(.A(d), .B(b), .Y(mai_mai_n265_));
  NA2        m237(.A(mai_mai_n75_), .B(mai_mai_n94_), .Y(mai_mai_n266_));
  NO2        m238(.A(mai_mai_n584_), .B(mai_mai_n266_), .Y(mai_mai_n267_));
  NAi31      m239(.An(m), .B(n), .C(k), .Y(mai_mai_n268_));
  INV        m240(.A(mai_mai_n109_), .Y(mai_mai_n269_));
  OAI210     m241(.A0(mai_mai_n269_), .A1(mai_mai_n267_), .B0(j), .Y(mai_mai_n270_));
  NA3        m242(.A(mai_mai_n270_), .B(mai_mai_n264_), .C(mai_mai_n261_), .Y(mai_mai_n271_));
  NO3        m243(.A(mai_mai_n271_), .B(mai_mai_n80_), .C(mai_mai_n255_), .Y(mai_mai_n272_));
  NAi31      m244(.An(m), .B(h), .C(f), .Y(mai_mai_n273_));
  NA3        m245(.A(h), .B(a), .C(mai_mai_n46_), .Y(mai_mai_n274_));
  INV        m246(.A(mai_mai_n274_), .Y(mai_mai_n275_));
  NO2        m247(.A(mai_mai_n274_), .B(mai_mai_n214_), .Y(mai_mai_n276_));
  NO2        m248(.A(mai_mai_n208_), .B(mai_mai_n47_), .Y(mai_mai_n277_));
  NA2        m249(.A(h), .B(m), .Y(mai_mai_n278_));
  NO2        m250(.A(mai_mai_n235_), .B(mai_mai_n38_), .Y(mai_mai_n279_));
  INV        m251(.A(mai_mai_n61_), .Y(mai_mai_n280_));
  OR2        m252(.A(mai_mai_n61_), .B(mai_mai_n226_), .Y(mai_mai_n281_));
  INV        m253(.A(mai_mai_n281_), .Y(mai_mai_n282_));
  NO3        m254(.A(m), .B(mai_mai_n78_), .C(i), .Y(mai_mai_n283_));
  NA2        m255(.A(mai_mai_n191_), .B(mai_mai_n46_), .Y(mai_mai_n284_));
  NO3        m256(.A(mai_mai_n282_), .B(mai_mai_n277_), .C(mai_mai_n276_), .Y(mai_mai_n285_));
  NA4        m257(.A(mai_mai_n285_), .B(mai_mai_n272_), .C(mai_mai_n251_), .D(mai_mai_n239_), .Y(mai08));
  NO2        m258(.A(k), .B(h), .Y(mai_mai_n287_));
  NO2        m259(.A(mai_mai_n575_), .B(mai_mai_n126_), .Y(mai_mai_n288_));
  NA2        m260(.A(c), .B(mai_mai_n288_), .Y(mai_mai_n289_));
  AOI210     m261(.A0(mai_mai_n237_), .A1(mai_mai_n73_), .B0(mai_mai_n46_), .Y(mai_mai_n290_));
  NA2        m262(.A(mai_mai_n95_), .B(mai_mai_n290_), .Y(mai_mai_n291_));
  NA2        m263(.A(mai_mai_n291_), .B(mai_mai_n289_), .Y(mai_mai_n292_));
  NA2        m264(.A(b), .B(mai_mai_n35_), .Y(mai_mai_n293_));
  NA2        m265(.A(mai_mai_n138_), .B(h), .Y(mai_mai_n294_));
  NA2        m266(.A(l), .B(mai_mai_n96_), .Y(mai_mai_n295_));
  NO2        m267(.A(mai_mai_n295_), .B(mai_mai_n135_), .Y(mai_mai_n296_));
  NA2        m268(.A(mai_mai_n296_), .B(i), .Y(mai_mai_n297_));
  NA3        m269(.A(m), .B(l), .C(k), .Y(mai_mai_n298_));
  NO2        m270(.A(mai_mai_n274_), .B(mai_mai_n298_), .Y(mai_mai_n299_));
  INV        m271(.A(mai_mai_n299_), .Y(mai_mai_n300_));
  NA4        m272(.A(mai_mai_n300_), .B(mai_mai_n297_), .C(mai_mai_n294_), .D(mai_mai_n293_), .Y(mai_mai_n301_));
  NO2        m273(.A(mai_mai_n301_), .B(mai_mai_n292_), .Y(mai_mai_n302_));
  INV        m274(.A(mai_mai_n109_), .Y(mai_mai_n303_));
  NA2        m275(.A(l), .B(mai_mai_n43_), .Y(mai_mai_n304_));
  NO2        m276(.A(mai_mai_n579_), .B(mai_mai_n304_), .Y(mai_mai_n305_));
  AOI210     m277(.A0(mai_mai_n303_), .A1(l), .B0(mai_mai_n305_), .Y(mai_mai_n306_));
  INV        m278(.A(mai_mai_n29_), .Y(mai_mai_n307_));
  NO2        m279(.A(mai_mai_n38_), .B(mai_mai_n55_), .Y(mai_mai_n308_));
  NO2        m280(.A(mai_mai_n126_), .B(mai_mai_n32_), .Y(mai_mai_n309_));
  AN3        m281(.A(b), .B(mai_mai_n309_), .C(m), .Y(mai_mai_n310_));
  NA2        m282(.A(mai_mai_n51_), .B(mai_mai_n46_), .Y(mai_mai_n311_));
  INV        m283(.A(mai_mai_n311_), .Y(mai_mai_n312_));
  NO2        m284(.A(mai_mai_n126_), .B(mai_mai_n62_), .Y(mai_mai_n313_));
  NA2        m285(.A(mai_mai_n313_), .B(b), .Y(mai_mai_n314_));
  INV        m286(.A(mai_mai_n314_), .Y(mai_mai_n315_));
  OR3        m287(.A(mai_mai_n315_), .B(mai_mai_n312_), .C(mai_mai_n310_), .Y(mai_mai_n316_));
  NA3        m288(.A(mai_mai_n95_), .B(mai_mai_n185_), .C(mai_mai_n30_), .Y(mai_mai_n317_));
  OAI210     m289(.A0(mai_mai_n298_), .A1(mai_mai_n273_), .B0(mai_mai_n209_), .Y(mai_mai_n318_));
  NA2        m290(.A(mai_mai_n108_), .B(b), .Y(mai_mai_n319_));
  AOI220     m291(.A0(mai_mai_n250_), .A1(a), .B0(mai_mai_n191_), .B1(mai_mai_n46_), .Y(mai_mai_n320_));
  NA2        m292(.A(mai_mai_n320_), .B(mai_mai_n319_), .Y(mai_mai_n321_));
  NA2        m293(.A(mai_mai_n321_), .B(mai_mai_n318_), .Y(mai_mai_n322_));
  INV        m294(.A(mai_mai_n322_), .Y(mai_mai_n323_));
  NO3        m295(.A(mai_mai_n323_), .B(mai_mai_n582_), .C(mai_mai_n316_), .Y(mai_mai_n324_));
  NO3        m296(.A(m), .B(mai_mai_n128_), .C(mai_mai_n56_), .Y(mai_mai_n325_));
  NO3        m297(.A(mai_mai_n572_), .B(mai_mai_n307_), .C(mai_mai_n118_), .Y(mai_mai_n326_));
  OR2        m298(.A(mai_mai_n273_), .B(mai_mai_n50_), .Y(mai_mai_n327_));
  NO2        m299(.A(mai_mai_n570_), .B(n), .Y(mai_mai_n328_));
  NO2        m300(.A(mai_mai_n320_), .B(mai_mai_n327_), .Y(mai_mai_n329_));
  NA2        m301(.A(mai_mai_n325_), .B(c), .Y(mai_mai_n330_));
  INV        m302(.A(mai_mai_n330_), .Y(mai_mai_n331_));
  INV        m303(.A(n), .Y(mai_mai_n332_));
  AOI220     m304(.A0(mai_mai_n313_), .A1(c), .B0(mai_mai_n332_), .B1(mai_mai_n288_), .Y(mai_mai_n333_));
  INV        m305(.A(mai_mai_n103_), .Y(mai_mai_n334_));
  NA2        m306(.A(mai_mai_n51_), .B(mai_mai_n334_), .Y(mai_mai_n335_));
  INV        m307(.A(mai_mai_n335_), .Y(mai_mai_n336_));
  INV        m308(.A(mai_mai_n333_), .Y(mai_mai_n337_));
  NO4        m309(.A(mai_mai_n337_), .B(mai_mai_n331_), .C(mai_mai_n329_), .D(mai_mai_n326_), .Y(mai_mai_n338_));
  NA4        m310(.A(mai_mai_n338_), .B(mai_mai_n324_), .C(mai_mai_n306_), .D(mai_mai_n302_), .Y(mai09));
  NO2        m311(.A(m), .B(m), .Y(mai_mai_n340_));
  INV        m312(.A(mai_mai_n340_), .Y(mai_mai_n341_));
  NA2        m313(.A(mai_mai_n181_), .B(e), .Y(mai_mai_n342_));
  NA3        m314(.A(mai_mai_n48_), .B(m), .C(f), .Y(mai_mai_n343_));
  INV        m315(.A(mai_mai_n327_), .Y(mai_mai_n344_));
  AN2        m316(.A(mai_mai_n344_), .B(mai_mai_n328_), .Y(mai_mai_n345_));
  INV        m317(.A(mai_mai_n143_), .Y(mai_mai_n346_));
  AOI210     m318(.A0(m), .A1(m), .B0(mai_mai_n249_), .Y(mai_mai_n347_));
  NA2        m319(.A(mai_mai_n319_), .B(mai_mai_n137_), .Y(mai_mai_n348_));
  AOI220     m320(.A0(m), .A1(mai_mai_n348_), .B0(mai_mai_n347_), .B1(mai_mai_n346_), .Y(mai_mai_n349_));
  NA3        m321(.A(mai_mai_n571_), .B(mai_mai_n87_), .C(e), .Y(mai_mai_n350_));
  NA2        m322(.A(mai_mai_n350_), .B(mai_mai_n349_), .Y(mai_mai_n351_));
  NA3        m323(.A(a), .B(f), .C(mai_mai_n46_), .Y(mai_mai_n352_));
  NO2        m324(.A(mai_mai_n268_), .B(mai_mai_n135_), .Y(mai_mai_n353_));
  AN2        m325(.A(mai_mai_n353_), .B(i), .Y(mai_mai_n354_));
  NA2        m326(.A(mai_mai_n75_), .B(i), .Y(mai_mai_n355_));
  OAI220     m327(.A0(mai_mai_n352_), .A1(mai_mai_n173_), .B0(mai_mai_n143_), .B1(mai_mai_n355_), .Y(mai_mai_n356_));
  NOi21      m328(.An(mai_mai_n98_), .B(mai_mai_n356_), .Y(mai_mai_n357_));
  INV        m329(.A(c), .Y(mai_mai_n358_));
  NO2        m330(.A(mai_mai_n358_), .B(mai_mai_n168_), .Y(mai_mai_n359_));
  NA2        m331(.A(mai_mai_n359_), .B(mai_mai_n207_), .Y(mai_mai_n360_));
  OR2        m332(.A(mai_mai_n273_), .B(mai_mai_n221_), .Y(mai_mai_n361_));
  NA3        m333(.A(mai_mai_n361_), .B(mai_mai_n360_), .C(mai_mai_n357_), .Y(mai_mai_n362_));
  NO3        m334(.A(mai_mai_n362_), .B(mai_mai_n351_), .C(mai_mai_n345_), .Y(mai_mai_n363_));
  BUFFER     m335(.A(mai_mai_n352_), .Y(mai_mai_n364_));
  INV        m336(.A(m), .Y(mai_mai_n365_));
  NO2        m337(.A(mai_mai_n365_), .B(mai_mai_n364_), .Y(mai_mai_n366_));
  INV        m338(.A(mai_mai_n173_), .Y(mai_mai_n367_));
  NA2        m339(.A(e), .B(d), .Y(mai_mai_n368_));
  NA3        m340(.A(e), .B(mai_mai_n186_), .C(mai_mai_n205_), .Y(mai_mai_n369_));
  NO2        m341(.A(mai_mai_n208_), .B(f), .Y(mai_mai_n370_));
  AOI210     m342(.A0(b), .A1(mai_mai_n146_), .B0(mai_mai_n370_), .Y(mai_mai_n371_));
  NA2        m343(.A(mai_mai_n371_), .B(mai_mai_n369_), .Y(mai_mai_n372_));
  NO2        m344(.A(mai_mai_n372_), .B(mai_mai_n366_), .Y(mai_mai_n373_));
  AOI220     m345(.A0(h), .A1(mai_mai_n353_), .B0(mai_mai_n252_), .B1(e), .Y(mai_mai_n374_));
  OAI210     m346(.A0(mai_mai_n80_), .A1(mai_mai_n189_), .B0(e), .Y(mai_mai_n375_));
  AN2        m347(.A(mai_mai_n375_), .B(mai_mai_n374_), .Y(mai_mai_n376_));
  NA4        m348(.A(mai_mai_n376_), .B(mai_mai_n373_), .C(mai_mai_n363_), .D(mai_mai_n342_), .Y(mai12));
  NO3        m349(.A(mai_mai_n180_), .B(mai_mai_n110_), .C(mai_mai_n94_), .Y(mai_mai_n378_));
  INV        m350(.A(mai_mai_n378_), .Y(mai_mai_n379_));
  NA2        m351(.A(h), .B(mai_mai_n222_), .Y(mai_mai_n380_));
  NA3        m352(.A(mai_mai_n380_), .B(mai_mai_n379_), .C(mai_mai_n179_), .Y(mai_mai_n381_));
  NO2        m353(.A(m), .B(mai_mai_n91_), .Y(mai_mai_n382_));
  INV        m354(.A(mai_mai_n103_), .Y(mai_mai_n383_));
  NO3        m355(.A(mai_mai_n274_), .B(mai_mai_n50_), .C(mai_mai_n36_), .Y(mai_mai_n384_));
  NO2        m356(.A(mai_mai_n384_), .B(mai_mai_n381_), .Y(mai_mai_n385_));
  INV        m357(.A(mai_mai_n242_), .Y(mai_mai_n386_));
  NOi21      m358(.An(mai_mai_n30_), .B(mai_mai_n268_), .Y(mai_mai_n387_));
  NA2        m359(.A(mai_mai_n386_), .B(mai_mai_n93_), .Y(mai_mai_n388_));
  INV        m360(.A(mai_mai_n388_), .Y(mai_mai_n389_));
  NO2        m361(.A(m), .B(mai_mai_n128_), .Y(mai_mai_n390_));
  INV        m362(.A(mai_mai_n149_), .Y(mai_mai_n391_));
  NO2        m363(.A(mai_mai_n391_), .B(mai_mai_n389_), .Y(mai_mai_n392_));
  NA2        m364(.A(mai_mai_n146_), .B(m), .Y(mai_mai_n393_));
  NA2        m365(.A(h), .B(i), .Y(mai_mai_n394_));
  OAI210     m366(.A0(mai_mai_n394_), .A1(mai_mai_n137_), .B0(mai_mai_n393_), .Y(mai_mai_n395_));
  OAI210     m367(.A0(mai_mai_n144_), .A1(h), .B0(mai_mai_n279_), .Y(mai_mai_n396_));
  NA2        m368(.A(a), .B(mai_mai_n57_), .Y(mai_mai_n397_));
  NA2        m369(.A(m), .B(i), .Y(mai_mai_n398_));
  OR2        m370(.A(mai_mai_n398_), .B(mai_mai_n397_), .Y(mai_mai_n399_));
  NO2        m371(.A(mai_mai_n278_), .B(m), .Y(mai_mai_n400_));
  INV        m372(.A(mai_mai_n343_), .Y(mai_mai_n401_));
  NA2        m373(.A(mai_mai_n401_), .B(mai_mai_n191_), .Y(mai_mai_n402_));
  NA3        m374(.A(mai_mai_n402_), .B(mai_mai_n399_), .C(mai_mai_n396_), .Y(mai_mai_n403_));
  NA2        m375(.A(mai_mai_n275_), .B(mai_mai_n48_), .Y(mai_mai_n404_));
  INV        m376(.A(mai_mai_n404_), .Y(mai_mai_n405_));
  NA2        m377(.A(mai_mai_n93_), .B(mai_mai_n219_), .Y(mai_mai_n406_));
  NA2        m378(.A(mai_mai_n400_), .B(b), .Y(mai_mai_n407_));
  NA2        m379(.A(mai_mai_n407_), .B(mai_mai_n406_), .Y(mai_mai_n408_));
  NO4        m380(.A(mai_mai_n408_), .B(mai_mai_n405_), .C(mai_mai_n403_), .D(mai_mai_n395_), .Y(mai_mai_n409_));
  INV        m381(.A(mai_mai_n116_), .Y(mai_mai_n410_));
  NA2        m382(.A(mai_mai_n410_), .B(mai_mai_n199_), .Y(mai_mai_n411_));
  INV        m383(.A(mai_mai_n411_), .Y(mai_mai_n412_));
  INV        m384(.A(mai_mai_n382_), .Y(mai_mai_n413_));
  NA2        m385(.A(mai_mai_n172_), .B(m), .Y(mai_mai_n414_));
  NA2        m386(.A(mai_mai_n414_), .B(mai_mai_n413_), .Y(mai_mai_n415_));
  NA3        m387(.A(c), .B(mai_mai_n576_), .C(mai_mai_n37_), .Y(mai_mai_n416_));
  OR2        m388(.A(mai_mai_n578_), .B(mai_mai_n415_), .Y(mai_mai_n417_));
  NO2        m389(.A(mai_mai_n417_), .B(mai_mai_n412_), .Y(mai_mai_n418_));
  NA4        m390(.A(mai_mai_n418_), .B(mai_mai_n409_), .C(mai_mai_n392_), .D(mai_mai_n385_), .Y(mai13));
  NA3        m391(.A(mai_mai_n108_), .B(b), .C(m), .Y(mai_mai_n420_));
  NA2        m392(.A(mai_mai_n198_), .B(f), .Y(mai_mai_n421_));
  NO4        m393(.A(mai_mai_n421_), .B(mai_mai_n420_), .C(j), .D(k), .Y(mai_mai_n422_));
  NO4        m394(.A(mai_mai_n59_), .B(mai_mai_n421_), .C(mai_mai_n394_), .D(a), .Y(mai_mai_n423_));
  NO3        m395(.A(d), .B(mai_mai_n245_), .C(mai_mai_n131_), .Y(mai_mai_n424_));
  AN2        m396(.A(d), .B(c), .Y(mai_mai_n425_));
  NA2        m397(.A(mai_mai_n425_), .B(mai_mai_n58_), .Y(mai_mai_n426_));
  NO3        m398(.A(mai_mai_n426_), .B(f), .C(mai_mai_n81_), .Y(mai_mai_n427_));
  NO2        m399(.A(mai_mai_n241_), .B(mai_mai_n131_), .Y(mai_mai_n428_));
  OR2        m400(.A(mai_mai_n427_), .B(mai_mai_n428_), .Y(mai_mai_n429_));
  OR4        m401(.A(mai_mai_n429_), .B(mai_mai_n424_), .C(mai_mai_n423_), .D(mai_mai_n422_), .Y(mai_mai_n430_));
  NO2        m402(.A(e), .B(mai_mai_n68_), .Y(mai_mai_n431_));
  NA2        m403(.A(mai_mai_n431_), .B(m), .Y(mai_mai_n432_));
  NO2        m404(.A(mai_mai_n81_), .B(mai_mai_n432_), .Y(mai_mai_n433_));
  NO2        m405(.A(e), .B(mai_mai_n131_), .Y(mai_mai_n434_));
  NOi21      m406(.An(mai_mai_n434_), .B(mai_mai_n114_), .Y(mai_mai_n435_));
  NOi41      m407(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n436_));
  NA2        m408(.A(mai_mai_n436_), .B(j), .Y(mai_mai_n437_));
  NO2        m409(.A(mai_mai_n437_), .B(mai_mai_n432_), .Y(mai_mai_n438_));
  NA3        m410(.A(k), .B(j), .C(i), .Y(mai_mai_n439_));
  NO2        m411(.A(mai_mai_n131_), .B(mai_mai_n49_), .Y(mai_mai_n440_));
  BUFFER     m412(.A(mai_mai_n440_), .Y(mai_mai_n441_));
  OR4        m413(.A(mai_mai_n441_), .B(mai_mai_n438_), .C(mai_mai_n435_), .D(mai_mai_n433_), .Y(mai_mai_n442_));
  INV        m414(.A(mai_mai_n138_), .Y(mai_mai_n443_));
  NO2        m415(.A(mai_mai_n443_), .B(mai_mai_n114_), .Y(mai_mai_n444_));
  NO3        m416(.A(mai_mai_n443_), .B(mai_mai_n241_), .C(mai_mai_n36_), .Y(mai_mai_n445_));
  NO2        m417(.A(f), .B(c), .Y(mai_mai_n446_));
  NOi21      m418(.An(mai_mai_n446_), .B(mai_mai_n180_), .Y(mai_mai_n447_));
  INV        m419(.A(mai_mai_n447_), .Y(mai_mai_n448_));
  OR3        m420(.A(mai_mai_n447_), .B(mai_mai_n442_), .C(mai_mai_n430_), .Y(mai02));
  OR3        m421(.A(n), .B(m), .C(i), .Y(mai_mai_n450_));
  NO4        m422(.A(mai_mai_n450_), .B(h), .C(l), .D(c), .Y(mai_mai_n451_));
  NO2        m423(.A(mai_mai_n440_), .B(mai_mai_n424_), .Y(mai_mai_n452_));
  NA3        m424(.A(m), .B(e), .C(h), .Y(mai_mai_n453_));
  BUFFER     m425(.A(mai_mai_n131_), .Y(mai_mai_n454_));
  OR2        m426(.A(mai_mai_n454_), .B(mai_mai_n453_), .Y(mai_mai_n455_));
  NO2        m427(.A(mai_mai_n443_), .B(mai_mai_n241_), .Y(mai_mai_n456_));
  NO2        m428(.A(mai_mai_n456_), .B(mai_mai_n433_), .Y(mai_mai_n457_));
  NA2        m429(.A(i), .B(h), .Y(mai_mai_n458_));
  INV        m430(.A(mai_mai_n61_), .Y(mai_mai_n459_));
  NO2        m431(.A(mai_mai_n65_), .B(mai_mai_n122_), .Y(mai_mai_n460_));
  NA2        m432(.A(mai_mai_n460_), .B(mai_mai_n459_), .Y(mai_mai_n461_));
  NA2        m433(.A(c), .B(b), .Y(mai_mai_n462_));
  NO2        m434(.A(mai_mai_n462_), .B(mai_mai_n368_), .Y(mai_mai_n463_));
  NO2        m435(.A(mai_mai_n439_), .B(mai_mai_n38_), .Y(mai_mai_n464_));
  AOI210     m436(.A0(mai_mai_n464_), .A1(mai_mai_n463_), .B0(mai_mai_n444_), .Y(mai_mai_n465_));
  AN4        m437(.A(mai_mai_n465_), .B(mai_mai_n461_), .C(mai_mai_n457_), .D(mai_mai_n455_), .Y(mai_mai_n466_));
  NO2        m438(.A(mai_mai_n426_), .B(f), .Y(mai_mai_n467_));
  NA2        m439(.A(mai_mai_n437_), .B(mai_mai_n81_), .Y(mai_mai_n468_));
  AOI210     m440(.A0(mai_mai_n468_), .A1(mai_mai_n467_), .B0(mai_mai_n422_), .Y(mai_mai_n469_));
  NAi41      m441(.An(mai_mai_n451_), .B(mai_mai_n469_), .C(mai_mai_n466_), .D(mai_mai_n452_), .Y(mai03));
  INV        m442(.A(mai_mai_n93_), .Y(mai_mai_n471_));
  NOi21      m443(.An(mai_mai_n327_), .B(m), .Y(mai_mai_n472_));
  OAI220     m444(.A0(mai_mai_n472_), .A1(mai_mai_n284_), .B0(mai_mai_n471_), .B1(mai_mai_n242_), .Y(mai_mai_n473_));
  NA4        m445(.A(i), .B(e), .C(mai_mai_n144_), .D(mai_mai_n138_), .Y(mai_mai_n474_));
  INV        m446(.A(mai_mai_n474_), .Y(mai_mai_n475_));
  NOi31      m447(.An(m), .B(n), .C(f), .Y(mai_mai_n476_));
  NA2        m448(.A(mai_mai_n476_), .B(h), .Y(mai_mai_n477_));
  NA2        m449(.A(c), .B(a), .Y(mai_mai_n478_));
  OAI220     m450(.A0(mai_mai_n478_), .A1(mai_mai_n477_), .B0(mai_mai_n361_), .B1(mai_mai_n171_), .Y(mai_mai_n479_));
  NO2        m451(.A(mai_mai_n479_), .B(mai_mai_n475_), .Y(mai_mai_n480_));
  INV        m452(.A(mai_mai_n424_), .Y(mai_mai_n481_));
  NA3        m453(.A(mai_mai_n448_), .B(mai_mai_n481_), .C(mai_mai_n480_), .Y(mai_mai_n482_));
  NO4        m454(.A(mai_mai_n482_), .B(mai_mai_n473_), .C(mai_mai_n336_), .D(mai_mai_n234_), .Y(mai_mai_n483_));
  NA2        m455(.A(c), .B(b), .Y(mai_mai_n484_));
  NO2        m456(.A(n), .B(mai_mai_n484_), .Y(mai_mai_n485_));
  OAI210     m457(.A0(m), .A1(h), .B0(mai_mai_n485_), .Y(mai_mai_n486_));
  NA2        m458(.A(mai_mai_n486_), .B(mai_mai_n483_), .Y(mai00));
  AOI210     m459(.A0(mai_mai_n367_), .A1(mai_mai_n383_), .B0(mai_mai_n475_), .Y(mai_mai_n488_));
  NA2        m460(.A(mai_mai_n488_), .B(mai_mai_n406_), .Y(mai_mai_n489_));
  INV        m461(.A(mai_mai_n207_), .Y(mai_mai_n490_));
  NO2        m462(.A(mai_mai_n490_), .B(mai_mai_n426_), .Y(mai_mai_n491_));
  NO3        m463(.A(mai_mai_n491_), .B(mai_mai_n489_), .C(mai_mai_n442_), .Y(mai_mai_n492_));
  NO2        m464(.A(h), .B(m), .Y(mai_mai_n493_));
  NA2        m465(.A(mai_mai_n82_), .B(mai_mai_n69_), .Y(mai_mai_n494_));
  NA2        m466(.A(n), .B(mai_mai_n146_), .Y(mai_mai_n495_));
  INV        m467(.A(mai_mai_n495_), .Y(mai_mai_n496_));
  NA3        m468(.A(mai_mai_n84_), .B(mai_mai_n56_), .C(m), .Y(mai_mai_n497_));
  NOi31      m469(.An(c), .B(h), .C(mai_mai_n497_), .Y(mai_mai_n498_));
  INV        m470(.A(mai_mai_n451_), .Y(mai_mai_n499_));
  NAi21      m471(.An(mai_mai_n428_), .B(mai_mai_n499_), .Y(mai_mai_n500_));
  NO3        m472(.A(mai_mai_n500_), .B(mai_mai_n498_), .C(mai_mai_n496_), .Y(mai_mai_n501_));
  AN2        m473(.A(mai_mai_n501_), .B(mai_mai_n494_), .Y(mai_mai_n502_));
  NA4        m474(.A(mai_mai_n265_), .B(k), .C(mai_mai_n96_), .D(h), .Y(mai_mai_n503_));
  AOI220     m475(.A0(mai_mai_n387_), .A1(d), .B0(mai_mai_n265_), .B1(mai_mai_n106_), .Y(mai_mai_n504_));
  NO3        m476(.A(mai_mai_n426_), .B(f), .C(mai_mai_n295_), .Y(mai_mai_n505_));
  INV        m477(.A(mai_mai_n61_), .Y(mai_mai_n506_));
  AN2        m478(.A(mai_mai_n506_), .B(mai_mai_n460_), .Y(mai_mai_n507_));
  NO2        m479(.A(mai_mai_n507_), .B(mai_mai_n505_), .Y(mai_mai_n508_));
  NA2        m480(.A(mai_mai_n508_), .B(mai_mai_n504_), .Y(mai_mai_n509_));
  NO2        m481(.A(mai_mai_n509_), .B(mai_mai_n574_), .Y(mai_mai_n510_));
  NA2        m482(.A(mai_mai_n341_), .B(mai_mai_n308_), .Y(mai_mai_n511_));
  NA4        m483(.A(mai_mai_n511_), .B(mai_mai_n510_), .C(mai_mai_n502_), .D(mai_mai_n492_), .Y(mai01));
  NA2        m484(.A(mai_mai_n390_), .B(c), .Y(mai_mai_n513_));
  NA2        m485(.A(mai_mai_n513_), .B(mai_mai_n374_), .Y(mai_mai_n514_));
  INV        m486(.A(mai_mai_n503_), .Y(mai_mai_n515_));
  INV        m487(.A(mai_mai_n515_), .Y(mai_mai_n516_));
  NAi31      m488(.An(mai_mai_n77_), .B(mai_mai_n240_), .C(mai_mai_n516_), .Y(mai_mai_n517_));
  NO2        m489(.A(mai_mai_n517_), .B(mai_mai_n514_), .Y(mai_mai_n518_));
  NA2        m490(.A(mai_mai_n328_), .B(m), .Y(mai_mai_n519_));
  INV        m491(.A(mai_mai_n519_), .Y(mai_mai_n520_));
  NO2        m492(.A(mai_mai_n580_), .B(mai_mai_n520_), .Y(mai_mai_n521_));
  NA2        m493(.A(mai_mai_n204_), .B(c), .Y(mai_mai_n522_));
  NO3        m494(.A(mai_mai_n458_), .B(mai_mai_n81_), .C(mai_mai_n47_), .Y(mai_mai_n523_));
  NO2        m495(.A(mai_mai_n458_), .B(mai_mai_n79_), .Y(mai_mai_n524_));
  NO3        m496(.A(mai_mai_n524_), .B(mai_mai_n523_), .C(mai_mai_n259_), .Y(mai_mai_n525_));
  NA4        m497(.A(mai_mai_n525_), .B(mai_mai_n522_), .C(mai_mai_n521_), .D(mai_mai_n518_), .Y(mai06));
  INV        m498(.A(mai_mai_n52_), .Y(mai_mai_n527_));
  OAI210     m499(.A0(mai_mai_n527_), .A1(mai_mai_n523_), .B0(c), .Y(mai_mai_n528_));
  NA2        m500(.A(mai_mai_n361_), .B(mai_mai_n528_), .Y(mai_mai_n529_));
  NO2        m501(.A(mai_mai_n529_), .B(mai_mai_n113_), .Y(mai_mai_n530_));
  AOI210     m502(.A0(i), .A1(mai_mai_n230_), .B0(mai_mai_n290_), .Y(mai_mai_n531_));
  NO2        m503(.A(mai_mai_n531_), .B(mai_mai_n142_), .Y(mai_mai_n532_));
  NA2        m504(.A(mai_mai_n37_), .B(mai_mai_n260_), .Y(mai_mai_n533_));
  INV        m505(.A(mai_mai_n533_), .Y(mai_mai_n534_));
  NO3        m506(.A(mai_mai_n387_), .B(mai_mai_n534_), .C(mai_mai_n532_), .Y(mai_mai_n535_));
  NO2        m507(.A(mai_mai_n99_), .B(mai_mai_n253_), .Y(mai_mai_n536_));
  NA2        m508(.A(a), .B(mai_mai_n536_), .Y(mai_mai_n537_));
  NA3        m509(.A(mai_mai_n208_), .B(mai_mai_n537_), .C(mai_mai_n504_), .Y(mai_mai_n538_));
  NO2        m510(.A(mai_mai_n354_), .B(mai_mai_n538_), .Y(mai_mai_n539_));
  NA4        m511(.A(mai_mai_n539_), .B(mai_mai_n535_), .C(mai_mai_n530_), .D(mai_mai_n525_), .Y(mai07));
  NOi31      m512(.An(n), .B(m), .C(b), .Y(mai_mai_n541_));
  NA3        m513(.A(mai_mai_n287_), .B(mai_mai_n280_), .C(mai_mai_n56_), .Y(mai_mai_n542_));
  NO2        m514(.A(mai_mai_n542_), .B(mai_mai_n36_), .Y(mai_mai_n543_));
  INV        m515(.A(mai_mai_n543_), .Y(mai_mai_n544_));
  NOi31      m516(.An(m), .B(n), .C(b), .Y(mai_mai_n545_));
  OAI210     m517(.A0(mai_mai_n85_), .A1(mai_mai_n213_), .B0(mai_mai_n436_), .Y(mai_mai_n546_));
  NO4        m518(.A(mai_mai_n61_), .B(m), .C(f), .D(e), .Y(mai_mai_n547_));
  NA2        m519(.A(mai_mai_n546_), .B(mai_mai_n544_), .Y(mai_mai_n548_));
  OR2        m520(.A(n), .B(i), .Y(mai_mai_n549_));
  OAI210     m521(.A0(mai_mai_n549_), .A1(mai_mai_n446_), .B0(mai_mai_n38_), .Y(mai_mai_n550_));
  NA2        m522(.A(mai_mai_n550_), .B(mai_mai_n493_), .Y(mai_mai_n551_));
  OAI210     m523(.A0(mai_mai_n547_), .A1(mai_mai_n541_), .B0(mai_mai_n358_), .Y(mai_mai_n552_));
  INV        m524(.A(mai_mai_n552_), .Y(mai_mai_n553_));
  NA2        m525(.A(mai_mai_n55_), .B(mai_mai_n545_), .Y(mai_mai_n554_));
  INV        m526(.A(mai_mai_n554_), .Y(mai_mai_n555_));
  NO2        m527(.A(mai_mai_n555_), .B(mai_mai_n553_), .Y(mai_mai_n556_));
  INV        m528(.A(mai_mai_n556_), .Y(mai_mai_n557_));
  OR3        m529(.A(mai_mai_n557_), .B(mai_mai_n577_), .C(mai_mai_n548_), .Y(mai04));
  NOi31      m530(.An(mai_mai_n547_), .B(k), .C(mai_mai_n426_), .Y(mai_mai_n559_));
  NO3        m531(.A(mai_mai_n116_), .B(mai_mai_n420_), .C(j), .Y(mai_mai_n560_));
  OR3        m532(.A(mai_mai_n560_), .B(mai_mai_n559_), .C(mai_mai_n438_), .Y(mai_mai_n561_));
  NO3        m533(.A(i), .B(mai_mai_n49_), .C(k), .Y(mai_mai_n562_));
  AOI210     m534(.A0(mai_mai_n562_), .A1(mai_mai_n434_), .B0(mai_mai_n498_), .Y(mai_mai_n563_));
  NA2        m535(.A(mai_mai_n563_), .B(mai_mai_n508_), .Y(mai_mai_n564_));
  NO4        m536(.A(mai_mai_n564_), .B(mai_mai_n561_), .C(mai_mai_n445_), .D(mai_mai_n430_), .Y(mai_mai_n565_));
  NA4        m537(.A(mai_mai_n565_), .B(mai_mai_n448_), .C(mai_mai_n474_), .D(mai_mai_n466_), .Y(mai05));
  INV        m538(.A(m), .Y(mai_mai_n569_));
  INV        m539(.A(b), .Y(mai_mai_n570_));
  INV        m540(.A(mai_mai_n287_), .Y(mai_mai_n571_));
  INV        m541(.A(m), .Y(mai_mai_n572_));
  INV        m542(.A(b), .Y(mai_mai_n573_));
  INV        m543(.A(mai_mai_n503_), .Y(mai_mai_n574_));
  INV        m544(.A(i), .Y(mai_mai_n575_));
  INV        m545(.A(m), .Y(mai_mai_n576_));
  INV        m546(.A(mai_mai_n551_), .Y(mai_mai_n577_));
  INV        m547(.A(mai_mai_n416_), .Y(mai_mai_n578_));
  INV        m548(.A(mai_mai_n283_), .Y(mai_mai_n579_));
  INV        m549(.A(mai_mai_n119_), .Y(mai_mai_n580_));
  INV        m550(.A(c), .Y(mai_mai_n581_));
  INV        m551(.A(mai_mai_n317_), .Y(mai_mai_n582_));
  INV        m552(.A(a), .Y(mai_mai_n583_));
  INV        m553(.A(b), .Y(mai_mai_n584_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA2        u0003(.A(men_men_n31_), .B(men_men_n30_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(u), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(u), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(u), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(u), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(u), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(u), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(u), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(u), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(u), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  INV        u0059(.A(men_men_n87_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(u), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(u), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(u), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n96_), .C(f), .Y(men_men_n98_));
  AN2        u0070(.A(j), .B(u), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(l), .C(i), .Y(men_men_n100_));
  NOi21      u0072(.An(u), .B(i), .Y(men_men_n101_));
  NOi32      u0073(.An(m), .Bn(j), .C(k), .Y(men_men_n102_));
  AOI220     u0074(.A0(men_men_n102_), .A1(men_men_n101_), .B0(men_men_n100_), .B1(men_men_n99_), .Y(men_men_n103_));
  NO2        u0075(.A(men_men_n103_), .B(f), .Y(men_men_n104_));
  NO4        u0076(.A(men_men_n104_), .B(men_men_n98_), .C(men_men_n95_), .D(men_men_n92_), .Y(men_men_n105_));
  NAi41      u0077(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n106_));
  AN2        u0078(.A(e), .B(b), .Y(men_men_n107_));
  NOi31      u0079(.An(c), .B(h), .C(f), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NO3        u0081(.A(men_men_n109_), .B(men_men_n106_), .C(u), .Y(men_men_n110_));
  NOi21      u0082(.An(u), .B(f), .Y(men_men_n111_));
  NOi21      u0083(.An(i), .B(h), .Y(men_men_n112_));
  NA3        u0084(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n36_), .Y(men_men_n113_));
  INV        u0085(.A(a), .Y(men_men_n114_));
  NA2        u0086(.A(men_men_n107_), .B(men_men_n114_), .Y(men_men_n115_));
  INV        u0087(.A(l), .Y(men_men_n116_));
  NOi21      u0088(.An(m), .B(n), .Y(men_men_n117_));
  AN2        u0089(.A(k), .B(h), .Y(men_men_n118_));
  NO2        u0090(.A(men_men_n113_), .B(men_men_n88_), .Y(men_men_n119_));
  INV        u0091(.A(b), .Y(men_men_n120_));
  NA2        u0092(.A(l), .B(j), .Y(men_men_n121_));
  AN2        u0093(.A(k), .B(i), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n121_), .Y(men_men_n123_));
  NA2        u0095(.A(u), .B(e), .Y(men_men_n124_));
  NOi32      u0096(.An(c), .Bn(a), .C(d), .Y(men_men_n125_));
  NA2        u0097(.A(men_men_n125_), .B(men_men_n117_), .Y(men_men_n126_));
  NO4        u0098(.A(men_men_n126_), .B(men_men_n124_), .C(men_men_n123_), .D(men_men_n120_), .Y(men_men_n127_));
  NO3        u0099(.A(men_men_n127_), .B(men_men_n119_), .C(men_men_n110_), .Y(men_men_n128_));
  OAI210     u0100(.A0(men_men_n105_), .A1(men_men_n88_), .B0(men_men_n128_), .Y(men_men_n129_));
  NOi31      u0101(.An(k), .B(m), .C(j), .Y(men_men_n130_));
  NA3        u0102(.A(men_men_n130_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n131_));
  NOi31      u0103(.An(k), .B(m), .C(i), .Y(men_men_n132_));
  NA3        u0104(.A(men_men_n132_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n133_));
  NA2        u0105(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n134_));
  NOi32      u0106(.An(f), .Bn(b), .C(e), .Y(men_men_n135_));
  NAi21      u0107(.An(u), .B(h), .Y(men_men_n136_));
  NAi21      u0108(.An(m), .B(n), .Y(men_men_n137_));
  NAi21      u0109(.An(j), .B(k), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n139_));
  NAi41      u0111(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n140_));
  NAi31      u0112(.An(j), .B(k), .C(h), .Y(men_men_n141_));
  NO3        u0113(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n137_), .Y(men_men_n142_));
  AOI210     u0114(.A0(men_men_n139_), .A1(men_men_n135_), .B0(men_men_n142_), .Y(men_men_n143_));
  NO2        u0115(.A(k), .B(j), .Y(men_men_n144_));
  NO2        u0116(.A(men_men_n144_), .B(men_men_n137_), .Y(men_men_n145_));
  AN2        u0117(.A(k), .B(j), .Y(men_men_n146_));
  NAi21      u0118(.An(c), .B(b), .Y(men_men_n147_));
  NA2        u0119(.A(f), .B(d), .Y(men_men_n148_));
  NO3        u0120(.A(men_men_n147_), .B(men_men_n146_), .C(men_men_n136_), .Y(men_men_n149_));
  NAi31      u0121(.An(f), .B(e), .C(b), .Y(men_men_n150_));
  NA2        u0122(.A(men_men_n149_), .B(men_men_n145_), .Y(men_men_n151_));
  NA2        u0123(.A(d), .B(b), .Y(men_men_n152_));
  NAi21      u0124(.An(e), .B(f), .Y(men_men_n153_));
  NO2        u0125(.A(men_men_n153_), .B(men_men_n152_), .Y(men_men_n154_));
  NA2        u0126(.A(b), .B(a), .Y(men_men_n155_));
  NAi21      u0127(.An(e), .B(u), .Y(men_men_n156_));
  NAi21      u0128(.An(c), .B(d), .Y(men_men_n157_));
  NAi31      u0129(.An(l), .B(k), .C(h), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n137_), .B(men_men_n158_), .Y(men_men_n159_));
  NA2        u0131(.A(men_men_n159_), .B(men_men_n154_), .Y(men_men_n160_));
  NAi41      u0132(.An(men_men_n134_), .B(men_men_n160_), .C(men_men_n151_), .D(men_men_n143_), .Y(men_men_n161_));
  NAi31      u0133(.An(e), .B(f), .C(b), .Y(men_men_n162_));
  NOi21      u0134(.An(u), .B(d), .Y(men_men_n163_));
  NO2        u0135(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  NOi21      u0136(.An(h), .B(i), .Y(men_men_n165_));
  NOi21      u0137(.An(k), .B(m), .Y(men_men_n166_));
  NA3        u0138(.A(men_men_n166_), .B(men_men_n165_), .C(n), .Y(men_men_n167_));
  NOi21      u0139(.An(men_men_n164_), .B(men_men_n167_), .Y(men_men_n168_));
  NOi21      u0140(.An(h), .B(u), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  NAi31      u0143(.An(l), .B(j), .C(h), .Y(men_men_n172_));
  NO2        u0144(.A(men_men_n172_), .B(men_men_n49_), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n67_), .Y(men_men_n174_));
  NOi32      u0146(.An(n), .Bn(k), .C(m), .Y(men_men_n175_));
  NA2        u0147(.A(l), .B(i), .Y(men_men_n176_));
  NA2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  OAI210     u0149(.A0(men_men_n177_), .A1(men_men_n171_), .B0(men_men_n174_), .Y(men_men_n178_));
  NAi31      u0150(.An(d), .B(f), .C(c), .Y(men_men_n179_));
  NAi31      u0151(.An(e), .B(f), .C(c), .Y(men_men_n180_));
  NA2        u0152(.A(men_men_n180_), .B(men_men_n179_), .Y(men_men_n181_));
  NA2        u0153(.A(j), .B(h), .Y(men_men_n182_));
  OR3        u0154(.A(n), .B(m), .C(k), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  NAi32      u0156(.An(m), .Bn(k), .C(n), .Y(men_men_n185_));
  NO2        u0157(.A(men_men_n185_), .B(men_men_n182_), .Y(men_men_n186_));
  AOI220     u0158(.A0(men_men_n186_), .A1(men_men_n164_), .B0(men_men_n184_), .B1(men_men_n181_), .Y(men_men_n187_));
  NO2        u0159(.A(n), .B(m), .Y(men_men_n188_));
  NA2        u0160(.A(men_men_n188_), .B(men_men_n50_), .Y(men_men_n189_));
  NAi21      u0161(.An(f), .B(e), .Y(men_men_n190_));
  NA2        u0162(.A(d), .B(c), .Y(men_men_n191_));
  NO2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NOi21      u0164(.An(men_men_n192_), .B(men_men_n189_), .Y(men_men_n193_));
  NAi21      u0165(.An(d), .B(c), .Y(men_men_n194_));
  NAi31      u0166(.An(m), .B(n), .C(b), .Y(men_men_n195_));
  NA2        u0167(.A(k), .B(i), .Y(men_men_n196_));
  NAi21      u0168(.An(h), .B(f), .Y(men_men_n197_));
  INV        u0169(.A(men_men_n197_), .Y(men_men_n198_));
  NO2        u0170(.A(men_men_n195_), .B(men_men_n157_), .Y(men_men_n199_));
  NA2        u0171(.A(men_men_n199_), .B(men_men_n198_), .Y(men_men_n200_));
  NOi32      u0172(.An(f), .Bn(c), .C(d), .Y(men_men_n201_));
  NOi32      u0173(.An(f), .Bn(c), .C(e), .Y(men_men_n202_));
  NO2        u0174(.A(men_men_n202_), .B(men_men_n201_), .Y(men_men_n203_));
  NO3        u0175(.A(n), .B(m), .C(j), .Y(men_men_n204_));
  NA2        u0176(.A(men_men_n204_), .B(men_men_n118_), .Y(men_men_n205_));
  AO210      u0177(.A0(men_men_n205_), .A1(men_men_n189_), .B0(men_men_n203_), .Y(men_men_n206_));
  NAi41      u0178(.An(men_men_n193_), .B(men_men_n206_), .C(men_men_n200_), .D(men_men_n187_), .Y(men_men_n207_));
  OR4        u0179(.A(men_men_n207_), .B(men_men_n178_), .C(men_men_n168_), .D(men_men_n161_), .Y(men_men_n208_));
  NO4        u0180(.A(men_men_n208_), .B(men_men_n129_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n209_));
  NA3        u0181(.A(m), .B(men_men_n116_), .C(j), .Y(men_men_n210_));
  NAi31      u0182(.An(n), .B(h), .C(u), .Y(men_men_n211_));
  NO2        u0183(.A(men_men_n211_), .B(men_men_n210_), .Y(men_men_n212_));
  NOi32      u0184(.An(m), .Bn(k), .C(l), .Y(men_men_n213_));
  NA3        u0185(.A(men_men_n213_), .B(men_men_n89_), .C(u), .Y(men_men_n214_));
  NO2        u0186(.A(men_men_n214_), .B(n), .Y(men_men_n215_));
  NOi21      u0187(.An(k), .B(j), .Y(men_men_n216_));
  NA4        u0188(.A(men_men_n216_), .B(men_men_n117_), .C(i), .D(u), .Y(men_men_n217_));
  AN2        u0189(.A(i), .B(u), .Y(men_men_n218_));
  NA3        u0190(.A(men_men_n76_), .B(men_men_n218_), .C(men_men_n117_), .Y(men_men_n219_));
  NA2        u0191(.A(men_men_n219_), .B(men_men_n217_), .Y(men_men_n220_));
  NO3        u0192(.A(men_men_n220_), .B(men_men_n215_), .C(men_men_n212_), .Y(men_men_n221_));
  NAi41      u0193(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n222_));
  INV        u0194(.A(men_men_n222_), .Y(men_men_n223_));
  INV        u0195(.A(f), .Y(men_men_n224_));
  INV        u0196(.A(u), .Y(men_men_n225_));
  NOi31      u0197(.An(i), .B(j), .C(h), .Y(men_men_n226_));
  NOi21      u0198(.An(l), .B(m), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n228_));
  NO3        u0200(.A(men_men_n228_), .B(men_men_n225_), .C(men_men_n224_), .Y(men_men_n229_));
  NA2        u0201(.A(men_men_n229_), .B(men_men_n223_), .Y(men_men_n230_));
  OAI210     u0202(.A0(men_men_n221_), .A1(men_men_n32_), .B0(men_men_n230_), .Y(men_men_n231_));
  NOi21      u0203(.An(n), .B(m), .Y(men_men_n232_));
  NOi32      u0204(.An(l), .Bn(i), .C(j), .Y(men_men_n233_));
  NA2        u0205(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n234_));
  OA220      u0206(.A0(men_men_n234_), .A1(men_men_n109_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n235_));
  NAi21      u0207(.An(j), .B(h), .Y(men_men_n236_));
  XN2        u0208(.A(i), .B(h), .Y(men_men_n237_));
  NA2        u0209(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  NOi31      u0210(.An(k), .B(n), .C(m), .Y(men_men_n239_));
  NOi31      u0211(.An(men_men_n239_), .B(men_men_n191_), .C(men_men_n190_), .Y(men_men_n240_));
  NA2        u0212(.A(men_men_n240_), .B(men_men_n238_), .Y(men_men_n241_));
  NAi31      u0213(.An(f), .B(e), .C(c), .Y(men_men_n242_));
  NO4        u0214(.A(men_men_n242_), .B(men_men_n183_), .C(men_men_n182_), .D(men_men_n59_), .Y(men_men_n243_));
  NA4        u0215(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n244_));
  NAi32      u0216(.An(m), .Bn(i), .C(k), .Y(men_men_n245_));
  NO3        u0217(.A(men_men_n245_), .B(men_men_n93_), .C(men_men_n244_), .Y(men_men_n246_));
  NA2        u0218(.A(k), .B(h), .Y(men_men_n247_));
  NO2        u0219(.A(men_men_n246_), .B(men_men_n243_), .Y(men_men_n248_));
  NAi21      u0220(.An(n), .B(a), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(men_men_n152_), .Y(men_men_n250_));
  NAi41      u0222(.An(u), .B(m), .C(k), .D(h), .Y(men_men_n251_));
  NO2        u0223(.A(men_men_n251_), .B(e), .Y(men_men_n252_));
  NO3        u0224(.A(men_men_n153_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n253_));
  OAI210     u0225(.A0(men_men_n253_), .A1(men_men_n252_), .B0(men_men_n250_), .Y(men_men_n254_));
  AN4        u0226(.A(men_men_n254_), .B(men_men_n248_), .C(men_men_n241_), .D(men_men_n235_), .Y(men_men_n255_));
  OR2        u0227(.A(h), .B(u), .Y(men_men_n256_));
  NO2        u0228(.A(men_men_n256_), .B(men_men_n106_), .Y(men_men_n257_));
  NA2        u0229(.A(men_men_n257_), .B(men_men_n135_), .Y(men_men_n258_));
  NAi41      u0230(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n259_), .B(men_men_n224_), .Y(men_men_n260_));
  NA2        u0232(.A(men_men_n166_), .B(men_men_n112_), .Y(men_men_n261_));
  NAi21      u0233(.An(men_men_n261_), .B(men_men_n260_), .Y(men_men_n262_));
  NO2        u0234(.A(n), .B(a), .Y(men_men_n263_));
  NAi31      u0235(.An(men_men_n251_), .B(men_men_n263_), .C(men_men_n107_), .Y(men_men_n264_));
  AN2        u0236(.A(men_men_n264_), .B(men_men_n262_), .Y(men_men_n265_));
  NAi21      u0237(.An(h), .B(i), .Y(men_men_n266_));
  NA2        u0238(.A(men_men_n188_), .B(k), .Y(men_men_n267_));
  NO2        u0239(.A(men_men_n267_), .B(men_men_n266_), .Y(men_men_n268_));
  NA2        u0240(.A(men_men_n268_), .B(men_men_n201_), .Y(men_men_n269_));
  NA3        u0241(.A(men_men_n269_), .B(men_men_n265_), .C(men_men_n258_), .Y(men_men_n270_));
  NOi21      u0242(.An(u), .B(e), .Y(men_men_n271_));
  NO2        u0243(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n272_));
  NA2        u0244(.A(men_men_n272_), .B(men_men_n271_), .Y(men_men_n273_));
  NOi32      u0245(.An(l), .Bn(j), .C(i), .Y(men_men_n274_));
  AOI210     u0246(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n274_), .Y(men_men_n275_));
  NO2        u0247(.A(men_men_n266_), .B(men_men_n44_), .Y(men_men_n276_));
  NAi21      u0248(.An(f), .B(u), .Y(men_men_n277_));
  NO2        u0249(.A(men_men_n277_), .B(men_men_n65_), .Y(men_men_n278_));
  NO2        u0250(.A(men_men_n69_), .B(men_men_n121_), .Y(men_men_n279_));
  AOI220     u0251(.A0(men_men_n279_), .A1(men_men_n278_), .B0(men_men_n276_), .B1(men_men_n67_), .Y(men_men_n280_));
  OAI210     u0252(.A0(men_men_n275_), .A1(men_men_n273_), .B0(men_men_n280_), .Y(men_men_n281_));
  NO3        u0253(.A(men_men_n138_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n282_));
  NOi41      u0254(.An(men_men_n255_), .B(men_men_n281_), .C(men_men_n270_), .D(men_men_n231_), .Y(men_men_n283_));
  NO4        u0255(.A(men_men_n212_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n284_));
  NO2        u0256(.A(men_men_n284_), .B(men_men_n115_), .Y(men_men_n285_));
  NA3        u0257(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n286_));
  NAi21      u0258(.An(h), .B(u), .Y(men_men_n287_));
  OR4        u0259(.A(men_men_n287_), .B(men_men_n286_), .C(men_men_n234_), .D(e), .Y(men_men_n288_));
  NO2        u0260(.A(men_men_n261_), .B(men_men_n277_), .Y(men_men_n289_));
  NA2        u0261(.A(men_men_n289_), .B(men_men_n78_), .Y(men_men_n290_));
  NAi31      u0262(.An(u), .B(k), .C(h), .Y(men_men_n291_));
  NO3        u0263(.A(men_men_n137_), .B(men_men_n291_), .C(l), .Y(men_men_n292_));
  NAi31      u0264(.An(e), .B(d), .C(a), .Y(men_men_n293_));
  NA2        u0265(.A(men_men_n292_), .B(men_men_n135_), .Y(men_men_n294_));
  NA3        u0266(.A(men_men_n294_), .B(men_men_n290_), .C(men_men_n288_), .Y(men_men_n295_));
  NA4        u0267(.A(men_men_n166_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n121_), .Y(men_men_n296_));
  NA3        u0268(.A(men_men_n166_), .B(men_men_n165_), .C(men_men_n86_), .Y(men_men_n297_));
  NO2        u0269(.A(men_men_n297_), .B(men_men_n203_), .Y(men_men_n298_));
  NOi21      u0270(.An(men_men_n296_), .B(men_men_n298_), .Y(men_men_n299_));
  NA3        u0271(.A(e), .B(c), .C(b), .Y(men_men_n300_));
  NO2        u0272(.A(men_men_n60_), .B(men_men_n300_), .Y(men_men_n301_));
  NAi32      u0273(.An(k), .Bn(i), .C(j), .Y(men_men_n302_));
  NAi31      u0274(.An(h), .B(l), .C(i), .Y(men_men_n303_));
  NA3        u0275(.A(men_men_n303_), .B(men_men_n302_), .C(men_men_n172_), .Y(men_men_n304_));
  NOi21      u0276(.An(men_men_n304_), .B(men_men_n49_), .Y(men_men_n305_));
  OAI210     u0277(.A0(men_men_n278_), .A1(men_men_n301_), .B0(men_men_n305_), .Y(men_men_n306_));
  NAi21      u0278(.An(l), .B(k), .Y(men_men_n307_));
  NO2        u0279(.A(men_men_n307_), .B(men_men_n49_), .Y(men_men_n308_));
  NOi21      u0280(.An(l), .B(j), .Y(men_men_n309_));
  NA2        u0281(.A(men_men_n169_), .B(men_men_n309_), .Y(men_men_n310_));
  NA3        u0282(.A(men_men_n122_), .B(men_men_n121_), .C(u), .Y(men_men_n311_));
  OR3        u0283(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n312_));
  AOI210     u0284(.A0(men_men_n311_), .A1(men_men_n310_), .B0(men_men_n312_), .Y(men_men_n313_));
  INV        u0285(.A(men_men_n313_), .Y(men_men_n314_));
  NAi32      u0286(.An(j), .Bn(h), .C(i), .Y(men_men_n315_));
  NAi21      u0287(.An(m), .B(l), .Y(men_men_n316_));
  NO3        u0288(.A(men_men_n316_), .B(men_men_n315_), .C(men_men_n86_), .Y(men_men_n317_));
  NA2        u0289(.A(h), .B(u), .Y(men_men_n318_));
  NA2        u0290(.A(men_men_n175_), .B(men_men_n45_), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n319_), .B(men_men_n318_), .Y(men_men_n320_));
  NA2        u0292(.A(men_men_n320_), .B(men_men_n170_), .Y(men_men_n321_));
  NA4        u0293(.A(men_men_n321_), .B(men_men_n314_), .C(men_men_n306_), .D(men_men_n299_), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n150_), .B(d), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n323_), .B(men_men_n53_), .Y(men_men_n324_));
  NO2        u0296(.A(men_men_n109_), .B(men_men_n106_), .Y(men_men_n325_));
  NAi32      u0297(.An(n), .Bn(m), .C(l), .Y(men_men_n326_));
  NO2        u0298(.A(men_men_n326_), .B(men_men_n315_), .Y(men_men_n327_));
  NA2        u0299(.A(men_men_n327_), .B(men_men_n192_), .Y(men_men_n328_));
  NO2        u0300(.A(men_men_n126_), .B(men_men_n120_), .Y(men_men_n329_));
  NAi31      u0301(.An(k), .B(l), .C(j), .Y(men_men_n330_));
  OAI210     u0302(.A0(men_men_n307_), .A1(j), .B0(men_men_n330_), .Y(men_men_n331_));
  NOi21      u0303(.An(men_men_n331_), .B(men_men_n124_), .Y(men_men_n332_));
  NA2        u0304(.A(men_men_n332_), .B(men_men_n329_), .Y(men_men_n333_));
  NA3        u0305(.A(men_men_n333_), .B(men_men_n328_), .C(men_men_n324_), .Y(men_men_n334_));
  NO4        u0306(.A(men_men_n334_), .B(men_men_n322_), .C(men_men_n295_), .D(men_men_n285_), .Y(men_men_n335_));
  NA2        u0307(.A(men_men_n268_), .B(men_men_n202_), .Y(men_men_n336_));
  NAi21      u0308(.An(m), .B(k), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n237_), .B(men_men_n337_), .Y(men_men_n338_));
  NAi41      u0310(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n339_), .B(men_men_n156_), .Y(men_men_n340_));
  NA2        u0312(.A(men_men_n340_), .B(men_men_n338_), .Y(men_men_n341_));
  NAi31      u0313(.An(i), .B(l), .C(h), .Y(men_men_n342_));
  NO4        u0314(.A(men_men_n342_), .B(men_men_n156_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n343_));
  NA2        u0315(.A(e), .B(c), .Y(men_men_n344_));
  NO3        u0316(.A(men_men_n344_), .B(n), .C(d), .Y(men_men_n345_));
  NOi21      u0317(.An(f), .B(h), .Y(men_men_n346_));
  NA2        u0318(.A(men_men_n346_), .B(men_men_n122_), .Y(men_men_n347_));
  NO2        u0319(.A(men_men_n347_), .B(men_men_n225_), .Y(men_men_n348_));
  NAi31      u0320(.An(d), .B(e), .C(b), .Y(men_men_n349_));
  NO2        u0321(.A(men_men_n137_), .B(men_men_n349_), .Y(men_men_n350_));
  NA2        u0322(.A(men_men_n350_), .B(men_men_n348_), .Y(men_men_n351_));
  NAi41      u0323(.An(men_men_n343_), .B(men_men_n351_), .C(men_men_n341_), .D(men_men_n336_), .Y(men_men_n352_));
  NO4        u0324(.A(men_men_n339_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n225_), .Y(men_men_n353_));
  NA2        u0325(.A(men_men_n263_), .B(men_men_n107_), .Y(men_men_n354_));
  OR2        u0326(.A(men_men_n354_), .B(men_men_n214_), .Y(men_men_n355_));
  NOi31      u0327(.An(l), .B(n), .C(m), .Y(men_men_n356_));
  NA2        u0328(.A(men_men_n356_), .B(men_men_n226_), .Y(men_men_n357_));
  NO2        u0329(.A(men_men_n357_), .B(men_men_n203_), .Y(men_men_n358_));
  NAi32      u0330(.An(men_men_n358_), .Bn(men_men_n353_), .C(men_men_n355_), .Y(men_men_n359_));
  NAi32      u0331(.An(m), .Bn(j), .C(k), .Y(men_men_n360_));
  NAi41      u0332(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n361_));
  OAI210     u0333(.A0(men_men_n222_), .A1(men_men_n360_), .B0(men_men_n361_), .Y(men_men_n362_));
  NOi31      u0334(.An(j), .B(m), .C(k), .Y(men_men_n363_));
  NO2        u0335(.A(men_men_n130_), .B(men_men_n363_), .Y(men_men_n364_));
  AN3        u0336(.A(h), .B(u), .C(f), .Y(men_men_n365_));
  NAi31      u0337(.An(men_men_n364_), .B(men_men_n365_), .C(men_men_n362_), .Y(men_men_n366_));
  NOi32      u0338(.An(m), .Bn(j), .C(l), .Y(men_men_n367_));
  NO2        u0339(.A(men_men_n367_), .B(men_men_n100_), .Y(men_men_n368_));
  NAi32      u0340(.An(men_men_n368_), .Bn(men_men_n211_), .C(men_men_n323_), .Y(men_men_n369_));
  NO2        u0341(.A(men_men_n316_), .B(men_men_n315_), .Y(men_men_n370_));
  NO2        u0342(.A(men_men_n228_), .B(u), .Y(men_men_n371_));
  NO2        u0343(.A(men_men_n162_), .B(men_men_n86_), .Y(men_men_n372_));
  AOI220     u0344(.A0(men_men_n372_), .A1(men_men_n371_), .B0(men_men_n260_), .B1(men_men_n370_), .Y(men_men_n373_));
  NA2        u0345(.A(men_men_n245_), .B(men_men_n81_), .Y(men_men_n374_));
  NA3        u0346(.A(men_men_n374_), .B(men_men_n365_), .C(men_men_n223_), .Y(men_men_n375_));
  NA4        u0347(.A(men_men_n375_), .B(men_men_n373_), .C(men_men_n369_), .D(men_men_n366_), .Y(men_men_n376_));
  NA3        u0348(.A(h), .B(u), .C(f), .Y(men_men_n377_));
  NO2        u0349(.A(men_men_n377_), .B(men_men_n77_), .Y(men_men_n378_));
  NA2        u0350(.A(men_men_n361_), .B(men_men_n222_), .Y(men_men_n379_));
  NA2        u0351(.A(men_men_n169_), .B(e), .Y(men_men_n380_));
  NO2        u0352(.A(men_men_n380_), .B(men_men_n41_), .Y(men_men_n381_));
  AOI220     u0353(.A0(men_men_n381_), .A1(men_men_n329_), .B0(men_men_n379_), .B1(men_men_n378_), .Y(men_men_n382_));
  NOi32      u0354(.An(j), .Bn(u), .C(i), .Y(men_men_n383_));
  NA3        u0355(.A(men_men_n383_), .B(men_men_n307_), .C(men_men_n117_), .Y(men_men_n384_));
  AO210      u0356(.A0(men_men_n115_), .A1(men_men_n32_), .B0(men_men_n384_), .Y(men_men_n385_));
  NOi32      u0357(.An(e), .Bn(b), .C(a), .Y(men_men_n386_));
  AN2        u0358(.A(l), .B(j), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n337_), .B(men_men_n387_), .Y(men_men_n388_));
  NO3        u0360(.A(men_men_n339_), .B(men_men_n72_), .C(men_men_n225_), .Y(men_men_n389_));
  NA3        u0361(.A(men_men_n219_), .B(men_men_n217_), .C(men_men_n35_), .Y(men_men_n390_));
  AOI220     u0362(.A0(men_men_n390_), .A1(men_men_n386_), .B0(men_men_n389_), .B1(men_men_n388_), .Y(men_men_n391_));
  NO2        u0363(.A(men_men_n349_), .B(n), .Y(men_men_n392_));
  NA2        u0364(.A(men_men_n218_), .B(k), .Y(men_men_n393_));
  NA3        u0365(.A(m), .B(men_men_n116_), .C(men_men_n224_), .Y(men_men_n394_));
  NA4        u0366(.A(men_men_n213_), .B(men_men_n89_), .C(u), .D(men_men_n224_), .Y(men_men_n395_));
  OAI210     u0367(.A0(men_men_n394_), .A1(men_men_n393_), .B0(men_men_n395_), .Y(men_men_n396_));
  NAi41      u0368(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n397_));
  NA2        u0369(.A(men_men_n51_), .B(men_men_n117_), .Y(men_men_n398_));
  NO2        u0370(.A(men_men_n398_), .B(men_men_n397_), .Y(men_men_n399_));
  AOI220     u0371(.A0(men_men_n399_), .A1(b), .B0(men_men_n396_), .B1(men_men_n392_), .Y(men_men_n400_));
  NA4        u0372(.A(men_men_n400_), .B(men_men_n391_), .C(men_men_n385_), .D(men_men_n382_), .Y(men_men_n401_));
  NO4        u0373(.A(men_men_n401_), .B(men_men_n376_), .C(men_men_n359_), .D(men_men_n352_), .Y(men_men_n402_));
  NA4        u0374(.A(men_men_n402_), .B(men_men_n335_), .C(men_men_n283_), .D(men_men_n209_), .Y(men10));
  NA3        u0375(.A(m), .B(k), .C(i), .Y(men_men_n404_));
  NO3        u0376(.A(men_men_n404_), .B(j), .C(men_men_n225_), .Y(men_men_n405_));
  NOi21      u0377(.An(e), .B(f), .Y(men_men_n406_));
  NO4        u0378(.A(men_men_n157_), .B(men_men_n406_), .C(n), .D(men_men_n114_), .Y(men_men_n407_));
  NAi31      u0379(.An(b), .B(f), .C(c), .Y(men_men_n408_));
  INV        u0380(.A(men_men_n408_), .Y(men_men_n409_));
  NOi32      u0381(.An(k), .Bn(h), .C(j), .Y(men_men_n410_));
  NA2        u0382(.A(men_men_n410_), .B(men_men_n232_), .Y(men_men_n411_));
  NA2        u0383(.A(men_men_n167_), .B(men_men_n411_), .Y(men_men_n412_));
  AOI220     u0384(.A0(men_men_n412_), .A1(men_men_n409_), .B0(men_men_n407_), .B1(men_men_n405_), .Y(men_men_n413_));
  AN2        u0385(.A(j), .B(h), .Y(men_men_n414_));
  NO3        u0386(.A(n), .B(m), .C(k), .Y(men_men_n415_));
  NA2        u0387(.A(men_men_n415_), .B(men_men_n414_), .Y(men_men_n416_));
  NO3        u0388(.A(men_men_n416_), .B(men_men_n157_), .C(men_men_n224_), .Y(men_men_n417_));
  OR2        u0389(.A(m), .B(k), .Y(men_men_n418_));
  NO2        u0390(.A(men_men_n182_), .B(men_men_n418_), .Y(men_men_n419_));
  NA4        u0391(.A(n), .B(f), .C(c), .D(men_men_n120_), .Y(men_men_n420_));
  NOi21      u0392(.An(men_men_n419_), .B(men_men_n420_), .Y(men_men_n421_));
  NOi32      u0393(.An(d), .Bn(a), .C(c), .Y(men_men_n422_));
  NA2        u0394(.A(men_men_n422_), .B(men_men_n190_), .Y(men_men_n423_));
  NAi21      u0395(.An(i), .B(u), .Y(men_men_n424_));
  NAi31      u0396(.An(k), .B(m), .C(j), .Y(men_men_n425_));
  NO3        u0397(.A(men_men_n425_), .B(men_men_n424_), .C(n), .Y(men_men_n426_));
  NOi21      u0398(.An(men_men_n426_), .B(men_men_n423_), .Y(men_men_n427_));
  NO3        u0399(.A(men_men_n427_), .B(men_men_n421_), .C(men_men_n417_), .Y(men_men_n428_));
  NO2        u0400(.A(men_men_n420_), .B(men_men_n316_), .Y(men_men_n429_));
  NOi32      u0401(.An(f), .Bn(d), .C(c), .Y(men_men_n430_));
  AOI220     u0402(.A0(men_men_n430_), .A1(men_men_n327_), .B0(men_men_n429_), .B1(men_men_n226_), .Y(men_men_n431_));
  NA3        u0403(.A(men_men_n431_), .B(men_men_n428_), .C(men_men_n413_), .Y(men_men_n432_));
  NO2        u0404(.A(men_men_n59_), .B(men_men_n120_), .Y(men_men_n433_));
  NA2        u0405(.A(men_men_n263_), .B(men_men_n433_), .Y(men_men_n434_));
  INV        u0406(.A(e), .Y(men_men_n435_));
  NA2        u0407(.A(men_men_n46_), .B(e), .Y(men_men_n436_));
  OAI220     u0408(.A0(men_men_n436_), .A1(men_men_n210_), .B0(men_men_n214_), .B1(men_men_n435_), .Y(men_men_n437_));
  AN2        u0409(.A(u), .B(e), .Y(men_men_n438_));
  NA3        u0410(.A(men_men_n438_), .B(men_men_n213_), .C(i), .Y(men_men_n439_));
  OAI210     u0411(.A0(men_men_n91_), .A1(men_men_n435_), .B0(men_men_n439_), .Y(men_men_n440_));
  NO2        u0412(.A(men_men_n103_), .B(men_men_n435_), .Y(men_men_n441_));
  NO3        u0413(.A(men_men_n441_), .B(men_men_n440_), .C(men_men_n437_), .Y(men_men_n442_));
  NOi32      u0414(.An(h), .Bn(e), .C(u), .Y(men_men_n443_));
  NA3        u0415(.A(men_men_n443_), .B(men_men_n309_), .C(m), .Y(men_men_n444_));
  NOi21      u0416(.An(u), .B(h), .Y(men_men_n445_));
  AN3        u0417(.A(m), .B(l), .C(i), .Y(men_men_n446_));
  NA3        u0418(.A(men_men_n446_), .B(men_men_n445_), .C(e), .Y(men_men_n447_));
  AN3        u0419(.A(h), .B(u), .C(e), .Y(men_men_n448_));
  NA2        u0420(.A(men_men_n448_), .B(men_men_n100_), .Y(men_men_n449_));
  AN3        u0421(.A(men_men_n449_), .B(men_men_n447_), .C(men_men_n444_), .Y(men_men_n450_));
  AOI210     u0422(.A0(men_men_n450_), .A1(men_men_n442_), .B0(men_men_n434_), .Y(men_men_n451_));
  NA3        u0423(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n452_));
  NO2        u0424(.A(men_men_n452_), .B(men_men_n434_), .Y(men_men_n453_));
  NA3        u0425(.A(men_men_n422_), .B(men_men_n190_), .C(men_men_n86_), .Y(men_men_n454_));
  NAi31      u0426(.An(b), .B(c), .C(a), .Y(men_men_n455_));
  NO2        u0427(.A(men_men_n455_), .B(n), .Y(men_men_n456_));
  OAI210     u0428(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n457_));
  NO2        u0429(.A(men_men_n457_), .B(men_men_n153_), .Y(men_men_n458_));
  NA2        u0430(.A(men_men_n458_), .B(men_men_n456_), .Y(men_men_n459_));
  INV        u0431(.A(men_men_n459_), .Y(men_men_n460_));
  NO4        u0432(.A(men_men_n460_), .B(men_men_n453_), .C(men_men_n451_), .D(men_men_n432_), .Y(men_men_n461_));
  NA2        u0433(.A(i), .B(u), .Y(men_men_n462_));
  NO3        u0434(.A(men_men_n293_), .B(men_men_n462_), .C(c), .Y(men_men_n463_));
  NOi21      u0435(.An(d), .B(c), .Y(men_men_n464_));
  NA2        u0436(.A(men_men_n464_), .B(a), .Y(men_men_n465_));
  NA3        u0437(.A(i), .B(u), .C(f), .Y(men_men_n466_));
  OR2        u0438(.A(men_men_n466_), .B(men_men_n71_), .Y(men_men_n467_));
  NA3        u0439(.A(men_men_n446_), .B(men_men_n445_), .C(men_men_n190_), .Y(men_men_n468_));
  AOI210     u0440(.A0(men_men_n468_), .A1(men_men_n467_), .B0(men_men_n465_), .Y(men_men_n469_));
  AOI210     u0441(.A0(men_men_n463_), .A1(men_men_n308_), .B0(men_men_n469_), .Y(men_men_n470_));
  OR2        u0442(.A(n), .B(m), .Y(men_men_n471_));
  NO2        u0443(.A(men_men_n471_), .B(men_men_n158_), .Y(men_men_n472_));
  NO2        u0444(.A(men_men_n191_), .B(men_men_n153_), .Y(men_men_n473_));
  OAI210     u0445(.A0(men_men_n472_), .A1(men_men_n184_), .B0(men_men_n473_), .Y(men_men_n474_));
  INV        u0446(.A(men_men_n398_), .Y(men_men_n475_));
  NA3        u0447(.A(men_men_n475_), .B(men_men_n386_), .C(d), .Y(men_men_n476_));
  NO2        u0448(.A(men_men_n455_), .B(men_men_n49_), .Y(men_men_n477_));
  NO3        u0449(.A(men_men_n66_), .B(men_men_n116_), .C(e), .Y(men_men_n478_));
  NAi21      u0450(.An(k), .B(j), .Y(men_men_n479_));
  NA2        u0451(.A(men_men_n266_), .B(men_men_n479_), .Y(men_men_n480_));
  NA3        u0452(.A(men_men_n480_), .B(men_men_n478_), .C(men_men_n477_), .Y(men_men_n481_));
  NAi21      u0453(.An(e), .B(d), .Y(men_men_n482_));
  NO2        u0454(.A(men_men_n267_), .B(men_men_n224_), .Y(men_men_n483_));
  NA3        u0455(.A(men_men_n483_), .B(men_men_n1667_), .C(men_men_n238_), .Y(men_men_n484_));
  NA4        u0456(.A(men_men_n484_), .B(men_men_n481_), .C(men_men_n476_), .D(men_men_n474_), .Y(men_men_n485_));
  NO2        u0457(.A(men_men_n357_), .B(men_men_n224_), .Y(men_men_n486_));
  NA2        u0458(.A(men_men_n486_), .B(men_men_n1667_), .Y(men_men_n487_));
  NOi31      u0459(.An(n), .B(m), .C(k), .Y(men_men_n488_));
  AOI220     u0460(.A0(men_men_n488_), .A1(men_men_n414_), .B0(men_men_n232_), .B1(men_men_n50_), .Y(men_men_n489_));
  NAi31      u0461(.An(u), .B(f), .C(c), .Y(men_men_n490_));
  OR3        u0462(.A(men_men_n490_), .B(men_men_n489_), .C(e), .Y(men_men_n491_));
  NA3        u0463(.A(men_men_n491_), .B(men_men_n487_), .C(men_men_n328_), .Y(men_men_n492_));
  NOi41      u0464(.An(men_men_n470_), .B(men_men_n492_), .C(men_men_n485_), .D(men_men_n281_), .Y(men_men_n493_));
  NOi32      u0465(.An(c), .Bn(a), .C(b), .Y(men_men_n494_));
  NA2        u0466(.A(men_men_n494_), .B(men_men_n117_), .Y(men_men_n495_));
  INV        u0467(.A(men_men_n291_), .Y(men_men_n496_));
  AN2        u0468(.A(e), .B(d), .Y(men_men_n497_));
  NA2        u0469(.A(men_men_n497_), .B(men_men_n496_), .Y(men_men_n498_));
  INV        u0470(.A(men_men_n153_), .Y(men_men_n499_));
  NO2        u0471(.A(men_men_n136_), .B(men_men_n41_), .Y(men_men_n500_));
  NO2        u0472(.A(men_men_n66_), .B(e), .Y(men_men_n501_));
  NOi31      u0473(.An(j), .B(k), .C(i), .Y(men_men_n502_));
  NOi21      u0474(.An(men_men_n172_), .B(men_men_n502_), .Y(men_men_n503_));
  NA4        u0475(.A(men_men_n342_), .B(men_men_n503_), .C(men_men_n275_), .D(men_men_n123_), .Y(men_men_n504_));
  AOI220     u0476(.A0(men_men_n504_), .A1(men_men_n501_), .B0(men_men_n500_), .B1(men_men_n499_), .Y(men_men_n505_));
  AOI210     u0477(.A0(men_men_n505_), .A1(men_men_n498_), .B0(men_men_n495_), .Y(men_men_n506_));
  NO2        u0478(.A(men_men_n220_), .B(men_men_n215_), .Y(men_men_n507_));
  NOi21      u0479(.An(a), .B(b), .Y(men_men_n508_));
  NA3        u0480(.A(e), .B(d), .C(c), .Y(men_men_n509_));
  NAi21      u0481(.An(men_men_n509_), .B(men_men_n508_), .Y(men_men_n510_));
  NO2        u0482(.A(men_men_n454_), .B(men_men_n214_), .Y(men_men_n511_));
  NOi21      u0483(.An(men_men_n510_), .B(men_men_n511_), .Y(men_men_n512_));
  AOI210     u0484(.A0(men_men_n284_), .A1(men_men_n507_), .B0(men_men_n512_), .Y(men_men_n513_));
  NO4        u0485(.A(men_men_n197_), .B(men_men_n106_), .C(men_men_n56_), .D(b), .Y(men_men_n514_));
  NA2        u0486(.A(men_men_n409_), .B(men_men_n159_), .Y(men_men_n515_));
  OR2        u0487(.A(k), .B(j), .Y(men_men_n516_));
  NA2        u0488(.A(l), .B(k), .Y(men_men_n517_));
  NA3        u0489(.A(men_men_n517_), .B(men_men_n516_), .C(men_men_n232_), .Y(men_men_n518_));
  AOI210     u0490(.A0(men_men_n245_), .A1(men_men_n360_), .B0(men_men_n86_), .Y(men_men_n519_));
  NOi21      u0491(.An(men_men_n518_), .B(men_men_n519_), .Y(men_men_n520_));
  NA3        u0492(.A(men_men_n296_), .B(men_men_n133_), .C(men_men_n131_), .Y(men_men_n521_));
  NA2        u0493(.A(men_men_n422_), .B(men_men_n117_), .Y(men_men_n522_));
  NO4        u0494(.A(men_men_n522_), .B(men_men_n97_), .C(men_men_n116_), .D(e), .Y(men_men_n523_));
  NO3        u0495(.A(men_men_n454_), .B(men_men_n94_), .C(men_men_n136_), .Y(men_men_n524_));
  NO4        u0496(.A(men_men_n524_), .B(men_men_n523_), .C(men_men_n521_), .D(men_men_n343_), .Y(men_men_n525_));
  NA2        u0497(.A(men_men_n525_), .B(men_men_n515_), .Y(men_men_n526_));
  NO4        u0498(.A(men_men_n526_), .B(men_men_n514_), .C(men_men_n513_), .D(men_men_n506_), .Y(men_men_n527_));
  NA2        u0499(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n528_));
  NOi21      u0500(.An(d), .B(e), .Y(men_men_n529_));
  NAi31      u0501(.An(j), .B(l), .C(i), .Y(men_men_n530_));
  OAI210     u0502(.A0(men_men_n530_), .A1(men_men_n137_), .B0(men_men_n106_), .Y(men_men_n531_));
  NO3        u0503(.A(men_men_n423_), .B(men_men_n368_), .C(men_men_n211_), .Y(men_men_n532_));
  NO2        u0504(.A(men_men_n423_), .B(men_men_n398_), .Y(men_men_n533_));
  NO4        u0505(.A(men_men_n533_), .B(men_men_n532_), .C(men_men_n193_), .D(men_men_n325_), .Y(men_men_n534_));
  NA3        u0506(.A(men_men_n534_), .B(men_men_n528_), .C(men_men_n255_), .Y(men_men_n535_));
  OAI210     u0507(.A0(men_men_n132_), .A1(men_men_n130_), .B0(n), .Y(men_men_n536_));
  NO2        u0508(.A(men_men_n536_), .B(men_men_n136_), .Y(men_men_n537_));
  OR2        u0509(.A(men_men_n317_), .B(men_men_n257_), .Y(men_men_n538_));
  OA210      u0510(.A0(men_men_n538_), .A1(men_men_n537_), .B0(men_men_n202_), .Y(men_men_n539_));
  XO2        u0511(.A(i), .B(h), .Y(men_men_n540_));
  NA3        u0512(.A(men_men_n540_), .B(men_men_n166_), .C(n), .Y(men_men_n541_));
  NAi41      u0513(.An(men_men_n317_), .B(men_men_n541_), .C(men_men_n489_), .D(men_men_n411_), .Y(men_men_n542_));
  AN2        u0514(.A(men_men_n542_), .B(men_men_n501_), .Y(men_men_n543_));
  NAi31      u0515(.An(c), .B(f), .C(d), .Y(men_men_n544_));
  AOI210     u0516(.A0(men_men_n297_), .A1(men_men_n205_), .B0(men_men_n544_), .Y(men_men_n545_));
  NOi21      u0517(.An(men_men_n84_), .B(men_men_n545_), .Y(men_men_n546_));
  NA3        u0518(.A(men_men_n407_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n547_));
  NA2        u0519(.A(men_men_n239_), .B(men_men_n112_), .Y(men_men_n548_));
  AOI210     u0520(.A0(men_men_n548_), .A1(men_men_n189_), .B0(men_men_n544_), .Y(men_men_n549_));
  AOI210     u0521(.A0(men_men_n384_), .A1(men_men_n35_), .B0(men_men_n510_), .Y(men_men_n550_));
  NOi31      u0522(.An(men_men_n547_), .B(men_men_n550_), .C(men_men_n549_), .Y(men_men_n551_));
  AO220      u0523(.A0(men_men_n305_), .A1(men_men_n278_), .B0(men_men_n173_), .B1(men_men_n67_), .Y(men_men_n552_));
  NA3        u0524(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n553_));
  NO2        u0525(.A(men_men_n553_), .B(men_men_n465_), .Y(men_men_n554_));
  NO2        u0526(.A(men_men_n554_), .B(men_men_n313_), .Y(men_men_n555_));
  NAi41      u0527(.An(men_men_n552_), .B(men_men_n555_), .C(men_men_n551_), .D(men_men_n546_), .Y(men_men_n556_));
  NO4        u0528(.A(men_men_n556_), .B(men_men_n543_), .C(men_men_n539_), .D(men_men_n535_), .Y(men_men_n557_));
  NA4        u0529(.A(men_men_n557_), .B(men_men_n527_), .C(men_men_n493_), .D(men_men_n461_), .Y(men11));
  NO2        u0530(.A(men_men_n73_), .B(f), .Y(men_men_n559_));
  NA2        u0531(.A(j), .B(u), .Y(men_men_n560_));
  NAi31      u0532(.An(i), .B(m), .C(l), .Y(men_men_n561_));
  NA3        u0533(.A(m), .B(k), .C(j), .Y(men_men_n562_));
  OAI220     u0534(.A0(men_men_n562_), .A1(men_men_n136_), .B0(men_men_n561_), .B1(men_men_n560_), .Y(men_men_n563_));
  NA2        u0535(.A(men_men_n563_), .B(men_men_n559_), .Y(men_men_n564_));
  NOi32      u0536(.An(e), .Bn(b), .C(f), .Y(men_men_n565_));
  NA2        u0537(.A(men_men_n274_), .B(men_men_n117_), .Y(men_men_n566_));
  NA2        u0538(.A(men_men_n46_), .B(j), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n567_), .B(men_men_n319_), .Y(men_men_n568_));
  NAi31      u0540(.An(d), .B(e), .C(a), .Y(men_men_n569_));
  NO2        u0541(.A(men_men_n569_), .B(n), .Y(men_men_n570_));
  AOI220     u0542(.A0(men_men_n570_), .A1(men_men_n104_), .B0(men_men_n568_), .B1(men_men_n565_), .Y(men_men_n571_));
  NAi41      u0543(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n572_));
  AN2        u0544(.A(men_men_n572_), .B(men_men_n397_), .Y(men_men_n573_));
  AOI210     u0545(.A0(men_men_n573_), .A1(men_men_n423_), .B0(men_men_n287_), .Y(men_men_n574_));
  NA2        u0546(.A(j), .B(i), .Y(men_men_n575_));
  NAi31      u0547(.An(n), .B(m), .C(k), .Y(men_men_n576_));
  NO3        u0548(.A(men_men_n576_), .B(men_men_n575_), .C(men_men_n116_), .Y(men_men_n577_));
  NO4        u0549(.A(n), .B(d), .C(men_men_n120_), .D(a), .Y(men_men_n578_));
  NO2        u0550(.A(c), .B(men_men_n155_), .Y(men_men_n579_));
  NO2        u0551(.A(men_men_n579_), .B(men_men_n578_), .Y(men_men_n580_));
  NOi32      u0552(.An(u), .Bn(f), .C(i), .Y(men_men_n581_));
  AOI220     u0553(.A0(men_men_n581_), .A1(men_men_n102_), .B0(men_men_n563_), .B1(f), .Y(men_men_n582_));
  NO2        u0554(.A(men_men_n291_), .B(men_men_n49_), .Y(men_men_n583_));
  NO2        u0555(.A(men_men_n582_), .B(men_men_n580_), .Y(men_men_n584_));
  AOI210     u0556(.A0(men_men_n577_), .A1(men_men_n574_), .B0(men_men_n584_), .Y(men_men_n585_));
  NA2        u0557(.A(men_men_n146_), .B(men_men_n34_), .Y(men_men_n586_));
  OAI220     u0558(.A0(men_men_n586_), .A1(m), .B0(men_men_n567_), .B1(men_men_n245_), .Y(men_men_n587_));
  NOi41      u0559(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n588_));
  NAi32      u0560(.An(e), .Bn(b), .C(c), .Y(men_men_n589_));
  OR2        u0561(.A(men_men_n589_), .B(men_men_n86_), .Y(men_men_n590_));
  AN2        u0562(.A(men_men_n361_), .B(men_men_n339_), .Y(men_men_n591_));
  NA2        u0563(.A(men_men_n591_), .B(men_men_n590_), .Y(men_men_n592_));
  OA210      u0564(.A0(men_men_n592_), .A1(men_men_n588_), .B0(men_men_n587_), .Y(men_men_n593_));
  OAI220     u0565(.A0(men_men_n425_), .A1(men_men_n424_), .B0(men_men_n561_), .B1(men_men_n560_), .Y(men_men_n594_));
  NAi31      u0566(.An(d), .B(c), .C(a), .Y(men_men_n595_));
  NO2        u0567(.A(men_men_n595_), .B(n), .Y(men_men_n596_));
  NA3        u0568(.A(men_men_n596_), .B(men_men_n594_), .C(e), .Y(men_men_n597_));
  NO3        u0569(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n225_), .Y(men_men_n598_));
  NO2        u0570(.A(men_men_n242_), .B(men_men_n114_), .Y(men_men_n599_));
  OAI210     u0571(.A0(men_men_n598_), .A1(men_men_n426_), .B0(men_men_n599_), .Y(men_men_n600_));
  NA2        u0572(.A(men_men_n600_), .B(men_men_n597_), .Y(men_men_n601_));
  NO2        u0573(.A(men_men_n293_), .B(n), .Y(men_men_n602_));
  NO2        u0574(.A(men_men_n456_), .B(men_men_n602_), .Y(men_men_n603_));
  NA2        u0575(.A(men_men_n594_), .B(f), .Y(men_men_n604_));
  NAi32      u0576(.An(d), .Bn(a), .C(b), .Y(men_men_n605_));
  NO2        u0577(.A(men_men_n605_), .B(men_men_n49_), .Y(men_men_n606_));
  NA2        u0578(.A(h), .B(f), .Y(men_men_n607_));
  NO2        u0579(.A(men_men_n607_), .B(men_men_n97_), .Y(men_men_n608_));
  NO3        u0580(.A(men_men_n185_), .B(men_men_n182_), .C(u), .Y(men_men_n609_));
  AOI220     u0581(.A0(men_men_n609_), .A1(men_men_n58_), .B0(men_men_n608_), .B1(men_men_n606_), .Y(men_men_n610_));
  OAI210     u0582(.A0(men_men_n604_), .A1(men_men_n603_), .B0(men_men_n610_), .Y(men_men_n611_));
  AN3        u0583(.A(j), .B(h), .C(u), .Y(men_men_n612_));
  NO2        u0584(.A(men_men_n152_), .B(c), .Y(men_men_n613_));
  NA3        u0585(.A(men_men_n613_), .B(men_men_n612_), .C(men_men_n488_), .Y(men_men_n614_));
  NA3        u0586(.A(f), .B(d), .C(b), .Y(men_men_n615_));
  NO4        u0587(.A(men_men_n615_), .B(men_men_n185_), .C(men_men_n182_), .D(u), .Y(men_men_n616_));
  NAi21      u0588(.An(men_men_n616_), .B(men_men_n614_), .Y(men_men_n617_));
  NO4        u0589(.A(men_men_n617_), .B(men_men_n611_), .C(men_men_n601_), .D(men_men_n593_), .Y(men_men_n618_));
  AN4        u0590(.A(men_men_n618_), .B(men_men_n585_), .C(men_men_n571_), .D(men_men_n564_), .Y(men_men_n619_));
  INV        u0591(.A(k), .Y(men_men_n620_));
  NA3        u0592(.A(l), .B(men_men_n620_), .C(i), .Y(men_men_n621_));
  INV        u0593(.A(men_men_n621_), .Y(men_men_n622_));
  NA4        u0594(.A(men_men_n422_), .B(men_men_n445_), .C(men_men_n190_), .D(men_men_n117_), .Y(men_men_n623_));
  NAi32      u0595(.An(h), .Bn(f), .C(u), .Y(men_men_n624_));
  NAi41      u0596(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n625_));
  OAI210     u0597(.A0(men_men_n569_), .A1(n), .B0(men_men_n625_), .Y(men_men_n626_));
  NA2        u0598(.A(men_men_n626_), .B(m), .Y(men_men_n627_));
  NAi31      u0599(.An(h), .B(u), .C(f), .Y(men_men_n628_));
  OR3        u0600(.A(men_men_n628_), .B(men_men_n293_), .C(men_men_n49_), .Y(men_men_n629_));
  NA4        u0601(.A(men_men_n445_), .B(men_men_n125_), .C(men_men_n117_), .D(e), .Y(men_men_n630_));
  AN2        u0602(.A(men_men_n630_), .B(men_men_n629_), .Y(men_men_n631_));
  OA210      u0603(.A0(men_men_n627_), .A1(men_men_n624_), .B0(men_men_n631_), .Y(men_men_n632_));
  NO3        u0604(.A(men_men_n624_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n633_));
  NO4        u0605(.A(men_men_n628_), .B(c), .C(men_men_n155_), .D(men_men_n75_), .Y(men_men_n634_));
  OR2        u0606(.A(men_men_n634_), .B(men_men_n633_), .Y(men_men_n635_));
  NAi31      u0607(.An(men_men_n635_), .B(men_men_n632_), .C(men_men_n623_), .Y(men_men_n636_));
  NAi31      u0608(.An(f), .B(h), .C(u), .Y(men_men_n637_));
  NO4        u0609(.A(men_men_n330_), .B(men_men_n637_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n638_));
  NOi32      u0610(.An(b), .Bn(a), .C(c), .Y(men_men_n639_));
  NOi41      u0611(.An(men_men_n639_), .B(men_men_n377_), .C(men_men_n69_), .D(men_men_n121_), .Y(men_men_n640_));
  OR2        u0612(.A(men_men_n640_), .B(men_men_n638_), .Y(men_men_n641_));
  NOi32      u0613(.An(d), .Bn(a), .C(e), .Y(men_men_n642_));
  NA2        u0614(.A(men_men_n642_), .B(men_men_n117_), .Y(men_men_n643_));
  NO2        u0615(.A(n), .B(c), .Y(men_men_n644_));
  NA3        u0616(.A(men_men_n644_), .B(men_men_n29_), .C(m), .Y(men_men_n645_));
  NAi32      u0617(.An(n), .Bn(f), .C(m), .Y(men_men_n646_));
  NA3        u0618(.A(men_men_n646_), .B(men_men_n645_), .C(men_men_n643_), .Y(men_men_n647_));
  NOi32      u0619(.An(e), .Bn(a), .C(d), .Y(men_men_n648_));
  AOI210     u0620(.A0(men_men_n29_), .A1(d), .B0(men_men_n648_), .Y(men_men_n649_));
  AOI210     u0621(.A0(men_men_n649_), .A1(men_men_n224_), .B0(men_men_n586_), .Y(men_men_n650_));
  AOI210     u0622(.A0(men_men_n650_), .A1(men_men_n647_), .B0(men_men_n641_), .Y(men_men_n651_));
  OAI210     u0623(.A0(men_men_n262_), .A1(men_men_n89_), .B0(men_men_n651_), .Y(men_men_n652_));
  AOI210     u0624(.A0(men_men_n636_), .A1(men_men_n622_), .B0(men_men_n652_), .Y(men_men_n653_));
  NO3        u0625(.A(men_men_n337_), .B(men_men_n61_), .C(n), .Y(men_men_n654_));
  NA3        u0626(.A(men_men_n544_), .B(men_men_n180_), .C(men_men_n179_), .Y(men_men_n655_));
  NA2        u0627(.A(men_men_n490_), .B(men_men_n242_), .Y(men_men_n656_));
  OR2        u0628(.A(men_men_n656_), .B(men_men_n655_), .Y(men_men_n657_));
  NA2        u0629(.A(men_men_n76_), .B(men_men_n117_), .Y(men_men_n658_));
  NO2        u0630(.A(men_men_n658_), .B(men_men_n45_), .Y(men_men_n659_));
  AOI220     u0631(.A0(men_men_n659_), .A1(men_men_n574_), .B0(men_men_n657_), .B1(men_men_n654_), .Y(men_men_n660_));
  NO2        u0632(.A(men_men_n660_), .B(men_men_n89_), .Y(men_men_n661_));
  NA3        u0633(.A(men_men_n588_), .B(men_men_n363_), .C(men_men_n46_), .Y(men_men_n662_));
  NOi32      u0634(.An(e), .Bn(c), .C(f), .Y(men_men_n663_));
  NOi21      u0635(.An(f), .B(u), .Y(men_men_n664_));
  NO2        u0636(.A(men_men_n664_), .B(men_men_n222_), .Y(men_men_n665_));
  AOI220     u0637(.A0(men_men_n665_), .A1(men_men_n419_), .B0(men_men_n663_), .B1(men_men_n184_), .Y(men_men_n666_));
  NA3        u0638(.A(men_men_n666_), .B(men_men_n662_), .C(men_men_n187_), .Y(men_men_n667_));
  AOI210     u0639(.A0(men_men_n573_), .A1(men_men_n423_), .B0(men_men_n318_), .Y(men_men_n668_));
  NA2        u0640(.A(men_men_n668_), .B(men_men_n279_), .Y(men_men_n669_));
  NOi21      u0641(.An(j), .B(l), .Y(men_men_n670_));
  NAi21      u0642(.An(k), .B(h), .Y(men_men_n671_));
  NO2        u0643(.A(men_men_n671_), .B(men_men_n277_), .Y(men_men_n672_));
  NA2        u0644(.A(men_men_n672_), .B(men_men_n670_), .Y(men_men_n673_));
  OR2        u0645(.A(men_men_n673_), .B(men_men_n627_), .Y(men_men_n674_));
  NOi31      u0646(.An(m), .B(n), .C(k), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n670_), .B(men_men_n675_), .Y(men_men_n676_));
  AOI210     u0648(.A0(men_men_n423_), .A1(men_men_n397_), .B0(men_men_n318_), .Y(men_men_n677_));
  NAi21      u0649(.An(men_men_n676_), .B(men_men_n677_), .Y(men_men_n678_));
  NO2        u0650(.A(men_men_n293_), .B(men_men_n49_), .Y(men_men_n679_));
  NO2        u0651(.A(men_men_n330_), .B(men_men_n637_), .Y(men_men_n680_));
  NO2        u0652(.A(men_men_n569_), .B(men_men_n49_), .Y(men_men_n681_));
  AOI220     u0653(.A0(men_men_n681_), .A1(men_men_n680_), .B0(men_men_n679_), .B1(men_men_n608_), .Y(men_men_n682_));
  NA4        u0654(.A(men_men_n682_), .B(men_men_n678_), .C(men_men_n674_), .D(men_men_n669_), .Y(men_men_n683_));
  NA2        u0655(.A(men_men_n112_), .B(men_men_n36_), .Y(men_men_n684_));
  NO2        u0656(.A(k), .B(men_men_n225_), .Y(men_men_n685_));
  NO2        u0657(.A(men_men_n565_), .B(men_men_n386_), .Y(men_men_n686_));
  NAi31      u0658(.An(men_men_n684_), .B(men_men_n386_), .C(men_men_n685_), .Y(men_men_n687_));
  NO2        u0659(.A(men_men_n567_), .B(men_men_n185_), .Y(men_men_n688_));
  NA3        u0660(.A(men_men_n589_), .B(men_men_n286_), .C(men_men_n150_), .Y(men_men_n689_));
  NA2        u0661(.A(men_men_n540_), .B(men_men_n166_), .Y(men_men_n690_));
  NO3        u0662(.A(men_men_n420_), .B(men_men_n690_), .C(men_men_n89_), .Y(men_men_n691_));
  AOI210     u0663(.A0(men_men_n689_), .A1(men_men_n688_), .B0(men_men_n691_), .Y(men_men_n692_));
  AN3        u0664(.A(f), .B(d), .C(b), .Y(men_men_n693_));
  OAI210     u0665(.A0(men_men_n693_), .A1(men_men_n135_), .B0(n), .Y(men_men_n694_));
  NA3        u0666(.A(men_men_n540_), .B(men_men_n166_), .C(men_men_n225_), .Y(men_men_n695_));
  AOI210     u0667(.A0(men_men_n694_), .A1(men_men_n244_), .B0(men_men_n695_), .Y(men_men_n696_));
  NAi31      u0668(.An(m), .B(n), .C(k), .Y(men_men_n697_));
  OR2        u0669(.A(men_men_n140_), .B(men_men_n61_), .Y(men_men_n698_));
  OAI210     u0670(.A0(men_men_n698_), .A1(men_men_n697_), .B0(men_men_n264_), .Y(men_men_n699_));
  OAI210     u0671(.A0(men_men_n699_), .A1(men_men_n696_), .B0(j), .Y(men_men_n700_));
  NA3        u0672(.A(men_men_n700_), .B(men_men_n692_), .C(men_men_n687_), .Y(men_men_n701_));
  NO4        u0673(.A(men_men_n701_), .B(men_men_n683_), .C(men_men_n667_), .D(men_men_n661_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n407_), .B(men_men_n169_), .Y(men_men_n703_));
  NAi31      u0675(.An(u), .B(h), .C(f), .Y(men_men_n704_));
  OR3        u0676(.A(men_men_n704_), .B(men_men_n293_), .C(n), .Y(men_men_n705_));
  OA210      u0677(.A0(men_men_n569_), .A1(n), .B0(men_men_n625_), .Y(men_men_n706_));
  NA2        u0678(.A(men_men_n443_), .B(men_men_n125_), .Y(men_men_n707_));
  OAI210     u0679(.A0(men_men_n706_), .A1(men_men_n93_), .B0(men_men_n707_), .Y(men_men_n708_));
  NOi21      u0680(.An(men_men_n705_), .B(men_men_n708_), .Y(men_men_n709_));
  AOI210     u0681(.A0(men_men_n709_), .A1(men_men_n703_), .B0(men_men_n562_), .Y(men_men_n710_));
  NO3        u0682(.A(u), .B(men_men_n224_), .C(men_men_n56_), .Y(men_men_n711_));
  NAi21      u0683(.An(h), .B(j), .Y(men_men_n712_));
  OAI210     u0684(.A0(men_men_n112_), .A1(men_men_n419_), .B0(men_men_n711_), .Y(men_men_n713_));
  OR2        u0685(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n639_), .B(men_men_n365_), .Y(men_men_n715_));
  OA220      u0687(.A0(men_men_n676_), .A1(men_men_n715_), .B0(men_men_n673_), .B1(men_men_n714_), .Y(men_men_n716_));
  NA3        u0688(.A(men_men_n559_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n717_));
  AN2        u0689(.A(h), .B(f), .Y(men_men_n718_));
  NA2        u0690(.A(men_men_n718_), .B(men_men_n37_), .Y(men_men_n719_));
  NA2        u0691(.A(men_men_n102_), .B(men_men_n46_), .Y(men_men_n720_));
  OAI220     u0692(.A0(men_men_n720_), .A1(men_men_n354_), .B0(men_men_n719_), .B1(men_men_n495_), .Y(men_men_n721_));
  AOI210     u0693(.A0(men_men_n605_), .A1(men_men_n455_), .B0(men_men_n49_), .Y(men_men_n722_));
  OAI220     u0694(.A0(men_men_n628_), .A1(men_men_n621_), .B0(men_men_n347_), .B1(men_men_n560_), .Y(men_men_n723_));
  AOI210     u0695(.A0(men_men_n723_), .A1(men_men_n722_), .B0(men_men_n721_), .Y(men_men_n724_));
  NA4        u0696(.A(men_men_n724_), .B(men_men_n717_), .C(men_men_n716_), .D(men_men_n713_), .Y(men_men_n725_));
  NO2        u0697(.A(men_men_n266_), .B(f), .Y(men_men_n726_));
  NO2        u0698(.A(men_men_n664_), .B(men_men_n61_), .Y(men_men_n727_));
  NO3        u0699(.A(men_men_n727_), .B(men_men_n726_), .C(men_men_n34_), .Y(men_men_n728_));
  NA2        u0700(.A(men_men_n350_), .B(men_men_n146_), .Y(men_men_n729_));
  NA2        u0701(.A(men_men_n137_), .B(men_men_n49_), .Y(men_men_n730_));
  AOI220     u0702(.A0(men_men_n730_), .A1(men_men_n565_), .B0(men_men_n386_), .B1(men_men_n117_), .Y(men_men_n731_));
  OA220      u0703(.A0(men_men_n731_), .A1(men_men_n586_), .B0(men_men_n384_), .B1(men_men_n115_), .Y(men_men_n732_));
  OAI210     u0704(.A0(men_men_n729_), .A1(men_men_n728_), .B0(men_men_n732_), .Y(men_men_n733_));
  NO3        u0705(.A(men_men_n430_), .B(men_men_n202_), .C(men_men_n201_), .Y(men_men_n734_));
  NA2        u0706(.A(men_men_n734_), .B(men_men_n242_), .Y(men_men_n735_));
  NA3        u0707(.A(men_men_n735_), .B(men_men_n268_), .C(j), .Y(men_men_n736_));
  NO3        u0708(.A(men_men_n490_), .B(men_men_n182_), .C(i), .Y(men_men_n737_));
  NA2        u0709(.A(men_men_n494_), .B(men_men_n86_), .Y(men_men_n738_));
  NO4        u0710(.A(men_men_n562_), .B(men_men_n738_), .C(men_men_n136_), .D(men_men_n224_), .Y(men_men_n739_));
  INV        u0711(.A(men_men_n739_), .Y(men_men_n740_));
  NA4        u0712(.A(men_men_n740_), .B(men_men_n736_), .C(men_men_n547_), .D(men_men_n428_), .Y(men_men_n741_));
  NO4        u0713(.A(men_men_n741_), .B(men_men_n733_), .C(men_men_n725_), .D(men_men_n710_), .Y(men_men_n742_));
  NA4        u0714(.A(men_men_n742_), .B(men_men_n702_), .C(men_men_n653_), .D(men_men_n619_), .Y(men08));
  NO2        u0715(.A(k), .B(h), .Y(men_men_n744_));
  AO210      u0716(.A0(men_men_n266_), .A1(men_men_n479_), .B0(men_men_n744_), .Y(men_men_n745_));
  NO2        u0717(.A(men_men_n745_), .B(men_men_n316_), .Y(men_men_n746_));
  NA2        u0718(.A(men_men_n663_), .B(men_men_n86_), .Y(men_men_n747_));
  NA2        u0719(.A(men_men_n747_), .B(men_men_n490_), .Y(men_men_n748_));
  AOI210     u0720(.A0(men_men_n748_), .A1(men_men_n746_), .B0(men_men_n524_), .Y(men_men_n749_));
  NO2        u0721(.A(a), .B(men_men_n57_), .Y(men_men_n750_));
  NO4        u0722(.A(men_men_n404_), .B(men_men_n116_), .C(j), .D(men_men_n225_), .Y(men_men_n751_));
  NA2        u0723(.A(men_men_n615_), .B(men_men_n244_), .Y(men_men_n752_));
  AOI220     u0724(.A0(men_men_n752_), .A1(men_men_n371_), .B0(men_men_n751_), .B1(men_men_n750_), .Y(men_men_n753_));
  AOI210     u0725(.A0(men_men_n615_), .A1(men_men_n162_), .B0(men_men_n86_), .Y(men_men_n754_));
  NA4        u0726(.A(men_men_n227_), .B(men_men_n146_), .C(men_men_n45_), .D(h), .Y(men_men_n755_));
  AN2        u0727(.A(l), .B(k), .Y(men_men_n756_));
  NA4        u0728(.A(men_men_n756_), .B(men_men_n112_), .C(men_men_n75_), .D(men_men_n225_), .Y(men_men_n757_));
  OAI210     u0729(.A0(men_men_n755_), .A1(u), .B0(men_men_n757_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n758_), .B(men_men_n754_), .Y(men_men_n759_));
  NA4        u0731(.A(men_men_n759_), .B(men_men_n753_), .C(men_men_n749_), .D(men_men_n373_), .Y(men_men_n760_));
  AN2        u0732(.A(men_men_n570_), .B(men_men_n98_), .Y(men_men_n761_));
  NO4        u0733(.A(men_men_n182_), .B(men_men_n418_), .C(men_men_n116_), .D(u), .Y(men_men_n762_));
  AOI210     u0734(.A0(men_men_n762_), .A1(men_men_n752_), .B0(men_men_n554_), .Y(men_men_n763_));
  NO2        u0735(.A(men_men_n38_), .B(men_men_n224_), .Y(men_men_n764_));
  AOI220     u0736(.A0(men_men_n665_), .A1(men_men_n370_), .B0(men_men_n764_), .B1(men_men_n602_), .Y(men_men_n765_));
  NAi31      u0737(.An(men_men_n761_), .B(men_men_n765_), .C(men_men_n763_), .Y(men_men_n766_));
  NO2        u0738(.A(men_men_n573_), .B(men_men_n35_), .Y(men_men_n767_));
  OAI210     u0739(.A0(men_men_n589_), .A1(men_men_n47_), .B0(men_men_n698_), .Y(men_men_n768_));
  AOI210     u0740(.A0(n), .A1(men_men_n768_), .B0(men_men_n767_), .Y(men_men_n769_));
  NO3        u0741(.A(men_men_n337_), .B(men_men_n136_), .C(men_men_n41_), .Y(men_men_n770_));
  NAi21      u0742(.An(men_men_n770_), .B(men_men_n757_), .Y(men_men_n771_));
  NA2        u0743(.A(men_men_n745_), .B(men_men_n141_), .Y(men_men_n772_));
  AOI220     u0744(.A0(men_men_n772_), .A1(men_men_n429_), .B0(men_men_n771_), .B1(men_men_n78_), .Y(men_men_n773_));
  OAI210     u0745(.A0(men_men_n769_), .A1(men_men_n89_), .B0(men_men_n773_), .Y(men_men_n774_));
  NA2        u0746(.A(men_men_n386_), .B(men_men_n43_), .Y(men_men_n775_));
  NA3        u0747(.A(men_men_n735_), .B(men_men_n356_), .C(men_men_n410_), .Y(men_men_n776_));
  NA2        u0748(.A(men_men_n756_), .B(men_men_n232_), .Y(men_men_n777_));
  NO2        u0749(.A(men_men_n777_), .B(men_men_n349_), .Y(men_men_n778_));
  AOI210     u0750(.A0(men_men_n778_), .A1(men_men_n726_), .B0(men_men_n523_), .Y(men_men_n779_));
  NA3        u0751(.A(m), .B(l), .C(k), .Y(men_men_n780_));
  AOI210     u0752(.A0(men_men_n707_), .A1(men_men_n705_), .B0(men_men_n780_), .Y(men_men_n781_));
  NO2        u0753(.A(men_men_n572_), .B(men_men_n287_), .Y(men_men_n782_));
  NOi21      u0754(.An(men_men_n782_), .B(men_men_n566_), .Y(men_men_n783_));
  NA4        u0755(.A(men_men_n117_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n784_));
  NA3        u0756(.A(men_men_n125_), .B(men_men_n438_), .C(i), .Y(men_men_n785_));
  NO2        u0757(.A(men_men_n785_), .B(men_men_n784_), .Y(men_men_n786_));
  NO3        u0758(.A(men_men_n786_), .B(men_men_n783_), .C(men_men_n781_), .Y(men_men_n787_));
  NA4        u0759(.A(men_men_n787_), .B(men_men_n779_), .C(men_men_n776_), .D(men_men_n775_), .Y(men_men_n788_));
  NO4        u0760(.A(men_men_n788_), .B(men_men_n774_), .C(men_men_n766_), .D(men_men_n760_), .Y(men_men_n789_));
  NA2        u0761(.A(men_men_n665_), .B(men_men_n419_), .Y(men_men_n790_));
  NOi31      u0762(.An(u), .B(h), .C(f), .Y(men_men_n791_));
  NA2        u0763(.A(men_men_n681_), .B(men_men_n791_), .Y(men_men_n792_));
  AO210      u0764(.A0(men_men_n792_), .A1(men_men_n629_), .B0(men_men_n575_), .Y(men_men_n793_));
  NO3        u0765(.A(men_men_n423_), .B(men_men_n560_), .C(h), .Y(men_men_n794_));
  AOI210     u0766(.A0(men_men_n794_), .A1(men_men_n117_), .B0(men_men_n533_), .Y(men_men_n795_));
  NA4        u0767(.A(men_men_n795_), .B(men_men_n793_), .C(men_men_n790_), .D(men_men_n265_), .Y(men_men_n796_));
  NA2        u0768(.A(men_men_n756_), .B(men_men_n75_), .Y(men_men_n797_));
  NO4        u0769(.A(men_men_n734_), .B(men_men_n182_), .C(n), .D(i), .Y(men_men_n798_));
  NOi21      u0770(.An(h), .B(j), .Y(men_men_n799_));
  NA2        u0771(.A(men_men_n799_), .B(f), .Y(men_men_n800_));
  NO2        u0772(.A(men_men_n800_), .B(men_men_n259_), .Y(men_men_n801_));
  NO3        u0773(.A(men_men_n801_), .B(men_men_n798_), .C(men_men_n737_), .Y(men_men_n802_));
  OAI220     u0774(.A0(men_men_n802_), .A1(men_men_n797_), .B0(men_men_n631_), .B1(men_men_n62_), .Y(men_men_n803_));
  NO2        u0775(.A(men_men_n796_), .B(men_men_n803_), .Y(men_men_n804_));
  NO2        u0776(.A(j), .B(i), .Y(men_men_n805_));
  NA3        u0777(.A(men_men_n805_), .B(men_men_n82_), .C(l), .Y(men_men_n806_));
  NA2        u0778(.A(men_men_n805_), .B(men_men_n33_), .Y(men_men_n807_));
  NA2        u0779(.A(men_men_n448_), .B(men_men_n125_), .Y(men_men_n808_));
  OA220      u0780(.A0(men_men_n808_), .A1(men_men_n807_), .B0(men_men_n806_), .B1(men_men_n627_), .Y(men_men_n809_));
  NO3        u0781(.A(men_men_n157_), .B(men_men_n49_), .C(men_men_n114_), .Y(men_men_n810_));
  NO3        u0782(.A(c), .B(men_men_n155_), .C(men_men_n75_), .Y(men_men_n811_));
  NO3        u0783(.A(men_men_n517_), .B(men_men_n466_), .C(j), .Y(men_men_n812_));
  OAI210     u0784(.A0(men_men_n811_), .A1(men_men_n810_), .B0(men_men_n812_), .Y(men_men_n813_));
  OAI210     u0785(.A0(men_men_n792_), .A1(men_men_n62_), .B0(men_men_n813_), .Y(men_men_n814_));
  NA2        u0786(.A(k), .B(j), .Y(men_men_n815_));
  NO3        u0787(.A(men_men_n316_), .B(men_men_n815_), .C(men_men_n40_), .Y(men_men_n816_));
  AOI210     u0788(.A0(men_men_n565_), .A1(n), .B0(men_men_n588_), .Y(men_men_n817_));
  NA2        u0789(.A(men_men_n817_), .B(men_men_n591_), .Y(men_men_n818_));
  AN3        u0790(.A(men_men_n818_), .B(men_men_n816_), .C(men_men_n101_), .Y(men_men_n819_));
  NO3        u0791(.A(men_men_n182_), .B(men_men_n418_), .C(men_men_n116_), .Y(men_men_n820_));
  AOI220     u0792(.A0(men_men_n820_), .A1(men_men_n260_), .B0(men_men_n656_), .B1(men_men_n327_), .Y(men_men_n821_));
  NAi21      u0793(.An(men_men_n649_), .B(men_men_n95_), .Y(men_men_n822_));
  NA2        u0794(.A(men_men_n822_), .B(men_men_n821_), .Y(men_men_n823_));
  NO2        u0795(.A(men_men_n316_), .B(men_men_n141_), .Y(men_men_n824_));
  AOI220     u0796(.A0(men_men_n824_), .A1(men_men_n665_), .B0(men_men_n770_), .B1(men_men_n754_), .Y(men_men_n825_));
  NO2        u0797(.A(men_men_n780_), .B(men_men_n93_), .Y(men_men_n826_));
  NA2        u0798(.A(men_men_n826_), .B(men_men_n626_), .Y(men_men_n827_));
  NO2        u0799(.A(men_men_n628_), .B(men_men_n121_), .Y(men_men_n828_));
  OAI210     u0800(.A0(men_men_n828_), .A1(men_men_n812_), .B0(men_men_n722_), .Y(men_men_n829_));
  NA3        u0801(.A(men_men_n829_), .B(men_men_n827_), .C(men_men_n825_), .Y(men_men_n830_));
  OR4        u0802(.A(men_men_n830_), .B(men_men_n823_), .C(men_men_n819_), .D(men_men_n814_), .Y(men_men_n831_));
  NA3        u0803(.A(men_men_n817_), .B(men_men_n591_), .C(men_men_n590_), .Y(men_men_n832_));
  NA4        u0804(.A(men_men_n832_), .B(men_men_n227_), .C(men_men_n479_), .D(men_men_n34_), .Y(men_men_n833_));
  NO4        u0805(.A(men_men_n517_), .B(men_men_n462_), .C(j), .D(f), .Y(men_men_n834_));
  OAI220     u0806(.A0(men_men_n755_), .A1(men_men_n747_), .B0(men_men_n354_), .B1(men_men_n38_), .Y(men_men_n835_));
  AOI210     u0807(.A0(men_men_n834_), .A1(men_men_n272_), .B0(men_men_n835_), .Y(men_men_n836_));
  NA3        u0808(.A(men_men_n581_), .B(men_men_n309_), .C(h), .Y(men_men_n837_));
  NOi21      u0809(.An(men_men_n722_), .B(men_men_n837_), .Y(men_men_n838_));
  NO2        u0810(.A(men_men_n94_), .B(men_men_n47_), .Y(men_men_n839_));
  OAI220     u0811(.A0(men_men_n837_), .A1(men_men_n645_), .B0(men_men_n806_), .B1(men_men_n714_), .Y(men_men_n840_));
  AOI210     u0812(.A0(men_men_n839_), .A1(men_men_n386_), .B0(men_men_n840_), .Y(men_men_n841_));
  NAi41      u0813(.An(men_men_n838_), .B(men_men_n841_), .C(men_men_n836_), .D(men_men_n833_), .Y(men_men_n842_));
  OR2        u0814(.A(men_men_n826_), .B(men_men_n98_), .Y(men_men_n843_));
  AOI220     u0815(.A0(men_men_n843_), .A1(men_men_n250_), .B0(men_men_n812_), .B1(men_men_n679_), .Y(men_men_n844_));
  NO2        u0816(.A(men_men_n706_), .B(men_men_n75_), .Y(men_men_n845_));
  AOI210     u0817(.A0(men_men_n834_), .A1(men_men_n845_), .B0(men_men_n358_), .Y(men_men_n846_));
  OAI210     u0818(.A0(men_men_n780_), .A1(men_men_n704_), .B0(men_men_n553_), .Y(men_men_n847_));
  NA3        u0819(.A(men_men_n263_), .B(men_men_n59_), .C(b), .Y(men_men_n848_));
  AOI220     u0820(.A0(men_men_n644_), .A1(men_men_n29_), .B0(men_men_n494_), .B1(men_men_n86_), .Y(men_men_n849_));
  NA2        u0821(.A(men_men_n849_), .B(men_men_n848_), .Y(men_men_n850_));
  NO2        u0822(.A(men_men_n837_), .B(men_men_n522_), .Y(men_men_n851_));
  AOI210     u0823(.A0(men_men_n850_), .A1(men_men_n847_), .B0(men_men_n851_), .Y(men_men_n852_));
  NA3        u0824(.A(men_men_n852_), .B(men_men_n846_), .C(men_men_n844_), .Y(men_men_n853_));
  NOi41      u0825(.An(men_men_n809_), .B(men_men_n853_), .C(men_men_n842_), .D(men_men_n831_), .Y(men_men_n854_));
  OR3        u0826(.A(men_men_n755_), .B(men_men_n244_), .C(u), .Y(men_men_n855_));
  NO3        u0827(.A(men_men_n364_), .B(men_men_n318_), .C(men_men_n116_), .Y(men_men_n856_));
  NA2        u0828(.A(men_men_n856_), .B(men_men_n818_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n858_));
  NO3        u0830(.A(men_men_n858_), .B(men_men_n807_), .C(men_men_n293_), .Y(men_men_n859_));
  NO3        u0831(.A(men_men_n560_), .B(men_men_n96_), .C(h), .Y(men_men_n860_));
  AOI210     u0832(.A0(men_men_n860_), .A1(men_men_n750_), .B0(men_men_n859_), .Y(men_men_n861_));
  NA4        u0833(.A(men_men_n861_), .B(men_men_n857_), .C(men_men_n855_), .D(men_men_n431_), .Y(men_men_n862_));
  OR2        u0834(.A(men_men_n704_), .B(men_men_n94_), .Y(men_men_n863_));
  NOi31      u0835(.An(b), .B(d), .C(a), .Y(men_men_n864_));
  NO2        u0836(.A(men_men_n864_), .B(men_men_n642_), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n865_), .B(n), .Y(men_men_n866_));
  NOi21      u0838(.An(men_men_n849_), .B(men_men_n866_), .Y(men_men_n867_));
  OAI220     u0839(.A0(men_men_n867_), .A1(men_men_n863_), .B0(men_men_n837_), .B1(men_men_n643_), .Y(men_men_n868_));
  NO2        u0840(.A(men_men_n589_), .B(men_men_n86_), .Y(men_men_n869_));
  NO3        u0841(.A(men_men_n664_), .B(men_men_n349_), .C(men_men_n121_), .Y(men_men_n870_));
  NOi21      u0842(.An(men_men_n870_), .B(men_men_n167_), .Y(men_men_n871_));
  AOI210     u0843(.A0(men_men_n856_), .A1(men_men_n869_), .B0(men_men_n871_), .Y(men_men_n872_));
  OAI210     u0844(.A0(men_men_n755_), .A1(men_men_n420_), .B0(men_men_n872_), .Y(men_men_n873_));
  NO2        u0845(.A(men_men_n734_), .B(n), .Y(men_men_n874_));
  AOI220     u0846(.A0(men_men_n824_), .A1(men_men_n711_), .B0(men_men_n874_), .B1(men_men_n746_), .Y(men_men_n875_));
  NO2        u0847(.A(men_men_n344_), .B(men_men_n249_), .Y(men_men_n876_));
  OAI210     u0848(.A0(men_men_n98_), .A1(men_men_n95_), .B0(men_men_n876_), .Y(men_men_n877_));
  NA2        u0849(.A(men_men_n125_), .B(men_men_n86_), .Y(men_men_n878_));
  AOI210     u0850(.A0(men_men_n452_), .A1(men_men_n444_), .B0(men_men_n878_), .Y(men_men_n879_));
  NAi21      u0851(.An(men_men_n879_), .B(men_men_n877_), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n778_), .B(men_men_n34_), .Y(men_men_n881_));
  NAi21      u0853(.An(men_men_n784_), .B(men_men_n463_), .Y(men_men_n882_));
  NO2        u0854(.A(men_men_n287_), .B(i), .Y(men_men_n883_));
  NA2        u0855(.A(men_men_n762_), .B(men_men_n372_), .Y(men_men_n884_));
  OAI210     u0856(.A0(men_men_n634_), .A1(men_men_n633_), .B0(men_men_n387_), .Y(men_men_n885_));
  AN3        u0857(.A(men_men_n885_), .B(men_men_n884_), .C(men_men_n882_), .Y(men_men_n886_));
  NAi41      u0858(.An(men_men_n880_), .B(men_men_n886_), .C(men_men_n881_), .D(men_men_n875_), .Y(men_men_n887_));
  NO4        u0859(.A(men_men_n887_), .B(men_men_n873_), .C(men_men_n868_), .D(men_men_n862_), .Y(men_men_n888_));
  NA4        u0860(.A(men_men_n888_), .B(men_men_n854_), .C(men_men_n804_), .D(men_men_n789_), .Y(men09));
  INV        u0861(.A(men_men_n126_), .Y(men_men_n890_));
  NA2        u0862(.A(f), .B(e), .Y(men_men_n891_));
  NO2        u0863(.A(men_men_n237_), .B(men_men_n116_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n892_), .B(u), .Y(men_men_n893_));
  NA4        u0865(.A(men_men_n330_), .B(men_men_n503_), .C(men_men_n275_), .D(men_men_n123_), .Y(men_men_n894_));
  AOI210     u0866(.A0(men_men_n894_), .A1(u), .B0(men_men_n500_), .Y(men_men_n895_));
  AOI210     u0867(.A0(men_men_n895_), .A1(men_men_n893_), .B0(men_men_n891_), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n472_), .B(e), .Y(men_men_n897_));
  NO2        u0869(.A(men_men_n897_), .B(men_men_n544_), .Y(men_men_n898_));
  AOI210     u0870(.A0(men_men_n896_), .A1(men_men_n890_), .B0(men_men_n898_), .Y(men_men_n899_));
  NO2        u0871(.A(men_men_n214_), .B(men_men_n224_), .Y(men_men_n900_));
  NA3        u0872(.A(m), .B(l), .C(i), .Y(men_men_n901_));
  OAI220     u0873(.A0(men_men_n628_), .A1(men_men_n901_), .B0(men_men_n377_), .B1(men_men_n561_), .Y(men_men_n902_));
  NA4        u0874(.A(men_men_n90_), .B(men_men_n89_), .C(u), .D(f), .Y(men_men_n903_));
  NAi31      u0875(.An(men_men_n902_), .B(men_men_n903_), .C(men_men_n467_), .Y(men_men_n904_));
  OA210      u0876(.A0(men_men_n904_), .A1(men_men_n900_), .B0(men_men_n602_), .Y(men_men_n905_));
  NA3        u0877(.A(men_men_n863_), .B(men_men_n604_), .C(men_men_n553_), .Y(men_men_n906_));
  OA210      u0878(.A0(men_men_n906_), .A1(men_men_n905_), .B0(men_men_n866_), .Y(men_men_n907_));
  INV        u0879(.A(men_men_n361_), .Y(men_men_n908_));
  NO2        u0880(.A(men_men_n132_), .B(men_men_n130_), .Y(men_men_n909_));
  NOi31      u0881(.An(k), .B(m), .C(l), .Y(men_men_n910_));
  NO2        u0882(.A(men_men_n363_), .B(men_men_n910_), .Y(men_men_n911_));
  AOI210     u0883(.A0(men_men_n911_), .A1(men_men_n909_), .B0(men_men_n637_), .Y(men_men_n912_));
  NA2        u0884(.A(men_men_n848_), .B(men_men_n354_), .Y(men_men_n913_));
  NA2        u0885(.A(men_men_n365_), .B(men_men_n367_), .Y(men_men_n914_));
  OAI210     u0886(.A0(men_men_n214_), .A1(men_men_n224_), .B0(men_men_n914_), .Y(men_men_n915_));
  AOI220     u0887(.A0(men_men_n915_), .A1(men_men_n913_), .B0(men_men_n912_), .B1(men_men_n908_), .Y(men_men_n916_));
  NA2        u0888(.A(men_men_n176_), .B(men_men_n118_), .Y(men_men_n917_));
  NA3        u0889(.A(men_men_n917_), .B(men_men_n745_), .C(men_men_n141_), .Y(men_men_n918_));
  NA3        u0890(.A(men_men_n918_), .B(men_men_n199_), .C(men_men_n31_), .Y(men_men_n919_));
  NA4        u0891(.A(men_men_n919_), .B(men_men_n916_), .C(men_men_n666_), .D(men_men_n84_), .Y(men_men_n920_));
  NO2        u0892(.A(men_men_n624_), .B(men_men_n530_), .Y(men_men_n921_));
  NA2        u0893(.A(men_men_n921_), .B(men_men_n199_), .Y(men_men_n922_));
  NOi21      u0894(.An(f), .B(d), .Y(men_men_n923_));
  NA2        u0895(.A(men_men_n923_), .B(m), .Y(men_men_n924_));
  NO2        u0896(.A(men_men_n924_), .B(men_men_n52_), .Y(men_men_n925_));
  NOi32      u0897(.An(u), .Bn(f), .C(d), .Y(men_men_n926_));
  NA4        u0898(.A(men_men_n926_), .B(men_men_n644_), .C(men_men_n29_), .D(m), .Y(men_men_n927_));
  NOi21      u0899(.An(men_men_n331_), .B(men_men_n927_), .Y(men_men_n928_));
  AOI210     u0900(.A0(men_men_n925_), .A1(men_men_n579_), .B0(men_men_n928_), .Y(men_men_n929_));
  NA3        u0901(.A(men_men_n330_), .B(men_men_n275_), .C(men_men_n123_), .Y(men_men_n930_));
  AN2        u0902(.A(f), .B(d), .Y(men_men_n931_));
  NA2        u0903(.A(men_men_n508_), .B(men_men_n931_), .Y(men_men_n932_));
  NO3        u0904(.A(men_men_n932_), .B(men_men_n75_), .C(men_men_n225_), .Y(men_men_n933_));
  NO2        u0905(.A(men_men_n302_), .B(men_men_n56_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n930_), .B(men_men_n933_), .Y(men_men_n935_));
  NAi41      u0907(.An(men_men_n521_), .B(men_men_n935_), .C(men_men_n929_), .D(men_men_n922_), .Y(men_men_n936_));
  NO4        u0908(.A(men_men_n664_), .B(men_men_n137_), .C(men_men_n349_), .D(men_men_n158_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n697_), .B(men_men_n349_), .Y(men_men_n938_));
  AN2        u0910(.A(men_men_n938_), .B(men_men_n726_), .Y(men_men_n939_));
  NO3        u0911(.A(men_men_n939_), .B(men_men_n937_), .C(men_men_n246_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n642_), .B(men_men_n86_), .Y(men_men_n941_));
  OAI220     u0913(.A0(men_men_n914_), .A1(men_men_n941_), .B0(men_men_n848_), .B1(men_men_n467_), .Y(men_men_n942_));
  NA3        u0914(.A(men_men_n166_), .B(men_men_n112_), .C(men_men_n111_), .Y(men_men_n943_));
  OAI220     u0915(.A0(men_men_n932_), .A1(men_men_n457_), .B0(men_men_n361_), .B1(men_men_n943_), .Y(men_men_n944_));
  NOi41      u0916(.An(men_men_n235_), .B(men_men_n944_), .C(men_men_n942_), .D(men_men_n325_), .Y(men_men_n945_));
  NA3        u0917(.A(men_men_n1666_), .B(men_men_n542_), .C(f), .Y(men_men_n946_));
  OR2        u0918(.A(men_men_n704_), .B(men_men_n576_), .Y(men_men_n947_));
  INV        u0919(.A(men_men_n947_), .Y(men_men_n948_));
  NA2        u0920(.A(men_men_n865_), .B(men_men_n115_), .Y(men_men_n949_));
  NA2        u0921(.A(men_men_n949_), .B(men_men_n948_), .Y(men_men_n950_));
  NA4        u0922(.A(men_men_n950_), .B(men_men_n946_), .C(men_men_n945_), .D(men_men_n940_), .Y(men_men_n951_));
  NO4        u0923(.A(men_men_n951_), .B(men_men_n936_), .C(men_men_n920_), .D(men_men_n907_), .Y(men_men_n952_));
  OR2        u0924(.A(men_men_n932_), .B(men_men_n75_), .Y(men_men_n953_));
  NA2        u0925(.A(men_men_n116_), .B(j), .Y(men_men_n954_));
  NA2        u0926(.A(men_men_n892_), .B(u), .Y(men_men_n955_));
  AOI210     u0927(.A0(men_men_n955_), .A1(men_men_n310_), .B0(men_men_n953_), .Y(men_men_n956_));
  AOI210     u0928(.A0(men_men_n848_), .A1(men_men_n354_), .B0(men_men_n903_), .Y(men_men_n957_));
  NO2        u0929(.A(men_men_n141_), .B(men_men_n137_), .Y(men_men_n958_));
  NO2        u0930(.A(men_men_n242_), .B(men_men_n236_), .Y(men_men_n959_));
  AOI220     u0931(.A0(men_men_n959_), .A1(men_men_n239_), .B0(men_men_n323_), .B1(men_men_n958_), .Y(men_men_n960_));
  NO2        u0932(.A(men_men_n457_), .B(men_men_n891_), .Y(men_men_n961_));
  NA2        u0933(.A(men_men_n961_), .B(men_men_n596_), .Y(men_men_n962_));
  NA2        u0934(.A(men_men_n962_), .B(men_men_n960_), .Y(men_men_n963_));
  NA2        u0935(.A(e), .B(d), .Y(men_men_n964_));
  OAI220     u0936(.A0(men_men_n964_), .A1(c), .B0(men_men_n344_), .B1(d), .Y(men_men_n965_));
  NA3        u0937(.A(men_men_n965_), .B(men_men_n483_), .C(men_men_n540_), .Y(men_men_n966_));
  AOI210     u0938(.A0(men_men_n548_), .A1(men_men_n189_), .B0(men_men_n242_), .Y(men_men_n967_));
  AOI210     u0939(.A0(men_men_n665_), .A1(men_men_n370_), .B0(men_men_n967_), .Y(men_men_n968_));
  NA2        u0940(.A(men_men_n302_), .B(men_men_n172_), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n933_), .B(men_men_n969_), .Y(men_men_n970_));
  NA3        u0942(.A(men_men_n175_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n971_));
  NA4        u0943(.A(men_men_n971_), .B(men_men_n970_), .C(men_men_n968_), .D(men_men_n966_), .Y(men_men_n972_));
  NO4        u0944(.A(men_men_n972_), .B(men_men_n963_), .C(men_men_n957_), .D(men_men_n956_), .Y(men_men_n973_));
  NA2        u0945(.A(men_men_n908_), .B(men_men_n31_), .Y(men_men_n974_));
  AO210      u0946(.A0(men_men_n974_), .A1(men_men_n747_), .B0(men_men_n228_), .Y(men_men_n975_));
  OAI220     u0947(.A0(men_men_n664_), .A1(men_men_n61_), .B0(men_men_n318_), .B1(j), .Y(men_men_n976_));
  AOI220     u0948(.A0(men_men_n976_), .A1(men_men_n938_), .B0(men_men_n654_), .B1(men_men_n663_), .Y(men_men_n977_));
  OAI210     u0949(.A0(men_men_n897_), .A1(men_men_n179_), .B0(men_men_n977_), .Y(men_men_n978_));
  OAI210     u0950(.A0(men_men_n892_), .A1(men_men_n969_), .B0(men_men_n926_), .Y(men_men_n979_));
  NO2        u0951(.A(men_men_n979_), .B(men_men_n645_), .Y(men_men_n980_));
  AOI210     u0952(.A0(men_men_n122_), .A1(men_men_n121_), .B0(men_men_n274_), .Y(men_men_n981_));
  NO2        u0953(.A(men_men_n981_), .B(men_men_n927_), .Y(men_men_n982_));
  AO210      u0954(.A0(men_men_n913_), .A1(men_men_n902_), .B0(men_men_n982_), .Y(men_men_n983_));
  NOi31      u0955(.An(men_men_n579_), .B(men_men_n924_), .C(men_men_n310_), .Y(men_men_n984_));
  NO4        u0956(.A(men_men_n984_), .B(men_men_n983_), .C(men_men_n980_), .D(men_men_n978_), .Y(men_men_n985_));
  AO220      u0957(.A0(men_men_n483_), .A1(men_men_n799_), .B0(men_men_n184_), .B1(f), .Y(men_men_n986_));
  OAI210     u0958(.A0(men_men_n986_), .A1(men_men_n486_), .B0(men_men_n965_), .Y(men_men_n987_));
  NO2        u0959(.A(men_men_n466_), .B(men_men_n71_), .Y(men_men_n988_));
  OAI210     u0960(.A0(men_men_n906_), .A1(men_men_n988_), .B0(men_men_n750_), .Y(men_men_n989_));
  AN4        u0961(.A(men_men_n989_), .B(men_men_n987_), .C(men_men_n985_), .D(men_men_n975_), .Y(men_men_n990_));
  NA4        u0962(.A(men_men_n990_), .B(men_men_n973_), .C(men_men_n952_), .D(men_men_n899_), .Y(men12));
  NO2        u0963(.A(men_men_n482_), .B(c), .Y(men_men_n992_));
  NO4        u0964(.A(men_men_n471_), .B(men_men_n266_), .C(men_men_n620_), .D(men_men_n225_), .Y(men_men_n993_));
  NA2        u0965(.A(men_men_n993_), .B(men_men_n992_), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n579_), .B(men_men_n988_), .Y(men_men_n995_));
  NO3        u0967(.A(men_men_n482_), .B(men_men_n86_), .C(men_men_n120_), .Y(men_men_n996_));
  NO2        u0968(.A(men_men_n909_), .B(men_men_n377_), .Y(men_men_n997_));
  NO2        u0969(.A(men_men_n704_), .B(men_men_n404_), .Y(men_men_n998_));
  AOI220     u0970(.A0(men_men_n998_), .A1(men_men_n578_), .B0(men_men_n997_), .B1(men_men_n996_), .Y(men_men_n999_));
  NA4        u0971(.A(men_men_n999_), .B(men_men_n995_), .C(men_men_n994_), .D(men_men_n470_), .Y(men_men_n1000_));
  AOI210     u0972(.A0(men_men_n245_), .A1(men_men_n360_), .B0(men_men_n211_), .Y(men_men_n1001_));
  OR2        u0973(.A(men_men_n1001_), .B(men_men_n993_), .Y(men_men_n1002_));
  AOI210     u0974(.A0(men_men_n357_), .A1(men_men_n416_), .B0(men_men_n225_), .Y(men_men_n1003_));
  OAI210     u0975(.A0(men_men_n1003_), .A1(men_men_n1002_), .B0(men_men_n430_), .Y(men_men_n1004_));
  NO2        u0976(.A(men_men_n684_), .B(men_men_n277_), .Y(men_men_n1005_));
  NO2        u0977(.A(men_men_n628_), .B(men_men_n901_), .Y(men_men_n1006_));
  AOI220     u0978(.A0(men_men_n1006_), .A1(men_men_n602_), .B0(men_men_n876_), .B1(men_men_n1005_), .Y(men_men_n1007_));
  INV        u0979(.A(men_men_n157_), .Y(men_men_n1008_));
  NA2        u0980(.A(men_men_n1008_), .B(men_men_n252_), .Y(men_men_n1009_));
  NA3        u0981(.A(men_men_n1009_), .B(men_men_n1007_), .C(men_men_n1004_), .Y(men_men_n1010_));
  OR2        u0982(.A(men_men_n345_), .B(men_men_n996_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n1011_), .B(men_men_n378_), .Y(men_men_n1012_));
  NO3        u0984(.A(men_men_n137_), .B(men_men_n158_), .C(men_men_n225_), .Y(men_men_n1013_));
  NA2        u0985(.A(men_men_n1013_), .B(men_men_n565_), .Y(men_men_n1014_));
  NA4        u0986(.A(men_men_n472_), .B(men_men_n464_), .C(men_men_n190_), .D(u), .Y(men_men_n1015_));
  NA3        u0987(.A(men_men_n1015_), .B(men_men_n1014_), .C(men_men_n1012_), .Y(men_men_n1016_));
  NO4        u0988(.A(men_men_n708_), .B(men_men_n1016_), .C(men_men_n1010_), .D(men_men_n1000_), .Y(men_men_n1017_));
  NO2        u0989(.A(men_men_n394_), .B(men_men_n393_), .Y(men_men_n1018_));
  NA2        u0990(.A(men_men_n625_), .B(men_men_n73_), .Y(men_men_n1019_));
  NA2        u0991(.A(men_men_n589_), .B(men_men_n150_), .Y(men_men_n1020_));
  NOi21      u0992(.An(men_men_n34_), .B(men_men_n697_), .Y(men_men_n1021_));
  AOI220     u0993(.A0(men_men_n1021_), .A1(men_men_n1020_), .B0(men_men_n1019_), .B1(men_men_n1018_), .Y(men_men_n1022_));
  OAI210     u0994(.A0(men_men_n264_), .A1(men_men_n45_), .B0(men_men_n1022_), .Y(men_men_n1023_));
  NA2        u0995(.A(men_men_n463_), .B(men_men_n279_), .Y(men_men_n1024_));
  NO3        u0996(.A(men_men_n878_), .B(men_men_n91_), .C(men_men_n435_), .Y(men_men_n1025_));
  NAi31      u0997(.An(men_men_n1025_), .B(men_men_n1024_), .C(men_men_n341_), .Y(men_men_n1026_));
  NO2        u0998(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n1027_));
  NO2        u0999(.A(men_men_n536_), .B(men_men_n318_), .Y(men_men_n1028_));
  NO2        u1000(.A(men_men_n536_), .B(men_men_n150_), .Y(men_men_n1029_));
  NA2        u1001(.A(men_men_n675_), .B(men_men_n387_), .Y(men_men_n1030_));
  OAI210     u1002(.A0(men_men_n785_), .A1(men_men_n1030_), .B0(men_men_n391_), .Y(men_men_n1031_));
  NO4        u1003(.A(men_men_n1031_), .B(men_men_n1029_), .C(men_men_n1026_), .D(men_men_n1023_), .Y(men_men_n1032_));
  NA2        u1004(.A(men_men_n370_), .B(u), .Y(men_men_n1033_));
  NA2        u1005(.A(men_men_n169_), .B(i), .Y(men_men_n1034_));
  NA2        u1006(.A(men_men_n46_), .B(i), .Y(men_men_n1035_));
  OAI220     u1007(.A0(men_men_n1035_), .A1(men_men_n210_), .B0(men_men_n1034_), .B1(men_men_n94_), .Y(men_men_n1036_));
  AOI210     u1008(.A0(men_men_n446_), .A1(men_men_n37_), .B0(men_men_n1036_), .Y(men_men_n1037_));
  NO2        u1009(.A(men_men_n150_), .B(men_men_n86_), .Y(men_men_n1038_));
  OR2        u1010(.A(men_men_n1038_), .B(men_men_n588_), .Y(men_men_n1039_));
  NA2        u1011(.A(men_men_n589_), .B(men_men_n408_), .Y(men_men_n1040_));
  AOI210     u1012(.A0(men_men_n1040_), .A1(n), .B0(men_men_n1039_), .Y(men_men_n1041_));
  OAI220     u1013(.A0(men_men_n1041_), .A1(men_men_n1033_), .B0(men_men_n1037_), .B1(men_men_n354_), .Y(men_men_n1042_));
  NO2        u1014(.A(men_men_n704_), .B(men_men_n530_), .Y(men_men_n1043_));
  NA3        u1015(.A(men_men_n365_), .B(men_men_n670_), .C(i), .Y(men_men_n1044_));
  OAI210     u1016(.A0(men_men_n466_), .A1(men_men_n330_), .B0(men_men_n1044_), .Y(men_men_n1045_));
  OAI220     u1017(.A0(men_men_n1045_), .A1(men_men_n1043_), .B0(men_men_n722_), .B1(men_men_n811_), .Y(men_men_n1046_));
  NA2        u1018(.A(men_men_n648_), .B(men_men_n117_), .Y(men_men_n1047_));
  OR3        u1019(.A(men_men_n330_), .B(men_men_n462_), .C(f), .Y(men_men_n1048_));
  NA3        u1020(.A(men_men_n670_), .B(men_men_n82_), .C(i), .Y(men_men_n1049_));
  OA220      u1021(.A0(men_men_n1049_), .A1(men_men_n1047_), .B0(men_men_n1048_), .B1(men_men_n627_), .Y(men_men_n1050_));
  NA3        u1022(.A(men_men_n346_), .B(men_men_n122_), .C(u), .Y(men_men_n1051_));
  AOI210     u1023(.A0(men_men_n719_), .A1(men_men_n1051_), .B0(m), .Y(men_men_n1052_));
  OAI210     u1024(.A0(men_men_n1052_), .A1(men_men_n997_), .B0(men_men_n345_), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n738_), .B(men_men_n941_), .Y(men_men_n1054_));
  NA2        u1026(.A(men_men_n903_), .B(men_men_n467_), .Y(men_men_n1055_));
  NA2        u1027(.A(men_men_n233_), .B(men_men_n79_), .Y(men_men_n1056_));
  NA3        u1028(.A(men_men_n1056_), .B(men_men_n1049_), .C(men_men_n1048_), .Y(men_men_n1057_));
  AOI220     u1029(.A0(men_men_n1057_), .A1(men_men_n272_), .B0(men_men_n1055_), .B1(men_men_n1054_), .Y(men_men_n1058_));
  NA4        u1030(.A(men_men_n1058_), .B(men_men_n1053_), .C(men_men_n1050_), .D(men_men_n1046_), .Y(men_men_n1059_));
  NO2        u1031(.A(men_men_n404_), .B(men_men_n93_), .Y(men_men_n1060_));
  OAI210     u1032(.A0(men_men_n1060_), .A1(men_men_n1005_), .B0(men_men_n250_), .Y(men_men_n1061_));
  NO2        u1033(.A(men_men_n489_), .B(men_men_n225_), .Y(men_men_n1062_));
  AOI220     u1034(.A0(men_men_n1062_), .A1(men_men_n409_), .B0(men_men_n1011_), .B1(men_men_n229_), .Y(men_men_n1063_));
  AOI220     u1035(.A0(men_men_n998_), .A1(men_men_n1008_), .B0(men_men_n626_), .B1(men_men_n92_), .Y(men_men_n1064_));
  NA3        u1036(.A(men_men_n1064_), .B(men_men_n1063_), .C(men_men_n1061_), .Y(men_men_n1065_));
  OAI210     u1037(.A0(men_men_n1055_), .A1(men_men_n1006_), .B0(men_men_n578_), .Y(men_men_n1066_));
  AOI210     u1038(.A0(men_men_n447_), .A1(men_men_n439_), .B0(men_men_n878_), .Y(men_men_n1067_));
  OAI210     u1039(.A0(men_men_n394_), .A1(men_men_n393_), .B0(men_men_n113_), .Y(men_men_n1068_));
  AOI210     u1040(.A0(men_men_n1068_), .A1(men_men_n570_), .B0(men_men_n1067_), .Y(men_men_n1069_));
  NA2        u1041(.A(men_men_n1052_), .B(men_men_n996_), .Y(men_men_n1070_));
  NO3        u1042(.A(men_men_n954_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1071_));
  AOI220     u1043(.A0(men_men_n1071_), .A1(men_men_n668_), .B0(men_men_n688_), .B1(men_men_n565_), .Y(men_men_n1072_));
  NA4        u1044(.A(men_men_n1072_), .B(men_men_n1070_), .C(men_men_n1069_), .D(men_men_n1066_), .Y(men_men_n1073_));
  NO4        u1045(.A(men_men_n1073_), .B(men_men_n1065_), .C(men_men_n1059_), .D(men_men_n1042_), .Y(men_men_n1074_));
  NAi31      u1046(.An(men_men_n147_), .B(men_men_n448_), .C(n), .Y(men_men_n1075_));
  NO3        u1047(.A(men_men_n130_), .B(men_men_n363_), .C(men_men_n910_), .Y(men_men_n1076_));
  NO2        u1048(.A(men_men_n1076_), .B(men_men_n1075_), .Y(men_men_n1077_));
  NO3        u1049(.A(men_men_n287_), .B(men_men_n147_), .C(men_men_n435_), .Y(men_men_n1078_));
  AOI210     u1050(.A0(men_men_n1078_), .A1(men_men_n531_), .B0(men_men_n1077_), .Y(men_men_n1079_));
  INV        u1051(.A(men_men_n524_), .Y(men_men_n1080_));
  NA2        u1052(.A(men_men_n1080_), .B(men_men_n1079_), .Y(men_men_n1081_));
  NA2        u1053(.A(men_men_n242_), .B(men_men_n180_), .Y(men_men_n1082_));
  NO3        u1054(.A(men_men_n327_), .B(men_men_n472_), .C(men_men_n184_), .Y(men_men_n1083_));
  NOi31      u1055(.An(men_men_n1082_), .B(men_men_n1083_), .C(men_men_n225_), .Y(men_men_n1084_));
  NAi21      u1056(.An(men_men_n589_), .B(men_men_n1062_), .Y(men_men_n1085_));
  NA2        u1057(.A(men_men_n465_), .B(men_men_n941_), .Y(men_men_n1086_));
  NO3        u1058(.A(men_men_n466_), .B(men_men_n330_), .C(men_men_n75_), .Y(men_men_n1087_));
  AOI220     u1059(.A0(men_men_n1087_), .A1(men_men_n1086_), .B0(men_men_n514_), .B1(u), .Y(men_men_n1088_));
  NA2        u1060(.A(men_men_n1088_), .B(men_men_n1085_), .Y(men_men_n1089_));
  OAI220     u1061(.A0(men_men_n1075_), .A1(men_men_n245_), .B0(men_men_n1044_), .B1(men_men_n643_), .Y(men_men_n1090_));
  INV        u1062(.A(men_men_n705_), .Y(men_men_n1091_));
  NA2        u1063(.A(men_men_n1001_), .B(men_men_n992_), .Y(men_men_n1092_));
  NO3        u1064(.A(c), .B(men_men_n155_), .C(men_men_n224_), .Y(men_men_n1093_));
  OAI210     u1065(.A0(men_men_n1093_), .A1(men_men_n559_), .B0(men_men_n405_), .Y(men_men_n1094_));
  OAI220     u1066(.A0(men_men_n998_), .A1(men_men_n1006_), .B0(men_men_n579_), .B1(men_men_n456_), .Y(men_men_n1095_));
  NA4        u1067(.A(men_men_n1095_), .B(men_men_n1094_), .C(men_men_n1092_), .D(men_men_n662_), .Y(men_men_n1096_));
  OAI210     u1068(.A0(men_men_n1001_), .A1(men_men_n993_), .B0(men_men_n1082_), .Y(men_men_n1097_));
  NA3        u1069(.A(men_men_n1040_), .B(men_men_n519_), .C(men_men_n46_), .Y(men_men_n1098_));
  AOI210     u1070(.A0(men_men_n407_), .A1(men_men_n405_), .B0(men_men_n353_), .Y(men_men_n1099_));
  NA4        u1071(.A(men_men_n1099_), .B(men_men_n1098_), .C(men_men_n1097_), .D(men_men_n288_), .Y(men_men_n1100_));
  OR4        u1072(.A(men_men_n1100_), .B(men_men_n1096_), .C(men_men_n1091_), .D(men_men_n1090_), .Y(men_men_n1101_));
  NO4        u1073(.A(men_men_n1101_), .B(men_men_n1089_), .C(men_men_n1084_), .D(men_men_n1081_), .Y(men_men_n1102_));
  NA4        u1074(.A(men_men_n1102_), .B(men_men_n1074_), .C(men_men_n1032_), .D(men_men_n1017_), .Y(men13));
  NA2        u1075(.A(men_men_n46_), .B(men_men_n89_), .Y(men_men_n1104_));
  AN2        u1076(.A(c), .B(b), .Y(men_men_n1105_));
  NA3        u1077(.A(men_men_n263_), .B(men_men_n1105_), .C(m), .Y(men_men_n1106_));
  NO4        u1078(.A(e), .B(men_men_n1106_), .C(men_men_n1104_), .D(men_men_n621_), .Y(men_men_n1107_));
  NA2        u1079(.A(men_men_n279_), .B(men_men_n1105_), .Y(men_men_n1108_));
  NO4        u1080(.A(men_men_n1108_), .B(e), .C(men_men_n1034_), .D(a), .Y(men_men_n1109_));
  NAi32      u1081(.An(d), .Bn(c), .C(e), .Y(men_men_n1110_));
  NA2        u1082(.A(men_men_n146_), .B(men_men_n45_), .Y(men_men_n1111_));
  NO4        u1083(.A(men_men_n1111_), .B(men_men_n1110_), .C(men_men_n628_), .D(men_men_n326_), .Y(men_men_n1112_));
  NA2        u1084(.A(men_men_n712_), .B(men_men_n236_), .Y(men_men_n1113_));
  NA2        u1085(.A(men_men_n438_), .B(men_men_n224_), .Y(men_men_n1114_));
  AN2        u1086(.A(d), .B(c), .Y(men_men_n1115_));
  NA2        u1087(.A(men_men_n1115_), .B(men_men_n120_), .Y(men_men_n1116_));
  NO4        u1088(.A(men_men_n1116_), .B(men_men_n1114_), .C(men_men_n185_), .D(men_men_n176_), .Y(men_men_n1117_));
  NA2        u1089(.A(men_men_n529_), .B(c), .Y(men_men_n1118_));
  NO4        u1090(.A(men_men_n1111_), .B(men_men_n624_), .C(men_men_n1118_), .D(men_men_n326_), .Y(men_men_n1119_));
  AO210      u1091(.A0(men_men_n1117_), .A1(men_men_n1113_), .B0(men_men_n1119_), .Y(men_men_n1120_));
  OR4        u1092(.A(men_men_n1120_), .B(men_men_n1112_), .C(men_men_n1109_), .D(men_men_n1107_), .Y(men_men_n1121_));
  NAi32      u1093(.An(f), .Bn(e), .C(c), .Y(men_men_n1122_));
  NO2        u1094(.A(men_men_n1122_), .B(men_men_n152_), .Y(men_men_n1123_));
  NA2        u1095(.A(men_men_n1123_), .B(u), .Y(men_men_n1124_));
  OR3        u1096(.A(men_men_n236_), .B(men_men_n185_), .C(men_men_n176_), .Y(men_men_n1125_));
  NO2        u1097(.A(men_men_n1125_), .B(men_men_n1124_), .Y(men_men_n1126_));
  NO2        u1098(.A(men_men_n1118_), .B(men_men_n326_), .Y(men_men_n1127_));
  NO2        u1099(.A(j), .B(men_men_n45_), .Y(men_men_n1128_));
  NA2        u1100(.A(men_men_n672_), .B(men_men_n1128_), .Y(men_men_n1129_));
  NOi21      u1101(.An(men_men_n1127_), .B(men_men_n1129_), .Y(men_men_n1130_));
  NO2        u1102(.A(men_men_n815_), .B(men_men_n116_), .Y(men_men_n1131_));
  NOi41      u1103(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1132_));
  NA2        u1104(.A(men_men_n1132_), .B(men_men_n1131_), .Y(men_men_n1133_));
  NO2        u1105(.A(men_men_n1133_), .B(men_men_n1124_), .Y(men_men_n1134_));
  OR3        u1106(.A(e), .B(d), .C(c), .Y(men_men_n1135_));
  NA3        u1107(.A(k), .B(j), .C(i), .Y(men_men_n1136_));
  NO3        u1108(.A(men_men_n1136_), .B(men_men_n326_), .C(men_men_n93_), .Y(men_men_n1137_));
  NOi21      u1109(.An(men_men_n1137_), .B(men_men_n1135_), .Y(men_men_n1138_));
  OR4        u1110(.A(men_men_n1138_), .B(men_men_n1134_), .C(men_men_n1130_), .D(men_men_n1126_), .Y(men_men_n1139_));
  NA3        u1111(.A(men_men_n497_), .B(men_men_n356_), .C(men_men_n56_), .Y(men_men_n1140_));
  NO2        u1112(.A(men_men_n1140_), .B(men_men_n1129_), .Y(men_men_n1141_));
  NO4        u1113(.A(men_men_n1140_), .B(men_men_n624_), .C(men_men_n479_), .D(men_men_n45_), .Y(men_men_n1142_));
  NO2        u1114(.A(f), .B(c), .Y(men_men_n1143_));
  NOi21      u1115(.An(men_men_n1143_), .B(men_men_n471_), .Y(men_men_n1144_));
  NA2        u1116(.A(men_men_n1144_), .B(men_men_n59_), .Y(men_men_n1145_));
  OR2        u1117(.A(k), .B(i), .Y(men_men_n1146_));
  NO3        u1118(.A(men_men_n1146_), .B(men_men_n256_), .C(l), .Y(men_men_n1147_));
  NOi31      u1119(.An(men_men_n1147_), .B(men_men_n1145_), .C(j), .Y(men_men_n1148_));
  OR3        u1120(.A(men_men_n1148_), .B(men_men_n1142_), .C(men_men_n1141_), .Y(men_men_n1149_));
  OR3        u1121(.A(men_men_n1149_), .B(men_men_n1139_), .C(men_men_n1121_), .Y(men02));
  OR2        u1122(.A(l), .B(k), .Y(men_men_n1151_));
  OR3        u1123(.A(h), .B(u), .C(f), .Y(men_men_n1152_));
  OR3        u1124(.A(n), .B(m), .C(i), .Y(men_men_n1153_));
  NO4        u1125(.A(men_men_n1153_), .B(men_men_n1152_), .C(men_men_n1151_), .D(men_men_n1135_), .Y(men_men_n1154_));
  NOi31      u1126(.An(e), .B(d), .C(c), .Y(men_men_n1155_));
  AOI210     u1127(.A0(men_men_n1137_), .A1(men_men_n1155_), .B0(men_men_n1112_), .Y(men_men_n1156_));
  AN3        u1128(.A(u), .B(f), .C(c), .Y(men_men_n1157_));
  NA3        u1129(.A(men_men_n1157_), .B(men_men_n497_), .C(h), .Y(men_men_n1158_));
  OR2        u1130(.A(men_men_n1136_), .B(men_men_n326_), .Y(men_men_n1159_));
  OR2        u1131(.A(men_men_n1159_), .B(men_men_n1158_), .Y(men_men_n1160_));
  NO3        u1132(.A(men_men_n1140_), .B(men_men_n1111_), .C(men_men_n624_), .Y(men_men_n1161_));
  NO2        u1133(.A(men_men_n1161_), .B(men_men_n1126_), .Y(men_men_n1162_));
  NA3        u1134(.A(l), .B(k), .C(j), .Y(men_men_n1163_));
  NA2        u1135(.A(i), .B(h), .Y(men_men_n1164_));
  NO3        u1136(.A(men_men_n1164_), .B(men_men_n1163_), .C(men_men_n137_), .Y(men_men_n1165_));
  NO3        u1137(.A(men_men_n148_), .B(men_men_n300_), .C(men_men_n225_), .Y(men_men_n1166_));
  AOI210     u1138(.A0(men_men_n1166_), .A1(men_men_n1165_), .B0(men_men_n1130_), .Y(men_men_n1167_));
  NA3        u1139(.A(c), .B(b), .C(a), .Y(men_men_n1168_));
  NO3        u1140(.A(men_men_n1168_), .B(men_men_n964_), .C(men_men_n224_), .Y(men_men_n1169_));
  NO4        u1141(.A(men_men_n1136_), .B(men_men_n318_), .C(men_men_n49_), .D(men_men_n116_), .Y(men_men_n1170_));
  AOI210     u1142(.A0(men_men_n1170_), .A1(men_men_n1169_), .B0(men_men_n1141_), .Y(men_men_n1171_));
  AN4        u1143(.A(men_men_n1171_), .B(men_men_n1167_), .C(men_men_n1162_), .D(men_men_n1160_), .Y(men_men_n1172_));
  INV        u1144(.A(men_men_n1114_), .Y(men_men_n1173_));
  NA2        u1145(.A(men_men_n1133_), .B(men_men_n1125_), .Y(men_men_n1174_));
  AOI210     u1146(.A0(men_men_n1174_), .A1(men_men_n1173_), .B0(men_men_n1107_), .Y(men_men_n1175_));
  NAi41      u1147(.An(men_men_n1154_), .B(men_men_n1175_), .C(men_men_n1172_), .D(men_men_n1156_), .Y(men03));
  NO2        u1148(.A(men_men_n561_), .B(men_men_n637_), .Y(men_men_n1177_));
  NA4        u1149(.A(men_men_n90_), .B(men_men_n89_), .C(u), .D(men_men_n224_), .Y(men_men_n1178_));
  NA4        u1150(.A(men_men_n612_), .B(m), .C(men_men_n116_), .D(men_men_n224_), .Y(men_men_n1179_));
  NA3        u1151(.A(men_men_n1179_), .B(men_men_n395_), .C(men_men_n1178_), .Y(men_men_n1180_));
  NO3        u1152(.A(men_men_n1180_), .B(men_men_n1177_), .C(men_men_n1068_), .Y(men_men_n1181_));
  NOi41      u1153(.An(men_men_n863_), .B(men_men_n915_), .C(men_men_n904_), .D(men_men_n764_), .Y(men_men_n1182_));
  OAI220     u1154(.A0(men_men_n1182_), .A1(men_men_n738_), .B0(men_men_n1181_), .B1(men_men_n625_), .Y(men_men_n1183_));
  NOi31      u1155(.An(i), .B(k), .C(j), .Y(men_men_n1184_));
  NA4        u1156(.A(men_men_n1184_), .B(men_men_n1155_), .C(men_men_n365_), .D(men_men_n356_), .Y(men_men_n1185_));
  OAI210     u1157(.A0(men_men_n878_), .A1(men_men_n449_), .B0(men_men_n1185_), .Y(men_men_n1186_));
  NOi31      u1158(.An(m), .B(n), .C(f), .Y(men_men_n1187_));
  NA2        u1159(.A(men_men_n1187_), .B(men_men_n51_), .Y(men_men_n1188_));
  AN2        u1160(.A(e), .B(c), .Y(men_men_n1189_));
  NA2        u1161(.A(men_men_n1189_), .B(a), .Y(men_men_n1190_));
  OAI220     u1162(.A0(men_men_n1190_), .A1(men_men_n1188_), .B0(men_men_n947_), .B1(men_men_n455_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n540_), .B(l), .Y(men_men_n1192_));
  NOi31      u1164(.An(men_men_n926_), .B(men_men_n1106_), .C(men_men_n1192_), .Y(men_men_n1193_));
  NO4        u1165(.A(men_men_n1193_), .B(men_men_n1191_), .C(men_men_n1186_), .D(men_men_n1067_), .Y(men_men_n1194_));
  NO2        u1166(.A(men_men_n300_), .B(a), .Y(men_men_n1195_));
  INV        u1167(.A(men_men_n1112_), .Y(men_men_n1196_));
  NO2        u1168(.A(men_men_n1164_), .B(men_men_n517_), .Y(men_men_n1197_));
  NO2        u1169(.A(men_men_n89_), .B(u), .Y(men_men_n1198_));
  AOI210     u1170(.A0(men_men_n1198_), .A1(men_men_n1197_), .B0(men_men_n1147_), .Y(men_men_n1199_));
  OR2        u1171(.A(men_men_n1199_), .B(men_men_n1145_), .Y(men_men_n1200_));
  NA3        u1172(.A(men_men_n1200_), .B(men_men_n1196_), .C(men_men_n1194_), .Y(men_men_n1201_));
  NO4        u1173(.A(men_men_n1201_), .B(men_men_n1183_), .C(men_men_n880_), .D(men_men_n601_), .Y(men_men_n1202_));
  NA2        u1174(.A(c), .B(b), .Y(men_men_n1203_));
  OAI210     u1175(.A0(men_men_n924_), .A1(men_men_n895_), .B0(men_men_n442_), .Y(men_men_n1204_));
  OAI210     u1176(.A0(men_men_n1204_), .A1(men_men_n925_), .B0(men_men_n1668_), .Y(men_men_n1205_));
  NAi21      u1177(.An(men_men_n450_), .B(men_men_n1668_), .Y(men_men_n1206_));
  NA3        u1178(.A(men_men_n456_), .B(men_men_n594_), .C(f), .Y(men_men_n1207_));
  OAI210     u1179(.A0(men_men_n583_), .A1(men_men_n39_), .B0(men_men_n1195_), .Y(men_men_n1208_));
  NA3        u1180(.A(men_men_n1208_), .B(men_men_n1207_), .C(men_men_n1206_), .Y(men_men_n1209_));
  NA2        u1181(.A(men_men_n275_), .B(men_men_n123_), .Y(men_men_n1210_));
  OAI210     u1182(.A0(men_men_n1210_), .A1(men_men_n304_), .B0(u), .Y(men_men_n1211_));
  NAi21      u1183(.An(f), .B(d), .Y(men_men_n1212_));
  NO2        u1184(.A(men_men_n1212_), .B(men_men_n1168_), .Y(men_men_n1213_));
  INV        u1185(.A(men_men_n1213_), .Y(men_men_n1214_));
  AOI210     u1186(.A0(men_men_n1211_), .A1(men_men_n310_), .B0(men_men_n1214_), .Y(men_men_n1215_));
  AOI210     u1187(.A0(men_men_n1215_), .A1(men_men_n117_), .B0(men_men_n1209_), .Y(men_men_n1216_));
  NA2        u1188(.A(men_men_n500_), .B(men_men_n499_), .Y(men_men_n1217_));
  NO2        u1189(.A(men_men_n191_), .B(men_men_n249_), .Y(men_men_n1218_));
  NA2        u1190(.A(men_men_n1218_), .B(m), .Y(men_men_n1219_));
  NA3        u1191(.A(men_men_n981_), .B(men_men_n1192_), .C(men_men_n503_), .Y(men_men_n1220_));
  OAI210     u1192(.A0(men_men_n1220_), .A1(men_men_n331_), .B0(men_men_n501_), .Y(men_men_n1221_));
  AOI210     u1193(.A0(men_men_n1221_), .A1(men_men_n1217_), .B0(men_men_n1219_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n596_), .B(men_men_n437_), .Y(men_men_n1223_));
  NA2        u1195(.A(men_men_n165_), .B(men_men_n33_), .Y(men_men_n1224_));
  AOI210     u1196(.A0(men_men_n1030_), .A1(men_men_n1224_), .B0(men_men_n225_), .Y(men_men_n1225_));
  OAI210     u1197(.A0(men_men_n1225_), .A1(men_men_n475_), .B0(men_men_n1213_), .Y(men_men_n1226_));
  NO2        u1198(.A(men_men_n398_), .B(men_men_n397_), .Y(men_men_n1227_));
  AOI210     u1199(.A0(men_men_n1218_), .A1(men_men_n458_), .B0(men_men_n1025_), .Y(men_men_n1228_));
  NAi41      u1200(.An(men_men_n1227_), .B(men_men_n1228_), .C(men_men_n1226_), .D(men_men_n1223_), .Y(men_men_n1229_));
  NO2        u1201(.A(men_men_n1229_), .B(men_men_n1222_), .Y(men_men_n1230_));
  NA4        u1202(.A(men_men_n1230_), .B(men_men_n1216_), .C(men_men_n1205_), .D(men_men_n1202_), .Y(men00));
  AOI210     u1203(.A0(men_men_n317_), .A1(men_men_n225_), .B0(men_men_n292_), .Y(men_men_n1232_));
  NO2        u1204(.A(men_men_n1232_), .B(men_men_n615_), .Y(men_men_n1233_));
  AOI210     u1205(.A0(men_men_n961_), .A1(men_men_n1008_), .B0(men_men_n1186_), .Y(men_men_n1234_));
  NO3        u1206(.A(men_men_n1161_), .B(men_men_n1025_), .C(men_men_n761_), .Y(men_men_n1235_));
  NA3        u1207(.A(men_men_n1235_), .B(men_men_n1234_), .C(men_men_n1069_), .Y(men_men_n1236_));
  NA2        u1208(.A(men_men_n542_), .B(f), .Y(men_men_n1237_));
  OAI210     u1209(.A0(men_men_n1076_), .A1(men_men_n40_), .B0(men_men_n690_), .Y(men_men_n1238_));
  NA3        u1210(.A(men_men_n1238_), .B(men_men_n271_), .C(n), .Y(men_men_n1239_));
  AOI210     u1211(.A0(men_men_n1239_), .A1(men_men_n1237_), .B0(men_men_n1116_), .Y(men_men_n1240_));
  NO4        u1212(.A(men_men_n1240_), .B(men_men_n1236_), .C(men_men_n1233_), .D(men_men_n1139_), .Y(men_men_n1241_));
  NA3        u1213(.A(men_men_n175_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1242_));
  NA3        u1214(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1243_));
  NOi31      u1215(.An(n), .B(m), .C(i), .Y(men_men_n1244_));
  NA3        u1216(.A(men_men_n1244_), .B(men_men_n693_), .C(men_men_n51_), .Y(men_men_n1245_));
  OAI210     u1217(.A0(men_men_n1243_), .A1(men_men_n1242_), .B0(men_men_n1245_), .Y(men_men_n1246_));
  INV        u1218(.A(men_men_n614_), .Y(men_men_n1247_));
  NO4        u1219(.A(men_men_n1247_), .B(men_men_n1246_), .C(men_men_n1227_), .D(men_men_n984_), .Y(men_men_n1248_));
  NO4        u1220(.A(men_men_n520_), .B(men_men_n380_), .C(men_men_n1203_), .D(men_men_n59_), .Y(men_men_n1249_));
  NA3        u1221(.A(men_men_n410_), .B(men_men_n232_), .C(u), .Y(men_men_n1250_));
  OA220      u1222(.A0(men_men_n1250_), .A1(men_men_n1243_), .B0(men_men_n411_), .B1(men_men_n140_), .Y(men_men_n1251_));
  NO2        u1223(.A(h), .B(u), .Y(men_men_n1252_));
  NA4        u1224(.A(men_men_n531_), .B(men_men_n497_), .C(men_men_n1252_), .D(men_men_n1105_), .Y(men_men_n1253_));
  OAI220     u1225(.A0(men_men_n561_), .A1(men_men_n637_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1254_));
  AOI220     u1226(.A0(men_men_n1254_), .A1(men_men_n570_), .B0(men_men_n1013_), .B1(men_men_n613_), .Y(men_men_n1255_));
  AOI220     u1227(.A0(men_men_n338_), .A1(men_men_n260_), .B0(men_men_n186_), .B1(men_men_n154_), .Y(men_men_n1256_));
  NA4        u1228(.A(men_men_n1256_), .B(men_men_n1255_), .C(men_men_n1253_), .D(men_men_n1251_), .Y(men_men_n1257_));
  NO3        u1229(.A(men_men_n1257_), .B(men_men_n1249_), .C(men_men_n281_), .Y(men_men_n1258_));
  INV        u1230(.A(men_men_n343_), .Y(men_men_n1259_));
  AOI210     u1231(.A0(men_men_n260_), .A1(men_men_n370_), .B0(men_men_n616_), .Y(men_men_n1260_));
  NA3        u1232(.A(men_men_n1260_), .B(men_men_n1259_), .C(men_men_n160_), .Y(men_men_n1261_));
  NO2        u1233(.A(men_men_n251_), .B(men_men_n190_), .Y(men_men_n1262_));
  NA2        u1234(.A(men_men_n1262_), .B(men_men_n456_), .Y(men_men_n1263_));
  NA3        u1235(.A(men_men_n188_), .B(men_men_n116_), .C(u), .Y(men_men_n1264_));
  NA3        u1236(.A(men_men_n497_), .B(men_men_n40_), .C(f), .Y(men_men_n1265_));
  NOi31      u1237(.An(men_men_n934_), .B(men_men_n1265_), .C(men_men_n1264_), .Y(men_men_n1266_));
  NAi31      u1238(.An(men_men_n195_), .B(men_men_n921_), .C(men_men_n497_), .Y(men_men_n1267_));
  NAi31      u1239(.An(men_men_n1266_), .B(men_men_n1267_), .C(men_men_n1263_), .Y(men_men_n1268_));
  NO2        u1240(.A(men_men_n291_), .B(men_men_n75_), .Y(men_men_n1269_));
  NO3        u1241(.A(men_men_n455_), .B(men_men_n891_), .C(n), .Y(men_men_n1270_));
  AOI210     u1242(.A0(men_men_n1270_), .A1(men_men_n1269_), .B0(men_men_n1154_), .Y(men_men_n1271_));
  NAi31      u1243(.An(men_men_n1119_), .B(men_men_n1271_), .C(men_men_n74_), .Y(men_men_n1272_));
  NO4        u1244(.A(men_men_n1272_), .B(men_men_n1268_), .C(men_men_n1261_), .D(men_men_n552_), .Y(men_men_n1273_));
  AN3        u1245(.A(men_men_n1273_), .B(men_men_n1258_), .C(men_men_n1248_), .Y(men_men_n1274_));
  NA2        u1246(.A(men_men_n570_), .B(men_men_n104_), .Y(men_men_n1275_));
  NA3        u1247(.A(men_men_n1187_), .B(men_men_n648_), .C(men_men_n496_), .Y(men_men_n1276_));
  NA4        u1248(.A(men_men_n1276_), .B(men_men_n597_), .C(men_men_n1275_), .D(men_men_n254_), .Y(men_men_n1277_));
  NA2        u1249(.A(men_men_n1180_), .B(men_men_n570_), .Y(men_men_n1278_));
  NA4        u1250(.A(men_men_n693_), .B(men_men_n216_), .C(men_men_n232_), .D(men_men_n169_), .Y(men_men_n1279_));
  NA3        u1251(.A(men_men_n1279_), .B(men_men_n1278_), .C(men_men_n314_), .Y(men_men_n1280_));
  OAI210     u1252(.A0(men_men_n495_), .A1(men_men_n124_), .B0(men_men_n927_), .Y(men_men_n1281_));
  AOI220     u1253(.A0(men_men_n1281_), .A1(men_men_n1220_), .B0(men_men_n596_), .B1(men_men_n437_), .Y(men_men_n1282_));
  OR4        u1254(.A(men_men_n1116_), .B(men_men_n287_), .C(men_men_n234_), .D(e), .Y(men_men_n1283_));
  NO2        u1255(.A(men_men_n228_), .B(men_men_n225_), .Y(men_men_n1284_));
  NA2        u1256(.A(n), .B(e), .Y(men_men_n1285_));
  NO2        u1257(.A(men_men_n1285_), .B(men_men_n152_), .Y(men_men_n1286_));
  AOI220     u1258(.A0(men_men_n1286_), .A1(men_men_n289_), .B0(men_men_n908_), .B1(men_men_n1284_), .Y(men_men_n1287_));
  OAI210     u1259(.A0(men_men_n381_), .A1(men_men_n332_), .B0(men_men_n477_), .Y(men_men_n1288_));
  NA4        u1260(.A(men_men_n1288_), .B(men_men_n1287_), .C(men_men_n1283_), .D(men_men_n1282_), .Y(men_men_n1289_));
  AOI210     u1261(.A0(men_men_n1286_), .A1(men_men_n912_), .B0(men_men_n879_), .Y(men_men_n1290_));
  AOI220     u1262(.A0(men_men_n1021_), .A1(men_men_n613_), .B0(men_men_n693_), .B1(men_men_n257_), .Y(men_men_n1291_));
  NO2        u1263(.A(men_men_n68_), .B(h), .Y(men_men_n1292_));
  NO3        u1264(.A(men_men_n1116_), .B(men_men_n1114_), .C(men_men_n777_), .Y(men_men_n1293_));
  NO2        u1265(.A(men_men_n1151_), .B(men_men_n137_), .Y(men_men_n1294_));
  AN2        u1266(.A(men_men_n1294_), .B(men_men_n1166_), .Y(men_men_n1295_));
  OAI210     u1267(.A0(men_men_n1295_), .A1(men_men_n1293_), .B0(men_men_n1292_), .Y(men_men_n1296_));
  NA4        u1268(.A(men_men_n1296_), .B(men_men_n1291_), .C(men_men_n1290_), .D(men_men_n929_), .Y(men_men_n1297_));
  NO4        u1269(.A(men_men_n1297_), .B(men_men_n1289_), .C(men_men_n1280_), .D(men_men_n1277_), .Y(men_men_n1298_));
  NA2        u1270(.A(men_men_n896_), .B(men_men_n810_), .Y(men_men_n1299_));
  NA4        u1271(.A(men_men_n1299_), .B(men_men_n1298_), .C(men_men_n1274_), .D(men_men_n1241_), .Y(men01));
  AN2        u1272(.A(men_men_n1094_), .B(men_men_n1092_), .Y(men_men_n1301_));
  NO4        u1273(.A(men_men_n859_), .B(men_men_n851_), .C(men_men_n511_), .D(men_men_n298_), .Y(men_men_n1302_));
  NO2        u1274(.A(men_men_n630_), .B(men_men_n307_), .Y(men_men_n1303_));
  OAI210     u1275(.A0(men_men_n1303_), .A1(men_men_n421_), .B0(i), .Y(men_men_n1304_));
  NA3        u1276(.A(men_men_n1304_), .B(men_men_n1302_), .C(men_men_n1301_), .Y(men_men_n1305_));
  NA2        u1277(.A(men_men_n626_), .B(men_men_n92_), .Y(men_men_n1306_));
  NA2        u1278(.A(men_men_n589_), .B(men_men_n286_), .Y(men_men_n1307_));
  NA2        u1279(.A(men_men_n1028_), .B(men_men_n1307_), .Y(men_men_n1308_));
  NA4        u1280(.A(men_men_n1308_), .B(men_men_n1306_), .C(men_men_n977_), .D(men_men_n355_), .Y(men_men_n1309_));
  NA2        u1281(.A(men_men_n45_), .B(f), .Y(men_men_n1310_));
  NA2        u1282(.A(men_men_n756_), .B(men_men_n99_), .Y(men_men_n1311_));
  NO2        u1283(.A(men_men_n1311_), .B(men_men_n1310_), .Y(men_men_n1312_));
  OAI210     u1284(.A0(men_men_n837_), .A1(men_men_n643_), .B0(men_men_n1279_), .Y(men_men_n1313_));
  AOI210     u1285(.A0(men_men_n1312_), .A1(men_men_n679_), .B0(men_men_n1313_), .Y(men_men_n1314_));
  NA2        u1286(.A(men_men_n122_), .B(l), .Y(men_men_n1315_));
  OA220      u1287(.A0(men_men_n1315_), .A1(men_men_n623_), .B0(men_men_n706_), .B1(men_men_n395_), .Y(men_men_n1316_));
  NAi41      u1288(.An(men_men_n168_), .B(men_men_n1316_), .C(men_men_n1314_), .D(men_men_n960_), .Y(men_men_n1317_));
  NO3        u1289(.A(men_men_n838_), .B(men_men_n721_), .C(men_men_n545_), .Y(men_men_n1318_));
  NA4        u1290(.A(men_men_n756_), .B(men_men_n99_), .C(men_men_n45_), .D(men_men_n224_), .Y(men_men_n1319_));
  OA220      u1291(.A0(men_men_n1319_), .A1(men_men_n714_), .B0(men_men_n205_), .B1(men_men_n203_), .Y(men_men_n1320_));
  NA3        u1292(.A(men_men_n1320_), .B(men_men_n1318_), .C(men_men_n143_), .Y(men_men_n1321_));
  NO4        u1293(.A(men_men_n1321_), .B(men_men_n1317_), .C(men_men_n1309_), .D(men_men_n1305_), .Y(men_men_n1322_));
  NA2        u1294(.A(men_men_n1250_), .B(men_men_n217_), .Y(men_men_n1323_));
  OAI210     u1295(.A0(men_men_n1323_), .A1(men_men_n320_), .B0(men_men_n565_), .Y(men_men_n1324_));
  NA2        u1296(.A(men_men_n573_), .B(men_men_n423_), .Y(men_men_n1325_));
  NA2        u1297(.A(men_men_n76_), .B(i), .Y(men_men_n1326_));
  AOI210     u1298(.A0(men_men_n629_), .A1(men_men_n623_), .B0(men_men_n1326_), .Y(men_men_n1327_));
  NOi21      u1299(.An(men_men_n598_), .B(men_men_n620_), .Y(men_men_n1328_));
  AOI210     u1300(.A0(men_men_n1328_), .A1(men_men_n1325_), .B0(men_men_n1327_), .Y(men_men_n1329_));
  AOI210     u1301(.A0(men_men_n214_), .A1(men_men_n91_), .B0(men_men_n224_), .Y(men_men_n1330_));
  OAI210     u1302(.A0(men_men_n866_), .A1(men_men_n456_), .B0(men_men_n1330_), .Y(men_men_n1331_));
  AN3        u1303(.A(m), .B(l), .C(k), .Y(men_men_n1332_));
  OAI210     u1304(.A0(men_men_n383_), .A1(men_men_n34_), .B0(men_men_n1332_), .Y(men_men_n1333_));
  NA2        u1305(.A(men_men_n213_), .B(men_men_n34_), .Y(men_men_n1334_));
  AO210      u1306(.A0(men_men_n1334_), .A1(men_men_n1333_), .B0(men_men_n354_), .Y(men_men_n1335_));
  NA4        u1307(.A(men_men_n1335_), .B(men_men_n1331_), .C(men_men_n1329_), .D(men_men_n1324_), .Y(men_men_n1336_));
  AOI210     u1308(.A0(men_men_n635_), .A1(men_men_n122_), .B0(men_men_n641_), .Y(men_men_n1337_));
  OAI210     u1309(.A0(men_men_n1315_), .A1(men_men_n632_), .B0(men_men_n1337_), .Y(men_men_n1338_));
  NA2        u1310(.A(men_men_n297_), .B(men_men_n205_), .Y(men_men_n1339_));
  OAI210     u1311(.A0(men_men_n1339_), .A1(men_men_n412_), .B0(men_men_n711_), .Y(men_men_n1340_));
  NO3        u1312(.A(men_men_n878_), .B(men_men_n214_), .C(men_men_n435_), .Y(men_men_n1341_));
  NO2        u1313(.A(men_men_n1341_), .B(men_men_n1025_), .Y(men_men_n1342_));
  OAI210     u1314(.A0(men_men_n1312_), .A1(men_men_n348_), .B0(men_men_n722_), .Y(men_men_n1343_));
  NA4        u1315(.A(men_men_n1343_), .B(men_men_n1342_), .C(men_men_n1340_), .D(men_men_n841_), .Y(men_men_n1344_));
  NO3        u1316(.A(men_men_n1344_), .B(men_men_n1338_), .C(men_men_n1336_), .Y(men_men_n1345_));
  NA3        u1317(.A(men_men_n644_), .B(men_men_n29_), .C(f), .Y(men_men_n1346_));
  NO2        u1318(.A(men_men_n1346_), .B(men_men_n214_), .Y(men_men_n1347_));
  AOI210     u1319(.A0(men_men_n537_), .A1(men_men_n58_), .B0(men_men_n1347_), .Y(men_men_n1348_));
  OR3        u1320(.A(men_men_n1311_), .B(men_men_n645_), .C(men_men_n1310_), .Y(men_men_n1349_));
  NA3        u1321(.A(men_men_n791_), .B(men_men_n76_), .C(i), .Y(men_men_n1350_));
  AOI210     u1322(.A0(men_men_n1350_), .A1(men_men_n1319_), .B0(men_men_n1047_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n217_), .B(men_men_n115_), .Y(men_men_n1352_));
  NO3        u1324(.A(men_men_n1352_), .B(men_men_n1351_), .C(men_men_n1246_), .Y(men_men_n1353_));
  NA4        u1325(.A(men_men_n1353_), .B(men_men_n1349_), .C(men_men_n1348_), .D(men_men_n809_), .Y(men_men_n1354_));
  NO2        u1326(.A(men_men_n1034_), .B(men_men_n244_), .Y(men_men_n1355_));
  NO2        u1327(.A(men_men_n1035_), .B(men_men_n591_), .Y(men_men_n1356_));
  OAI210     u1328(.A0(men_men_n1356_), .A1(men_men_n1355_), .B0(men_men_n363_), .Y(men_men_n1357_));
  NA2        u1329(.A(men_men_n608_), .B(men_men_n606_), .Y(men_men_n1358_));
  NO3        u1330(.A(men_men_n81_), .B(men_men_n318_), .C(men_men_n45_), .Y(men_men_n1359_));
  NA2        u1331(.A(men_men_n1359_), .B(men_men_n588_), .Y(men_men_n1360_));
  NA3        u1332(.A(men_men_n1360_), .B(men_men_n1358_), .C(men_men_n716_), .Y(men_men_n1361_));
  OR2        u1333(.A(men_men_n1250_), .B(men_men_n1243_), .Y(men_men_n1362_));
  NO2        u1334(.A(men_men_n395_), .B(men_men_n73_), .Y(men_men_n1363_));
  AOI210     u1335(.A0(men_men_n782_), .A1(men_men_n659_), .B0(men_men_n1363_), .Y(men_men_n1364_));
  NA2        u1336(.A(men_men_n1359_), .B(men_men_n869_), .Y(men_men_n1365_));
  NA4        u1337(.A(men_men_n1365_), .B(men_men_n1364_), .C(men_men_n1362_), .D(men_men_n413_), .Y(men_men_n1366_));
  NOi41      u1338(.An(men_men_n1357_), .B(men_men_n1366_), .C(men_men_n1361_), .D(men_men_n1354_), .Y(men_men_n1367_));
  NO2        u1339(.A(men_men_n136_), .B(men_men_n45_), .Y(men_men_n1368_));
  AO220      u1340(.A0(i), .A1(men_men_n665_), .B0(men_men_n1368_), .B1(men_men_n754_), .Y(men_men_n1369_));
  NA2        u1341(.A(men_men_n1369_), .B(men_men_n363_), .Y(men_men_n1370_));
  NA2        u1342(.A(men_men_n490_), .B(men_men_n140_), .Y(men_men_n1371_));
  NO3        u1343(.A(men_men_n1164_), .B(men_men_n185_), .C(men_men_n89_), .Y(men_men_n1372_));
  AOI220     u1344(.A0(men_men_n1372_), .A1(men_men_n1371_), .B0(men_men_n1359_), .B1(men_men_n1038_), .Y(men_men_n1373_));
  NA2        u1345(.A(men_men_n1373_), .B(men_men_n1370_), .Y(men_men_n1374_));
  NO2        u1346(.A(men_men_n656_), .B(men_men_n655_), .Y(men_men_n1375_));
  NO4        u1347(.A(men_men_n1164_), .B(men_men_n1375_), .C(men_men_n183_), .D(men_men_n89_), .Y(men_men_n1376_));
  NO3        u1348(.A(men_men_n1376_), .B(men_men_n1374_), .C(men_men_n683_), .Y(men_men_n1377_));
  NA4        u1349(.A(men_men_n1377_), .B(men_men_n1367_), .C(men_men_n1345_), .D(men_men_n1322_), .Y(men06));
  NO2        u1350(.A(men_men_n436_), .B(men_men_n595_), .Y(men_men_n1379_));
  NO2        u1351(.A(men_men_n784_), .B(i), .Y(men_men_n1380_));
  OAI210     u1352(.A0(men_men_n1380_), .A1(men_men_n282_), .B0(men_men_n1379_), .Y(men_men_n1381_));
  NO2        u1353(.A(men_men_n236_), .B(men_men_n106_), .Y(men_men_n1382_));
  OAI210     u1354(.A0(men_men_n1382_), .A1(men_men_n1372_), .B0(men_men_n409_), .Y(men_men_n1383_));
  NO3        u1355(.A(men_men_n639_), .B(men_men_n864_), .C(men_men_n642_), .Y(men_men_n1384_));
  OR2        u1356(.A(men_men_n1384_), .B(men_men_n947_), .Y(men_men_n1385_));
  NA4        u1357(.A(men_men_n1385_), .B(men_men_n1383_), .C(men_men_n1381_), .D(men_men_n1357_), .Y(men_men_n1386_));
  NO3        u1358(.A(men_men_n1386_), .B(men_men_n1361_), .C(men_men_n270_), .Y(men_men_n1387_));
  NO2        u1359(.A(men_men_n318_), .B(men_men_n45_), .Y(men_men_n1388_));
  AOI210     u1360(.A0(men_men_n1388_), .A1(men_men_n1039_), .B0(men_men_n1355_), .Y(men_men_n1389_));
  AOI210     u1361(.A0(men_men_n1388_), .A1(men_men_n592_), .B0(men_men_n1369_), .Y(men_men_n1390_));
  AOI210     u1362(.A0(men_men_n1390_), .A1(men_men_n1389_), .B0(men_men_n360_), .Y(men_men_n1391_));
  OAI210     u1363(.A0(men_men_n91_), .A1(men_men_n40_), .B0(men_men_n720_), .Y(men_men_n1392_));
  NA2        u1364(.A(men_men_n1392_), .B(men_men_n386_), .Y(men_men_n1393_));
  NO2        u1365(.A(men_men_n548_), .B(men_men_n180_), .Y(men_men_n1394_));
  NOi21      u1366(.An(men_men_n142_), .B(men_men_n45_), .Y(men_men_n1395_));
  NO2        u1367(.A(men_men_n649_), .B(men_men_n1188_), .Y(men_men_n1396_));
  OAI210     u1368(.A0(men_men_n490_), .A1(men_men_n261_), .B0(men_men_n971_), .Y(men_men_n1397_));
  NO4        u1369(.A(men_men_n1397_), .B(men_men_n1396_), .C(men_men_n1395_), .D(men_men_n1394_), .Y(men_men_n1398_));
  OR2        u1370(.A(men_men_n640_), .B(men_men_n638_), .Y(men_men_n1399_));
  NO2        u1371(.A(men_men_n394_), .B(men_men_n141_), .Y(men_men_n1400_));
  AOI210     u1372(.A0(men_men_n1400_), .A1(men_men_n626_), .B0(men_men_n1399_), .Y(men_men_n1401_));
  NA3        u1373(.A(men_men_n1401_), .B(men_men_n1398_), .C(men_men_n1393_), .Y(men_men_n1402_));
  NO2        u1374(.A(men_men_n800_), .B(men_men_n393_), .Y(men_men_n1403_));
  NO3        u1375(.A(men_men_n722_), .B(men_men_n811_), .C(men_men_n679_), .Y(men_men_n1404_));
  NOi21      u1376(.An(men_men_n1403_), .B(men_men_n1404_), .Y(men_men_n1405_));
  AN2        u1377(.A(men_men_n1021_), .B(men_men_n689_), .Y(men_men_n1406_));
  NO4        u1378(.A(men_men_n1406_), .B(men_men_n1405_), .C(men_men_n1402_), .D(men_men_n1391_), .Y(men_men_n1407_));
  NO2        u1379(.A(men_men_n858_), .B(men_men_n293_), .Y(men_men_n1408_));
  OAI220     u1380(.A0(men_men_n784_), .A1(men_men_n47_), .B0(men_men_n236_), .B1(men_men_n658_), .Y(men_men_n1409_));
  OAI210     u1381(.A0(men_men_n293_), .A1(c), .B0(men_men_n686_), .Y(men_men_n1410_));
  AOI220     u1382(.A0(men_men_n1410_), .A1(men_men_n1409_), .B0(men_men_n1408_), .B1(men_men_n282_), .Y(men_men_n1411_));
  NO3        u1383(.A(men_men_n256_), .B(men_men_n106_), .C(men_men_n300_), .Y(men_men_n1412_));
  OAI220     u1384(.A0(men_men_n747_), .A1(men_men_n261_), .B0(men_men_n544_), .B1(men_men_n548_), .Y(men_men_n1413_));
  OAI210     u1385(.A0(l), .A1(i), .B0(k), .Y(men_men_n1414_));
  NO3        u1386(.A(men_men_n1414_), .B(men_men_n637_), .C(j), .Y(men_men_n1415_));
  NOi21      u1387(.An(men_men_n1415_), .B(men_men_n714_), .Y(men_men_n1416_));
  NO4        u1388(.A(men_men_n1416_), .B(men_men_n1413_), .C(men_men_n1412_), .D(men_men_n1191_), .Y(men_men_n1417_));
  NA4        u1389(.A(men_men_n849_), .B(men_men_n848_), .C(men_men_n465_), .D(men_men_n941_), .Y(men_men_n1418_));
  NAi31      u1390(.An(men_men_n800_), .B(men_men_n1418_), .C(men_men_n213_), .Y(men_men_n1419_));
  NA4        u1391(.A(men_men_n1419_), .B(men_men_n1417_), .C(men_men_n1411_), .D(men_men_n1291_), .Y(men_men_n1420_));
  NOi31      u1392(.An(men_men_n1384_), .B(men_men_n494_), .C(men_men_n422_), .Y(men_men_n1421_));
  OR3        u1393(.A(men_men_n1421_), .B(men_men_n837_), .C(men_men_n576_), .Y(men_men_n1422_));
  OR3        u1394(.A(men_men_n397_), .B(men_men_n236_), .C(men_men_n658_), .Y(men_men_n1423_));
  AOI210     u1395(.A0(men_men_n608_), .A1(men_men_n477_), .B0(men_men_n399_), .Y(men_men_n1424_));
  NA2        u1396(.A(men_men_n1415_), .B(men_men_n845_), .Y(men_men_n1425_));
  NA4        u1397(.A(men_men_n1425_), .B(men_men_n1424_), .C(men_men_n1423_), .D(men_men_n1422_), .Y(men_men_n1426_));
  AOI220     u1398(.A0(men_men_n1403_), .A1(men_men_n810_), .B0(men_men_n1400_), .B1(men_men_n250_), .Y(men_men_n1427_));
  AO220      u1399(.A0(men_men_n1382_), .A1(men_men_n711_), .B0(men_men_n993_), .B1(men_men_n992_), .Y(men_men_n1428_));
  NO4        u1400(.A(men_men_n1428_), .B(men_men_n939_), .C(men_men_n533_), .D(men_men_n514_), .Y(men_men_n1429_));
  NA3        u1401(.A(men_men_n1429_), .B(men_men_n1427_), .C(men_men_n1365_), .Y(men_men_n1430_));
  NAi21      u1402(.An(j), .B(i), .Y(men_men_n1431_));
  NO4        u1403(.A(men_men_n1375_), .B(men_men_n1431_), .C(men_men_n471_), .D(men_men_n247_), .Y(men_men_n1432_));
  NO4        u1404(.A(men_men_n1432_), .B(men_men_n1430_), .C(men_men_n1426_), .D(men_men_n1420_), .Y(men_men_n1433_));
  NA4        u1405(.A(men_men_n1433_), .B(men_men_n1407_), .C(men_men_n1387_), .D(men_men_n1377_), .Y(men07));
  NOi21      u1406(.An(j), .B(k), .Y(men_men_n1435_));
  NA4        u1407(.A(men_men_n188_), .B(men_men_n112_), .C(men_men_n1435_), .D(f), .Y(men_men_n1436_));
  NAi32      u1408(.An(m), .Bn(b), .C(n), .Y(men_men_n1437_));
  NO3        u1409(.A(men_men_n1437_), .B(u), .C(f), .Y(men_men_n1438_));
  OAI210     u1410(.A0(men_men_n342_), .A1(men_men_n516_), .B0(men_men_n1438_), .Y(men_men_n1439_));
  NAi21      u1411(.An(f), .B(c), .Y(men_men_n1440_));
  OR2        u1412(.A(e), .B(d), .Y(men_men_n1441_));
  OAI220     u1413(.A0(men_men_n1441_), .A1(men_men_n1440_), .B0(men_men_n671_), .B1(men_men_n344_), .Y(men_men_n1442_));
  NA3        u1414(.A(men_men_n1442_), .B(men_men_n1128_), .C(men_men_n188_), .Y(men_men_n1443_));
  NOi31      u1415(.An(n), .B(m), .C(b), .Y(men_men_n1444_));
  NO3        u1416(.A(men_men_n137_), .B(men_men_n479_), .C(h), .Y(men_men_n1445_));
  NA3        u1417(.A(men_men_n1443_), .B(men_men_n1439_), .C(men_men_n1436_), .Y(men_men_n1446_));
  NOi41      u1418(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1447_));
  NA3        u1419(.A(men_men_n1447_), .B(men_men_n931_), .C(men_men_n438_), .Y(men_men_n1448_));
  NOi21      u1420(.An(h), .B(k), .Y(men_men_n1449_));
  NO2        u1421(.A(men_men_n1448_), .B(men_men_n56_), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1166_), .B(men_men_n232_), .Y(men_men_n1451_));
  NO2        u1423(.A(men_men_n1451_), .B(men_men_n61_), .Y(men_men_n1452_));
  NO2        u1424(.A(k), .B(i), .Y(men_men_n1453_));
  NA3        u1425(.A(men_men_n1453_), .B(men_men_n959_), .C(men_men_n188_), .Y(men_men_n1454_));
  NA2        u1426(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1455_));
  NO2        u1427(.A(men_men_n1122_), .B(men_men_n471_), .Y(men_men_n1456_));
  NA3        u1428(.A(men_men_n1456_), .B(men_men_n1455_), .C(men_men_n225_), .Y(men_men_n1457_));
  NO2        u1429(.A(men_men_n1136_), .B(men_men_n326_), .Y(men_men_n1458_));
  NA2        u1430(.A(men_men_n577_), .B(men_men_n82_), .Y(men_men_n1459_));
  NA2        u1431(.A(men_men_n1292_), .B(men_men_n308_), .Y(men_men_n1460_));
  NA4        u1432(.A(men_men_n1460_), .B(men_men_n1459_), .C(men_men_n1457_), .D(men_men_n1454_), .Y(men_men_n1461_));
  NO4        u1433(.A(men_men_n1461_), .B(men_men_n1452_), .C(men_men_n1450_), .D(men_men_n1446_), .Y(men_men_n1462_));
  NO3        u1434(.A(e), .B(d), .C(c), .Y(men_men_n1463_));
  OAI210     u1435(.A0(men_men_n137_), .A1(men_men_n225_), .B0(men_men_n646_), .Y(men_men_n1464_));
  NA2        u1436(.A(men_men_n1464_), .B(men_men_n1463_), .Y(men_men_n1465_));
  INV        u1437(.A(men_men_n1465_), .Y(men_men_n1466_));
  OR2        u1438(.A(h), .B(f), .Y(men_men_n1467_));
  NO3        u1439(.A(n), .B(m), .C(i), .Y(men_men_n1468_));
  OAI210     u1440(.A0(men_men_n1189_), .A1(men_men_n163_), .B0(men_men_n1468_), .Y(men_men_n1469_));
  NO2        u1441(.A(i), .B(u), .Y(men_men_n1470_));
  OR3        u1442(.A(men_men_n1470_), .B(men_men_n1437_), .C(men_men_n72_), .Y(men_men_n1471_));
  OAI220     u1443(.A0(men_men_n1471_), .A1(men_men_n516_), .B0(men_men_n1469_), .B1(men_men_n1467_), .Y(men_men_n1472_));
  NA3        u1444(.A(men_men_n744_), .B(men_men_n730_), .C(men_men_n116_), .Y(men_men_n1473_));
  NA3        u1445(.A(men_men_n1444_), .B(men_men_n1131_), .C(men_men_n718_), .Y(men_men_n1474_));
  AOI210     u1446(.A0(men_men_n1474_), .A1(men_men_n1473_), .B0(men_men_n45_), .Y(men_men_n1475_));
  NA2        u1447(.A(men_men_n1468_), .B(men_men_n685_), .Y(men_men_n1476_));
  NO2        u1448(.A(l), .B(k), .Y(men_men_n1477_));
  NOi41      u1449(.An(men_men_n581_), .B(men_men_n1477_), .C(men_men_n509_), .D(men_men_n471_), .Y(men_men_n1478_));
  NO3        u1450(.A(men_men_n471_), .B(d), .C(c), .Y(men_men_n1479_));
  NO4        u1451(.A(men_men_n1478_), .B(men_men_n1475_), .C(men_men_n1472_), .D(men_men_n1466_), .Y(men_men_n1480_));
  NO2        u1452(.A(men_men_n153_), .B(h), .Y(men_men_n1481_));
  NO2        u1453(.A(u), .B(c), .Y(men_men_n1482_));
  NA3        u1454(.A(men_men_n1482_), .B(men_men_n148_), .C(men_men_n196_), .Y(men_men_n1483_));
  NO2        u1455(.A(men_men_n1483_), .B(men_men_n1665_), .Y(men_men_n1484_));
  NA2        u1456(.A(men_men_n1484_), .B(men_men_n188_), .Y(men_men_n1485_));
  OAI210     u1457(.A0(men_men_n1449_), .A1(men_men_n224_), .B0(men_men_n1146_), .Y(men_men_n1486_));
  NO2        u1458(.A(men_men_n482_), .B(a), .Y(men_men_n1487_));
  NA3        u1459(.A(men_men_n1487_), .B(men_men_n1486_), .C(men_men_n117_), .Y(men_men_n1488_));
  NO2        u1460(.A(i), .B(h), .Y(men_men_n1489_));
  NA2        u1461(.A(men_men_n1489_), .B(men_men_n232_), .Y(men_men_n1490_));
  AOI210     u1462(.A0(men_men_n1212_), .A1(h), .B0(men_men_n443_), .Y(men_men_n1491_));
  NA2        u1463(.A(men_men_n144_), .B(men_men_n232_), .Y(men_men_n1492_));
  AOI210     u1464(.A0(men_men_n271_), .A1(men_men_n120_), .B0(men_men_n565_), .Y(men_men_n1493_));
  OAI220     u1465(.A0(men_men_n1493_), .A1(men_men_n1490_), .B0(men_men_n1492_), .B1(men_men_n1491_), .Y(men_men_n1494_));
  NO2        u1466(.A(men_men_n807_), .B(men_men_n197_), .Y(men_men_n1495_));
  NOi31      u1467(.An(m), .B(n), .C(b), .Y(men_men_n1496_));
  NOi31      u1468(.An(f), .B(d), .C(c), .Y(men_men_n1497_));
  NA2        u1469(.A(men_men_n1497_), .B(men_men_n1496_), .Y(men_men_n1498_));
  INV        u1470(.A(men_men_n1498_), .Y(men_men_n1499_));
  NO3        u1471(.A(men_men_n1499_), .B(men_men_n1495_), .C(men_men_n1494_), .Y(men_men_n1500_));
  NA2        u1472(.A(men_men_n1157_), .B(men_men_n497_), .Y(men_men_n1501_));
  NO4        u1473(.A(men_men_n1501_), .B(men_men_n1131_), .C(men_men_n471_), .D(men_men_n45_), .Y(men_men_n1502_));
  NO3        u1474(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1503_));
  INV        u1475(.A(men_men_n1502_), .Y(men_men_n1504_));
  AN4        u1476(.A(men_men_n1504_), .B(men_men_n1500_), .C(men_men_n1488_), .D(men_men_n1485_), .Y(men_men_n1505_));
  NA2        u1477(.A(men_men_n1444_), .B(men_men_n406_), .Y(men_men_n1506_));
  NO2        u1478(.A(men_men_n1506_), .B(men_men_n1113_), .Y(men_men_n1507_));
  NA2        u1479(.A(men_men_n1479_), .B(men_men_n226_), .Y(men_men_n1508_));
  NO2        u1480(.A(men_men_n197_), .B(b), .Y(men_men_n1509_));
  AOI220     u1481(.A0(men_men_n1244_), .A1(men_men_n1509_), .B0(men_men_n1165_), .B1(men_men_n1501_), .Y(men_men_n1510_));
  NO2        u1482(.A(i), .B(men_men_n224_), .Y(men_men_n1511_));
  NA4        u1483(.A(men_men_n1218_), .B(men_men_n1511_), .C(men_men_n107_), .D(m), .Y(men_men_n1512_));
  NAi41      u1484(.An(men_men_n1507_), .B(men_men_n1512_), .C(men_men_n1510_), .D(men_men_n1508_), .Y(men_men_n1513_));
  NO4        u1485(.A(men_men_n137_), .B(u), .C(f), .D(e), .Y(men_men_n1514_));
  NA3        u1486(.A(men_men_n1453_), .B(men_men_n309_), .C(h), .Y(men_men_n1515_));
  NA2        u1487(.A(men_men_n204_), .B(men_men_n101_), .Y(men_men_n1516_));
  OR2        u1488(.A(e), .B(a), .Y(men_men_n1517_));
  NO2        u1489(.A(men_men_n1441_), .B(men_men_n1440_), .Y(men_men_n1518_));
  AOI210     u1490(.A0(men_men_n30_), .A1(h), .B0(men_men_n1518_), .Y(men_men_n1519_));
  NO2        u1491(.A(men_men_n1519_), .B(men_men_n1153_), .Y(men_men_n1520_));
  NOi41      u1492(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1521_));
  NA2        u1493(.A(men_men_n1521_), .B(men_men_n117_), .Y(men_men_n1522_));
  NA2        u1494(.A(men_men_n1447_), .B(men_men_n1477_), .Y(men_men_n1523_));
  NA2        u1495(.A(men_men_n1523_), .B(men_men_n1522_), .Y(men_men_n1524_));
  OR3        u1496(.A(men_men_n576_), .B(men_men_n575_), .C(men_men_n116_), .Y(men_men_n1525_));
  NA2        u1497(.A(men_men_n1187_), .B(men_men_n435_), .Y(men_men_n1526_));
  OAI220     u1498(.A0(men_men_n1526_), .A1(men_men_n464_), .B0(men_men_n1525_), .B1(men_men_n318_), .Y(men_men_n1527_));
  AO210      u1499(.A0(men_men_n1527_), .A1(men_men_n120_), .B0(men_men_n1524_), .Y(men_men_n1528_));
  NO3        u1500(.A(men_men_n1528_), .B(men_men_n1520_), .C(men_men_n1513_), .Y(men_men_n1529_));
  NA4        u1501(.A(men_men_n1529_), .B(men_men_n1505_), .C(men_men_n1480_), .D(men_men_n1462_), .Y(men_men_n1530_));
  NO2        u1502(.A(men_men_n1203_), .B(men_men_n114_), .Y(men_men_n1531_));
  NA2        u1503(.A(men_men_n406_), .B(men_men_n56_), .Y(men_men_n1532_));
  AOI210     u1504(.A0(men_men_n1532_), .A1(men_men_n1122_), .B0(men_men_n1476_), .Y(men_men_n1533_));
  NA2        u1505(.A(men_men_n226_), .B(men_men_n188_), .Y(men_men_n1534_));
  AOI210     u1506(.A0(men_men_n1534_), .A1(men_men_n1264_), .B0(men_men_n1532_), .Y(men_men_n1535_));
  NO2        u1507(.A(men_men_n1158_), .B(men_men_n1153_), .Y(men_men_n1536_));
  NO3        u1508(.A(men_men_n1536_), .B(men_men_n1535_), .C(men_men_n1533_), .Y(men_men_n1537_));
  NO2        u1509(.A(men_men_n418_), .B(j), .Y(men_men_n1538_));
  NA3        u1510(.A(men_men_n1503_), .B(men_men_n1441_), .C(men_men_n1187_), .Y(men_men_n1539_));
  NAi41      u1511(.An(men_men_n1489_), .B(men_men_n1144_), .C(men_men_n176_), .D(men_men_n156_), .Y(men_men_n1540_));
  NA2        u1512(.A(men_men_n1540_), .B(men_men_n1539_), .Y(men_men_n1541_));
  NA3        u1513(.A(u), .B(men_men_n1538_), .C(men_men_n165_), .Y(men_men_n1542_));
  INV        u1514(.A(men_men_n1542_), .Y(men_men_n1543_));
  NO3        u1515(.A(men_men_n800_), .B(men_men_n183_), .C(men_men_n438_), .Y(men_men_n1544_));
  NO3        u1516(.A(men_men_n1544_), .B(men_men_n1543_), .C(men_men_n1541_), .Y(men_men_n1545_));
  NO3        u1517(.A(men_men_n1153_), .B(men_men_n620_), .C(u), .Y(men_men_n1546_));
  NOi21      u1518(.An(men_men_n1534_), .B(men_men_n1546_), .Y(men_men_n1547_));
  AOI210     u1519(.A0(men_men_n1547_), .A1(men_men_n1516_), .B0(men_men_n1122_), .Y(men_men_n1548_));
  NA2        u1520(.A(men_men_n883_), .B(men_men_n204_), .Y(men_men_n1549_));
  INV        u1521(.A(men_men_n1549_), .Y(men_men_n1550_));
  OAI220     u1522(.A0(men_men_n712_), .A1(u), .B0(men_men_n236_), .B1(c), .Y(men_men_n1551_));
  AOI210     u1523(.A0(men_men_n1509_), .A1(men_men_n41_), .B0(men_men_n1551_), .Y(men_men_n1552_));
  NO2        u1524(.A(men_men_n137_), .B(l), .Y(men_men_n1553_));
  NO2        u1525(.A(men_men_n236_), .B(k), .Y(men_men_n1554_));
  OAI210     u1526(.A0(men_men_n1554_), .A1(men_men_n1489_), .B0(men_men_n1553_), .Y(men_men_n1555_));
  OAI220     u1527(.A0(men_men_n1555_), .A1(men_men_n31_), .B0(men_men_n1552_), .B1(men_men_n185_), .Y(men_men_n1556_));
  NO3        u1528(.A(men_men_n1525_), .B(men_men_n497_), .C(men_men_n377_), .Y(men_men_n1557_));
  NO4        u1529(.A(men_men_n1557_), .B(men_men_n1556_), .C(men_men_n1550_), .D(men_men_n1548_), .Y(men_men_n1558_));
  NO2        u1530(.A(men_men_n49_), .B(men_men_n620_), .Y(men_men_n1559_));
  NO3        u1531(.A(men_men_n1168_), .B(men_men_n1441_), .C(men_men_n49_), .Y(men_men_n1560_));
  AOI220     u1532(.A0(men_men_n1560_), .A1(men_men_n225_), .B0(men_men_n1169_), .B1(men_men_n1559_), .Y(men_men_n1561_));
  NO2        u1533(.A(men_men_n1153_), .B(h), .Y(men_men_n1562_));
  NA3        u1534(.A(men_men_n1562_), .B(d), .C(men_men_n1114_), .Y(men_men_n1563_));
  OAI220     u1535(.A0(men_men_n1563_), .A1(c), .B0(men_men_n1561_), .B1(j), .Y(men_men_n1564_));
  NA3        u1536(.A(men_men_n1531_), .B(men_men_n497_), .C(f), .Y(men_men_n1565_));
  NA2        u1537(.A(men_men_n188_), .B(men_men_n116_), .Y(men_men_n1566_));
  NO2        u1538(.A(men_men_n1435_), .B(men_men_n42_), .Y(men_men_n1567_));
  AOI210     u1539(.A0(men_men_n117_), .A1(men_men_n40_), .B0(men_men_n1567_), .Y(men_men_n1568_));
  NO2        u1540(.A(men_men_n1568_), .B(men_men_n1565_), .Y(men_men_n1569_));
  AOI210     u1541(.A0(men_men_n560_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1570_));
  NA2        u1542(.A(men_men_n1570_), .B(men_men_n1487_), .Y(men_men_n1571_));
  NO2        u1543(.A(men_men_n1431_), .B(men_men_n183_), .Y(men_men_n1572_));
  NOi21      u1544(.An(d), .B(f), .Y(men_men_n1573_));
  NO3        u1545(.A(men_men_n1497_), .B(men_men_n1573_), .C(men_men_n40_), .Y(men_men_n1574_));
  NA2        u1546(.A(men_men_n1574_), .B(men_men_n1572_), .Y(men_men_n1575_));
  NO2        u1547(.A(men_men_n1441_), .B(f), .Y(men_men_n1576_));
  NA2        u1548(.A(men_men_n1487_), .B(men_men_n1567_), .Y(men_men_n1577_));
  NO2        u1549(.A(men_men_n318_), .B(c), .Y(men_men_n1578_));
  NA2        u1550(.A(men_men_n1578_), .B(men_men_n577_), .Y(men_men_n1579_));
  NA4        u1551(.A(men_men_n1579_), .B(men_men_n1577_), .C(men_men_n1575_), .D(men_men_n1571_), .Y(men_men_n1580_));
  NO3        u1552(.A(men_men_n1580_), .B(men_men_n1569_), .C(men_men_n1564_), .Y(men_men_n1581_));
  NA4        u1553(.A(men_men_n1581_), .B(men_men_n1558_), .C(men_men_n1545_), .D(men_men_n1537_), .Y(men_men_n1582_));
  NO3        u1554(.A(men_men_n1157_), .B(men_men_n1143_), .C(men_men_n40_), .Y(men_men_n1583_));
  OAI220     u1555(.A0(men_men_n497_), .A1(men_men_n318_), .B0(men_men_n136_), .B1(men_men_n59_), .Y(men_men_n1584_));
  OAI210     u1556(.A0(men_men_n1584_), .A1(men_men_n1583_), .B0(men_men_n1458_), .Y(men_men_n1585_));
  NA2        u1557(.A(men_men_n1514_), .B(b), .Y(men_men_n1586_));
  NO2        u1558(.A(men_men_n1110_), .B(men_men_n137_), .Y(men_men_n1587_));
  NA2        u1559(.A(men_men_n1587_), .B(men_men_n664_), .Y(men_men_n1588_));
  NA3        u1560(.A(men_men_n1588_), .B(men_men_n1586_), .C(men_men_n1585_), .Y(men_men_n1589_));
  NA2        u1561(.A(men_men_n1482_), .B(men_men_n1573_), .Y(men_men_n1590_));
  NO2        u1562(.A(men_men_n1590_), .B(m), .Y(men_men_n1591_));
  NA3        u1563(.A(men_men_n1166_), .B(men_men_n112_), .C(men_men_n232_), .Y(men_men_n1592_));
  OAI220     u1564(.A0(men_men_n157_), .A1(men_men_n190_), .B0(men_men_n479_), .B1(u), .Y(men_men_n1593_));
  OAI210     u1565(.A0(men_men_n1593_), .A1(men_men_n114_), .B0(men_men_n1496_), .Y(men_men_n1594_));
  NA2        u1566(.A(men_men_n1594_), .B(men_men_n1592_), .Y(men_men_n1595_));
  NO3        u1567(.A(men_men_n1595_), .B(men_men_n1591_), .C(men_men_n1589_), .Y(men_men_n1596_));
  NO2        u1568(.A(men_men_n1440_), .B(e), .Y(men_men_n1597_));
  NA2        u1569(.A(men_men_n1597_), .B(men_men_n433_), .Y(men_men_n1598_));
  NA2        u1570(.A(men_men_n1198_), .B(men_men_n675_), .Y(men_men_n1599_));
  OR3        u1571(.A(men_men_n1554_), .B(men_men_n1292_), .C(men_men_n137_), .Y(men_men_n1600_));
  OAI220     u1572(.A0(men_men_n1600_), .A1(men_men_n1598_), .B0(men_men_n1599_), .B1(men_men_n473_), .Y(men_men_n1601_));
  NO3        u1573(.A(men_men_n1525_), .B(men_men_n377_), .C(a), .Y(men_men_n1602_));
  NO2        u1574(.A(men_men_n1602_), .B(men_men_n1601_), .Y(men_men_n1603_));
  NO2        u1575(.A(men_men_n190_), .B(c), .Y(men_men_n1604_));
  OAI210     u1576(.A0(men_men_n1604_), .A1(men_men_n1597_), .B0(men_men_n188_), .Y(men_men_n1605_));
  AOI220     u1577(.A0(men_men_n1605_), .A1(men_men_n1145_), .B0(men_men_n567_), .B1(men_men_n393_), .Y(men_men_n1606_));
  NA2        u1578(.A(men_men_n575_), .B(u), .Y(men_men_n1607_));
  AOI210     u1579(.A0(men_men_n1607_), .A1(men_men_n1479_), .B0(men_men_n1560_), .Y(men_men_n1608_));
  NO2        u1580(.A(men_men_n1517_), .B(f), .Y(men_men_n1609_));
  AOI210     u1581(.A0(men_men_n1198_), .A1(a), .B0(men_men_n1609_), .Y(men_men_n1610_));
  OAI220     u1582(.A0(men_men_n1610_), .A1(men_men_n69_), .B0(men_men_n1608_), .B1(men_men_n224_), .Y(men_men_n1611_));
  AOI210     u1583(.A0(men_men_n964_), .A1(men_men_n445_), .B0(men_men_n108_), .Y(men_men_n1612_));
  OR2        u1584(.A(men_men_n1612_), .B(men_men_n575_), .Y(men_men_n1613_));
  NA2        u1585(.A(men_men_n1609_), .B(men_men_n1455_), .Y(men_men_n1614_));
  OAI220     u1586(.A0(men_men_n1614_), .A1(men_men_n49_), .B0(men_men_n1613_), .B1(men_men_n183_), .Y(men_men_n1615_));
  NA4        u1587(.A(men_men_n1166_), .B(men_men_n1163_), .C(men_men_n232_), .D(men_men_n68_), .Y(men_men_n1616_));
  NA2        u1588(.A(men_men_n1445_), .B(men_men_n191_), .Y(men_men_n1617_));
  NO2        u1589(.A(men_men_n49_), .B(l), .Y(men_men_n1618_));
  OAI210     u1590(.A0(men_men_n1517_), .A1(men_men_n923_), .B0(men_men_n516_), .Y(men_men_n1619_));
  OAI210     u1591(.A0(men_men_n1619_), .A1(men_men_n1169_), .B0(men_men_n1618_), .Y(men_men_n1620_));
  NO2        u1592(.A(men_men_n266_), .B(u), .Y(men_men_n1621_));
  NO2        u1593(.A(m), .B(i), .Y(men_men_n1622_));
  AOI220     u1594(.A0(men_men_n1622_), .A1(men_men_n1481_), .B0(men_men_n1144_), .B1(men_men_n1621_), .Y(men_men_n1623_));
  NA4        u1595(.A(men_men_n1623_), .B(men_men_n1620_), .C(men_men_n1617_), .D(men_men_n1616_), .Y(men_men_n1624_));
  NO4        u1596(.A(men_men_n1624_), .B(men_men_n1615_), .C(men_men_n1611_), .D(men_men_n1606_), .Y(men_men_n1625_));
  NA3        u1597(.A(men_men_n1625_), .B(men_men_n1603_), .C(men_men_n1596_), .Y(men_men_n1626_));
  NA3        u1598(.A(men_men_n1027_), .B(men_men_n144_), .C(men_men_n46_), .Y(men_men_n1627_));
  AOI210     u1599(.A0(men_men_n154_), .A1(c), .B0(men_men_n1627_), .Y(men_men_n1628_));
  OAI210     u1600(.A0(men_men_n620_), .A1(u), .B0(men_men_n194_), .Y(men_men_n1629_));
  NA2        u1601(.A(men_men_n1629_), .B(men_men_n1562_), .Y(men_men_n1630_));
  AO210      u1602(.A0(men_men_n138_), .A1(l), .B0(men_men_n1506_), .Y(men_men_n1631_));
  NO2        u1603(.A(men_men_n72_), .B(c), .Y(men_men_n1632_));
  NO4        u1604(.A(men_men_n1467_), .B(men_men_n195_), .C(men_men_n479_), .D(men_men_n45_), .Y(men_men_n1633_));
  AOI210     u1605(.A0(men_men_n1572_), .A1(men_men_n1632_), .B0(men_men_n1633_), .Y(men_men_n1634_));
  NA3        u1606(.A(men_men_n1634_), .B(men_men_n1631_), .C(men_men_n1630_), .Y(men_men_n1635_));
  NO2        u1607(.A(men_men_n1635_), .B(men_men_n1628_), .Y(men_men_n1636_));
  NO4        u1608(.A(men_men_n236_), .B(men_men_n195_), .C(men_men_n271_), .D(k), .Y(men_men_n1637_));
  AOI210     u1609(.A0(men_men_n163_), .A1(men_men_n56_), .B0(men_men_n1597_), .Y(men_men_n1638_));
  NO2        u1610(.A(men_men_n1638_), .B(men_men_n1566_), .Y(men_men_n1639_));
  NO2        u1611(.A(men_men_n1627_), .B(men_men_n114_), .Y(men_men_n1640_));
  NOi21      u1612(.An(men_men_n1445_), .B(e), .Y(men_men_n1641_));
  NO4        u1613(.A(men_men_n1641_), .B(men_men_n1640_), .C(men_men_n1639_), .D(men_men_n1637_), .Y(men_men_n1642_));
  AN2        u1614(.A(men_men_n1166_), .B(men_men_n1151_), .Y(men_men_n1643_));
  AOI220     u1615(.A0(men_men_n1622_), .A1(men_men_n685_), .B0(men_men_n1128_), .B1(men_men_n166_), .Y(men_men_n1644_));
  NOi31      u1616(.An(men_men_n30_), .B(men_men_n1644_), .C(n), .Y(men_men_n1645_));
  AOI210     u1617(.A0(men_men_n1643_), .A1(men_men_n1244_), .B0(men_men_n1645_), .Y(men_men_n1646_));
  NO2        u1618(.A(men_men_n1565_), .B(men_men_n69_), .Y(men_men_n1647_));
  NA2        u1619(.A(men_men_n59_), .B(a), .Y(men_men_n1648_));
  NO2        u1620(.A(men_men_n1453_), .B(men_men_n122_), .Y(men_men_n1649_));
  OAI220     u1621(.A0(men_men_n1649_), .A1(men_men_n1506_), .B0(men_men_n1526_), .B1(men_men_n1648_), .Y(men_men_n1650_));
  NO2        u1622(.A(men_men_n1650_), .B(men_men_n1647_), .Y(men_men_n1651_));
  NA4        u1623(.A(men_men_n1651_), .B(men_men_n1646_), .C(men_men_n1642_), .D(men_men_n1636_), .Y(men_men_n1652_));
  OR4        u1624(.A(men_men_n1652_), .B(men_men_n1626_), .C(men_men_n1582_), .D(men_men_n1530_), .Y(men04));
  NOi31      u1625(.An(men_men_n1514_), .B(men_men_n1515_), .C(men_men_n1116_), .Y(men_men_n1654_));
  NA2        u1626(.A(men_men_n1576_), .B(men_men_n883_), .Y(men_men_n1655_));
  NO4        u1627(.A(men_men_n1655_), .B(men_men_n1106_), .C(men_men_n517_), .D(j), .Y(men_men_n1656_));
  OR3        u1628(.A(men_men_n1656_), .B(men_men_n1654_), .C(men_men_n1134_), .Y(men_men_n1657_));
  NO3        u1629(.A(men_men_n1455_), .B(men_men_n93_), .C(k), .Y(men_men_n1658_));
  AOI210     u1630(.A0(men_men_n1658_), .A1(men_men_n1127_), .B0(men_men_n1266_), .Y(men_men_n1659_));
  NA2        u1631(.A(men_men_n1659_), .B(men_men_n1296_), .Y(men_men_n1660_));
  NO4        u1632(.A(men_men_n1660_), .B(men_men_n1657_), .C(men_men_n1142_), .D(men_men_n1121_), .Y(men_men_n1661_));
  NA4        u1633(.A(men_men_n1661_), .B(men_men_n1200_), .C(men_men_n1185_), .D(men_men_n1172_), .Y(men05));
  INV        u1634(.A(l), .Y(men_men_n1665_));
  INV        u1635(.A(b), .Y(men_men_n1666_));
  INV        u1636(.A(e), .Y(men_men_n1667_));
  INV        u1637(.A(a), .Y(men_men_n1668_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule