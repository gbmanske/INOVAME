// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n133_, new_new_n134_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n583_, new_new_n584_, new_new_n585_, new_new_n586_,
    new_new_n587_, new_new_n588_, new_new_n589_, new_new_n590_,
    new_new_n591_, new_new_n592_, new_new_n593_, new_new_n594_,
    new_new_n595_, new_new_n596_, new_new_n597_, new_new_n598_,
    new_new_n599_, new_new_n600_, new_new_n601_, new_new_n602_,
    new_new_n603_, new_new_n604_, new_new_n605_, new_new_n606_,
    new_new_n607_, new_new_n608_, new_new_n609_, new_new_n610_,
    new_new_n611_, new_new_n612_, new_new_n613_, new_new_n614_,
    new_new_n615_, new_new_n616_, new_new_n617_, new_new_n618_,
    new_new_n619_, new_new_n620_, new_new_n621_, new_new_n622_,
    new_new_n623_, new_new_n624_, new_new_n625_, new_new_n626_,
    new_new_n627_, new_new_n629_, new_new_n630_, new_new_n631_,
    new_new_n632_, new_new_n633_, new_new_n634_, new_new_n635_,
    new_new_n636_, new_new_n637_, new_new_n638_, new_new_n639_,
    new_new_n640_, new_new_n641_, new_new_n642_, new_new_n643_,
    new_new_n644_, new_new_n645_, new_new_n646_, new_new_n647_,
    new_new_n648_, new_new_n649_, new_new_n650_, new_new_n651_,
    new_new_n652_, new_new_n653_, new_new_n654_, new_new_n655_,
    new_new_n656_, new_new_n657_, new_new_n658_, new_new_n659_,
    new_new_n660_, new_new_n661_, new_new_n662_, new_new_n663_,
    new_new_n664_, new_new_n665_, new_new_n666_, new_new_n667_,
    new_new_n668_, new_new_n669_, new_new_n670_, new_new_n671_,
    new_new_n672_, new_new_n674_, new_new_n675_, new_new_n676_,
    new_new_n677_, new_new_n678_, new_new_n679_, new_new_n680_,
    new_new_n681_, new_new_n682_, new_new_n683_, new_new_n684_,
    new_new_n685_, new_new_n686_, new_new_n687_, new_new_n688_,
    new_new_n689_, new_new_n690_, new_new_n691_, new_new_n692_,
    new_new_n693_, new_new_n694_, new_new_n695_, new_new_n696_,
    new_new_n697_, new_new_n698_, new_new_n699_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n703_, new_new_n704_,
    new_new_n705_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n827_,
    new_new_n828_, new_new_n829_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n55_));
  NO2        g033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  NAi21      g035(.An(i_2_), .B(i_7_), .Y(new_new_n58_));
  INV        g036(.A(i_1_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_6_), .Y(new_new_n60_));
  NA3        g038(.A(new_new_n60_), .B(new_new_n58_), .C(new_new_n31_), .Y(new_new_n61_));
  NA2        g039(.A(i_1_), .B(i_10_), .Y(new_new_n62_));
  NO2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NAi21      g041(.An(new_new_n63_), .B(new_new_n61_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n50_), .B(i_2_), .Y(new_new_n65_));
  AOI210     g043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_6_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(new_new_n25_), .Y(new_new_n68_));
  INV        g046(.A(i_0_), .Y(new_new_n69_));
  NAi21      g047(.An(i_5_), .B(i_10_), .Y(new_new_n70_));
  NA2        g048(.A(i_5_), .B(i_9_), .Y(new_new_n71_));
  AOI210     g049(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n69_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n72_), .B(new_new_n68_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n66_), .A1(new_new_n65_), .B0(new_new_n73_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n74_), .A1(new_new_n64_), .B0(i_0_), .Y(new_new_n75_));
  NA2        g053(.A(i_12_), .B(i_5_), .Y(new_new_n76_));
  NA2        g054(.A(i_2_), .B(i_8_), .Y(new_new_n77_));
  NO2        g055(.A(new_new_n77_), .B(new_new_n56_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_7_), .Y(new_new_n79_));
  INV        g057(.A(i_6_), .Y(new_new_n80_));
  OR4        g058(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n81_));
  INV        g059(.A(new_new_n81_), .Y(new_new_n82_));
  NO2        g060(.A(i_2_), .B(i_7_), .Y(new_new_n83_));
  INV        g061(.A(new_new_n78_), .Y(new_new_n84_));
  NAi21      g062(.An(i_6_), .B(i_10_), .Y(new_new_n85_));
  NA2        g063(.A(i_6_), .B(i_9_), .Y(new_new_n86_));
  AOI210     g064(.A0(new_new_n86_), .A1(new_new_n85_), .B0(new_new_n59_), .Y(new_new_n87_));
  NA2        g065(.A(i_2_), .B(i_6_), .Y(new_new_n88_));
  NO2        g066(.A(new_new_n88_), .B(new_new_n25_), .Y(new_new_n89_));
  NO2        g067(.A(new_new_n89_), .B(new_new_n87_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n84_), .B0(new_new_n76_), .Y(new_new_n91_));
  AN3        g069(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n92_));
  NAi21      g070(.An(i_6_), .B(i_11_), .Y(new_new_n93_));
  NA2        g071(.A(new_new_n92_), .B(new_new_n32_), .Y(new_new_n94_));
  INV        g072(.A(i_7_), .Y(new_new_n95_));
  NA2        g073(.A(new_new_n46_), .B(new_new_n95_), .Y(new_new_n96_));
  NO2        g074(.A(i_0_), .B(i_5_), .Y(new_new_n97_));
  NO2        g075(.A(new_new_n97_), .B(new_new_n80_), .Y(new_new_n98_));
  NA2        g076(.A(i_12_), .B(i_3_), .Y(new_new_n99_));
  INV        g077(.A(new_new_n99_), .Y(new_new_n100_));
  NA3        g078(.A(new_new_n100_), .B(new_new_n98_), .C(new_new_n96_), .Y(new_new_n101_));
  NAi21      g079(.An(i_7_), .B(i_11_), .Y(new_new_n102_));
  NO3        g080(.A(new_new_n102_), .B(new_new_n85_), .C(new_new_n53_), .Y(new_new_n103_));
  AN2        g081(.A(i_2_), .B(i_10_), .Y(new_new_n104_));
  NO2        g082(.A(new_new_n104_), .B(i_7_), .Y(new_new_n105_));
  OR2        g083(.A(new_new_n76_), .B(new_new_n56_), .Y(new_new_n106_));
  NO2        g084(.A(i_8_), .B(new_new_n95_), .Y(new_new_n107_));
  NO3        g085(.A(new_new_n107_), .B(new_new_n106_), .C(new_new_n105_), .Y(new_new_n108_));
  NA2        g086(.A(i_12_), .B(i_7_), .Y(new_new_n109_));
  NO2        g087(.A(new_new_n59_), .B(new_new_n26_), .Y(new_new_n110_));
  NA2        g088(.A(new_new_n110_), .B(i_0_), .Y(new_new_n111_));
  NA2        g089(.A(i_11_), .B(i_12_), .Y(new_new_n112_));
  OAI210     g090(.A0(new_new_n111_), .A1(new_new_n109_), .B0(new_new_n112_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n113_), .B(new_new_n108_), .Y(new_new_n114_));
  NAi41      g092(.An(new_new_n103_), .B(new_new_n114_), .C(new_new_n101_), .D(new_new_n94_), .Y(new_new_n115_));
  NOi21      g093(.An(i_1_), .B(i_5_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(i_11_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n95_), .B(new_new_n37_), .Y(new_new_n118_));
  NA2        g096(.A(i_7_), .B(new_new_n25_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(new_new_n118_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(new_new_n46_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n86_), .B(new_new_n85_), .Y(new_new_n122_));
  NAi21      g100(.An(i_3_), .B(i_8_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n58_), .Y(new_new_n124_));
  NOi31      g102(.An(new_new_n124_), .B(new_new_n122_), .C(new_new_n121_), .Y(new_new_n125_));
  NO2        g103(.A(i_1_), .B(new_new_n80_), .Y(new_new_n126_));
  NO2        g104(.A(i_6_), .B(i_5_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(i_3_), .Y(new_new_n128_));
  AO210      g106(.A0(new_new_n128_), .A1(new_new_n47_), .B0(new_new_n126_), .Y(new_new_n129_));
  OAI220     g107(.A0(new_new_n129_), .A1(new_new_n102_), .B0(new_new_n125_), .B1(new_new_n117_), .Y(new_new_n130_));
  NO3        g108(.A(new_new_n130_), .B(new_new_n115_), .C(new_new_n91_), .Y(new_new_n131_));
  NA3        g109(.A(new_new_n131_), .B(new_new_n75_), .C(new_new_n55_), .Y(ori2));
  NO2        g110(.A(new_new_n59_), .B(new_new_n37_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n828_), .B(new_new_n133_), .Y(new_new_n134_));
  NA4        g112(.A(new_new_n134_), .B(new_new_n73_), .C(new_new_n65_), .D(new_new_n30_), .Y(ori0));
  AN2        g113(.A(i_8_), .B(i_7_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(i_6_), .Y(new_new_n137_));
  NO2        g115(.A(i_12_), .B(i_13_), .Y(new_new_n138_));
  NAi21      g116(.An(i_5_), .B(i_11_), .Y(new_new_n139_));
  NOi21      g117(.An(new_new_n138_), .B(new_new_n139_), .Y(new_new_n140_));
  NO2        g118(.A(i_0_), .B(i_1_), .Y(new_new_n141_));
  NA2        g119(.A(i_2_), .B(i_3_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n142_), .B(i_4_), .Y(new_new_n143_));
  NA3        g121(.A(new_new_n143_), .B(new_new_n141_), .C(new_new_n140_), .Y(new_new_n144_));
  NA2        g122(.A(i_1_), .B(i_5_), .Y(new_new_n145_));
  OR2        g123(.A(i_0_), .B(i_1_), .Y(new_new_n146_));
  NAi32      g124(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n147_));
  NOi21      g125(.An(i_4_), .B(i_10_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n40_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n69_), .B(i_2_), .C(i_1_), .Y(new_new_n150_));
  INV        g128(.A(new_new_n150_), .Y(new_new_n151_));
  NOi21      g129(.An(i_4_), .B(i_9_), .Y(new_new_n152_));
  NOi21      g130(.An(i_11_), .B(i_13_), .Y(new_new_n153_));
  NA2        g131(.A(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  NO2        g132(.A(i_4_), .B(i_5_), .Y(new_new_n155_));
  NAi21      g133(.An(i_12_), .B(i_11_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n156_), .B(i_13_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n69_), .B(new_new_n59_), .Y(new_new_n158_));
  NA2        g136(.A(i_3_), .B(i_5_), .Y(new_new_n159_));
  NO2        g137(.A(new_new_n69_), .B(i_5_), .Y(new_new_n160_));
  NO2        g138(.A(i_13_), .B(i_10_), .Y(new_new_n161_));
  NA3        g139(.A(new_new_n161_), .B(new_new_n160_), .C(new_new_n44_), .Y(new_new_n162_));
  NO2        g140(.A(i_2_), .B(i_1_), .Y(new_new_n163_));
  NA2        g141(.A(new_new_n163_), .B(i_3_), .Y(new_new_n164_));
  NAi21      g142(.An(i_4_), .B(i_12_), .Y(new_new_n165_));
  INV        g143(.A(i_8_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n166_), .B(i_7_), .Y(new_new_n167_));
  NO3        g145(.A(i_3_), .B(new_new_n80_), .C(new_new_n48_), .Y(new_new_n168_));
  NA2        g146(.A(new_new_n168_), .B(new_new_n107_), .Y(new_new_n169_));
  NO3        g147(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n170_));
  NO3        g148(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n171_));
  NO2        g149(.A(i_3_), .B(i_8_), .Y(new_new_n172_));
  NO3        g150(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n173_));
  NA3        g151(.A(new_new_n173_), .B(new_new_n172_), .C(new_new_n40_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n97_), .B(new_new_n56_), .Y(new_new_n175_));
  INV        g153(.A(new_new_n175_), .Y(new_new_n176_));
  NO2        g154(.A(i_13_), .B(i_9_), .Y(new_new_n177_));
  NAi21      g155(.An(i_12_), .B(i_3_), .Y(new_new_n178_));
  NO2        g156(.A(new_new_n44_), .B(i_5_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n176_), .B(new_new_n174_), .Y(new_new_n180_));
  NA2        g158(.A(new_new_n180_), .B(i_7_), .Y(new_new_n181_));
  NO2        g159(.A(new_new_n181_), .B(i_4_), .Y(new_new_n182_));
  NAi21      g160(.An(i_12_), .B(i_7_), .Y(new_new_n183_));
  NA3        g161(.A(i_13_), .B(new_new_n166_), .C(i_10_), .Y(new_new_n184_));
  NO2        g162(.A(new_new_n184_), .B(new_new_n183_), .Y(new_new_n185_));
  NA2        g163(.A(i_0_), .B(i_5_), .Y(new_new_n186_));
  OAI220     g164(.A0(new_new_n80_), .A1(new_new_n164_), .B0(i_2_), .B1(new_new_n128_), .Y(new_new_n187_));
  NAi31      g165(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n36_), .B(i_13_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n46_), .B(new_new_n59_), .Y(new_new_n190_));
  NA3        g168(.A(new_new_n190_), .B(i_3_), .C(new_new_n189_), .Y(new_new_n191_));
  INV        g169(.A(i_13_), .Y(new_new_n192_));
  NO2        g170(.A(i_12_), .B(new_new_n192_), .Y(new_new_n193_));
  NA3        g171(.A(new_new_n193_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n194_));
  OAI210     g172(.A0(new_new_n191_), .A1(new_new_n188_), .B0(new_new_n194_), .Y(new_new_n195_));
  AOI220     g173(.A0(new_new_n195_), .A1(new_new_n136_), .B0(new_new_n187_), .B1(new_new_n185_), .Y(new_new_n196_));
  NO2        g174(.A(i_12_), .B(new_new_n37_), .Y(new_new_n197_));
  OR2        g175(.A(i_8_), .B(i_7_), .Y(new_new_n198_));
  INV        g176(.A(i_12_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n44_), .B(new_new_n199_), .Y(new_new_n200_));
  NO3        g178(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n201_));
  NA2        g179(.A(i_2_), .B(i_1_), .Y(new_new_n202_));
  NO3        g180(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n203_));
  NAi21      g181(.An(i_4_), .B(i_3_), .Y(new_new_n204_));
  NO2        g182(.A(i_0_), .B(i_6_), .Y(new_new_n205_));
  NOi41      g183(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n202_), .B(new_new_n159_), .Y(new_new_n207_));
  NO2        g185(.A(i_11_), .B(new_new_n192_), .Y(new_new_n208_));
  NOi21      g186(.An(i_1_), .B(i_6_), .Y(new_new_n209_));
  NAi21      g187(.An(i_3_), .B(i_7_), .Y(new_new_n210_));
  NA2        g188(.A(new_new_n199_), .B(i_9_), .Y(new_new_n211_));
  OR4        g189(.A(new_new_n211_), .B(new_new_n210_), .C(new_new_n209_), .D(new_new_n160_), .Y(new_new_n212_));
  NO2        g190(.A(i_12_), .B(i_3_), .Y(new_new_n213_));
  NA2        g191(.A(new_new_n69_), .B(i_5_), .Y(new_new_n214_));
  NA2        g192(.A(i_3_), .B(i_9_), .Y(new_new_n215_));
  NAi21      g193(.An(i_7_), .B(i_10_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NA3        g195(.A(new_new_n217_), .B(new_new_n214_), .C(new_new_n60_), .Y(new_new_n218_));
  NA2        g196(.A(new_new_n218_), .B(new_new_n212_), .Y(new_new_n219_));
  INV        g197(.A(new_new_n137_), .Y(new_new_n220_));
  NA2        g198(.A(new_new_n199_), .B(i_13_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n221_), .B(new_new_n71_), .Y(new_new_n222_));
  AOI220     g200(.A0(new_new_n222_), .A1(new_new_n220_), .B0(new_new_n219_), .B1(new_new_n208_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n198_), .B(new_new_n37_), .Y(new_new_n224_));
  NA2        g202(.A(i_12_), .B(i_6_), .Y(new_new_n225_));
  OR2        g203(.A(i_13_), .B(i_9_), .Y(new_new_n226_));
  NO3        g204(.A(new_new_n226_), .B(new_new_n225_), .C(new_new_n48_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n204_), .B(i_2_), .Y(new_new_n228_));
  NA3        g206(.A(new_new_n228_), .B(new_new_n227_), .C(new_new_n44_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n208_), .B(i_9_), .Y(new_new_n230_));
  NA2        g208(.A(new_new_n214_), .B(new_new_n60_), .Y(new_new_n231_));
  OAI210     g209(.A0(new_new_n231_), .A1(new_new_n230_), .B0(new_new_n229_), .Y(new_new_n232_));
  NO3        g210(.A(i_11_), .B(new_new_n192_), .C(new_new_n25_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n210_), .B(i_8_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n232_), .B(new_new_n224_), .Y(new_new_n235_));
  NA3        g213(.A(new_new_n235_), .B(new_new_n223_), .C(new_new_n196_), .Y(new_new_n236_));
  NO3        g214(.A(i_12_), .B(new_new_n192_), .C(new_new_n37_), .Y(new_new_n237_));
  INV        g215(.A(new_new_n237_), .Y(new_new_n238_));
  NO3        g216(.A(i_0_), .B(i_2_), .C(new_new_n59_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n202_), .B(i_0_), .Y(new_new_n240_));
  AOI220     g218(.A0(new_new_n240_), .A1(new_new_n167_), .B0(new_new_n239_), .B1(new_new_n136_), .Y(new_new_n241_));
  NA2        g219(.A(i_5_), .B(new_new_n26_), .Y(new_new_n242_));
  NO2        g220(.A(new_new_n242_), .B(new_new_n241_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n151_), .B(new_new_n137_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n244_), .B(new_new_n243_), .Y(new_new_n245_));
  NO2        g223(.A(i_3_), .B(i_10_), .Y(new_new_n246_));
  NO2        g224(.A(i_2_), .B(new_new_n95_), .Y(new_new_n247_));
  AN2        g225(.A(i_3_), .B(i_10_), .Y(new_new_n248_));
  NO2        g226(.A(i_5_), .B(new_new_n37_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n245_), .B(new_new_n238_), .Y(new_new_n251_));
  NO3        g229(.A(new_new_n251_), .B(new_new_n236_), .C(new_new_n182_), .Y(new_new_n252_));
  NO3        g230(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n253_));
  NO3        g231(.A(i_6_), .B(new_new_n166_), .C(i_7_), .Y(new_new_n254_));
  NO2        g232(.A(i_2_), .B(i_3_), .Y(new_new_n255_));
  OR2        g233(.A(i_0_), .B(i_5_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n146_), .B(new_new_n46_), .Y(new_new_n257_));
  NO2        g235(.A(i_12_), .B(i_10_), .Y(new_new_n258_));
  NOi21      g236(.An(i_5_), .B(i_0_), .Y(new_new_n259_));
  NO2        g237(.A(i_2_), .B(new_new_n95_), .Y(new_new_n260_));
  NO4        g238(.A(new_new_n260_), .B(i_4_), .C(new_new_n259_), .D(new_new_n123_), .Y(new_new_n261_));
  NA4        g239(.A(new_new_n79_), .B(new_new_n36_), .C(new_new_n80_), .D(i_8_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n261_), .B(new_new_n258_), .Y(new_new_n263_));
  NO2        g241(.A(i_6_), .B(i_8_), .Y(new_new_n264_));
  NOi21      g242(.An(i_0_), .B(i_2_), .Y(new_new_n265_));
  AN2        g243(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n266_));
  NO2        g244(.A(i_1_), .B(i_7_), .Y(new_new_n267_));
  INV        g245(.A(new_new_n263_), .Y(new_new_n268_));
  NA3        g246(.A(new_new_n209_), .B(new_new_n247_), .C(new_new_n166_), .Y(new_new_n269_));
  NO2        g247(.A(new_new_n166_), .B(i_9_), .Y(new_new_n270_));
  NA2        g248(.A(new_new_n270_), .B(new_new_n175_), .Y(new_new_n271_));
  INV        g249(.A(new_new_n243_), .Y(new_new_n272_));
  AOI210     g250(.A0(new_new_n272_), .A1(new_new_n269_), .B0(new_new_n149_), .Y(new_new_n273_));
  AOI210     g251(.A0(new_new_n268_), .A1(new_new_n253_), .B0(new_new_n273_), .Y(new_new_n274_));
  NOi32      g252(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n275_));
  INV        g253(.A(new_new_n275_), .Y(new_new_n276_));
  NAi21      g254(.An(i_0_), .B(i_6_), .Y(new_new_n277_));
  NAi21      g255(.An(i_1_), .B(i_5_), .Y(new_new_n278_));
  NA2        g256(.A(new_new_n278_), .B(new_new_n277_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n279_), .B(new_new_n25_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(new_new_n147_), .Y(new_new_n281_));
  NAi41      g259(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n282_));
  OAI220     g260(.A0(new_new_n282_), .A1(new_new_n278_), .B0(new_new_n188_), .B1(new_new_n147_), .Y(new_new_n283_));
  AOI210     g261(.A0(new_new_n282_), .A1(new_new_n147_), .B0(new_new_n146_), .Y(new_new_n284_));
  NOi32      g262(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n285_));
  NAi21      g263(.An(i_6_), .B(i_1_), .Y(new_new_n286_));
  NA3        g264(.A(new_new_n286_), .B(new_new_n285_), .C(new_new_n46_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n287_), .B(i_0_), .Y(new_new_n288_));
  OR3        g266(.A(new_new_n288_), .B(new_new_n284_), .C(new_new_n283_), .Y(new_new_n289_));
  NO2        g267(.A(i_1_), .B(new_new_n95_), .Y(new_new_n290_));
  NAi21      g268(.An(i_3_), .B(i_4_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n291_), .B(i_9_), .Y(new_new_n292_));
  AN2        g270(.A(i_6_), .B(i_7_), .Y(new_new_n293_));
  OAI210     g271(.A0(new_new_n293_), .A1(new_new_n290_), .B0(new_new_n292_), .Y(new_new_n294_));
  NA2        g272(.A(i_2_), .B(i_7_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n291_), .B(i_10_), .Y(new_new_n296_));
  NA3        g274(.A(new_new_n296_), .B(new_new_n295_), .C(new_new_n205_), .Y(new_new_n297_));
  AOI210     g275(.A0(new_new_n297_), .A1(new_new_n294_), .B0(new_new_n160_), .Y(new_new_n298_));
  AOI210     g276(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n299_));
  OAI210     g277(.A0(new_new_n299_), .A1(new_new_n163_), .B0(new_new_n296_), .Y(new_new_n300_));
  AOI220     g278(.A0(new_new_n296_), .A1(new_new_n267_), .B0(new_new_n201_), .B1(new_new_n163_), .Y(new_new_n301_));
  AOI210     g279(.A0(new_new_n301_), .A1(new_new_n300_), .B0(i_5_), .Y(new_new_n302_));
  NO4        g280(.A(new_new_n302_), .B(new_new_n298_), .C(new_new_n289_), .D(new_new_n281_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n303_), .B(new_new_n276_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n305_));
  AN2        g283(.A(i_12_), .B(i_5_), .Y(new_new_n306_));
  NA2        g284(.A(new_new_n829_), .B(new_new_n306_), .Y(new_new_n307_));
  NO2        g285(.A(i_11_), .B(i_6_), .Y(new_new_n308_));
  NA3        g286(.A(new_new_n308_), .B(new_new_n257_), .C(new_new_n192_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n309_), .B(new_new_n307_), .Y(new_new_n310_));
  NO2        g288(.A(i_5_), .B(i_10_), .Y(new_new_n311_));
  NA2        g289(.A(new_new_n311_), .B(new_new_n228_), .Y(new_new_n312_));
  NA2        g290(.A(new_new_n138_), .B(new_new_n45_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n313_), .B(new_new_n312_), .Y(new_new_n314_));
  OAI210     g292(.A0(new_new_n314_), .A1(new_new_n310_), .B0(new_new_n305_), .Y(new_new_n315_));
  NO2        g293(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n316_));
  NO2        g294(.A(new_new_n144_), .B(new_new_n80_), .Y(new_new_n317_));
  OAI210     g295(.A0(new_new_n317_), .A1(new_new_n310_), .B0(new_new_n316_), .Y(new_new_n318_));
  NO3        g296(.A(new_new_n80_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n319_));
  NA3        g297(.A(new_new_n246_), .B(new_new_n71_), .C(new_new_n54_), .Y(new_new_n320_));
  NO2        g298(.A(i_11_), .B(i_12_), .Y(new_new_n321_));
  NA2        g299(.A(new_new_n321_), .B(new_new_n36_), .Y(new_new_n322_));
  NO2        g300(.A(new_new_n320_), .B(new_new_n322_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n311_), .B(new_new_n199_), .Y(new_new_n324_));
  NAi21      g302(.An(i_13_), .B(i_0_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n325_), .B(new_new_n202_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n323_), .B(new_new_n326_), .Y(new_new_n327_));
  NA3        g305(.A(new_new_n327_), .B(new_new_n318_), .C(new_new_n315_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n44_), .B(new_new_n192_), .Y(new_new_n329_));
  NO3        g307(.A(i_1_), .B(i_12_), .C(new_new_n80_), .Y(new_new_n330_));
  NO2        g308(.A(i_0_), .B(i_11_), .Y(new_new_n331_));
  NOi21      g309(.An(i_2_), .B(i_12_), .Y(new_new_n332_));
  OR2        g310(.A(i_13_), .B(i_10_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n154_), .B(new_new_n118_), .Y(new_new_n334_));
  NO2        g312(.A(new_new_n95_), .B(new_new_n25_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n159_), .B(new_new_n80_), .Y(new_new_n336_));
  NA2        g314(.A(new_new_n166_), .B(i_10_), .Y(new_new_n337_));
  NA3        g315(.A(new_new_n214_), .B(new_new_n60_), .C(i_2_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n338_), .B(new_new_n337_), .Y(new_new_n339_));
  NO2        g317(.A(i_3_), .B(new_new_n48_), .Y(new_new_n340_));
  NA3        g318(.A(new_new_n267_), .B(new_new_n266_), .C(new_new_n340_), .Y(new_new_n341_));
  INV        g319(.A(new_new_n254_), .Y(new_new_n342_));
  OAI210     g320(.A0(new_new_n342_), .A1(new_new_n164_), .B0(new_new_n341_), .Y(new_new_n343_));
  NO2        g321(.A(new_new_n343_), .B(new_new_n339_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n344_), .B(new_new_n230_), .Y(new_new_n345_));
  NO3        g323(.A(new_new_n345_), .B(new_new_n328_), .C(new_new_n304_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n69_), .B(i_13_), .Y(new_new_n347_));
  NO2        g325(.A(i_10_), .B(i_9_), .Y(new_new_n348_));
  NAi21      g326(.An(i_12_), .B(i_8_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(i_3_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n46_), .B(i_4_), .Y(new_new_n351_));
  NA2        g329(.A(new_new_n351_), .B(new_new_n98_), .Y(new_new_n352_));
  NO2        g330(.A(new_new_n352_), .B(new_new_n174_), .Y(new_new_n353_));
  NA2        g331(.A(new_new_n250_), .B(i_0_), .Y(new_new_n354_));
  NO3        g332(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n355_));
  NA2        g333(.A(new_new_n225_), .B(new_new_n93_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n356_), .B(new_new_n355_), .Y(new_new_n357_));
  NA2        g335(.A(i_8_), .B(i_9_), .Y(new_new_n358_));
  AOI210     g336(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n359_));
  OR2        g337(.A(new_new_n359_), .B(new_new_n358_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n237_), .B(new_new_n175_), .Y(new_new_n361_));
  OAI220     g339(.A0(new_new_n361_), .A1(new_new_n360_), .B0(new_new_n357_), .B1(new_new_n354_), .Y(new_new_n362_));
  NA2        g340(.A(new_new_n208_), .B(new_new_n249_), .Y(new_new_n363_));
  NO3        g341(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n364_));
  INV        g342(.A(new_new_n364_), .Y(new_new_n365_));
  NA3        g343(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n366_));
  NA4        g344(.A(new_new_n139_), .B(new_new_n110_), .C(new_new_n76_), .D(new_new_n23_), .Y(new_new_n367_));
  OAI220     g345(.A0(new_new_n367_), .A1(new_new_n366_), .B0(new_new_n365_), .B1(new_new_n363_), .Y(new_new_n368_));
  NO3        g346(.A(new_new_n368_), .B(new_new_n362_), .C(new_new_n353_), .Y(new_new_n369_));
  OR2        g347(.A(new_new_n271_), .B(new_new_n149_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n92_), .B(i_13_), .Y(new_new_n371_));
  NA2        g349(.A(new_new_n336_), .B(new_new_n305_), .Y(new_new_n372_));
  NO2        g350(.A(i_2_), .B(i_13_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n372_), .B(new_new_n371_), .Y(new_new_n374_));
  NO3        g352(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n375_));
  NO2        g353(.A(i_6_), .B(i_7_), .Y(new_new_n376_));
  NO2        g354(.A(i_11_), .B(i_1_), .Y(new_new_n377_));
  OR2        g355(.A(i_11_), .B(i_8_), .Y(new_new_n378_));
  NOi21      g356(.An(i_2_), .B(i_7_), .Y(new_new_n379_));
  NO2        g357(.A(i_3_), .B(new_new_n166_), .Y(new_new_n380_));
  NO2        g358(.A(i_6_), .B(i_10_), .Y(new_new_n381_));
  NA3        g359(.A(new_new_n206_), .B(new_new_n153_), .C(new_new_n127_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n146_), .B(i_3_), .Y(new_new_n384_));
  NAi31      g362(.An(new_new_n383_), .B(new_new_n384_), .C(new_new_n193_), .Y(new_new_n385_));
  NA3        g363(.A(new_new_n316_), .B(new_new_n158_), .C(new_new_n143_), .Y(new_new_n386_));
  NA3        g364(.A(new_new_n386_), .B(new_new_n385_), .C(new_new_n382_), .Y(new_new_n387_));
  NO2        g365(.A(new_new_n387_), .B(new_new_n374_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n355_), .B(new_new_n306_), .Y(new_new_n389_));
  NA2        g367(.A(new_new_n364_), .B(new_new_n311_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n191_), .Y(new_new_n391_));
  NAi21      g369(.An(new_new_n184_), .B(new_new_n321_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n267_), .B(new_new_n186_), .Y(new_new_n393_));
  NO2        g371(.A(new_new_n393_), .B(new_new_n392_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n253_), .B(new_new_n201_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n395_), .B(new_new_n338_), .Y(new_new_n396_));
  NO3        g374(.A(new_new_n396_), .B(new_new_n394_), .C(new_new_n391_), .Y(new_new_n397_));
  NA4        g375(.A(new_new_n397_), .B(new_new_n388_), .C(new_new_n370_), .D(new_new_n369_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n117_), .B(new_new_n106_), .Y(new_new_n399_));
  AN2        g377(.A(new_new_n399_), .B(new_new_n355_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n400_), .B(new_new_n250_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n275_), .B(new_new_n69_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n36_), .B(i_8_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n39_), .B(i_13_), .Y(new_new_n404_));
  OAI210     g382(.A0(i_8_), .A1(new_new_n59_), .B0(new_new_n129_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n405_), .B(new_new_n334_), .Y(new_new_n406_));
  NA3        g384(.A(new_new_n406_), .B(new_new_n404_), .C(new_new_n401_), .Y(new_new_n407_));
  NO2        g385(.A(i_12_), .B(new_new_n166_), .Y(new_new_n408_));
  NO2        g386(.A(i_8_), .B(i_7_), .Y(new_new_n409_));
  AOI220     g387(.A0(new_new_n336_), .A1(new_new_n257_), .B0(new_new_n207_), .B1(new_new_n205_), .Y(new_new_n410_));
  OAI220     g388(.A0(new_new_n410_), .A1(new_new_n221_), .B0(new_new_n371_), .B1(new_new_n128_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n411_), .B(new_new_n224_), .Y(new_new_n412_));
  NA3        g390(.A(new_new_n248_), .B(new_new_n155_), .C(new_new_n92_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n146_), .B(i_5_), .Y(new_new_n414_));
  NA3        g392(.A(new_new_n414_), .B(new_new_n329_), .C(new_new_n255_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n415_), .B(new_new_n413_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n416_), .B(new_new_n364_), .Y(new_new_n417_));
  NA2        g395(.A(new_new_n417_), .B(new_new_n412_), .Y(new_new_n418_));
  AOI210     g396(.A0(new_new_n286_), .A1(new_new_n46_), .B0(new_new_n290_), .Y(new_new_n419_));
  NA2        g397(.A(i_0_), .B(new_new_n48_), .Y(new_new_n420_));
  NA3        g398(.A(new_new_n408_), .B(new_new_n233_), .C(new_new_n420_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n419_), .B(new_new_n421_), .Y(new_new_n422_));
  INV        g400(.A(new_new_n422_), .Y(new_new_n423_));
  NO4        g401(.A(new_new_n209_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n424_));
  NO3        g402(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n198_), .B(new_new_n36_), .Y(new_new_n426_));
  NO2        g404(.A(new_new_n333_), .B(i_1_), .Y(new_new_n427_));
  NOi31      g405(.An(new_new_n427_), .B(new_new_n356_), .C(new_new_n69_), .Y(new_new_n428_));
  NOi21      g406(.An(i_10_), .B(i_6_), .Y(new_new_n429_));
  NO2        g407(.A(new_new_n80_), .B(new_new_n25_), .Y(new_new_n430_));
  AOI220     g408(.A0(new_new_n237_), .A1(new_new_n430_), .B0(new_new_n233_), .B1(new_new_n429_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n431_), .B(new_new_n354_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n109_), .B(new_new_n23_), .Y(new_new_n433_));
  NOi21      g411(.An(new_new_n140_), .B(new_new_n262_), .Y(new_new_n434_));
  NO2        g412(.A(new_new_n434_), .B(new_new_n432_), .Y(new_new_n435_));
  NO2        g413(.A(new_new_n402_), .B(new_new_n301_), .Y(new_new_n436_));
  INV        g414(.A(new_new_n255_), .Y(new_new_n437_));
  NO2        g415(.A(i_12_), .B(new_new_n80_), .Y(new_new_n438_));
  NA3        g416(.A(new_new_n438_), .B(new_new_n233_), .C(new_new_n420_), .Y(new_new_n439_));
  NA3        g417(.A(new_new_n308_), .B(new_new_n237_), .C(new_new_n186_), .Y(new_new_n440_));
  AOI210     g418(.A0(new_new_n440_), .A1(new_new_n439_), .B0(new_new_n437_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n295_), .B(new_new_n205_), .Y(new_new_n442_));
  NO2        g420(.A(new_new_n442_), .B(new_new_n392_), .Y(new_new_n443_));
  NO3        g421(.A(new_new_n443_), .B(new_new_n441_), .C(new_new_n436_), .Y(new_new_n444_));
  NA3        g422(.A(new_new_n444_), .B(new_new_n435_), .C(new_new_n423_), .Y(new_new_n445_));
  NO4        g423(.A(new_new_n445_), .B(new_new_n418_), .C(new_new_n407_), .D(new_new_n398_), .Y(new_new_n446_));
  NA4        g424(.A(new_new_n446_), .B(new_new_n346_), .C(new_new_n274_), .D(new_new_n252_), .Y(ori7));
  NO2        g425(.A(new_new_n88_), .B(new_new_n54_), .Y(new_new_n448_));
  NO2        g426(.A(new_new_n102_), .B(new_new_n85_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n829_), .B(new_new_n449_), .Y(new_new_n450_));
  NA2        g428(.A(new_new_n381_), .B(new_new_n79_), .Y(new_new_n451_));
  NA2        g429(.A(i_11_), .B(new_new_n166_), .Y(new_new_n452_));
  NA2        g430(.A(new_new_n138_), .B(new_new_n452_), .Y(new_new_n453_));
  OAI210     g431(.A0(new_new_n453_), .A1(new_new_n451_), .B0(new_new_n450_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n199_), .B(i_4_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n455_), .B(i_8_), .Y(new_new_n456_));
  NA2        g434(.A(i_2_), .B(new_new_n80_), .Y(new_new_n457_));
  OAI210     g435(.A0(new_new_n83_), .A1(new_new_n172_), .B0(new_new_n173_), .Y(new_new_n458_));
  NO2        g436(.A(i_7_), .B(new_new_n37_), .Y(new_new_n459_));
  NA2        g437(.A(i_4_), .B(i_8_), .Y(new_new_n460_));
  AOI210     g438(.A0(new_new_n460_), .A1(new_new_n248_), .B0(new_new_n459_), .Y(new_new_n461_));
  OAI220     g439(.A0(new_new_n461_), .A1(new_new_n457_), .B0(new_new_n458_), .B1(i_13_), .Y(new_new_n462_));
  NO3        g440(.A(new_new_n462_), .B(new_new_n454_), .C(new_new_n448_), .Y(new_new_n463_));
  AOI210     g441(.A0(new_new_n123_), .A1(new_new_n58_), .B0(i_10_), .Y(new_new_n464_));
  AOI210     g442(.A0(new_new_n464_), .A1(new_new_n199_), .B0(new_new_n148_), .Y(new_new_n465_));
  OR2        g443(.A(i_6_), .B(i_10_), .Y(new_new_n466_));
  INV        g444(.A(new_new_n171_), .Y(new_new_n467_));
  OR2        g445(.A(new_new_n465_), .B(new_new_n226_), .Y(new_new_n468_));
  AOI210     g446(.A0(new_new_n468_), .A1(new_new_n463_), .B0(new_new_n59_), .Y(new_new_n469_));
  NOi21      g447(.An(i_11_), .B(i_7_), .Y(new_new_n470_));
  AO210      g448(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n471_), .B(new_new_n470_), .Y(new_new_n472_));
  NA2        g450(.A(new_new_n472_), .B(new_new_n177_), .Y(new_new_n473_));
  NA3        g451(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n474_));
  NAi31      g452(.An(new_new_n474_), .B(new_new_n183_), .C(i_11_), .Y(new_new_n475_));
  AOI210     g453(.A0(new_new_n475_), .A1(new_new_n473_), .B0(new_new_n59_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n477_));
  AO210      g455(.A0(new_new_n477_), .A1(new_new_n301_), .B0(new_new_n41_), .Y(new_new_n478_));
  NO3        g456(.A(new_new_n216_), .B(new_new_n178_), .C(new_new_n452_), .Y(new_new_n479_));
  OAI210     g457(.A0(new_new_n479_), .A1(new_new_n193_), .B0(new_new_n59_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n332_), .B(new_new_n31_), .Y(new_new_n481_));
  OR2        g459(.A(new_new_n178_), .B(new_new_n102_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n482_), .B(new_new_n481_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n59_), .B(i_9_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n484_), .B(i_4_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n485_), .B(new_new_n483_), .Y(new_new_n486_));
  NO2        g464(.A(i_1_), .B(i_12_), .Y(new_new_n487_));
  NA3        g465(.A(new_new_n487_), .B(new_new_n104_), .C(new_new_n24_), .Y(new_new_n488_));
  BUFFER     g466(.A(new_new_n488_), .Y(new_new_n489_));
  NA4        g467(.A(new_new_n489_), .B(new_new_n486_), .C(new_new_n480_), .D(new_new_n478_), .Y(new_new_n490_));
  OAI210     g468(.A0(new_new_n490_), .A1(new_new_n476_), .B0(i_6_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n474_), .B(new_new_n102_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n492_), .B(new_new_n438_), .Y(new_new_n493_));
  NO2        g471(.A(new_new_n199_), .B(new_new_n80_), .Y(new_new_n494_));
  NO2        g472(.A(new_new_n494_), .B(i_11_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n493_), .B(new_new_n357_), .Y(new_new_n496_));
  NO3        g474(.A(new_new_n466_), .B(new_new_n198_), .C(new_new_n23_), .Y(new_new_n497_));
  AOI210     g475(.A0(i_1_), .A1(new_new_n217_), .B0(new_new_n497_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n498_), .B(new_new_n44_), .Y(new_new_n499_));
  NA3        g477(.A(new_new_n409_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n500_));
  INV        g478(.A(i_2_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n133_), .B(i_9_), .Y(new_new_n502_));
  NA3        g480(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n46_), .B(i_1_), .Y(new_new_n504_));
  NA3        g482(.A(new_new_n504_), .B(new_new_n225_), .C(new_new_n44_), .Y(new_new_n505_));
  OAI220     g483(.A0(new_new_n505_), .A1(new_new_n503_), .B0(new_new_n502_), .B1(new_new_n501_), .Y(new_new_n506_));
  NA3        g484(.A(new_new_n484_), .B(new_new_n255_), .C(i_6_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(new_new_n23_), .Y(new_new_n508_));
  AOI210     g486(.A0(new_new_n377_), .A1(new_new_n335_), .B0(new_new_n203_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n509_), .B(new_new_n457_), .Y(new_new_n510_));
  NO2        g488(.A(i_11_), .B(new_new_n37_), .Y(new_new_n511_));
  OR3        g489(.A(new_new_n510_), .B(new_new_n508_), .C(new_new_n506_), .Y(new_new_n512_));
  NO3        g490(.A(new_new_n512_), .B(new_new_n499_), .C(new_new_n496_), .Y(new_new_n513_));
  NO2        g491(.A(new_new_n199_), .B(new_new_n95_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n514_), .B(new_new_n470_), .Y(new_new_n515_));
  NO2        g493(.A(new_new_n198_), .B(new_new_n44_), .Y(new_new_n516_));
  NO3        g494(.A(new_new_n516_), .B(new_new_n250_), .C(new_new_n200_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n112_), .B(new_new_n37_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n518_), .B(i_6_), .Y(new_new_n519_));
  NO2        g497(.A(new_new_n80_), .B(i_9_), .Y(new_new_n520_));
  NO2        g498(.A(new_new_n520_), .B(new_new_n59_), .Y(new_new_n521_));
  NO2        g499(.A(new_new_n521_), .B(new_new_n487_), .Y(new_new_n522_));
  NO4        g500(.A(new_new_n522_), .B(new_new_n519_), .C(new_new_n517_), .D(i_4_), .Y(new_new_n523_));
  NA2        g501(.A(i_1_), .B(i_3_), .Y(new_new_n524_));
  INV        g502(.A(new_new_n523_), .Y(new_new_n525_));
  NA3        g503(.A(new_new_n525_), .B(new_new_n513_), .C(new_new_n491_), .Y(new_new_n526_));
  NO3        g504(.A(new_new_n378_), .B(i_3_), .C(i_7_), .Y(new_new_n527_));
  NOi21      g505(.An(new_new_n527_), .B(i_10_), .Y(new_new_n528_));
  OA210      g506(.A0(new_new_n528_), .A1(new_new_n206_), .B0(new_new_n80_), .Y(new_new_n529_));
  NA3        g507(.A(new_new_n381_), .B(new_new_n403_), .C(new_new_n46_), .Y(new_new_n530_));
  NO3        g508(.A(new_new_n379_), .B(new_new_n460_), .C(new_new_n80_), .Y(new_new_n531_));
  NA2        g509(.A(new_new_n531_), .B(new_new_n25_), .Y(new_new_n532_));
  NA3        g510(.A(new_new_n148_), .B(new_new_n79_), .C(new_new_n80_), .Y(new_new_n533_));
  NA3        g511(.A(new_new_n533_), .B(new_new_n532_), .C(new_new_n530_), .Y(new_new_n534_));
  OAI210     g512(.A0(new_new_n534_), .A1(new_new_n529_), .B0(i_1_), .Y(new_new_n535_));
  AOI210     g513(.A0(new_new_n225_), .A1(new_new_n93_), .B0(i_1_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n291_), .B(i_2_), .Y(new_new_n537_));
  NA2        g515(.A(new_new_n537_), .B(new_new_n536_), .Y(new_new_n538_));
  OAI210     g516(.A0(new_new_n507_), .A1(new_new_n349_), .B0(new_new_n538_), .Y(new_new_n539_));
  INV        g517(.A(new_new_n539_), .Y(new_new_n540_));
  AOI210     g518(.A0(new_new_n540_), .A1(new_new_n535_), .B0(i_13_), .Y(new_new_n541_));
  NA2        g519(.A(new_new_n100_), .B(new_new_n133_), .Y(new_new_n542_));
  AOI220     g520(.A0(new_new_n373_), .A1(new_new_n148_), .B0(new_new_n351_), .B1(new_new_n133_), .Y(new_new_n543_));
  OAI210     g521(.A0(new_new_n543_), .A1(new_new_n44_), .B0(new_new_n542_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n54_), .B(i_12_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n379_), .B(new_new_n24_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n827_), .B(new_new_n88_), .Y(new_new_n547_));
  AOI210     g525(.A0(new_new_n544_), .A1(new_new_n264_), .B0(new_new_n547_), .Y(new_new_n548_));
  INV        g526(.A(new_new_n109_), .Y(new_new_n549_));
  AOI220     g527(.A0(new_new_n549_), .A1(new_new_n68_), .B0(new_new_n308_), .B1(new_new_n504_), .Y(new_new_n550_));
  NO2        g528(.A(new_new_n550_), .B(new_new_n204_), .Y(new_new_n551_));
  AOI210     g529(.A0(new_new_n349_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n552_));
  NOi31      g530(.An(new_new_n552_), .B(new_new_n451_), .C(new_new_n44_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n122_), .B(i_13_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n503_), .B(new_new_n109_), .Y(new_new_n555_));
  INV        g533(.A(new_new_n555_), .Y(new_new_n556_));
  OAI220     g534(.A0(new_new_n556_), .A1(new_new_n67_), .B0(new_new_n554_), .B1(new_new_n536_), .Y(new_new_n557_));
  NO3        g535(.A(new_new_n67_), .B(new_new_n32_), .C(new_new_n95_), .Y(new_new_n558_));
  NA2        g536(.A(new_new_n26_), .B(new_new_n166_), .Y(new_new_n559_));
  INV        g537(.A(i_7_), .Y(new_new_n560_));
  INV        g538(.A(new_new_n558_), .Y(new_new_n561_));
  AOI220     g539(.A0(new_new_n308_), .A1(new_new_n504_), .B0(new_new_n87_), .B1(new_new_n96_), .Y(new_new_n562_));
  OAI220     g540(.A0(new_new_n562_), .A1(new_new_n456_), .B0(new_new_n561_), .B1(new_new_n467_), .Y(new_new_n563_));
  NO4        g541(.A(new_new_n563_), .B(new_new_n557_), .C(new_new_n553_), .D(new_new_n551_), .Y(new_new_n564_));
  OR2        g542(.A(i_11_), .B(i_6_), .Y(new_new_n565_));
  NA3        g543(.A(new_new_n455_), .B(new_new_n559_), .C(i_7_), .Y(new_new_n566_));
  AOI210     g544(.A0(new_new_n566_), .A1(new_new_n556_), .B0(new_new_n565_), .Y(new_new_n567_));
  NA3        g545(.A(new_new_n332_), .B(new_new_n459_), .C(new_new_n93_), .Y(new_new_n568_));
  NA2        g546(.A(new_new_n495_), .B(i_13_), .Y(new_new_n569_));
  NA2        g547(.A(new_new_n96_), .B(new_new_n559_), .Y(new_new_n570_));
  NAi21      g548(.An(i_11_), .B(i_12_), .Y(new_new_n571_));
  NOi41      g549(.An(new_new_n105_), .B(new_new_n571_), .C(i_13_), .D(new_new_n80_), .Y(new_new_n572_));
  NO3        g550(.A(new_new_n379_), .B(new_new_n438_), .C(new_new_n460_), .Y(new_new_n573_));
  AOI220     g551(.A0(new_new_n573_), .A1(new_new_n253_), .B0(new_new_n572_), .B1(new_new_n570_), .Y(new_new_n574_));
  NA3        g552(.A(new_new_n574_), .B(new_new_n569_), .C(new_new_n568_), .Y(new_new_n575_));
  OAI210     g553(.A0(new_new_n575_), .A1(new_new_n567_), .B0(new_new_n59_), .Y(new_new_n576_));
  NO2        g554(.A(i_2_), .B(i_12_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n290_), .B(new_new_n577_), .Y(new_new_n578_));
  INV        g556(.A(new_new_n578_), .Y(new_new_n579_));
  NA3        g557(.A(new_new_n579_), .B(new_new_n45_), .C(new_new_n192_), .Y(new_new_n580_));
  NA4        g558(.A(new_new_n580_), .B(new_new_n576_), .C(new_new_n564_), .D(new_new_n548_), .Y(new_new_n581_));
  OR4        g559(.A(new_new_n581_), .B(new_new_n541_), .C(new_new_n526_), .D(new_new_n469_), .Y(ori5));
  NA2        g560(.A(new_new_n515_), .B(new_new_n228_), .Y(new_new_n583_));
  AN2        g561(.A(new_new_n24_), .B(i_10_), .Y(new_new_n584_));
  NA3        g562(.A(new_new_n584_), .B(new_new_n577_), .C(new_new_n102_), .Y(new_new_n585_));
  NO2        g563(.A(new_new_n456_), .B(i_11_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n83_), .B(new_new_n586_), .Y(new_new_n587_));
  NA3        g565(.A(new_new_n587_), .B(new_new_n585_), .C(new_new_n583_), .Y(new_new_n588_));
  NO3        g566(.A(i_11_), .B(new_new_n199_), .C(i_13_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n590_));
  NA2        g568(.A(i_12_), .B(i_8_), .Y(new_new_n591_));
  OAI210     g569(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n591_), .Y(new_new_n592_));
  INV        g570(.A(new_new_n348_), .Y(new_new_n593_));
  AOI220     g571(.A0(new_new_n255_), .A1(new_new_n433_), .B0(new_new_n592_), .B1(new_new_n590_), .Y(new_new_n594_));
  INV        g572(.A(new_new_n594_), .Y(new_new_n595_));
  NO2        g573(.A(new_new_n595_), .B(new_new_n588_), .Y(new_new_n596_));
  INV        g574(.A(new_new_n153_), .Y(new_new_n597_));
  INV        g575(.A(new_new_n206_), .Y(new_new_n598_));
  OAI210     g576(.A0(new_new_n537_), .A1(new_new_n350_), .B0(new_new_n105_), .Y(new_new_n599_));
  AOI210     g577(.A0(new_new_n599_), .A1(new_new_n598_), .B0(new_new_n597_), .Y(new_new_n600_));
  NO2        g578(.A(new_new_n358_), .B(new_new_n26_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n601_), .B(new_new_n335_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n602_), .B(i_2_), .Y(new_new_n603_));
  INV        g581(.A(new_new_n603_), .Y(new_new_n604_));
  AOI210     g582(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n333_), .Y(new_new_n605_));
  AOI210     g583(.A0(new_new_n605_), .A1(new_new_n604_), .B0(new_new_n600_), .Y(new_new_n606_));
  NO2        g584(.A(new_new_n165_), .B(new_new_n120_), .Y(new_new_n607_));
  OAI210     g585(.A0(new_new_n607_), .A1(new_new_n590_), .B0(i_2_), .Y(new_new_n608_));
  INV        g586(.A(new_new_n154_), .Y(new_new_n609_));
  NO3        g587(.A(new_new_n471_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n610_));
  AOI210     g588(.A0(new_new_n609_), .A1(new_new_n83_), .B0(new_new_n610_), .Y(new_new_n611_));
  AOI210     g589(.A0(new_new_n611_), .A1(new_new_n608_), .B0(new_new_n166_), .Y(new_new_n612_));
  OA210      g590(.A0(new_new_n472_), .A1(new_new_n121_), .B0(i_13_), .Y(new_new_n613_));
  AOI210     g591(.A0(new_new_n178_), .A1(new_new_n142_), .B0(new_new_n403_), .Y(new_new_n614_));
  NA2        g592(.A(new_new_n614_), .B(new_new_n335_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n96_), .B(new_new_n44_), .Y(new_new_n616_));
  INV        g594(.A(new_new_n247_), .Y(new_new_n617_));
  NA4        g595(.A(new_new_n617_), .B(new_new_n248_), .C(new_new_n119_), .D(new_new_n42_), .Y(new_new_n618_));
  OAI210     g596(.A0(new_new_n618_), .A1(new_new_n616_), .B0(new_new_n615_), .Y(new_new_n619_));
  NO3        g597(.A(new_new_n619_), .B(new_new_n613_), .C(new_new_n612_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n433_), .B(new_new_n28_), .Y(new_new_n621_));
  NA2        g599(.A(new_new_n589_), .B(new_new_n234_), .Y(new_new_n622_));
  NA2        g600(.A(new_new_n622_), .B(new_new_n621_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n58_), .B(i_12_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n624_), .B(new_new_n121_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n452_), .Y(new_new_n626_));
  AOI220     g604(.A0(new_new_n626_), .A1(new_new_n36_), .B0(new_new_n623_), .B1(new_new_n46_), .Y(new_new_n627_));
  NA4        g605(.A(new_new_n627_), .B(new_new_n620_), .C(new_new_n606_), .D(new_new_n596_), .Y(ori6));
  NA4        g606(.A(new_new_n311_), .B(new_new_n380_), .C(new_new_n67_), .D(new_new_n95_), .Y(new_new_n629_));
  INV        g607(.A(new_new_n629_), .Y(new_new_n630_));
  NO2        g608(.A(new_new_n188_), .B(new_new_n383_), .Y(new_new_n631_));
  NO2        g609(.A(i_11_), .B(i_9_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n630_), .B(new_new_n259_), .Y(new_new_n633_));
  OR2        g611(.A(new_new_n633_), .B(i_12_), .Y(new_new_n634_));
  NA2        g612(.A(new_new_n296_), .B(new_new_n267_), .Y(new_new_n635_));
  NA2        g613(.A(new_new_n438_), .B(new_new_n59_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n528_), .B(new_new_n67_), .Y(new_new_n637_));
  BUFFER     g615(.A(new_new_n477_), .Y(new_new_n638_));
  NA4        g616(.A(new_new_n638_), .B(new_new_n637_), .C(new_new_n636_), .D(new_new_n635_), .Y(new_new_n639_));
  INV        g617(.A(new_new_n169_), .Y(new_new_n640_));
  AOI220     g618(.A0(new_new_n640_), .A1(new_new_n632_), .B0(new_new_n639_), .B1(new_new_n69_), .Y(new_new_n641_));
  INV        g619(.A(new_new_n258_), .Y(new_new_n642_));
  NA2        g620(.A(new_new_n71_), .B(new_new_n126_), .Y(new_new_n643_));
  INV        g621(.A(new_new_n119_), .Y(new_new_n644_));
  NA2        g622(.A(new_new_n644_), .B(new_new_n46_), .Y(new_new_n645_));
  AOI210     g623(.A0(new_new_n645_), .A1(new_new_n643_), .B0(new_new_n642_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n32_), .B(i_11_), .Y(new_new_n647_));
  NA3        g625(.A(new_new_n647_), .B(new_new_n376_), .C(new_new_n311_), .Y(new_new_n648_));
  NAi32      g626(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n565_), .B(new_new_n649_), .Y(new_new_n650_));
  OAI210     g628(.A0(new_new_n527_), .A1(new_new_n426_), .B0(new_new_n425_), .Y(new_new_n651_));
  NAi31      g629(.An(new_new_n650_), .B(new_new_n651_), .C(new_new_n648_), .Y(new_new_n652_));
  OR2        g630(.A(new_new_n652_), .B(new_new_n646_), .Y(new_new_n653_));
  AO220      g631(.A0(new_new_n279_), .A1(new_new_n270_), .B0(new_new_n319_), .B1(new_new_n452_), .Y(new_new_n654_));
  NA3        g632(.A(new_new_n654_), .B(new_new_n213_), .C(i_7_), .Y(new_new_n655_));
  BUFFER     g633(.A(new_new_n472_), .Y(new_new_n656_));
  NA3        g634(.A(new_new_n656_), .B(new_new_n141_), .C(new_new_n65_), .Y(new_new_n657_));
  AO210      g635(.A0(new_new_n390_), .A1(new_new_n593_), .B0(new_new_n36_), .Y(new_new_n658_));
  NA3        g636(.A(new_new_n658_), .B(new_new_n657_), .C(new_new_n655_), .Y(new_new_n659_));
  OAI210     g637(.A0(new_new_n494_), .A1(i_11_), .B0(new_new_n81_), .Y(new_new_n660_));
  AOI220     g638(.A0(new_new_n660_), .A1(new_new_n425_), .B0(new_new_n631_), .B1(new_new_n560_), .Y(new_new_n661_));
  NA3        g639(.A(new_new_n295_), .B(new_new_n201_), .C(new_new_n141_), .Y(new_new_n662_));
  NA2        g640(.A(new_new_n319_), .B(new_new_n66_), .Y(new_new_n663_));
  NA4        g641(.A(new_new_n663_), .B(new_new_n662_), .C(new_new_n661_), .D(new_new_n458_), .Y(new_new_n664_));
  AO210      g642(.A0(new_new_n403_), .A1(new_new_n46_), .B0(new_new_n82_), .Y(new_new_n665_));
  NA3        g643(.A(new_new_n665_), .B(new_new_n381_), .C(new_new_n186_), .Y(new_new_n666_));
  AOI210     g644(.A0(new_new_n350_), .A1(new_new_n348_), .B0(new_new_n424_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n466_), .B(new_new_n96_), .Y(new_new_n668_));
  OAI210     g646(.A0(new_new_n668_), .A1(new_new_n106_), .B0(new_new_n331_), .Y(new_new_n669_));
  NA2        g647(.A(new_new_n205_), .B(new_new_n46_), .Y(new_new_n670_));
  NA3        g648(.A(new_new_n669_), .B(new_new_n667_), .C(new_new_n666_), .Y(new_new_n671_));
  NO4        g649(.A(new_new_n671_), .B(new_new_n664_), .C(new_new_n659_), .D(new_new_n653_), .Y(new_new_n672_));
  NA4        g650(.A(new_new_n672_), .B(new_new_n641_), .C(new_new_n634_), .D(new_new_n303_), .Y(ori3));
  NA2        g651(.A(i_12_), .B(i_10_), .Y(new_new_n674_));
  NO2        g652(.A(i_11_), .B(new_new_n199_), .Y(new_new_n675_));
  NA3        g653(.A(new_new_n662_), .B(new_new_n458_), .C(new_new_n294_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n676_), .B(new_new_n40_), .Y(new_new_n677_));
  NOi21      g655(.An(new_new_n92_), .B(new_new_n602_), .Y(new_new_n678_));
  NO3        g656(.A(new_new_n482_), .B(new_new_n358_), .C(new_new_n126_), .Y(new_new_n679_));
  NA2        g657(.A(new_new_n332_), .B(new_new_n45_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n679_), .B(new_new_n678_), .Y(new_new_n681_));
  AOI210     g659(.A0(new_new_n681_), .A1(new_new_n677_), .B0(new_new_n48_), .Y(new_new_n682_));
  NO4        g660(.A(new_new_n299_), .B(new_new_n306_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n160_), .B(new_new_n429_), .Y(new_new_n684_));
  NOi21      g662(.An(new_new_n684_), .B(new_new_n683_), .Y(new_new_n685_));
  NO2        g663(.A(new_new_n685_), .B(new_new_n59_), .Y(new_new_n686_));
  NOi21      g664(.An(i_5_), .B(i_9_), .Y(new_new_n687_));
  NA2        g665(.A(new_new_n687_), .B(new_new_n347_), .Y(new_new_n688_));
  BUFFER     g666(.A(new_new_n225_), .Y(new_new_n689_));
  AOI210     g667(.A0(new_new_n689_), .A1(new_new_n377_), .B0(new_new_n531_), .Y(new_new_n690_));
  NO2        g668(.A(new_new_n690_), .B(new_new_n688_), .Y(new_new_n691_));
  NO3        g669(.A(new_new_n691_), .B(new_new_n686_), .C(new_new_n682_), .Y(new_new_n692_));
  NA2        g670(.A(new_new_n160_), .B(new_new_n24_), .Y(new_new_n693_));
  NO2        g671(.A(new_new_n518_), .B(new_new_n449_), .Y(new_new_n694_));
  NO2        g672(.A(new_new_n694_), .B(new_new_n693_), .Y(new_new_n695_));
  NA2        g673(.A(new_new_n253_), .B(new_new_n124_), .Y(new_new_n696_));
  NAi21      g674(.An(new_new_n149_), .B(new_new_n340_), .Y(new_new_n697_));
  OAI220     g675(.A0(new_new_n697_), .A1(new_new_n670_), .B0(new_new_n696_), .B1(new_new_n324_), .Y(new_new_n698_));
  NO2        g676(.A(new_new_n698_), .B(new_new_n695_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n430_), .B(i_0_), .Y(new_new_n700_));
  NO3        g678(.A(new_new_n700_), .B(new_new_n307_), .C(new_new_n83_), .Y(new_new_n701_));
  INV        g679(.A(new_new_n701_), .Y(new_new_n702_));
  NA2        g680(.A(new_new_n589_), .B(new_new_n259_), .Y(new_new_n703_));
  AOI210     g681(.A0(new_new_n381_), .A1(new_new_n83_), .B0(new_new_n56_), .Y(new_new_n704_));
  NO2        g682(.A(new_new_n704_), .B(new_new_n703_), .Y(new_new_n705_));
  NA2        g683(.A(i_0_), .B(i_10_), .Y(new_new_n706_));
  INV        g684(.A(new_new_n705_), .Y(new_new_n707_));
  NA3        g685(.A(new_new_n707_), .B(new_new_n702_), .C(new_new_n699_), .Y(new_new_n708_));
  NO2        g686(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n709_));
  NA2        g687(.A(i_11_), .B(i_9_), .Y(new_new_n710_));
  NO3        g688(.A(i_12_), .B(new_new_n710_), .C(new_new_n457_), .Y(new_new_n711_));
  AN2        g689(.A(new_new_n711_), .B(new_new_n709_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n316_), .B(new_new_n158_), .Y(new_new_n713_));
  INV        g691(.A(new_new_n713_), .Y(new_new_n714_));
  NO2        g692(.A(new_new_n710_), .B(new_new_n69_), .Y(new_new_n715_));
  NO2        g693(.A(new_new_n156_), .B(i_0_), .Y(new_new_n716_));
  INV        g694(.A(new_new_n330_), .Y(new_new_n717_));
  NO2        g695(.A(new_new_n717_), .B(new_new_n688_), .Y(new_new_n718_));
  NO3        g696(.A(new_new_n718_), .B(new_new_n714_), .C(new_new_n712_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n511_), .B(new_new_n116_), .Y(new_new_n720_));
  NO2        g698(.A(i_6_), .B(new_new_n720_), .Y(new_new_n721_));
  NA2        g699(.A(new_new_n153_), .B(new_new_n97_), .Y(new_new_n722_));
  NA2        g700(.A(new_new_n459_), .B(new_new_n259_), .Y(new_new_n723_));
  NO2        g701(.A(new_new_n723_), .B(new_new_n680_), .Y(new_new_n724_));
  NO2        g702(.A(new_new_n724_), .B(new_new_n721_), .Y(new_new_n725_));
  NOi21      g703(.An(i_7_), .B(i_5_), .Y(new_new_n726_));
  NOi31      g704(.An(new_new_n726_), .B(i_0_), .C(new_new_n571_), .Y(new_new_n727_));
  NA3        g705(.A(new_new_n727_), .B(new_new_n829_), .C(i_6_), .Y(new_new_n728_));
  BUFFER     g706(.A(new_new_n728_), .Y(new_new_n729_));
  INV        g707(.A(new_new_n256_), .Y(new_new_n730_));
  NA3        g708(.A(new_new_n729_), .B(new_new_n725_), .C(new_new_n719_), .Y(new_new_n731_));
  NO2        g709(.A(new_new_n674_), .B(new_new_n255_), .Y(new_new_n732_));
  OA210      g710(.A0(new_new_n376_), .A1(new_new_n190_), .B0(new_new_n375_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n732_), .B(new_new_n715_), .Y(new_new_n734_));
  NA3        g712(.A(new_new_n375_), .B(new_new_n332_), .C(new_new_n45_), .Y(new_new_n735_));
  OAI210     g713(.A0(new_new_n697_), .A1(i_7_), .B0(new_new_n735_), .Y(new_new_n736_));
  NA2        g714(.A(new_new_n715_), .B(new_new_n248_), .Y(new_new_n737_));
  OAI210     g715(.A0(i_3_), .A1(new_new_n162_), .B0(new_new_n737_), .Y(new_new_n738_));
  AOI220     g716(.A0(new_new_n738_), .A1(new_new_n376_), .B0(new_new_n736_), .B1(new_new_n69_), .Y(new_new_n739_));
  NA3        g717(.A(i_5_), .B(new_new_n305_), .C(new_new_n494_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n88_), .B(new_new_n44_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n71_), .B(new_new_n591_), .Y(new_new_n742_));
  AOI220     g720(.A0(new_new_n742_), .A1(new_new_n741_), .B0(new_new_n155_), .B1(new_new_n449_), .Y(new_new_n743_));
  AOI210     g721(.A0(new_new_n743_), .A1(new_new_n740_), .B0(new_new_n47_), .Y(new_new_n744_));
  NO3        g722(.A(i_5_), .B(new_new_n277_), .C(new_new_n24_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n546_), .A1(new_new_n414_), .B0(new_new_n745_), .Y(new_new_n746_));
  NAi21      g724(.An(i_9_), .B(i_5_), .Y(new_new_n747_));
  NO2        g725(.A(new_new_n747_), .B(new_new_n325_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n748_), .B(new_new_n472_), .Y(new_new_n749_));
  OAI220     g727(.A0(new_new_n749_), .A1(new_new_n80_), .B0(new_new_n746_), .B1(new_new_n154_), .Y(new_new_n750_));
  NO2        g728(.A(new_new_n750_), .B(new_new_n744_), .Y(new_new_n751_));
  NA3        g729(.A(new_new_n751_), .B(new_new_n739_), .C(new_new_n734_), .Y(new_new_n752_));
  NO3        g730(.A(new_new_n752_), .B(new_new_n731_), .C(new_new_n708_), .Y(new_new_n753_));
  NO2        g731(.A(i_0_), .B(new_new_n571_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n636_), .B(new_new_n722_), .Y(new_new_n755_));
  INV        g733(.A(new_new_n755_), .Y(new_new_n756_));
  NO2        g734(.A(new_new_n651_), .B(new_new_n325_), .Y(new_new_n757_));
  NA2        g735(.A(new_new_n205_), .B(new_new_n197_), .Y(new_new_n758_));
  AOI210     g736(.A0(new_new_n758_), .A1(new_new_n700_), .B0(new_new_n145_), .Y(new_new_n759_));
  NO2        g737(.A(new_new_n759_), .B(new_new_n757_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n760_), .B(new_new_n756_), .Y(new_new_n761_));
  NO3        g739(.A(new_new_n706_), .B(new_new_n687_), .C(new_new_n165_), .Y(new_new_n762_));
  AOI220     g740(.A0(new_new_n762_), .A1(i_11_), .B0(new_new_n428_), .B1(new_new_n71_), .Y(new_new_n763_));
  NO3        g741(.A(new_new_n179_), .B(new_new_n306_), .C(i_0_), .Y(new_new_n764_));
  OAI210     g742(.A0(new_new_n764_), .A1(new_new_n72_), .B0(i_13_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n765_), .B(new_new_n763_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n204_), .B(new_new_n88_), .Y(new_new_n767_));
  AOI210     g745(.A0(new_new_n767_), .A1(new_new_n754_), .B0(new_new_n103_), .Y(new_new_n768_));
  OR2        g746(.A(new_new_n768_), .B(i_5_), .Y(new_new_n769_));
  AOI210     g747(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n156_), .Y(new_new_n770_));
  NA2        g748(.A(new_new_n770_), .B(new_new_n733_), .Y(new_new_n771_));
  NO3        g749(.A(new_new_n680_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n772_));
  NA2        g750(.A(new_new_n389_), .B(new_new_n382_), .Y(new_new_n773_));
  NO2        g751(.A(new_new_n773_), .B(new_new_n772_), .Y(new_new_n774_));
  NA3        g752(.A(new_new_n311_), .B(new_new_n153_), .C(new_new_n152_), .Y(new_new_n775_));
  NA3        g753(.A(i_5_), .B(new_new_n240_), .C(new_new_n197_), .Y(new_new_n776_));
  NA2        g754(.A(new_new_n776_), .B(new_new_n775_), .Y(new_new_n777_));
  NA3        g755(.A(new_new_n311_), .B(new_new_n266_), .C(new_new_n189_), .Y(new_new_n778_));
  INV        g756(.A(new_new_n778_), .Y(new_new_n779_));
  NO3        g757(.A(new_new_n710_), .B(new_new_n186_), .C(new_new_n165_), .Y(new_new_n780_));
  NO3        g758(.A(new_new_n780_), .B(new_new_n779_), .C(new_new_n777_), .Y(new_new_n781_));
  NA4        g759(.A(new_new_n781_), .B(new_new_n774_), .C(new_new_n771_), .D(new_new_n769_), .Y(new_new_n782_));
  NO2        g760(.A(new_new_n80_), .B(i_5_), .Y(new_new_n783_));
  NA3        g761(.A(new_new_n675_), .B(new_new_n104_), .C(new_new_n119_), .Y(new_new_n784_));
  INV        g762(.A(new_new_n784_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n785_), .B(new_new_n783_), .Y(new_new_n786_));
  NA3        g764(.A(new_new_n248_), .B(i_5_), .C(new_new_n166_), .Y(new_new_n787_));
  NAi31      g765(.An(new_new_n203_), .B(new_new_n787_), .C(new_new_n204_), .Y(new_new_n788_));
  NO4        g766(.A(new_new_n202_), .B(new_new_n179_), .C(i_0_), .D(i_12_), .Y(new_new_n789_));
  AOI220     g767(.A0(new_new_n789_), .A1(new_new_n788_), .B0(new_new_n630_), .B1(new_new_n157_), .Y(new_new_n790_));
  AN2        g768(.A(new_new_n706_), .B(new_new_n145_), .Y(new_new_n791_));
  NO4        g769(.A(new_new_n791_), .B(i_12_), .C(new_new_n500_), .D(new_new_n126_), .Y(new_new_n792_));
  NA2        g770(.A(new_new_n792_), .B(new_new_n186_), .Y(new_new_n793_));
  NA2        g771(.A(new_new_n726_), .B(new_new_n373_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n60_), .B(new_new_n95_), .Y(new_new_n795_));
  OAI220     g773(.A0(new_new_n795_), .A1(new_new_n787_), .B0(new_new_n794_), .B1(new_new_n521_), .Y(new_new_n796_));
  NA2        g774(.A(new_new_n796_), .B(new_new_n716_), .Y(new_new_n797_));
  NA4        g775(.A(new_new_n797_), .B(new_new_n793_), .C(new_new_n790_), .D(new_new_n786_), .Y(new_new_n798_));
  NO4        g776(.A(new_new_n798_), .B(new_new_n782_), .C(new_new_n766_), .D(new_new_n761_), .Y(new_new_n799_));
  NA2        g777(.A(new_new_n647_), .B(new_new_n37_), .Y(new_new_n800_));
  NA2        g778(.A(new_new_n800_), .B(new_new_n465_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n801_), .B(new_new_n177_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n497_), .B(new_new_n48_), .Y(new_new_n803_));
  AOI210     g781(.A0(new_new_n803_), .A1(new_new_n802_), .B0(new_new_n69_), .Y(new_new_n804_));
  INV        g782(.A(new_new_n302_), .Y(new_new_n805_));
  NO2        g783(.A(new_new_n805_), .B(new_new_n597_), .Y(new_new_n806_));
  INV        g784(.A(new_new_n72_), .Y(new_new_n807_));
  AOI210     g785(.A0(new_new_n770_), .A1(i_5_), .B0(new_new_n727_), .Y(new_new_n808_));
  AOI210     g786(.A0(new_new_n808_), .A1(new_new_n807_), .B0(new_new_n524_), .Y(new_new_n809_));
  INV        g787(.A(new_new_n809_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n227_), .B(new_new_n83_), .Y(new_new_n811_));
  NA3        g789(.A(new_new_n601_), .B(new_new_n240_), .C(new_new_n76_), .Y(new_new_n812_));
  AOI210     g790(.A0(new_new_n812_), .A1(new_new_n811_), .B0(i_11_), .Y(new_new_n813_));
  NO3        g791(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n814_));
  OAI210     g792(.A0(new_new_n730_), .A1(new_new_n249_), .B0(new_new_n814_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n815_), .B(new_new_n571_), .Y(new_new_n816_));
  NO4        g794(.A(new_new_n747_), .B(new_new_n378_), .C(new_new_n210_), .D(new_new_n209_), .Y(new_new_n817_));
  NO2        g795(.A(new_new_n817_), .B(new_new_n424_), .Y(new_new_n818_));
  INV        g796(.A(new_new_n283_), .Y(new_new_n819_));
  AOI210     g797(.A0(new_new_n819_), .A1(new_new_n818_), .B0(new_new_n41_), .Y(new_new_n820_));
  NO3        g798(.A(new_new_n820_), .B(new_new_n816_), .C(new_new_n813_), .Y(new_new_n821_));
  OAI210     g799(.A0(new_new_n810_), .A1(i_4_), .B0(new_new_n821_), .Y(new_new_n822_));
  NO3        g800(.A(new_new_n822_), .B(new_new_n806_), .C(new_new_n804_), .Y(new_new_n823_));
  NA4        g801(.A(new_new_n823_), .B(new_new_n799_), .C(new_new_n753_), .D(new_new_n692_), .Y(ori4));
  INV        g802(.A(new_new_n545_), .Y(new_new_n827_));
  INV        g803(.A(i_6_), .Y(new_new_n828_));
  INV        g804(.A(i_4_), .Y(new_new_n829_));
endmodule


