// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n133_, new_new_n134_, new_new_n135_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1022_, new_new_n1023_,
    new_new_n1024_, new_new_n1025_, new_new_n1026_, new_new_n1027_,
    new_new_n1028_, new_new_n1029_, new_new_n1030_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g0016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g0017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g0018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(men1));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g0028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g0029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g0032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  INV        g0037(.A(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(new_new_n65_), .B(new_new_n61_), .Y(new_new_n66_));
  NA2        g0044(.A(new_new_n50_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g0046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g0047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g0048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g0049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g0050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g0051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g0052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  OAI210     g0053(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n75_), .Y(new_new_n76_));
  OAI210     g0054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g0055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g0056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g0057(.A(i_3_), .B(i_9_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_7_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n63_), .Y(new_new_n82_));
  INV        g0060(.A(i_6_), .Y(new_new_n83_));
  OR4        g0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n84_));
  NO2        g0062(.A(i_2_), .B(i_7_), .Y(new_new_n85_));
  NA2        g0063(.A(new_new_n82_), .B(new_new_n84_), .Y(new_new_n86_));
  NAi21      g0064(.An(i_6_), .B(i_10_), .Y(new_new_n87_));
  NA2        g0065(.A(i_6_), .B(i_9_), .Y(new_new_n88_));
  NO2        g0066(.A(new_new_n87_), .B(new_new_n63_), .Y(new_new_n89_));
  NA2        g0067(.A(i_2_), .B(i_6_), .Y(new_new_n90_));
  NO3        g0068(.A(new_new_n90_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n91_));
  INV        g0069(.A(new_new_n91_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n92_), .A1(new_new_n86_), .B0(new_new_n78_), .Y(new_new_n93_));
  AN3        g0071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n94_));
  NAi21      g0072(.An(i_6_), .B(i_11_), .Y(new_new_n95_));
  NO2        g0073(.A(i_5_), .B(i_8_), .Y(new_new_n96_));
  NOi21      g0074(.An(new_new_n96_), .B(new_new_n95_), .Y(new_new_n97_));
  NA2        g0075(.A(new_new_n94_), .B(new_new_n32_), .Y(new_new_n98_));
  INV        g0076(.A(i_7_), .Y(new_new_n99_));
  NO2        g0077(.A(i_0_), .B(i_5_), .Y(new_new_n100_));
  NO2        g0078(.A(new_new_n100_), .B(new_new_n83_), .Y(new_new_n101_));
  NA2        g0079(.A(i_12_), .B(i_3_), .Y(new_new_n102_));
  INV        g0080(.A(new_new_n102_), .Y(new_new_n103_));
  NAi21      g0081(.An(i_7_), .B(i_11_), .Y(new_new_n104_));
  NO3        g0082(.A(new_new_n104_), .B(new_new_n87_), .C(new_new_n53_), .Y(new_new_n105_));
  AN2        g0083(.A(i_2_), .B(i_10_), .Y(new_new_n106_));
  NO2        g0084(.A(new_new_n106_), .B(i_7_), .Y(new_new_n107_));
  OR2        g0085(.A(new_new_n78_), .B(new_new_n58_), .Y(new_new_n108_));
  NO2        g0086(.A(i_8_), .B(new_new_n99_), .Y(new_new_n109_));
  NO3        g0087(.A(new_new_n109_), .B(new_new_n108_), .C(new_new_n107_), .Y(new_new_n110_));
  NA2        g0088(.A(i_12_), .B(i_7_), .Y(new_new_n111_));
  NA2        g0089(.A(i_1_), .B(i_0_), .Y(new_new_n112_));
  NA2        g0090(.A(i_11_), .B(i_12_), .Y(new_new_n113_));
  OAI210     g0091(.A0(new_new_n112_), .A1(new_new_n111_), .B0(new_new_n113_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n114_), .B(new_new_n110_), .Y(new_new_n115_));
  NAi31      g0093(.An(new_new_n105_), .B(new_new_n115_), .C(new_new_n98_), .Y(new_new_n116_));
  NOi21      g0094(.An(i_1_), .B(i_5_), .Y(new_new_n117_));
  NA2        g0095(.A(new_new_n117_), .B(i_11_), .Y(new_new_n118_));
  NA2        g0096(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n119_));
  NA2        g0097(.A(i_7_), .B(new_new_n25_), .Y(new_new_n120_));
  NA2        g0098(.A(new_new_n120_), .B(new_new_n119_), .Y(new_new_n121_));
  NO2        g0099(.A(new_new_n121_), .B(new_new_n46_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n88_), .B(new_new_n87_), .Y(new_new_n123_));
  NAi21      g0101(.An(i_3_), .B(i_8_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(new_new_n62_), .Y(new_new_n125_));
  NOi31      g0103(.An(new_new_n125_), .B(new_new_n123_), .C(new_new_n122_), .Y(new_new_n126_));
  NO2        g0104(.A(i_1_), .B(new_new_n83_), .Y(new_new_n127_));
  NO2        g0105(.A(i_6_), .B(i_5_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(i_3_), .Y(new_new_n129_));
  NO2        g0107(.A(new_new_n126_), .B(new_new_n118_), .Y(new_new_n130_));
  NO3        g0108(.A(new_new_n130_), .B(new_new_n116_), .C(new_new_n93_), .Y(new_new_n131_));
  NA3        g0109(.A(new_new_n131_), .B(new_new_n77_), .C(new_new_n56_), .Y(men2));
  NO2        g0110(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n133_));
  INV        g0111(.A(i_6_), .Y(new_new_n134_));
  NA2        g0112(.A(new_new_n134_), .B(new_new_n133_), .Y(new_new_n135_));
  NA4        g0113(.A(new_new_n135_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(men0));
  AN2        g0114(.A(i_8_), .B(i_7_), .Y(new_new_n137_));
  NA2        g0115(.A(new_new_n137_), .B(i_6_), .Y(new_new_n138_));
  NO2        g0116(.A(i_12_), .B(i_13_), .Y(new_new_n139_));
  NAi21      g0117(.An(i_5_), .B(i_11_), .Y(new_new_n140_));
  NOi21      g0118(.An(new_new_n139_), .B(new_new_n140_), .Y(new_new_n141_));
  NO2        g0119(.A(i_0_), .B(i_1_), .Y(new_new_n142_));
  NA2        g0120(.A(i_2_), .B(i_3_), .Y(new_new_n143_));
  NO2        g0121(.A(new_new_n143_), .B(i_4_), .Y(new_new_n144_));
  NA3        g0122(.A(new_new_n144_), .B(new_new_n142_), .C(new_new_n141_), .Y(new_new_n145_));
  OR2        g0123(.A(new_new_n145_), .B(new_new_n25_), .Y(new_new_n146_));
  AN2        g0124(.A(new_new_n139_), .B(new_new_n80_), .Y(new_new_n147_));
  NO2        g0125(.A(new_new_n147_), .B(new_new_n27_), .Y(new_new_n148_));
  NA2        g0126(.A(i_1_), .B(i_5_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n71_), .B(new_new_n46_), .Y(new_new_n150_));
  NA2        g0128(.A(new_new_n150_), .B(new_new_n36_), .Y(new_new_n151_));
  NO3        g0129(.A(new_new_n151_), .B(new_new_n149_), .C(new_new_n148_), .Y(new_new_n152_));
  OR2        g0130(.A(i_0_), .B(i_1_), .Y(new_new_n153_));
  NO3        g0131(.A(new_new_n153_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n154_));
  NAi32      g0132(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n155_));
  NAi21      g0133(.An(new_new_n155_), .B(new_new_n154_), .Y(new_new_n156_));
  NOi21      g0134(.An(i_4_), .B(i_10_), .Y(new_new_n157_));
  NA2        g0135(.A(new_new_n157_), .B(new_new_n39_), .Y(new_new_n158_));
  NO2        g0136(.A(i_3_), .B(i_5_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n71_), .B(i_2_), .C(i_1_), .Y(new_new_n160_));
  OAI210     g0138(.A0(i_2_), .A1(new_new_n158_), .B0(new_new_n156_), .Y(new_new_n161_));
  NO2        g0139(.A(new_new_n161_), .B(new_new_n152_), .Y(new_new_n162_));
  AOI210     g0140(.A0(new_new_n162_), .A1(new_new_n146_), .B0(new_new_n138_), .Y(new_new_n163_));
  NOi21      g0141(.An(i_4_), .B(i_9_), .Y(new_new_n164_));
  NOi21      g0142(.An(i_11_), .B(i_13_), .Y(new_new_n165_));
  NA2        g0143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  NO2        g0144(.A(i_4_), .B(i_5_), .Y(new_new_n167_));
  NAi21      g0145(.An(i_12_), .B(i_11_), .Y(new_new_n168_));
  NO2        g0146(.A(new_new_n168_), .B(i_13_), .Y(new_new_n169_));
  NA3        g0147(.A(new_new_n169_), .B(new_new_n167_), .C(new_new_n80_), .Y(new_new_n170_));
  AOI210     g0148(.A0(new_new_n170_), .A1(new_new_n166_), .B0(i_2_), .Y(new_new_n171_));
  NO2        g0149(.A(new_new_n71_), .B(new_new_n63_), .Y(new_new_n172_));
  NA2        g0150(.A(new_new_n172_), .B(new_new_n46_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n36_), .B(i_5_), .Y(new_new_n174_));
  NAi31      g0152(.An(new_new_n174_), .B(new_new_n147_), .C(i_11_), .Y(new_new_n175_));
  NA2        g0153(.A(i_3_), .B(i_5_), .Y(new_new_n176_));
  AOI210     g0154(.A0(new_new_n166_), .A1(new_new_n175_), .B0(new_new_n173_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n71_), .B(i_5_), .Y(new_new_n178_));
  NO2        g0156(.A(i_13_), .B(i_10_), .Y(new_new_n179_));
  NA3        g0157(.A(new_new_n179_), .B(new_new_n178_), .C(new_new_n44_), .Y(new_new_n180_));
  NO2        g0158(.A(i_2_), .B(i_1_), .Y(new_new_n181_));
  NA2        g0159(.A(new_new_n181_), .B(i_3_), .Y(new_new_n182_));
  NAi21      g0160(.An(i_4_), .B(i_12_), .Y(new_new_n183_));
  NO4        g0161(.A(new_new_n183_), .B(new_new_n182_), .C(new_new_n180_), .D(new_new_n25_), .Y(new_new_n184_));
  NO3        g0162(.A(new_new_n184_), .B(new_new_n177_), .C(new_new_n171_), .Y(new_new_n185_));
  INV        g0163(.A(i_8_), .Y(new_new_n186_));
  NO2        g0164(.A(new_new_n186_), .B(i_7_), .Y(new_new_n187_));
  NA2        g0165(.A(new_new_n187_), .B(i_6_), .Y(new_new_n188_));
  NO3        g0166(.A(i_3_), .B(new_new_n83_), .C(new_new_n48_), .Y(new_new_n189_));
  NA2        g0167(.A(new_new_n189_), .B(new_new_n109_), .Y(new_new_n190_));
  NO3        g0168(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n191_));
  NA3        g0169(.A(new_new_n191_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n192_));
  NO3        g0170(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n193_));
  OAI210     g0171(.A0(new_new_n94_), .A1(i_12_), .B0(new_new_n193_), .Y(new_new_n194_));
  AOI210     g0172(.A0(new_new_n194_), .A1(new_new_n192_), .B0(new_new_n190_), .Y(new_new_n195_));
  NO2        g0173(.A(i_3_), .B(i_8_), .Y(new_new_n196_));
  NO3        g0174(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n197_));
  NA3        g0175(.A(new_new_n197_), .B(new_new_n196_), .C(new_new_n39_), .Y(new_new_n198_));
  NO2        g0176(.A(new_new_n100_), .B(new_new_n58_), .Y(new_new_n199_));
  NO2        g0177(.A(i_13_), .B(i_9_), .Y(new_new_n200_));
  NA3        g0178(.A(new_new_n200_), .B(i_6_), .C(new_new_n186_), .Y(new_new_n201_));
  NAi21      g0179(.An(i_12_), .B(i_3_), .Y(new_new_n202_));
  OR2        g0180(.A(new_new_n202_), .B(new_new_n201_), .Y(new_new_n203_));
  NO2        g0181(.A(new_new_n44_), .B(i_5_), .Y(new_new_n204_));
  NO3        g0182(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n205_));
  OAI220     g0183(.A0(i_2_), .A1(new_new_n203_), .B0(new_new_n100_), .B1(new_new_n198_), .Y(new_new_n206_));
  AOI210     g0184(.A0(new_new_n206_), .A1(i_7_), .B0(new_new_n195_), .Y(new_new_n207_));
  OAI220     g0185(.A0(new_new_n207_), .A1(i_4_), .B0(new_new_n188_), .B1(new_new_n185_), .Y(new_new_n208_));
  NAi21      g0186(.An(i_12_), .B(i_7_), .Y(new_new_n209_));
  NA3        g0187(.A(i_13_), .B(new_new_n186_), .C(i_10_), .Y(new_new_n210_));
  NO2        g0188(.A(new_new_n210_), .B(new_new_n209_), .Y(new_new_n211_));
  NA2        g0189(.A(i_0_), .B(i_5_), .Y(new_new_n212_));
  NA2        g0190(.A(new_new_n212_), .B(new_new_n101_), .Y(new_new_n213_));
  OAI220     g0191(.A0(new_new_n213_), .A1(new_new_n182_), .B0(new_new_n173_), .B1(new_new_n129_), .Y(new_new_n214_));
  NAi31      g0192(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n215_));
  NO2        g0193(.A(new_new_n36_), .B(i_13_), .Y(new_new_n216_));
  NO2        g0194(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n218_));
  NA3        g0196(.A(new_new_n218_), .B(new_new_n217_), .C(new_new_n216_), .Y(new_new_n219_));
  INV        g0197(.A(i_13_), .Y(new_new_n220_));
  NO2        g0198(.A(i_12_), .B(new_new_n220_), .Y(new_new_n221_));
  NA3        g0199(.A(new_new_n221_), .B(new_new_n191_), .C(new_new_n189_), .Y(new_new_n222_));
  OAI210     g0200(.A0(new_new_n219_), .A1(new_new_n215_), .B0(new_new_n222_), .Y(new_new_n223_));
  AOI220     g0201(.A0(new_new_n223_), .A1(new_new_n137_), .B0(new_new_n214_), .B1(new_new_n211_), .Y(new_new_n224_));
  NO2        g0202(.A(i_12_), .B(new_new_n37_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n176_), .B(i_4_), .Y(new_new_n226_));
  INV        g0204(.A(new_new_n226_), .Y(new_new_n227_));
  OR2        g0205(.A(i_8_), .B(i_7_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n228_), .B(new_new_n83_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n53_), .B(i_1_), .Y(new_new_n230_));
  NA2        g0208(.A(new_new_n230_), .B(new_new_n229_), .Y(new_new_n231_));
  INV        g0209(.A(i_12_), .Y(new_new_n232_));
  NO3        g0210(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n233_));
  NA2        g0211(.A(i_2_), .B(i_1_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n231_), .B(new_new_n227_), .Y(new_new_n235_));
  NAi21      g0213(.An(i_4_), .B(i_3_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n236_), .B(new_new_n73_), .Y(new_new_n237_));
  NO2        g0215(.A(i_0_), .B(i_6_), .Y(new_new_n238_));
  NOi41      g0216(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n234_), .B(new_new_n176_), .Y(new_new_n241_));
  NAi21      g0219(.An(new_new_n240_), .B(new_new_n241_), .Y(new_new_n242_));
  INV        g0220(.A(new_new_n242_), .Y(new_new_n243_));
  AOI220     g0221(.A0(new_new_n243_), .A1(new_new_n39_), .B0(new_new_n235_), .B1(new_new_n200_), .Y(new_new_n244_));
  NO2        g0222(.A(i_11_), .B(new_new_n220_), .Y(new_new_n245_));
  NOi21      g0223(.An(i_1_), .B(i_6_), .Y(new_new_n246_));
  NAi21      g0224(.An(i_3_), .B(i_7_), .Y(new_new_n247_));
  NA2        g0225(.A(new_new_n232_), .B(i_9_), .Y(new_new_n248_));
  OR4        g0226(.A(new_new_n248_), .B(new_new_n247_), .C(new_new_n246_), .D(new_new_n178_), .Y(new_new_n249_));
  NO2        g0227(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n250_));
  NO2        g0228(.A(i_12_), .B(i_3_), .Y(new_new_n251_));
  NA2        g0229(.A(new_new_n71_), .B(i_5_), .Y(new_new_n252_));
  NA2        g0230(.A(i_3_), .B(i_9_), .Y(new_new_n253_));
  NAi21      g0231(.An(i_7_), .B(i_10_), .Y(new_new_n254_));
  NO2        g0232(.A(new_new_n254_), .B(new_new_n253_), .Y(new_new_n255_));
  NA3        g0233(.A(new_new_n255_), .B(new_new_n252_), .C(new_new_n64_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n256_), .B(new_new_n249_), .Y(new_new_n257_));
  NA3        g0235(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n258_));
  NA2        g0236(.A(new_new_n257_), .B(new_new_n245_), .Y(new_new_n259_));
  NO2        g0237(.A(new_new_n228_), .B(new_new_n37_), .Y(new_new_n260_));
  NA2        g0238(.A(i_12_), .B(i_6_), .Y(new_new_n261_));
  OR2        g0239(.A(i_13_), .B(i_9_), .Y(new_new_n262_));
  NO3        g0240(.A(new_new_n262_), .B(new_new_n261_), .C(new_new_n48_), .Y(new_new_n263_));
  NO2        g0241(.A(new_new_n236_), .B(i_2_), .Y(new_new_n264_));
  NA3        g0242(.A(new_new_n264_), .B(new_new_n263_), .C(new_new_n44_), .Y(new_new_n265_));
  NA2        g0243(.A(new_new_n245_), .B(i_9_), .Y(new_new_n266_));
  OAI210     g0244(.A0(new_new_n71_), .A1(new_new_n266_), .B0(new_new_n265_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n150_), .B(new_new_n63_), .Y(new_new_n268_));
  NO3        g0246(.A(i_11_), .B(new_new_n220_), .C(new_new_n25_), .Y(new_new_n269_));
  NO2        g0247(.A(new_new_n247_), .B(i_8_), .Y(new_new_n270_));
  NO2        g0248(.A(i_6_), .B(new_new_n48_), .Y(new_new_n271_));
  NA3        g0249(.A(new_new_n271_), .B(new_new_n270_), .C(new_new_n269_), .Y(new_new_n272_));
  NO3        g0250(.A(new_new_n26_), .B(new_new_n83_), .C(i_5_), .Y(new_new_n273_));
  NA3        g0251(.A(new_new_n273_), .B(new_new_n260_), .C(new_new_n221_), .Y(new_new_n274_));
  AOI210     g0252(.A0(new_new_n274_), .A1(new_new_n272_), .B0(new_new_n268_), .Y(new_new_n275_));
  AOI210     g0253(.A0(new_new_n267_), .A1(new_new_n260_), .B0(new_new_n275_), .Y(new_new_n276_));
  NA4        g0254(.A(new_new_n276_), .B(new_new_n259_), .C(new_new_n244_), .D(new_new_n224_), .Y(new_new_n277_));
  NO3        g0255(.A(i_12_), .B(new_new_n220_), .C(new_new_n37_), .Y(new_new_n278_));
  INV        g0256(.A(new_new_n278_), .Y(new_new_n279_));
  NOi21      g0257(.An(new_new_n159_), .B(new_new_n83_), .Y(new_new_n280_));
  NO3        g0258(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n281_));
  AOI220     g0259(.A0(new_new_n281_), .A1(new_new_n189_), .B0(new_new_n280_), .B1(new_new_n230_), .Y(new_new_n282_));
  NO2        g0260(.A(new_new_n282_), .B(i_7_), .Y(new_new_n283_));
  NO3        g0261(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n284_));
  NO2        g0262(.A(new_new_n234_), .B(i_0_), .Y(new_new_n285_));
  AOI220     g0263(.A0(new_new_n285_), .A1(new_new_n187_), .B0(new_new_n284_), .B1(new_new_n137_), .Y(new_new_n286_));
  NA2        g0264(.A(new_new_n271_), .B(new_new_n26_), .Y(new_new_n287_));
  NO2        g0265(.A(new_new_n287_), .B(new_new_n286_), .Y(new_new_n288_));
  NA2        g0266(.A(i_0_), .B(i_1_), .Y(new_new_n289_));
  NO2        g0267(.A(new_new_n289_), .B(i_2_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n59_), .B(i_6_), .Y(new_new_n291_));
  NA3        g0269(.A(new_new_n291_), .B(new_new_n290_), .C(new_new_n159_), .Y(new_new_n292_));
  OAI210     g0270(.A0(i_2_), .A1(new_new_n138_), .B0(new_new_n292_), .Y(new_new_n293_));
  NO3        g0271(.A(new_new_n293_), .B(new_new_n288_), .C(new_new_n283_), .Y(new_new_n294_));
  NO2        g0272(.A(i_3_), .B(i_10_), .Y(new_new_n295_));
  NA3        g0273(.A(new_new_n295_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n296_));
  NO2        g0274(.A(i_2_), .B(new_new_n99_), .Y(new_new_n297_));
  NOi21      g0275(.An(new_new_n212_), .B(new_new_n100_), .Y(new_new_n298_));
  NA3        g0276(.A(new_new_n298_), .B(i_1_), .C(new_new_n297_), .Y(new_new_n299_));
  AN2        g0277(.A(i_3_), .B(i_10_), .Y(new_new_n300_));
  NA4        g0278(.A(new_new_n300_), .B(new_new_n191_), .C(new_new_n169_), .D(new_new_n167_), .Y(new_new_n301_));
  NO2        g0279(.A(i_5_), .B(new_new_n37_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n303_));
  OR2        g0281(.A(new_new_n299_), .B(new_new_n296_), .Y(new_new_n304_));
  OAI220     g0282(.A0(new_new_n304_), .A1(i_6_), .B0(new_new_n294_), .B1(new_new_n279_), .Y(new_new_n305_));
  NO4        g0283(.A(new_new_n305_), .B(new_new_n277_), .C(new_new_n208_), .D(new_new_n163_), .Y(new_new_n306_));
  NO3        g0284(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n307_));
  NO2        g0285(.A(new_new_n59_), .B(new_new_n83_), .Y(new_new_n308_));
  NA2        g0286(.A(new_new_n285_), .B(new_new_n308_), .Y(new_new_n309_));
  NO3        g0287(.A(i_6_), .B(new_new_n186_), .C(i_7_), .Y(new_new_n310_));
  AOI210     g0288(.A0(new_new_n1030_), .A1(new_new_n309_), .B0(i_5_), .Y(new_new_n311_));
  NO2        g0289(.A(i_2_), .B(i_3_), .Y(new_new_n312_));
  OR2        g0290(.A(i_0_), .B(i_5_), .Y(new_new_n313_));
  NA2        g0291(.A(new_new_n212_), .B(new_new_n313_), .Y(new_new_n314_));
  NA4        g0292(.A(new_new_n314_), .B(new_new_n229_), .C(new_new_n312_), .D(i_1_), .Y(new_new_n315_));
  NA2        g0293(.A(new_new_n285_), .B(new_new_n280_), .Y(new_new_n316_));
  NO2        g0294(.A(new_new_n153_), .B(new_new_n46_), .Y(new_new_n317_));
  NA2        g0295(.A(new_new_n317_), .B(new_new_n159_), .Y(new_new_n318_));
  NA3        g0296(.A(new_new_n318_), .B(new_new_n316_), .C(new_new_n315_), .Y(new_new_n319_));
  OAI210     g0297(.A0(new_new_n319_), .A1(new_new_n311_), .B0(i_4_), .Y(new_new_n320_));
  NO2        g0298(.A(i_12_), .B(i_10_), .Y(new_new_n321_));
  NOi21      g0299(.An(i_5_), .B(i_0_), .Y(new_new_n322_));
  AOI210     g0300(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n99_), .Y(new_new_n323_));
  NO4        g0301(.A(new_new_n323_), .B(i_4_), .C(new_new_n322_), .D(new_new_n124_), .Y(new_new_n324_));
  NA4        g0302(.A(new_new_n81_), .B(new_new_n36_), .C(new_new_n83_), .D(i_8_), .Y(new_new_n325_));
  NA2        g0303(.A(new_new_n324_), .B(new_new_n321_), .Y(new_new_n326_));
  NO2        g0304(.A(i_6_), .B(i_8_), .Y(new_new_n327_));
  AN2        g0305(.A(i_0_), .B(new_new_n327_), .Y(new_new_n328_));
  NO2        g0306(.A(i_1_), .B(i_7_), .Y(new_new_n329_));
  NA3        g0307(.A(i_0_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n330_));
  NA3        g0308(.A(new_new_n330_), .B(new_new_n326_), .C(new_new_n320_), .Y(new_new_n331_));
  NA2        g0309(.A(new_new_n1026_), .B(i_6_), .Y(new_new_n332_));
  NA3        g0310(.A(new_new_n246_), .B(new_new_n297_), .C(new_new_n186_), .Y(new_new_n333_));
  AOI210     g0311(.A0(new_new_n333_), .A1(new_new_n332_), .B0(new_new_n314_), .Y(new_new_n334_));
  NOi21      g0312(.An(new_new_n149_), .B(new_new_n101_), .Y(new_new_n335_));
  NO2        g0313(.A(new_new_n335_), .B(new_new_n120_), .Y(new_new_n336_));
  OAI210     g0314(.A0(new_new_n336_), .A1(new_new_n334_), .B0(i_3_), .Y(new_new_n337_));
  NO2        g0315(.A(new_new_n289_), .B(new_new_n79_), .Y(new_new_n338_));
  NA2        g0316(.A(new_new_n338_), .B(new_new_n128_), .Y(new_new_n339_));
  NO2        g0317(.A(new_new_n90_), .B(new_new_n186_), .Y(new_new_n340_));
  NA3        g0318(.A(new_new_n298_), .B(new_new_n340_), .C(new_new_n63_), .Y(new_new_n341_));
  AOI210     g0319(.A0(new_new_n341_), .A1(new_new_n339_), .B0(i_3_), .Y(new_new_n342_));
  NO2        g0320(.A(new_new_n186_), .B(i_9_), .Y(new_new_n343_));
  NA2        g0321(.A(new_new_n343_), .B(new_new_n199_), .Y(new_new_n344_));
  NO2        g0322(.A(new_new_n342_), .B(new_new_n288_), .Y(new_new_n345_));
  AOI210     g0323(.A0(new_new_n345_), .A1(new_new_n337_), .B0(new_new_n158_), .Y(new_new_n346_));
  AOI210     g0324(.A0(new_new_n331_), .A1(new_new_n307_), .B0(new_new_n346_), .Y(new_new_n347_));
  NOi32      g0325(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n348_));
  INV        g0326(.A(new_new_n348_), .Y(new_new_n349_));
  NAi21      g0327(.An(i_0_), .B(i_6_), .Y(new_new_n350_));
  INV        g0328(.A(new_new_n350_), .Y(new_new_n351_));
  NA2        g0329(.A(new_new_n351_), .B(new_new_n25_), .Y(new_new_n352_));
  OAI210     g0330(.A0(new_new_n352_), .A1(new_new_n155_), .B0(new_new_n240_), .Y(new_new_n353_));
  NAi41      g0331(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n354_));
  NO2        g0332(.A(new_new_n215_), .B(new_new_n155_), .Y(new_new_n355_));
  AOI210     g0333(.A0(new_new_n354_), .A1(new_new_n155_), .B0(new_new_n153_), .Y(new_new_n356_));
  NOi32      g0334(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n357_));
  NAi21      g0335(.An(i_6_), .B(i_1_), .Y(new_new_n358_));
  NA3        g0336(.A(new_new_n358_), .B(new_new_n357_), .C(new_new_n46_), .Y(new_new_n359_));
  NO2        g0337(.A(new_new_n359_), .B(i_0_), .Y(new_new_n360_));
  OR3        g0338(.A(new_new_n360_), .B(new_new_n356_), .C(new_new_n355_), .Y(new_new_n361_));
  NO2        g0339(.A(i_1_), .B(new_new_n99_), .Y(new_new_n362_));
  NAi21      g0340(.An(i_3_), .B(i_4_), .Y(new_new_n363_));
  NO2        g0341(.A(new_new_n363_), .B(i_9_), .Y(new_new_n364_));
  AN2        g0342(.A(i_6_), .B(i_7_), .Y(new_new_n365_));
  OAI210     g0343(.A0(new_new_n365_), .A1(new_new_n362_), .B0(new_new_n364_), .Y(new_new_n366_));
  NA2        g0344(.A(i_2_), .B(i_7_), .Y(new_new_n367_));
  NO2        g0345(.A(new_new_n363_), .B(i_10_), .Y(new_new_n368_));
  NA3        g0346(.A(new_new_n368_), .B(new_new_n367_), .C(new_new_n238_), .Y(new_new_n369_));
  AOI210     g0347(.A0(new_new_n369_), .A1(new_new_n366_), .B0(new_new_n178_), .Y(new_new_n370_));
  AOI220     g0348(.A0(new_new_n368_), .A1(new_new_n329_), .B0(new_new_n233_), .B1(new_new_n181_), .Y(new_new_n371_));
  NO2        g0349(.A(new_new_n371_), .B(i_5_), .Y(new_new_n372_));
  NO4        g0350(.A(new_new_n372_), .B(new_new_n370_), .C(new_new_n361_), .D(new_new_n353_), .Y(new_new_n373_));
  NO2        g0351(.A(new_new_n373_), .B(new_new_n349_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n375_));
  AN2        g0353(.A(i_12_), .B(i_5_), .Y(new_new_n376_));
  NO2        g0354(.A(i_4_), .B(new_new_n26_), .Y(new_new_n377_));
  NA2        g0355(.A(new_new_n377_), .B(new_new_n376_), .Y(new_new_n378_));
  NO2        g0356(.A(i_11_), .B(i_6_), .Y(new_new_n379_));
  NA3        g0357(.A(new_new_n379_), .B(new_new_n317_), .C(new_new_n220_), .Y(new_new_n380_));
  NO2        g0358(.A(new_new_n380_), .B(new_new_n378_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n236_), .B(i_5_), .Y(new_new_n382_));
  NO2        g0360(.A(i_5_), .B(i_10_), .Y(new_new_n383_));
  AOI220     g0361(.A0(new_new_n383_), .A1(new_new_n264_), .B0(new_new_n382_), .B1(new_new_n191_), .Y(new_new_n384_));
  INV        g0362(.A(new_new_n45_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n385_), .B(new_new_n384_), .Y(new_new_n386_));
  OAI210     g0364(.A0(new_new_n386_), .A1(new_new_n381_), .B0(new_new_n375_), .Y(new_new_n387_));
  NO2        g0365(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n388_));
  NO2        g0366(.A(new_new_n145_), .B(new_new_n83_), .Y(new_new_n389_));
  OAI210     g0367(.A0(new_new_n389_), .A1(new_new_n381_), .B0(new_new_n388_), .Y(new_new_n390_));
  NO3        g0368(.A(new_new_n83_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n391_));
  INV        g0369(.A(i_3_), .Y(new_new_n392_));
  NO2        g0370(.A(i_11_), .B(i_12_), .Y(new_new_n393_));
  NAi21      g0371(.An(i_13_), .B(i_0_), .Y(new_new_n394_));
  NA2        g0372(.A(new_new_n390_), .B(new_new_n387_), .Y(new_new_n395_));
  NA2        g0373(.A(new_new_n44_), .B(new_new_n220_), .Y(new_new_n396_));
  NO3        g0374(.A(i_1_), .B(i_12_), .C(new_new_n83_), .Y(new_new_n397_));
  NO2        g0375(.A(i_0_), .B(i_11_), .Y(new_new_n398_));
  AN2        g0376(.A(i_1_), .B(i_6_), .Y(new_new_n399_));
  NOi21      g0377(.An(i_2_), .B(i_12_), .Y(new_new_n400_));
  NA2        g0378(.A(new_new_n400_), .B(new_new_n399_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n401_), .B(new_new_n1022_), .Y(new_new_n402_));
  NA2        g0380(.A(new_new_n137_), .B(i_9_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(i_4_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n402_), .B(new_new_n404_), .Y(new_new_n405_));
  NAi21      g0383(.An(i_9_), .B(i_4_), .Y(new_new_n406_));
  OR2        g0384(.A(i_13_), .B(i_10_), .Y(new_new_n407_));
  NO3        g0385(.A(new_new_n407_), .B(new_new_n113_), .C(new_new_n406_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n166_), .B(new_new_n119_), .Y(new_new_n409_));
  OR2        g0387(.A(new_new_n210_), .B(new_new_n209_), .Y(new_new_n410_));
  NO2        g0388(.A(new_new_n99_), .B(new_new_n25_), .Y(new_new_n411_));
  NA2        g0389(.A(new_new_n278_), .B(new_new_n411_), .Y(new_new_n412_));
  NA2        g0390(.A(new_new_n271_), .B(new_new_n205_), .Y(new_new_n413_));
  OAI220     g0391(.A0(new_new_n413_), .A1(new_new_n410_), .B0(new_new_n412_), .B1(new_new_n335_), .Y(new_new_n414_));
  INV        g0392(.A(new_new_n414_), .Y(new_new_n415_));
  AOI210     g0393(.A0(new_new_n415_), .A1(new_new_n405_), .B0(new_new_n26_), .Y(new_new_n416_));
  NA2        g0394(.A(new_new_n316_), .B(new_new_n315_), .Y(new_new_n417_));
  AOI220     g0395(.A0(new_new_n291_), .A1(new_new_n281_), .B0(new_new_n285_), .B1(new_new_n308_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n418_), .B(i_5_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n176_), .B(new_new_n83_), .Y(new_new_n420_));
  AOI220     g0398(.A0(new_new_n420_), .A1(new_new_n290_), .B0(new_new_n273_), .B1(new_new_n205_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n421_), .B(i_7_), .Y(new_new_n422_));
  NO3        g0400(.A(new_new_n422_), .B(new_new_n419_), .C(new_new_n417_), .Y(new_new_n423_));
  NA2        g0401(.A(new_new_n189_), .B(new_new_n94_), .Y(new_new_n424_));
  NA3        g0402(.A(new_new_n317_), .B(new_new_n159_), .C(new_new_n83_), .Y(new_new_n425_));
  AOI210     g0403(.A0(new_new_n425_), .A1(new_new_n424_), .B0(i_8_), .Y(new_new_n426_));
  NA3        g0404(.A(new_new_n252_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n291_), .B(new_new_n230_), .Y(new_new_n428_));
  OAI220     g0406(.A0(new_new_n428_), .A1(new_new_n176_), .B0(new_new_n427_), .B1(new_new_n1029_), .Y(new_new_n429_));
  NO2        g0407(.A(i_3_), .B(new_new_n48_), .Y(new_new_n430_));
  NA3        g0408(.A(new_new_n329_), .B(new_new_n328_), .C(new_new_n430_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n310_), .B(new_new_n314_), .Y(new_new_n432_));
  OAI210     g0410(.A0(new_new_n432_), .A1(new_new_n182_), .B0(new_new_n431_), .Y(new_new_n433_));
  NO3        g0411(.A(new_new_n433_), .B(new_new_n429_), .C(new_new_n426_), .Y(new_new_n434_));
  AOI210     g0412(.A0(new_new_n434_), .A1(new_new_n423_), .B0(new_new_n266_), .Y(new_new_n435_));
  NO4        g0413(.A(new_new_n435_), .B(new_new_n416_), .C(new_new_n395_), .D(new_new_n374_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n63_), .B(i_4_), .Y(new_new_n437_));
  NO2        g0415(.A(new_new_n71_), .B(i_13_), .Y(new_new_n438_));
  NA3        g0416(.A(new_new_n438_), .B(new_new_n437_), .C(i_2_), .Y(new_new_n439_));
  NO2        g0417(.A(i_10_), .B(i_9_), .Y(new_new_n440_));
  NAi21      g0418(.An(i_12_), .B(i_8_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n441_), .B(i_3_), .Y(new_new_n442_));
  NA2        g0420(.A(new_new_n442_), .B(new_new_n440_), .Y(new_new_n443_));
  NO2        g0421(.A(new_new_n46_), .B(i_4_), .Y(new_new_n444_));
  NA2        g0422(.A(new_new_n444_), .B(new_new_n101_), .Y(new_new_n445_));
  OAI220     g0423(.A0(new_new_n445_), .A1(new_new_n198_), .B0(new_new_n443_), .B1(new_new_n439_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n303_), .B(i_0_), .Y(new_new_n447_));
  NO3        g0425(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n261_), .B(new_new_n95_), .Y(new_new_n449_));
  NA2        g0427(.A(i_8_), .B(i_9_), .Y(new_new_n450_));
  NA2        g0428(.A(new_new_n278_), .B(new_new_n199_), .Y(new_new_n451_));
  NO2        g0429(.A(new_new_n451_), .B(new_new_n450_), .Y(new_new_n452_));
  NO3        g0430(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n453_));
  NA3        g0431(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n452_), .B(new_new_n446_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n290_), .B(new_new_n104_), .Y(new_new_n456_));
  OR2        g0434(.A(new_new_n456_), .B(new_new_n201_), .Y(new_new_n457_));
  OA220      g0435(.A0(new_new_n344_), .A1(new_new_n158_), .B0(new_new_n457_), .B1(new_new_n227_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n94_), .B(i_13_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n420_), .B(new_new_n375_), .Y(new_new_n460_));
  NO2        g0438(.A(i_2_), .B(i_13_), .Y(new_new_n461_));
  NA3        g0439(.A(new_new_n461_), .B(new_new_n157_), .C(new_new_n97_), .Y(new_new_n462_));
  OAI220     g0440(.A0(new_new_n462_), .A1(new_new_n232_), .B0(new_new_n460_), .B1(new_new_n459_), .Y(new_new_n463_));
  NO3        g0441(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n464_));
  NO2        g0442(.A(i_6_), .B(i_7_), .Y(new_new_n465_));
  NOi21      g0443(.An(i_2_), .B(i_7_), .Y(new_new_n466_));
  NAi31      g0444(.An(i_11_), .B(new_new_n466_), .C(new_new_n1023_), .Y(new_new_n467_));
  NO2        g0445(.A(new_new_n407_), .B(i_6_), .Y(new_new_n468_));
  NA3        g0446(.A(new_new_n468_), .B(new_new_n437_), .C(new_new_n73_), .Y(new_new_n469_));
  NO2        g0447(.A(new_new_n469_), .B(new_new_n467_), .Y(new_new_n470_));
  NO2        g0448(.A(i_3_), .B(new_new_n186_), .Y(new_new_n471_));
  NO2        g0449(.A(i_6_), .B(i_10_), .Y(new_new_n472_));
  NA3        g0450(.A(new_new_n239_), .B(new_new_n165_), .C(new_new_n128_), .Y(new_new_n473_));
  NA2        g0451(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n474_));
  NO2        g0452(.A(new_new_n153_), .B(i_3_), .Y(new_new_n475_));
  NAi31      g0453(.An(new_new_n474_), .B(new_new_n475_), .C(new_new_n221_), .Y(new_new_n476_));
  NA3        g0454(.A(new_new_n388_), .B(new_new_n172_), .C(new_new_n144_), .Y(new_new_n477_));
  NA3        g0455(.A(new_new_n477_), .B(new_new_n476_), .C(new_new_n473_), .Y(new_new_n478_));
  NO3        g0456(.A(new_new_n478_), .B(new_new_n470_), .C(new_new_n463_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n448_), .B(new_new_n376_), .Y(new_new_n480_));
  NA2        g0458(.A(new_new_n453_), .B(new_new_n383_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n481_), .B(new_new_n219_), .Y(new_new_n482_));
  NAi21      g0460(.An(new_new_n210_), .B(new_new_n393_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n329_), .B(new_new_n212_), .Y(new_new_n484_));
  NO2        g0462(.A(i_0_), .B(new_new_n83_), .Y(new_new_n485_));
  NA3        g0463(.A(new_new_n485_), .B(i_3_), .C(new_new_n137_), .Y(new_new_n486_));
  OAI220     g0464(.A0(new_new_n38_), .A1(new_new_n486_), .B0(new_new_n484_), .B1(new_new_n483_), .Y(new_new_n487_));
  NA2        g0465(.A(new_new_n27_), .B(i_10_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n307_), .B(new_new_n233_), .Y(new_new_n489_));
  OAI220     g0467(.A0(new_new_n489_), .A1(new_new_n427_), .B0(new_new_n488_), .B1(new_new_n459_), .Y(new_new_n490_));
  NO3        g0468(.A(new_new_n490_), .B(new_new_n487_), .C(new_new_n482_), .Y(new_new_n491_));
  NA4        g0469(.A(new_new_n491_), .B(new_new_n479_), .C(new_new_n458_), .D(new_new_n455_), .Y(new_new_n492_));
  NA3        g0470(.A(new_new_n300_), .B(new_new_n169_), .C(new_new_n167_), .Y(new_new_n493_));
  OAI210     g0471(.A0(new_new_n296_), .A1(new_new_n174_), .B0(new_new_n493_), .Y(new_new_n494_));
  AN2        g0472(.A(new_new_n281_), .B(new_new_n229_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n495_), .B(new_new_n494_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n118_), .B(new_new_n108_), .Y(new_new_n497_));
  AN2        g0475(.A(new_new_n497_), .B(new_new_n448_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n307_), .B(new_new_n160_), .Y(new_new_n499_));
  OAI210     g0477(.A0(new_new_n499_), .A1(new_new_n227_), .B0(new_new_n301_), .Y(new_new_n500_));
  AOI210     g0478(.A0(new_new_n498_), .A1(new_new_n303_), .B0(new_new_n500_), .Y(new_new_n501_));
  NA4        g0479(.A(new_new_n438_), .B(new_new_n437_), .C(new_new_n196_), .D(i_2_), .Y(new_new_n502_));
  INV        g0480(.A(new_new_n502_), .Y(new_new_n503_));
  NA2        g0481(.A(new_new_n376_), .B(new_new_n220_), .Y(new_new_n504_));
  NA2        g0482(.A(new_new_n348_), .B(new_new_n71_), .Y(new_new_n505_));
  NA2        g0483(.A(new_new_n365_), .B(new_new_n357_), .Y(new_new_n506_));
  AO210      g0484(.A0(new_new_n505_), .A1(new_new_n504_), .B0(new_new_n506_), .Y(new_new_n507_));
  NO2        g0485(.A(new_new_n36_), .B(i_8_), .Y(new_new_n508_));
  INV        g0486(.A(new_new_n408_), .Y(new_new_n509_));
  NA2        g0487(.A(new_new_n509_), .B(new_new_n507_), .Y(new_new_n510_));
  AOI210     g0488(.A0(new_new_n503_), .A1(new_new_n197_), .B0(new_new_n510_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n252_), .B(new_new_n64_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n512_), .B(new_new_n129_), .Y(new_new_n513_));
  AOI210     g0491(.A0(new_new_n187_), .A1(i_9_), .B0(new_new_n260_), .Y(new_new_n514_));
  NO2        g0492(.A(new_new_n514_), .B(new_new_n192_), .Y(new_new_n515_));
  AOI220     g0493(.A0(i_3_), .A1(new_new_n515_), .B0(new_new_n513_), .B1(new_new_n409_), .Y(new_new_n516_));
  NA4        g0494(.A(new_new_n516_), .B(new_new_n511_), .C(new_new_n501_), .D(new_new_n496_), .Y(new_new_n517_));
  NO2        g0495(.A(i_12_), .B(new_new_n186_), .Y(new_new_n518_));
  NA3        g0496(.A(new_new_n472_), .B(new_new_n167_), .C(new_new_n27_), .Y(new_new_n519_));
  NO3        g0497(.A(new_new_n519_), .B(i_13_), .C(new_new_n456_), .Y(new_new_n520_));
  NOi31      g0498(.An(new_new_n310_), .B(new_new_n407_), .C(new_new_n38_), .Y(new_new_n521_));
  OAI210     g0499(.A0(new_new_n521_), .A1(new_new_n520_), .B0(new_new_n377_), .Y(new_new_n522_));
  NO2        g0500(.A(i_8_), .B(i_7_), .Y(new_new_n523_));
  OAI210     g0501(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n524_), .B(new_new_n218_), .Y(new_new_n525_));
  AOI220     g0503(.A0(new_new_n317_), .A1(new_new_n39_), .B0(new_new_n230_), .B1(new_new_n200_), .Y(new_new_n526_));
  OAI220     g0504(.A0(new_new_n526_), .A1(new_new_n176_), .B0(new_new_n525_), .B1(new_new_n236_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n44_), .B(i_10_), .Y(new_new_n528_));
  NO2        g0506(.A(new_new_n528_), .B(i_6_), .Y(new_new_n529_));
  NA3        g0507(.A(new_new_n529_), .B(new_new_n527_), .C(new_new_n523_), .Y(new_new_n530_));
  AOI220     g0508(.A0(new_new_n420_), .A1(new_new_n317_), .B0(new_new_n241_), .B1(new_new_n238_), .Y(new_new_n531_));
  OAI220     g0509(.A0(new_new_n531_), .A1(i_12_), .B0(new_new_n459_), .B1(new_new_n129_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n532_), .B(new_new_n260_), .Y(new_new_n533_));
  NOi31      g0511(.An(new_new_n285_), .B(new_new_n296_), .C(new_new_n174_), .Y(new_new_n534_));
  NA3        g0512(.A(new_new_n300_), .B(new_new_n167_), .C(new_new_n94_), .Y(new_new_n535_));
  NO2        g0513(.A(new_new_n153_), .B(i_5_), .Y(new_new_n536_));
  NA3        g0514(.A(new_new_n536_), .B(new_new_n396_), .C(new_new_n312_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n537_), .B(new_new_n535_), .Y(new_new_n538_));
  OAI210     g0516(.A0(new_new_n538_), .A1(new_new_n534_), .B0(new_new_n453_), .Y(new_new_n539_));
  NA4        g0517(.A(new_new_n539_), .B(new_new_n533_), .C(new_new_n530_), .D(new_new_n522_), .Y(new_new_n540_));
  NA3        g0518(.A(new_new_n212_), .B(new_new_n69_), .C(new_new_n44_), .Y(new_new_n541_));
  NA2        g0519(.A(new_new_n278_), .B(new_new_n81_), .Y(new_new_n542_));
  AOI210     g0520(.A0(new_new_n541_), .A1(new_new_n339_), .B0(new_new_n542_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n291_), .B(new_new_n281_), .Y(new_new_n544_));
  NO2        g0522(.A(new_new_n544_), .B(new_new_n166_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n440_), .B(new_new_n216_), .Y(new_new_n547_));
  NO2        g0525(.A(new_new_n546_), .B(new_new_n547_), .Y(new_new_n548_));
  AOI210     g0526(.A0(new_new_n358_), .A1(new_new_n46_), .B0(new_new_n362_), .Y(new_new_n549_));
  NA2        g0527(.A(i_0_), .B(new_new_n48_), .Y(new_new_n550_));
  NA3        g0528(.A(new_new_n518_), .B(new_new_n269_), .C(new_new_n550_), .Y(new_new_n551_));
  NO2        g0529(.A(new_new_n549_), .B(new_new_n551_), .Y(new_new_n552_));
  NO4        g0530(.A(new_new_n552_), .B(new_new_n548_), .C(new_new_n545_), .D(new_new_n543_), .Y(new_new_n553_));
  NO4        g0531(.A(new_new_n246_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n554_));
  NO3        g0532(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n555_));
  NO2        g0533(.A(new_new_n228_), .B(new_new_n36_), .Y(new_new_n556_));
  AN2        g0534(.A(new_new_n556_), .B(new_new_n555_), .Y(new_new_n557_));
  OA210      g0535(.A0(new_new_n557_), .A1(new_new_n554_), .B0(new_new_n348_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n407_), .B(i_1_), .Y(new_new_n559_));
  NOi31      g0537(.An(new_new_n559_), .B(new_new_n449_), .C(new_new_n71_), .Y(new_new_n560_));
  AN3        g0538(.A(new_new_n560_), .B(new_new_n404_), .C(i_2_), .Y(new_new_n561_));
  NO2        g0539(.A(new_new_n418_), .B(new_new_n170_), .Y(new_new_n562_));
  NO3        g0540(.A(new_new_n562_), .B(new_new_n561_), .C(new_new_n558_), .Y(new_new_n563_));
  NOi21      g0541(.An(i_10_), .B(i_6_), .Y(new_new_n564_));
  NO2        g0542(.A(new_new_n83_), .B(new_new_n25_), .Y(new_new_n565_));
  NA2        g0543(.A(new_new_n278_), .B(new_new_n565_), .Y(new_new_n566_));
  NO2        g0544(.A(new_new_n566_), .B(new_new_n447_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n111_), .B(new_new_n23_), .Y(new_new_n568_));
  NA2        g0546(.A(new_new_n310_), .B(new_new_n160_), .Y(new_new_n569_));
  AOI220     g0547(.A0(new_new_n569_), .A1(new_new_n428_), .B0(new_new_n166_), .B1(new_new_n175_), .Y(new_new_n570_));
  NO2        g0548(.A(new_new_n191_), .B(new_new_n37_), .Y(new_new_n571_));
  NOi31      g0549(.An(new_new_n141_), .B(new_new_n571_), .C(new_new_n325_), .Y(new_new_n572_));
  NO3        g0550(.A(new_new_n572_), .B(new_new_n570_), .C(new_new_n567_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n505_), .B(new_new_n371_), .Y(new_new_n574_));
  INV        g0552(.A(new_new_n312_), .Y(new_new_n575_));
  NO2        g0553(.A(i_12_), .B(new_new_n83_), .Y(new_new_n576_));
  NA3        g0554(.A(new_new_n576_), .B(new_new_n269_), .C(new_new_n550_), .Y(new_new_n577_));
  NA3        g0555(.A(new_new_n379_), .B(new_new_n278_), .C(new_new_n212_), .Y(new_new_n578_));
  AOI210     g0556(.A0(new_new_n578_), .A1(new_new_n577_), .B0(new_new_n575_), .Y(new_new_n579_));
  NA2        g0557(.A(new_new_n167_), .B(i_0_), .Y(new_new_n580_));
  NO2        g0558(.A(new_new_n580_), .B(new_new_n296_), .Y(new_new_n581_));
  OR2        g0559(.A(i_2_), .B(i_5_), .Y(new_new_n582_));
  OR2        g0560(.A(new_new_n582_), .B(new_new_n399_), .Y(new_new_n583_));
  NA2        g0561(.A(new_new_n367_), .B(new_new_n238_), .Y(new_new_n584_));
  AOI210     g0562(.A0(new_new_n584_), .A1(new_new_n583_), .B0(new_new_n483_), .Y(new_new_n585_));
  NO4        g0563(.A(new_new_n585_), .B(new_new_n581_), .C(new_new_n579_), .D(new_new_n574_), .Y(new_new_n586_));
  NA4        g0564(.A(new_new_n586_), .B(new_new_n573_), .C(new_new_n563_), .D(new_new_n553_), .Y(new_new_n587_));
  NO4        g0565(.A(new_new_n587_), .B(new_new_n540_), .C(new_new_n517_), .D(new_new_n492_), .Y(new_new_n588_));
  NA4        g0566(.A(new_new_n588_), .B(new_new_n436_), .C(new_new_n347_), .D(new_new_n306_), .Y(men7));
  NO2        g0567(.A(new_new_n104_), .B(new_new_n87_), .Y(new_new_n590_));
  NA2        g0568(.A(new_new_n377_), .B(new_new_n590_), .Y(new_new_n591_));
  NA2        g0569(.A(new_new_n472_), .B(new_new_n81_), .Y(new_new_n592_));
  NA2        g0570(.A(i_11_), .B(new_new_n186_), .Y(new_new_n593_));
  INV        g0571(.A(new_new_n591_), .Y(new_new_n594_));
  NA3        g0572(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n232_), .B(i_4_), .Y(new_new_n596_));
  NA2        g0574(.A(new_new_n596_), .B(i_8_), .Y(new_new_n597_));
  AOI210     g0575(.A0(new_new_n597_), .A1(new_new_n102_), .B0(new_new_n595_), .Y(new_new_n598_));
  NA2        g0576(.A(i_2_), .B(new_new_n83_), .Y(new_new_n599_));
  OAI210     g0577(.A0(new_new_n85_), .A1(new_new_n196_), .B0(new_new_n197_), .Y(new_new_n600_));
  NO2        g0578(.A(i_7_), .B(new_new_n37_), .Y(new_new_n601_));
  NA2        g0579(.A(i_4_), .B(i_8_), .Y(new_new_n602_));
  AOI210     g0580(.A0(new_new_n602_), .A1(new_new_n300_), .B0(new_new_n601_), .Y(new_new_n603_));
  OAI220     g0581(.A0(new_new_n603_), .A1(new_new_n599_), .B0(new_new_n600_), .B1(i_13_), .Y(new_new_n604_));
  NO3        g0582(.A(new_new_n604_), .B(new_new_n598_), .C(new_new_n594_), .Y(new_new_n605_));
  AOI210     g0583(.A0(new_new_n124_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n606_));
  AOI210     g0584(.A0(new_new_n606_), .A1(new_new_n232_), .B0(new_new_n157_), .Y(new_new_n607_));
  OR2        g0585(.A(i_6_), .B(i_10_), .Y(new_new_n608_));
  NO2        g0586(.A(new_new_n608_), .B(new_new_n23_), .Y(new_new_n609_));
  OR3        g0587(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n610_));
  NO3        g0588(.A(new_new_n610_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n611_));
  INV        g0589(.A(new_new_n193_), .Y(new_new_n612_));
  OA220      g0590(.A0(new_new_n610_), .A1(new_new_n575_), .B0(new_new_n607_), .B1(new_new_n262_), .Y(new_new_n613_));
  AOI210     g0591(.A0(new_new_n613_), .A1(new_new_n605_), .B0(new_new_n63_), .Y(new_new_n614_));
  NOi21      g0592(.An(i_11_), .B(i_7_), .Y(new_new_n615_));
  AO210      g0593(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n616_));
  NO2        g0594(.A(new_new_n616_), .B(new_new_n615_), .Y(new_new_n617_));
  NA2        g0595(.A(new_new_n617_), .B(new_new_n200_), .Y(new_new_n618_));
  NA3        g0596(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n619_));
  AOI210     g0597(.A0(new_new_n619_), .A1(new_new_n618_), .B0(new_new_n63_), .Y(new_new_n620_));
  AO210      g0598(.A0(new_new_n84_), .A1(new_new_n371_), .B0(new_new_n40_), .Y(new_new_n621_));
  NO3        g0599(.A(new_new_n254_), .B(new_new_n202_), .C(new_new_n593_), .Y(new_new_n622_));
  OAI210     g0600(.A0(new_new_n622_), .A1(new_new_n221_), .B0(new_new_n63_), .Y(new_new_n623_));
  NA2        g0601(.A(new_new_n400_), .B(new_new_n31_), .Y(new_new_n624_));
  OR2        g0602(.A(new_new_n202_), .B(new_new_n104_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n625_), .B(new_new_n624_), .Y(new_new_n626_));
  NO2        g0604(.A(new_new_n63_), .B(i_9_), .Y(new_new_n627_));
  NO2        g0605(.A(new_new_n627_), .B(i_4_), .Y(new_new_n628_));
  NA2        g0606(.A(new_new_n628_), .B(new_new_n626_), .Y(new_new_n629_));
  NO2        g0607(.A(i_1_), .B(i_12_), .Y(new_new_n630_));
  NA3        g0608(.A(new_new_n630_), .B(new_new_n106_), .C(new_new_n24_), .Y(new_new_n631_));
  NA4        g0609(.A(new_new_n631_), .B(new_new_n629_), .C(new_new_n623_), .D(new_new_n621_), .Y(new_new_n632_));
  OAI210     g0610(.A0(new_new_n632_), .A1(new_new_n620_), .B0(i_6_), .Y(new_new_n633_));
  INV        g0611(.A(new_new_n619_), .Y(new_new_n634_));
  NA2        g0612(.A(new_new_n634_), .B(new_new_n576_), .Y(new_new_n635_));
  NO2        g0613(.A(new_new_n232_), .B(new_new_n83_), .Y(new_new_n636_));
  NO2        g0614(.A(new_new_n636_), .B(i_11_), .Y(new_new_n637_));
  INV        g0615(.A(new_new_n635_), .Y(new_new_n638_));
  NO4        g0616(.A(new_new_n209_), .B(new_new_n124_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n639_));
  NA2        g0617(.A(new_new_n639_), .B(new_new_n627_), .Y(new_new_n640_));
  NO3        g0618(.A(new_new_n608_), .B(new_new_n228_), .C(new_new_n23_), .Y(new_new_n641_));
  AOI210     g0619(.A0(i_1_), .A1(new_new_n255_), .B0(new_new_n641_), .Y(new_new_n642_));
  OAI210     g0620(.A0(new_new_n642_), .A1(new_new_n44_), .B0(new_new_n640_), .Y(new_new_n643_));
  NA3        g0621(.A(new_new_n523_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n644_));
  NA3        g0622(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n645_));
  NO2        g0623(.A(new_new_n46_), .B(i_1_), .Y(new_new_n646_));
  NA3        g0624(.A(new_new_n646_), .B(new_new_n261_), .C(new_new_n44_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n647_), .B(new_new_n645_), .Y(new_new_n648_));
  NA3        g0626(.A(new_new_n627_), .B(new_new_n312_), .C(i_6_), .Y(new_new_n649_));
  NAi21      g0627(.An(new_new_n644_), .B(new_new_n89_), .Y(new_new_n650_));
  NO2        g0628(.A(i_11_), .B(new_new_n37_), .Y(new_new_n651_));
  NA2        g0629(.A(new_new_n651_), .B(new_new_n24_), .Y(new_new_n652_));
  OAI210     g0630(.A0(new_new_n652_), .A1(i_6_), .B0(new_new_n650_), .Y(new_new_n653_));
  OR2        g0631(.A(new_new_n653_), .B(new_new_n648_), .Y(new_new_n654_));
  NO3        g0632(.A(new_new_n654_), .B(new_new_n643_), .C(new_new_n638_), .Y(new_new_n655_));
  NO2        g0633(.A(new_new_n406_), .B(new_new_n83_), .Y(new_new_n656_));
  NA2        g0634(.A(i_3_), .B(new_new_n186_), .Y(new_new_n657_));
  NO2        g0635(.A(new_new_n228_), .B(new_new_n44_), .Y(new_new_n658_));
  NO3        g0636(.A(new_new_n658_), .B(new_new_n303_), .C(i_12_), .Y(new_new_n659_));
  NO2        g0637(.A(new_new_n113_), .B(new_new_n37_), .Y(new_new_n660_));
  NO2        g0638(.A(new_new_n660_), .B(i_6_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n83_), .B(i_9_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n662_), .B(new_new_n63_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n663_), .B(new_new_n630_), .Y(new_new_n664_));
  NO4        g0642(.A(new_new_n664_), .B(new_new_n661_), .C(new_new_n659_), .D(i_4_), .Y(new_new_n665_));
  NA2        g0643(.A(i_1_), .B(i_3_), .Y(new_new_n666_));
  NA2        g0644(.A(new_new_n658_), .B(new_new_n564_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n667_), .B(new_new_n666_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n668_), .B(new_new_n665_), .Y(new_new_n669_));
  NA3        g0647(.A(new_new_n669_), .B(new_new_n655_), .C(new_new_n633_), .Y(new_new_n670_));
  NO3        g0648(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n671_));
  OA210      g0649(.A0(new_new_n671_), .A1(new_new_n239_), .B0(new_new_n83_), .Y(new_new_n672_));
  NA2        g0650(.A(new_new_n365_), .B(new_new_n364_), .Y(new_new_n673_));
  NA3        g0651(.A(new_new_n472_), .B(new_new_n508_), .C(new_new_n46_), .Y(new_new_n674_));
  NO3        g0652(.A(new_new_n466_), .B(new_new_n602_), .C(new_new_n83_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n675_), .B(new_new_n25_), .Y(new_new_n676_));
  NA3        g0654(.A(new_new_n676_), .B(new_new_n674_), .C(new_new_n673_), .Y(new_new_n677_));
  OAI210     g0655(.A0(new_new_n677_), .A1(new_new_n672_), .B0(i_1_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n363_), .B(i_2_), .Y(new_new_n679_));
  AOI210     g0657(.A0(new_new_n649_), .A1(new_new_n678_), .B0(i_13_), .Y(new_new_n680_));
  OR2        g0658(.A(i_11_), .B(i_7_), .Y(new_new_n681_));
  NA2        g0659(.A(new_new_n103_), .B(new_new_n133_), .Y(new_new_n682_));
  AOI220     g0660(.A0(new_new_n461_), .A1(new_new_n157_), .B0(new_new_n444_), .B1(new_new_n133_), .Y(new_new_n683_));
  OAI210     g0661(.A0(new_new_n683_), .A1(new_new_n44_), .B0(new_new_n682_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n466_), .B(new_new_n24_), .Y(new_new_n685_));
  AOI210     g0663(.A0(new_new_n685_), .A1(new_new_n656_), .B0(new_new_n239_), .Y(new_new_n686_));
  OAI220     g0664(.A0(new_new_n686_), .A1(new_new_n40_), .B0(new_new_n54_), .B1(new_new_n90_), .Y(new_new_n687_));
  AOI210     g0665(.A0(new_new_n684_), .A1(new_new_n327_), .B0(new_new_n687_), .Y(new_new_n688_));
  AOI220     g0666(.A0(i_12_), .A1(new_new_n70_), .B0(new_new_n379_), .B1(new_new_n646_), .Y(new_new_n689_));
  NO2        g0667(.A(new_new_n689_), .B(new_new_n236_), .Y(new_new_n690_));
  AOI210     g0668(.A0(new_new_n441_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n691_));
  NOi31      g0669(.An(new_new_n691_), .B(new_new_n592_), .C(new_new_n44_), .Y(new_new_n692_));
  NA2        g0670(.A(new_new_n123_), .B(i_13_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n645_), .B(new_new_n111_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n693_), .B(new_new_n1028_), .Y(new_new_n695_));
  NO3        g0673(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n99_), .Y(new_new_n696_));
  NA2        g0674(.A(i_3_), .B(i_7_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n232_), .B(new_new_n83_), .Y(new_new_n698_));
  AOI210     g0676(.A0(new_new_n698_), .A1(new_new_n697_), .B0(new_new_n696_), .Y(new_new_n699_));
  AOI210     g0677(.A0(new_new_n379_), .A1(new_new_n646_), .B0(new_new_n89_), .Y(new_new_n700_));
  OAI220     g0678(.A0(new_new_n700_), .A1(new_new_n597_), .B0(new_new_n699_), .B1(new_new_n612_), .Y(new_new_n701_));
  NO4        g0679(.A(new_new_n701_), .B(new_new_n695_), .C(new_new_n692_), .D(new_new_n690_), .Y(new_new_n702_));
  NA3        g0680(.A(new_new_n400_), .B(new_new_n601_), .C(new_new_n95_), .Y(new_new_n703_));
  NA2        g0681(.A(new_new_n637_), .B(i_13_), .Y(new_new_n704_));
  NAi21      g0682(.An(i_11_), .B(i_12_), .Y(new_new_n705_));
  NOi41      g0683(.An(new_new_n107_), .B(new_new_n705_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n706_));
  NO2        g0684(.A(new_new_n576_), .B(new_new_n602_), .Y(new_new_n707_));
  AOI210     g0685(.A0(new_new_n707_), .A1(new_new_n307_), .B0(new_new_n706_), .Y(new_new_n708_));
  NA3        g0686(.A(new_new_n708_), .B(new_new_n704_), .C(new_new_n703_), .Y(new_new_n709_));
  OAI210     g0687(.A0(new_new_n709_), .A1(new_new_n694_), .B0(new_new_n63_), .Y(new_new_n710_));
  NA2        g0688(.A(i_8_), .B(new_new_n25_), .Y(new_new_n711_));
  NO3        g0689(.A(new_new_n711_), .B(new_new_n377_), .C(new_new_n596_), .Y(new_new_n712_));
  OAI210     g0690(.A0(new_new_n712_), .A1(new_new_n364_), .B0(new_new_n362_), .Y(new_new_n713_));
  NO2        g0691(.A(new_new_n124_), .B(i_2_), .Y(new_new_n714_));
  INV        g0692(.A(new_new_n714_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n715_), .B(new_new_n713_), .Y(new_new_n716_));
  NA3        g0694(.A(new_new_n716_), .B(new_new_n45_), .C(new_new_n220_), .Y(new_new_n717_));
  NA4        g0695(.A(new_new_n717_), .B(new_new_n710_), .C(new_new_n702_), .D(new_new_n688_), .Y(new_new_n718_));
  OR4        g0696(.A(new_new_n718_), .B(new_new_n680_), .C(new_new_n670_), .D(new_new_n614_), .Y(men5));
  NO2        g0697(.A(new_new_n597_), .B(i_11_), .Y(new_new_n720_));
  NA2        g0698(.A(new_new_n85_), .B(new_new_n720_), .Y(new_new_n721_));
  INV        g0699(.A(new_new_n721_), .Y(new_new_n722_));
  NO3        g0700(.A(i_11_), .B(new_new_n232_), .C(i_13_), .Y(new_new_n723_));
  NO2        g0701(.A(new_new_n120_), .B(new_new_n23_), .Y(new_new_n724_));
  NA2        g0702(.A(i_12_), .B(i_8_), .Y(new_new_n725_));
  OAI210     g0703(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n725_), .Y(new_new_n726_));
  INV        g0704(.A(new_new_n440_), .Y(new_new_n727_));
  AOI220     g0705(.A0(new_new_n312_), .A1(new_new_n568_), .B0(new_new_n726_), .B1(new_new_n724_), .Y(new_new_n728_));
  INV        g0706(.A(new_new_n728_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n729_), .B(new_new_n722_), .Y(new_new_n730_));
  INV        g0708(.A(new_new_n165_), .Y(new_new_n731_));
  INV        g0709(.A(new_new_n239_), .Y(new_new_n732_));
  OAI210     g0710(.A0(new_new_n679_), .A1(new_new_n442_), .B0(new_new_n107_), .Y(new_new_n733_));
  AOI210     g0711(.A0(new_new_n733_), .A1(new_new_n732_), .B0(new_new_n731_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n450_), .B(new_new_n26_), .Y(new_new_n735_));
  NO2        g0713(.A(new_new_n735_), .B(new_new_n411_), .Y(new_new_n736_));
  NA2        g0714(.A(new_new_n736_), .B(i_2_), .Y(new_new_n737_));
  INV        g0715(.A(new_new_n737_), .Y(new_new_n738_));
  AOI210     g0716(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n407_), .Y(new_new_n739_));
  AOI210     g0717(.A0(new_new_n739_), .A1(new_new_n738_), .B0(new_new_n734_), .Y(new_new_n740_));
  NO2        g0718(.A(new_new_n183_), .B(new_new_n121_), .Y(new_new_n741_));
  OAI210     g0719(.A0(new_new_n741_), .A1(new_new_n724_), .B0(i_2_), .Y(new_new_n742_));
  NO2        g0720(.A(new_new_n742_), .B(new_new_n186_), .Y(new_new_n743_));
  OA210      g0721(.A0(new_new_n617_), .A1(new_new_n122_), .B0(i_13_), .Y(new_new_n744_));
  NA2        g0722(.A(new_new_n193_), .B(new_new_n196_), .Y(new_new_n745_));
  NO2        g0723(.A(new_new_n745_), .B(new_new_n367_), .Y(new_new_n746_));
  AOI210     g0724(.A0(new_new_n202_), .A1(new_new_n143_), .B0(new_new_n508_), .Y(new_new_n747_));
  NA2        g0725(.A(new_new_n747_), .B(new_new_n411_), .Y(new_new_n748_));
  NO2        g0726(.A(i_2_), .B(new_new_n44_), .Y(new_new_n749_));
  NA3        g0727(.A(new_new_n300_), .B(new_new_n120_), .C(new_new_n42_), .Y(new_new_n750_));
  OAI210     g0728(.A0(new_new_n750_), .A1(new_new_n749_), .B0(new_new_n748_), .Y(new_new_n751_));
  NO4        g0729(.A(new_new_n751_), .B(new_new_n746_), .C(new_new_n744_), .D(new_new_n743_), .Y(new_new_n752_));
  NA2        g0730(.A(new_new_n568_), .B(new_new_n28_), .Y(new_new_n753_));
  NA2        g0731(.A(new_new_n723_), .B(new_new_n270_), .Y(new_new_n754_));
  NA2        g0732(.A(new_new_n754_), .B(new_new_n753_), .Y(new_new_n755_));
  NO2        g0733(.A(new_new_n62_), .B(i_12_), .Y(new_new_n756_));
  NO2        g0734(.A(new_new_n756_), .B(new_new_n122_), .Y(new_new_n757_));
  NO2        g0735(.A(new_new_n757_), .B(new_new_n593_), .Y(new_new_n758_));
  AOI220     g0736(.A0(new_new_n758_), .A1(new_new_n36_), .B0(new_new_n755_), .B1(new_new_n46_), .Y(new_new_n759_));
  NA4        g0737(.A(new_new_n759_), .B(new_new_n752_), .C(new_new_n740_), .D(new_new_n730_), .Y(men6));
  NA2        g0738(.A(new_new_n25_), .B(new_new_n714_), .Y(new_new_n761_));
  NA4        g0739(.A(new_new_n383_), .B(new_new_n471_), .C(new_new_n69_), .D(new_new_n99_), .Y(new_new_n762_));
  INV        g0740(.A(new_new_n762_), .Y(new_new_n763_));
  NO2        g0741(.A(new_new_n215_), .B(new_new_n474_), .Y(new_new_n764_));
  NO2        g0742(.A(i_11_), .B(i_9_), .Y(new_new_n765_));
  NO2        g0743(.A(new_new_n763_), .B(new_new_n322_), .Y(new_new_n766_));
  AO210      g0744(.A0(new_new_n766_), .A1(new_new_n761_), .B0(i_12_), .Y(new_new_n767_));
  NA2        g0745(.A(new_new_n368_), .B(new_new_n329_), .Y(new_new_n768_));
  NA2        g0746(.A(new_new_n576_), .B(new_new_n63_), .Y(new_new_n769_));
  NA2        g0747(.A(new_new_n671_), .B(new_new_n69_), .Y(new_new_n770_));
  NA4        g0748(.A(new_new_n84_), .B(new_new_n770_), .C(new_new_n769_), .D(new_new_n768_), .Y(new_new_n771_));
  AOI220     g0749(.A0(new_new_n189_), .A1(new_new_n765_), .B0(new_new_n771_), .B1(new_new_n71_), .Y(new_new_n772_));
  NA2        g0750(.A(new_new_n1025_), .B(new_new_n756_), .Y(new_new_n773_));
  AOI210     g0751(.A0(new_new_n773_), .A1(new_new_n506_), .B0(new_new_n178_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n32_), .B(i_11_), .Y(new_new_n775_));
  NA3        g0753(.A(new_new_n775_), .B(new_new_n465_), .C(new_new_n383_), .Y(new_new_n776_));
  NAi32      g0754(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n777_));
  AOI210     g0755(.A0(i_6_), .A1(new_new_n84_), .B0(new_new_n777_), .Y(new_new_n778_));
  OAI210     g0756(.A0(new_new_n671_), .A1(new_new_n556_), .B0(new_new_n555_), .Y(new_new_n779_));
  NAi31      g0757(.An(new_new_n778_), .B(new_new_n779_), .C(new_new_n776_), .Y(new_new_n780_));
  OR2        g0758(.A(new_new_n780_), .B(new_new_n774_), .Y(new_new_n781_));
  NA3        g0759(.A(new_new_n343_), .B(new_new_n251_), .C(i_7_), .Y(new_new_n782_));
  NA3        g0760(.A(new_new_n442_), .B(new_new_n142_), .C(new_new_n67_), .Y(new_new_n783_));
  AO210      g0761(.A0(new_new_n481_), .A1(new_new_n727_), .B0(new_new_n36_), .Y(new_new_n784_));
  NA3        g0762(.A(new_new_n784_), .B(new_new_n783_), .C(new_new_n782_), .Y(new_new_n785_));
  AOI210     g0763(.A0(new_new_n1027_), .A1(new_new_n555_), .B0(new_new_n764_), .Y(new_new_n786_));
  NA3        g0764(.A(new_new_n367_), .B(new_new_n233_), .C(new_new_n142_), .Y(new_new_n787_));
  NA2        g0765(.A(new_new_n391_), .B(new_new_n68_), .Y(new_new_n788_));
  NA3        g0766(.A(new_new_n788_), .B(new_new_n787_), .C(new_new_n786_), .Y(new_new_n789_));
  NA3        g0767(.A(new_new_n46_), .B(new_new_n472_), .C(new_new_n212_), .Y(new_new_n790_));
  AOI210     g0768(.A0(new_new_n442_), .A1(new_new_n440_), .B0(new_new_n554_), .Y(new_new_n791_));
  NA2        g0769(.A(new_new_n108_), .B(new_new_n398_), .Y(new_new_n792_));
  NA3        g0770(.A(new_new_n792_), .B(new_new_n791_), .C(new_new_n790_), .Y(new_new_n793_));
  NO4        g0771(.A(new_new_n793_), .B(new_new_n789_), .C(new_new_n785_), .D(new_new_n781_), .Y(new_new_n794_));
  NA4        g0772(.A(new_new_n794_), .B(new_new_n772_), .C(new_new_n767_), .D(new_new_n373_), .Y(men3));
  NA2        g0773(.A(i_12_), .B(i_10_), .Y(new_new_n796_));
  NA2        g0774(.A(i_6_), .B(i_7_), .Y(new_new_n797_));
  NO2        g0775(.A(new_new_n797_), .B(i_0_), .Y(new_new_n798_));
  NO2        g0776(.A(i_11_), .B(new_new_n232_), .Y(new_new_n799_));
  OAI210     g0777(.A0(new_new_n798_), .A1(new_new_n285_), .B0(new_new_n799_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n800_), .B(new_new_n186_), .Y(new_new_n801_));
  NO3        g0779(.A(new_new_n447_), .B(new_new_n87_), .C(new_new_n44_), .Y(new_new_n802_));
  OA210      g0780(.A0(new_new_n802_), .A1(new_new_n801_), .B0(new_new_n167_), .Y(new_new_n803_));
  NA3        g0781(.A(new_new_n787_), .B(new_new_n600_), .C(new_new_n366_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n804_), .B(new_new_n39_), .Y(new_new_n805_));
  NOi21      g0783(.An(new_new_n94_), .B(new_new_n736_), .Y(new_new_n806_));
  NO3        g0784(.A(new_new_n625_), .B(new_new_n450_), .C(new_new_n127_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n400_), .B(new_new_n45_), .Y(new_new_n808_));
  AN2        g0786(.A(new_new_n449_), .B(new_new_n55_), .Y(new_new_n809_));
  NO3        g0787(.A(new_new_n809_), .B(new_new_n807_), .C(new_new_n806_), .Y(new_new_n810_));
  AOI210     g0788(.A0(new_new_n810_), .A1(new_new_n805_), .B0(new_new_n48_), .Y(new_new_n811_));
  NA2        g0789(.A(new_new_n178_), .B(new_new_n564_), .Y(new_new_n812_));
  NA2        g0790(.A(new_new_n691_), .B(new_new_n662_), .Y(new_new_n813_));
  NA2        g0791(.A(i_0_), .B(new_new_n430_), .Y(new_new_n814_));
  OAI220     g0792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n812_), .B1(new_new_n63_), .Y(new_new_n815_));
  NOi21      g0793(.An(i_5_), .B(i_9_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n816_), .B(new_new_n438_), .Y(new_new_n817_));
  NO3        g0795(.A(new_new_n403_), .B(new_new_n261_), .C(new_new_n71_), .Y(new_new_n818_));
  NO2        g0796(.A(new_new_n168_), .B(new_new_n143_), .Y(new_new_n819_));
  AOI210     g0797(.A0(new_new_n819_), .A1(new_new_n238_), .B0(new_new_n818_), .Y(new_new_n820_));
  OAI220     g0798(.A0(new_new_n820_), .A1(new_new_n174_), .B0(new_new_n602_), .B1(new_new_n817_), .Y(new_new_n821_));
  NO4        g0799(.A(new_new_n821_), .B(new_new_n815_), .C(new_new_n811_), .D(new_new_n803_), .Y(new_new_n822_));
  NA2        g0800(.A(new_new_n178_), .B(new_new_n24_), .Y(new_new_n823_));
  NO2        g0801(.A(new_new_n660_), .B(new_new_n590_), .Y(new_new_n824_));
  NO2        g0802(.A(new_new_n824_), .B(new_new_n823_), .Y(new_new_n825_));
  NA2        g0803(.A(new_new_n307_), .B(new_new_n125_), .Y(new_new_n826_));
  NAi21      g0804(.An(new_new_n158_), .B(new_new_n430_), .Y(new_new_n827_));
  OAI220     g0805(.A0(new_new_n827_), .A1(i_2_), .B0(new_new_n826_), .B1(i_10_), .Y(new_new_n828_));
  NO2        g0806(.A(new_new_n828_), .B(new_new_n825_), .Y(new_new_n829_));
  NO2        g0807(.A(new_new_n383_), .B(new_new_n289_), .Y(new_new_n830_));
  NA2        g0808(.A(new_new_n830_), .B(new_new_n694_), .Y(new_new_n831_));
  NA2        g0809(.A(new_new_n565_), .B(i_0_), .Y(new_new_n832_));
  NO3        g0810(.A(new_new_n832_), .B(new_new_n378_), .C(new_new_n85_), .Y(new_new_n833_));
  NO4        g0811(.A(new_new_n582_), .B(new_new_n209_), .C(new_new_n407_), .D(new_new_n399_), .Y(new_new_n834_));
  AOI210     g0812(.A0(new_new_n834_), .A1(i_11_), .B0(new_new_n833_), .Y(new_new_n835_));
  AN2        g0813(.A(new_new_n94_), .B(new_new_n237_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n723_), .B(new_new_n322_), .Y(new_new_n837_));
  AOI210     g0815(.A0(new_new_n472_), .A1(new_new_n85_), .B0(new_new_n58_), .Y(new_new_n838_));
  OAI220     g0816(.A0(new_new_n838_), .A1(new_new_n837_), .B0(new_new_n652_), .B1(new_new_n525_), .Y(new_new_n839_));
  NO2        g0817(.A(new_new_n248_), .B(new_new_n149_), .Y(new_new_n840_));
  NA2        g0818(.A(i_0_), .B(i_10_), .Y(new_new_n841_));
  OAI210     g0819(.A0(new_new_n841_), .A1(new_new_n83_), .B0(new_new_n528_), .Y(new_new_n842_));
  NO4        g0820(.A(new_new_n111_), .B(new_new_n58_), .C(new_new_n657_), .D(i_5_), .Y(new_new_n843_));
  AO220      g0821(.A0(new_new_n843_), .A1(new_new_n842_), .B0(new_new_n840_), .B1(i_6_), .Y(new_new_n844_));
  AOI220     g0822(.A0(i_0_), .A1(new_new_n96_), .B0(new_new_n178_), .B1(new_new_n81_), .Y(new_new_n845_));
  NA2        g0823(.A(new_new_n559_), .B(i_4_), .Y(new_new_n846_));
  OAI220     g0824(.A0(i_1_), .A1(new_new_n837_), .B0(new_new_n846_), .B1(new_new_n845_), .Y(new_new_n847_));
  NO4        g0825(.A(new_new_n847_), .B(new_new_n844_), .C(new_new_n839_), .D(new_new_n836_), .Y(new_new_n848_));
  NA4        g0826(.A(new_new_n848_), .B(new_new_n835_), .C(new_new_n831_), .D(new_new_n829_), .Y(new_new_n849_));
  NO2        g0827(.A(new_new_n100_), .B(new_new_n37_), .Y(new_new_n850_));
  NA2        g0828(.A(i_11_), .B(i_9_), .Y(new_new_n851_));
  NO3        g0829(.A(i_12_), .B(new_new_n851_), .C(new_new_n599_), .Y(new_new_n852_));
  AN2        g0830(.A(new_new_n852_), .B(new_new_n850_), .Y(new_new_n853_));
  NO2        g0831(.A(new_new_n48_), .B(i_7_), .Y(new_new_n854_));
  INV        g0832(.A(new_new_n156_), .Y(new_new_n855_));
  NO2        g0833(.A(new_new_n851_), .B(new_new_n71_), .Y(new_new_n856_));
  NO2        g0834(.A(new_new_n168_), .B(i_0_), .Y(new_new_n857_));
  INV        g0835(.A(new_new_n857_), .Y(new_new_n858_));
  NA2        g0836(.A(new_new_n465_), .B(new_new_n226_), .Y(new_new_n859_));
  INV        g0837(.A(new_new_n397_), .Y(new_new_n860_));
  OAI220     g0838(.A0(new_new_n860_), .A1(new_new_n817_), .B0(new_new_n859_), .B1(new_new_n858_), .Y(new_new_n861_));
  NO3        g0839(.A(new_new_n861_), .B(new_new_n855_), .C(new_new_n853_), .Y(new_new_n862_));
  NA2        g0840(.A(new_new_n651_), .B(new_new_n117_), .Y(new_new_n863_));
  NO2        g0841(.A(i_6_), .B(new_new_n863_), .Y(new_new_n864_));
  AOI210     g0842(.A0(new_new_n441_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n165_), .B(new_new_n100_), .Y(new_new_n866_));
  NOi32      g0844(.An(new_new_n865_), .Bn(new_new_n181_), .C(new_new_n866_), .Y(new_new_n867_));
  AOI210     g0845(.A0(new_new_n601_), .A1(new_new_n322_), .B0(new_new_n237_), .Y(new_new_n868_));
  NO2        g0846(.A(new_new_n868_), .B(new_new_n808_), .Y(new_new_n869_));
  NO3        g0847(.A(new_new_n869_), .B(new_new_n867_), .C(new_new_n864_), .Y(new_new_n870_));
  NOi21      g0848(.An(i_7_), .B(i_5_), .Y(new_new_n871_));
  NOi31      g0849(.An(new_new_n871_), .B(i_0_), .C(new_new_n705_), .Y(new_new_n872_));
  NA3        g0850(.A(new_new_n872_), .B(new_new_n377_), .C(i_6_), .Y(new_new_n873_));
  OA210      g0851(.A0(new_new_n866_), .A1(new_new_n506_), .B0(new_new_n873_), .Y(new_new_n874_));
  NO2        g0852(.A(new_new_n258_), .B(new_new_n313_), .Y(new_new_n875_));
  NO2        g0853(.A(new_new_n705_), .B(new_new_n253_), .Y(new_new_n876_));
  NA2        g0854(.A(new_new_n876_), .B(new_new_n875_), .Y(new_new_n877_));
  NA4        g0855(.A(new_new_n877_), .B(new_new_n874_), .C(new_new_n870_), .D(new_new_n862_), .Y(new_new_n878_));
  NO2        g0856(.A(new_new_n823_), .B(new_new_n234_), .Y(new_new_n879_));
  AN2        g0857(.A(new_new_n327_), .B(new_new_n322_), .Y(new_new_n880_));
  NA2        g0858(.A(new_new_n879_), .B(i_10_), .Y(new_new_n881_));
  NO2        g0859(.A(new_new_n796_), .B(new_new_n312_), .Y(new_new_n882_));
  OA210      g0860(.A0(new_new_n465_), .A1(new_new_n218_), .B0(new_new_n464_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n882_), .B(new_new_n856_), .Y(new_new_n884_));
  NA3        g0862(.A(new_new_n464_), .B(new_new_n400_), .C(new_new_n45_), .Y(new_new_n885_));
  OAI210     g0863(.A0(new_new_n827_), .A1(i_7_), .B0(new_new_n885_), .Y(new_new_n886_));
  NO2        g0864(.A(new_new_n251_), .B(new_new_n46_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n856_), .B(new_new_n300_), .Y(new_new_n888_));
  OAI210     g0866(.A0(new_new_n887_), .A1(new_new_n180_), .B0(new_new_n888_), .Y(new_new_n889_));
  AOI220     g0867(.A0(new_new_n889_), .A1(new_new_n465_), .B0(new_new_n886_), .B1(new_new_n71_), .Y(new_new_n890_));
  NA3        g0868(.A(i_5_), .B(new_new_n375_), .C(new_new_n636_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n90_), .B(new_new_n44_), .Y(new_new_n892_));
  NO2        g0870(.A(new_new_n73_), .B(new_new_n725_), .Y(new_new_n893_));
  AOI220     g0871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n167_), .B1(new_new_n590_), .Y(new_new_n894_));
  AOI210     g0872(.A0(new_new_n894_), .A1(new_new_n891_), .B0(new_new_n47_), .Y(new_new_n895_));
  NO3        g0873(.A(new_new_n582_), .B(new_new_n350_), .C(new_new_n24_), .Y(new_new_n896_));
  AOI210     g0874(.A0(new_new_n685_), .A1(new_new_n536_), .B0(new_new_n896_), .Y(new_new_n897_));
  NAi21      g0875(.An(i_9_), .B(i_5_), .Y(new_new_n898_));
  NO2        g0876(.A(new_new_n898_), .B(new_new_n394_), .Y(new_new_n899_));
  NO2        g0877(.A(new_new_n595_), .B(new_new_n102_), .Y(new_new_n900_));
  AOI220     g0878(.A0(new_new_n900_), .A1(i_0_), .B0(new_new_n899_), .B1(new_new_n617_), .Y(new_new_n901_));
  OAI220     g0879(.A0(new_new_n901_), .A1(new_new_n83_), .B0(new_new_n897_), .B1(new_new_n166_), .Y(new_new_n902_));
  NO3        g0880(.A(new_new_n902_), .B(new_new_n895_), .C(new_new_n510_), .Y(new_new_n903_));
  NA4        g0881(.A(new_new_n903_), .B(new_new_n890_), .C(new_new_n884_), .D(new_new_n881_), .Y(new_new_n904_));
  NO3        g0882(.A(new_new_n904_), .B(new_new_n878_), .C(new_new_n849_), .Y(new_new_n905_));
  NO2        g0883(.A(i_0_), .B(new_new_n705_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n71_), .B(new_new_n44_), .Y(new_new_n907_));
  NO3        g0885(.A(new_new_n102_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n908_));
  AO220      g0886(.A0(new_new_n908_), .A1(new_new_n44_), .B0(new_new_n906_), .B1(new_new_n167_), .Y(new_new_n909_));
  AOI210     g0887(.A0(new_new_n769_), .A1(new_new_n673_), .B0(new_new_n866_), .Y(new_new_n910_));
  AOI210     g0888(.A0(new_new_n909_), .A1(new_new_n340_), .B0(new_new_n910_), .Y(new_new_n911_));
  NA2        g0889(.A(new_new_n714_), .B(new_new_n141_), .Y(new_new_n912_));
  INV        g0890(.A(new_new_n912_), .Y(new_new_n913_));
  NA2        g0891(.A(new_new_n913_), .B(new_new_n662_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n779_), .B(new_new_n394_), .Y(new_new_n915_));
  NA3        g0893(.A(new_new_n798_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n916_));
  NA2        g0894(.A(new_new_n799_), .B(i_9_), .Y(new_new_n917_));
  AOI210     g0895(.A0(new_new_n916_), .A1(new_new_n486_), .B0(new_new_n917_), .Y(new_new_n918_));
  OAI210     g0896(.A0(new_new_n238_), .A1(i_9_), .B0(new_new_n225_), .Y(new_new_n919_));
  AOI210     g0897(.A0(new_new_n919_), .A1(new_new_n832_), .B0(new_new_n149_), .Y(new_new_n920_));
  NO3        g0898(.A(new_new_n920_), .B(new_new_n918_), .C(new_new_n915_), .Y(new_new_n921_));
  NA3        g0899(.A(new_new_n921_), .B(new_new_n914_), .C(new_new_n911_), .Y(new_new_n922_));
  NA2        g0900(.A(new_new_n880_), .B(new_new_n367_), .Y(new_new_n923_));
  AOI210     g0901(.A0(new_new_n296_), .A1(new_new_n158_), .B0(new_new_n923_), .Y(new_new_n924_));
  INV        g0902(.A(new_new_n924_), .Y(new_new_n925_));
  NO3        g0903(.A(new_new_n841_), .B(new_new_n816_), .C(new_new_n183_), .Y(new_new_n926_));
  NA2        g0904(.A(new_new_n926_), .B(i_11_), .Y(new_new_n927_));
  NO3        g0905(.A(new_new_n204_), .B(new_new_n376_), .C(i_0_), .Y(new_new_n928_));
  OAI210     g0906(.A0(new_new_n928_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n929_));
  INV        g0907(.A(new_new_n212_), .Y(new_new_n930_));
  NO2        g0908(.A(i_12_), .B(new_new_n612_), .Y(new_new_n931_));
  NA3        g0909(.A(new_new_n931_), .B(new_new_n392_), .C(new_new_n930_), .Y(new_new_n932_));
  NA4        g0910(.A(new_new_n932_), .B(new_new_n929_), .C(new_new_n927_), .D(new_new_n925_), .Y(new_new_n933_));
  NO2        g0911(.A(new_new_n236_), .B(new_new_n90_), .Y(new_new_n934_));
  AOI210     g0912(.A0(new_new_n934_), .A1(new_new_n906_), .B0(new_new_n105_), .Y(new_new_n935_));
  AOI220     g0913(.A0(new_new_n871_), .A1(new_new_n475_), .B0(new_new_n798_), .B1(new_new_n159_), .Y(new_new_n936_));
  NA2        g0914(.A(new_new_n343_), .B(new_new_n169_), .Y(new_new_n937_));
  OA220      g0915(.A0(new_new_n937_), .A1(new_new_n936_), .B0(new_new_n935_), .B1(i_5_), .Y(new_new_n938_));
  AOI210     g0916(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n168_), .Y(new_new_n939_));
  NA2        g0917(.A(new_new_n939_), .B(new_new_n883_), .Y(new_new_n940_));
  NA3        g0918(.A(new_new_n609_), .B(new_new_n178_), .C(new_new_n81_), .Y(new_new_n941_));
  NA2        g0919(.A(new_new_n941_), .B(new_new_n535_), .Y(new_new_n942_));
  NO3        g0920(.A(new_new_n808_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n943_));
  NA3        g0921(.A(new_new_n480_), .B(new_new_n473_), .C(new_new_n462_), .Y(new_new_n944_));
  NO3        g0922(.A(new_new_n944_), .B(new_new_n943_), .C(new_new_n942_), .Y(new_new_n945_));
  NA3        g0923(.A(new_new_n383_), .B(new_new_n165_), .C(new_new_n164_), .Y(new_new_n946_));
  NA3        g0924(.A(new_new_n383_), .B(new_new_n328_), .C(new_new_n216_), .Y(new_new_n947_));
  INV        g0925(.A(new_new_n947_), .Y(new_new_n948_));
  NOi31      g0926(.An(new_new_n382_), .B(new_new_n907_), .C(new_new_n234_), .Y(new_new_n949_));
  NO3        g0927(.A(new_new_n949_), .B(new_new_n948_), .C(new_new_n1024_), .Y(new_new_n950_));
  NA4        g0928(.A(new_new_n950_), .B(new_new_n945_), .C(new_new_n940_), .D(new_new_n938_), .Y(new_new_n951_));
  INV        g0929(.A(new_new_n611_), .Y(new_new_n952_));
  NO3        g0930(.A(new_new_n952_), .B(new_new_n550_), .C(i_3_), .Y(new_new_n953_));
  NO2        g0931(.A(new_new_n83_), .B(i_5_), .Y(new_new_n954_));
  NA3        g0932(.A(new_new_n799_), .B(new_new_n106_), .C(new_new_n120_), .Y(new_new_n955_));
  INV        g0933(.A(new_new_n955_), .Y(new_new_n956_));
  AOI210     g0934(.A0(new_new_n956_), .A1(new_new_n954_), .B0(new_new_n953_), .Y(new_new_n957_));
  NA3        g0935(.A(new_new_n300_), .B(i_5_), .C(new_new_n186_), .Y(new_new_n958_));
  NO4        g0936(.A(new_new_n234_), .B(new_new_n204_), .C(i_0_), .D(i_12_), .Y(new_new_n959_));
  AOI220     g0937(.A0(new_new_n959_), .A1(i_10_), .B0(new_new_n763_), .B1(new_new_n169_), .Y(new_new_n960_));
  AN2        g0938(.A(new_new_n841_), .B(new_new_n149_), .Y(new_new_n961_));
  NO4        g0939(.A(new_new_n961_), .B(i_12_), .C(new_new_n644_), .D(new_new_n127_), .Y(new_new_n962_));
  NA2        g0940(.A(new_new_n962_), .B(new_new_n212_), .Y(new_new_n963_));
  NA3        g0941(.A(new_new_n96_), .B(new_new_n564_), .C(i_11_), .Y(new_new_n964_));
  NO2        g0942(.A(new_new_n964_), .B(new_new_n151_), .Y(new_new_n965_));
  NA2        g0943(.A(new_new_n871_), .B(new_new_n461_), .Y(new_new_n966_));
  INV        g0944(.A(new_new_n64_), .Y(new_new_n967_));
  OAI220     g0945(.A0(new_new_n967_), .A1(new_new_n958_), .B0(new_new_n966_), .B1(new_new_n663_), .Y(new_new_n968_));
  AOI210     g0946(.A0(new_new_n968_), .A1(new_new_n857_), .B0(new_new_n965_), .Y(new_new_n969_));
  NA4        g0947(.A(new_new_n969_), .B(new_new_n963_), .C(new_new_n960_), .D(new_new_n957_), .Y(new_new_n970_));
  NO4        g0948(.A(new_new_n970_), .B(new_new_n951_), .C(new_new_n933_), .D(new_new_n922_), .Y(new_new_n971_));
  NA2        g0949(.A(new_new_n775_), .B(new_new_n37_), .Y(new_new_n972_));
  NA3        g0950(.A(new_new_n865_), .B(new_new_n362_), .C(i_5_), .Y(new_new_n973_));
  NA3        g0951(.A(new_new_n973_), .B(new_new_n972_), .C(new_new_n607_), .Y(new_new_n974_));
  NA2        g0952(.A(new_new_n974_), .B(new_new_n200_), .Y(new_new_n975_));
  AN2        g0953(.A(new_new_n681_), .B(new_new_n363_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n179_), .B(new_new_n181_), .Y(new_new_n977_));
  AO210      g0955(.A0(new_new_n976_), .A1(new_new_n33_), .B0(new_new_n977_), .Y(new_new_n978_));
  OAI210     g0956(.A0(new_new_n611_), .A1(new_new_n609_), .B0(new_new_n312_), .Y(new_new_n979_));
  NAi31      g0957(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n980_));
  NO2        g0958(.A(new_new_n68_), .B(new_new_n980_), .Y(new_new_n981_));
  NO2        g0959(.A(new_new_n981_), .B(new_new_n641_), .Y(new_new_n982_));
  NA3        g0960(.A(new_new_n982_), .B(new_new_n979_), .C(new_new_n978_), .Y(new_new_n983_));
  NO2        g0961(.A(new_new_n454_), .B(new_new_n261_), .Y(new_new_n984_));
  NO4        g0962(.A(new_new_n228_), .B(new_new_n140_), .C(new_new_n666_), .D(new_new_n37_), .Y(new_new_n985_));
  NO3        g0963(.A(new_new_n985_), .B(new_new_n984_), .C(new_new_n834_), .Y(new_new_n986_));
  OAI210     g0964(.A0(new_new_n964_), .A1(new_new_n143_), .B0(new_new_n986_), .Y(new_new_n987_));
  AOI210     g0965(.A0(new_new_n983_), .A1(new_new_n48_), .B0(new_new_n987_), .Y(new_new_n988_));
  AOI210     g0966(.A0(new_new_n988_), .A1(new_new_n975_), .B0(new_new_n71_), .Y(new_new_n989_));
  NO2        g0967(.A(new_new_n557_), .B(new_new_n372_), .Y(new_new_n990_));
  NO2        g0968(.A(new_new_n990_), .B(new_new_n731_), .Y(new_new_n991_));
  OAI210     g0969(.A0(new_new_n78_), .A1(new_new_n54_), .B0(new_new_n104_), .Y(new_new_n992_));
  NA2        g0970(.A(new_new_n992_), .B(new_new_n74_), .Y(new_new_n993_));
  AOI210     g0971(.A0(new_new_n939_), .A1(new_new_n854_), .B0(new_new_n872_), .Y(new_new_n994_));
  AOI210     g0972(.A0(new_new_n994_), .A1(new_new_n993_), .B0(new_new_n666_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n258_), .B(new_new_n57_), .Y(new_new_n996_));
  AOI220     g0974(.A0(new_new_n996_), .A1(new_new_n74_), .B0(new_new_n338_), .B1(new_new_n250_), .Y(new_new_n997_));
  NO2        g0975(.A(new_new_n997_), .B(new_new_n232_), .Y(new_new_n998_));
  NA3        g0976(.A(new_new_n94_), .B(new_new_n302_), .C(new_new_n31_), .Y(new_new_n999_));
  INV        g0977(.A(new_new_n999_), .Y(new_new_n1000_));
  NO3        g0978(.A(new_new_n1000_), .B(new_new_n998_), .C(new_new_n995_), .Y(new_new_n1001_));
  OAI210     g0979(.A0(new_new_n263_), .A1(new_new_n154_), .B0(new_new_n85_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n735_), .B(new_new_n285_), .C(new_new_n78_), .Y(new_new_n1003_));
  AOI210     g0981(.A0(new_new_n1003_), .A1(new_new_n1002_), .B0(i_11_), .Y(new_new_n1004_));
  NA2        g0982(.A(new_new_n602_), .B(new_new_n209_), .Y(new_new_n1005_));
  OAI210     g0983(.A0(new_new_n1005_), .A1(new_new_n865_), .B0(new_new_n200_), .Y(new_new_n1006_));
  NA2        g0984(.A(new_new_n160_), .B(i_5_), .Y(new_new_n1007_));
  NO2        g0985(.A(new_new_n1006_), .B(new_new_n1007_), .Y(new_new_n1008_));
  NO3        g0986(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1009_));
  OAI210     g0987(.A0(new_new_n875_), .A1(new_new_n302_), .B0(new_new_n1009_), .Y(new_new_n1010_));
  NO2        g0988(.A(new_new_n1010_), .B(new_new_n705_), .Y(new_new_n1011_));
  NO4        g0989(.A(new_new_n898_), .B(i_11_), .C(new_new_n247_), .D(new_new_n246_), .Y(new_new_n1012_));
  NO2        g0990(.A(new_new_n1012_), .B(new_new_n554_), .Y(new_new_n1013_));
  NO2        g0991(.A(new_new_n778_), .B(new_new_n355_), .Y(new_new_n1014_));
  AOI210     g0992(.A0(new_new_n1014_), .A1(new_new_n1013_), .B0(new_new_n40_), .Y(new_new_n1015_));
  NO4        g0993(.A(new_new_n1015_), .B(new_new_n1011_), .C(new_new_n1008_), .D(new_new_n1004_), .Y(new_new_n1016_));
  OAI210     g0994(.A0(new_new_n1001_), .A1(i_4_), .B0(new_new_n1016_), .Y(new_new_n1017_));
  NO3        g0995(.A(new_new_n1017_), .B(new_new_n991_), .C(new_new_n989_), .Y(new_new_n1018_));
  NA4        g0996(.A(new_new_n1018_), .B(new_new_n971_), .C(new_new_n905_), .D(new_new_n822_), .Y(men4));
  INV        g0997(.A(i_5_), .Y(new_new_n1022_));
  INV        g0998(.A(i_3_), .Y(new_new_n1023_));
  INV        g0999(.A(new_new_n946_), .Y(new_new_n1024_));
  INV        g1000(.A(i_9_), .Y(new_new_n1025_));
  INV        g1001(.A(i_1_), .Y(new_new_n1026_));
  INV        g1002(.A(i_11_), .Y(new_new_n1027_));
  INV        g1003(.A(i_1_), .Y(new_new_n1028_));
  INV        g1004(.A(i_10_), .Y(new_new_n1029_));
  INV        g1005(.A(new_new_n191_), .Y(new_new_n1030_));
endmodule


