//Benchmark atmr_alu4_1266_0.5

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n112_, ori_ori_n113_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n125_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  BUFFER     o008(.A(i_11_), .Y(ori_ori_n31_));
  BUFFER     o009(.A(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n35_), .Y(ori1));
  INV        o019(.A(i_11_), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(i_6_), .Y(ori_ori_n43_));
  INV        o021(.A(i_2_), .Y(ori_ori_n44_));
  INV        o022(.A(i_5_), .Y(ori_ori_n45_));
  NO2        o023(.A(i_7_), .B(i_10_), .Y(ori_ori_n46_));
  AOI210     o024(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n46_), .Y(ori_ori_n47_));
  NA2        o025(.A(i_0_), .B(i_2_), .Y(ori_ori_n48_));
  NA2        o026(.A(i_7_), .B(i_9_), .Y(ori_ori_n49_));
  NO2        o027(.A(ori_ori_n49_), .B(ori_ori_n48_), .Y(ori_ori_n50_));
  NA2        o028(.A(i_2_), .B(ori_ori_n43_), .Y(ori_ori_n51_));
  NO2        o029(.A(i_1_), .B(i_6_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_8_), .B(i_7_), .Y(ori_ori_n53_));
  NAi21      o031(.An(i_2_), .B(i_7_), .Y(ori_ori_n54_));
  INV        o032(.A(i_1_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n55_), .B(i_6_), .Y(ori_ori_n56_));
  NA3        o034(.A(ori_ori_n56_), .B(ori_ori_n54_), .C(ori_ori_n31_), .Y(ori_ori_n57_));
  NA2        o035(.A(i_1_), .B(i_10_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(i_6_), .Y(ori_ori_n59_));
  NAi21      o037(.An(ori_ori_n59_), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n47_), .B(i_2_), .Y(ori_ori_n61_));
  AOI210     o039(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n62_));
  NA2        o040(.A(i_1_), .B(i_6_), .Y(ori_ori_n63_));
  NO2        o041(.A(ori_ori_n63_), .B(ori_ori_n25_), .Y(ori_ori_n64_));
  INV        o042(.A(i_0_), .Y(ori_ori_n65_));
  NA2        o043(.A(i_5_), .B(i_9_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  NO2        o045(.A(ori_ori_n67_), .B(ori_ori_n64_), .Y(ori_ori_n68_));
  OAI210     o046(.A0(ori_ori_n62_), .A1(ori_ori_n61_), .B0(ori_ori_n68_), .Y(ori_ori_n69_));
  OAI210     o047(.A0(ori_ori_n69_), .A1(ori_ori_n60_), .B0(i_0_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_12_), .B(i_5_), .Y(ori_ori_n71_));
  NO2        o049(.A(i_3_), .B(i_7_), .Y(ori_ori_n72_));
  INV        o050(.A(i_6_), .Y(ori_ori_n73_));
  NO2        o051(.A(i_2_), .B(i_7_), .Y(ori_ori_n74_));
  INV        o052(.A(ori_ori_n74_), .Y(ori_ori_n75_));
  NA2        o053(.A(i_1_), .B(ori_ori_n75_), .Y(ori_ori_n76_));
  NAi21      o054(.An(i_6_), .B(i_10_), .Y(ori_ori_n77_));
  NA2        o055(.A(i_6_), .B(i_9_), .Y(ori_ori_n78_));
  AOI210     o056(.A0(ori_ori_n78_), .A1(ori_ori_n77_), .B0(ori_ori_n55_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_2_), .B(i_6_), .Y(ori_ori_n80_));
  INV        o058(.A(ori_ori_n79_), .Y(ori_ori_n81_));
  AOI210     o059(.A0(ori_ori_n81_), .A1(ori_ori_n76_), .B0(ori_ori_n71_), .Y(ori_ori_n82_));
  AN3        o060(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n83_));
  NAi21      o061(.An(i_6_), .B(i_11_), .Y(ori_ori_n84_));
  INV        o062(.A(i_7_), .Y(ori_ori_n85_));
  NA2        o063(.A(ori_ori_n44_), .B(ori_ori_n85_), .Y(ori_ori_n86_));
  NO2        o064(.A(i_0_), .B(i_5_), .Y(ori_ori_n87_));
  NO2        o065(.A(ori_ori_n87_), .B(ori_ori_n73_), .Y(ori_ori_n88_));
  NA2        o066(.A(i_12_), .B(i_3_), .Y(ori_ori_n89_));
  NA3        o067(.A(i_12_), .B(ori_ori_n88_), .C(ori_ori_n86_), .Y(ori_ori_n90_));
  NAi21      o068(.An(i_7_), .B(i_11_), .Y(ori_ori_n91_));
  AN2        o069(.A(i_2_), .B(i_10_), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n92_), .B(i_7_), .Y(ori_ori_n93_));
  BUFFER     o071(.A(ori_ori_n71_), .Y(ori_ori_n94_));
  NA2        o072(.A(i_12_), .B(i_7_), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n55_), .B(ori_ori_n26_), .Y(ori_ori_n96_));
  NA2        o074(.A(i_11_), .B(i_12_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n97_), .B(ori_ori_n90_), .Y(ori_ori_n98_));
  BUFFER     o076(.A(i_1_), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n99_), .B(i_11_), .Y(ori_ori_n100_));
  NA2        o078(.A(ori_ori_n85_), .B(ori_ori_n37_), .Y(ori_ori_n101_));
  NA2        o079(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n102_), .B(ori_ori_n101_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n103_), .B(ori_ori_n44_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n78_), .B(ori_ori_n77_), .Y(ori_ori_n105_));
  NAi21      o083(.An(i_3_), .B(i_8_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n105_), .B(ori_ori_n104_), .Y(ori_ori_n107_));
  NO2        o085(.A(i_6_), .B(i_5_), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n107_), .B(ori_ori_n100_), .Y(ori_ori_n109_));
  NO3        o087(.A(ori_ori_n109_), .B(ori_ori_n98_), .C(ori_ori_n82_), .Y(ori_ori_n110_));
  NA3        o088(.A(ori_ori_n110_), .B(ori_ori_n70_), .C(ori_ori_n51_), .Y(ori2));
  NO2        o089(.A(ori_ori_n55_), .B(ori_ori_n37_), .Y(ori_ori_n112_));
  INV        o090(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  NA4        o091(.A(ori_ori_n113_), .B(ori_ori_n68_), .C(ori_ori_n61_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o092(.A(i_12_), .B(i_13_), .Y(ori_ori_n115_));
  NAi21      o093(.An(i_5_), .B(i_11_), .Y(ori_ori_n116_));
  NO2        o094(.A(i_0_), .B(i_1_), .Y(ori_ori_n117_));
  NA2        o095(.A(i_1_), .B(i_5_), .Y(ori_ori_n118_));
  OR2        o096(.A(i_0_), .B(i_1_), .Y(ori_ori_n119_));
  NOi21      o097(.An(i_4_), .B(i_10_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(ori_ori_n40_), .Y(ori_ori_n121_));
  NOi21      o099(.An(i_4_), .B(i_9_), .Y(ori_ori_n122_));
  NOi21      o100(.An(i_11_), .B(i_13_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(ori_ori_n122_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n65_), .B(i_5_), .Y(ori_ori_n125_));
  NO2        o103(.A(i_2_), .B(i_1_), .Y(ori_ori_n126_));
  NAi21      o104(.An(i_4_), .B(i_12_), .Y(ori_ori_n127_));
  INV        o105(.A(i_8_), .Y(ori_ori_n128_));
  NO2        o106(.A(i_3_), .B(i_8_), .Y(ori_ori_n129_));
  NO3        o107(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n130_));
  NO2        o108(.A(ori_ori_n87_), .B(ori_ori_n52_), .Y(ori_ori_n131_));
  NO2        o109(.A(i_13_), .B(i_9_), .Y(ori_ori_n132_));
  NAi21      o110(.An(i_12_), .B(i_3_), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n42_), .B(i_5_), .Y(ori_ori_n134_));
  NA3        o112(.A(i_13_), .B(ori_ori_n128_), .C(i_10_), .Y(ori_ori_n135_));
  NA2        o113(.A(i_0_), .B(i_5_), .Y(ori_ori_n136_));
  NAi31      o114(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n65_), .B(ori_ori_n26_), .Y(ori_ori_n138_));
  NO2        o116(.A(ori_ori_n44_), .B(ori_ori_n55_), .Y(ori_ori_n139_));
  INV        o117(.A(i_13_), .Y(ori_ori_n140_));
  NO2        o118(.A(i_12_), .B(ori_ori_n140_), .Y(ori_ori_n141_));
  OR2        o119(.A(i_8_), .B(i_7_), .Y(ori_ori_n142_));
  INV        o120(.A(i_12_), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n42_), .B(ori_ori_n143_), .Y(ori_ori_n144_));
  NO3        o122(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n145_));
  NA2        o123(.A(i_2_), .B(i_1_), .Y(ori_ori_n146_));
  NAi21      o124(.An(i_4_), .B(i_3_), .Y(ori_ori_n147_));
  NO2        o125(.A(i_0_), .B(i_6_), .Y(ori_ori_n148_));
  NOi41      o126(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n149_));
  NO2        o127(.A(i_11_), .B(ori_ori_n140_), .Y(ori_ori_n150_));
  NOi21      o128(.An(i_1_), .B(i_6_), .Y(ori_ori_n151_));
  NAi21      o129(.An(i_3_), .B(i_7_), .Y(ori_ori_n152_));
  NA2        o130(.A(ori_ori_n143_), .B(i_9_), .Y(ori_ori_n153_));
  OR4        o131(.A(ori_ori_n153_), .B(ori_ori_n152_), .C(ori_ori_n151_), .D(ori_ori_n125_), .Y(ori_ori_n154_));
  NA2        o132(.A(ori_ori_n65_), .B(i_5_), .Y(ori_ori_n155_));
  NA2        o133(.A(i_3_), .B(i_9_), .Y(ori_ori_n156_));
  NAi21      o134(.An(i_7_), .B(i_10_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n157_), .B(ori_ori_n156_), .Y(ori_ori_n158_));
  NA3        o136(.A(ori_ori_n158_), .B(ori_ori_n155_), .C(ori_ori_n56_), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n159_), .B(ori_ori_n154_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(ori_ori_n150_), .Y(ori_ori_n161_));
  NA2        o139(.A(i_12_), .B(i_6_), .Y(ori_ori_n162_));
  OR2        o140(.A(i_13_), .B(i_9_), .Y(ori_ori_n163_));
  NO2        o141(.A(ori_ori_n147_), .B(i_2_), .Y(ori_ori_n164_));
  NA2        o142(.A(ori_ori_n150_), .B(i_9_), .Y(ori_ori_n165_));
  NO3        o143(.A(i_11_), .B(ori_ori_n140_), .C(ori_ori_n25_), .Y(ori_ori_n166_));
  NO3        o144(.A(i_12_), .B(ori_ori_n140_), .C(ori_ori_n37_), .Y(ori_ori_n167_));
  AN2        o145(.A(i_3_), .B(i_10_), .Y(ori_ori_n168_));
  NO2        o146(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n169_));
  NO3        o147(.A(ori_ori_n42_), .B(i_13_), .C(i_9_), .Y(ori_ori_n170_));
  NO2        o148(.A(i_2_), .B(i_3_), .Y(ori_ori_n171_));
  NO2        o149(.A(i_12_), .B(i_10_), .Y(ori_ori_n172_));
  NOi21      o150(.An(i_5_), .B(i_0_), .Y(ori_ori_n173_));
  NO2        o151(.A(i_1_), .B(i_7_), .Y(ori_ori_n174_));
  NOi21      o152(.An(ori_ori_n118_), .B(ori_ori_n88_), .Y(ori_ori_n175_));
  NO2        o153(.A(ori_ori_n175_), .B(ori_ori_n102_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(i_3_), .Y(ori_ori_n177_));
  NO2        o155(.A(ori_ori_n128_), .B(i_9_), .Y(ori_ori_n178_));
  NA2        o156(.A(ori_ori_n178_), .B(ori_ori_n131_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n179_), .B(ori_ori_n44_), .Y(ori_ori_n180_));
  INV        o158(.A(ori_ori_n180_), .Y(ori_ori_n181_));
  AOI210     o159(.A0(ori_ori_n181_), .A1(ori_ori_n177_), .B0(ori_ori_n121_), .Y(ori_ori_n182_));
  INV        o160(.A(ori_ori_n182_), .Y(ori_ori_n183_));
  NOi32      o161(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n184_));
  INV        o162(.A(ori_ori_n184_), .Y(ori_ori_n185_));
  NOi32      o163(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n186_));
  NAi21      o164(.An(i_6_), .B(i_1_), .Y(ori_ori_n187_));
  NA3        o165(.A(ori_ori_n187_), .B(ori_ori_n186_), .C(ori_ori_n44_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n188_), .B(i_0_), .Y(ori_ori_n189_));
  NO2        o167(.A(i_1_), .B(ori_ori_n85_), .Y(ori_ori_n190_));
  NAi21      o168(.An(i_3_), .B(i_4_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n191_), .B(i_9_), .Y(ori_ori_n192_));
  AN2        o170(.A(i_6_), .B(i_7_), .Y(ori_ori_n193_));
  OAI210     o171(.A0(ori_ori_n193_), .A1(ori_ori_n190_), .B0(ori_ori_n192_), .Y(ori_ori_n194_));
  NA2        o172(.A(i_2_), .B(i_7_), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n191_), .B(i_10_), .Y(ori_ori_n196_));
  NA3        o174(.A(ori_ori_n196_), .B(ori_ori_n195_), .C(ori_ori_n148_), .Y(ori_ori_n197_));
  AOI210     o175(.A0(ori_ori_n197_), .A1(ori_ori_n194_), .B0(ori_ori_n125_), .Y(ori_ori_n198_));
  AOI210     o176(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n199_));
  OAI210     o177(.A0(ori_ori_n199_), .A1(ori_ori_n126_), .B0(ori_ori_n196_), .Y(ori_ori_n200_));
  AOI220     o178(.A0(ori_ori_n196_), .A1(ori_ori_n174_), .B0(ori_ori_n145_), .B1(ori_ori_n126_), .Y(ori_ori_n201_));
  AOI210     o179(.A0(ori_ori_n201_), .A1(ori_ori_n200_), .B0(i_5_), .Y(ori_ori_n202_));
  NO3        o180(.A(ori_ori_n202_), .B(ori_ori_n198_), .C(ori_ori_n189_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n203_), .B(ori_ori_n185_), .Y(ori_ori_n204_));
  AN2        o182(.A(i_12_), .B(i_5_), .Y(ori_ori_n205_));
  NO2        o183(.A(i_5_), .B(i_10_), .Y(ori_ori_n206_));
  NO3        o184(.A(ori_ori_n73_), .B(ori_ori_n45_), .C(i_9_), .Y(ori_ori_n207_));
  NO2        o185(.A(i_11_), .B(i_12_), .Y(ori_ori_n208_));
  NAi21      o186(.An(i_13_), .B(i_0_), .Y(ori_ori_n209_));
  NO3        o187(.A(i_1_), .B(i_12_), .C(ori_ori_n73_), .Y(ori_ori_n210_));
  NO2        o188(.A(i_0_), .B(i_11_), .Y(ori_ori_n211_));
  AN2        o189(.A(i_1_), .B(i_6_), .Y(ori_ori_n212_));
  NAi21      o190(.An(i_9_), .B(i_4_), .Y(ori_ori_n213_));
  OR2        o191(.A(i_13_), .B(i_10_), .Y(ori_ori_n214_));
  NO3        o192(.A(ori_ori_n214_), .B(ori_ori_n97_), .C(ori_ori_n213_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n216_));
  NA2        o194(.A(ori_ori_n167_), .B(ori_ori_n216_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n217_), .B(ori_ori_n175_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n128_), .B(i_10_), .Y(ori_ori_n219_));
  NA3        o197(.A(ori_ori_n155_), .B(ori_ori_n56_), .C(i_2_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n220_), .B(ori_ori_n219_), .Y(ori_ori_n221_));
  INV        o199(.A(ori_ori_n221_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n222_), .B(ori_ori_n165_), .Y(ori_ori_n223_));
  NO3        o201(.A(ori_ori_n223_), .B(ori_ori_n218_), .C(ori_ori_n204_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n65_), .B(i_13_), .Y(ori_ori_n225_));
  NO2        o203(.A(i_10_), .B(i_9_), .Y(ori_ori_n226_));
  NAi21      o204(.An(i_12_), .B(i_8_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n227_), .B(i_3_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n162_), .B(ori_ori_n84_), .Y(ori_ori_n229_));
  NA2        o207(.A(i_8_), .B(i_9_), .Y(ori_ori_n230_));
  NA2        o208(.A(ori_ori_n167_), .B(ori_ori_n131_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NA3        o210(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n233_));
  NA4        o211(.A(ori_ori_n116_), .B(ori_ori_n96_), .C(ori_ori_n71_), .D(ori_ori_n23_), .Y(ori_ori_n234_));
  NO2        o212(.A(ori_ori_n234_), .B(ori_ori_n233_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n235_), .B(ori_ori_n232_), .Y(ori_ori_n236_));
  NA2        o214(.A(ori_ori_n83_), .B(i_13_), .Y(ori_ori_n237_));
  NO3        o215(.A(i_4_), .B(ori_ori_n45_), .C(i_8_), .Y(ori_ori_n238_));
  NO2        o216(.A(i_6_), .B(i_7_), .Y(ori_ori_n239_));
  NO2        o217(.A(i_11_), .B(i_1_), .Y(ori_ori_n240_));
  NOi21      o218(.An(i_2_), .B(i_7_), .Y(ori_ori_n241_));
  NO2        o219(.A(i_6_), .B(i_10_), .Y(ori_ori_n242_));
  NA3        o220(.A(ori_ori_n149_), .B(ori_ori_n123_), .C(ori_ori_n108_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n44_), .B(ori_ori_n42_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n119_), .B(i_3_), .Y(ori_ori_n245_));
  NAi31      o223(.An(ori_ori_n244_), .B(ori_ori_n245_), .C(ori_ori_n141_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n246_), .B(ori_ori_n243_), .Y(ori_ori_n247_));
  INV        o225(.A(ori_ori_n247_), .Y(ori_ori_n248_));
  NAi21      o226(.An(ori_ori_n135_), .B(ori_ori_n208_), .Y(ori_ori_n249_));
  NA2        o227(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n170_), .B(ori_ori_n145_), .Y(ori_ori_n251_));
  OAI220     o229(.A0(ori_ori_n251_), .A1(ori_ori_n220_), .B0(ori_ori_n250_), .B1(ori_ori_n237_), .Y(ori_ori_n252_));
  INV        o230(.A(ori_ori_n252_), .Y(ori_ori_n253_));
  NA3        o231(.A(ori_ori_n253_), .B(ori_ori_n248_), .C(ori_ori_n236_), .Y(ori_ori_n254_));
  NA2        o232(.A(ori_ori_n205_), .B(ori_ori_n140_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n193_), .B(ori_ori_n186_), .Y(ori_ori_n256_));
  OR2        o234(.A(ori_ori_n255_), .B(ori_ori_n256_), .Y(ori_ori_n257_));
  AOI210     o235(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n215_), .Y(ori_ori_n258_));
  NA2        o236(.A(ori_ori_n258_), .B(ori_ori_n257_), .Y(ori_ori_n259_));
  NO2        o237(.A(i_12_), .B(ori_ori_n128_), .Y(ori_ori_n260_));
  NA2        o238(.A(ori_ori_n42_), .B(i_10_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n119_), .B(i_5_), .Y(ori_ori_n262_));
  NA3        o240(.A(ori_ori_n136_), .B(ori_ori_n63_), .C(ori_ori_n42_), .Y(ori_ori_n263_));
  NA2        o241(.A(ori_ori_n167_), .B(ori_ori_n72_), .Y(ori_ori_n264_));
  NO2        o242(.A(ori_ori_n263_), .B(ori_ori_n264_), .Y(ori_ori_n265_));
  NA2        o243(.A(ori_ori_n139_), .B(ori_ori_n138_), .Y(ori_ori_n266_));
  NA2        o244(.A(ori_ori_n226_), .B(i_4_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n266_), .B(ori_ori_n267_), .Y(ori_ori_n268_));
  AOI210     o246(.A0(ori_ori_n187_), .A1(ori_ori_n44_), .B0(ori_ori_n190_), .Y(ori_ori_n269_));
  NA2        o247(.A(i_0_), .B(ori_ori_n45_), .Y(ori_ori_n270_));
  NA3        o248(.A(ori_ori_n260_), .B(ori_ori_n166_), .C(ori_ori_n270_), .Y(ori_ori_n271_));
  NO2        o249(.A(ori_ori_n269_), .B(ori_ori_n271_), .Y(ori_ori_n272_));
  NO3        o250(.A(ori_ori_n272_), .B(ori_ori_n268_), .C(ori_ori_n265_), .Y(ori_ori_n273_));
  NOi21      o251(.An(i_10_), .B(i_6_), .Y(ori_ori_n274_));
  OR2        o252(.A(i_2_), .B(i_5_), .Y(ori_ori_n275_));
  OR2        o253(.A(ori_ori_n275_), .B(ori_ori_n212_), .Y(ori_ori_n276_));
  INV        o254(.A(ori_ori_n148_), .Y(ori_ori_n277_));
  AOI210     o255(.A0(ori_ori_n277_), .A1(ori_ori_n276_), .B0(ori_ori_n249_), .Y(ori_ori_n278_));
  INV        o256(.A(ori_ori_n278_), .Y(ori_ori_n279_));
  NA2        o257(.A(ori_ori_n279_), .B(ori_ori_n273_), .Y(ori_ori_n280_));
  NO3        o258(.A(ori_ori_n280_), .B(ori_ori_n259_), .C(ori_ori_n254_), .Y(ori_ori_n281_));
  NA4        o259(.A(ori_ori_n281_), .B(ori_ori_n224_), .C(ori_ori_n183_), .D(ori_ori_n161_), .Y(ori7));
  NO2        o260(.A(ori_ori_n80_), .B(ori_ori_n49_), .Y(ori_ori_n283_));
  NA2        o261(.A(ori_ori_n242_), .B(ori_ori_n72_), .Y(ori_ori_n284_));
  INV        o262(.A(i_11_), .Y(ori_ori_n285_));
  INV        o263(.A(ori_ori_n115_), .Y(ori_ori_n286_));
  NO2        o264(.A(ori_ori_n286_), .B(ori_ori_n284_), .Y(ori_ori_n287_));
  NA3        o265(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n288_));
  NA2        o266(.A(i_12_), .B(i_8_), .Y(ori_ori_n289_));
  NO2        o267(.A(ori_ori_n89_), .B(ori_ori_n288_), .Y(ori_ori_n290_));
  NA2        o268(.A(i_2_), .B(ori_ori_n73_), .Y(ori_ori_n291_));
  OAI210     o269(.A0(ori_ori_n74_), .A1(ori_ori_n129_), .B0(ori_ori_n130_), .Y(ori_ori_n292_));
  NA2        o270(.A(i_4_), .B(i_8_), .Y(ori_ori_n293_));
  INV        o271(.A(ori_ori_n168_), .Y(ori_ori_n294_));
  NO2        o272(.A(ori_ori_n294_), .B(ori_ori_n291_), .Y(ori_ori_n295_));
  NO4        o273(.A(ori_ori_n295_), .B(ori_ori_n290_), .C(ori_ori_n287_), .D(ori_ori_n283_), .Y(ori_ori_n296_));
  AOI210     o274(.A0(ori_ori_n106_), .A1(ori_ori_n54_), .B0(i_10_), .Y(ori_ori_n297_));
  AOI210     o275(.A0(ori_ori_n297_), .A1(ori_ori_n143_), .B0(ori_ori_n120_), .Y(ori_ori_n298_));
  OR2        o276(.A(i_6_), .B(i_10_), .Y(ori_ori_n299_));
  OR3        o277(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n300_));
  OR2        o278(.A(ori_ori_n298_), .B(ori_ori_n163_), .Y(ori_ori_n301_));
  AOI210     o279(.A0(ori_ori_n301_), .A1(ori_ori_n296_), .B0(ori_ori_n55_), .Y(ori_ori_n302_));
  NOi21      o280(.An(i_11_), .B(i_7_), .Y(ori_ori_n303_));
  AO210      o281(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n304_), .B(ori_ori_n303_), .Y(ori_ori_n305_));
  NA2        o283(.A(ori_ori_n305_), .B(ori_ori_n132_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n306_), .B(ori_ori_n55_), .Y(ori_ori_n307_));
  OR2        o285(.A(ori_ori_n133_), .B(ori_ori_n91_), .Y(ori_ori_n308_));
  NO2        o286(.A(i_1_), .B(i_12_), .Y(ori_ori_n309_));
  NA3        o287(.A(ori_ori_n309_), .B(ori_ori_n92_), .C(ori_ori_n24_), .Y(ori_ori_n310_));
  BUFFER     o288(.A(ori_ori_n310_), .Y(ori_ori_n311_));
  NA2        o289(.A(ori_ori_n311_), .B(ori_ori_n308_), .Y(ori_ori_n312_));
  OAI210     o290(.A0(ori_ori_n312_), .A1(ori_ori_n307_), .B0(i_6_), .Y(ori_ori_n313_));
  NO3        o291(.A(ori_ori_n299_), .B(ori_ori_n142_), .C(ori_ori_n23_), .Y(ori_ori_n314_));
  AOI210     o292(.A0(i_1_), .A1(ori_ori_n158_), .B0(ori_ori_n314_), .Y(ori_ori_n315_));
  NO2        o293(.A(ori_ori_n315_), .B(ori_ori_n42_), .Y(ori_ori_n316_));
  NO2        o294(.A(ori_ori_n44_), .B(i_1_), .Y(ori_ori_n317_));
  NA3        o295(.A(ori_ori_n317_), .B(ori_ori_n162_), .C(ori_ori_n42_), .Y(ori_ori_n318_));
  NO2        o296(.A(ori_ori_n515_), .B(ori_ori_n316_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n143_), .B(ori_ori_n85_), .Y(ori_ori_n320_));
  NO2        o298(.A(ori_ori_n320_), .B(ori_ori_n303_), .Y(ori_ori_n321_));
  NA2        o299(.A(ori_ori_n321_), .B(i_1_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n322_), .B(ori_ori_n300_), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n213_), .B(ori_ori_n73_), .Y(ori_ori_n324_));
  NA2        o302(.A(ori_ori_n323_), .B(ori_ori_n44_), .Y(ori_ori_n325_));
  NA2        o303(.A(i_3_), .B(ori_ori_n128_), .Y(ori_ori_n326_));
  NO2        o304(.A(ori_ori_n142_), .B(ori_ori_n42_), .Y(ori_ori_n327_));
  NO3        o305(.A(ori_ori_n327_), .B(i_2_), .C(ori_ori_n144_), .Y(ori_ori_n328_));
  NO2        o306(.A(ori_ori_n97_), .B(ori_ori_n37_), .Y(ori_ori_n329_));
  NO2        o307(.A(ori_ori_n329_), .B(i_6_), .Y(ori_ori_n330_));
  NO2        o308(.A(ori_ori_n73_), .B(i_9_), .Y(ori_ori_n331_));
  NO2        o309(.A(ori_ori_n331_), .B(ori_ori_n55_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n332_), .B(ori_ori_n309_), .Y(ori_ori_n333_));
  NO4        o311(.A(ori_ori_n333_), .B(ori_ori_n330_), .C(ori_ori_n328_), .D(i_4_), .Y(ori_ori_n334_));
  NA2        o312(.A(i_1_), .B(i_3_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n230_), .B(ori_ori_n80_), .Y(ori_ori_n336_));
  NO2        o314(.A(ori_ori_n327_), .B(ori_ori_n336_), .Y(ori_ori_n337_));
  NO2        o315(.A(ori_ori_n337_), .B(ori_ori_n335_), .Y(ori_ori_n338_));
  NO2        o316(.A(ori_ori_n338_), .B(ori_ori_n334_), .Y(ori_ori_n339_));
  NA4        o317(.A(ori_ori_n339_), .B(ori_ori_n325_), .C(ori_ori_n319_), .D(ori_ori_n313_), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n341_));
  AOI210     o319(.A0(ori_ori_n162_), .A1(ori_ori_n84_), .B0(i_1_), .Y(ori_ori_n342_));
  NO2        o320(.A(ori_ori_n191_), .B(i_2_), .Y(ori_ori_n343_));
  NA2        o321(.A(ori_ori_n343_), .B(ori_ori_n342_), .Y(ori_ori_n344_));
  AOI210     o322(.A0(ori_ori_n344_), .A1(ori_ori_n341_), .B0(i_13_), .Y(ori_ori_n345_));
  OR2        o323(.A(i_11_), .B(i_7_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n241_), .B(ori_ori_n24_), .Y(ori_ori_n347_));
  NA2        o325(.A(ori_ori_n347_), .B(ori_ori_n324_), .Y(ori_ori_n348_));
  NO2        o326(.A(ori_ori_n348_), .B(i_13_), .Y(ori_ori_n349_));
  INV        o327(.A(ori_ori_n349_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n284_), .B(ori_ori_n42_), .Y(ori_ori_n351_));
  NA2        o329(.A(ori_ori_n105_), .B(i_13_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n352_), .B(ori_ori_n342_), .Y(ori_ori_n353_));
  INV        o331(.A(i_7_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n79_), .B(ori_ori_n86_), .Y(ori_ori_n355_));
  NO2        o333(.A(ori_ori_n355_), .B(ori_ori_n289_), .Y(ori_ori_n356_));
  NO3        o334(.A(ori_ori_n356_), .B(ori_ori_n353_), .C(ori_ori_n351_), .Y(ori_ori_n357_));
  OR2        o335(.A(i_11_), .B(i_6_), .Y(ori_ori_n358_));
  NA2        o336(.A(i_12_), .B(i_7_), .Y(ori_ori_n359_));
  NO2        o337(.A(ori_ori_n359_), .B(ori_ori_n358_), .Y(ori_ori_n360_));
  NAi21      o338(.An(i_11_), .B(i_12_), .Y(ori_ori_n361_));
  NOi41      o339(.An(ori_ori_n93_), .B(ori_ori_n361_), .C(i_13_), .D(ori_ori_n73_), .Y(ori_ori_n362_));
  NO2        o340(.A(i_6_), .B(ori_ori_n293_), .Y(ori_ori_n363_));
  AOI210     o341(.A0(ori_ori_n363_), .A1(ori_ori_n170_), .B0(ori_ori_n362_), .Y(ori_ori_n364_));
  INV        o342(.A(ori_ori_n364_), .Y(ori_ori_n365_));
  OAI210     o343(.A0(ori_ori_n365_), .A1(ori_ori_n360_), .B0(ori_ori_n55_), .Y(ori_ori_n366_));
  NO2        o344(.A(i_2_), .B(i_12_), .Y(ori_ori_n367_));
  NA2        o345(.A(ori_ori_n190_), .B(ori_ori_n367_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n192_), .B(ori_ori_n190_), .Y(ori_ori_n369_));
  NA2        o347(.A(ori_ori_n369_), .B(ori_ori_n368_), .Y(ori_ori_n370_));
  NA2        o348(.A(ori_ori_n370_), .B(ori_ori_n43_), .Y(ori_ori_n371_));
  NA4        o349(.A(ori_ori_n371_), .B(ori_ori_n366_), .C(ori_ori_n357_), .D(ori_ori_n350_), .Y(ori_ori_n372_));
  OR4        o350(.A(ori_ori_n372_), .B(ori_ori_n345_), .C(ori_ori_n340_), .D(ori_ori_n302_), .Y(ori5));
  NA2        o351(.A(ori_ori_n321_), .B(ori_ori_n164_), .Y(ori_ori_n374_));
  AN2        o352(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n375_));
  NA2        o353(.A(ori_ori_n375_), .B(ori_ori_n367_), .Y(ori_ori_n376_));
  NO2        o354(.A(ori_ori_n289_), .B(i_11_), .Y(ori_ori_n377_));
  NA2        o355(.A(ori_ori_n74_), .B(ori_ori_n377_), .Y(ori_ori_n378_));
  NA3        o356(.A(ori_ori_n378_), .B(ori_ori_n376_), .C(ori_ori_n374_), .Y(ori_ori_n379_));
  NO3        o357(.A(i_11_), .B(ori_ori_n143_), .C(i_13_), .Y(ori_ori_n380_));
  NO2        o358(.A(ori_ori_n102_), .B(ori_ori_n23_), .Y(ori_ori_n381_));
  NA2        o359(.A(i_12_), .B(ori_ori_n381_), .Y(ori_ori_n382_));
  INV        o360(.A(ori_ori_n382_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n383_), .B(ori_ori_n379_), .Y(ori_ori_n384_));
  INV        o362(.A(ori_ori_n123_), .Y(ori_ori_n385_));
  INV        o363(.A(ori_ori_n149_), .Y(ori_ori_n386_));
  NO2        o364(.A(ori_ori_n343_), .B(ori_ori_n228_), .Y(ori_ori_n387_));
  AOI210     o365(.A0(ori_ori_n387_), .A1(ori_ori_n386_), .B0(ori_ori_n385_), .Y(ori_ori_n388_));
  NO2        o366(.A(ori_ori_n230_), .B(ori_ori_n26_), .Y(ori_ori_n389_));
  NO2        o367(.A(ori_ori_n389_), .B(ori_ori_n216_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n124_), .B(ori_ori_n128_), .Y(ori_ori_n391_));
  OA210      o369(.A0(ori_ori_n305_), .A1(ori_ori_n104_), .B0(i_13_), .Y(ori_ori_n392_));
  NO2        o370(.A(ori_ori_n133_), .B(ori_ori_n514_), .Y(ori_ori_n393_));
  NA2        o371(.A(ori_ori_n393_), .B(ori_ori_n216_), .Y(ori_ori_n394_));
  NA2        o372(.A(ori_ori_n85_), .B(ori_ori_n168_), .Y(ori_ori_n395_));
  OAI210     o373(.A0(ori_ori_n395_), .A1(i_11_), .B0(ori_ori_n394_), .Y(ori_ori_n396_));
  NO3        o374(.A(ori_ori_n396_), .B(ori_ori_n392_), .C(ori_ori_n391_), .Y(ori_ori_n397_));
  NO2        o375(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n398_));
  NO2        o376(.A(ori_ori_n398_), .B(ori_ori_n104_), .Y(ori_ori_n399_));
  NO2        o377(.A(ori_ori_n399_), .B(ori_ori_n285_), .Y(ori_ori_n400_));
  NA2        o378(.A(ori_ori_n400_), .B(ori_ori_n36_), .Y(ori_ori_n401_));
  NA4        o379(.A(ori_ori_n401_), .B(ori_ori_n397_), .C(ori_ori_n516_), .D(ori_ori_n384_), .Y(ori6));
  NO2        o380(.A(ori_ori_n137_), .B(ori_ori_n244_), .Y(ori_ori_n403_));
  NO2        o381(.A(ori_ori_n151_), .B(i_9_), .Y(ori_ori_n404_));
  NA2        o382(.A(ori_ori_n404_), .B(ori_ori_n398_), .Y(ori_ori_n405_));
  AOI210     o383(.A0(ori_ori_n405_), .A1(ori_ori_n256_), .B0(ori_ori_n125_), .Y(ori_ori_n406_));
  NAi32      o384(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n407_));
  NO2        o385(.A(ori_ori_n358_), .B(ori_ori_n407_), .Y(ori_ori_n408_));
  OR2        o386(.A(ori_ori_n408_), .B(ori_ori_n406_), .Y(ori_ori_n409_));
  NO2        o387(.A(ori_ori_n346_), .B(i_2_), .Y(ori_ori_n410_));
  NA2        o388(.A(ori_ori_n45_), .B(ori_ori_n37_), .Y(ori_ori_n411_));
  INV        o389(.A(ori_ori_n411_), .Y(ori_ori_n412_));
  NA2        o390(.A(ori_ori_n412_), .B(ori_ori_n410_), .Y(ori_ori_n413_));
  BUFFER     o391(.A(ori_ori_n305_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n414_), .B(ori_ori_n117_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n415_), .B(ori_ori_n413_), .Y(ori_ori_n416_));
  NA2        o394(.A(ori_ori_n403_), .B(ori_ori_n354_), .Y(ori_ori_n417_));
  NA3        o395(.A(ori_ori_n195_), .B(ori_ori_n145_), .C(ori_ori_n117_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n207_), .B(ori_ori_n62_), .Y(ori_ori_n419_));
  NA4        o397(.A(ori_ori_n419_), .B(ori_ori_n418_), .C(ori_ori_n417_), .D(ori_ori_n292_), .Y(ori_ori_n420_));
  NA2        o398(.A(ori_ori_n228_), .B(ori_ori_n226_), .Y(ori_ori_n421_));
  NO2        o399(.A(ori_ori_n299_), .B(ori_ori_n86_), .Y(ori_ori_n422_));
  OAI210     o400(.A0(ori_ori_n422_), .A1(ori_ori_n94_), .B0(ori_ori_n211_), .Y(ori_ori_n423_));
  INV        o401(.A(ori_ori_n276_), .Y(ori_ori_n424_));
  NA2        o402(.A(ori_ori_n424_), .B(ori_ori_n172_), .Y(ori_ori_n425_));
  NA3        o403(.A(ori_ori_n425_), .B(ori_ori_n423_), .C(ori_ori_n421_), .Y(ori_ori_n426_));
  NO4        o404(.A(ori_ori_n426_), .B(ori_ori_n420_), .C(ori_ori_n416_), .D(ori_ori_n409_), .Y(ori_ori_n427_));
  NA2        o405(.A(ori_ori_n427_), .B(ori_ori_n203_), .Y(ori3));
  NA2        o406(.A(i_12_), .B(i_10_), .Y(ori_ori_n429_));
  NO2        o407(.A(i_11_), .B(ori_ori_n143_), .Y(ori_ori_n430_));
  NA3        o408(.A(ori_ori_n418_), .B(ori_ori_n292_), .C(ori_ori_n194_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n431_), .B(ori_ori_n40_), .Y(ori_ori_n432_));
  NOi21      o410(.An(ori_ori_n83_), .B(ori_ori_n390_), .Y(ori_ori_n433_));
  NO2        o411(.A(ori_ori_n308_), .B(ori_ori_n230_), .Y(ori_ori_n434_));
  AN2        o412(.A(ori_ori_n229_), .B(ori_ori_n50_), .Y(ori_ori_n435_));
  NO3        o413(.A(ori_ori_n435_), .B(ori_ori_n434_), .C(ori_ori_n433_), .Y(ori_ori_n436_));
  AOI210     o414(.A0(ori_ori_n436_), .A1(ori_ori_n432_), .B0(ori_ori_n45_), .Y(ori_ori_n437_));
  NO4        o415(.A(ori_ori_n199_), .B(ori_ori_n205_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n438_));
  NA2        o416(.A(ori_ori_n125_), .B(ori_ori_n274_), .Y(ori_ori_n439_));
  NOi21      o417(.An(ori_ori_n439_), .B(ori_ori_n438_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n440_), .B(ori_ori_n55_), .Y(ori_ori_n441_));
  NOi21      o419(.An(i_5_), .B(i_9_), .Y(ori_ori_n442_));
  NA2        o420(.A(ori_ori_n442_), .B(ori_ori_n225_), .Y(ori_ori_n443_));
  BUFFER     o421(.A(ori_ori_n162_), .Y(ori_ori_n444_));
  NA2        o422(.A(ori_ori_n444_), .B(ori_ori_n240_), .Y(ori_ori_n445_));
  NO2        o423(.A(ori_ori_n445_), .B(ori_ori_n443_), .Y(ori_ori_n446_));
  NO3        o424(.A(ori_ori_n446_), .B(ori_ori_n441_), .C(ori_ori_n437_), .Y(ori_ori_n447_));
  NO4        o425(.A(ori_ori_n275_), .B(i_12_), .C(ori_ori_n214_), .D(ori_ori_n212_), .Y(ori_ori_n448_));
  NA2        o426(.A(ori_ori_n448_), .B(i_11_), .Y(ori_ori_n449_));
  NA2        o427(.A(ori_ori_n380_), .B(ori_ori_n173_), .Y(ori_ori_n450_));
  NO2        o428(.A(ori_ori_n74_), .B(ori_ori_n52_), .Y(ori_ori_n451_));
  NO2        o429(.A(ori_ori_n451_), .B(ori_ori_n450_), .Y(ori_ori_n452_));
  NO2        o430(.A(ori_ori_n153_), .B(ori_ori_n118_), .Y(ori_ori_n453_));
  INV        o431(.A(ori_ori_n261_), .Y(ori_ori_n454_));
  NO4        o432(.A(ori_ori_n95_), .B(ori_ori_n52_), .C(ori_ori_n326_), .D(i_5_), .Y(ori_ori_n455_));
  AO220      o433(.A0(ori_ori_n455_), .A1(ori_ori_n454_), .B0(ori_ori_n453_), .B1(i_6_), .Y(ori_ori_n456_));
  NO2        o434(.A(ori_ori_n456_), .B(ori_ori_n452_), .Y(ori_ori_n457_));
  NA2        o435(.A(ori_ori_n457_), .B(ori_ori_n449_), .Y(ori_ori_n458_));
  NO2        o436(.A(ori_ori_n87_), .B(ori_ori_n37_), .Y(ori_ori_n459_));
  NA2        o437(.A(i_11_), .B(i_9_), .Y(ori_ori_n460_));
  NO3        o438(.A(i_12_), .B(ori_ori_n460_), .C(ori_ori_n291_), .Y(ori_ori_n461_));
  AN2        o439(.A(ori_ori_n461_), .B(ori_ori_n459_), .Y(ori_ori_n462_));
  NO2        o440(.A(ori_ori_n460_), .B(ori_ori_n65_), .Y(ori_ori_n463_));
  INV        o441(.A(ori_ori_n210_), .Y(ori_ori_n464_));
  NO2        o442(.A(ori_ori_n464_), .B(ori_ori_n443_), .Y(ori_ori_n465_));
  NO2        o443(.A(ori_ori_n465_), .B(ori_ori_n462_), .Y(ori_ori_n466_));
  INV        o444(.A(ori_ori_n466_), .Y(ori_ori_n467_));
  NO2        o445(.A(ori_ori_n429_), .B(ori_ori_n171_), .Y(ori_ori_n468_));
  OA210      o446(.A0(ori_ori_n239_), .A1(ori_ori_n139_), .B0(ori_ori_n238_), .Y(ori_ori_n469_));
  OAI210     o447(.A0(ori_ori_n469_), .A1(ori_ori_n468_), .B0(ori_ori_n463_), .Y(ori_ori_n470_));
  NA2        o448(.A(ori_ori_n347_), .B(ori_ori_n262_), .Y(ori_ori_n471_));
  NAi21      o449(.An(i_9_), .B(i_5_), .Y(ori_ori_n472_));
  NO2        o450(.A(ori_ori_n472_), .B(ori_ori_n209_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n473_), .B(ori_ori_n305_), .Y(ori_ori_n474_));
  OAI220     o452(.A0(ori_ori_n474_), .A1(ori_ori_n73_), .B0(ori_ori_n471_), .B1(ori_ori_n124_), .Y(ori_ori_n475_));
  NO2        o453(.A(ori_ori_n475_), .B(ori_ori_n259_), .Y(ori_ori_n476_));
  NA2        o454(.A(ori_ori_n476_), .B(ori_ori_n470_), .Y(ori_ori_n477_));
  NO3        o455(.A(ori_ori_n477_), .B(ori_ori_n467_), .C(ori_ori_n458_), .Y(ori_ori_n478_));
  NO3        o456(.A(ori_ori_n134_), .B(ori_ori_n205_), .C(i_0_), .Y(ori_ori_n479_));
  OAI210     o457(.A0(ori_ori_n479_), .A1(ori_ori_n67_), .B0(i_13_), .Y(ori_ori_n480_));
  INV        o458(.A(ori_ori_n480_), .Y(ori_ori_n481_));
  NO2        o459(.A(i_0_), .B(i_12_), .Y(ori_ori_n482_));
  NA2        o460(.A(ori_ori_n482_), .B(ori_ori_n469_), .Y(ori_ori_n483_));
  NA3        o461(.A(ori_ori_n206_), .B(ori_ori_n123_), .C(ori_ori_n122_), .Y(ori_ori_n484_));
  INV        o462(.A(ori_ori_n484_), .Y(ori_ori_n485_));
  NO3        o463(.A(ori_ori_n460_), .B(ori_ori_n136_), .C(ori_ori_n127_), .Y(ori_ori_n486_));
  NO2        o464(.A(ori_ori_n486_), .B(ori_ori_n485_), .Y(ori_ori_n487_));
  NA3        o465(.A(ori_ori_n487_), .B(ori_ori_n243_), .C(ori_ori_n483_), .Y(ori_ori_n488_));
  NO2        o466(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n489_));
  NA3        o467(.A(ori_ori_n430_), .B(ori_ori_n92_), .C(ori_ori_n102_), .Y(ori_ori_n490_));
  INV        o468(.A(ori_ori_n490_), .Y(ori_ori_n491_));
  NA2        o469(.A(ori_ori_n491_), .B(ori_ori_n489_), .Y(ori_ori_n492_));
  NAi21      o470(.An(i_10_), .B(ori_ori_n147_), .Y(ori_ori_n493_));
  NO4        o471(.A(ori_ori_n146_), .B(ori_ori_n134_), .C(i_0_), .D(i_12_), .Y(ori_ori_n494_));
  NA2        o472(.A(ori_ori_n494_), .B(ori_ori_n493_), .Y(ori_ori_n495_));
  NA2        o473(.A(ori_ori_n495_), .B(ori_ori_n492_), .Y(ori_ori_n496_));
  NO3        o474(.A(ori_ori_n496_), .B(ori_ori_n488_), .C(ori_ori_n481_), .Y(ori_ori_n497_));
  NA2        o475(.A(ori_ori_n410_), .B(ori_ori_n37_), .Y(ori_ori_n498_));
  NA2        o476(.A(ori_ori_n498_), .B(ori_ori_n298_), .Y(ori_ori_n499_));
  NA2        o477(.A(ori_ori_n499_), .B(ori_ori_n132_), .Y(ori_ori_n500_));
  NAi31      o478(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n501_));
  NO2        o479(.A(ori_ori_n62_), .B(ori_ori_n501_), .Y(ori_ori_n502_));
  AOI210     o480(.A0(ori_ori_n502_), .A1(ori_ori_n45_), .B0(ori_ori_n448_), .Y(ori_ori_n503_));
  AOI210     o481(.A0(ori_ori_n503_), .A1(ori_ori_n500_), .B0(ori_ori_n65_), .Y(ori_ori_n504_));
  INV        o482(.A(ori_ori_n202_), .Y(ori_ori_n505_));
  NO2        o483(.A(ori_ori_n505_), .B(ori_ori_n385_), .Y(ori_ori_n506_));
  NO3        o484(.A(ori_ori_n53_), .B(ori_ori_n52_), .C(i_4_), .Y(ori_ori_n507_));
  NA2        o485(.A(ori_ori_n169_), .B(ori_ori_n507_), .Y(ori_ori_n508_));
  NO2        o486(.A(ori_ori_n508_), .B(ori_ori_n361_), .Y(ori_ori_n509_));
  NO3        o487(.A(ori_ori_n509_), .B(ori_ori_n506_), .C(ori_ori_n504_), .Y(ori_ori_n510_));
  NA4        o488(.A(ori_ori_n510_), .B(ori_ori_n497_), .C(ori_ori_n478_), .D(ori_ori_n447_), .Y(ori4));
  INV        o489(.A(i_8_), .Y(ori_ori_n514_));
  INV        o490(.A(ori_ori_n318_), .Y(ori_ori_n515_));
  INV        o491(.A(ori_ori_n388_), .Y(ori_ori_n516_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  OAI210     m028(.A0(mai_mai_n50_), .A1(i_3_), .B0(mai_mai_n48_), .Y(mai_mai_n51_));
  AOI210     m029(.A0(mai_mai_n51_), .A1(mai_mai_n47_), .B0(mai_mai_n46_), .Y(mai_mai_n52_));
  NA2        m030(.A(i_0_), .B(i_2_), .Y(mai_mai_n53_));
  NA2        m031(.A(i_7_), .B(i_9_), .Y(mai_mai_n54_));
  NA2        m032(.A(mai_mai_n52_), .B(mai_mai_n45_), .Y(mai_mai_n55_));
  NA3        m033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n56_));
  NO2        m034(.A(i_1_), .B(i_6_), .Y(mai_mai_n57_));
  NA2        m035(.A(i_8_), .B(i_7_), .Y(mai_mai_n58_));
  OAI210     m036(.A0(mai_mai_n58_), .A1(mai_mai_n57_), .B0(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n59_), .B(i_12_), .Y(mai_mai_n60_));
  NAi21      m038(.An(i_2_), .B(i_7_), .Y(mai_mai_n61_));
  INV        m039(.A(i_1_), .Y(mai_mai_n62_));
  NA2        m040(.A(i_1_), .B(i_10_), .Y(mai_mai_n63_));
  NO2        m041(.A(mai_mai_n63_), .B(i_6_), .Y(mai_mai_n64_));
  NAi21      m042(.An(mai_mai_n64_), .B(mai_mai_n60_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n66_));
  NA2        m044(.A(i_1_), .B(i_6_), .Y(mai_mai_n67_));
  NO2        m045(.A(mai_mai_n67_), .B(mai_mai_n25_), .Y(mai_mai_n68_));
  INV        m046(.A(i_0_), .Y(mai_mai_n69_));
  NAi21      m047(.An(i_5_), .B(i_10_), .Y(mai_mai_n70_));
  NA2        m048(.A(i_5_), .B(i_9_), .Y(mai_mai_n71_));
  AOI210     m049(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n69_), .Y(mai_mai_n72_));
  INV        m050(.A(mai_mai_n72_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n72_), .A1(mai_mai_n65_), .B0(i_0_), .Y(mai_mai_n74_));
  NA2        m052(.A(i_12_), .B(i_5_), .Y(mai_mai_n75_));
  NA2        m053(.A(i_2_), .B(i_8_), .Y(mai_mai_n76_));
  NO2        m054(.A(i_3_), .B(i_9_), .Y(mai_mai_n77_));
  NO2        m055(.A(i_3_), .B(i_7_), .Y(mai_mai_n78_));
  NO3        m056(.A(mai_mai_n78_), .B(mai_mai_n77_), .C(mai_mai_n62_), .Y(mai_mai_n79_));
  INV        m057(.A(i_6_), .Y(mai_mai_n80_));
  OR4        m058(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n81_));
  INV        m059(.A(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m060(.A(i_2_), .B(i_7_), .Y(mai_mai_n83_));
  NA2        m061(.A(mai_mai_n79_), .B(i_2_), .Y(mai_mai_n84_));
  NAi21      m062(.An(i_6_), .B(i_10_), .Y(mai_mai_n85_));
  NA2        m063(.A(i_2_), .B(i_6_), .Y(mai_mai_n86_));
  NO2        m064(.A(mai_mai_n84_), .B(mai_mai_n75_), .Y(mai_mai_n87_));
  AN3        m065(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n88_));
  NAi21      m066(.An(i_6_), .B(i_11_), .Y(mai_mai_n89_));
  NO2        m067(.A(i_5_), .B(i_8_), .Y(mai_mai_n90_));
  NOi21      m068(.An(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n91_));
  AOI220     m069(.A0(mai_mai_n91_), .A1(mai_mai_n61_), .B0(mai_mai_n88_), .B1(mai_mai_n32_), .Y(mai_mai_n92_));
  INV        m070(.A(i_7_), .Y(mai_mai_n93_));
  NO2        m071(.A(i_0_), .B(i_5_), .Y(mai_mai_n94_));
  NA2        m072(.A(i_12_), .B(i_3_), .Y(mai_mai_n95_));
  INV        m073(.A(mai_mai_n95_), .Y(mai_mai_n96_));
  NAi21      m074(.An(i_7_), .B(i_11_), .Y(mai_mai_n97_));
  NO3        m075(.A(mai_mai_n97_), .B(mai_mai_n85_), .C(mai_mai_n53_), .Y(mai_mai_n98_));
  AN2        m076(.A(i_2_), .B(i_10_), .Y(mai_mai_n99_));
  NO2        m077(.A(mai_mai_n99_), .B(i_7_), .Y(mai_mai_n100_));
  OR2        m078(.A(mai_mai_n75_), .B(mai_mai_n57_), .Y(mai_mai_n101_));
  NO2        m079(.A(i_8_), .B(mai_mai_n93_), .Y(mai_mai_n102_));
  NO3        m080(.A(mai_mai_n102_), .B(mai_mai_n101_), .C(mai_mai_n100_), .Y(mai_mai_n103_));
  NA2        m081(.A(i_12_), .B(i_7_), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n62_), .B(mai_mai_n26_), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n105_), .B(i_0_), .Y(mai_mai_n106_));
  NA2        m084(.A(i_11_), .B(i_12_), .Y(mai_mai_n107_));
  OAI210     m085(.A0(mai_mai_n106_), .A1(mai_mai_n104_), .B0(mai_mai_n107_), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n108_), .B(mai_mai_n103_), .Y(mai_mai_n109_));
  NAi31      m087(.An(mai_mai_n98_), .B(mai_mai_n109_), .C(mai_mai_n92_), .Y(mai_mai_n110_));
  NOi21      m088(.An(i_1_), .B(i_5_), .Y(mai_mai_n111_));
  NA2        m089(.A(mai_mai_n111_), .B(i_11_), .Y(mai_mai_n112_));
  NA2        m090(.A(mai_mai_n93_), .B(mai_mai_n37_), .Y(mai_mai_n113_));
  NA2        m091(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n114_), .B(mai_mai_n113_), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n115_), .B(mai_mai_n46_), .Y(mai_mai_n116_));
  NAi21      m094(.An(i_3_), .B(i_8_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n117_), .B(mai_mai_n61_), .Y(mai_mai_n118_));
  BUFFER     m096(.A(mai_mai_n118_), .Y(mai_mai_n119_));
  NO2        m097(.A(i_1_), .B(mai_mai_n80_), .Y(mai_mai_n120_));
  NO2        m098(.A(i_6_), .B(i_5_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n121_), .B(i_3_), .Y(mai_mai_n122_));
  AO210      m100(.A0(mai_mai_n122_), .A1(mai_mai_n47_), .B0(mai_mai_n120_), .Y(mai_mai_n123_));
  OAI220     m101(.A0(mai_mai_n123_), .A1(mai_mai_n97_), .B0(mai_mai_n119_), .B1(mai_mai_n112_), .Y(mai_mai_n124_));
  NO3        m102(.A(mai_mai_n124_), .B(mai_mai_n110_), .C(mai_mai_n87_), .Y(mai_mai_n125_));
  NA3        m103(.A(mai_mai_n125_), .B(mai_mai_n74_), .C(mai_mai_n55_), .Y(mai2));
  NO2        m104(.A(mai_mai_n62_), .B(mai_mai_n37_), .Y(mai_mai_n127_));
  NA2        m105(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n129_));
  NA4        m107(.A(mai_mai_n129_), .B(mai_mai_n73_), .C(mai_mai_n66_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m108(.A(i_8_), .B(i_7_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n131_), .B(i_6_), .Y(mai_mai_n132_));
  NO2        m110(.A(i_12_), .B(i_13_), .Y(mai_mai_n133_));
  NAi21      m111(.An(i_5_), .B(i_11_), .Y(mai_mai_n134_));
  NOi21      m112(.An(mai_mai_n133_), .B(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m113(.A(i_0_), .B(i_1_), .Y(mai_mai_n136_));
  NA2        m114(.A(i_2_), .B(i_3_), .Y(mai_mai_n137_));
  NO2        m115(.A(mai_mai_n137_), .B(i_4_), .Y(mai_mai_n138_));
  NA3        m116(.A(mai_mai_n138_), .B(mai_mai_n136_), .C(mai_mai_n135_), .Y(mai_mai_n139_));
  NA2        m117(.A(i_1_), .B(i_5_), .Y(mai_mai_n140_));
  NO2        m118(.A(mai_mai_n69_), .B(mai_mai_n46_), .Y(mai_mai_n141_));
  NA2        m119(.A(mai_mai_n141_), .B(mai_mai_n36_), .Y(mai_mai_n142_));
  NO3        m120(.A(mai_mai_n142_), .B(mai_mai_n140_), .C(i_13_), .Y(mai_mai_n143_));
  OR2        m121(.A(i_0_), .B(i_1_), .Y(mai_mai_n144_));
  NO3        m122(.A(mai_mai_n144_), .B(mai_mai_n75_), .C(i_13_), .Y(mai_mai_n145_));
  NAi32      m123(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n146_));
  NAi21      m124(.An(mai_mai_n146_), .B(mai_mai_n145_), .Y(mai_mai_n147_));
  NOi21      m125(.An(i_4_), .B(i_10_), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n40_), .Y(mai_mai_n149_));
  NO2        m127(.A(i_3_), .B(i_5_), .Y(mai_mai_n150_));
  NO3        m128(.A(mai_mai_n69_), .B(i_2_), .C(i_1_), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n151_), .B(mai_mai_n150_), .Y(mai_mai_n152_));
  OAI210     m130(.A0(mai_mai_n152_), .A1(mai_mai_n149_), .B0(mai_mai_n147_), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n153_), .B(mai_mai_n143_), .Y(mai_mai_n154_));
  NO2        m132(.A(mai_mai_n154_), .B(mai_mai_n132_), .Y(mai_mai_n155_));
  NA2        m133(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n156_));
  NOi21      m134(.An(i_4_), .B(i_9_), .Y(mai_mai_n157_));
  NOi21      m135(.An(i_11_), .B(i_13_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  OR2        m137(.A(mai_mai_n159_), .B(mai_mai_n156_), .Y(mai_mai_n160_));
  NO2        m138(.A(i_4_), .B(i_5_), .Y(mai_mai_n161_));
  NAi21      m139(.An(i_12_), .B(i_11_), .Y(mai_mai_n162_));
  NA3        m140(.A(mai_mai_n883_), .B(mai_mai_n161_), .C(mai_mai_n77_), .Y(mai_mai_n163_));
  NA2        m141(.A(mai_mai_n163_), .B(mai_mai_n160_), .Y(mai_mai_n164_));
  NO2        m142(.A(mai_mai_n69_), .B(mai_mai_n62_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n46_), .Y(mai_mai_n166_));
  NA2        m144(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n167_));
  NAi31      m145(.An(mai_mai_n167_), .B(mai_mai_n77_), .C(i_11_), .Y(mai_mai_n168_));
  NA2        m146(.A(i_3_), .B(i_5_), .Y(mai_mai_n169_));
  AOI210     m147(.A0(mai_mai_n159_), .A1(mai_mai_n168_), .B0(mai_mai_n166_), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n69_), .B(i_5_), .Y(mai_mai_n171_));
  NA2        m149(.A(mai_mai_n171_), .B(mai_mai_n44_), .Y(mai_mai_n172_));
  NO2        m150(.A(i_2_), .B(i_1_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n173_), .B(i_3_), .Y(mai_mai_n174_));
  NAi21      m152(.An(i_4_), .B(i_12_), .Y(mai_mai_n175_));
  NO3        m153(.A(mai_mai_n175_), .B(mai_mai_n174_), .C(mai_mai_n172_), .Y(mai_mai_n176_));
  NO3        m154(.A(mai_mai_n176_), .B(mai_mai_n170_), .C(mai_mai_n164_), .Y(mai_mai_n177_));
  INV        m155(.A(i_8_), .Y(mai_mai_n178_));
  NO2        m156(.A(mai_mai_n178_), .B(i_7_), .Y(mai_mai_n179_));
  NA2        m157(.A(mai_mai_n179_), .B(i_6_), .Y(mai_mai_n180_));
  NO3        m158(.A(i_3_), .B(mai_mai_n80_), .C(mai_mai_n48_), .Y(mai_mai_n181_));
  NA2        m159(.A(mai_mai_n181_), .B(mai_mai_n102_), .Y(mai_mai_n182_));
  NO3        m160(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n183_));
  NA3        m161(.A(mai_mai_n183_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n184_));
  NO2        m162(.A(i_11_), .B(mai_mai_n182_), .Y(mai_mai_n185_));
  NO2        m163(.A(i_3_), .B(i_8_), .Y(mai_mai_n186_));
  NO3        m164(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n187_));
  NA3        m165(.A(mai_mai_n187_), .B(mai_mai_n186_), .C(mai_mai_n40_), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n94_), .B(mai_mai_n57_), .Y(mai_mai_n189_));
  NO2        m167(.A(i_13_), .B(i_9_), .Y(mai_mai_n190_));
  NA3        m168(.A(mai_mai_n190_), .B(i_6_), .C(mai_mai_n178_), .Y(mai_mai_n191_));
  BUFFER     m169(.A(mai_mai_n191_), .Y(mai_mai_n192_));
  NO2        m170(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n193_));
  NO3        m171(.A(i_0_), .B(i_2_), .C(mai_mai_n62_), .Y(mai_mai_n194_));
  NA3        m172(.A(mai_mai_n194_), .B(mai_mai_n193_), .C(i_10_), .Y(mai_mai_n195_));
  OAI220     m173(.A0(mai_mai_n195_), .A1(mai_mai_n192_), .B0(mai_mai_n57_), .B1(mai_mai_n188_), .Y(mai_mai_n196_));
  AOI210     m174(.A0(mai_mai_n196_), .A1(i_7_), .B0(mai_mai_n185_), .Y(mai_mai_n197_));
  OAI220     m175(.A0(mai_mai_n197_), .A1(i_4_), .B0(mai_mai_n180_), .B1(mai_mai_n177_), .Y(mai_mai_n198_));
  NA3        m176(.A(i_13_), .B(mai_mai_n178_), .C(i_10_), .Y(mai_mai_n199_));
  NO2        m177(.A(mai_mai_n199_), .B(i_12_), .Y(mai_mai_n200_));
  NA2        m178(.A(i_0_), .B(i_5_), .Y(mai_mai_n201_));
  OAI220     m179(.A0(mai_mai_n80_), .A1(mai_mai_n174_), .B0(mai_mai_n166_), .B1(mai_mai_n122_), .Y(mai_mai_n202_));
  NAi31      m180(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n203_));
  INV        m181(.A(i_13_), .Y(mai_mai_n204_));
  NO2        m182(.A(i_12_), .B(mai_mai_n204_), .Y(mai_mai_n205_));
  NA3        m183(.A(mai_mai_n205_), .B(mai_mai_n183_), .C(mai_mai_n181_), .Y(mai_mai_n206_));
  INV        m184(.A(mai_mai_n206_), .Y(mai_mai_n207_));
  AOI220     m185(.A0(mai_mai_n207_), .A1(mai_mai_n131_), .B0(mai_mai_n202_), .B1(mai_mai_n200_), .Y(mai_mai_n208_));
  NO2        m186(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n169_), .B(i_4_), .Y(mai_mai_n210_));
  NA2        m188(.A(mai_mai_n210_), .B(mai_mai_n209_), .Y(mai_mai_n211_));
  OR2        m189(.A(i_8_), .B(i_7_), .Y(mai_mai_n212_));
  NO2        m190(.A(mai_mai_n212_), .B(mai_mai_n80_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n53_), .B(i_1_), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n214_), .B(mai_mai_n213_), .Y(mai_mai_n215_));
  INV        m193(.A(i_12_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n44_), .B(mai_mai_n216_), .Y(mai_mai_n217_));
  NO3        m195(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n218_));
  NA2        m196(.A(i_2_), .B(i_1_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n215_), .B(mai_mai_n211_), .Y(mai_mai_n220_));
  NO3        m198(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n221_));
  NAi21      m199(.An(i_4_), .B(i_3_), .Y(mai_mai_n222_));
  NO2        m200(.A(i_0_), .B(i_6_), .Y(mai_mai_n223_));
  NOi41      m201(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n224_), .B(mai_mai_n223_), .Y(mai_mai_n225_));
  NO2        m203(.A(mai_mai_n219_), .B(mai_mai_n169_), .Y(mai_mai_n226_));
  NAi21      m204(.An(mai_mai_n225_), .B(mai_mai_n226_), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n227_), .Y(mai_mai_n228_));
  AOI210     m206(.A0(mai_mai_n228_), .A1(mai_mai_n40_), .B0(mai_mai_n220_), .Y(mai_mai_n229_));
  NO2        m207(.A(i_11_), .B(mai_mai_n204_), .Y(mai_mai_n230_));
  NOi21      m208(.An(i_1_), .B(i_6_), .Y(mai_mai_n231_));
  NAi21      m209(.An(i_3_), .B(i_7_), .Y(mai_mai_n232_));
  NA2        m210(.A(mai_mai_n216_), .B(i_9_), .Y(mai_mai_n233_));
  NA2        m211(.A(mai_mai_n69_), .B(i_5_), .Y(mai_mai_n234_));
  NA3        m212(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n235_));
  INV        m213(.A(mai_mai_n132_), .Y(mai_mai_n236_));
  NA2        m214(.A(mai_mai_n216_), .B(i_13_), .Y(mai_mai_n237_));
  NO2        m215(.A(mai_mai_n237_), .B(mai_mai_n71_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n238_), .B(mai_mai_n236_), .Y(mai_mai_n239_));
  NO2        m217(.A(mai_mai_n212_), .B(mai_mai_n37_), .Y(mai_mai_n240_));
  NA2        m218(.A(i_12_), .B(i_6_), .Y(mai_mai_n241_));
  OR2        m219(.A(i_13_), .B(i_9_), .Y(mai_mai_n242_));
  NO3        m220(.A(mai_mai_n242_), .B(mai_mai_n241_), .C(mai_mai_n48_), .Y(mai_mai_n243_));
  NO2        m221(.A(mai_mai_n222_), .B(i_2_), .Y(mai_mai_n244_));
  NA3        m222(.A(mai_mai_n244_), .B(mai_mai_n243_), .C(mai_mai_n44_), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n230_), .B(i_9_), .Y(mai_mai_n246_));
  OAI210     m224(.A0(mai_mai_n62_), .A1(mai_mai_n246_), .B0(mai_mai_n245_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n141_), .B(mai_mai_n62_), .Y(mai_mai_n248_));
  NO3        m226(.A(i_11_), .B(mai_mai_n204_), .C(mai_mai_n25_), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n232_), .B(i_8_), .Y(mai_mai_n250_));
  NO2        m228(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n250_), .B(mai_mai_n249_), .Y(mai_mai_n252_));
  NA3        m230(.A(i_6_), .B(mai_mai_n240_), .C(mai_mai_n205_), .Y(mai_mai_n253_));
  AOI210     m231(.A0(mai_mai_n253_), .A1(mai_mai_n252_), .B0(mai_mai_n248_), .Y(mai_mai_n254_));
  AOI210     m232(.A0(mai_mai_n247_), .A1(mai_mai_n240_), .B0(mai_mai_n254_), .Y(mai_mai_n255_));
  NA4        m233(.A(mai_mai_n255_), .B(mai_mai_n239_), .C(mai_mai_n229_), .D(mai_mai_n208_), .Y(mai_mai_n256_));
  NO3        m234(.A(i_12_), .B(mai_mai_n204_), .C(mai_mai_n37_), .Y(mai_mai_n257_));
  INV        m235(.A(mai_mai_n257_), .Y(mai_mai_n258_));
  NO3        m236(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n259_));
  NO3        m237(.A(i_0_), .B(i_2_), .C(mai_mai_n62_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n219_), .B(i_0_), .Y(mai_mai_n261_));
  AOI220     m239(.A0(mai_mai_n261_), .A1(mai_mai_n179_), .B0(mai_mai_n260_), .B1(mai_mai_n131_), .Y(mai_mai_n262_));
  NA2        m240(.A(mai_mai_n251_), .B(mai_mai_n26_), .Y(mai_mai_n263_));
  NO2        m241(.A(mai_mai_n263_), .B(mai_mai_n262_), .Y(mai_mai_n264_));
  NA2        m242(.A(i_0_), .B(i_1_), .Y(mai_mai_n265_));
  NO2        m243(.A(mai_mai_n265_), .B(i_2_), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n58_), .B(i_6_), .Y(mai_mai_n267_));
  NA3        m245(.A(mai_mai_n267_), .B(mai_mai_n266_), .C(mai_mai_n150_), .Y(mai_mai_n268_));
  OAI210     m246(.A0(mai_mai_n152_), .A1(mai_mai_n132_), .B0(mai_mai_n268_), .Y(mai_mai_n269_));
  NO2        m247(.A(mai_mai_n269_), .B(mai_mai_n264_), .Y(mai_mai_n270_));
  NO2        m248(.A(i_3_), .B(i_10_), .Y(mai_mai_n271_));
  NA3        m249(.A(mai_mai_n271_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n272_));
  NO2        m250(.A(i_2_), .B(mai_mai_n93_), .Y(mai_mai_n273_));
  NA2        m251(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n274_), .B(i_8_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n275_), .B(mai_mai_n273_), .Y(mai_mai_n276_));
  AN2        m254(.A(i_3_), .B(i_10_), .Y(mai_mai_n277_));
  NA3        m255(.A(mai_mai_n183_), .B(mai_mai_n883_), .C(mai_mai_n161_), .Y(mai_mai_n278_));
  NO2        m256(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n280_));
  OR2        m258(.A(mai_mai_n276_), .B(mai_mai_n272_), .Y(mai_mai_n281_));
  OAI220     m259(.A0(mai_mai_n281_), .A1(i_6_), .B0(mai_mai_n270_), .B1(mai_mai_n258_), .Y(mai_mai_n282_));
  NO4        m260(.A(mai_mai_n282_), .B(mai_mai_n256_), .C(mai_mai_n198_), .D(mai_mai_n155_), .Y(mai_mai_n283_));
  NO3        m261(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n284_));
  NO3        m262(.A(i_6_), .B(mai_mai_n178_), .C(i_7_), .Y(mai_mai_n285_));
  AOI210     m263(.A0(i_1_), .A1(mai_mai_n219_), .B0(mai_mai_n156_), .Y(mai_mai_n286_));
  NO2        m264(.A(i_2_), .B(i_3_), .Y(mai_mai_n287_));
  OR2        m265(.A(i_0_), .B(i_5_), .Y(mai_mai_n288_));
  NA2        m266(.A(mai_mai_n201_), .B(mai_mai_n288_), .Y(mai_mai_n289_));
  NA4        m267(.A(mai_mai_n289_), .B(mai_mai_n213_), .C(mai_mai_n287_), .D(i_1_), .Y(mai_mai_n290_));
  NA3        m268(.A(mai_mai_n261_), .B(mai_mai_n150_), .C(mai_mai_n102_), .Y(mai_mai_n291_));
  NAi21      m269(.An(i_8_), .B(i_7_), .Y(mai_mai_n292_));
  NO2        m270(.A(mai_mai_n292_), .B(i_6_), .Y(mai_mai_n293_));
  NA3        m271(.A(i_2_), .B(mai_mai_n293_), .C(mai_mai_n150_), .Y(mai_mai_n294_));
  NA3        m272(.A(mai_mai_n294_), .B(mai_mai_n291_), .C(mai_mai_n290_), .Y(mai_mai_n295_));
  OAI210     m273(.A0(mai_mai_n295_), .A1(mai_mai_n286_), .B0(i_4_), .Y(mai_mai_n296_));
  NO2        m274(.A(i_12_), .B(i_10_), .Y(mai_mai_n297_));
  NOi21      m275(.An(i_5_), .B(i_0_), .Y(mai_mai_n298_));
  NO3        m276(.A(mai_mai_n274_), .B(mai_mai_n298_), .C(mai_mai_n117_), .Y(mai_mai_n299_));
  NA4        m277(.A(mai_mai_n78_), .B(mai_mai_n36_), .C(mai_mai_n80_), .D(i_8_), .Y(mai_mai_n300_));
  NA2        m278(.A(mai_mai_n299_), .B(mai_mai_n297_), .Y(mai_mai_n301_));
  NO2        m279(.A(i_6_), .B(i_8_), .Y(mai_mai_n302_));
  NOi21      m280(.An(i_0_), .B(i_2_), .Y(mai_mai_n303_));
  AN2        m281(.A(mai_mai_n303_), .B(mai_mai_n302_), .Y(mai_mai_n304_));
  NO2        m282(.A(i_1_), .B(i_7_), .Y(mai_mai_n305_));
  AO220      m283(.A0(mai_mai_n305_), .A1(mai_mai_n304_), .B0(mai_mai_n293_), .B1(mai_mai_n214_), .Y(mai_mai_n306_));
  NA2        m284(.A(mai_mai_n306_), .B(i_4_), .Y(mai_mai_n307_));
  NA3        m285(.A(mai_mai_n307_), .B(mai_mai_n301_), .C(mai_mai_n296_), .Y(mai_mai_n308_));
  NO3        m286(.A(mai_mai_n212_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n309_));
  NO3        m287(.A(mai_mai_n292_), .B(i_2_), .C(i_1_), .Y(mai_mai_n310_));
  OAI210     m288(.A0(mai_mai_n310_), .A1(mai_mai_n309_), .B0(i_6_), .Y(mai_mai_n311_));
  NA2        m289(.A(mai_mai_n231_), .B(mai_mai_n273_), .Y(mai_mai_n312_));
  AOI210     m290(.A0(mai_mai_n312_), .A1(mai_mai_n311_), .B0(mai_mai_n289_), .Y(mai_mai_n313_));
  NA2        m291(.A(mai_mai_n313_), .B(i_3_), .Y(mai_mai_n314_));
  NO2        m292(.A(mai_mai_n86_), .B(mai_mai_n178_), .Y(mai_mai_n315_));
  NA2        m293(.A(mai_mai_n315_), .B(mai_mai_n62_), .Y(mai_mai_n316_));
  NO2        m294(.A(mai_mai_n316_), .B(i_7_), .Y(mai_mai_n317_));
  NO2        m295(.A(mai_mai_n178_), .B(i_9_), .Y(mai_mai_n318_));
  NA2        m296(.A(mai_mai_n318_), .B(mai_mai_n189_), .Y(mai_mai_n319_));
  NO2        m297(.A(mai_mai_n317_), .B(mai_mai_n264_), .Y(mai_mai_n320_));
  AOI210     m298(.A0(mai_mai_n320_), .A1(mai_mai_n314_), .B0(mai_mai_n149_), .Y(mai_mai_n321_));
  AOI210     m299(.A0(mai_mai_n308_), .A1(mai_mai_n284_), .B0(mai_mai_n321_), .Y(mai_mai_n322_));
  NOi32      m300(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n323_));
  INV        m301(.A(mai_mai_n323_), .Y(mai_mai_n324_));
  NAi21      m302(.An(i_0_), .B(i_6_), .Y(mai_mai_n325_));
  NAi21      m303(.An(i_1_), .B(i_5_), .Y(mai_mai_n326_));
  NA2        m304(.A(mai_mai_n326_), .B(mai_mai_n325_), .Y(mai_mai_n327_));
  NA2        m305(.A(mai_mai_n327_), .B(mai_mai_n25_), .Y(mai_mai_n328_));
  OAI210     m306(.A0(mai_mai_n328_), .A1(mai_mai_n146_), .B0(mai_mai_n225_), .Y(mai_mai_n329_));
  NAi41      m307(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n330_));
  OAI220     m308(.A0(mai_mai_n330_), .A1(mai_mai_n326_), .B0(mai_mai_n203_), .B1(mai_mai_n146_), .Y(mai_mai_n331_));
  NO2        m309(.A(mai_mai_n146_), .B(mai_mai_n144_), .Y(mai_mai_n332_));
  OR2        m310(.A(mai_mai_n332_), .B(mai_mai_n331_), .Y(mai_mai_n333_));
  NO2        m311(.A(i_1_), .B(mai_mai_n93_), .Y(mai_mai_n334_));
  NAi21      m312(.An(i_3_), .B(i_4_), .Y(mai_mai_n335_));
  NA2        m313(.A(i_2_), .B(i_7_), .Y(mai_mai_n336_));
  NO2        m314(.A(mai_mai_n335_), .B(i_10_), .Y(mai_mai_n337_));
  AOI210     m315(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n338_));
  OAI210     m316(.A0(mai_mai_n338_), .A1(mai_mai_n173_), .B0(mai_mai_n337_), .Y(mai_mai_n339_));
  AOI220     m317(.A0(mai_mai_n337_), .A1(mai_mai_n305_), .B0(mai_mai_n218_), .B1(mai_mai_n173_), .Y(mai_mai_n340_));
  AOI210     m318(.A0(mai_mai_n340_), .A1(mai_mai_n339_), .B0(i_5_), .Y(mai_mai_n341_));
  NO3        m319(.A(mai_mai_n341_), .B(mai_mai_n333_), .C(mai_mai_n329_), .Y(mai_mai_n342_));
  NO2        m320(.A(mai_mai_n342_), .B(mai_mai_n324_), .Y(mai_mai_n343_));
  NO2        m321(.A(mai_mai_n58_), .B(mai_mai_n25_), .Y(mai_mai_n344_));
  AN2        m322(.A(i_12_), .B(i_5_), .Y(mai_mai_n345_));
  NO2        m323(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n346_));
  NA2        m324(.A(mai_mai_n346_), .B(mai_mai_n345_), .Y(mai_mai_n347_));
  NO2        m325(.A(i_11_), .B(i_6_), .Y(mai_mai_n348_));
  NA3        m326(.A(mai_mai_n348_), .B(i_2_), .C(mai_mai_n204_), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n349_), .B(mai_mai_n347_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n222_), .B(i_5_), .Y(mai_mai_n351_));
  NO2        m329(.A(i_5_), .B(i_10_), .Y(mai_mai_n352_));
  AOI220     m330(.A0(mai_mai_n352_), .A1(mai_mai_n244_), .B0(mai_mai_n351_), .B1(mai_mai_n183_), .Y(mai_mai_n353_));
  NA2        m331(.A(mai_mai_n133_), .B(mai_mai_n45_), .Y(mai_mai_n354_));
  NO2        m332(.A(mai_mai_n354_), .B(mai_mai_n353_), .Y(mai_mai_n355_));
  OAI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n350_), .B0(mai_mai_n344_), .Y(mai_mai_n356_));
  NO2        m334(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n357_));
  NO2        m335(.A(mai_mai_n139_), .B(mai_mai_n80_), .Y(mai_mai_n358_));
  NO2        m336(.A(mai_mai_n358_), .B(mai_mai_n350_), .Y(mai_mai_n359_));
  NO2        m337(.A(i_11_), .B(i_12_), .Y(mai_mai_n360_));
  NA2        m338(.A(mai_mai_n352_), .B(mai_mai_n216_), .Y(mai_mai_n361_));
  NAi21      m339(.An(i_13_), .B(i_0_), .Y(mai_mai_n362_));
  NO2        m340(.A(mai_mai_n362_), .B(mai_mai_n219_), .Y(mai_mai_n363_));
  NA2        m341(.A(mai_mai_n877_), .B(mai_mai_n363_), .Y(mai_mai_n364_));
  NA3        m342(.A(mai_mai_n364_), .B(mai_mai_n359_), .C(mai_mai_n356_), .Y(mai_mai_n365_));
  NA2        m343(.A(mai_mai_n44_), .B(mai_mai_n204_), .Y(mai_mai_n366_));
  NO2        m344(.A(i_0_), .B(i_11_), .Y(mai_mai_n367_));
  AN2        m345(.A(i_1_), .B(i_6_), .Y(mai_mai_n368_));
  NOi21      m346(.An(i_2_), .B(i_12_), .Y(mai_mai_n369_));
  NA2        m347(.A(mai_mai_n369_), .B(mai_mai_n368_), .Y(mai_mai_n370_));
  INV        m348(.A(mai_mai_n370_), .Y(mai_mai_n371_));
  NO2        m349(.A(mai_mai_n881_), .B(i_4_), .Y(mai_mai_n372_));
  NA2        m350(.A(mai_mai_n371_), .B(mai_mai_n372_), .Y(mai_mai_n373_));
  OR2        m351(.A(i_13_), .B(i_10_), .Y(mai_mai_n374_));
  NO3        m352(.A(mai_mai_n374_), .B(mai_mai_n107_), .C(i_9_), .Y(mai_mai_n375_));
  NO2        m353(.A(mai_mai_n159_), .B(mai_mai_n113_), .Y(mai_mai_n376_));
  NO2        m354(.A(mai_mai_n93_), .B(mai_mai_n25_), .Y(mai_mai_n377_));
  NA2        m355(.A(mai_mai_n251_), .B(mai_mai_n194_), .Y(mai_mai_n378_));
  NO2        m356(.A(mai_mai_n378_), .B(mai_mai_n199_), .Y(mai_mai_n379_));
  INV        m357(.A(mai_mai_n379_), .Y(mai_mai_n380_));
  AOI210     m358(.A0(mai_mai_n380_), .A1(mai_mai_n373_), .B0(mai_mai_n26_), .Y(mai_mai_n381_));
  NA2        m359(.A(mai_mai_n291_), .B(mai_mai_n290_), .Y(mai_mai_n382_));
  AOI220     m360(.A0(mai_mai_n267_), .A1(mai_mai_n259_), .B0(mai_mai_n261_), .B1(i_6_), .Y(mai_mai_n383_));
  NO2        m361(.A(mai_mai_n383_), .B(mai_mai_n156_), .Y(mai_mai_n384_));
  NO2        m362(.A(mai_mai_n169_), .B(mai_mai_n80_), .Y(mai_mai_n385_));
  AOI220     m363(.A0(mai_mai_n385_), .A1(mai_mai_n266_), .B0(i_6_), .B1(mai_mai_n194_), .Y(mai_mai_n386_));
  NO2        m364(.A(mai_mai_n386_), .B(i_7_), .Y(mai_mai_n387_));
  NO3        m365(.A(mai_mai_n387_), .B(mai_mai_n384_), .C(mai_mai_n382_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n181_), .B(mai_mai_n88_), .Y(mai_mai_n389_));
  NA3        m367(.A(i_2_), .B(mai_mai_n150_), .C(mai_mai_n80_), .Y(mai_mai_n390_));
  AOI210     m368(.A0(mai_mai_n390_), .A1(mai_mai_n389_), .B0(mai_mai_n292_), .Y(mai_mai_n391_));
  NA2        m369(.A(mai_mai_n267_), .B(mai_mai_n214_), .Y(mai_mai_n392_));
  NO2        m370(.A(mai_mai_n392_), .B(mai_mai_n169_), .Y(mai_mai_n393_));
  NA3        m371(.A(mai_mai_n305_), .B(mai_mai_n304_), .C(i_5_), .Y(mai_mai_n394_));
  INV        m372(.A(mai_mai_n285_), .Y(mai_mai_n395_));
  OAI210     m373(.A0(mai_mai_n395_), .A1(mai_mai_n174_), .B0(mai_mai_n394_), .Y(mai_mai_n396_));
  NO3        m374(.A(mai_mai_n396_), .B(mai_mai_n393_), .C(mai_mai_n391_), .Y(mai_mai_n397_));
  AOI210     m375(.A0(mai_mai_n397_), .A1(mai_mai_n388_), .B0(mai_mai_n246_), .Y(mai_mai_n398_));
  NO4        m376(.A(mai_mai_n398_), .B(mai_mai_n381_), .C(mai_mai_n365_), .D(mai_mai_n343_), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n69_), .B(i_13_), .Y(mai_mai_n400_));
  NA3        m378(.A(mai_mai_n400_), .B(i_1_), .C(i_2_), .Y(mai_mai_n401_));
  NO2        m379(.A(i_10_), .B(i_9_), .Y(mai_mai_n402_));
  NAi21      m380(.An(i_12_), .B(i_8_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n403_), .B(i_3_), .Y(mai_mai_n404_));
  NA2        m382(.A(i_2_), .B(i_6_), .Y(mai_mai_n405_));
  OAI220     m383(.A0(mai_mai_n405_), .A1(mai_mai_n188_), .B0(mai_mai_n880_), .B1(mai_mai_n401_), .Y(mai_mai_n406_));
  NA2        m384(.A(mai_mai_n280_), .B(i_0_), .Y(mai_mai_n407_));
  NO3        m385(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n408_));
  NA2        m386(.A(mai_mai_n241_), .B(mai_mai_n89_), .Y(mai_mai_n409_));
  NA2        m387(.A(mai_mai_n409_), .B(mai_mai_n408_), .Y(mai_mai_n410_));
  NA2        m388(.A(i_8_), .B(i_9_), .Y(mai_mai_n411_));
  NO2        m389(.A(i_7_), .B(i_2_), .Y(mai_mai_n412_));
  OR2        m390(.A(mai_mai_n412_), .B(mai_mai_n411_), .Y(mai_mai_n413_));
  NA2        m391(.A(mai_mai_n257_), .B(mai_mai_n189_), .Y(mai_mai_n414_));
  NO2        m392(.A(mai_mai_n414_), .B(mai_mai_n413_), .Y(mai_mai_n415_));
  NA2        m393(.A(mai_mai_n230_), .B(mai_mai_n279_), .Y(mai_mai_n416_));
  NO3        m394(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n417_));
  INV        m395(.A(mai_mai_n417_), .Y(mai_mai_n418_));
  NA3        m396(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n419_));
  NA3        m397(.A(mai_mai_n134_), .B(mai_mai_n105_), .C(mai_mai_n23_), .Y(mai_mai_n420_));
  OAI220     m398(.A0(mai_mai_n420_), .A1(mai_mai_n419_), .B0(mai_mai_n418_), .B1(mai_mai_n416_), .Y(mai_mai_n421_));
  NO3        m399(.A(mai_mai_n421_), .B(mai_mai_n415_), .C(mai_mai_n406_), .Y(mai_mai_n422_));
  OR2        m400(.A(mai_mai_n265_), .B(mai_mai_n191_), .Y(mai_mai_n423_));
  OA210      m401(.A0(mai_mai_n319_), .A1(mai_mai_n93_), .B0(mai_mai_n268_), .Y(mai_mai_n424_));
  OA220      m402(.A0(mai_mai_n424_), .A1(mai_mai_n149_), .B0(mai_mai_n423_), .B1(mai_mai_n211_), .Y(mai_mai_n425_));
  NA2        m403(.A(mai_mai_n88_), .B(i_13_), .Y(mai_mai_n426_));
  NA2        m404(.A(mai_mai_n385_), .B(mai_mai_n344_), .Y(mai_mai_n427_));
  NO2        m405(.A(i_2_), .B(i_13_), .Y(mai_mai_n428_));
  NO2        m406(.A(mai_mai_n427_), .B(mai_mai_n426_), .Y(mai_mai_n429_));
  NO3        m407(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n430_));
  NO2        m408(.A(i_6_), .B(i_7_), .Y(mai_mai_n431_));
  NA2        m409(.A(mai_mai_n431_), .B(mai_mai_n430_), .Y(mai_mai_n432_));
  NO2        m410(.A(i_11_), .B(i_1_), .Y(mai_mai_n433_));
  NOi21      m411(.An(i_2_), .B(i_7_), .Y(mai_mai_n434_));
  NAi31      m412(.An(i_11_), .B(mai_mai_n434_), .C(i_0_), .Y(mai_mai_n435_));
  NO2        m413(.A(mai_mai_n374_), .B(i_6_), .Y(mai_mai_n436_));
  NA3        m414(.A(mai_mai_n436_), .B(i_1_), .C(mai_mai_n71_), .Y(mai_mai_n437_));
  NO2        m415(.A(mai_mai_n437_), .B(mai_mai_n435_), .Y(mai_mai_n438_));
  NO2        m416(.A(i_3_), .B(mai_mai_n178_), .Y(mai_mai_n439_));
  NO2        m417(.A(i_6_), .B(i_10_), .Y(mai_mai_n440_));
  NA3        m418(.A(mai_mai_n440_), .B(mai_mai_n284_), .C(mai_mai_n439_), .Y(mai_mai_n441_));
  NO2        m419(.A(mai_mai_n441_), .B(mai_mai_n142_), .Y(mai_mai_n442_));
  NA2        m420(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n443_));
  NO2        m421(.A(mai_mai_n144_), .B(i_3_), .Y(mai_mai_n444_));
  NAi31      m422(.An(mai_mai_n443_), .B(mai_mai_n444_), .C(mai_mai_n205_), .Y(mai_mai_n445_));
  NA3        m423(.A(mai_mai_n357_), .B(mai_mai_n165_), .C(mai_mai_n138_), .Y(mai_mai_n446_));
  NA2        m424(.A(mai_mai_n446_), .B(mai_mai_n445_), .Y(mai_mai_n447_));
  NO4        m425(.A(mai_mai_n447_), .B(mai_mai_n442_), .C(mai_mai_n438_), .D(mai_mai_n429_), .Y(mai_mai_n448_));
  NA2        m426(.A(mai_mai_n408_), .B(mai_mai_n345_), .Y(mai_mai_n449_));
  NA2        m427(.A(mai_mai_n417_), .B(mai_mai_n352_), .Y(mai_mai_n450_));
  NAi21      m428(.An(mai_mai_n199_), .B(mai_mai_n360_), .Y(mai_mai_n451_));
  INV        m429(.A(mai_mai_n305_), .Y(mai_mai_n452_));
  NO2        m430(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n453_));
  NA3        m431(.A(i_6_), .B(mai_mai_n453_), .C(mai_mai_n131_), .Y(mai_mai_n454_));
  OR3        m432(.A(mai_mai_n274_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n455_));
  OAI220     m433(.A0(mai_mai_n455_), .A1(mai_mai_n454_), .B0(mai_mai_n452_), .B1(mai_mai_n451_), .Y(mai_mai_n456_));
  NA3        m434(.A(mai_mai_n277_), .B(i_1_), .C(mai_mai_n69_), .Y(mai_mai_n457_));
  NO2        m435(.A(mai_mai_n457_), .B(mai_mai_n432_), .Y(mai_mai_n458_));
  NO2        m436(.A(mai_mai_n458_), .B(mai_mai_n456_), .Y(mai_mai_n459_));
  NA4        m437(.A(mai_mai_n459_), .B(mai_mai_n448_), .C(mai_mai_n425_), .D(mai_mai_n422_), .Y(mai_mai_n460_));
  NA2        m438(.A(mai_mai_n112_), .B(mai_mai_n101_), .Y(mai_mai_n461_));
  AN2        m439(.A(mai_mai_n461_), .B(mai_mai_n408_), .Y(mai_mai_n462_));
  INV        m440(.A(mai_mai_n151_), .Y(mai_mai_n463_));
  OAI210     m441(.A0(mai_mai_n463_), .A1(mai_mai_n211_), .B0(mai_mai_n278_), .Y(mai_mai_n464_));
  AOI220     m442(.A0(mai_mai_n464_), .A1(mai_mai_n293_), .B0(mai_mai_n462_), .B1(mai_mai_n280_), .Y(mai_mai_n465_));
  NA2        m443(.A(mai_mai_n323_), .B(mai_mai_n69_), .Y(mai_mai_n466_));
  NO2        m444(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n467_));
  NAi41      m445(.An(mai_mai_n466_), .B(mai_mai_n440_), .C(mai_mai_n467_), .D(mai_mai_n46_), .Y(mai_mai_n468_));
  AOI210     m446(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n375_), .Y(mai_mai_n469_));
  NA2        m447(.A(mai_mai_n469_), .B(mai_mai_n468_), .Y(mai_mai_n470_));
  INV        m448(.A(mai_mai_n470_), .Y(mai_mai_n471_));
  NA2        m449(.A(mai_mai_n234_), .B(i_1_), .Y(mai_mai_n472_));
  OAI210     m450(.A0(i_8_), .A1(mai_mai_n472_), .B0(mai_mai_n123_), .Y(mai_mai_n473_));
  INV        m451(.A(mai_mai_n184_), .Y(mai_mai_n474_));
  OR2        m452(.A(mai_mai_n169_), .B(i_4_), .Y(mai_mai_n475_));
  INV        m453(.A(mai_mai_n475_), .Y(mai_mai_n476_));
  AOI220     m454(.A0(mai_mai_n476_), .A1(mai_mai_n474_), .B0(mai_mai_n473_), .B1(mai_mai_n376_), .Y(mai_mai_n477_));
  NA3        m455(.A(mai_mai_n477_), .B(mai_mai_n471_), .C(mai_mai_n465_), .Y(mai_mai_n478_));
  NA2        m456(.A(mai_mai_n351_), .B(mai_mai_n266_), .Y(mai_mai_n479_));
  NA2        m457(.A(mai_mai_n347_), .B(mai_mai_n479_), .Y(mai_mai_n480_));
  NO2        m458(.A(mai_mai_n374_), .B(mai_mai_n38_), .Y(mai_mai_n481_));
  NA2        m459(.A(mai_mai_n481_), .B(mai_mai_n480_), .Y(mai_mai_n482_));
  NO2        m460(.A(i_8_), .B(i_7_), .Y(mai_mai_n483_));
  OAI220     m461(.A0(mai_mai_n46_), .A1(mai_mai_n475_), .B0(i_5_), .B1(mai_mai_n222_), .Y(mai_mai_n484_));
  NO2        m462(.A(i_11_), .B(i_6_), .Y(mai_mai_n485_));
  NA3        m463(.A(mai_mai_n485_), .B(mai_mai_n484_), .C(mai_mai_n483_), .Y(mai_mai_n486_));
  AOI220     m464(.A0(mai_mai_n385_), .A1(i_2_), .B0(mai_mai_n226_), .B1(mai_mai_n223_), .Y(mai_mai_n487_));
  OAI220     m465(.A0(mai_mai_n487_), .A1(mai_mai_n237_), .B0(mai_mai_n426_), .B1(mai_mai_n122_), .Y(mai_mai_n488_));
  NA2        m466(.A(mai_mai_n488_), .B(mai_mai_n240_), .Y(mai_mai_n489_));
  NO2        m467(.A(mai_mai_n272_), .B(mai_mai_n167_), .Y(mai_mai_n490_));
  NA2        m468(.A(mai_mai_n161_), .B(mai_mai_n88_), .Y(mai_mai_n491_));
  NO2        m469(.A(mai_mai_n144_), .B(i_5_), .Y(mai_mai_n492_));
  NA3        m470(.A(mai_mai_n492_), .B(mai_mai_n366_), .C(mai_mai_n287_), .Y(mai_mai_n493_));
  NA2        m471(.A(mai_mai_n493_), .B(mai_mai_n491_), .Y(mai_mai_n494_));
  OAI210     m472(.A0(mai_mai_n494_), .A1(mai_mai_n490_), .B0(mai_mai_n417_), .Y(mai_mai_n495_));
  NA4        m473(.A(mai_mai_n495_), .B(mai_mai_n489_), .C(mai_mai_n486_), .D(mai_mai_n482_), .Y(mai_mai_n496_));
  NA2        m474(.A(mai_mai_n257_), .B(mai_mai_n78_), .Y(mai_mai_n497_));
  NO2        m475(.A(mai_mai_n76_), .B(mai_mai_n497_), .Y(mai_mai_n498_));
  NO2        m476(.A(mai_mai_n46_), .B(mai_mai_n160_), .Y(mai_mai_n499_));
  NO2        m477(.A(mai_mai_n499_), .B(mai_mai_n498_), .Y(mai_mai_n500_));
  NO4        m478(.A(mai_mai_n231_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n501_));
  NO3        m479(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n502_));
  NO2        m480(.A(mai_mai_n212_), .B(mai_mai_n36_), .Y(mai_mai_n503_));
  AN2        m481(.A(mai_mai_n503_), .B(mai_mai_n502_), .Y(mai_mai_n504_));
  OA210      m482(.A0(mai_mai_n504_), .A1(mai_mai_n501_), .B0(mai_mai_n323_), .Y(mai_mai_n505_));
  NO2        m483(.A(mai_mai_n374_), .B(i_1_), .Y(mai_mai_n506_));
  NOi31      m484(.An(mai_mai_n506_), .B(mai_mai_n409_), .C(mai_mai_n69_), .Y(mai_mai_n507_));
  AN4        m485(.A(mai_mai_n507_), .B(mai_mai_n372_), .C(mai_mai_n453_), .D(i_2_), .Y(mai_mai_n508_));
  NO2        m486(.A(mai_mai_n383_), .B(mai_mai_n163_), .Y(mai_mai_n509_));
  NO3        m487(.A(mai_mai_n509_), .B(mai_mai_n508_), .C(mai_mai_n505_), .Y(mai_mai_n510_));
  NOi21      m488(.An(i_10_), .B(i_6_), .Y(mai_mai_n511_));
  NA2        m489(.A(mai_mai_n249_), .B(mai_mai_n511_), .Y(mai_mai_n512_));
  NO2        m490(.A(mai_mai_n512_), .B(mai_mai_n407_), .Y(mai_mai_n513_));
  NO2        m491(.A(mai_mai_n104_), .B(mai_mai_n23_), .Y(mai_mai_n514_));
  NA2        m492(.A(mai_mai_n285_), .B(mai_mai_n151_), .Y(mai_mai_n515_));
  AOI220     m493(.A0(mai_mai_n515_), .A1(mai_mai_n392_), .B0(mai_mai_n159_), .B1(mai_mai_n168_), .Y(mai_mai_n516_));
  NO2        m494(.A(mai_mai_n183_), .B(mai_mai_n37_), .Y(mai_mai_n517_));
  NOi31      m495(.An(mai_mai_n135_), .B(mai_mai_n517_), .C(mai_mai_n300_), .Y(mai_mai_n518_));
  NO3        m496(.A(mai_mai_n518_), .B(mai_mai_n516_), .C(mai_mai_n513_), .Y(mai_mai_n519_));
  NO2        m497(.A(mai_mai_n466_), .B(mai_mai_n340_), .Y(mai_mai_n520_));
  INV        m498(.A(mai_mai_n287_), .Y(mai_mai_n521_));
  NO2        m499(.A(i_12_), .B(mai_mai_n80_), .Y(mai_mai_n522_));
  NA3        m500(.A(mai_mai_n522_), .B(mai_mai_n249_), .C(i_5_), .Y(mai_mai_n523_));
  NA3        m501(.A(mai_mai_n348_), .B(mai_mai_n257_), .C(mai_mai_n201_), .Y(mai_mai_n524_));
  AOI210     m502(.A0(mai_mai_n524_), .A1(mai_mai_n523_), .B0(mai_mai_n521_), .Y(mai_mai_n525_));
  NO3        m503(.A(i_4_), .B(mai_mai_n311_), .C(mai_mai_n272_), .Y(mai_mai_n526_));
  NO3        m504(.A(mai_mai_n526_), .B(mai_mai_n525_), .C(mai_mai_n520_), .Y(mai_mai_n527_));
  NA4        m505(.A(mai_mai_n527_), .B(mai_mai_n519_), .C(mai_mai_n510_), .D(mai_mai_n500_), .Y(mai_mai_n528_));
  NO4        m506(.A(mai_mai_n528_), .B(mai_mai_n496_), .C(mai_mai_n478_), .D(mai_mai_n460_), .Y(mai_mai_n529_));
  NA4        m507(.A(mai_mai_n529_), .B(mai_mai_n399_), .C(mai_mai_n322_), .D(mai_mai_n283_), .Y(mai7));
  NO2        m508(.A(mai_mai_n86_), .B(mai_mai_n54_), .Y(mai_mai_n531_));
  NO2        m509(.A(mai_mai_n97_), .B(mai_mai_n85_), .Y(mai_mai_n532_));
  NA2        m510(.A(mai_mai_n440_), .B(mai_mai_n78_), .Y(mai_mai_n533_));
  NA2        m511(.A(i_11_), .B(mai_mai_n178_), .Y(mai_mai_n534_));
  NA3        m512(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n535_));
  NO2        m513(.A(mai_mai_n216_), .B(i_4_), .Y(mai_mai_n536_));
  NO2        m514(.A(mai_mai_n95_), .B(mai_mai_n535_), .Y(mai_mai_n537_));
  NA2        m515(.A(i_2_), .B(mai_mai_n80_), .Y(mai_mai_n538_));
  NO2        m516(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n539_));
  NA2        m517(.A(i_4_), .B(i_8_), .Y(mai_mai_n540_));
  NO4        m518(.A(mai_mai_n187_), .B(mai_mai_n537_), .C(mai_mai_n532_), .D(mai_mai_n531_), .Y(mai_mai_n541_));
  AOI210     m519(.A0(mai_mai_n117_), .A1(mai_mai_n61_), .B0(i_10_), .Y(mai_mai_n542_));
  AOI210     m520(.A0(mai_mai_n542_), .A1(mai_mai_n216_), .B0(mai_mai_n148_), .Y(mai_mai_n543_));
  OR2        m521(.A(i_6_), .B(i_10_), .Y(mai_mai_n544_));
  NO2        m522(.A(mai_mai_n544_), .B(mai_mai_n23_), .Y(mai_mai_n545_));
  NO3        m523(.A(i_10_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n546_));
  NO2        m524(.A(mai_mai_n546_), .B(mai_mai_n545_), .Y(mai_mai_n547_));
  OA220      m525(.A0(mai_mai_n547_), .A1(mai_mai_n521_), .B0(mai_mai_n543_), .B1(mai_mai_n242_), .Y(mai_mai_n548_));
  AOI210     m526(.A0(mai_mai_n548_), .A1(mai_mai_n541_), .B0(mai_mai_n62_), .Y(mai_mai_n549_));
  NOi21      m527(.An(i_11_), .B(i_7_), .Y(mai_mai_n550_));
  NO2        m528(.A(i_2_), .B(mai_mai_n550_), .Y(mai_mai_n551_));
  NA3        m529(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n552_));
  NAi21      m530(.An(mai_mai_n552_), .B(i_11_), .Y(mai_mai_n553_));
  NO2        m531(.A(mai_mai_n553_), .B(mai_mai_n62_), .Y(mai_mai_n554_));
  NA2        m532(.A(mai_mai_n82_), .B(mai_mai_n62_), .Y(mai_mai_n555_));
  AO210      m533(.A0(mai_mai_n555_), .A1(mai_mai_n340_), .B0(mai_mai_n41_), .Y(mai_mai_n556_));
  NA2        m534(.A(mai_mai_n205_), .B(mai_mai_n62_), .Y(mai_mai_n557_));
  NO2        m535(.A(mai_mai_n62_), .B(i_9_), .Y(mai_mai_n558_));
  NO2        m536(.A(i_1_), .B(i_12_), .Y(mai_mai_n559_));
  NA2        m537(.A(mai_mai_n557_), .B(mai_mai_n556_), .Y(mai_mai_n560_));
  OAI210     m538(.A0(mai_mai_n560_), .A1(mai_mai_n554_), .B0(i_6_), .Y(mai_mai_n561_));
  NO2        m539(.A(i_6_), .B(i_11_), .Y(mai_mai_n562_));
  INV        m540(.A(mai_mai_n410_), .Y(mai_mai_n563_));
  NO4        m541(.A(i_12_), .B(mai_mai_n117_), .C(i_13_), .D(mai_mai_n80_), .Y(mai_mai_n564_));
  NA2        m542(.A(mai_mai_n564_), .B(mai_mai_n558_), .Y(mai_mai_n565_));
  INV        m543(.A(mai_mai_n565_), .Y(mai_mai_n566_));
  NA3        m544(.A(mai_mai_n483_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n567_));
  NA2        m545(.A(mai_mai_n127_), .B(i_9_), .Y(mai_mai_n568_));
  NA3        m546(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n569_));
  NO2        m547(.A(mai_mai_n568_), .B(mai_mai_n875_), .Y(mai_mai_n570_));
  NA3        m548(.A(mai_mai_n558_), .B(mai_mai_n287_), .C(i_6_), .Y(mai_mai_n571_));
  NO2        m549(.A(mai_mai_n571_), .B(mai_mai_n23_), .Y(mai_mai_n572_));
  AOI210     m550(.A0(mai_mai_n433_), .A1(mai_mai_n377_), .B0(mai_mai_n221_), .Y(mai_mai_n573_));
  NO2        m551(.A(mai_mai_n573_), .B(mai_mai_n538_), .Y(mai_mai_n574_));
  NO2        m552(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n575_));
  NA2        m553(.A(mai_mai_n575_), .B(mai_mai_n24_), .Y(mai_mai_n576_));
  NO2        m554(.A(mai_mai_n576_), .B(i_6_), .Y(mai_mai_n577_));
  OR4        m555(.A(mai_mai_n577_), .B(mai_mai_n574_), .C(mai_mai_n572_), .D(mai_mai_n570_), .Y(mai_mai_n578_));
  NO3        m556(.A(mai_mai_n578_), .B(mai_mai_n566_), .C(mai_mai_n563_), .Y(mai_mai_n579_));
  NO2        m557(.A(mai_mai_n212_), .B(mai_mai_n44_), .Y(mai_mai_n580_));
  NO3        m558(.A(mai_mai_n580_), .B(mai_mai_n280_), .C(mai_mai_n217_), .Y(mai_mai_n581_));
  NO2        m559(.A(i_10_), .B(i_6_), .Y(mai_mai_n582_));
  NO2        m560(.A(mai_mai_n80_), .B(i_9_), .Y(mai_mai_n583_));
  NO2        m561(.A(mai_mai_n583_), .B(mai_mai_n62_), .Y(mai_mai_n584_));
  NO2        m562(.A(mai_mai_n584_), .B(mai_mai_n559_), .Y(mai_mai_n585_));
  NO4        m563(.A(mai_mai_n585_), .B(mai_mai_n582_), .C(mai_mai_n581_), .D(i_4_), .Y(mai_mai_n586_));
  NA2        m564(.A(i_1_), .B(i_3_), .Y(mai_mai_n587_));
  INV        m565(.A(mai_mai_n586_), .Y(mai_mai_n588_));
  NA3        m566(.A(mai_mai_n588_), .B(mai_mai_n579_), .C(mai_mai_n561_), .Y(mai_mai_n589_));
  NO3        m567(.A(i_11_), .B(i_3_), .C(i_7_), .Y(mai_mai_n590_));
  NOi21      m568(.An(mai_mai_n590_), .B(i_10_), .Y(mai_mai_n591_));
  OA210      m569(.A0(mai_mai_n591_), .A1(mai_mai_n224_), .B0(mai_mai_n80_), .Y(mai_mai_n592_));
  NA3        m570(.A(mai_mai_n440_), .B(mai_mai_n467_), .C(mai_mai_n46_), .Y(mai_mai_n593_));
  NO3        m571(.A(mai_mai_n434_), .B(mai_mai_n540_), .C(mai_mai_n80_), .Y(mai_mai_n594_));
  NA2        m572(.A(mai_mai_n594_), .B(mai_mai_n25_), .Y(mai_mai_n595_));
  NA2        m573(.A(mai_mai_n595_), .B(mai_mai_n593_), .Y(mai_mai_n596_));
  OAI210     m574(.A0(mai_mai_n596_), .A1(mai_mai_n592_), .B0(i_1_), .Y(mai_mai_n597_));
  AOI210     m575(.A0(mai_mai_n241_), .A1(mai_mai_n89_), .B0(i_1_), .Y(mai_mai_n598_));
  NO2        m576(.A(mai_mai_n335_), .B(i_2_), .Y(mai_mai_n599_));
  NA2        m577(.A(mai_mai_n599_), .B(mai_mai_n598_), .Y(mai_mai_n600_));
  AOI210     m578(.A0(mai_mai_n600_), .A1(mai_mai_n597_), .B0(i_13_), .Y(mai_mai_n601_));
  NA2        m579(.A(mai_mai_n96_), .B(mai_mai_n127_), .Y(mai_mai_n602_));
  AOI220     m580(.A0(mai_mai_n428_), .A1(mai_mai_n148_), .B0(i_2_), .B1(mai_mai_n127_), .Y(mai_mai_n603_));
  OAI210     m581(.A0(mai_mai_n603_), .A1(mai_mai_n44_), .B0(mai_mai_n602_), .Y(mai_mai_n604_));
  NO2        m582(.A(mai_mai_n54_), .B(i_12_), .Y(mai_mai_n605_));
  NA2        m583(.A(mai_mai_n224_), .B(mai_mai_n120_), .Y(mai_mai_n606_));
  OAI220     m584(.A0(mai_mai_n606_), .A1(mai_mai_n41_), .B0(mai_mai_n874_), .B1(mai_mai_n86_), .Y(mai_mai_n607_));
  AOI210     m585(.A0(mai_mai_n604_), .A1(mai_mai_n302_), .B0(mai_mai_n607_), .Y(mai_mai_n608_));
  AOI220     m586(.A0(i_7_), .A1(mai_mai_n68_), .B0(mai_mai_n348_), .B1(i_2_), .Y(mai_mai_n609_));
  NO2        m587(.A(mai_mai_n609_), .B(mai_mai_n222_), .Y(mai_mai_n610_));
  AOI210     m588(.A0(mai_mai_n403_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n611_));
  NOi31      m589(.An(mai_mai_n611_), .B(mai_mai_n533_), .C(mai_mai_n44_), .Y(mai_mai_n612_));
  NO3        m590(.A(mai_mai_n67_), .B(mai_mai_n32_), .C(mai_mai_n93_), .Y(mai_mai_n613_));
  NA2        m591(.A(mai_mai_n26_), .B(mai_mai_n178_), .Y(mai_mai_n614_));
  NO3        m592(.A(mai_mai_n434_), .B(mai_mai_n216_), .C(mai_mai_n80_), .Y(mai_mai_n615_));
  AOI210     m593(.A0(mai_mai_n615_), .A1(mai_mai_n26_), .B0(mai_mai_n613_), .Y(mai_mai_n616_));
  NO2        m594(.A(mai_mai_n616_), .B(i_9_), .Y(mai_mai_n617_));
  NO3        m595(.A(mai_mai_n617_), .B(mai_mai_n612_), .C(mai_mai_n610_), .Y(mai_mai_n618_));
  OR2        m596(.A(i_11_), .B(i_6_), .Y(mai_mai_n619_));
  NA3        m597(.A(mai_mai_n536_), .B(mai_mai_n614_), .C(i_7_), .Y(mai_mai_n620_));
  AOI210     m598(.A0(mai_mai_n620_), .A1(mai_mai_n569_), .B0(mai_mai_n619_), .Y(mai_mai_n621_));
  NA3        m599(.A(mai_mai_n369_), .B(mai_mai_n539_), .C(mai_mai_n89_), .Y(mai_mai_n622_));
  NA2        m600(.A(mai_mai_n562_), .B(i_13_), .Y(mai_mai_n623_));
  NA2        m601(.A(i_2_), .B(mai_mai_n614_), .Y(mai_mai_n624_));
  NAi21      m602(.An(i_11_), .B(i_12_), .Y(mai_mai_n625_));
  NOi41      m603(.An(mai_mai_n100_), .B(mai_mai_n625_), .C(i_13_), .D(mai_mai_n80_), .Y(mai_mai_n626_));
  NA2        m604(.A(mai_mai_n626_), .B(mai_mai_n624_), .Y(mai_mai_n627_));
  NA3        m605(.A(mai_mai_n627_), .B(mai_mai_n623_), .C(mai_mai_n622_), .Y(mai_mai_n628_));
  OAI210     m606(.A0(mai_mai_n628_), .A1(mai_mai_n621_), .B0(mai_mai_n62_), .Y(mai_mai_n629_));
  NA2        m607(.A(mai_mai_n216_), .B(mai_mai_n334_), .Y(mai_mai_n630_));
  NO2        m608(.A(mai_mai_n117_), .B(i_2_), .Y(mai_mai_n631_));
  NA2        m609(.A(mai_mai_n631_), .B(mai_mai_n559_), .Y(mai_mai_n632_));
  NA2        m610(.A(mai_mai_n632_), .B(mai_mai_n630_), .Y(mai_mai_n633_));
  NA3        m611(.A(mai_mai_n633_), .B(mai_mai_n45_), .C(mai_mai_n204_), .Y(mai_mai_n634_));
  NA4        m612(.A(mai_mai_n634_), .B(mai_mai_n629_), .C(mai_mai_n618_), .D(mai_mai_n608_), .Y(mai_mai_n635_));
  OR4        m613(.A(mai_mai_n635_), .B(mai_mai_n601_), .C(mai_mai_n589_), .D(mai_mai_n549_), .Y(mai5));
  NO2        m614(.A(i_4_), .B(i_11_), .Y(mai_mai_n637_));
  NA2        m615(.A(mai_mai_n83_), .B(mai_mai_n637_), .Y(mai_mai_n638_));
  INV        m616(.A(mai_mai_n638_), .Y(mai_mai_n639_));
  NO3        m617(.A(i_11_), .B(mai_mai_n216_), .C(i_13_), .Y(mai_mai_n640_));
  NO2        m618(.A(mai_mai_n114_), .B(mai_mai_n23_), .Y(mai_mai_n641_));
  NA2        m619(.A(i_12_), .B(i_8_), .Y(mai_mai_n642_));
  INV        m620(.A(mai_mai_n402_), .Y(mai_mai_n643_));
  NA2        m621(.A(mai_mai_n287_), .B(mai_mai_n514_), .Y(mai_mai_n644_));
  INV        m622(.A(mai_mai_n644_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n645_), .B(mai_mai_n639_), .Y(mai_mai_n646_));
  INV        m624(.A(mai_mai_n158_), .Y(mai_mai_n647_));
  OAI210     m625(.A0(mai_mai_n599_), .A1(mai_mai_n404_), .B0(mai_mai_n100_), .Y(mai_mai_n648_));
  NO2        m626(.A(mai_mai_n648_), .B(mai_mai_n647_), .Y(mai_mai_n649_));
  NO2        m627(.A(mai_mai_n411_), .B(mai_mai_n26_), .Y(mai_mai_n650_));
  INV        m628(.A(mai_mai_n377_), .Y(mai_mai_n651_));
  NA2        m629(.A(mai_mai_n651_), .B(i_2_), .Y(mai_mai_n652_));
  INV        m630(.A(mai_mai_n652_), .Y(mai_mai_n653_));
  INV        m631(.A(mai_mai_n374_), .Y(mai_mai_n654_));
  AOI210     m632(.A0(mai_mai_n654_), .A1(mai_mai_n653_), .B0(mai_mai_n649_), .Y(mai_mai_n655_));
  OAI210     m633(.A0(mai_mai_n884_), .A1(mai_mai_n641_), .B0(i_2_), .Y(mai_mai_n656_));
  NO2        m634(.A(mai_mai_n38_), .B(mai_mai_n26_), .Y(mai_mai_n657_));
  AOI210     m635(.A0(mai_mai_n876_), .A1(mai_mai_n656_), .B0(mai_mai_n178_), .Y(mai_mai_n658_));
  OA210      m636(.A0(mai_mai_n551_), .A1(mai_mai_n116_), .B0(i_13_), .Y(mai_mai_n659_));
  INV        m637(.A(mai_mai_n77_), .Y(mai_mai_n660_));
  NO2        m638(.A(mai_mai_n660_), .B(mai_mai_n336_), .Y(mai_mai_n661_));
  NO2        m639(.A(mai_mai_n137_), .B(mai_mai_n467_), .Y(mai_mai_n662_));
  NA2        m640(.A(mai_mai_n662_), .B(mai_mai_n377_), .Y(mai_mai_n663_));
  NO2        m641(.A(i_2_), .B(mai_mai_n44_), .Y(mai_mai_n664_));
  NA3        m642(.A(mai_mai_n277_), .B(mai_mai_n114_), .C(mai_mai_n42_), .Y(mai_mai_n665_));
  OAI210     m643(.A0(mai_mai_n665_), .A1(mai_mai_n664_), .B0(mai_mai_n663_), .Y(mai_mai_n666_));
  NO4        m644(.A(mai_mai_n666_), .B(mai_mai_n661_), .C(mai_mai_n659_), .D(mai_mai_n658_), .Y(mai_mai_n667_));
  NA2        m645(.A(mai_mai_n514_), .B(mai_mai_n28_), .Y(mai_mai_n668_));
  NA2        m646(.A(mai_mai_n640_), .B(mai_mai_n250_), .Y(mai_mai_n669_));
  NA2        m647(.A(mai_mai_n669_), .B(mai_mai_n668_), .Y(mai_mai_n670_));
  NO2        m648(.A(i_7_), .B(mai_mai_n116_), .Y(mai_mai_n671_));
  NO2        m649(.A(mai_mai_n671_), .B(mai_mai_n534_), .Y(mai_mai_n672_));
  AOI220     m650(.A0(mai_mai_n672_), .A1(mai_mai_n36_), .B0(mai_mai_n670_), .B1(mai_mai_n46_), .Y(mai_mai_n673_));
  NA4        m651(.A(mai_mai_n673_), .B(mai_mai_n667_), .C(mai_mai_n655_), .D(mai_mai_n646_), .Y(mai6));
  NO2        m652(.A(mai_mai_n279_), .B(i_1_), .Y(mai_mai_n675_));
  NO2        m653(.A(mai_mai_n171_), .B(mai_mai_n128_), .Y(mai_mai_n676_));
  OAI210     m654(.A0(mai_mai_n676_), .A1(mai_mai_n675_), .B0(mai_mai_n631_), .Y(mai_mai_n677_));
  NA4        m655(.A(mai_mai_n352_), .B(mai_mai_n439_), .C(mai_mai_n67_), .D(mai_mai_n93_), .Y(mai_mai_n678_));
  INV        m656(.A(mai_mai_n678_), .Y(mai_mai_n679_));
  NO2        m657(.A(mai_mai_n679_), .B(mai_mai_n298_), .Y(mai_mai_n680_));
  AO210      m658(.A0(mai_mai_n680_), .A1(mai_mai_n677_), .B0(i_12_), .Y(mai_mai_n681_));
  NA2        m659(.A(mai_mai_n337_), .B(mai_mai_n305_), .Y(mai_mai_n682_));
  NA2        m660(.A(mai_mai_n522_), .B(mai_mai_n62_), .Y(mai_mai_n683_));
  INV        m661(.A(mai_mai_n591_), .Y(mai_mai_n684_));
  NA3        m662(.A(mai_mai_n684_), .B(mai_mai_n683_), .C(mai_mai_n682_), .Y(mai_mai_n685_));
  NA2        m663(.A(mai_mai_n685_), .B(mai_mai_n69_), .Y(mai_mai_n686_));
  INV        m664(.A(mai_mai_n297_), .Y(mai_mai_n687_));
  NA2        m665(.A(mai_mai_n71_), .B(mai_mai_n120_), .Y(mai_mai_n688_));
  AOI210     m666(.A0(mai_mai_n114_), .A1(mai_mai_n688_), .B0(mai_mai_n687_), .Y(mai_mai_n689_));
  NO2        m667(.A(mai_mai_n231_), .B(i_9_), .Y(mai_mai_n690_));
  NA2        m668(.A(mai_mai_n690_), .B(i_7_), .Y(mai_mai_n691_));
  NO2        m669(.A(mai_mai_n691_), .B(mai_mai_n171_), .Y(mai_mai_n692_));
  NA3        m670(.A(mai_mai_n879_), .B(mai_mai_n431_), .C(mai_mai_n352_), .Y(mai_mai_n693_));
  NAi32      m671(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n694_));
  AOI210     m672(.A0(mai_mai_n619_), .A1(mai_mai_n81_), .B0(mai_mai_n694_), .Y(mai_mai_n695_));
  NA2        m673(.A(mai_mai_n503_), .B(mai_mai_n502_), .Y(mai_mai_n696_));
  NAi31      m674(.An(mai_mai_n695_), .B(mai_mai_n696_), .C(mai_mai_n693_), .Y(mai_mai_n697_));
  OR3        m675(.A(mai_mai_n697_), .B(mai_mai_n692_), .C(mai_mai_n689_), .Y(mai_mai_n698_));
  OR2        m676(.A(mai_mai_n551_), .B(mai_mai_n404_), .Y(mai_mai_n699_));
  NA3        m677(.A(mai_mai_n699_), .B(mai_mai_n136_), .C(mai_mai_n66_), .Y(mai_mai_n700_));
  AO210      m678(.A0(mai_mai_n450_), .A1(mai_mai_n643_), .B0(mai_mai_n36_), .Y(mai_mai_n701_));
  NA2        m679(.A(mai_mai_n701_), .B(mai_mai_n700_), .Y(mai_mai_n702_));
  NA2        m680(.A(mai_mai_n878_), .B(mai_mai_n502_), .Y(mai_mai_n703_));
  INV        m681(.A(mai_mai_n703_), .Y(mai_mai_n704_));
  AO210      m682(.A0(mai_mai_n467_), .A1(mai_mai_n46_), .B0(mai_mai_n82_), .Y(mai_mai_n705_));
  NA2        m683(.A(mai_mai_n705_), .B(mai_mai_n440_), .Y(mai_mai_n706_));
  AOI210     m684(.A0(mai_mai_n404_), .A1(mai_mai_n402_), .B0(mai_mai_n501_), .Y(mai_mai_n707_));
  NA2        m685(.A(mai_mai_n101_), .B(mai_mai_n367_), .Y(mai_mai_n708_));
  NA2        m686(.A(mai_mai_n223_), .B(mai_mai_n46_), .Y(mai_mai_n709_));
  NA3        m687(.A(mai_mai_n708_), .B(mai_mai_n707_), .C(mai_mai_n706_), .Y(mai_mai_n710_));
  NO4        m688(.A(mai_mai_n710_), .B(mai_mai_n704_), .C(mai_mai_n702_), .D(mai_mai_n698_), .Y(mai_mai_n711_));
  NA4        m689(.A(mai_mai_n711_), .B(mai_mai_n686_), .C(mai_mai_n681_), .D(mai_mai_n342_), .Y(mai3));
  NO2        m690(.A(i_11_), .B(mai_mai_n216_), .Y(mai_mai_n713_));
  OAI210     m691(.A0(i_6_), .A1(mai_mai_n261_), .B0(mai_mai_n713_), .Y(mai_mai_n714_));
  NO2        m692(.A(mai_mai_n714_), .B(mai_mai_n178_), .Y(mai_mai_n715_));
  NO2        m693(.A(mai_mai_n407_), .B(mai_mai_n44_), .Y(mai_mai_n716_));
  OA210      m694(.A0(mai_mai_n716_), .A1(mai_mai_n715_), .B0(mai_mai_n161_), .Y(mai_mai_n717_));
  NA2        m695(.A(mai_mai_n369_), .B(mai_mai_n45_), .Y(mai_mai_n718_));
  NO4        m696(.A(mai_mai_n338_), .B(mai_mai_n345_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n719_));
  NA2        m697(.A(mai_mai_n171_), .B(mai_mai_n511_), .Y(mai_mai_n720_));
  NOi21      m698(.An(mai_mai_n720_), .B(mai_mai_n719_), .Y(mai_mai_n721_));
  NA2        m699(.A(mai_mai_n611_), .B(mai_mai_n583_), .Y(mai_mai_n722_));
  NA2        m700(.A(mai_mai_n303_), .B(i_5_), .Y(mai_mai_n723_));
  OAI220     m701(.A0(mai_mai_n723_), .A1(mai_mai_n722_), .B0(mai_mai_n721_), .B1(mai_mai_n62_), .Y(mai_mai_n724_));
  NOi21      m702(.An(i_5_), .B(i_9_), .Y(mai_mai_n725_));
  NA2        m703(.A(mai_mai_n725_), .B(mai_mai_n400_), .Y(mai_mai_n726_));
  NO2        m704(.A(mai_mai_n162_), .B(mai_mai_n137_), .Y(mai_mai_n727_));
  NA2        m705(.A(mai_mai_n727_), .B(mai_mai_n223_), .Y(mai_mai_n728_));
  OAI220     m706(.A0(mai_mai_n728_), .A1(mai_mai_n167_), .B0(i_1_), .B1(mai_mai_n726_), .Y(mai_mai_n729_));
  NO3        m707(.A(mai_mai_n729_), .B(mai_mai_n724_), .C(mai_mai_n717_), .Y(mai_mai_n730_));
  NA2        m708(.A(mai_mai_n171_), .B(mai_mai_n24_), .Y(mai_mai_n731_));
  NO2        m709(.A(mai_mai_n37_), .B(mai_mai_n731_), .Y(mai_mai_n732_));
  NA2        m710(.A(mai_mai_n284_), .B(mai_mai_n118_), .Y(mai_mai_n733_));
  NAi21      m711(.An(mai_mai_n149_), .B(i_5_), .Y(mai_mai_n734_));
  OAI220     m712(.A0(mai_mai_n734_), .A1(mai_mai_n709_), .B0(mai_mai_n733_), .B1(mai_mai_n361_), .Y(mai_mai_n735_));
  NO2        m713(.A(mai_mai_n735_), .B(mai_mai_n732_), .Y(mai_mai_n736_));
  NA2        m714(.A(i_9_), .B(i_0_), .Y(mai_mai_n737_));
  NO3        m715(.A(mai_mai_n737_), .B(mai_mai_n347_), .C(mai_mai_n83_), .Y(mai_mai_n738_));
  INV        m716(.A(mai_mai_n738_), .Y(mai_mai_n739_));
  INV        m717(.A(mai_mai_n431_), .Y(mai_mai_n740_));
  NA2        m718(.A(mai_mai_n640_), .B(mai_mai_n298_), .Y(mai_mai_n741_));
  NO2        m719(.A(mai_mai_n576_), .B(i_5_), .Y(mai_mai_n742_));
  NO2        m720(.A(mai_mai_n233_), .B(mai_mai_n140_), .Y(mai_mai_n743_));
  NA2        m721(.A(i_0_), .B(i_10_), .Y(mai_mai_n744_));
  AN2        m722(.A(mai_mai_n743_), .B(i_6_), .Y(mai_mai_n745_));
  NO2        m723(.A(i_1_), .B(mai_mai_n741_), .Y(mai_mai_n746_));
  NO3        m724(.A(mai_mai_n746_), .B(mai_mai_n745_), .C(mai_mai_n742_), .Y(mai_mai_n747_));
  NA3        m725(.A(mai_mai_n747_), .B(mai_mai_n739_), .C(mai_mai_n736_), .Y(mai_mai_n748_));
  NA2        m726(.A(i_11_), .B(i_9_), .Y(mai_mai_n749_));
  NO2        m727(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n750_));
  NA2        m728(.A(mai_mai_n357_), .B(mai_mai_n165_), .Y(mai_mai_n751_));
  NA2        m729(.A(mai_mai_n751_), .B(mai_mai_n147_), .Y(mai_mai_n752_));
  NO2        m730(.A(mai_mai_n162_), .B(i_0_), .Y(mai_mai_n753_));
  NA2        m731(.A(mai_mai_n431_), .B(mai_mai_n210_), .Y(mai_mai_n754_));
  NO2        m732(.A(mai_mai_n754_), .B(mai_mai_n162_), .Y(mai_mai_n755_));
  NO2        m733(.A(mai_mai_n755_), .B(mai_mai_n752_), .Y(mai_mai_n756_));
  NA2        m734(.A(mai_mai_n575_), .B(mai_mai_n111_), .Y(mai_mai_n757_));
  NO2        m735(.A(i_6_), .B(mai_mai_n757_), .Y(mai_mai_n758_));
  AOI210     m736(.A0(mai_mai_n403_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n759_));
  INV        m737(.A(mai_mai_n94_), .Y(mai_mai_n760_));
  NOi32      m738(.An(mai_mai_n759_), .Bn(mai_mai_n173_), .C(mai_mai_n760_), .Y(mai_mai_n761_));
  NA2        m739(.A(mai_mai_n539_), .B(mai_mai_n298_), .Y(mai_mai_n762_));
  NO2        m740(.A(mai_mai_n762_), .B(mai_mai_n718_), .Y(mai_mai_n763_));
  NO3        m741(.A(mai_mai_n763_), .B(mai_mai_n761_), .C(mai_mai_n758_), .Y(mai_mai_n764_));
  NOi21      m742(.An(i_7_), .B(i_5_), .Y(mai_mai_n765_));
  NOi31      m743(.An(mai_mai_n765_), .B(i_0_), .C(mai_mai_n625_), .Y(mai_mai_n766_));
  NO2        m744(.A(mai_mai_n235_), .B(mai_mai_n288_), .Y(mai_mai_n767_));
  INV        m745(.A(mai_mai_n625_), .Y(mai_mai_n768_));
  NA2        m746(.A(mai_mai_n768_), .B(mai_mai_n767_), .Y(mai_mai_n769_));
  NA3        m747(.A(mai_mai_n769_), .B(mai_mai_n764_), .C(mai_mai_n756_), .Y(mai_mai_n770_));
  NO2        m748(.A(mai_mai_n731_), .B(mai_mai_n219_), .Y(mai_mai_n771_));
  AN2        m749(.A(mai_mai_n302_), .B(mai_mai_n298_), .Y(mai_mai_n772_));
  AN2        m750(.A(mai_mai_n772_), .B(mai_mai_n727_), .Y(mai_mai_n773_));
  OAI210     m751(.A0(mai_mai_n773_), .A1(mai_mai_n771_), .B0(i_10_), .Y(mai_mai_n774_));
  NA3        m752(.A(mai_mai_n430_), .B(mai_mai_n369_), .C(mai_mai_n45_), .Y(mai_mai_n775_));
  OAI210     m753(.A0(mai_mai_n734_), .A1(mai_mai_n740_), .B0(mai_mai_n775_), .Y(mai_mai_n776_));
  NA2        m754(.A(i_0_), .B(mai_mai_n277_), .Y(mai_mai_n777_));
  NA2        m755(.A(mai_mai_n172_), .B(mai_mai_n777_), .Y(mai_mai_n778_));
  AOI220     m756(.A0(mai_mai_n778_), .A1(mai_mai_n431_), .B0(mai_mai_n776_), .B1(mai_mai_n69_), .Y(mai_mai_n779_));
  NO2        m757(.A(mai_mai_n71_), .B(mai_mai_n642_), .Y(mai_mai_n780_));
  AOI210     m758(.A0(mai_mai_n161_), .A1(mai_mai_n532_), .B0(mai_mai_n780_), .Y(mai_mai_n781_));
  NO2        m759(.A(mai_mai_n781_), .B(mai_mai_n47_), .Y(mai_mai_n782_));
  NO3        m760(.A(i_5_), .B(mai_mai_n325_), .C(mai_mai_n24_), .Y(mai_mai_n783_));
  INV        m761(.A(mai_mai_n783_), .Y(mai_mai_n784_));
  NO2        m762(.A(mai_mai_n535_), .B(mai_mai_n95_), .Y(mai_mai_n785_));
  NA2        m763(.A(mai_mai_n785_), .B(i_0_), .Y(mai_mai_n786_));
  OAI220     m764(.A0(mai_mai_n786_), .A1(mai_mai_n80_), .B0(mai_mai_n784_), .B1(mai_mai_n159_), .Y(mai_mai_n787_));
  NO3        m765(.A(mai_mai_n787_), .B(mai_mai_n782_), .C(mai_mai_n470_), .Y(mai_mai_n788_));
  NA3        m766(.A(mai_mai_n788_), .B(mai_mai_n779_), .C(mai_mai_n774_), .Y(mai_mai_n789_));
  NO3        m767(.A(mai_mai_n789_), .B(mai_mai_n770_), .C(mai_mai_n748_), .Y(mai_mai_n790_));
  NO2        m768(.A(i_0_), .B(mai_mai_n625_), .Y(mai_mai_n791_));
  NO2        m769(.A(mai_mai_n683_), .B(mai_mai_n760_), .Y(mai_mai_n792_));
  INV        m770(.A(mai_mai_n792_), .Y(mai_mai_n793_));
  NA3        m771(.A(mai_mai_n135_), .B(mai_mai_n583_), .C(mai_mai_n69_), .Y(mai_mai_n794_));
  NA3        m772(.A(i_6_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n795_));
  NA2        m773(.A(mai_mai_n713_), .B(i_9_), .Y(mai_mai_n796_));
  AOI210     m774(.A0(mai_mai_n795_), .A1(mai_mai_n454_), .B0(mai_mai_n796_), .Y(mai_mai_n797_));
  NA2        m775(.A(mai_mai_n223_), .B(mai_mai_n209_), .Y(mai_mai_n798_));
  AOI210     m776(.A0(mai_mai_n798_), .A1(mai_mai_n737_), .B0(mai_mai_n140_), .Y(mai_mai_n799_));
  NO2        m777(.A(mai_mai_n799_), .B(mai_mai_n797_), .Y(mai_mai_n800_));
  NA3        m778(.A(mai_mai_n800_), .B(mai_mai_n794_), .C(mai_mai_n793_), .Y(mai_mai_n801_));
  NA2        m779(.A(mai_mai_n772_), .B(mai_mai_n336_), .Y(mai_mai_n802_));
  AOI210     m780(.A0(mai_mai_n272_), .A1(mai_mai_n149_), .B0(mai_mai_n802_), .Y(mai_mai_n803_));
  NA2        m781(.A(mai_mai_n750_), .B(mai_mai_n444_), .Y(mai_mai_n804_));
  NO2        m782(.A(mai_mai_n149_), .B(mai_mai_n804_), .Y(mai_mai_n805_));
  NO2        m783(.A(mai_mai_n805_), .B(mai_mai_n803_), .Y(mai_mai_n806_));
  NO2        m784(.A(mai_mai_n744_), .B(mai_mai_n175_), .Y(mai_mai_n807_));
  AOI220     m785(.A0(mai_mai_n807_), .A1(i_11_), .B0(mai_mai_n507_), .B1(mai_mai_n71_), .Y(mai_mai_n808_));
  NO3        m786(.A(mai_mai_n193_), .B(mai_mai_n345_), .C(i_0_), .Y(mai_mai_n809_));
  OAI210     m787(.A0(mai_mai_n809_), .A1(mai_mai_n72_), .B0(i_13_), .Y(mai_mai_n810_));
  INV        m788(.A(mai_mai_n201_), .Y(mai_mai_n811_));
  NO2        m789(.A(i_13_), .B(mai_mai_n128_), .Y(mai_mai_n812_));
  NA3        m790(.A(mai_mai_n812_), .B(i_7_), .C(mai_mai_n811_), .Y(mai_mai_n813_));
  NA4        m791(.A(mai_mai_n813_), .B(mai_mai_n810_), .C(mai_mai_n808_), .D(mai_mai_n806_), .Y(mai_mai_n814_));
  AOI210     m792(.A0(i_6_), .A1(mai_mai_n791_), .B0(mai_mai_n98_), .Y(mai_mai_n815_));
  NA2        m793(.A(mai_mai_n765_), .B(mai_mai_n444_), .Y(mai_mai_n816_));
  OA220      m794(.A0(mai_mai_n162_), .A1(mai_mai_n816_), .B0(mai_mai_n815_), .B1(i_5_), .Y(mai_mai_n817_));
  NO2        m795(.A(i_0_), .B(mai_mai_n162_), .Y(mai_mai_n818_));
  NO3        m796(.A(mai_mai_n718_), .B(mai_mai_n54_), .C(mai_mai_n48_), .Y(mai_mai_n819_));
  INV        m797(.A(mai_mai_n449_), .Y(mai_mai_n820_));
  NO2        m798(.A(mai_mai_n820_), .B(mai_mai_n819_), .Y(mai_mai_n821_));
  NA3        m799(.A(mai_mai_n750_), .B(mai_mai_n261_), .C(mai_mai_n209_), .Y(mai_mai_n822_));
  INV        m800(.A(mai_mai_n822_), .Y(mai_mai_n823_));
  NA3        m801(.A(mai_mai_n352_), .B(mai_mai_n304_), .C(i_4_), .Y(mai_mai_n824_));
  INV        m802(.A(mai_mai_n824_), .Y(mai_mai_n825_));
  NOi31      m803(.An(mai_mai_n351_), .B(i_11_), .C(mai_mai_n219_), .Y(mai_mai_n826_));
  NO3        m804(.A(mai_mai_n749_), .B(mai_mai_n201_), .C(mai_mai_n175_), .Y(mai_mai_n827_));
  NO4        m805(.A(mai_mai_n827_), .B(mai_mai_n826_), .C(mai_mai_n825_), .D(mai_mai_n823_), .Y(mai_mai_n828_));
  NA3        m806(.A(mai_mai_n828_), .B(mai_mai_n821_), .C(mai_mai_n817_), .Y(mai_mai_n829_));
  NA3        m807(.A(mai_mai_n277_), .B(i_5_), .C(mai_mai_n178_), .Y(mai_mai_n830_));
  NA2        m808(.A(mai_mai_n830_), .B(mai_mai_n222_), .Y(mai_mai_n831_));
  NO3        m809(.A(mai_mai_n219_), .B(i_0_), .C(i_12_), .Y(mai_mai_n832_));
  AOI210     m810(.A0(mai_mai_n832_), .A1(mai_mai_n831_), .B0(mai_mai_n679_), .Y(mai_mai_n833_));
  AN2        m811(.A(mai_mai_n744_), .B(mai_mai_n140_), .Y(mai_mai_n834_));
  NO3        m812(.A(mai_mai_n834_), .B(i_12_), .C(mai_mai_n567_), .Y(mai_mai_n835_));
  INV        m813(.A(mai_mai_n835_), .Y(mai_mai_n836_));
  NA3        m814(.A(mai_mai_n90_), .B(mai_mai_n511_), .C(i_11_), .Y(mai_mai_n837_));
  NO2        m815(.A(mai_mai_n837_), .B(mai_mai_n142_), .Y(mai_mai_n838_));
  NA2        m816(.A(mai_mai_n765_), .B(mai_mai_n428_), .Y(mai_mai_n839_));
  OAI220     m817(.A0(i_7_), .A1(mai_mai_n830_), .B0(mai_mai_n839_), .B1(mai_mai_n584_), .Y(mai_mai_n840_));
  AOI210     m818(.A0(mai_mai_n840_), .A1(mai_mai_n753_), .B0(mai_mai_n838_), .Y(mai_mai_n841_));
  NA3        m819(.A(mai_mai_n841_), .B(mai_mai_n836_), .C(mai_mai_n833_), .Y(mai_mai_n842_));
  NO4        m820(.A(mai_mai_n842_), .B(mai_mai_n829_), .C(mai_mai_n814_), .D(mai_mai_n801_), .Y(mai_mai_n843_));
  NA2        m821(.A(mai_mai_n879_), .B(mai_mai_n37_), .Y(mai_mai_n844_));
  NA2        m822(.A(mai_mai_n844_), .B(mai_mai_n543_), .Y(mai_mai_n845_));
  NA2        m823(.A(mai_mai_n845_), .B(mai_mai_n190_), .Y(mai_mai_n846_));
  OR2        m824(.A(i_11_), .B(i_2_), .Y(mai_mai_n847_));
  NO2        m825(.A(mai_mai_n419_), .B(mai_mai_n241_), .Y(mai_mai_n848_));
  AOI210     m826(.A0(mai_mai_n882_), .A1(mai_mai_n48_), .B0(mai_mai_n848_), .Y(mai_mai_n849_));
  AOI210     m827(.A0(mai_mai_n849_), .A1(mai_mai_n846_), .B0(mai_mai_n69_), .Y(mai_mai_n850_));
  NO2        m828(.A(mai_mai_n504_), .B(mai_mai_n341_), .Y(mai_mai_n851_));
  NO2        m829(.A(mai_mai_n851_), .B(mai_mai_n647_), .Y(mai_mai_n852_));
  INV        m830(.A(mai_mai_n72_), .Y(mai_mai_n853_));
  AOI210     m831(.A0(mai_mai_n818_), .A1(mai_mai_n750_), .B0(mai_mai_n766_), .Y(mai_mai_n854_));
  AOI210     m832(.A0(mai_mai_n854_), .A1(mai_mai_n853_), .B0(mai_mai_n587_), .Y(mai_mai_n855_));
  NA2        m833(.A(i_8_), .B(mai_mai_n72_), .Y(mai_mai_n856_));
  NO2        m834(.A(mai_mai_n856_), .B(mai_mai_n216_), .Y(mai_mai_n857_));
  NA2        m835(.A(mai_mai_n88_), .B(mai_mai_n279_), .Y(mai_mai_n858_));
  INV        m836(.A(mai_mai_n858_), .Y(mai_mai_n859_));
  NO3        m837(.A(mai_mai_n859_), .B(mai_mai_n857_), .C(mai_mai_n855_), .Y(mai_mai_n860_));
  OAI210     m838(.A0(mai_mai_n243_), .A1(mai_mai_n145_), .B0(mai_mai_n83_), .Y(mai_mai_n861_));
  NA2        m839(.A(mai_mai_n650_), .B(mai_mai_n261_), .Y(mai_mai_n862_));
  AOI210     m840(.A0(mai_mai_n862_), .A1(mai_mai_n861_), .B0(i_11_), .Y(mai_mai_n863_));
  NO4        m841(.A(i_9_), .B(i_11_), .C(mai_mai_n232_), .D(mai_mai_n231_), .Y(mai_mai_n864_));
  NO2        m842(.A(mai_mai_n864_), .B(mai_mai_n501_), .Y(mai_mai_n865_));
  INV        m843(.A(mai_mai_n331_), .Y(mai_mai_n866_));
  AOI210     m844(.A0(mai_mai_n866_), .A1(mai_mai_n865_), .B0(mai_mai_n41_), .Y(mai_mai_n867_));
  NO2        m845(.A(mai_mai_n867_), .B(mai_mai_n863_), .Y(mai_mai_n868_));
  OAI210     m846(.A0(mai_mai_n860_), .A1(i_4_), .B0(mai_mai_n868_), .Y(mai_mai_n869_));
  NO3        m847(.A(mai_mai_n869_), .B(mai_mai_n852_), .C(mai_mai_n850_), .Y(mai_mai_n870_));
  NA4        m848(.A(mai_mai_n870_), .B(mai_mai_n843_), .C(mai_mai_n790_), .D(mai_mai_n730_), .Y(mai4));
  INV        m849(.A(mai_mai_n605_), .Y(mai_mai_n874_));
  INV        m850(.A(i_2_), .Y(mai_mai_n875_));
  INV        m851(.A(mai_mai_n657_), .Y(mai_mai_n876_));
  INV        m852(.A(mai_mai_n203_), .Y(mai_mai_n877_));
  INV        m853(.A(i_11_), .Y(mai_mai_n878_));
  INV        m854(.A(i_11_), .Y(mai_mai_n879_));
  INV        m855(.A(mai_mai_n402_), .Y(mai_mai_n880_));
  INV        m856(.A(i_7_), .Y(mai_mai_n881_));
  INV        m857(.A(mai_mai_n847_), .Y(mai_mai_n882_));
  INV        m858(.A(i_13_), .Y(mai_mai_n883_));
  INV        m859(.A(mai_mai_n175_), .Y(mai_mai_n884_));
  NAi21      u000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u002(.A(i_9_), .Y(men_men_n25_));
  INV        u003(.A(i_3_), .Y(men_men_n26_));
  NO2        u004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u013(.A(i_4_), .Y(men_men_n36_));
  INV        u014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u020(.A(men_men_n35_), .Y(men1));
  INV        u021(.A(i_11_), .Y(men_men_n44_));
  NO2        u022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u023(.A(i_2_), .Y(men_men_n46_));
  NA2        u024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u025(.A(i_5_), .Y(men_men_n48_));
  NO2        u026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  NA2        u028(.A(i_0_), .B(i_2_), .Y(men_men_n51_));
  NA2        u029(.A(i_7_), .B(i_9_), .Y(men_men_n52_));
  NO2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(i_1_), .B(i_6_), .Y(men_men_n54_));
  NA2        u032(.A(i_8_), .B(i_7_), .Y(men_men_n55_));
  NA2        u033(.A(i_8_), .B(i_12_), .Y(men_men_n56_));
  INV        u034(.A(i_1_), .Y(men_men_n57_));
  NA2        u035(.A(men_men_n57_), .B(i_6_), .Y(men_men_n58_));
  INV        u036(.A(men_men_n31_), .Y(men_men_n59_));
  NA2        u037(.A(men_men_n59_), .B(men_men_n56_), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n50_), .B(i_2_), .Y(men_men_n61_));
  AOI210     u039(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n62_));
  NA2        u040(.A(i_1_), .B(i_6_), .Y(men_men_n63_));
  NO2        u041(.A(men_men_n63_), .B(men_men_n25_), .Y(men_men_n64_));
  INV        u042(.A(i_0_), .Y(men_men_n65_));
  NAi21      u043(.An(i_5_), .B(i_10_), .Y(men_men_n66_));
  NA2        u044(.A(i_5_), .B(i_9_), .Y(men_men_n67_));
  AOI210     u045(.A0(men_men_n67_), .A1(men_men_n66_), .B0(men_men_n65_), .Y(men_men_n68_));
  NO2        u046(.A(men_men_n68_), .B(men_men_n64_), .Y(men_men_n69_));
  NA2        u047(.A(men_men_n61_), .B(men_men_n69_), .Y(men_men_n70_));
  OAI210     u048(.A0(men_men_n70_), .A1(men_men_n60_), .B0(i_0_), .Y(men_men_n71_));
  NA2        u049(.A(i_12_), .B(i_5_), .Y(men_men_n72_));
  NA2        u050(.A(i_2_), .B(i_8_), .Y(men_men_n73_));
  NO2        u051(.A(i_3_), .B(i_9_), .Y(men_men_n74_));
  NO2        u052(.A(i_3_), .B(i_7_), .Y(men_men_n75_));
  NO3        u053(.A(men_men_n75_), .B(men_men_n74_), .C(men_men_n57_), .Y(men_men_n76_));
  INV        u054(.A(i_6_), .Y(men_men_n77_));
  OR4        u055(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n78_));
  INV        u056(.A(men_men_n78_), .Y(men_men_n79_));
  NO2        u057(.A(i_2_), .B(i_7_), .Y(men_men_n80_));
  OAI210     u058(.A0(men_men_n76_), .A1(i_8_), .B0(men_men_n78_), .Y(men_men_n81_));
  NAi21      u059(.An(i_6_), .B(i_10_), .Y(men_men_n82_));
  NA2        u060(.A(i_6_), .B(i_9_), .Y(men_men_n83_));
  AOI210     u061(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n57_), .Y(men_men_n84_));
  NA2        u062(.A(i_2_), .B(i_6_), .Y(men_men_n85_));
  NO3        u063(.A(men_men_n85_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n86_));
  NO2        u064(.A(men_men_n86_), .B(men_men_n84_), .Y(men_men_n87_));
  AOI210     u065(.A0(men_men_n87_), .A1(men_men_n81_), .B0(men_men_n72_), .Y(men_men_n88_));
  AN3        u066(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n89_));
  NAi21      u067(.An(i_6_), .B(i_11_), .Y(men_men_n90_));
  NO2        u068(.A(i_5_), .B(i_8_), .Y(men_men_n91_));
  NOi21      u069(.An(men_men_n91_), .B(men_men_n90_), .Y(men_men_n92_));
  AOI210     u070(.A0(men_men_n89_), .A1(men_men_n32_), .B0(men_men_n92_), .Y(men_men_n93_));
  INV        u071(.A(i_7_), .Y(men_men_n94_));
  NO2        u072(.A(i_0_), .B(i_5_), .Y(men_men_n95_));
  NO2        u073(.A(men_men_n95_), .B(men_men_n77_), .Y(men_men_n96_));
  NA2        u074(.A(i_12_), .B(i_3_), .Y(men_men_n97_));
  INV        u075(.A(men_men_n97_), .Y(men_men_n98_));
  NAi21      u076(.An(i_7_), .B(i_11_), .Y(men_men_n99_));
  NO3        u077(.A(men_men_n99_), .B(men_men_n82_), .C(men_men_n51_), .Y(men_men_n100_));
  AN2        u078(.A(i_2_), .B(i_10_), .Y(men_men_n101_));
  OR2        u079(.A(men_men_n72_), .B(men_men_n54_), .Y(men_men_n102_));
  NO2        u080(.A(i_8_), .B(men_men_n94_), .Y(men_men_n103_));
  NO3        u081(.A(men_men_n103_), .B(men_men_n102_), .C(men_men_n1008_), .Y(men_men_n104_));
  NA2        u082(.A(i_12_), .B(i_7_), .Y(men_men_n105_));
  NA2        u083(.A(i_11_), .B(i_12_), .Y(men_men_n106_));
  INV        u084(.A(men_men_n104_), .Y(men_men_n107_));
  NA3        u085(.A(men_men_n107_), .B(men_men_n97_), .C(men_men_n93_), .Y(men_men_n108_));
  NOi21      u086(.An(i_1_), .B(i_5_), .Y(men_men_n109_));
  NA2        u087(.A(men_men_n109_), .B(i_11_), .Y(men_men_n110_));
  NA2        u088(.A(men_men_n94_), .B(men_men_n37_), .Y(men_men_n111_));
  NA2        u089(.A(i_7_), .B(men_men_n25_), .Y(men_men_n112_));
  NA2        u090(.A(men_men_n112_), .B(men_men_n111_), .Y(men_men_n113_));
  NA2        u091(.A(men_men_n83_), .B(men_men_n82_), .Y(men_men_n114_));
  NAi21      u092(.An(i_3_), .B(i_8_), .Y(men_men_n115_));
  INV        u093(.A(men_men_n115_), .Y(men_men_n116_));
  NOi31      u094(.An(men_men_n116_), .B(men_men_n114_), .C(i_10_), .Y(men_men_n117_));
  NO2        u095(.A(i_1_), .B(men_men_n77_), .Y(men_men_n118_));
  NO2        u096(.A(i_6_), .B(i_5_), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n119_), .B(i_3_), .Y(men_men_n120_));
  AO210      u098(.A0(men_men_n120_), .A1(men_men_n47_), .B0(men_men_n118_), .Y(men_men_n121_));
  OAI220     u099(.A0(men_men_n121_), .A1(men_men_n99_), .B0(men_men_n117_), .B1(men_men_n110_), .Y(men_men_n122_));
  NO3        u100(.A(men_men_n122_), .B(men_men_n108_), .C(men_men_n88_), .Y(men_men_n123_));
  NA2        u101(.A(men_men_n123_), .B(men_men_n71_), .Y(men2));
  NO2        u102(.A(men_men_n57_), .B(men_men_n37_), .Y(men_men_n125_));
  NA3        u103(.A(men_men_n69_), .B(men_men_n61_), .C(men_men_n30_), .Y(men0));
  AN2        u104(.A(i_8_), .B(i_7_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n127_), .B(i_6_), .Y(men_men_n128_));
  NO2        u106(.A(i_12_), .B(i_13_), .Y(men_men_n129_));
  NAi21      u107(.An(i_5_), .B(i_11_), .Y(men_men_n130_));
  NOi21      u108(.An(men_men_n129_), .B(men_men_n130_), .Y(men_men_n131_));
  NO2        u109(.A(i_0_), .B(i_1_), .Y(men_men_n132_));
  NA2        u110(.A(i_2_), .B(i_3_), .Y(men_men_n133_));
  NO2        u111(.A(men_men_n133_), .B(i_4_), .Y(men_men_n134_));
  NA3        u112(.A(men_men_n134_), .B(men_men_n132_), .C(men_men_n131_), .Y(men_men_n135_));
  OR2        u113(.A(men_men_n135_), .B(men_men_n25_), .Y(men_men_n136_));
  AN2        u114(.A(men_men_n129_), .B(men_men_n74_), .Y(men_men_n137_));
  NO2        u115(.A(men_men_n137_), .B(men_men_n27_), .Y(men_men_n138_));
  NA2        u116(.A(i_1_), .B(i_5_), .Y(men_men_n139_));
  NO2        u117(.A(men_men_n65_), .B(men_men_n46_), .Y(men_men_n140_));
  NA2        u118(.A(men_men_n140_), .B(men_men_n36_), .Y(men_men_n141_));
  NO3        u119(.A(men_men_n141_), .B(men_men_n139_), .C(men_men_n138_), .Y(men_men_n142_));
  OR2        u120(.A(i_0_), .B(i_1_), .Y(men_men_n143_));
  NO3        u121(.A(men_men_n143_), .B(men_men_n72_), .C(i_13_), .Y(men_men_n144_));
  NAi32      u122(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n145_));
  NAi21      u123(.An(men_men_n145_), .B(men_men_n144_), .Y(men_men_n146_));
  NOi21      u124(.An(i_4_), .B(i_10_), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n147_), .B(men_men_n39_), .Y(men_men_n148_));
  NO2        u126(.A(i_3_), .B(i_5_), .Y(men_men_n149_));
  NO3        u127(.A(men_men_n65_), .B(i_2_), .C(i_1_), .Y(men_men_n150_));
  NO2        u128(.A(men_men_n1011_), .B(men_men_n142_), .Y(men_men_n151_));
  AOI210     u129(.A0(men_men_n151_), .A1(men_men_n136_), .B0(men_men_n128_), .Y(men_men_n152_));
  NA3        u130(.A(men_men_n65_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n153_));
  NOi21      u131(.An(i_4_), .B(i_9_), .Y(men_men_n154_));
  NOi21      u132(.An(i_11_), .B(i_13_), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  NO2        u134(.A(i_4_), .B(i_5_), .Y(men_men_n157_));
  NAi21      u135(.An(i_12_), .B(i_11_), .Y(men_men_n158_));
  NO2        u136(.A(men_men_n158_), .B(i_13_), .Y(men_men_n159_));
  NA3        u137(.A(men_men_n159_), .B(men_men_n157_), .C(men_men_n74_), .Y(men_men_n160_));
  AOI210     u138(.A0(men_men_n160_), .A1(men_men_n156_), .B0(men_men_n153_), .Y(men_men_n161_));
  NO2        u139(.A(men_men_n65_), .B(men_men_n57_), .Y(men_men_n162_));
  NA2        u140(.A(men_men_n36_), .B(i_5_), .Y(men_men_n163_));
  NAi31      u141(.An(men_men_n163_), .B(men_men_n137_), .C(i_11_), .Y(men_men_n164_));
  NA2        u142(.A(i_3_), .B(i_5_), .Y(men_men_n165_));
  OR2        u143(.A(men_men_n165_), .B(men_men_n156_), .Y(men_men_n166_));
  AOI210     u144(.A0(men_men_n166_), .A1(men_men_n164_), .B0(i_2_), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n65_), .B(i_5_), .Y(men_men_n168_));
  NO2        u146(.A(i_13_), .B(i_10_), .Y(men_men_n169_));
  NA3        u147(.A(men_men_n169_), .B(men_men_n168_), .C(men_men_n44_), .Y(men_men_n170_));
  NO2        u148(.A(i_2_), .B(i_1_), .Y(men_men_n171_));
  NA2        u149(.A(men_men_n171_), .B(i_3_), .Y(men_men_n172_));
  NAi21      u150(.An(i_4_), .B(i_12_), .Y(men_men_n173_));
  NO4        u151(.A(men_men_n173_), .B(men_men_n172_), .C(men_men_n170_), .D(men_men_n25_), .Y(men_men_n174_));
  NO3        u152(.A(men_men_n174_), .B(men_men_n167_), .C(men_men_n161_), .Y(men_men_n175_));
  INV        u153(.A(i_8_), .Y(men_men_n176_));
  NO2        u154(.A(men_men_n176_), .B(i_7_), .Y(men_men_n177_));
  NA2        u155(.A(men_men_n177_), .B(i_6_), .Y(men_men_n178_));
  NO3        u156(.A(i_3_), .B(men_men_n77_), .C(men_men_n48_), .Y(men_men_n179_));
  NA2        u157(.A(men_men_n179_), .B(men_men_n103_), .Y(men_men_n180_));
  NO3        u158(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n181_));
  NA3        u159(.A(men_men_n181_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n182_));
  NO3        u160(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n183_));
  OAI210     u161(.A0(men_men_n89_), .A1(i_12_), .B0(men_men_n183_), .Y(men_men_n184_));
  AOI210     u162(.A0(men_men_n184_), .A1(men_men_n182_), .B0(men_men_n180_), .Y(men_men_n185_));
  NO2        u163(.A(i_3_), .B(i_8_), .Y(men_men_n186_));
  NO3        u164(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n187_));
  NA3        u165(.A(men_men_n187_), .B(men_men_n186_), .C(men_men_n39_), .Y(men_men_n188_));
  NO2        u166(.A(i_13_), .B(i_9_), .Y(men_men_n189_));
  NAi21      u167(.An(i_12_), .B(i_3_), .Y(men_men_n190_));
  NO3        u168(.A(i_0_), .B(i_2_), .C(men_men_n57_), .Y(men_men_n191_));
  NA2        u169(.A(men_men_n191_), .B(i_10_), .Y(men_men_n192_));
  OAI220     u170(.A0(men_men_n192_), .A1(men_men_n190_), .B0(men_men_n95_), .B1(men_men_n188_), .Y(men_men_n193_));
  AOI210     u171(.A0(men_men_n193_), .A1(i_7_), .B0(men_men_n185_), .Y(men_men_n194_));
  OAI220     u172(.A0(men_men_n194_), .A1(i_4_), .B0(men_men_n178_), .B1(men_men_n175_), .Y(men_men_n195_));
  NAi21      u173(.An(i_12_), .B(i_7_), .Y(men_men_n196_));
  NA3        u174(.A(i_13_), .B(men_men_n176_), .C(i_10_), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n197_), .B(men_men_n196_), .Y(men_men_n198_));
  NA2        u176(.A(i_0_), .B(i_5_), .Y(men_men_n199_));
  NA2        u177(.A(men_men_n199_), .B(men_men_n96_), .Y(men_men_n200_));
  OAI220     u178(.A0(men_men_n200_), .A1(men_men_n172_), .B0(i_2_), .B1(men_men_n120_), .Y(men_men_n201_));
  NAi31      u179(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n36_), .B(i_13_), .Y(men_men_n203_));
  NO2        u181(.A(men_men_n46_), .B(men_men_n57_), .Y(men_men_n204_));
  NA3        u182(.A(men_men_n204_), .B(i_3_), .C(men_men_n203_), .Y(men_men_n205_));
  INV        u183(.A(i_13_), .Y(men_men_n206_));
  NO2        u184(.A(i_12_), .B(men_men_n206_), .Y(men_men_n207_));
  NA3        u185(.A(men_men_n207_), .B(men_men_n181_), .C(men_men_n179_), .Y(men_men_n208_));
  OAI210     u186(.A0(men_men_n205_), .A1(men_men_n202_), .B0(men_men_n208_), .Y(men_men_n209_));
  AOI220     u187(.A0(men_men_n209_), .A1(men_men_n127_), .B0(men_men_n201_), .B1(men_men_n198_), .Y(men_men_n210_));
  NO2        u188(.A(i_12_), .B(men_men_n37_), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n165_), .B(i_4_), .Y(men_men_n212_));
  NA2        u190(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n213_));
  OR2        u191(.A(i_8_), .B(i_7_), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n214_), .B(men_men_n77_), .Y(men_men_n215_));
  NO2        u193(.A(men_men_n51_), .B(i_1_), .Y(men_men_n216_));
  NA2        u194(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  INV        u195(.A(i_12_), .Y(men_men_n218_));
  NO3        u196(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n219_));
  NA2        u197(.A(i_2_), .B(i_1_), .Y(men_men_n220_));
  NO2        u198(.A(men_men_n217_), .B(men_men_n213_), .Y(men_men_n221_));
  NO3        u199(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n222_));
  NAi21      u200(.An(i_4_), .B(i_3_), .Y(men_men_n223_));
  NO2        u201(.A(men_men_n223_), .B(men_men_n67_), .Y(men_men_n224_));
  NO2        u202(.A(i_0_), .B(i_6_), .Y(men_men_n225_));
  NOi41      u203(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n226_));
  NA2        u204(.A(men_men_n226_), .B(men_men_n225_), .Y(men_men_n227_));
  NA2        u205(.A(men_men_n221_), .B(men_men_n189_), .Y(men_men_n228_));
  NO2        u206(.A(i_11_), .B(men_men_n206_), .Y(men_men_n229_));
  NOi21      u207(.An(i_1_), .B(i_6_), .Y(men_men_n230_));
  NAi21      u208(.An(i_3_), .B(i_7_), .Y(men_men_n231_));
  NA2        u209(.A(men_men_n218_), .B(i_9_), .Y(men_men_n232_));
  OR4        u210(.A(men_men_n232_), .B(men_men_n231_), .C(men_men_n230_), .D(men_men_n168_), .Y(men_men_n233_));
  NO2        u211(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n234_));
  NO2        u212(.A(i_12_), .B(i_3_), .Y(men_men_n235_));
  NA2        u213(.A(i_3_), .B(i_9_), .Y(men_men_n236_));
  NAi21      u214(.An(i_7_), .B(i_10_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  NA3        u216(.A(men_men_n238_), .B(men_men_n1010_), .C(men_men_n58_), .Y(men_men_n239_));
  NA2        u217(.A(men_men_n239_), .B(men_men_n233_), .Y(men_men_n240_));
  NA3        u218(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n241_));
  NA2        u219(.A(men_men_n218_), .B(i_13_), .Y(men_men_n242_));
  NO2        u220(.A(men_men_n242_), .B(men_men_n67_), .Y(men_men_n243_));
  AOI220     u221(.A0(men_men_n243_), .A1(men_men_n127_), .B0(men_men_n240_), .B1(men_men_n229_), .Y(men_men_n244_));
  NO2        u222(.A(men_men_n214_), .B(men_men_n37_), .Y(men_men_n245_));
  NA2        u223(.A(i_12_), .B(i_6_), .Y(men_men_n246_));
  NO3        u224(.A(i_9_), .B(men_men_n246_), .C(men_men_n48_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n223_), .B(i_2_), .Y(men_men_n248_));
  NA3        u226(.A(men_men_n248_), .B(men_men_n247_), .C(men_men_n44_), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n229_), .B(i_9_), .Y(men_men_n250_));
  OAI210     u228(.A0(men_men_n65_), .A1(men_men_n250_), .B0(men_men_n249_), .Y(men_men_n251_));
  NO3        u229(.A(i_11_), .B(men_men_n206_), .C(men_men_n25_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n231_), .B(i_8_), .Y(men_men_n253_));
  NO2        u231(.A(i_6_), .B(men_men_n48_), .Y(men_men_n254_));
  NA3        u232(.A(men_men_n254_), .B(men_men_n253_), .C(men_men_n252_), .Y(men_men_n255_));
  NO3        u233(.A(men_men_n26_), .B(men_men_n77_), .C(i_5_), .Y(men_men_n256_));
  NA3        u234(.A(men_men_n256_), .B(men_men_n245_), .C(men_men_n207_), .Y(men_men_n257_));
  AOI210     u235(.A0(men_men_n257_), .A1(men_men_n255_), .B0(men_men_n46_), .Y(men_men_n258_));
  AOI210     u236(.A0(men_men_n251_), .A1(men_men_n245_), .B0(men_men_n258_), .Y(men_men_n259_));
  NA4        u237(.A(men_men_n259_), .B(men_men_n244_), .C(men_men_n228_), .D(men_men_n210_), .Y(men_men_n260_));
  NO3        u238(.A(i_12_), .B(men_men_n206_), .C(men_men_n37_), .Y(men_men_n261_));
  INV        u239(.A(men_men_n261_), .Y(men_men_n262_));
  INV        u240(.A(i_8_), .Y(men_men_n263_));
  NOi21      u241(.An(men_men_n149_), .B(men_men_n77_), .Y(men_men_n264_));
  NO3        u242(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n265_));
  AOI220     u243(.A0(men_men_n265_), .A1(men_men_n179_), .B0(men_men_n264_), .B1(men_men_n216_), .Y(men_men_n266_));
  NO2        u244(.A(men_men_n266_), .B(men_men_n263_), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n220_), .B(i_0_), .Y(men_men_n268_));
  AOI220     u246(.A0(men_men_n268_), .A1(men_men_n177_), .B0(i_1_), .B1(men_men_n127_), .Y(men_men_n269_));
  NA2        u247(.A(men_men_n254_), .B(men_men_n26_), .Y(men_men_n270_));
  NO2        u248(.A(men_men_n270_), .B(men_men_n269_), .Y(men_men_n271_));
  NA2        u249(.A(i_0_), .B(i_1_), .Y(men_men_n272_));
  NO2        u250(.A(men_men_n272_), .B(i_2_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n55_), .B(i_6_), .Y(men_men_n274_));
  NA3        u252(.A(men_men_n274_), .B(men_men_n273_), .C(men_men_n149_), .Y(men_men_n275_));
  OAI210     u253(.A0(i_3_), .A1(men_men_n128_), .B0(men_men_n275_), .Y(men_men_n276_));
  NO3        u254(.A(men_men_n276_), .B(men_men_n271_), .C(men_men_n267_), .Y(men_men_n277_));
  NO2        u255(.A(i_3_), .B(i_10_), .Y(men_men_n278_));
  NA3        u256(.A(men_men_n278_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n279_));
  NO2        u257(.A(i_2_), .B(men_men_n94_), .Y(men_men_n280_));
  NA2        u258(.A(i_1_), .B(men_men_n36_), .Y(men_men_n281_));
  NOi21      u259(.An(men_men_n199_), .B(men_men_n95_), .Y(men_men_n282_));
  NA3        u260(.A(men_men_n282_), .B(i_1_), .C(men_men_n280_), .Y(men_men_n283_));
  AN2        u261(.A(i_3_), .B(i_10_), .Y(men_men_n284_));
  NA4        u262(.A(men_men_n284_), .B(men_men_n181_), .C(men_men_n159_), .D(men_men_n157_), .Y(men_men_n285_));
  NO2        u263(.A(i_5_), .B(men_men_n37_), .Y(men_men_n286_));
  NO2        u264(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n287_));
  OR2        u265(.A(men_men_n283_), .B(men_men_n279_), .Y(men_men_n288_));
  OAI220     u266(.A0(men_men_n288_), .A1(i_6_), .B0(men_men_n277_), .B1(men_men_n262_), .Y(men_men_n289_));
  NO4        u267(.A(men_men_n289_), .B(men_men_n260_), .C(men_men_n195_), .D(men_men_n152_), .Y(men_men_n290_));
  NO3        u268(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n291_));
  NO2        u269(.A(men_men_n55_), .B(men_men_n77_), .Y(men_men_n292_));
  NA2        u270(.A(men_men_n268_), .B(men_men_n292_), .Y(men_men_n293_));
  NO3        u271(.A(i_6_), .B(men_men_n176_), .C(i_7_), .Y(men_men_n294_));
  NA2        u272(.A(men_men_n294_), .B(men_men_n181_), .Y(men_men_n295_));
  AOI210     u273(.A0(men_men_n295_), .A1(men_men_n293_), .B0(i_5_), .Y(men_men_n296_));
  NO2        u274(.A(i_2_), .B(i_3_), .Y(men_men_n297_));
  OR2        u275(.A(i_0_), .B(i_5_), .Y(men_men_n298_));
  NA2        u276(.A(men_men_n199_), .B(men_men_n298_), .Y(men_men_n299_));
  NA4        u277(.A(men_men_n299_), .B(men_men_n215_), .C(men_men_n297_), .D(i_1_), .Y(men_men_n300_));
  NA3        u278(.A(men_men_n268_), .B(men_men_n264_), .C(men_men_n103_), .Y(men_men_n301_));
  NO2        u279(.A(men_men_n143_), .B(men_men_n46_), .Y(men_men_n302_));
  NA3        u280(.A(men_men_n302_), .B(i_7_), .C(men_men_n149_), .Y(men_men_n303_));
  NA3        u281(.A(men_men_n303_), .B(men_men_n301_), .C(men_men_n300_), .Y(men_men_n304_));
  OAI210     u282(.A0(men_men_n304_), .A1(men_men_n296_), .B0(i_4_), .Y(men_men_n305_));
  NO2        u283(.A(i_12_), .B(i_10_), .Y(men_men_n306_));
  NOi21      u284(.An(i_5_), .B(i_0_), .Y(men_men_n307_));
  AOI210     u285(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n94_), .Y(men_men_n308_));
  NO3        u286(.A(men_men_n308_), .B(men_men_n281_), .C(men_men_n115_), .Y(men_men_n309_));
  NA4        u287(.A(men_men_n75_), .B(men_men_n36_), .C(men_men_n77_), .D(i_8_), .Y(men_men_n310_));
  NA2        u288(.A(men_men_n309_), .B(men_men_n306_), .Y(men_men_n311_));
  NO2        u289(.A(i_6_), .B(i_8_), .Y(men_men_n312_));
  NOi21      u290(.An(i_0_), .B(i_2_), .Y(men_men_n313_));
  AN2        u291(.A(men_men_n313_), .B(men_men_n312_), .Y(men_men_n314_));
  NO2        u292(.A(i_1_), .B(i_7_), .Y(men_men_n315_));
  NA3        u293(.A(men_men_n312_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n316_));
  NA3        u294(.A(men_men_n316_), .B(men_men_n311_), .C(men_men_n305_), .Y(men_men_n317_));
  INV        u295(.A(i_8_), .Y(men_men_n318_));
  NOi21      u296(.An(men_men_n139_), .B(men_men_n96_), .Y(men_men_n319_));
  NA2        u297(.A(men_men_n318_), .B(i_3_), .Y(men_men_n320_));
  NO2        u298(.A(men_men_n272_), .B(men_men_n73_), .Y(men_men_n321_));
  NA2        u299(.A(men_men_n321_), .B(men_men_n119_), .Y(men_men_n322_));
  NO2        u300(.A(men_men_n85_), .B(men_men_n176_), .Y(men_men_n323_));
  NA3        u301(.A(men_men_n282_), .B(men_men_n323_), .C(men_men_n57_), .Y(men_men_n324_));
  AOI210     u302(.A0(men_men_n324_), .A1(men_men_n322_), .B0(i_3_), .Y(men_men_n325_));
  NO2        u303(.A(men_men_n176_), .B(i_9_), .Y(men_men_n326_));
  NA2        u304(.A(men_men_n326_), .B(i_1_), .Y(men_men_n327_));
  NO2        u305(.A(men_men_n325_), .B(men_men_n271_), .Y(men_men_n328_));
  AOI210     u306(.A0(men_men_n328_), .A1(men_men_n320_), .B0(men_men_n148_), .Y(men_men_n329_));
  AOI210     u307(.A0(men_men_n317_), .A1(men_men_n291_), .B0(men_men_n329_), .Y(men_men_n330_));
  NOi32      u308(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n331_));
  INV        u309(.A(men_men_n331_), .Y(men_men_n332_));
  NAi21      u310(.An(i_1_), .B(i_5_), .Y(men_men_n333_));
  NA2        u311(.A(men_men_n333_), .B(i_0_), .Y(men_men_n334_));
  NA2        u312(.A(men_men_n334_), .B(men_men_n25_), .Y(men_men_n335_));
  OAI210     u313(.A0(men_men_n335_), .A1(men_men_n145_), .B0(men_men_n227_), .Y(men_men_n336_));
  NAi41      u314(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n337_));
  OAI220     u315(.A0(men_men_n337_), .A1(men_men_n333_), .B0(men_men_n202_), .B1(men_men_n145_), .Y(men_men_n338_));
  AOI210     u316(.A0(men_men_n337_), .A1(men_men_n145_), .B0(men_men_n143_), .Y(men_men_n339_));
  NOi32      u317(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n340_));
  NA2        u318(.A(men_men_n340_), .B(men_men_n46_), .Y(men_men_n341_));
  NO2        u319(.A(men_men_n341_), .B(i_0_), .Y(men_men_n342_));
  OR3        u320(.A(men_men_n342_), .B(men_men_n339_), .C(men_men_n338_), .Y(men_men_n343_));
  NO2        u321(.A(i_1_), .B(men_men_n94_), .Y(men_men_n344_));
  NAi21      u322(.An(i_3_), .B(i_4_), .Y(men_men_n345_));
  NO2        u323(.A(men_men_n345_), .B(i_9_), .Y(men_men_n346_));
  AN2        u324(.A(i_6_), .B(i_7_), .Y(men_men_n347_));
  OAI210     u325(.A0(men_men_n347_), .A1(men_men_n344_), .B0(men_men_n346_), .Y(men_men_n348_));
  NA2        u326(.A(i_2_), .B(i_7_), .Y(men_men_n349_));
  NO2        u327(.A(men_men_n345_), .B(i_10_), .Y(men_men_n350_));
  NA3        u328(.A(men_men_n350_), .B(men_men_n349_), .C(men_men_n225_), .Y(men_men_n351_));
  AOI210     u329(.A0(men_men_n351_), .A1(men_men_n348_), .B0(men_men_n168_), .Y(men_men_n352_));
  AOI220     u330(.A0(men_men_n350_), .A1(men_men_n315_), .B0(men_men_n219_), .B1(men_men_n171_), .Y(men_men_n353_));
  NO3        u331(.A(men_men_n352_), .B(men_men_n343_), .C(men_men_n336_), .Y(men_men_n354_));
  NO2        u332(.A(men_men_n354_), .B(men_men_n332_), .Y(men_men_n355_));
  NO2        u333(.A(men_men_n55_), .B(men_men_n25_), .Y(men_men_n356_));
  AN2        u334(.A(i_12_), .B(i_5_), .Y(men_men_n357_));
  NO2        u335(.A(i_4_), .B(men_men_n26_), .Y(men_men_n358_));
  NO2        u336(.A(i_11_), .B(i_6_), .Y(men_men_n359_));
  NA3        u337(.A(men_men_n359_), .B(men_men_n302_), .C(men_men_n206_), .Y(men_men_n360_));
  NO2        u338(.A(men_men_n360_), .B(men_men_n1007_), .Y(men_men_n361_));
  NO2        u339(.A(men_men_n223_), .B(i_5_), .Y(men_men_n362_));
  NO2        u340(.A(i_5_), .B(i_10_), .Y(men_men_n363_));
  NA2        u341(.A(men_men_n129_), .B(men_men_n45_), .Y(men_men_n364_));
  NO2        u342(.A(men_men_n364_), .B(men_men_n223_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n365_), .A1(men_men_n361_), .B0(men_men_n356_), .Y(men_men_n366_));
  NO2        u344(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n367_));
  INV        u345(.A(men_men_n135_), .Y(men_men_n368_));
  OAI210     u346(.A0(men_men_n368_), .A1(men_men_n361_), .B0(men_men_n367_), .Y(men_men_n369_));
  NO3        u347(.A(men_men_n77_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n370_));
  NO2        u348(.A(i_3_), .B(men_men_n94_), .Y(men_men_n371_));
  NO2        u349(.A(i_11_), .B(i_12_), .Y(men_men_n372_));
  NA2        u350(.A(men_men_n363_), .B(men_men_n218_), .Y(men_men_n373_));
  NA3        u351(.A(men_men_n103_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n374_));
  OAI220     u352(.A0(men_men_n374_), .A1(men_men_n202_), .B0(men_men_n373_), .B1(men_men_n310_), .Y(men_men_n375_));
  NAi21      u353(.An(i_13_), .B(i_0_), .Y(men_men_n376_));
  INV        u354(.A(men_men_n375_), .Y(men_men_n377_));
  NA3        u355(.A(men_men_n377_), .B(men_men_n369_), .C(men_men_n366_), .Y(men_men_n378_));
  NO3        u356(.A(i_1_), .B(i_12_), .C(men_men_n77_), .Y(men_men_n379_));
  NO2        u357(.A(i_0_), .B(i_11_), .Y(men_men_n380_));
  INV        u358(.A(i_5_), .Y(men_men_n381_));
  NOi21      u359(.An(i_2_), .B(i_12_), .Y(men_men_n382_));
  NO2        u360(.A(i_12_), .B(men_men_n381_), .Y(men_men_n383_));
  NA2        u361(.A(men_men_n127_), .B(i_9_), .Y(men_men_n384_));
  NO2        u362(.A(men_men_n384_), .B(i_4_), .Y(men_men_n385_));
  NA2        u363(.A(men_men_n383_), .B(men_men_n385_), .Y(men_men_n386_));
  NAi21      u364(.An(i_9_), .B(i_4_), .Y(men_men_n387_));
  OR2        u365(.A(i_13_), .B(i_10_), .Y(men_men_n388_));
  NO2        u366(.A(men_men_n156_), .B(men_men_n111_), .Y(men_men_n389_));
  NO2        u367(.A(men_men_n94_), .B(men_men_n25_), .Y(men_men_n390_));
  NA2        u368(.A(men_men_n261_), .B(men_men_n390_), .Y(men_men_n391_));
  INV        u369(.A(men_men_n191_), .Y(men_men_n392_));
  OAI220     u370(.A0(men_men_n392_), .A1(men_men_n196_), .B0(men_men_n391_), .B1(men_men_n319_), .Y(men_men_n393_));
  INV        u371(.A(men_men_n393_), .Y(men_men_n394_));
  AOI210     u372(.A0(men_men_n394_), .A1(men_men_n386_), .B0(men_men_n26_), .Y(men_men_n395_));
  NA2        u373(.A(men_men_n301_), .B(men_men_n300_), .Y(men_men_n396_));
  AOI220     u374(.A0(men_men_n274_), .A1(men_men_n265_), .B0(men_men_n268_), .B1(men_men_n292_), .Y(men_men_n397_));
  NO2        u375(.A(men_men_n165_), .B(men_men_n77_), .Y(men_men_n398_));
  AOI220     u376(.A0(men_men_n398_), .A1(men_men_n273_), .B0(men_men_n256_), .B1(men_men_n191_), .Y(men_men_n399_));
  NO2        u377(.A(men_men_n399_), .B(men_men_n263_), .Y(men_men_n400_));
  NO2        u378(.A(men_men_n400_), .B(men_men_n396_), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n179_), .B(men_men_n89_), .Y(men_men_n402_));
  NA3        u380(.A(men_men_n302_), .B(men_men_n149_), .C(men_men_n77_), .Y(men_men_n403_));
  AOI210     u381(.A0(men_men_n403_), .A1(men_men_n402_), .B0(i_8_), .Y(men_men_n404_));
  NA3        u382(.A(men_men_n1010_), .B(men_men_n58_), .C(i_2_), .Y(men_men_n405_));
  NA2        u383(.A(men_men_n274_), .B(men_men_n216_), .Y(men_men_n406_));
  OAI220     u384(.A0(men_men_n406_), .A1(men_men_n165_), .B0(men_men_n405_), .B1(men_men_n1004_), .Y(men_men_n407_));
  NO2        u385(.A(i_3_), .B(men_men_n48_), .Y(men_men_n408_));
  NA3        u386(.A(men_men_n315_), .B(men_men_n314_), .C(men_men_n408_), .Y(men_men_n409_));
  NA2        u387(.A(men_men_n294_), .B(men_men_n299_), .Y(men_men_n410_));
  NA2        u388(.A(men_men_n410_), .B(men_men_n409_), .Y(men_men_n411_));
  NO3        u389(.A(men_men_n411_), .B(men_men_n407_), .C(men_men_n404_), .Y(men_men_n412_));
  AOI210     u390(.A0(men_men_n412_), .A1(men_men_n401_), .B0(men_men_n250_), .Y(men_men_n413_));
  NO4        u391(.A(men_men_n413_), .B(men_men_n395_), .C(men_men_n378_), .D(men_men_n355_), .Y(men_men_n414_));
  NO2        u392(.A(men_men_n57_), .B(i_4_), .Y(men_men_n415_));
  NO2        u393(.A(men_men_n65_), .B(i_13_), .Y(men_men_n416_));
  NA3        u394(.A(men_men_n416_), .B(men_men_n415_), .C(i_2_), .Y(men_men_n417_));
  NO2        u395(.A(i_10_), .B(i_9_), .Y(men_men_n418_));
  NAi21      u396(.An(i_12_), .B(i_8_), .Y(men_men_n419_));
  NO2        u397(.A(men_men_n419_), .B(i_3_), .Y(men_men_n420_));
  NA2        u398(.A(men_men_n420_), .B(men_men_n418_), .Y(men_men_n421_));
  NA2        u399(.A(men_men_n1002_), .B(men_men_n96_), .Y(men_men_n422_));
  OAI220     u400(.A0(men_men_n422_), .A1(men_men_n188_), .B0(men_men_n421_), .B1(men_men_n417_), .Y(men_men_n423_));
  NA2        u401(.A(men_men_n287_), .B(i_0_), .Y(men_men_n424_));
  NO3        u402(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n425_));
  NA2        u403(.A(men_men_n246_), .B(men_men_n90_), .Y(men_men_n426_));
  NA2        u404(.A(men_men_n426_), .B(men_men_n425_), .Y(men_men_n427_));
  NA2        u405(.A(i_8_), .B(i_9_), .Y(men_men_n428_));
  NO2        u406(.A(men_men_n427_), .B(men_men_n424_), .Y(men_men_n429_));
  NA2        u407(.A(men_men_n229_), .B(men_men_n286_), .Y(men_men_n430_));
  NO3        u408(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n431_));
  AOI210     u409(.A0(men_men_n235_), .A1(men_men_n171_), .B0(men_men_n431_), .Y(men_men_n432_));
  NO2        u410(.A(men_men_n432_), .B(men_men_n430_), .Y(men_men_n433_));
  NO3        u411(.A(men_men_n433_), .B(men_men_n429_), .C(men_men_n423_), .Y(men_men_n434_));
  NA2        u412(.A(men_men_n273_), .B(men_men_n99_), .Y(men_men_n435_));
  OA220      u413(.A0(men_men_n327_), .A1(men_men_n148_), .B0(men_men_n435_), .B1(men_men_n213_), .Y(men_men_n436_));
  NA2        u414(.A(men_men_n89_), .B(i_13_), .Y(men_men_n437_));
  NA2        u415(.A(men_men_n398_), .B(men_men_n356_), .Y(men_men_n438_));
  NO2        u416(.A(i_2_), .B(i_13_), .Y(men_men_n439_));
  NA3        u417(.A(men_men_n439_), .B(men_men_n147_), .C(men_men_n92_), .Y(men_men_n440_));
  NO2        u418(.A(men_men_n438_), .B(men_men_n437_), .Y(men_men_n441_));
  NO3        u419(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n442_));
  NO2        u420(.A(i_6_), .B(i_7_), .Y(men_men_n443_));
  NA2        u421(.A(men_men_n443_), .B(men_men_n442_), .Y(men_men_n444_));
  OR2        u422(.A(i_11_), .B(i_8_), .Y(men_men_n445_));
  NOi21      u423(.An(i_2_), .B(i_7_), .Y(men_men_n446_));
  NAi31      u424(.An(men_men_n445_), .B(men_men_n446_), .C(men_men_n999_), .Y(men_men_n447_));
  NO2        u425(.A(men_men_n388_), .B(i_6_), .Y(men_men_n448_));
  NA3        u426(.A(men_men_n448_), .B(men_men_n415_), .C(men_men_n67_), .Y(men_men_n449_));
  NO2        u427(.A(men_men_n449_), .B(men_men_n447_), .Y(men_men_n450_));
  NO2        u428(.A(i_3_), .B(men_men_n176_), .Y(men_men_n451_));
  NO2        u429(.A(i_6_), .B(i_10_), .Y(men_men_n452_));
  NA4        u430(.A(men_men_n452_), .B(men_men_n291_), .C(men_men_n451_), .D(men_men_n218_), .Y(men_men_n453_));
  NO2        u431(.A(men_men_n453_), .B(men_men_n141_), .Y(men_men_n454_));
  NA3        u432(.A(men_men_n226_), .B(men_men_n155_), .C(men_men_n119_), .Y(men_men_n455_));
  NO2        u433(.A(men_men_n143_), .B(i_3_), .Y(men_men_n456_));
  NA3        u434(.A(men_men_n367_), .B(men_men_n162_), .C(men_men_n134_), .Y(men_men_n457_));
  NA2        u435(.A(men_men_n457_), .B(men_men_n455_), .Y(men_men_n458_));
  NO4        u436(.A(men_men_n458_), .B(men_men_n454_), .C(men_men_n450_), .D(men_men_n441_), .Y(men_men_n459_));
  NA2        u437(.A(men_men_n425_), .B(men_men_n357_), .Y(men_men_n460_));
  NA2        u438(.A(men_men_n431_), .B(men_men_n363_), .Y(men_men_n461_));
  NO2        u439(.A(men_men_n461_), .B(men_men_n205_), .Y(men_men_n462_));
  NAi21      u440(.An(men_men_n197_), .B(men_men_n372_), .Y(men_men_n463_));
  NO2        u441(.A(men_men_n26_), .B(i_5_), .Y(men_men_n464_));
  NA3        u442(.A(men_men_n1001_), .B(men_men_n464_), .C(men_men_n127_), .Y(men_men_n465_));
  NO2        u443(.A(men_men_n38_), .B(men_men_n465_), .Y(men_men_n466_));
  NA2        u444(.A(men_men_n27_), .B(i_10_), .Y(men_men_n467_));
  NA2        u445(.A(men_men_n291_), .B(men_men_n219_), .Y(men_men_n468_));
  OAI220     u446(.A0(men_men_n468_), .A1(men_men_n405_), .B0(men_men_n467_), .B1(men_men_n437_), .Y(men_men_n469_));
  NA4        u447(.A(men_men_n284_), .B(men_men_n204_), .C(men_men_n65_), .D(men_men_n218_), .Y(men_men_n470_));
  NO2        u448(.A(men_men_n470_), .B(men_men_n444_), .Y(men_men_n471_));
  NO4        u449(.A(men_men_n471_), .B(men_men_n469_), .C(men_men_n466_), .D(men_men_n462_), .Y(men_men_n472_));
  NA4        u450(.A(men_men_n472_), .B(men_men_n459_), .C(men_men_n436_), .D(men_men_n434_), .Y(men_men_n473_));
  NA3        u451(.A(men_men_n284_), .B(men_men_n159_), .C(men_men_n157_), .Y(men_men_n474_));
  OAI210     u452(.A0(men_men_n279_), .A1(men_men_n163_), .B0(men_men_n474_), .Y(men_men_n475_));
  AN2        u453(.A(men_men_n265_), .B(men_men_n215_), .Y(men_men_n476_));
  NA2        u454(.A(men_men_n476_), .B(men_men_n475_), .Y(men_men_n477_));
  NA2        u455(.A(men_men_n291_), .B(men_men_n150_), .Y(men_men_n478_));
  OAI210     u456(.A0(men_men_n478_), .A1(men_men_n213_), .B0(men_men_n285_), .Y(men_men_n479_));
  INV        u457(.A(men_men_n479_), .Y(men_men_n480_));
  NA4        u458(.A(men_men_n416_), .B(men_men_n415_), .C(men_men_n186_), .D(i_2_), .Y(men_men_n481_));
  INV        u459(.A(men_men_n481_), .Y(men_men_n482_));
  NA2        u460(.A(men_men_n357_), .B(men_men_n206_), .Y(men_men_n483_));
  NA2        u461(.A(men_men_n331_), .B(men_men_n65_), .Y(men_men_n484_));
  NA2        u462(.A(men_men_n347_), .B(men_men_n340_), .Y(men_men_n485_));
  AO210      u463(.A0(men_men_n484_), .A1(men_men_n483_), .B0(men_men_n485_), .Y(men_men_n486_));
  NO2        u464(.A(men_men_n36_), .B(i_8_), .Y(men_men_n487_));
  INV        u465(.A(men_men_n486_), .Y(men_men_n488_));
  AOI210     u466(.A0(men_men_n482_), .A1(men_men_n187_), .B0(men_men_n488_), .Y(men_men_n489_));
  OAI210     u467(.A0(i_8_), .A1(men_men_n57_), .B0(men_men_n121_), .Y(men_men_n490_));
  AOI210     u468(.A0(men_men_n177_), .A1(i_9_), .B0(men_men_n245_), .Y(men_men_n491_));
  NO2        u469(.A(men_men_n491_), .B(men_men_n182_), .Y(men_men_n492_));
  AOI220     u470(.A0(i_6_), .A1(men_men_n492_), .B0(men_men_n490_), .B1(men_men_n389_), .Y(men_men_n493_));
  NA4        u471(.A(men_men_n493_), .B(men_men_n489_), .C(men_men_n480_), .D(men_men_n477_), .Y(men_men_n494_));
  NA2        u472(.A(men_men_n362_), .B(men_men_n273_), .Y(men_men_n495_));
  NA2        u473(.A(men_men_n153_), .B(men_men_n495_), .Y(men_men_n496_));
  NO2        u474(.A(i_12_), .B(men_men_n176_), .Y(men_men_n497_));
  NA2        u475(.A(men_men_n497_), .B(men_men_n206_), .Y(men_men_n498_));
  NO3        u476(.A(i_6_), .B(men_men_n498_), .C(men_men_n435_), .Y(men_men_n499_));
  NOi21      u477(.An(men_men_n294_), .B(men_men_n38_), .Y(men_men_n500_));
  OAI210     u478(.A0(men_men_n500_), .A1(men_men_n499_), .B0(men_men_n496_), .Y(men_men_n501_));
  NO2        u479(.A(i_8_), .B(i_7_), .Y(men_men_n502_));
  OAI210     u480(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n503_));
  NA2        u481(.A(men_men_n503_), .B(men_men_n204_), .Y(men_men_n504_));
  AOI220     u482(.A0(men_men_n302_), .A1(men_men_n39_), .B0(men_men_n216_), .B1(men_men_n189_), .Y(men_men_n505_));
  OAI220     u483(.A0(men_men_n505_), .A1(men_men_n165_), .B0(men_men_n504_), .B1(men_men_n223_), .Y(men_men_n506_));
  NA2        u484(.A(men_men_n44_), .B(i_10_), .Y(men_men_n507_));
  NO2        u485(.A(men_men_n507_), .B(i_6_), .Y(men_men_n508_));
  NA3        u486(.A(men_men_n508_), .B(men_men_n506_), .C(men_men_n502_), .Y(men_men_n509_));
  AOI220     u487(.A0(men_men_n398_), .A1(men_men_n302_), .B0(i_2_), .B1(men_men_n225_), .Y(men_men_n510_));
  OAI220     u488(.A0(men_men_n510_), .A1(men_men_n242_), .B0(men_men_n437_), .B1(men_men_n120_), .Y(men_men_n511_));
  NA2        u489(.A(men_men_n511_), .B(men_men_n245_), .Y(men_men_n512_));
  NOi21      u490(.An(men_men_n268_), .B(men_men_n279_), .Y(men_men_n513_));
  NA3        u491(.A(men_men_n284_), .B(men_men_n157_), .C(men_men_n89_), .Y(men_men_n514_));
  NO2        u492(.A(men_men_n203_), .B(men_men_n44_), .Y(men_men_n515_));
  NO2        u493(.A(men_men_n143_), .B(i_5_), .Y(men_men_n516_));
  NA2        u494(.A(men_men_n516_), .B(men_men_n297_), .Y(men_men_n517_));
  OAI210     u495(.A0(men_men_n517_), .A1(men_men_n515_), .B0(men_men_n514_), .Y(men_men_n518_));
  OAI210     u496(.A0(men_men_n518_), .A1(men_men_n513_), .B0(men_men_n431_), .Y(men_men_n519_));
  NA4        u497(.A(men_men_n519_), .B(men_men_n512_), .C(men_men_n509_), .D(men_men_n501_), .Y(men_men_n520_));
  NA3        u498(.A(men_men_n199_), .B(men_men_n63_), .C(men_men_n44_), .Y(men_men_n521_));
  NA2        u499(.A(men_men_n261_), .B(men_men_n75_), .Y(men_men_n522_));
  AOI210     u500(.A0(men_men_n521_), .A1(men_men_n322_), .B0(men_men_n522_), .Y(men_men_n523_));
  NA2        u501(.A(men_men_n274_), .B(men_men_n265_), .Y(men_men_n524_));
  NO2        u502(.A(men_men_n524_), .B(men_men_n156_), .Y(men_men_n525_));
  NA2        u503(.A(men_men_n204_), .B(i_3_), .Y(men_men_n526_));
  NA2        u504(.A(men_men_n418_), .B(men_men_n203_), .Y(men_men_n527_));
  NO2        u505(.A(men_men_n526_), .B(men_men_n527_), .Y(men_men_n528_));
  NA2        u506(.A(i_0_), .B(men_men_n48_), .Y(men_men_n529_));
  NA3        u507(.A(men_men_n497_), .B(men_men_n252_), .C(men_men_n529_), .Y(men_men_n530_));
  NO2        u508(.A(i_2_), .B(men_men_n530_), .Y(men_men_n531_));
  NO4        u509(.A(men_men_n531_), .B(men_men_n528_), .C(men_men_n525_), .D(men_men_n523_), .Y(men_men_n532_));
  NO4        u510(.A(men_men_n230_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n533_));
  NO3        u511(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n534_));
  NO2        u512(.A(men_men_n214_), .B(men_men_n36_), .Y(men_men_n535_));
  AN2        u513(.A(men_men_n535_), .B(men_men_n534_), .Y(men_men_n536_));
  NO2        u514(.A(men_men_n388_), .B(i_1_), .Y(men_men_n537_));
  NOi31      u515(.An(men_men_n537_), .B(men_men_n426_), .C(men_men_n65_), .Y(men_men_n538_));
  AN4        u516(.A(men_men_n538_), .B(men_men_n385_), .C(men_men_n464_), .D(i_2_), .Y(men_men_n539_));
  NO2        u517(.A(men_men_n397_), .B(men_men_n160_), .Y(men_men_n540_));
  NO2        u518(.A(men_men_n540_), .B(men_men_n539_), .Y(men_men_n541_));
  NOi21      u519(.An(i_10_), .B(i_6_), .Y(men_men_n542_));
  NO2        u520(.A(men_men_n77_), .B(men_men_n25_), .Y(men_men_n543_));
  NA2        u521(.A(men_men_n261_), .B(men_men_n543_), .Y(men_men_n544_));
  NO2        u522(.A(men_men_n544_), .B(men_men_n424_), .Y(men_men_n545_));
  NO2        u523(.A(men_men_n105_), .B(men_men_n23_), .Y(men_men_n546_));
  NA2        u524(.A(men_men_n294_), .B(men_men_n150_), .Y(men_men_n547_));
  AOI220     u525(.A0(men_men_n547_), .A1(men_men_n406_), .B0(men_men_n166_), .B1(men_men_n164_), .Y(men_men_n548_));
  NOi21      u526(.An(men_men_n131_), .B(men_men_n310_), .Y(men_men_n549_));
  NO3        u527(.A(men_men_n549_), .B(men_men_n548_), .C(men_men_n545_), .Y(men_men_n550_));
  NO2        u528(.A(men_men_n484_), .B(men_men_n353_), .Y(men_men_n551_));
  INV        u529(.A(men_men_n297_), .Y(men_men_n552_));
  NO2        u530(.A(i_12_), .B(men_men_n77_), .Y(men_men_n553_));
  NA2        u531(.A(men_men_n553_), .B(men_men_n252_), .Y(men_men_n554_));
  NA3        u532(.A(men_men_n359_), .B(men_men_n261_), .C(men_men_n199_), .Y(men_men_n555_));
  AOI210     u533(.A0(men_men_n555_), .A1(men_men_n554_), .B0(men_men_n552_), .Y(men_men_n556_));
  NA2        u534(.A(men_men_n157_), .B(i_0_), .Y(men_men_n557_));
  NO3        u535(.A(men_men_n557_), .B(i_8_), .C(men_men_n279_), .Y(men_men_n558_));
  OR2        u536(.A(i_2_), .B(i_5_), .Y(men_men_n559_));
  AOI210     u537(.A0(men_men_n349_), .A1(men_men_n225_), .B0(men_men_n181_), .Y(men_men_n560_));
  NO2        u538(.A(men_men_n560_), .B(men_men_n463_), .Y(men_men_n561_));
  NO4        u539(.A(men_men_n561_), .B(men_men_n558_), .C(men_men_n556_), .D(men_men_n551_), .Y(men_men_n562_));
  NA4        u540(.A(men_men_n562_), .B(men_men_n550_), .C(men_men_n541_), .D(men_men_n532_), .Y(men_men_n563_));
  NO4        u541(.A(men_men_n563_), .B(men_men_n520_), .C(men_men_n494_), .D(men_men_n473_), .Y(men_men_n564_));
  NA4        u542(.A(men_men_n564_), .B(men_men_n414_), .C(men_men_n330_), .D(men_men_n290_), .Y(men7));
  NO2        u543(.A(men_men_n99_), .B(men_men_n82_), .Y(men_men_n566_));
  NA2        u544(.A(men_men_n358_), .B(men_men_n566_), .Y(men_men_n567_));
  NA2        u545(.A(men_men_n452_), .B(men_men_n75_), .Y(men_men_n568_));
  NA2        u546(.A(men_men_n129_), .B(i_8_), .Y(men_men_n569_));
  OAI210     u547(.A0(men_men_n569_), .A1(men_men_n568_), .B0(men_men_n567_), .Y(men_men_n570_));
  NA3        u548(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n571_));
  NO2        u549(.A(men_men_n218_), .B(i_4_), .Y(men_men_n572_));
  NA2        u550(.A(men_men_n572_), .B(i_8_), .Y(men_men_n573_));
  NA2        u551(.A(i_2_), .B(men_men_n77_), .Y(men_men_n574_));
  OAI210     u552(.A0(men_men_n80_), .A1(men_men_n186_), .B0(men_men_n187_), .Y(men_men_n575_));
  NO2        u553(.A(i_7_), .B(men_men_n37_), .Y(men_men_n576_));
  NA2        u554(.A(i_4_), .B(i_8_), .Y(men_men_n577_));
  AOI210     u555(.A0(men_men_n577_), .A1(men_men_n284_), .B0(men_men_n576_), .Y(men_men_n578_));
  OAI220     u556(.A0(men_men_n578_), .A1(men_men_n574_), .B0(men_men_n575_), .B1(i_13_), .Y(men_men_n579_));
  NO2        u557(.A(men_men_n579_), .B(men_men_n570_), .Y(men_men_n580_));
  OR2        u558(.A(i_6_), .B(i_10_), .Y(men_men_n581_));
  NO2        u559(.A(men_men_n581_), .B(men_men_n23_), .Y(men_men_n582_));
  OR3        u560(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n583_));
  NO3        u561(.A(men_men_n583_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n584_));
  INV        u562(.A(men_men_n183_), .Y(men_men_n585_));
  INV        u563(.A(men_men_n584_), .Y(men_men_n586_));
  OR2        u564(.A(men_men_n586_), .B(men_men_n552_), .Y(men_men_n587_));
  AOI210     u565(.A0(men_men_n587_), .A1(men_men_n580_), .B0(men_men_n57_), .Y(men_men_n588_));
  NOi21      u566(.An(i_11_), .B(i_7_), .Y(men_men_n589_));
  AO210      u567(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n590_));
  NO2        u568(.A(men_men_n590_), .B(men_men_n589_), .Y(men_men_n591_));
  NA2        u569(.A(men_men_n591_), .B(men_men_n189_), .Y(men_men_n592_));
  NA3        u570(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n593_));
  NAi31      u571(.An(men_men_n593_), .B(men_men_n196_), .C(i_11_), .Y(men_men_n594_));
  AOI210     u572(.A0(men_men_n594_), .A1(men_men_n592_), .B0(men_men_n57_), .Y(men_men_n595_));
  NA2        u573(.A(men_men_n79_), .B(men_men_n57_), .Y(men_men_n596_));
  AO210      u574(.A0(men_men_n596_), .A1(men_men_n353_), .B0(men_men_n40_), .Y(men_men_n597_));
  NO3        u575(.A(men_men_n237_), .B(men_men_n190_), .C(i_8_), .Y(men_men_n598_));
  OAI210     u576(.A0(men_men_n598_), .A1(men_men_n207_), .B0(men_men_n57_), .Y(men_men_n599_));
  NA2        u577(.A(men_men_n382_), .B(men_men_n31_), .Y(men_men_n600_));
  OR2        u578(.A(men_men_n190_), .B(men_men_n99_), .Y(men_men_n601_));
  NA2        u579(.A(men_men_n601_), .B(men_men_n600_), .Y(men_men_n602_));
  NO2        u580(.A(men_men_n57_), .B(i_9_), .Y(men_men_n603_));
  NO2        u581(.A(men_men_n603_), .B(i_4_), .Y(men_men_n604_));
  NA2        u582(.A(men_men_n604_), .B(men_men_n602_), .Y(men_men_n605_));
  NO2        u583(.A(i_1_), .B(i_12_), .Y(men_men_n606_));
  NA3        u584(.A(men_men_n606_), .B(men_men_n101_), .C(men_men_n24_), .Y(men_men_n607_));
  NA4        u585(.A(men_men_n607_), .B(men_men_n605_), .C(men_men_n599_), .D(men_men_n597_), .Y(men_men_n608_));
  OAI210     u586(.A0(men_men_n608_), .A1(men_men_n595_), .B0(i_6_), .Y(men_men_n609_));
  NO2        u587(.A(men_men_n593_), .B(men_men_n99_), .Y(men_men_n610_));
  NA2        u588(.A(men_men_n610_), .B(men_men_n553_), .Y(men_men_n611_));
  NO2        u589(.A(i_6_), .B(i_11_), .Y(men_men_n612_));
  NA2        u590(.A(men_men_n611_), .B(men_men_n427_), .Y(men_men_n613_));
  NO4        u591(.A(men_men_n196_), .B(men_men_n115_), .C(i_13_), .D(men_men_n77_), .Y(men_men_n614_));
  NA2        u592(.A(men_men_n614_), .B(men_men_n603_), .Y(men_men_n615_));
  NO3        u593(.A(men_men_n581_), .B(men_men_n214_), .C(men_men_n23_), .Y(men_men_n616_));
  AOI210     u594(.A0(i_1_), .A1(men_men_n238_), .B0(men_men_n616_), .Y(men_men_n617_));
  OAI210     u595(.A0(men_men_n617_), .A1(men_men_n44_), .B0(men_men_n615_), .Y(men_men_n618_));
  NA3        u596(.A(men_men_n502_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n619_));
  NA2        u597(.A(men_men_n125_), .B(i_9_), .Y(men_men_n620_));
  NA3        u598(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n621_));
  NO2        u599(.A(men_men_n46_), .B(i_1_), .Y(men_men_n622_));
  NA3        u600(.A(men_men_n622_), .B(men_men_n246_), .C(men_men_n44_), .Y(men_men_n623_));
  OAI220     u601(.A0(men_men_n623_), .A1(men_men_n621_), .B0(men_men_n620_), .B1(men_men_n997_), .Y(men_men_n624_));
  NA3        u602(.A(men_men_n603_), .B(men_men_n297_), .C(i_6_), .Y(men_men_n625_));
  NO2        u603(.A(men_men_n625_), .B(men_men_n23_), .Y(men_men_n626_));
  NO2        u604(.A(i_11_), .B(men_men_n37_), .Y(men_men_n627_));
  NA2        u605(.A(men_men_n627_), .B(men_men_n24_), .Y(men_men_n628_));
  NO2        u606(.A(men_men_n628_), .B(men_men_n46_), .Y(men_men_n629_));
  OR3        u607(.A(men_men_n629_), .B(men_men_n626_), .C(men_men_n624_), .Y(men_men_n630_));
  NO3        u608(.A(men_men_n630_), .B(men_men_n618_), .C(men_men_n613_), .Y(men_men_n631_));
  NO2        u609(.A(men_men_n218_), .B(men_men_n94_), .Y(men_men_n632_));
  NO2        u610(.A(men_men_n632_), .B(men_men_n589_), .Y(men_men_n633_));
  NA2        u611(.A(men_men_n633_), .B(i_1_), .Y(men_men_n634_));
  NO2        u612(.A(men_men_n634_), .B(men_men_n583_), .Y(men_men_n635_));
  NO2        u613(.A(men_men_n387_), .B(men_men_n77_), .Y(men_men_n636_));
  NA2        u614(.A(men_men_n635_), .B(men_men_n46_), .Y(men_men_n637_));
  NA2        u615(.A(i_3_), .B(men_men_n176_), .Y(men_men_n638_));
  NO2        u616(.A(men_men_n638_), .B(men_men_n105_), .Y(men_men_n639_));
  AN2        u617(.A(men_men_n639_), .B(men_men_n508_), .Y(men_men_n640_));
  NO2        u618(.A(men_men_n214_), .B(men_men_n44_), .Y(men_men_n641_));
  NO2        u619(.A(men_men_n106_), .B(men_men_n37_), .Y(men_men_n642_));
  NA2        u620(.A(i_1_), .B(i_3_), .Y(men_men_n643_));
  NO2        u621(.A(men_men_n428_), .B(men_men_n85_), .Y(men_men_n644_));
  AOI210     u622(.A0(men_men_n641_), .A1(men_men_n542_), .B0(men_men_n644_), .Y(men_men_n645_));
  NO2        u623(.A(men_men_n645_), .B(men_men_n643_), .Y(men_men_n646_));
  NO2        u624(.A(men_men_n646_), .B(men_men_n640_), .Y(men_men_n647_));
  NA4        u625(.A(men_men_n647_), .B(men_men_n637_), .C(men_men_n631_), .D(men_men_n609_), .Y(men_men_n648_));
  NO3        u626(.A(men_men_n445_), .B(i_3_), .C(i_7_), .Y(men_men_n649_));
  NOi21      u627(.An(men_men_n649_), .B(i_10_), .Y(men_men_n650_));
  AN2        u628(.A(men_men_n650_), .B(men_men_n77_), .Y(men_men_n651_));
  NA2        u629(.A(men_men_n347_), .B(men_men_n346_), .Y(men_men_n652_));
  NO3        u630(.A(men_men_n446_), .B(men_men_n577_), .C(men_men_n77_), .Y(men_men_n653_));
  NA2        u631(.A(men_men_n653_), .B(men_men_n25_), .Y(men_men_n654_));
  NA2        u632(.A(men_men_n147_), .B(men_men_n77_), .Y(men_men_n655_));
  NA3        u633(.A(men_men_n655_), .B(men_men_n654_), .C(men_men_n652_), .Y(men_men_n656_));
  OAI210     u634(.A0(men_men_n656_), .A1(men_men_n651_), .B0(i_1_), .Y(men_men_n657_));
  NO2        u635(.A(men_men_n625_), .B(men_men_n419_), .Y(men_men_n658_));
  INV        u636(.A(men_men_n658_), .Y(men_men_n659_));
  AOI210     u637(.A0(men_men_n659_), .A1(men_men_n657_), .B0(i_13_), .Y(men_men_n660_));
  OR2        u638(.A(i_11_), .B(i_7_), .Y(men_men_n661_));
  NA3        u639(.A(men_men_n661_), .B(men_men_n98_), .C(men_men_n125_), .Y(men_men_n662_));
  AOI220     u640(.A0(men_men_n439_), .A1(men_men_n147_), .B0(men_men_n1002_), .B1(men_men_n125_), .Y(men_men_n663_));
  OAI210     u641(.A0(men_men_n663_), .A1(men_men_n44_), .B0(men_men_n662_), .Y(men_men_n664_));
  AOI220     u642(.A0(i_7_), .A1(men_men_n636_), .B0(men_men_n226_), .B1(men_men_n118_), .Y(men_men_n665_));
  OAI220     u643(.A0(men_men_n665_), .A1(men_men_n40_), .B0(men_men_n52_), .B1(men_men_n85_), .Y(men_men_n666_));
  AOI210     u644(.A0(men_men_n664_), .A1(men_men_n312_), .B0(men_men_n666_), .Y(men_men_n667_));
  AOI220     u645(.A0(i_12_), .A1(men_men_n64_), .B0(men_men_n359_), .B1(men_men_n622_), .Y(men_men_n668_));
  NO2        u646(.A(men_men_n668_), .B(men_men_n223_), .Y(men_men_n669_));
  AOI210     u647(.A0(men_men_n419_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n670_));
  NA2        u648(.A(men_men_n114_), .B(i_13_), .Y(men_men_n671_));
  NO2        u649(.A(men_men_n621_), .B(men_men_n105_), .Y(men_men_n672_));
  INV        u650(.A(men_men_n672_), .Y(men_men_n673_));
  OAI220     u651(.A0(men_men_n673_), .A1(men_men_n63_), .B0(men_men_n671_), .B1(men_men_n1006_), .Y(men_men_n674_));
  NO3        u652(.A(men_men_n63_), .B(men_men_n32_), .C(men_men_n94_), .Y(men_men_n675_));
  NA2        u653(.A(men_men_n26_), .B(men_men_n176_), .Y(men_men_n676_));
  INV        u654(.A(men_men_n675_), .Y(men_men_n677_));
  AOI210     u655(.A0(men_men_n359_), .A1(men_men_n622_), .B0(men_men_n84_), .Y(men_men_n678_));
  OAI220     u656(.A0(men_men_n678_), .A1(men_men_n573_), .B0(men_men_n677_), .B1(men_men_n585_), .Y(men_men_n679_));
  NO3        u657(.A(men_men_n679_), .B(men_men_n674_), .C(men_men_n669_), .Y(men_men_n680_));
  NA3        u658(.A(men_men_n382_), .B(men_men_n576_), .C(men_men_n90_), .Y(men_men_n681_));
  NA2        u659(.A(men_men_n612_), .B(i_13_), .Y(men_men_n682_));
  INV        u660(.A(men_men_n676_), .Y(men_men_n683_));
  NAi21      u661(.An(i_11_), .B(i_12_), .Y(men_men_n684_));
  NO3        u662(.A(men_men_n684_), .B(i_13_), .C(men_men_n77_), .Y(men_men_n685_));
  NO3        u663(.A(men_men_n446_), .B(men_men_n553_), .C(men_men_n577_), .Y(men_men_n686_));
  AOI220     u664(.A0(men_men_n686_), .A1(men_men_n291_), .B0(men_men_n685_), .B1(men_men_n683_), .Y(men_men_n687_));
  NA3        u665(.A(men_men_n687_), .B(men_men_n682_), .C(men_men_n681_), .Y(men_men_n688_));
  NA2        u666(.A(men_men_n688_), .B(men_men_n57_), .Y(men_men_n689_));
  NO2        u667(.A(i_2_), .B(i_12_), .Y(men_men_n690_));
  NA2        u668(.A(men_men_n344_), .B(men_men_n690_), .Y(men_men_n691_));
  NA2        u669(.A(i_8_), .B(men_men_n25_), .Y(men_men_n692_));
  NO2        u670(.A(men_men_n692_), .B(men_men_n358_), .Y(men_men_n693_));
  OAI210     u671(.A0(men_men_n693_), .A1(men_men_n346_), .B0(men_men_n344_), .Y(men_men_n694_));
  NO2        u672(.A(men_men_n115_), .B(i_2_), .Y(men_men_n695_));
  NA2        u673(.A(men_men_n695_), .B(men_men_n606_), .Y(men_men_n696_));
  NA3        u674(.A(men_men_n696_), .B(men_men_n694_), .C(men_men_n691_), .Y(men_men_n697_));
  NA3        u675(.A(men_men_n697_), .B(men_men_n45_), .C(men_men_n206_), .Y(men_men_n698_));
  NA4        u676(.A(men_men_n698_), .B(men_men_n689_), .C(men_men_n680_), .D(men_men_n667_), .Y(men_men_n699_));
  OR4        u677(.A(men_men_n699_), .B(men_men_n660_), .C(men_men_n648_), .D(men_men_n588_), .Y(men5));
  AOI210     u678(.A0(men_men_n633_), .A1(men_men_n248_), .B0(men_men_n389_), .Y(men_men_n701_));
  NA3        u679(.A(men_men_n24_), .B(men_men_n690_), .C(men_men_n99_), .Y(men_men_n702_));
  NA2        u680(.A(men_men_n702_), .B(men_men_n701_), .Y(men_men_n703_));
  NO3        u681(.A(i_11_), .B(men_men_n218_), .C(i_13_), .Y(men_men_n704_));
  NO2        u682(.A(men_men_n112_), .B(men_men_n23_), .Y(men_men_n705_));
  NA2        u683(.A(i_12_), .B(i_8_), .Y(men_men_n706_));
  OAI210     u684(.A0(men_men_n46_), .A1(i_3_), .B0(men_men_n706_), .Y(men_men_n707_));
  INV        u685(.A(men_men_n418_), .Y(men_men_n708_));
  AOI220     u686(.A0(men_men_n297_), .A1(men_men_n546_), .B0(men_men_n707_), .B1(men_men_n705_), .Y(men_men_n709_));
  INV        u687(.A(men_men_n709_), .Y(men_men_n710_));
  NO2        u688(.A(men_men_n710_), .B(men_men_n703_), .Y(men_men_n711_));
  INV        u689(.A(men_men_n155_), .Y(men_men_n712_));
  NO2        u690(.A(men_men_n428_), .B(men_men_n26_), .Y(men_men_n713_));
  NO2        u691(.A(men_men_n713_), .B(men_men_n390_), .Y(men_men_n714_));
  NA2        u692(.A(men_men_n714_), .B(i_2_), .Y(men_men_n715_));
  INV        u693(.A(men_men_n715_), .Y(men_men_n716_));
  AOI210     u694(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n388_), .Y(men_men_n717_));
  AOI210     u695(.A0(men_men_n717_), .A1(men_men_n716_), .B0(men_men_n226_), .Y(men_men_n718_));
  NO2        u696(.A(men_men_n173_), .B(men_men_n113_), .Y(men_men_n719_));
  OAI210     u697(.A0(men_men_n719_), .A1(men_men_n705_), .B0(i_2_), .Y(men_men_n720_));
  NO3        u698(.A(men_men_n590_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n721_));
  AOI210     u699(.A0(men_men_n155_), .A1(men_men_n80_), .B0(men_men_n721_), .Y(men_men_n722_));
  AOI210     u700(.A0(men_men_n722_), .A1(men_men_n720_), .B0(men_men_n176_), .Y(men_men_n723_));
  NA2        u701(.A(men_men_n183_), .B(men_men_n186_), .Y(men_men_n724_));
  NA2        u702(.A(men_men_n137_), .B(i_8_), .Y(men_men_n725_));
  AOI210     u703(.A0(men_men_n725_), .A1(men_men_n724_), .B0(men_men_n349_), .Y(men_men_n726_));
  NA2        u704(.A(men_men_n190_), .B(men_men_n133_), .Y(men_men_n727_));
  NA2        u705(.A(men_men_n727_), .B(men_men_n390_), .Y(men_men_n728_));
  NA3        u706(.A(men_men_n284_), .B(men_men_n112_), .C(men_men_n42_), .Y(men_men_n729_));
  OAI210     u707(.A0(men_men_n729_), .A1(men_men_n46_), .B0(men_men_n728_), .Y(men_men_n730_));
  NO3        u708(.A(men_men_n730_), .B(men_men_n726_), .C(men_men_n723_), .Y(men_men_n731_));
  NA2        u709(.A(men_men_n546_), .B(men_men_n28_), .Y(men_men_n732_));
  NA2        u710(.A(men_men_n704_), .B(men_men_n253_), .Y(men_men_n733_));
  NA2        u711(.A(men_men_n733_), .B(men_men_n732_), .Y(men_men_n734_));
  INV        u712(.A(men_men_n734_), .Y(men_men_n735_));
  NA4        u713(.A(men_men_n735_), .B(men_men_n731_), .C(men_men_n718_), .D(men_men_n711_), .Y(men6));
  NA2        u714(.A(men_men_n25_), .B(men_men_n695_), .Y(men_men_n737_));
  NA4        u715(.A(men_men_n363_), .B(men_men_n451_), .C(men_men_n63_), .D(men_men_n94_), .Y(men_men_n738_));
  INV        u716(.A(men_men_n738_), .Y(men_men_n739_));
  NO2        u717(.A(men_men_n202_), .B(i_2_), .Y(men_men_n740_));
  NO2        u718(.A(i_11_), .B(i_9_), .Y(men_men_n741_));
  NO2        u719(.A(men_men_n739_), .B(men_men_n307_), .Y(men_men_n742_));
  AO210      u720(.A0(men_men_n742_), .A1(men_men_n737_), .B0(i_12_), .Y(men_men_n743_));
  NA2        u721(.A(men_men_n350_), .B(men_men_n315_), .Y(men_men_n744_));
  NA2        u722(.A(men_men_n553_), .B(men_men_n57_), .Y(men_men_n745_));
  NA2        u723(.A(men_men_n650_), .B(men_men_n63_), .Y(men_men_n746_));
  NA4        u724(.A(men_men_n596_), .B(men_men_n746_), .C(men_men_n745_), .D(men_men_n744_), .Y(men_men_n747_));
  INV        u725(.A(men_men_n180_), .Y(men_men_n748_));
  AOI220     u726(.A0(men_men_n748_), .A1(men_men_n741_), .B0(men_men_n747_), .B1(men_men_n65_), .Y(men_men_n749_));
  INV        u727(.A(men_men_n306_), .Y(men_men_n750_));
  NA2        u728(.A(men_men_n67_), .B(men_men_n118_), .Y(men_men_n751_));
  INV        u729(.A(men_men_n112_), .Y(men_men_n752_));
  NA2        u730(.A(men_men_n752_), .B(men_men_n46_), .Y(men_men_n753_));
  AOI210     u731(.A0(men_men_n753_), .A1(men_men_n751_), .B0(men_men_n750_), .Y(men_men_n754_));
  INV        u732(.A(men_men_n485_), .Y(men_men_n755_));
  NO2        u733(.A(men_men_n32_), .B(i_11_), .Y(men_men_n756_));
  NA3        u734(.A(men_men_n756_), .B(men_men_n443_), .C(men_men_n363_), .Y(men_men_n757_));
  OAI210     u735(.A0(men_men_n649_), .A1(men_men_n535_), .B0(men_men_n534_), .Y(men_men_n758_));
  NA2        u736(.A(men_men_n758_), .B(men_men_n757_), .Y(men_men_n759_));
  OR3        u737(.A(men_men_n759_), .B(men_men_n755_), .C(men_men_n754_), .Y(men_men_n760_));
  NA3        u738(.A(men_men_n326_), .B(men_men_n235_), .C(i_7_), .Y(men_men_n761_));
  NA2        u739(.A(men_men_n420_), .B(men_men_n132_), .Y(men_men_n762_));
  AO210      u740(.A0(men_men_n461_), .A1(men_men_n708_), .B0(men_men_n36_), .Y(men_men_n763_));
  NA3        u741(.A(men_men_n763_), .B(men_men_n762_), .C(men_men_n761_), .Y(men_men_n764_));
  OAI210     u742(.A0(i_6_), .A1(i_11_), .B0(men_men_n78_), .Y(men_men_n765_));
  AOI220     u743(.A0(men_men_n765_), .A1(men_men_n534_), .B0(men_men_n740_), .B1(men_men_n1009_), .Y(men_men_n766_));
  NA3        u744(.A(men_men_n349_), .B(men_men_n219_), .C(men_men_n132_), .Y(men_men_n767_));
  OAI210     u745(.A0(men_men_n370_), .A1(men_men_n187_), .B0(men_men_n62_), .Y(men_men_n768_));
  NA4        u746(.A(men_men_n768_), .B(men_men_n767_), .C(men_men_n766_), .D(men_men_n575_), .Y(men_men_n769_));
  AO210      u747(.A0(men_men_n487_), .A1(men_men_n46_), .B0(men_men_n79_), .Y(men_men_n770_));
  NA3        u748(.A(men_men_n770_), .B(men_men_n452_), .C(men_men_n199_), .Y(men_men_n771_));
  INV        u749(.A(men_men_n533_), .Y(men_men_n772_));
  NO2        u750(.A(men_men_n581_), .B(i_2_), .Y(men_men_n773_));
  OAI210     u751(.A0(men_men_n773_), .A1(men_men_n102_), .B0(men_men_n380_), .Y(men_men_n774_));
  INV        u752(.A(men_men_n559_), .Y(men_men_n775_));
  NA3        u753(.A(men_men_n775_), .B(men_men_n306_), .C(i_7_), .Y(men_men_n776_));
  NA4        u754(.A(men_men_n776_), .B(men_men_n774_), .C(men_men_n772_), .D(men_men_n771_), .Y(men_men_n777_));
  NO4        u755(.A(men_men_n777_), .B(men_men_n769_), .C(men_men_n764_), .D(men_men_n760_), .Y(men_men_n778_));
  NA4        u756(.A(men_men_n778_), .B(men_men_n749_), .C(men_men_n743_), .D(men_men_n354_), .Y(men3));
  NA2        u757(.A(i_12_), .B(i_10_), .Y(men_men_n780_));
  NA2        u758(.A(i_6_), .B(i_7_), .Y(men_men_n781_));
  NO2        u759(.A(men_men_n781_), .B(i_0_), .Y(men_men_n782_));
  NO2        u760(.A(i_11_), .B(men_men_n218_), .Y(men_men_n783_));
  NA2        u761(.A(men_men_n268_), .B(men_men_n783_), .Y(men_men_n784_));
  NO2        u762(.A(men_men_n784_), .B(men_men_n176_), .Y(men_men_n785_));
  NO3        u763(.A(men_men_n424_), .B(men_men_n82_), .C(men_men_n44_), .Y(men_men_n786_));
  OA210      u764(.A0(men_men_n786_), .A1(men_men_n785_), .B0(men_men_n157_), .Y(men_men_n787_));
  NA3        u765(.A(men_men_n767_), .B(men_men_n575_), .C(men_men_n348_), .Y(men_men_n788_));
  NA2        u766(.A(men_men_n788_), .B(men_men_n39_), .Y(men_men_n789_));
  NO3        u767(.A(men_men_n601_), .B(men_men_n428_), .C(men_men_n118_), .Y(men_men_n790_));
  NA2        u768(.A(men_men_n382_), .B(men_men_n45_), .Y(men_men_n791_));
  AN2        u769(.A(men_men_n426_), .B(men_men_n53_), .Y(men_men_n792_));
  NO2        u770(.A(men_men_n792_), .B(men_men_n790_), .Y(men_men_n793_));
  AOI210     u771(.A0(men_men_n793_), .A1(men_men_n789_), .B0(men_men_n48_), .Y(men_men_n794_));
  NA2        u772(.A(men_men_n670_), .B(men_men_n1003_), .Y(men_men_n795_));
  NA2        u773(.A(men_men_n313_), .B(men_men_n408_), .Y(men_men_n796_));
  NO2        u774(.A(men_men_n796_), .B(men_men_n795_), .Y(men_men_n797_));
  NOi21      u775(.An(i_5_), .B(i_9_), .Y(men_men_n798_));
  NA2        u776(.A(men_men_n798_), .B(men_men_n416_), .Y(men_men_n799_));
  INV        u777(.A(men_men_n653_), .Y(men_men_n800_));
  NO2        u778(.A(men_men_n800_), .B(men_men_n799_), .Y(men_men_n801_));
  NO4        u779(.A(men_men_n801_), .B(men_men_n797_), .C(men_men_n794_), .D(men_men_n787_), .Y(men_men_n802_));
  NA2        u780(.A(men_men_n168_), .B(men_men_n24_), .Y(men_men_n803_));
  NO2        u781(.A(men_men_n642_), .B(men_men_n566_), .Y(men_men_n804_));
  NO2        u782(.A(men_men_n804_), .B(men_men_n803_), .Y(men_men_n805_));
  NA2        u783(.A(men_men_n291_), .B(men_men_n116_), .Y(men_men_n806_));
  NAi21      u784(.An(men_men_n148_), .B(men_men_n408_), .Y(men_men_n807_));
  NO2        u785(.A(men_men_n806_), .B(men_men_n373_), .Y(men_men_n808_));
  NO2        u786(.A(men_men_n808_), .B(men_men_n805_), .Y(men_men_n809_));
  NO2        u787(.A(men_men_n363_), .B(men_men_n272_), .Y(men_men_n810_));
  NA2        u788(.A(men_men_n810_), .B(men_men_n672_), .Y(men_men_n811_));
  NA2        u789(.A(men_men_n543_), .B(i_0_), .Y(men_men_n812_));
  NO3        u790(.A(men_men_n812_), .B(men_men_n1007_), .C(men_men_n80_), .Y(men_men_n813_));
  NO4        u791(.A(men_men_n559_), .B(men_men_n196_), .C(men_men_n388_), .D(i_6_), .Y(men_men_n814_));
  INV        u792(.A(men_men_n813_), .Y(men_men_n815_));
  AN2        u793(.A(men_men_n89_), .B(men_men_n224_), .Y(men_men_n816_));
  NA2        u794(.A(men_men_n704_), .B(men_men_n307_), .Y(men_men_n817_));
  AOI210     u795(.A0(men_men_n452_), .A1(men_men_n80_), .B0(men_men_n54_), .Y(men_men_n818_));
  OAI220     u796(.A0(men_men_n818_), .A1(men_men_n817_), .B0(men_men_n628_), .B1(men_men_n504_), .Y(men_men_n819_));
  NA2        u797(.A(i_0_), .B(i_10_), .Y(men_men_n820_));
  NO4        u798(.A(men_men_n105_), .B(men_men_n54_), .C(men_men_n638_), .D(i_5_), .Y(men_men_n821_));
  AN2        u799(.A(men_men_n821_), .B(i_10_), .Y(men_men_n822_));
  AOI220     u800(.A0(men_men_n313_), .A1(men_men_n91_), .B0(men_men_n168_), .B1(men_men_n75_), .Y(men_men_n823_));
  NA2        u801(.A(men_men_n537_), .B(i_4_), .Y(men_men_n824_));
  NA2        u802(.A(men_men_n171_), .B(men_men_n186_), .Y(men_men_n825_));
  OAI220     u803(.A0(men_men_n825_), .A1(men_men_n817_), .B0(men_men_n824_), .B1(men_men_n823_), .Y(men_men_n826_));
  NO4        u804(.A(men_men_n826_), .B(men_men_n822_), .C(men_men_n819_), .D(men_men_n816_), .Y(men_men_n827_));
  NA4        u805(.A(men_men_n827_), .B(men_men_n815_), .C(men_men_n811_), .D(men_men_n809_), .Y(men_men_n828_));
  NO2        u806(.A(men_men_n95_), .B(men_men_n37_), .Y(men_men_n829_));
  NA2        u807(.A(i_11_), .B(i_9_), .Y(men_men_n830_));
  NO3        u808(.A(i_12_), .B(men_men_n830_), .C(men_men_n574_), .Y(men_men_n831_));
  AN2        u809(.A(men_men_n831_), .B(men_men_n829_), .Y(men_men_n832_));
  NO2        u810(.A(men_men_n48_), .B(i_7_), .Y(men_men_n833_));
  NA2        u811(.A(men_men_n367_), .B(men_men_n162_), .Y(men_men_n834_));
  NA2        u812(.A(men_men_n834_), .B(men_men_n146_), .Y(men_men_n835_));
  NO2        u813(.A(men_men_n830_), .B(men_men_n65_), .Y(men_men_n836_));
  NO2        u814(.A(men_men_n158_), .B(i_0_), .Y(men_men_n837_));
  INV        u815(.A(men_men_n837_), .Y(men_men_n838_));
  NA2        u816(.A(men_men_n443_), .B(men_men_n212_), .Y(men_men_n839_));
  AOI210     u817(.A0(men_men_n347_), .A1(men_men_n41_), .B0(men_men_n379_), .Y(men_men_n840_));
  OAI220     u818(.A0(men_men_n840_), .A1(men_men_n799_), .B0(men_men_n839_), .B1(men_men_n838_), .Y(men_men_n841_));
  NO3        u819(.A(men_men_n841_), .B(men_men_n835_), .C(men_men_n832_), .Y(men_men_n842_));
  NA2        u820(.A(men_men_n627_), .B(men_men_n109_), .Y(men_men_n843_));
  NO2        u821(.A(i_6_), .B(men_men_n843_), .Y(men_men_n844_));
  AOI210     u822(.A0(men_men_n419_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n845_));
  NA2        u823(.A(men_men_n155_), .B(men_men_n95_), .Y(men_men_n846_));
  NOi32      u824(.An(men_men_n845_), .Bn(men_men_n171_), .C(men_men_n846_), .Y(men_men_n847_));
  NO2        u825(.A(men_men_n1000_), .B(men_men_n791_), .Y(men_men_n848_));
  NO3        u826(.A(men_men_n848_), .B(men_men_n847_), .C(men_men_n844_), .Y(men_men_n849_));
  NOi21      u827(.An(i_7_), .B(i_5_), .Y(men_men_n850_));
  NOi31      u828(.An(men_men_n850_), .B(i_0_), .C(men_men_n684_), .Y(men_men_n851_));
  NA3        u829(.A(men_men_n851_), .B(men_men_n358_), .C(i_6_), .Y(men_men_n852_));
  OA210      u830(.A0(men_men_n846_), .A1(men_men_n485_), .B0(men_men_n852_), .Y(men_men_n853_));
  NO3        u831(.A(men_men_n376_), .B(men_men_n337_), .C(men_men_n333_), .Y(men_men_n854_));
  INV        u832(.A(men_men_n298_), .Y(men_men_n855_));
  INV        u833(.A(men_men_n854_), .Y(men_men_n856_));
  NA4        u834(.A(men_men_n856_), .B(men_men_n853_), .C(men_men_n849_), .D(men_men_n842_), .Y(men_men_n857_));
  NO2        u835(.A(men_men_n803_), .B(men_men_n220_), .Y(men_men_n858_));
  AN2        u836(.A(men_men_n312_), .B(men_men_n307_), .Y(men_men_n859_));
  NA2        u837(.A(men_men_n858_), .B(i_10_), .Y(men_men_n860_));
  NO2        u838(.A(men_men_n780_), .B(men_men_n297_), .Y(men_men_n861_));
  OA210      u839(.A0(men_men_n443_), .A1(men_men_n204_), .B0(men_men_n442_), .Y(men_men_n862_));
  NA2        u840(.A(men_men_n861_), .B(men_men_n836_), .Y(men_men_n863_));
  NO2        u841(.A(men_men_n807_), .B(i_6_), .Y(men_men_n864_));
  NO2        u842(.A(men_men_n235_), .B(men_men_n46_), .Y(men_men_n865_));
  NA2        u843(.A(men_men_n836_), .B(men_men_n284_), .Y(men_men_n866_));
  OAI210     u844(.A0(men_men_n865_), .A1(men_men_n170_), .B0(men_men_n866_), .Y(men_men_n867_));
  AOI220     u845(.A0(men_men_n867_), .A1(men_men_n443_), .B0(men_men_n864_), .B1(men_men_n65_), .Y(men_men_n868_));
  NO2        u846(.A(men_men_n67_), .B(men_men_n706_), .Y(men_men_n869_));
  AOI220     u847(.A0(men_men_n869_), .A1(i_11_), .B0(men_men_n157_), .B1(men_men_n566_), .Y(men_men_n870_));
  NO2        u848(.A(men_men_n870_), .B(men_men_n47_), .Y(men_men_n871_));
  NO3        u849(.A(men_men_n559_), .B(i_0_), .C(men_men_n24_), .Y(men_men_n872_));
  AOI210     u850(.A0(i_7_), .A1(men_men_n516_), .B0(men_men_n872_), .Y(men_men_n873_));
  NAi21      u851(.An(i_9_), .B(i_5_), .Y(men_men_n874_));
  NO2        u852(.A(men_men_n874_), .B(men_men_n376_), .Y(men_men_n875_));
  NO2        u853(.A(men_men_n571_), .B(men_men_n97_), .Y(men_men_n876_));
  AOI220     u854(.A0(men_men_n876_), .A1(i_0_), .B0(men_men_n875_), .B1(men_men_n591_), .Y(men_men_n877_));
  OAI220     u855(.A0(men_men_n877_), .A1(men_men_n77_), .B0(men_men_n873_), .B1(men_men_n156_), .Y(men_men_n878_));
  NO3        u856(.A(men_men_n878_), .B(men_men_n871_), .C(men_men_n488_), .Y(men_men_n879_));
  NA4        u857(.A(men_men_n879_), .B(men_men_n868_), .C(men_men_n863_), .D(men_men_n860_), .Y(men_men_n880_));
  NO3        u858(.A(men_men_n880_), .B(men_men_n857_), .C(men_men_n828_), .Y(men_men_n881_));
  NO2        u859(.A(i_0_), .B(men_men_n684_), .Y(men_men_n882_));
  NA2        u860(.A(men_men_n65_), .B(men_men_n44_), .Y(men_men_n883_));
  NO3        u861(.A(men_men_n97_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n884_));
  AO220      u862(.A0(men_men_n884_), .A1(men_men_n65_), .B0(men_men_n882_), .B1(men_men_n157_), .Y(men_men_n885_));
  AOI210     u863(.A0(men_men_n745_), .A1(men_men_n652_), .B0(men_men_n846_), .Y(men_men_n886_));
  AOI210     u864(.A0(men_men_n885_), .A1(men_men_n323_), .B0(men_men_n886_), .Y(men_men_n887_));
  NA2        u865(.A(men_men_n695_), .B(men_men_n131_), .Y(men_men_n888_));
  NO2        u866(.A(men_men_n758_), .B(men_men_n376_), .Y(men_men_n889_));
  NA3        u867(.A(men_men_n782_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n890_));
  NA2        u868(.A(men_men_n783_), .B(i_9_), .Y(men_men_n891_));
  AOI210     u869(.A0(men_men_n890_), .A1(men_men_n465_), .B0(men_men_n891_), .Y(men_men_n892_));
  OAI210     u870(.A0(men_men_n225_), .A1(i_9_), .B0(men_men_n211_), .Y(men_men_n893_));
  AOI210     u871(.A0(men_men_n893_), .A1(men_men_n812_), .B0(men_men_n139_), .Y(men_men_n894_));
  NO3        u872(.A(men_men_n894_), .B(men_men_n892_), .C(men_men_n889_), .Y(men_men_n895_));
  NA3        u873(.A(men_men_n895_), .B(men_men_n888_), .C(men_men_n887_), .Y(men_men_n896_));
  INV        u874(.A(men_men_n859_), .Y(men_men_n897_));
  AOI210     u875(.A0(men_men_n279_), .A1(men_men_n148_), .B0(men_men_n897_), .Y(men_men_n898_));
  NA3        u876(.A(men_men_n39_), .B(men_men_n28_), .C(men_men_n44_), .Y(men_men_n899_));
  NA2        u877(.A(men_men_n833_), .B(men_men_n456_), .Y(men_men_n900_));
  AOI210     u878(.A0(men_men_n899_), .A1(men_men_n148_), .B0(men_men_n900_), .Y(men_men_n901_));
  NO2        u879(.A(men_men_n901_), .B(men_men_n898_), .Y(men_men_n902_));
  NO3        u880(.A(men_men_n820_), .B(men_men_n798_), .C(men_men_n173_), .Y(men_men_n903_));
  AOI220     u881(.A0(men_men_n903_), .A1(i_11_), .B0(men_men_n538_), .B1(men_men_n67_), .Y(men_men_n904_));
  NA2        u882(.A(men_men_n68_), .B(i_13_), .Y(men_men_n905_));
  INV        u883(.A(men_men_n199_), .Y(men_men_n906_));
  OAI220     u884(.A0(men_men_n498_), .A1(men_men_n1005_), .B0(i_12_), .B1(men_men_n585_), .Y(men_men_n907_));
  NA3        u885(.A(men_men_n907_), .B(men_men_n371_), .C(men_men_n906_), .Y(men_men_n908_));
  NA4        u886(.A(men_men_n908_), .B(men_men_n905_), .C(men_men_n904_), .D(men_men_n902_), .Y(men_men_n909_));
  NO2        u887(.A(men_men_n223_), .B(men_men_n85_), .Y(men_men_n910_));
  AOI210     u888(.A0(men_men_n910_), .A1(men_men_n882_), .B0(men_men_n100_), .Y(men_men_n911_));
  AOI220     u889(.A0(men_men_n850_), .A1(men_men_n456_), .B0(men_men_n782_), .B1(men_men_n149_), .Y(men_men_n912_));
  NA2        u890(.A(men_men_n326_), .B(men_men_n159_), .Y(men_men_n913_));
  OA220      u891(.A0(men_men_n913_), .A1(men_men_n912_), .B0(men_men_n911_), .B1(i_5_), .Y(men_men_n914_));
  AOI210     u892(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n158_), .Y(men_men_n915_));
  NA2        u893(.A(men_men_n915_), .B(men_men_n862_), .Y(men_men_n916_));
  NA3        u894(.A(men_men_n582_), .B(men_men_n168_), .C(men_men_n75_), .Y(men_men_n917_));
  NA2        u895(.A(men_men_n917_), .B(men_men_n514_), .Y(men_men_n918_));
  NA3        u896(.A(men_men_n460_), .B(men_men_n455_), .C(men_men_n440_), .Y(men_men_n919_));
  NO2        u897(.A(men_men_n919_), .B(men_men_n918_), .Y(men_men_n920_));
  NA3        u898(.A(men_men_n363_), .B(men_men_n155_), .C(men_men_n154_), .Y(men_men_n921_));
  NA3        u899(.A(men_men_n833_), .B(men_men_n268_), .C(men_men_n211_), .Y(men_men_n922_));
  NA2        u900(.A(men_men_n922_), .B(men_men_n921_), .Y(men_men_n923_));
  NA3        u901(.A(men_men_n363_), .B(men_men_n314_), .C(men_men_n203_), .Y(men_men_n924_));
  INV        u902(.A(men_men_n924_), .Y(men_men_n925_));
  NOi31      u903(.An(men_men_n362_), .B(men_men_n883_), .C(men_men_n220_), .Y(men_men_n926_));
  NO3        u904(.A(men_men_n926_), .B(men_men_n925_), .C(men_men_n923_), .Y(men_men_n927_));
  NA4        u905(.A(men_men_n927_), .B(men_men_n920_), .C(men_men_n916_), .D(men_men_n914_), .Y(men_men_n928_));
  INV        u906(.A(men_men_n584_), .Y(men_men_n929_));
  NO3        u907(.A(men_men_n929_), .B(men_men_n529_), .C(i_3_), .Y(men_men_n930_));
  NO2        u908(.A(men_men_n77_), .B(i_5_), .Y(men_men_n931_));
  NA3        u909(.A(men_men_n783_), .B(men_men_n101_), .C(men_men_n112_), .Y(men_men_n932_));
  INV        u910(.A(men_men_n932_), .Y(men_men_n933_));
  AOI210     u911(.A0(men_men_n933_), .A1(men_men_n931_), .B0(men_men_n930_), .Y(men_men_n934_));
  NA3        u912(.A(men_men_n284_), .B(i_5_), .C(men_men_n176_), .Y(men_men_n935_));
  NO3        u913(.A(men_men_n220_), .B(i_0_), .C(i_12_), .Y(men_men_n936_));
  AOI220     u914(.A0(men_men_n936_), .A1(men_men_n222_), .B0(men_men_n739_), .B1(men_men_n159_), .Y(men_men_n937_));
  AN2        u915(.A(men_men_n820_), .B(men_men_n139_), .Y(men_men_n938_));
  NO4        u916(.A(men_men_n938_), .B(i_12_), .C(men_men_n619_), .D(men_men_n118_), .Y(men_men_n939_));
  NA2        u917(.A(men_men_n939_), .B(men_men_n199_), .Y(men_men_n940_));
  NA3        u918(.A(men_men_n91_), .B(men_men_n542_), .C(i_11_), .Y(men_men_n941_));
  NO2        u919(.A(men_men_n941_), .B(men_men_n141_), .Y(men_men_n942_));
  NA2        u920(.A(men_men_n850_), .B(men_men_n439_), .Y(men_men_n943_));
  INV        u921(.A(men_men_n58_), .Y(men_men_n944_));
  OAI210     u922(.A0(men_men_n944_), .A1(men_men_n935_), .B0(men_men_n943_), .Y(men_men_n945_));
  AOI210     u923(.A0(men_men_n945_), .A1(men_men_n837_), .B0(men_men_n942_), .Y(men_men_n946_));
  NA4        u924(.A(men_men_n946_), .B(men_men_n940_), .C(men_men_n937_), .D(men_men_n934_), .Y(men_men_n947_));
  NO4        u925(.A(men_men_n947_), .B(men_men_n928_), .C(men_men_n909_), .D(men_men_n896_), .Y(men_men_n948_));
  NA2        u926(.A(men_men_n756_), .B(men_men_n37_), .Y(men_men_n949_));
  NA3        u927(.A(men_men_n845_), .B(men_men_n344_), .C(i_5_), .Y(men_men_n950_));
  NA2        u928(.A(men_men_n950_), .B(men_men_n949_), .Y(men_men_n951_));
  NA2        u929(.A(men_men_n951_), .B(men_men_n189_), .Y(men_men_n952_));
  AN2        u930(.A(men_men_n661_), .B(men_men_n345_), .Y(men_men_n953_));
  NA2        u931(.A(men_men_n169_), .B(men_men_n171_), .Y(men_men_n954_));
  AO210      u932(.A0(men_men_n953_), .A1(men_men_n33_), .B0(men_men_n954_), .Y(men_men_n955_));
  OAI210     u933(.A0(men_men_n584_), .A1(men_men_n582_), .B0(men_men_n297_), .Y(men_men_n956_));
  NAi31      u934(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n957_));
  NO2        u935(.A(men_men_n62_), .B(men_men_n957_), .Y(men_men_n958_));
  NO2        u936(.A(men_men_n958_), .B(men_men_n616_), .Y(men_men_n959_));
  NA3        u937(.A(men_men_n959_), .B(men_men_n956_), .C(men_men_n955_), .Y(men_men_n960_));
  NO4        u938(.A(men_men_n214_), .B(men_men_n130_), .C(men_men_n643_), .D(men_men_n37_), .Y(men_men_n961_));
  NO2        u939(.A(men_men_n961_), .B(men_men_n814_), .Y(men_men_n962_));
  OAI210     u940(.A0(men_men_n941_), .A1(men_men_n133_), .B0(men_men_n962_), .Y(men_men_n963_));
  AOI210     u941(.A0(men_men_n960_), .A1(men_men_n48_), .B0(men_men_n963_), .Y(men_men_n964_));
  AOI210     u942(.A0(men_men_n964_), .A1(men_men_n952_), .B0(men_men_n65_), .Y(men_men_n965_));
  NO2        u943(.A(men_men_n998_), .B(men_men_n712_), .Y(men_men_n966_));
  OAI210     u944(.A0(men_men_n72_), .A1(men_men_n52_), .B0(men_men_n99_), .Y(men_men_n967_));
  NA2        u945(.A(men_men_n967_), .B(men_men_n68_), .Y(men_men_n968_));
  AOI210     u946(.A0(men_men_n915_), .A1(men_men_n833_), .B0(men_men_n851_), .Y(men_men_n969_));
  AOI210     u947(.A0(men_men_n969_), .A1(men_men_n968_), .B0(men_men_n643_), .Y(men_men_n970_));
  INV        u948(.A(men_men_n241_), .Y(men_men_n971_));
  AOI220     u949(.A0(men_men_n971_), .A1(men_men_n68_), .B0(men_men_n321_), .B1(men_men_n234_), .Y(men_men_n972_));
  NO2        u950(.A(men_men_n972_), .B(men_men_n218_), .Y(men_men_n973_));
  NA3        u951(.A(men_men_n89_), .B(men_men_n286_), .C(men_men_n31_), .Y(men_men_n974_));
  INV        u952(.A(men_men_n974_), .Y(men_men_n975_));
  NO3        u953(.A(men_men_n975_), .B(men_men_n973_), .C(men_men_n970_), .Y(men_men_n976_));
  OAI210     u954(.A0(men_men_n247_), .A1(men_men_n144_), .B0(men_men_n80_), .Y(men_men_n977_));
  NA3        u955(.A(men_men_n713_), .B(men_men_n268_), .C(men_men_n72_), .Y(men_men_n978_));
  AOI210     u956(.A0(men_men_n978_), .A1(men_men_n977_), .B0(i_11_), .Y(men_men_n979_));
  NA2        u957(.A(men_men_n577_), .B(men_men_n196_), .Y(men_men_n980_));
  NA2        u958(.A(men_men_n980_), .B(men_men_n189_), .Y(men_men_n981_));
  NA2        u959(.A(men_men_n150_), .B(i_5_), .Y(men_men_n982_));
  AOI210     u960(.A0(men_men_n981_), .A1(men_men_n724_), .B0(men_men_n982_), .Y(men_men_n983_));
  NO3        u961(.A(men_men_n55_), .B(men_men_n54_), .C(i_4_), .Y(men_men_n984_));
  OAI210     u962(.A0(men_men_n855_), .A1(men_men_n286_), .B0(men_men_n984_), .Y(men_men_n985_));
  NO2        u963(.A(men_men_n985_), .B(men_men_n684_), .Y(men_men_n986_));
  NO4        u964(.A(men_men_n874_), .B(men_men_n445_), .C(men_men_n231_), .D(men_men_n230_), .Y(men_men_n987_));
  NO2        u965(.A(men_men_n987_), .B(men_men_n533_), .Y(men_men_n988_));
  INV        u966(.A(men_men_n338_), .Y(men_men_n989_));
  AOI210     u967(.A0(men_men_n989_), .A1(men_men_n988_), .B0(men_men_n40_), .Y(men_men_n990_));
  NO4        u968(.A(men_men_n990_), .B(men_men_n986_), .C(men_men_n983_), .D(men_men_n979_), .Y(men_men_n991_));
  OAI210     u969(.A0(men_men_n976_), .A1(i_4_), .B0(men_men_n991_), .Y(men_men_n992_));
  NO3        u970(.A(men_men_n992_), .B(men_men_n966_), .C(men_men_n965_), .Y(men_men_n993_));
  NA4        u971(.A(men_men_n993_), .B(men_men_n948_), .C(men_men_n881_), .D(men_men_n802_), .Y(men4));
  INV        u972(.A(i_2_), .Y(men_men_n997_));
  INV        u973(.A(men_men_n536_), .Y(men_men_n998_));
  INV        u974(.A(i_3_), .Y(men_men_n999_));
  INV        u975(.A(men_men_n307_), .Y(men_men_n1000_));
  INV        u976(.A(i_0_), .Y(men_men_n1001_));
  INV        u977(.A(i_4_), .Y(men_men_n1002_));
  INV        u978(.A(i_9_), .Y(men_men_n1003_));
  INV        u979(.A(i_10_), .Y(men_men_n1004_));
  INV        u980(.A(i_6_), .Y(men_men_n1005_));
  INV        u981(.A(i_1_), .Y(men_men_n1006_));
  INV        u982(.A(men_men_n357_), .Y(men_men_n1007_));
  INV        u983(.A(i_10_), .Y(men_men_n1008_));
  INV        u984(.A(i_7_), .Y(men_men_n1009_));
  INV        u985(.A(i_5_), .Y(men_men_n1010_));
  INV        u986(.A(men_men_n145_), .Y(men_men_n1011_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule