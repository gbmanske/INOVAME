//Benchmark atmr_9sym_175_0.0625

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  NA2        o002(.A(i_4_), .B(ori_ori_n12_), .Y(ori_ori_n13_));
  INV        o003(.A(i_5_), .Y(ori_ori_n14_));
  NOi21      o004(.An(i_3_), .B(i_7_), .Y(ori_ori_n15_));
  NA3        o005(.A(ori_ori_n15_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n16_));
  INV        o006(.A(i_0_), .Y(ori_ori_n17_));
  NOi21      o007(.An(i_1_), .B(i_3_), .Y(ori_ori_n18_));
  NA2        o008(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  AOI210     o009(.A0(ori_ori_n19_), .A1(ori_ori_n16_), .B0(ori_ori_n13_), .Y(ori_ori_n20_));
  INV        o010(.A(i_4_), .Y(ori_ori_n21_));
  NA2        o011(.A(i_0_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  INV        o012(.A(i_7_), .Y(ori_ori_n23_));
  NA3        o013(.A(i_6_), .B(i_5_), .C(ori_ori_n23_), .Y(ori_ori_n24_));
  AOI220     o014(.A0(i_1_), .A1(i_2_), .B0(i_8_), .B1(i_5_), .Y(ori_ori_n25_));
  AOI210     o015(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n22_), .Y(ori_ori_n26_));
  AOI210     o016(.A0(ori_ori_n26_), .A1(ori_ori_n11_), .B0(ori_ori_n20_), .Y(ori_ori_n27_));
  NA2        o017(.A(i_0_), .B(ori_ori_n14_), .Y(ori_ori_n28_));
  NA2        o018(.A(ori_ori_n17_), .B(i_5_), .Y(ori_ori_n29_));
  NO2        o019(.A(i_2_), .B(i_4_), .Y(ori_ori_n30_));
  NA3        o020(.A(ori_ori_n30_), .B(i_6_), .C(i_8_), .Y(ori_ori_n31_));
  AOI210     o021(.A0(ori_ori_n29_), .A1(ori_ori_n28_), .B0(ori_ori_n31_), .Y(ori_ori_n32_));
  INV        o022(.A(i_2_), .Y(ori_ori_n33_));
  NOi21      o023(.An(i_5_), .B(i_0_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_6_), .B(i_8_), .Y(ori_ori_n35_));
  NOi21      o025(.An(i_5_), .B(i_6_), .Y(ori_ori_n36_));
  AOI220     o026(.A0(ori_ori_n36_), .A1(i_7_), .B0(ori_ori_n35_), .B1(ori_ori_n34_), .Y(ori_ori_n37_));
  NO3        o027(.A(ori_ori_n37_), .B(ori_ori_n33_), .C(i_4_), .Y(ori_ori_n38_));
  NOi21      o028(.An(i_0_), .B(i_4_), .Y(ori_ori_n39_));
  INV        o029(.A(i_1_), .Y(ori_ori_n40_));
  NOi21      o030(.An(i_3_), .B(i_0_), .Y(ori_ori_n41_));
  NA2        o031(.A(ori_ori_n41_), .B(ori_ori_n40_), .Y(ori_ori_n42_));
  NO2        o032(.A(ori_ori_n24_), .B(ori_ori_n42_), .Y(ori_ori_n43_));
  NO3        o033(.A(ori_ori_n43_), .B(ori_ori_n38_), .C(ori_ori_n32_), .Y(ori_ori_n44_));
  NA2        o034(.A(i_1_), .B(ori_ori_n11_), .Y(ori_ori_n45_));
  NOi21      o035(.An(i_4_), .B(i_0_), .Y(ori_ori_n46_));
  NA2        o036(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n47_));
  NOi21      o037(.An(i_2_), .B(i_8_), .Y(ori_ori_n48_));
  NOi31      o038(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n49_));
  NA2        o039(.A(ori_ori_n49_), .B(i_0_), .Y(ori_ori_n50_));
  NOi21      o040(.An(i_4_), .B(i_3_), .Y(ori_ori_n51_));
  NOi21      o041(.An(i_1_), .B(i_4_), .Y(ori_ori_n52_));
  NA2        o042(.A(ori_ori_n51_), .B(ori_ori_n48_), .Y(ori_ori_n53_));
  NA2        o043(.A(ori_ori_n53_), .B(ori_ori_n50_), .Y(ori_ori_n54_));
  AN2        o044(.A(i_8_), .B(i_7_), .Y(ori_ori_n55_));
  INV        o045(.A(ori_ori_n55_), .Y(ori_ori_n56_));
  NOi21      o046(.An(i_8_), .B(i_7_), .Y(ori_ori_n57_));
  NA2        o047(.A(ori_ori_n57_), .B(ori_ori_n51_), .Y(ori_ori_n58_));
  OAI210     o048(.A0(ori_ori_n56_), .A1(ori_ori_n47_), .B0(ori_ori_n58_), .Y(ori_ori_n59_));
  AOI220     o049(.A0(ori_ori_n59_), .A1(ori_ori_n33_), .B0(ori_ori_n54_), .B1(ori_ori_n36_), .Y(ori_ori_n60_));
  NA3        o050(.A(ori_ori_n60_), .B(ori_ori_n44_), .C(ori_ori_n27_), .Y(ori_ori_n61_));
  INV        o051(.A(i_8_), .Y(ori_ori_n62_));
  NO3        o052(.A(ori_ori_n62_), .B(ori_ori_n13_), .C(i_1_), .Y(ori_ori_n63_));
  NOi21      o053(.An(i_1_), .B(i_2_), .Y(ori_ori_n64_));
  NA2        o054(.A(ori_ori_n63_), .B(ori_ori_n14_), .Y(ori_ori_n65_));
  NA3        o055(.A(ori_ori_n57_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n66_));
  NOi32      o056(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(ori_ori_n67_));
  NA2        o057(.A(ori_ori_n67_), .B(i_3_), .Y(ori_ori_n68_));
  NA2        o058(.A(ori_ori_n18_), .B(i_6_), .Y(ori_ori_n69_));
  NA2        o059(.A(ori_ori_n69_), .B(ori_ori_n68_), .Y(ori_ori_n70_));
  INV        o060(.A(i_0_), .Y(ori_ori_n71_));
  NA2        o061(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n72_));
  NA2        o062(.A(ori_ori_n72_), .B(ori_ori_n65_), .Y(ori_ori_n73_));
  NAi21      o063(.An(i_3_), .B(i_6_), .Y(ori_ori_n74_));
  NA2        o064(.A(ori_ori_n35_), .B(ori_ori_n34_), .Y(ori_ori_n75_));
  NOi21      o065(.An(i_7_), .B(i_8_), .Y(ori_ori_n76_));
  OAI210     o066(.A0(i_5_), .A1(ori_ori_n11_), .B0(ori_ori_n75_), .Y(ori_ori_n77_));
  NA2        o067(.A(ori_ori_n77_), .B(ori_ori_n64_), .Y(ori_ori_n78_));
  NA3        o068(.A(i_8_), .B(i_2_), .C(ori_ori_n14_), .Y(ori_ori_n79_));
  AOI210     o069(.A0(ori_ori_n22_), .A1(ori_ori_n45_), .B0(ori_ori_n79_), .Y(ori_ori_n80_));
  INV        o070(.A(ori_ori_n80_), .Y(ori_ori_n81_));
  NA3        o071(.A(ori_ori_n57_), .B(ori_ori_n33_), .C(i_3_), .Y(ori_ori_n82_));
  NA2        o072(.A(ori_ori_n40_), .B(i_6_), .Y(ori_ori_n83_));
  NO2        o073(.A(ori_ori_n83_), .B(ori_ori_n82_), .Y(ori_ori_n84_));
  NOi21      o074(.An(i_2_), .B(i_1_), .Y(ori_ori_n85_));
  AN3        o075(.A(ori_ori_n76_), .B(ori_ori_n85_), .C(ori_ori_n46_), .Y(ori_ori_n86_));
  NAi21      o076(.An(i_6_), .B(i_0_), .Y(ori_ori_n87_));
  NA3        o077(.A(ori_ori_n52_), .B(i_5_), .C(ori_ori_n23_), .Y(ori_ori_n88_));
  NOi21      o078(.An(i_4_), .B(i_6_), .Y(ori_ori_n89_));
  BUFFER     o079(.A(i_5_), .Y(ori_ori_n90_));
  NA2        o080(.A(ori_ori_n64_), .B(ori_ori_n89_), .Y(ori_ori_n91_));
  NA2        o081(.A(ori_ori_n88_), .B(ori_ori_n91_), .Y(ori_ori_n92_));
  NA2        o082(.A(ori_ori_n64_), .B(ori_ori_n35_), .Y(ori_ori_n93_));
  NO3        o083(.A(ori_ori_n92_), .B(ori_ori_n86_), .C(ori_ori_n84_), .Y(ori_ori_n94_));
  NA2        o084(.A(ori_ori_n57_), .B(ori_ori_n12_), .Y(ori_ori_n95_));
  NA2        o085(.A(ori_ori_n35_), .B(ori_ori_n14_), .Y(ori_ori_n96_));
  NOi21      o086(.An(i_3_), .B(i_1_), .Y(ori_ori_n97_));
  NA2        o087(.A(ori_ori_n97_), .B(i_4_), .Y(ori_ori_n98_));
  AOI210     o088(.A0(ori_ori_n96_), .A1(ori_ori_n95_), .B0(ori_ori_n98_), .Y(ori_ori_n99_));
  NOi31      o089(.An(ori_ori_n41_), .B(i_5_), .C(ori_ori_n33_), .Y(ori_ori_n100_));
  NO2        o090(.A(ori_ori_n100_), .B(ori_ori_n99_), .Y(ori_ori_n101_));
  NA4        o091(.A(ori_ori_n101_), .B(ori_ori_n94_), .C(ori_ori_n81_), .D(ori_ori_n78_), .Y(ori_ori_n102_));
  NOi31      o092(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n103_));
  NA3        o093(.A(ori_ori_n35_), .B(i_2_), .C(ori_ori_n14_), .Y(ori_ori_n104_));
  NA2        o094(.A(ori_ori_n104_), .B(ori_ori_n93_), .Y(ori_ori_n105_));
  NA2        o095(.A(ori_ori_n105_), .B(ori_ori_n39_), .Y(ori_ori_n106_));
  NA2        o096(.A(ori_ori_n51_), .B(i_7_), .Y(ori_ori_n107_));
  AOI210     o097(.A0(ori_ori_n107_), .A1(ori_ori_n66_), .B0(ori_ori_n29_), .Y(ori_ori_n108_));
  NA4        o098(.A(ori_ori_n55_), .B(ori_ori_n85_), .C(ori_ori_n17_), .D(ori_ori_n12_), .Y(ori_ori_n109_));
  NAi31      o099(.An(ori_ori_n87_), .B(ori_ori_n76_), .C(ori_ori_n85_), .Y(ori_ori_n110_));
  NA3        o100(.A(ori_ori_n57_), .B(ori_ori_n49_), .C(i_6_), .Y(ori_ori_n111_));
  NA3        o101(.A(ori_ori_n111_), .B(ori_ori_n110_), .C(ori_ori_n109_), .Y(ori_ori_n112_));
  NOi21      o102(.An(i_0_), .B(i_2_), .Y(ori_ori_n113_));
  NA3        o103(.A(ori_ori_n113_), .B(i_7_), .C(ori_ori_n89_), .Y(ori_ori_n114_));
  NOi32      o104(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n115_));
  NA2        o105(.A(ori_ori_n115_), .B(ori_ori_n103_), .Y(ori_ori_n116_));
  NA3        o106(.A(ori_ori_n113_), .B(ori_ori_n51_), .C(ori_ori_n35_), .Y(ori_ori_n117_));
  NA3        o107(.A(ori_ori_n117_), .B(ori_ori_n116_), .C(ori_ori_n114_), .Y(ori_ori_n118_));
  NA4        o108(.A(ori_ori_n49_), .B(i_6_), .C(ori_ori_n14_), .D(i_7_), .Y(ori_ori_n119_));
  NA2        o109(.A(ori_ori_n52_), .B(ori_ori_n36_), .Y(ori_ori_n120_));
  NA2        o110(.A(ori_ori_n120_), .B(ori_ori_n119_), .Y(ori_ori_n121_));
  NO4        o111(.A(ori_ori_n121_), .B(ori_ori_n118_), .C(ori_ori_n112_), .D(ori_ori_n108_), .Y(ori_ori_n122_));
  INV        o112(.A(i_2_), .Y(ori_ori_n123_));
  AOI220     o113(.A0(ori_ori_n123_), .A1(ori_ori_n76_), .B0(ori_ori_n55_), .B1(ori_ori_n30_), .Y(ori_ori_n124_));
  NO2        o114(.A(ori_ori_n124_), .B(ori_ori_n83_), .Y(ori_ori_n125_));
  NO4        o115(.A(i_2_), .B(ori_ori_n21_), .C(ori_ori_n11_), .D(ori_ori_n14_), .Y(ori_ori_n126_));
  NA2        o116(.A(i_2_), .B(i_4_), .Y(ori_ori_n127_));
  AOI210     o117(.A0(ori_ori_n87_), .A1(ori_ori_n74_), .B0(ori_ori_n127_), .Y(ori_ori_n128_));
  NO2        o118(.A(i_8_), .B(i_7_), .Y(ori_ori_n129_));
  OA210      o119(.A0(ori_ori_n128_), .A1(ori_ori_n126_), .B0(ori_ori_n129_), .Y(ori_ori_n130_));
  NA2        o120(.A(ori_ori_n97_), .B(i_0_), .Y(ori_ori_n131_));
  NO2        o121(.A(ori_ori_n131_), .B(i_4_), .Y(ori_ori_n132_));
  NO3        o122(.A(ori_ori_n132_), .B(ori_ori_n130_), .C(ori_ori_n125_), .Y(ori_ori_n133_));
  NA2        o123(.A(ori_ori_n76_), .B(ori_ori_n12_), .Y(ori_ori_n134_));
  NA2        o124(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n135_));
  NA2        o125(.A(ori_ori_n46_), .B(i_3_), .Y(ori_ori_n136_));
  AOI210     o126(.A0(ori_ori_n136_), .A1(ori_ori_n135_), .B0(ori_ori_n134_), .Y(ori_ori_n137_));
  NO2        o127(.A(ori_ori_n82_), .B(ori_ori_n29_), .Y(ori_ori_n138_));
  NA4        o128(.A(ori_ori_n90_), .B(ori_ori_n55_), .C(ori_ori_n40_), .D(ori_ori_n21_), .Y(ori_ori_n139_));
  NA3        o129(.A(ori_ori_n48_), .B(ori_ori_n34_), .C(ori_ori_n15_), .Y(ori_ori_n140_));
  NOi31      o130(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n141_));
  OAI210     o131(.A0(ori_ori_n115_), .A1(ori_ori_n67_), .B0(ori_ori_n141_), .Y(ori_ori_n142_));
  NA3        o132(.A(ori_ori_n142_), .B(ori_ori_n140_), .C(ori_ori_n139_), .Y(ori_ori_n143_));
  NO3        o133(.A(ori_ori_n143_), .B(ori_ori_n138_), .C(ori_ori_n137_), .Y(ori_ori_n144_));
  NA4        o134(.A(ori_ori_n144_), .B(ori_ori_n133_), .C(ori_ori_n122_), .D(ori_ori_n106_), .Y(ori_ori_n145_));
  OR4        o135(.A(ori_ori_n145_), .B(ori_ori_n102_), .C(ori_ori_n73_), .D(ori_ori_n61_), .Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  INV        m002(.A(i_5_), .Y(mai_mai_n13_));
  NOi21      m003(.An(i_3_), .B(i_7_), .Y(mai_mai_n14_));
  INV        m004(.A(i_0_), .Y(mai_mai_n15_));
  NOi21      m005(.An(i_1_), .B(i_3_), .Y(mai_mai_n16_));
  INV        m006(.A(i_4_), .Y(mai_mai_n17_));
  NA2        m007(.A(i_0_), .B(mai_mai_n17_), .Y(mai_mai_n18_));
  INV        m008(.A(i_7_), .Y(mai_mai_n19_));
  NA3        m009(.A(i_6_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n20_));
  NOi21      m010(.An(i_8_), .B(i_6_), .Y(mai_mai_n21_));
  NOi21      m011(.An(i_1_), .B(i_8_), .Y(mai_mai_n22_));
  AOI220     m012(.A0(mai_mai_n22_), .A1(i_2_), .B0(mai_mai_n21_), .B1(i_5_), .Y(mai_mai_n23_));
  AOI210     m013(.A0(mai_mai_n23_), .A1(mai_mai_n20_), .B0(mai_mai_n18_), .Y(mai_mai_n24_));
  NA2        m014(.A(mai_mai_n24_), .B(mai_mai_n11_), .Y(mai_mai_n25_));
  NA2        m015(.A(i_0_), .B(mai_mai_n13_), .Y(mai_mai_n26_));
  NA2        m016(.A(mai_mai_n15_), .B(i_5_), .Y(mai_mai_n27_));
  NO2        m017(.A(i_2_), .B(i_4_), .Y(mai_mai_n28_));
  NA3        m018(.A(mai_mai_n28_), .B(i_6_), .C(i_8_), .Y(mai_mai_n29_));
  AOI210     m019(.A0(mai_mai_n27_), .A1(mai_mai_n26_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  INV        m020(.A(i_2_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_6_), .B(i_8_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_7_), .B(i_1_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_5_), .B(i_6_), .Y(mai_mai_n34_));
  AOI220     m024(.A0(mai_mai_n34_), .A1(mai_mai_n33_), .B0(mai_mai_n32_), .B1(i_5_), .Y(mai_mai_n35_));
  NO3        m025(.A(mai_mai_n35_), .B(mai_mai_n31_), .C(i_4_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_0_), .B(i_4_), .Y(mai_mai_n37_));
  XO2        m027(.A(i_1_), .B(i_3_), .Y(mai_mai_n38_));
  NOi21      m028(.An(i_7_), .B(i_5_), .Y(mai_mai_n39_));
  AN3        m029(.A(mai_mai_n39_), .B(mai_mai_n38_), .C(mai_mai_n37_), .Y(mai_mai_n40_));
  INV        m030(.A(i_1_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_3_), .B(i_0_), .Y(mai_mai_n42_));
  NA2        m032(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA3        m033(.A(i_6_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n44_));
  AOI210     m034(.A0(mai_mai_n44_), .A1(mai_mai_n20_), .B0(mai_mai_n43_), .Y(mai_mai_n45_));
  NO4        m035(.A(mai_mai_n45_), .B(mai_mai_n40_), .C(mai_mai_n36_), .D(mai_mai_n30_), .Y(mai_mai_n46_));
  INV        m036(.A(i_8_), .Y(mai_mai_n47_));
  NA2        m037(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n48_));
  NO4        m038(.A(mai_mai_n48_), .B(mai_mai_n26_), .C(i_2_), .D(mai_mai_n47_), .Y(mai_mai_n49_));
  NOi21      m039(.An(i_4_), .B(i_0_), .Y(mai_mai_n50_));
  AOI210     m040(.A0(mai_mai_n50_), .A1(mai_mai_n21_), .B0(mai_mai_n14_), .Y(mai_mai_n51_));
  NA2        m041(.A(i_1_), .B(mai_mai_n13_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_2_), .B(i_8_), .Y(mai_mai_n53_));
  NO3        m043(.A(mai_mai_n53_), .B(mai_mai_n50_), .C(mai_mai_n37_), .Y(mai_mai_n54_));
  NO3        m044(.A(mai_mai_n54_), .B(mai_mai_n52_), .C(mai_mai_n51_), .Y(mai_mai_n55_));
  NO2        m045(.A(mai_mai_n55_), .B(mai_mai_n49_), .Y(mai_mai_n56_));
  NOi31      m046(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n57_));
  NA2        m047(.A(mai_mai_n57_), .B(i_0_), .Y(mai_mai_n58_));
  NOi21      m048(.An(i_4_), .B(i_3_), .Y(mai_mai_n59_));
  NOi21      m049(.An(i_1_), .B(i_4_), .Y(mai_mai_n60_));
  OAI210     m050(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n53_), .Y(mai_mai_n61_));
  NA2        m051(.A(mai_mai_n61_), .B(mai_mai_n58_), .Y(mai_mai_n62_));
  AN2        m052(.A(i_8_), .B(i_7_), .Y(mai_mai_n63_));
  NA2        m053(.A(mai_mai_n63_), .B(mai_mai_n12_), .Y(mai_mai_n64_));
  NOi21      m054(.An(i_8_), .B(i_7_), .Y(mai_mai_n65_));
  NA3        m055(.A(mai_mai_n65_), .B(mai_mai_n59_), .C(i_6_), .Y(mai_mai_n66_));
  OAI210     m056(.A0(mai_mai_n64_), .A1(mai_mai_n52_), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  AOI220     m057(.A0(mai_mai_n67_), .A1(mai_mai_n31_), .B0(mai_mai_n62_), .B1(mai_mai_n34_), .Y(mai_mai_n68_));
  NA4        m058(.A(mai_mai_n68_), .B(mai_mai_n56_), .C(mai_mai_n46_), .D(mai_mai_n25_), .Y(mai_mai_n69_));
  NA2        m059(.A(i_8_), .B(mai_mai_n19_), .Y(mai_mai_n70_));
  AOI220     m060(.A0(mai_mai_n42_), .A1(i_1_), .B0(mai_mai_n38_), .B1(i_2_), .Y(mai_mai_n71_));
  NOi21      m061(.An(i_1_), .B(i_2_), .Y(mai_mai_n72_));
  NA3        m062(.A(mai_mai_n72_), .B(mai_mai_n50_), .C(i_6_), .Y(mai_mai_n73_));
  OAI210     m063(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n73_), .Y(mai_mai_n74_));
  NA2        m064(.A(mai_mai_n74_), .B(mai_mai_n13_), .Y(mai_mai_n75_));
  NA3        m065(.A(mai_mai_n65_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n76_));
  NA3        m066(.A(mai_mai_n22_), .B(i_0_), .C(mai_mai_n13_), .Y(mai_mai_n77_));
  NA2        m067(.A(mai_mai_n77_), .B(mai_mai_n76_), .Y(mai_mai_n78_));
  NOi32      m068(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n79_));
  NA2        m069(.A(mai_mai_n79_), .B(i_3_), .Y(mai_mai_n80_));
  NA3        m070(.A(mai_mai_n16_), .B(i_2_), .C(i_6_), .Y(mai_mai_n81_));
  NA2        m071(.A(mai_mai_n81_), .B(mai_mai_n80_), .Y(mai_mai_n82_));
  NO2        m072(.A(i_0_), .B(i_4_), .Y(mai_mai_n83_));
  AOI220     m073(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n78_), .B1(mai_mai_n59_), .Y(mai_mai_n84_));
  NA2        m074(.A(mai_mai_n84_), .B(mai_mai_n75_), .Y(mai_mai_n85_));
  NO3        m075(.A(i_3_), .B(i_0_), .C(mai_mai_n47_), .Y(mai_mai_n86_));
  NA2        m076(.A(mai_mai_n32_), .B(i_5_), .Y(mai_mai_n87_));
  NOi21      m077(.An(i_7_), .B(i_8_), .Y(mai_mai_n88_));
  INV        m078(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  OAI210     m079(.A0(mai_mai_n89_), .A1(mai_mai_n11_), .B0(mai_mai_n87_), .Y(mai_mai_n90_));
  OAI210     m080(.A0(mai_mai_n90_), .A1(mai_mai_n86_), .B0(mai_mai_n72_), .Y(mai_mai_n91_));
  NA3        m081(.A(mai_mai_n21_), .B(i_2_), .C(mai_mai_n13_), .Y(mai_mai_n92_));
  AOI210     m082(.A0(mai_mai_n18_), .A1(mai_mai_n48_), .B0(mai_mai_n92_), .Y(mai_mai_n93_));
  AOI220     m083(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n16_), .B1(mai_mai_n31_), .Y(mai_mai_n94_));
  NA3        m084(.A(mai_mai_n17_), .B(i_5_), .C(i_7_), .Y(mai_mai_n95_));
  NO2        m085(.A(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  NO2        m086(.A(mai_mai_n96_), .B(mai_mai_n93_), .Y(mai_mai_n97_));
  NA3        m087(.A(mai_mai_n65_), .B(mai_mai_n31_), .C(i_3_), .Y(mai_mai_n98_));
  NA2        m088(.A(mai_mai_n41_), .B(i_6_), .Y(mai_mai_n99_));
  AOI210     m089(.A0(mai_mai_n99_), .A1(mai_mai_n18_), .B0(mai_mai_n98_), .Y(mai_mai_n100_));
  NOi21      m090(.An(i_4_), .B(i_6_), .Y(mai_mai_n101_));
  NOi21      m091(.An(i_5_), .B(i_3_), .Y(mai_mai_n102_));
  NA3        m092(.A(mai_mai_n102_), .B(mai_mai_n72_), .C(mai_mai_n101_), .Y(mai_mai_n103_));
  INV        m093(.A(mai_mai_n103_), .Y(mai_mai_n104_));
  NO2        m094(.A(mai_mai_n104_), .B(mai_mai_n100_), .Y(mai_mai_n105_));
  NOi21      m095(.An(i_6_), .B(i_1_), .Y(mai_mai_n106_));
  AOI220     m096(.A0(mai_mai_n106_), .A1(i_7_), .B0(mai_mai_n21_), .B1(i_5_), .Y(mai_mai_n107_));
  NOi31      m097(.An(mai_mai_n50_), .B(mai_mai_n107_), .C(i_2_), .Y(mai_mai_n108_));
  NOi21      m098(.An(i_3_), .B(i_1_), .Y(mai_mai_n109_));
  NA2        m099(.A(mai_mai_n109_), .B(i_4_), .Y(mai_mai_n110_));
  NO2        m100(.A(i_6_), .B(mai_mai_n110_), .Y(mai_mai_n111_));
  NO2        m101(.A(mai_mai_n111_), .B(mai_mai_n108_), .Y(mai_mai_n112_));
  NA4        m102(.A(mai_mai_n112_), .B(mai_mai_n105_), .C(mai_mai_n97_), .D(mai_mai_n91_), .Y(mai_mai_n113_));
  NOi31      m103(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n114_));
  INV        m104(.A(mai_mai_n114_), .Y(mai_mai_n115_));
  NA2        m105(.A(mai_mai_n32_), .B(mai_mai_n13_), .Y(mai_mai_n116_));
  NA2        m106(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NA2        m107(.A(mai_mai_n117_), .B(mai_mai_n37_), .Y(mai_mai_n118_));
  NA2        m108(.A(mai_mai_n59_), .B(mai_mai_n33_), .Y(mai_mai_n119_));
  AOI210     m109(.A0(mai_mai_n119_), .A1(mai_mai_n76_), .B0(mai_mai_n27_), .Y(mai_mai_n120_));
  NA3        m110(.A(mai_mai_n65_), .B(mai_mai_n57_), .C(i_6_), .Y(mai_mai_n121_));
  INV        m111(.A(mai_mai_n121_), .Y(mai_mai_n122_));
  NA3        m112(.A(mai_mai_n57_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n123_));
  NA4        m113(.A(mai_mai_n60_), .B(mai_mai_n34_), .C(mai_mai_n15_), .D(i_8_), .Y(mai_mai_n124_));
  NA2        m114(.A(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n125_));
  NO3        m115(.A(mai_mai_n125_), .B(mai_mai_n122_), .C(mai_mai_n120_), .Y(mai_mai_n126_));
  BUFFER     m116(.A(i_5_), .Y(mai_mai_n127_));
  AOI220     m117(.A0(mai_mai_n127_), .A1(mai_mai_n88_), .B0(mai_mai_n63_), .B1(mai_mai_n28_), .Y(mai_mai_n128_));
  NO2        m118(.A(mai_mai_n128_), .B(mai_mai_n99_), .Y(mai_mai_n129_));
  NO3        m119(.A(i_2_), .B(mai_mai_n17_), .C(mai_mai_n11_), .Y(mai_mai_n130_));
  NA2        m120(.A(i_2_), .B(i_4_), .Y(mai_mai_n131_));
  INV        m121(.A(mai_mai_n131_), .Y(mai_mai_n132_));
  NO2        m122(.A(i_8_), .B(i_7_), .Y(mai_mai_n133_));
  OA210      m123(.A0(mai_mai_n132_), .A1(mai_mai_n130_), .B0(mai_mai_n133_), .Y(mai_mai_n134_));
  NA4        m124(.A(mai_mai_n109_), .B(i_0_), .C(i_5_), .D(mai_mai_n19_), .Y(mai_mai_n135_));
  NO2        m125(.A(mai_mai_n135_), .B(i_4_), .Y(mai_mai_n136_));
  NO3        m126(.A(mai_mai_n136_), .B(mai_mai_n134_), .C(mai_mai_n129_), .Y(mai_mai_n137_));
  INV        m127(.A(mai_mai_n88_), .Y(mai_mai_n138_));
  NA2        m128(.A(i_2_), .B(mai_mai_n13_), .Y(mai_mai_n139_));
  NO2        m129(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n140_));
  NA3        m130(.A(i_0_), .B(mai_mai_n65_), .C(mai_mai_n101_), .Y(mai_mai_n141_));
  OAI210     m131(.A0(mai_mai_n98_), .A1(mai_mai_n27_), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  NA4        m132(.A(mai_mai_n102_), .B(mai_mai_n63_), .C(mai_mai_n41_), .D(mai_mai_n17_), .Y(mai_mai_n143_));
  NOi31      m133(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n144_));
  OAI210     m134(.A0(i_4_), .A1(mai_mai_n79_), .B0(mai_mai_n144_), .Y(mai_mai_n145_));
  NA2        m135(.A(mai_mai_n145_), .B(mai_mai_n143_), .Y(mai_mai_n146_));
  NO3        m136(.A(mai_mai_n146_), .B(mai_mai_n142_), .C(mai_mai_n140_), .Y(mai_mai_n147_));
  NA4        m137(.A(mai_mai_n147_), .B(mai_mai_n137_), .C(mai_mai_n126_), .D(mai_mai_n118_), .Y(mai_mai_n148_));
  OR4        m138(.A(mai_mai_n148_), .B(mai_mai_n113_), .C(mai_mai_n85_), .D(mai_mai_n69_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  INV        u011(.A(i_7_), .Y(men_men_n22_));
  NA3        u012(.A(i_6_), .B(i_5_), .C(men_men_n22_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  NOi21      u014(.An(i_1_), .B(i_8_), .Y(men_men_n25_));
  AOI220     u015(.A0(men_men_n25_), .A1(i_2_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n26_));
  AOI210     u016(.A0(men_men_n26_), .A1(men_men_n23_), .B0(i_4_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n28_));
  NA2        u018(.A(i_0_), .B(men_men_n14_), .Y(men_men_n29_));
  INV        u019(.A(i_2_), .Y(men_men_n30_));
  NOi21      u020(.An(i_5_), .B(i_0_), .Y(men_men_n31_));
  NOi21      u021(.An(i_6_), .B(i_8_), .Y(men_men_n32_));
  NOi21      u022(.An(i_7_), .B(i_1_), .Y(men_men_n33_));
  NOi21      u023(.An(i_5_), .B(i_6_), .Y(men_men_n34_));
  AOI220     u024(.A0(men_men_n34_), .A1(men_men_n33_), .B0(men_men_n32_), .B1(men_men_n31_), .Y(men_men_n35_));
  NO3        u025(.A(men_men_n35_), .B(men_men_n30_), .C(i_4_), .Y(men_men_n36_));
  NOi21      u026(.An(i_0_), .B(i_4_), .Y(men_men_n37_));
  XO2        u027(.A(i_1_), .B(i_3_), .Y(men_men_n38_));
  NOi21      u028(.An(i_7_), .B(i_5_), .Y(men_men_n39_));
  AN3        u029(.A(men_men_n39_), .B(men_men_n38_), .C(men_men_n37_), .Y(men_men_n40_));
  INV        u030(.A(i_1_), .Y(men_men_n41_));
  NOi21      u031(.An(i_3_), .B(i_0_), .Y(men_men_n42_));
  NO2        u032(.A(men_men_n23_), .B(i_0_), .Y(men_men_n43_));
  NO3        u033(.A(men_men_n43_), .B(men_men_n40_), .C(men_men_n36_), .Y(men_men_n44_));
  INV        u034(.A(i_8_), .Y(men_men_n45_));
  NO4        u035(.A(i_3_), .B(men_men_n29_), .C(i_2_), .D(men_men_n45_), .Y(men_men_n46_));
  NOi21      u036(.An(i_4_), .B(i_0_), .Y(men_men_n47_));
  AOI210     u037(.A0(men_men_n47_), .A1(men_men_n24_), .B0(men_men_n15_), .Y(men_men_n48_));
  NA2        u038(.A(i_1_), .B(men_men_n14_), .Y(men_men_n49_));
  NOi21      u039(.An(i_2_), .B(i_8_), .Y(men_men_n50_));
  NO3        u040(.A(men_men_n50_), .B(men_men_n47_), .C(men_men_n37_), .Y(men_men_n51_));
  NO3        u041(.A(men_men_n51_), .B(men_men_n49_), .C(men_men_n48_), .Y(men_men_n52_));
  NO2        u042(.A(men_men_n52_), .B(men_men_n46_), .Y(men_men_n53_));
  NOi31      u043(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n54_));
  NOi21      u044(.An(i_4_), .B(i_3_), .Y(men_men_n55_));
  NOi21      u045(.An(i_1_), .B(i_4_), .Y(men_men_n56_));
  AN2        u046(.A(i_8_), .B(i_7_), .Y(men_men_n57_));
  NA2        u047(.A(men_men_n57_), .B(men_men_n12_), .Y(men_men_n58_));
  NOi21      u048(.An(i_8_), .B(i_7_), .Y(men_men_n59_));
  NA3        u049(.A(men_men_n59_), .B(men_men_n55_), .C(i_6_), .Y(men_men_n60_));
  OAI210     u050(.A0(men_men_n58_), .A1(men_men_n49_), .B0(men_men_n60_), .Y(men_men_n61_));
  AOI220     u051(.A0(men_men_n61_), .A1(men_men_n30_), .B0(men_men_n50_), .B1(men_men_n34_), .Y(men_men_n62_));
  NA4        u052(.A(men_men_n62_), .B(men_men_n53_), .C(men_men_n44_), .D(men_men_n28_), .Y(men_men_n63_));
  NA2        u053(.A(i_8_), .B(i_7_), .Y(men_men_n64_));
  NO2        u054(.A(men_men_n64_), .B(i_1_), .Y(men_men_n65_));
  NA2        u055(.A(i_8_), .B(men_men_n22_), .Y(men_men_n66_));
  AOI220     u056(.A0(men_men_n42_), .A1(i_1_), .B0(men_men_n38_), .B1(i_2_), .Y(men_men_n67_));
  NOi21      u057(.An(i_1_), .B(i_2_), .Y(men_men_n68_));
  NA3        u058(.A(men_men_n68_), .B(men_men_n47_), .C(i_6_), .Y(men_men_n69_));
  OAI210     u059(.A0(men_men_n67_), .A1(men_men_n66_), .B0(men_men_n69_), .Y(men_men_n70_));
  OAI210     u060(.A0(men_men_n70_), .A1(men_men_n65_), .B0(men_men_n14_), .Y(men_men_n71_));
  NA3        u061(.A(men_men_n59_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n72_));
  NA3        u062(.A(men_men_n25_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n73_));
  NA2        u063(.A(men_men_n73_), .B(men_men_n72_), .Y(men_men_n74_));
  NA2        u064(.A(men_men_n74_), .B(men_men_n55_), .Y(men_men_n75_));
  NA2        u065(.A(men_men_n75_), .B(men_men_n71_), .Y(men_men_n76_));
  NAi21      u066(.An(i_3_), .B(i_6_), .Y(men_men_n77_));
  NO3        u067(.A(men_men_n77_), .B(i_0_), .C(men_men_n45_), .Y(men_men_n78_));
  NOi21      u068(.An(i_7_), .B(i_8_), .Y(men_men_n79_));
  NOi31      u069(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n80_));
  AOI210     u070(.A0(men_men_n79_), .A1(men_men_n12_), .B0(men_men_n80_), .Y(men_men_n81_));
  NO2        u071(.A(men_men_n81_), .B(men_men_n11_), .Y(men_men_n82_));
  OAI210     u072(.A0(men_men_n82_), .A1(men_men_n78_), .B0(men_men_n68_), .Y(men_men_n83_));
  NA3        u073(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n84_));
  AOI210     u074(.A0(i_4_), .A1(i_3_), .B0(men_men_n84_), .Y(men_men_n85_));
  NA3        u075(.A(men_men_n21_), .B(i_5_), .C(i_7_), .Y(men_men_n86_));
  NO2        u076(.A(men_men_n86_), .B(i_2_), .Y(men_men_n87_));
  NO2        u077(.A(men_men_n87_), .B(men_men_n85_), .Y(men_men_n88_));
  NA3        u078(.A(men_men_n59_), .B(men_men_n30_), .C(i_3_), .Y(men_men_n89_));
  AOI210     u079(.A0(i_1_), .A1(i_4_), .B0(men_men_n89_), .Y(men_men_n90_));
  NAi21      u080(.An(i_6_), .B(i_0_), .Y(men_men_n91_));
  NA3        u081(.A(men_men_n56_), .B(i_5_), .C(men_men_n22_), .Y(men_men_n92_));
  NOi21      u082(.An(i_4_), .B(i_6_), .Y(men_men_n93_));
  NOi21      u083(.An(i_5_), .B(i_3_), .Y(men_men_n94_));
  NA3        u084(.A(men_men_n94_), .B(men_men_n68_), .C(men_men_n93_), .Y(men_men_n95_));
  OAI210     u085(.A0(men_men_n92_), .A1(men_men_n91_), .B0(men_men_n95_), .Y(men_men_n96_));
  NA2        u086(.A(men_men_n68_), .B(men_men_n32_), .Y(men_men_n97_));
  NOi21      u087(.An(men_men_n39_), .B(men_men_n97_), .Y(men_men_n98_));
  NO3        u088(.A(men_men_n98_), .B(men_men_n96_), .C(men_men_n90_), .Y(men_men_n99_));
  NOi21      u089(.An(i_6_), .B(i_1_), .Y(men_men_n100_));
  AOI220     u090(.A0(men_men_n100_), .A1(i_7_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n101_));
  NOi21      u091(.An(men_men_n47_), .B(men_men_n101_), .Y(men_men_n102_));
  NA2        u092(.A(men_men_n32_), .B(men_men_n14_), .Y(men_men_n103_));
  NOi21      u093(.An(i_3_), .B(i_1_), .Y(men_men_n104_));
  INV        u094(.A(men_men_n104_), .Y(men_men_n105_));
  NO2        u095(.A(men_men_n103_), .B(men_men_n105_), .Y(men_men_n106_));
  AOI210     u096(.A0(men_men_n79_), .A1(men_men_n14_), .B0(men_men_n93_), .Y(men_men_n107_));
  NOi31      u097(.An(men_men_n42_), .B(men_men_n107_), .C(men_men_n30_), .Y(men_men_n108_));
  NO3        u098(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n102_), .Y(men_men_n109_));
  NA4        u099(.A(men_men_n109_), .B(men_men_n99_), .C(men_men_n88_), .D(men_men_n83_), .Y(men_men_n110_));
  NA2        u100(.A(men_men_n50_), .B(men_men_n15_), .Y(men_men_n111_));
  NOi31      u101(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n112_));
  NA2        u102(.A(men_men_n112_), .B(i_7_), .Y(men_men_n113_));
  NA3        u103(.A(men_men_n32_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n114_));
  NA4        u104(.A(men_men_n114_), .B(men_men_n113_), .C(men_men_n111_), .D(men_men_n97_), .Y(men_men_n115_));
  NA2        u105(.A(men_men_n115_), .B(men_men_n37_), .Y(men_men_n116_));
  NAi31      u106(.An(men_men_n91_), .B(men_men_n79_), .C(i_2_), .Y(men_men_n117_));
  NA2        u107(.A(men_men_n59_), .B(men_men_n54_), .Y(men_men_n118_));
  NA2        u108(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n119_));
  NOi21      u109(.An(i_0_), .B(i_2_), .Y(men_men_n120_));
  NA3        u110(.A(men_men_n120_), .B(men_men_n33_), .C(men_men_n93_), .Y(men_men_n121_));
  NA3        u111(.A(men_men_n47_), .B(men_men_n39_), .C(men_men_n18_), .Y(men_men_n122_));
  NA3        u112(.A(men_men_n120_), .B(men_men_n55_), .C(men_men_n32_), .Y(men_men_n123_));
  NA3        u113(.A(men_men_n123_), .B(men_men_n122_), .C(men_men_n121_), .Y(men_men_n124_));
  NA4        u114(.A(men_men_n56_), .B(men_men_n34_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n125_));
  INV        u115(.A(men_men_n125_), .Y(men_men_n126_));
  NO3        u116(.A(men_men_n126_), .B(men_men_n124_), .C(men_men_n119_), .Y(men_men_n127_));
  NO3        u117(.A(i_2_), .B(men_men_n11_), .C(men_men_n14_), .Y(men_men_n128_));
  NA2        u118(.A(i_2_), .B(i_4_), .Y(men_men_n129_));
  AOI210     u119(.A0(men_men_n91_), .A1(men_men_n77_), .B0(men_men_n129_), .Y(men_men_n130_));
  NO2        u120(.A(i_8_), .B(i_7_), .Y(men_men_n131_));
  OA210      u121(.A0(men_men_n130_), .A1(men_men_n128_), .B0(men_men_n131_), .Y(men_men_n132_));
  NA3        u122(.A(men_men_n104_), .B(i_5_), .C(men_men_n22_), .Y(men_men_n133_));
  INV        u123(.A(men_men_n133_), .Y(men_men_n134_));
  NO2        u124(.A(men_men_n134_), .B(men_men_n132_), .Y(men_men_n135_));
  INV        u125(.A(men_men_n79_), .Y(men_men_n136_));
  INV        u126(.A(men_men_n47_), .Y(men_men_n137_));
  NO2        u127(.A(men_men_n137_), .B(men_men_n136_), .Y(men_men_n138_));
  NA3        u128(.A(men_men_n120_), .B(men_men_n59_), .C(men_men_n93_), .Y(men_men_n139_));
  INV        u129(.A(men_men_n139_), .Y(men_men_n140_));
  NA3        u130(.A(men_men_n94_), .B(men_men_n57_), .C(men_men_n41_), .Y(men_men_n141_));
  INV        u131(.A(men_men_n141_), .Y(men_men_n142_));
  NO3        u132(.A(men_men_n142_), .B(men_men_n140_), .C(men_men_n138_), .Y(men_men_n143_));
  NA4        u133(.A(men_men_n143_), .B(men_men_n135_), .C(men_men_n127_), .D(men_men_n116_), .Y(men_men_n144_));
  OR4        u134(.A(men_men_n144_), .B(men_men_n110_), .C(men_men_n76_), .D(men_men_n63_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule