library verilog;
use verilog.vl_types.all;
entity latchDSR_vlg_vec_tst is
end latchDSR_vlg_vec_tst;
