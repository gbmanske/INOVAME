library verilog;
use verilog.vl_types.all;
entity shiftreg4bitsbib_vlg_vec_tst is
end shiftreg4bitsbib_vlg_vec_tst;
