library verilog;
use verilog.vl_types.all;
entity ChaveCarro_vlg_vec_tst is
end ChaveCarro_vlg_vec_tst;
