library verilog;
use verilog.vl_types.all;
entity freqdiv4 is
    port(
        clk             : in     vl_logic;
        q               : out    vl_logic
    );
end freqdiv4;
