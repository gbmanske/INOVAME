//Benchmark atmr_misex3_1774_0.0156

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1374_, ori_ori_n1375_, ori_ori_n1376_, ori_ori_n1377_, ori_ori_n1378_, ori_ori_n1379_, ori_ori_n1380_, ori_ori_n1381_, ori_ori_n1382_, ori_ori_n1383_, ori_ori_n1384_, ori_ori_n1385_, ori_ori_n1386_, ori_ori_n1387_, ori_ori_n1388_, ori_ori_n1389_, ori_ori_n1390_, ori_ori_n1391_, ori_ori_n1392_, ori_ori_n1393_, ori_ori_n1394_, ori_ori_n1395_, ori_ori_n1396_, ori_ori_n1397_, ori_ori_n1398_, ori_ori_n1399_, ori_ori_n1404_, ori_ori_n1405_, ori_ori_n1406_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1533_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1540_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1544_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1549_, mai_mai_n1550_, mai_mai_n1551_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(g), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(g), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o0010(.A(ori_ori_n38_), .B(n), .Y(ori_ori_n39_));
  INV        o0011(.A(h), .Y(ori_ori_n40_));
  NAi21      o0012(.An(j), .B(l), .Y(ori_ori_n41_));
  NAi32      o0013(.An(n), .Bn(g), .C(m), .Y(ori_ori_n42_));
  NO3        o0014(.A(ori_ori_n42_), .B(ori_ori_n41_), .C(ori_ori_n40_), .Y(ori_ori_n43_));
  NAi31      o0015(.An(n), .B(m), .C(l), .Y(ori_ori_n44_));
  INV        o0016(.A(i), .Y(ori_ori_n45_));
  AN2        o0017(.A(h), .B(g), .Y(ori_ori_n46_));
  NA2        o0018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NAi21      o0020(.An(n), .B(m), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(l), .Y(ori_ori_n50_));
  NOi32      o0022(.An(k), .Bn(h), .C(g), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NO2        o0024(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  NO4        o0025(.A(ori_ori_n53_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n54_));
  AOI210     o0026(.A0(ori_ori_n54_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n55_));
  INV        o0027(.A(c), .Y(ori_ori_n56_));
  NA2        o0028(.A(e), .B(b), .Y(ori_ori_n57_));
  NO2        o0029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0030(.A(d), .Y(ori_ori_n59_));
  NA2        o0031(.A(g), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NAi21      o0032(.An(i), .B(h), .Y(ori_ori_n61_));
  NAi31      o0033(.An(i), .B(l), .C(j), .Y(ori_ori_n62_));
  OAI220     o0034(.A0(ori_ori_n62_), .A1(ori_ori_n49_), .B0(ori_ori_n61_), .B1(ori_ori_n44_), .Y(ori_ori_n63_));
  NAi31      o0035(.An(ori_ori_n60_), .B(ori_ori_n63_), .C(ori_ori_n58_), .Y(ori_ori_n64_));
  NAi41      o0036(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n65_));
  NA2        o0037(.A(g), .B(f), .Y(ori_ori_n66_));
  NO2        o0038(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  NAi21      o0039(.An(i), .B(j), .Y(ori_ori_n68_));
  NAi32      o0040(.An(n), .Bn(k), .C(m), .Y(ori_ori_n69_));
  NAi21      o0041(.An(e), .B(h), .Y(ori_ori_n70_));
  NAi41      o0042(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n71_));
  INV        o0043(.A(m), .Y(ori_ori_n72_));
  NOi21      o0044(.An(k), .B(l), .Y(ori_ori_n73_));
  NA2        o0045(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  AN4        o0046(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n75_));
  NOi31      o0047(.An(h), .B(g), .C(f), .Y(ori_ori_n76_));
  NA2        o0048(.A(ori_ori_n76_), .B(ori_ori_n75_), .Y(ori_ori_n77_));
  NAi32      o0049(.An(m), .Bn(k), .C(j), .Y(ori_ori_n78_));
  NOi32      o0050(.An(h), .Bn(g), .C(f), .Y(ori_ori_n79_));
  NA2        o0051(.A(ori_ori_n79_), .B(ori_ori_n75_), .Y(ori_ori_n80_));
  OA220      o0052(.A0(ori_ori_n80_), .A1(ori_ori_n78_), .B0(ori_ori_n77_), .B1(ori_ori_n74_), .Y(ori_ori_n81_));
  NA2        o0053(.A(ori_ori_n81_), .B(ori_ori_n64_), .Y(ori_ori_n82_));
  INV        o0054(.A(n), .Y(ori_ori_n83_));
  NOi32      o0055(.An(e), .Bn(b), .C(d), .Y(ori_ori_n84_));
  NA2        o0056(.A(ori_ori_n84_), .B(ori_ori_n83_), .Y(ori_ori_n85_));
  INV        o0057(.A(j), .Y(ori_ori_n86_));
  AN3        o0058(.A(m), .B(k), .C(i), .Y(ori_ori_n87_));
  NA3        o0059(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(g), .Y(ori_ori_n88_));
  NO2        o0060(.A(ori_ori_n88_), .B(f), .Y(ori_ori_n89_));
  NAi32      o0061(.An(g), .Bn(f), .C(h), .Y(ori_ori_n90_));
  NAi31      o0062(.An(j), .B(m), .C(l), .Y(ori_ori_n91_));
  NO2        o0063(.A(ori_ori_n91_), .B(ori_ori_n90_), .Y(ori_ori_n92_));
  NA2        o0064(.A(m), .B(l), .Y(ori_ori_n93_));
  NAi31      o0065(.An(k), .B(j), .C(g), .Y(ori_ori_n94_));
  NO3        o0066(.A(ori_ori_n94_), .B(ori_ori_n93_), .C(f), .Y(ori_ori_n95_));
  AN2        o0067(.A(j), .B(g), .Y(ori_ori_n96_));
  NOi32      o0068(.An(m), .Bn(l), .C(i), .Y(ori_ori_n97_));
  NOi21      o0069(.An(g), .B(i), .Y(ori_ori_n98_));
  NOi32      o0070(.An(m), .Bn(j), .C(k), .Y(ori_ori_n99_));
  AOI220     o0071(.A0(ori_ori_n99_), .A1(ori_ori_n98_), .B0(ori_ori_n97_), .B1(ori_ori_n96_), .Y(ori_ori_n100_));
  NO2        o0072(.A(ori_ori_n100_), .B(f), .Y(ori_ori_n101_));
  NO3        o0073(.A(ori_ori_n101_), .B(ori_ori_n95_), .C(ori_ori_n89_), .Y(ori_ori_n102_));
  NAi41      o0074(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n103_));
  AN2        o0075(.A(e), .B(b), .Y(ori_ori_n104_));
  NOi31      o0076(.An(c), .B(h), .C(f), .Y(ori_ori_n105_));
  NA2        o0077(.A(ori_ori_n105_), .B(ori_ori_n104_), .Y(ori_ori_n106_));
  NO2        o0078(.A(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n107_));
  NOi21      o0079(.An(g), .B(f), .Y(ori_ori_n108_));
  NOi21      o0080(.An(i), .B(h), .Y(ori_ori_n109_));
  NA3        o0081(.A(ori_ori_n109_), .B(ori_ori_n108_), .C(ori_ori_n36_), .Y(ori_ori_n110_));
  INV        o0082(.A(a), .Y(ori_ori_n111_));
  NA2        o0083(.A(ori_ori_n104_), .B(ori_ori_n111_), .Y(ori_ori_n112_));
  INV        o0084(.A(l), .Y(ori_ori_n113_));
  NOi21      o0085(.An(m), .B(n), .Y(ori_ori_n114_));
  AN2        o0086(.A(k), .B(h), .Y(ori_ori_n115_));
  NO2        o0087(.A(ori_ori_n110_), .B(ori_ori_n85_), .Y(ori_ori_n116_));
  INV        o0088(.A(b), .Y(ori_ori_n117_));
  NA2        o0089(.A(l), .B(j), .Y(ori_ori_n118_));
  AN2        o0090(.A(k), .B(i), .Y(ori_ori_n119_));
  NA2        o0091(.A(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n120_));
  NA2        o0092(.A(g), .B(e), .Y(ori_ori_n121_));
  NOi32      o0093(.An(c), .Bn(a), .C(d), .Y(ori_ori_n122_));
  NA2        o0094(.A(ori_ori_n122_), .B(ori_ori_n114_), .Y(ori_ori_n123_));
  NO2        o0095(.A(ori_ori_n116_), .B(ori_ori_n107_), .Y(ori_ori_n124_));
  OAI210     o0096(.A0(ori_ori_n102_), .A1(ori_ori_n85_), .B0(ori_ori_n124_), .Y(ori_ori_n125_));
  NOi31      o0097(.An(k), .B(m), .C(j), .Y(ori_ori_n126_));
  NA3        o0098(.A(ori_ori_n126_), .B(ori_ori_n76_), .C(ori_ori_n75_), .Y(ori_ori_n127_));
  NOi31      o0099(.An(k), .B(m), .C(i), .Y(ori_ori_n128_));
  NA3        o0100(.A(ori_ori_n128_), .B(ori_ori_n79_), .C(ori_ori_n75_), .Y(ori_ori_n129_));
  NA2        o0101(.A(ori_ori_n129_), .B(ori_ori_n127_), .Y(ori_ori_n130_));
  NOi32      o0102(.An(f), .Bn(b), .C(e), .Y(ori_ori_n131_));
  NAi21      o0103(.An(g), .B(h), .Y(ori_ori_n132_));
  NAi21      o0104(.An(m), .B(n), .Y(ori_ori_n133_));
  NAi21      o0105(.An(j), .B(k), .Y(ori_ori_n134_));
  NO3        o0106(.A(ori_ori_n134_), .B(ori_ori_n133_), .C(ori_ori_n132_), .Y(ori_ori_n135_));
  NAi41      o0107(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n136_));
  NAi31      o0108(.An(j), .B(k), .C(h), .Y(ori_ori_n137_));
  NO3        o0109(.A(ori_ori_n137_), .B(ori_ori_n136_), .C(ori_ori_n133_), .Y(ori_ori_n138_));
  AOI210     o0110(.A0(ori_ori_n135_), .A1(ori_ori_n131_), .B0(ori_ori_n138_), .Y(ori_ori_n139_));
  NO2        o0111(.A(k), .B(j), .Y(ori_ori_n140_));
  NO2        o0112(.A(ori_ori_n140_), .B(ori_ori_n133_), .Y(ori_ori_n141_));
  AN2        o0113(.A(k), .B(j), .Y(ori_ori_n142_));
  NAi21      o0114(.An(c), .B(b), .Y(ori_ori_n143_));
  NA2        o0115(.A(f), .B(d), .Y(ori_ori_n144_));
  NO4        o0116(.A(ori_ori_n144_), .B(ori_ori_n143_), .C(ori_ori_n142_), .D(ori_ori_n132_), .Y(ori_ori_n145_));
  NA2        o0117(.A(h), .B(c), .Y(ori_ori_n146_));
  NAi31      o0118(.An(f), .B(e), .C(b), .Y(ori_ori_n147_));
  NA2        o0119(.A(ori_ori_n145_), .B(ori_ori_n141_), .Y(ori_ori_n148_));
  NA2        o0120(.A(d), .B(b), .Y(ori_ori_n149_));
  NAi21      o0121(.An(e), .B(f), .Y(ori_ori_n150_));
  NO2        o0122(.A(ori_ori_n150_), .B(ori_ori_n149_), .Y(ori_ori_n151_));
  NA2        o0123(.A(b), .B(a), .Y(ori_ori_n152_));
  NAi21      o0124(.An(e), .B(g), .Y(ori_ori_n153_));
  NAi21      o0125(.An(c), .B(d), .Y(ori_ori_n154_));
  NAi31      o0126(.An(l), .B(k), .C(h), .Y(ori_ori_n155_));
  NO2        o0127(.A(ori_ori_n133_), .B(ori_ori_n155_), .Y(ori_ori_n156_));
  NA2        o0128(.A(ori_ori_n156_), .B(ori_ori_n151_), .Y(ori_ori_n157_));
  NAi41      o0129(.An(ori_ori_n130_), .B(ori_ori_n157_), .C(ori_ori_n148_), .D(ori_ori_n139_), .Y(ori_ori_n158_));
  NAi31      o0130(.An(e), .B(f), .C(b), .Y(ori_ori_n159_));
  NOi21      o0131(.An(g), .B(d), .Y(ori_ori_n160_));
  NO2        o0132(.A(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  NOi21      o0133(.An(h), .B(i), .Y(ori_ori_n162_));
  NOi21      o0134(.An(k), .B(m), .Y(ori_ori_n163_));
  NA3        o0135(.A(ori_ori_n163_), .B(ori_ori_n162_), .C(n), .Y(ori_ori_n164_));
  NOi21      o0136(.An(ori_ori_n161_), .B(ori_ori_n164_), .Y(ori_ori_n165_));
  NOi21      o0137(.An(h), .B(g), .Y(ori_ori_n166_));
  NO2        o0138(.A(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n167_));
  NAi31      o0139(.An(l), .B(j), .C(h), .Y(ori_ori_n168_));
  NO2        o0140(.A(ori_ori_n168_), .B(ori_ori_n49_), .Y(ori_ori_n169_));
  NA2        o0141(.A(ori_ori_n169_), .B(ori_ori_n67_), .Y(ori_ori_n170_));
  NOi32      o0142(.An(n), .Bn(k), .C(m), .Y(ori_ori_n171_));
  NA2        o0143(.A(l), .B(i), .Y(ori_ori_n172_));
  INV        o0144(.A(ori_ori_n170_), .Y(ori_ori_n173_));
  NAi31      o0145(.An(d), .B(f), .C(c), .Y(ori_ori_n174_));
  NAi31      o0146(.An(e), .B(f), .C(c), .Y(ori_ori_n175_));
  NA2        o0147(.A(ori_ori_n175_), .B(ori_ori_n174_), .Y(ori_ori_n176_));
  NA2        o0148(.A(j), .B(h), .Y(ori_ori_n177_));
  OR3        o0149(.A(n), .B(m), .C(k), .Y(ori_ori_n178_));
  NO2        o0150(.A(ori_ori_n178_), .B(ori_ori_n177_), .Y(ori_ori_n179_));
  NAi32      o0151(.An(m), .Bn(k), .C(n), .Y(ori_ori_n180_));
  NO2        o0152(.A(ori_ori_n180_), .B(ori_ori_n177_), .Y(ori_ori_n181_));
  AOI220     o0153(.A0(ori_ori_n181_), .A1(ori_ori_n161_), .B0(ori_ori_n179_), .B1(ori_ori_n176_), .Y(ori_ori_n182_));
  NO2        o0154(.A(n), .B(m), .Y(ori_ori_n183_));
  NA2        o0155(.A(ori_ori_n183_), .B(ori_ori_n50_), .Y(ori_ori_n184_));
  NAi21      o0156(.An(f), .B(e), .Y(ori_ori_n185_));
  NA2        o0157(.A(d), .B(c), .Y(ori_ori_n186_));
  NO2        o0158(.A(ori_ori_n186_), .B(ori_ori_n185_), .Y(ori_ori_n187_));
  NOi21      o0159(.An(ori_ori_n187_), .B(ori_ori_n184_), .Y(ori_ori_n188_));
  NAi31      o0160(.An(m), .B(n), .C(b), .Y(ori_ori_n189_));
  NA2        o0161(.A(k), .B(i), .Y(ori_ori_n190_));
  NAi21      o0162(.An(h), .B(f), .Y(ori_ori_n191_));
  NO2        o0163(.A(ori_ori_n191_), .B(ori_ori_n190_), .Y(ori_ori_n192_));
  NO2        o0164(.A(ori_ori_n189_), .B(ori_ori_n154_), .Y(ori_ori_n193_));
  NA2        o0165(.A(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n194_));
  NOi32      o0166(.An(f), .Bn(c), .C(d), .Y(ori_ori_n195_));
  NOi32      o0167(.An(f), .Bn(c), .C(e), .Y(ori_ori_n196_));
  NO2        o0168(.A(ori_ori_n196_), .B(ori_ori_n195_), .Y(ori_ori_n197_));
  NO3        o0169(.A(n), .B(m), .C(j), .Y(ori_ori_n198_));
  NA2        o0170(.A(ori_ori_n198_), .B(ori_ori_n115_), .Y(ori_ori_n199_));
  AO210      o0171(.A0(ori_ori_n199_), .A1(ori_ori_n184_), .B0(ori_ori_n197_), .Y(ori_ori_n200_));
  NAi41      o0172(.An(ori_ori_n188_), .B(ori_ori_n200_), .C(ori_ori_n194_), .D(ori_ori_n182_), .Y(ori_ori_n201_));
  OR4        o0173(.A(ori_ori_n201_), .B(ori_ori_n173_), .C(ori_ori_n165_), .D(ori_ori_n158_), .Y(ori_ori_n202_));
  NO4        o0174(.A(ori_ori_n202_), .B(ori_ori_n125_), .C(ori_ori_n82_), .D(ori_ori_n55_), .Y(ori_ori_n203_));
  NA3        o0175(.A(m), .B(ori_ori_n113_), .C(j), .Y(ori_ori_n204_));
  NAi31      o0176(.An(n), .B(h), .C(g), .Y(ori_ori_n205_));
  NO2        o0177(.A(ori_ori_n205_), .B(ori_ori_n204_), .Y(ori_ori_n206_));
  NOi32      o0178(.An(m), .Bn(k), .C(l), .Y(ori_ori_n207_));
  NA3        o0179(.A(ori_ori_n207_), .B(ori_ori_n86_), .C(g), .Y(ori_ori_n208_));
  NO2        o0180(.A(ori_ori_n208_), .B(n), .Y(ori_ori_n209_));
  NOi21      o0181(.An(k), .B(j), .Y(ori_ori_n210_));
  NA4        o0182(.A(ori_ori_n210_), .B(ori_ori_n114_), .C(i), .D(g), .Y(ori_ori_n211_));
  AN2        o0183(.A(i), .B(g), .Y(ori_ori_n212_));
  NA3        o0184(.A(ori_ori_n73_), .B(ori_ori_n212_), .C(ori_ori_n114_), .Y(ori_ori_n213_));
  NA2        o0185(.A(ori_ori_n213_), .B(ori_ori_n211_), .Y(ori_ori_n214_));
  NO3        o0186(.A(ori_ori_n214_), .B(ori_ori_n209_), .C(ori_ori_n206_), .Y(ori_ori_n215_));
  NAi41      o0187(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n216_));
  INV        o0188(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  INV        o0189(.A(f), .Y(ori_ori_n218_));
  INV        o0190(.A(g), .Y(ori_ori_n219_));
  NOi31      o0191(.An(i), .B(j), .C(h), .Y(ori_ori_n220_));
  NOi21      o0192(.An(l), .B(m), .Y(ori_ori_n221_));
  NA2        o0193(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NO3        o0194(.A(ori_ori_n222_), .B(ori_ori_n219_), .C(ori_ori_n218_), .Y(ori_ori_n223_));
  NA2        o0195(.A(ori_ori_n223_), .B(ori_ori_n217_), .Y(ori_ori_n224_));
  OAI210     o0196(.A0(ori_ori_n215_), .A1(ori_ori_n32_), .B0(ori_ori_n224_), .Y(ori_ori_n225_));
  NOi21      o0197(.An(n), .B(m), .Y(ori_ori_n226_));
  NOi32      o0198(.An(l), .Bn(i), .C(j), .Y(ori_ori_n227_));
  NA2        o0199(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  OA220      o0200(.A0(ori_ori_n228_), .A1(ori_ori_n106_), .B0(ori_ori_n78_), .B1(ori_ori_n77_), .Y(ori_ori_n229_));
  NAi21      o0201(.An(j), .B(h), .Y(ori_ori_n230_));
  XN2        o0202(.A(i), .B(h), .Y(ori_ori_n231_));
  NA2        o0203(.A(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NOi31      o0204(.An(k), .B(n), .C(m), .Y(ori_ori_n233_));
  NOi31      o0205(.An(ori_ori_n233_), .B(ori_ori_n186_), .C(ori_ori_n185_), .Y(ori_ori_n234_));
  NA2        o0206(.A(ori_ori_n234_), .B(ori_ori_n232_), .Y(ori_ori_n235_));
  NAi31      o0207(.An(f), .B(e), .C(c), .Y(ori_ori_n236_));
  NO4        o0208(.A(ori_ori_n236_), .B(ori_ori_n178_), .C(ori_ori_n177_), .D(ori_ori_n59_), .Y(ori_ori_n237_));
  NA4        o0209(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n238_));
  NAi32      o0210(.An(m), .Bn(i), .C(k), .Y(ori_ori_n239_));
  NO3        o0211(.A(ori_ori_n239_), .B(ori_ori_n90_), .C(ori_ori_n238_), .Y(ori_ori_n240_));
  INV        o0212(.A(k), .Y(ori_ori_n241_));
  NO2        o0213(.A(ori_ori_n240_), .B(ori_ori_n237_), .Y(ori_ori_n242_));
  NAi21      o0214(.An(n), .B(a), .Y(ori_ori_n243_));
  NO2        o0215(.A(ori_ori_n243_), .B(ori_ori_n149_), .Y(ori_ori_n244_));
  NAi41      o0216(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n245_), .B(e), .Y(ori_ori_n246_));
  NA2        o0218(.A(ori_ori_n246_), .B(ori_ori_n244_), .Y(ori_ori_n247_));
  AN4        o0219(.A(ori_ori_n247_), .B(ori_ori_n242_), .C(ori_ori_n235_), .D(ori_ori_n229_), .Y(ori_ori_n248_));
  OR2        o0220(.A(h), .B(g), .Y(ori_ori_n249_));
  NO2        o0221(.A(ori_ori_n249_), .B(ori_ori_n103_), .Y(ori_ori_n250_));
  NA2        o0222(.A(ori_ori_n250_), .B(ori_ori_n131_), .Y(ori_ori_n251_));
  NAi41      o0223(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n252_));
  NO2        o0224(.A(ori_ori_n252_), .B(ori_ori_n218_), .Y(ori_ori_n253_));
  NA2        o0225(.A(ori_ori_n163_), .B(ori_ori_n109_), .Y(ori_ori_n254_));
  NAi21      o0226(.An(ori_ori_n254_), .B(ori_ori_n253_), .Y(ori_ori_n255_));
  NO2        o0227(.A(n), .B(a), .Y(ori_ori_n256_));
  NAi31      o0228(.An(ori_ori_n245_), .B(ori_ori_n256_), .C(ori_ori_n104_), .Y(ori_ori_n257_));
  AN2        o0229(.A(ori_ori_n257_), .B(ori_ori_n255_), .Y(ori_ori_n258_));
  NAi21      o0230(.An(h), .B(i), .Y(ori_ori_n259_));
  NA2        o0231(.A(ori_ori_n183_), .B(k), .Y(ori_ori_n260_));
  NO2        o0232(.A(ori_ori_n260_), .B(ori_ori_n259_), .Y(ori_ori_n261_));
  NA2        o0233(.A(ori_ori_n261_), .B(ori_ori_n195_), .Y(ori_ori_n262_));
  NA3        o0234(.A(ori_ori_n262_), .B(ori_ori_n258_), .C(ori_ori_n251_), .Y(ori_ori_n263_));
  NOi21      o0235(.An(g), .B(e), .Y(ori_ori_n264_));
  NO2        o0236(.A(ori_ori_n71_), .B(ori_ori_n72_), .Y(ori_ori_n265_));
  NA2        o0237(.A(ori_ori_n265_), .B(ori_ori_n264_), .Y(ori_ori_n266_));
  NOi32      o0238(.An(l), .Bn(j), .C(i), .Y(ori_ori_n267_));
  AOI210     o0239(.A0(ori_ori_n73_), .A1(ori_ori_n86_), .B0(ori_ori_n267_), .Y(ori_ori_n268_));
  NO2        o0240(.A(ori_ori_n259_), .B(ori_ori_n44_), .Y(ori_ori_n269_));
  NAi21      o0241(.An(f), .B(g), .Y(ori_ori_n270_));
  NO2        o0242(.A(ori_ori_n270_), .B(ori_ori_n65_), .Y(ori_ori_n271_));
  NO2        o0243(.A(ori_ori_n69_), .B(ori_ori_n118_), .Y(ori_ori_n272_));
  AOI220     o0244(.A0(ori_ori_n272_), .A1(ori_ori_n271_), .B0(ori_ori_n269_), .B1(ori_ori_n67_), .Y(ori_ori_n273_));
  OAI210     o0245(.A0(ori_ori_n268_), .A1(ori_ori_n266_), .B0(ori_ori_n273_), .Y(ori_ori_n274_));
  NO2        o0246(.A(ori_ori_n134_), .B(ori_ori_n49_), .Y(ori_ori_n275_));
  NOi41      o0247(.An(ori_ori_n248_), .B(ori_ori_n274_), .C(ori_ori_n263_), .D(ori_ori_n225_), .Y(ori_ori_n276_));
  NO4        o0248(.A(ori_ori_n206_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n277_));
  NO2        o0249(.A(ori_ori_n277_), .B(ori_ori_n112_), .Y(ori_ori_n278_));
  NA3        o0250(.A(ori_ori_n59_), .B(c), .C(b), .Y(ori_ori_n279_));
  NAi21      o0251(.An(h), .B(g), .Y(ori_ori_n280_));
  OR4        o0252(.A(ori_ori_n280_), .B(ori_ori_n279_), .C(ori_ori_n228_), .D(e), .Y(ori_ori_n281_));
  NO2        o0253(.A(ori_ori_n254_), .B(ori_ori_n270_), .Y(ori_ori_n282_));
  NAi31      o0254(.An(g), .B(k), .C(h), .Y(ori_ori_n283_));
  NAi31      o0255(.An(e), .B(d), .C(a), .Y(ori_ori_n284_));
  INV        o0256(.A(ori_ori_n281_), .Y(ori_ori_n285_));
  NA4        o0257(.A(ori_ori_n163_), .B(ori_ori_n79_), .C(ori_ori_n75_), .D(ori_ori_n118_), .Y(ori_ori_n286_));
  NA3        o0258(.A(ori_ori_n163_), .B(ori_ori_n162_), .C(ori_ori_n83_), .Y(ori_ori_n287_));
  NO2        o0259(.A(ori_ori_n287_), .B(ori_ori_n197_), .Y(ori_ori_n288_));
  NOi21      o0260(.An(ori_ori_n286_), .B(ori_ori_n288_), .Y(ori_ori_n289_));
  NA3        o0261(.A(e), .B(c), .C(b), .Y(ori_ori_n290_));
  NO2        o0262(.A(ori_ori_n60_), .B(ori_ori_n290_), .Y(ori_ori_n291_));
  NAi32      o0263(.An(k), .Bn(i), .C(j), .Y(ori_ori_n292_));
  NAi31      o0264(.An(h), .B(l), .C(i), .Y(ori_ori_n293_));
  NA3        o0265(.A(ori_ori_n293_), .B(ori_ori_n292_), .C(ori_ori_n168_), .Y(ori_ori_n294_));
  NOi21      o0266(.An(ori_ori_n294_), .B(ori_ori_n49_), .Y(ori_ori_n295_));
  OAI210     o0267(.A0(ori_ori_n271_), .A1(ori_ori_n291_), .B0(ori_ori_n295_), .Y(ori_ori_n296_));
  NAi21      o0268(.An(l), .B(k), .Y(ori_ori_n297_));
  NO2        o0269(.A(ori_ori_n297_), .B(ori_ori_n49_), .Y(ori_ori_n298_));
  NOi21      o0270(.An(l), .B(j), .Y(ori_ori_n299_));
  NA2        o0271(.A(ori_ori_n166_), .B(ori_ori_n299_), .Y(ori_ori_n300_));
  NA3        o0272(.A(ori_ori_n119_), .B(ori_ori_n118_), .C(g), .Y(ori_ori_n301_));
  OR3        o0273(.A(ori_ori_n71_), .B(ori_ori_n72_), .C(e), .Y(ori_ori_n302_));
  AOI210     o0274(.A0(ori_ori_n301_), .A1(ori_ori_n300_), .B0(ori_ori_n302_), .Y(ori_ori_n303_));
  INV        o0275(.A(ori_ori_n303_), .Y(ori_ori_n304_));
  NAi32      o0276(.An(j), .Bn(h), .C(i), .Y(ori_ori_n305_));
  NAi21      o0277(.An(m), .B(l), .Y(ori_ori_n306_));
  NO3        o0278(.A(ori_ori_n306_), .B(ori_ori_n305_), .C(ori_ori_n83_), .Y(ori_ori_n307_));
  NA2        o0279(.A(h), .B(g), .Y(ori_ori_n308_));
  NA2        o0280(.A(ori_ori_n171_), .B(ori_ori_n45_), .Y(ori_ori_n309_));
  NO2        o0281(.A(ori_ori_n309_), .B(ori_ori_n308_), .Y(ori_ori_n310_));
  NA2        o0282(.A(ori_ori_n310_), .B(ori_ori_n167_), .Y(ori_ori_n311_));
  NA4        o0283(.A(ori_ori_n311_), .B(ori_ori_n304_), .C(ori_ori_n296_), .D(ori_ori_n289_), .Y(ori_ori_n312_));
  NO2        o0284(.A(ori_ori_n147_), .B(d), .Y(ori_ori_n313_));
  NA2        o0285(.A(ori_ori_n313_), .B(ori_ori_n53_), .Y(ori_ori_n314_));
  NO2        o0286(.A(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n315_));
  NAi32      o0287(.An(n), .Bn(m), .C(l), .Y(ori_ori_n316_));
  NO2        o0288(.A(ori_ori_n316_), .B(ori_ori_n305_), .Y(ori_ori_n317_));
  NA2        o0289(.A(ori_ori_n317_), .B(ori_ori_n187_), .Y(ori_ori_n318_));
  NO2        o0290(.A(ori_ori_n123_), .B(ori_ori_n117_), .Y(ori_ori_n319_));
  NAi31      o0291(.An(k), .B(l), .C(j), .Y(ori_ori_n320_));
  OAI210     o0292(.A0(ori_ori_n297_), .A1(j), .B0(ori_ori_n320_), .Y(ori_ori_n321_));
  NOi21      o0293(.An(ori_ori_n321_), .B(ori_ori_n121_), .Y(ori_ori_n322_));
  NA2        o0294(.A(ori_ori_n322_), .B(ori_ori_n319_), .Y(ori_ori_n323_));
  NA3        o0295(.A(ori_ori_n323_), .B(ori_ori_n318_), .C(ori_ori_n314_), .Y(ori_ori_n324_));
  NO4        o0296(.A(ori_ori_n324_), .B(ori_ori_n312_), .C(ori_ori_n285_), .D(ori_ori_n278_), .Y(ori_ori_n325_));
  NA2        o0297(.A(ori_ori_n261_), .B(ori_ori_n196_), .Y(ori_ori_n326_));
  NAi21      o0298(.An(m), .B(k), .Y(ori_ori_n327_));
  NO2        o0299(.A(ori_ori_n231_), .B(ori_ori_n327_), .Y(ori_ori_n328_));
  NAi41      o0300(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n329_));
  NO2        o0301(.A(ori_ori_n329_), .B(ori_ori_n153_), .Y(ori_ori_n330_));
  NA2        o0302(.A(ori_ori_n330_), .B(ori_ori_n328_), .Y(ori_ori_n331_));
  NAi31      o0303(.An(i), .B(l), .C(h), .Y(ori_ori_n332_));
  NO4        o0304(.A(ori_ori_n332_), .B(ori_ori_n153_), .C(ori_ori_n71_), .D(ori_ori_n72_), .Y(ori_ori_n333_));
  NA2        o0305(.A(e), .B(c), .Y(ori_ori_n334_));
  NO3        o0306(.A(ori_ori_n334_), .B(n), .C(d), .Y(ori_ori_n335_));
  NOi21      o0307(.An(f), .B(h), .Y(ori_ori_n336_));
  NA2        o0308(.A(ori_ori_n336_), .B(ori_ori_n119_), .Y(ori_ori_n337_));
  NO2        o0309(.A(ori_ori_n337_), .B(ori_ori_n219_), .Y(ori_ori_n338_));
  NAi31      o0310(.An(d), .B(e), .C(b), .Y(ori_ori_n339_));
  NO2        o0311(.A(ori_ori_n133_), .B(ori_ori_n339_), .Y(ori_ori_n340_));
  NA2        o0312(.A(ori_ori_n340_), .B(ori_ori_n338_), .Y(ori_ori_n341_));
  NAi41      o0313(.An(ori_ori_n333_), .B(ori_ori_n341_), .C(ori_ori_n331_), .D(ori_ori_n326_), .Y(ori_ori_n342_));
  NO4        o0314(.A(ori_ori_n329_), .B(ori_ori_n78_), .C(ori_ori_n70_), .D(ori_ori_n219_), .Y(ori_ori_n343_));
  NA2        o0315(.A(ori_ori_n256_), .B(ori_ori_n104_), .Y(ori_ori_n344_));
  OR2        o0316(.A(ori_ori_n344_), .B(ori_ori_n208_), .Y(ori_ori_n345_));
  NOi31      o0317(.An(l), .B(n), .C(m), .Y(ori_ori_n346_));
  NA2        o0318(.A(ori_ori_n346_), .B(ori_ori_n220_), .Y(ori_ori_n347_));
  NO2        o0319(.A(ori_ori_n347_), .B(ori_ori_n197_), .Y(ori_ori_n348_));
  NAi32      o0320(.An(ori_ori_n348_), .Bn(ori_ori_n343_), .C(ori_ori_n345_), .Y(ori_ori_n349_));
  NAi32      o0321(.An(m), .Bn(j), .C(k), .Y(ori_ori_n350_));
  NAi41      o0322(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n351_));
  OAI210     o0323(.A0(ori_ori_n216_), .A1(ori_ori_n350_), .B0(ori_ori_n351_), .Y(ori_ori_n352_));
  NOi31      o0324(.An(j), .B(m), .C(k), .Y(ori_ori_n353_));
  NO2        o0325(.A(ori_ori_n126_), .B(ori_ori_n353_), .Y(ori_ori_n354_));
  AN3        o0326(.A(h), .B(g), .C(f), .Y(ori_ori_n355_));
  NAi31      o0327(.An(ori_ori_n354_), .B(ori_ori_n355_), .C(ori_ori_n352_), .Y(ori_ori_n356_));
  NOi32      o0328(.An(m), .Bn(j), .C(l), .Y(ori_ori_n357_));
  NO2        o0329(.A(ori_ori_n357_), .B(ori_ori_n97_), .Y(ori_ori_n358_));
  NO2        o0330(.A(ori_ori_n306_), .B(ori_ori_n305_), .Y(ori_ori_n359_));
  NO2        o0331(.A(ori_ori_n222_), .B(g), .Y(ori_ori_n360_));
  NO2        o0332(.A(ori_ori_n159_), .B(ori_ori_n83_), .Y(ori_ori_n361_));
  AOI220     o0333(.A0(ori_ori_n361_), .A1(ori_ori_n360_), .B0(ori_ori_n253_), .B1(ori_ori_n359_), .Y(ori_ori_n362_));
  NA2        o0334(.A(ori_ori_n239_), .B(ori_ori_n78_), .Y(ori_ori_n363_));
  NA3        o0335(.A(ori_ori_n363_), .B(ori_ori_n355_), .C(ori_ori_n217_), .Y(ori_ori_n364_));
  NA3        o0336(.A(ori_ori_n364_), .B(ori_ori_n362_), .C(ori_ori_n356_), .Y(ori_ori_n365_));
  NA3        o0337(.A(h), .B(g), .C(f), .Y(ori_ori_n366_));
  NO2        o0338(.A(ori_ori_n366_), .B(ori_ori_n74_), .Y(ori_ori_n367_));
  NA2        o0339(.A(ori_ori_n351_), .B(ori_ori_n216_), .Y(ori_ori_n368_));
  NA2        o0340(.A(ori_ori_n166_), .B(e), .Y(ori_ori_n369_));
  NO2        o0341(.A(ori_ori_n369_), .B(ori_ori_n41_), .Y(ori_ori_n370_));
  AOI220     o0342(.A0(ori_ori_n370_), .A1(ori_ori_n319_), .B0(ori_ori_n368_), .B1(ori_ori_n367_), .Y(ori_ori_n371_));
  NOi32      o0343(.An(j), .Bn(g), .C(i), .Y(ori_ori_n372_));
  NA3        o0344(.A(ori_ori_n372_), .B(ori_ori_n297_), .C(ori_ori_n114_), .Y(ori_ori_n373_));
  AO210      o0345(.A0(ori_ori_n112_), .A1(ori_ori_n32_), .B0(ori_ori_n373_), .Y(ori_ori_n374_));
  NOi32      o0346(.An(e), .Bn(b), .C(a), .Y(ori_ori_n375_));
  AN2        o0347(.A(l), .B(j), .Y(ori_ori_n376_));
  NO2        o0348(.A(ori_ori_n327_), .B(ori_ori_n376_), .Y(ori_ori_n377_));
  NO3        o0349(.A(ori_ori_n329_), .B(ori_ori_n70_), .C(ori_ori_n219_), .Y(ori_ori_n378_));
  NA3        o0350(.A(ori_ori_n213_), .B(ori_ori_n211_), .C(ori_ori_n35_), .Y(ori_ori_n379_));
  AOI220     o0351(.A0(ori_ori_n379_), .A1(ori_ori_n375_), .B0(ori_ori_n378_), .B1(ori_ori_n377_), .Y(ori_ori_n380_));
  NO2        o0352(.A(ori_ori_n339_), .B(n), .Y(ori_ori_n381_));
  NA2        o0353(.A(ori_ori_n212_), .B(k), .Y(ori_ori_n382_));
  NA3        o0354(.A(m), .B(ori_ori_n113_), .C(ori_ori_n218_), .Y(ori_ori_n383_));
  NA4        o0355(.A(ori_ori_n207_), .B(ori_ori_n86_), .C(g), .D(ori_ori_n218_), .Y(ori_ori_n384_));
  OAI210     o0356(.A0(ori_ori_n383_), .A1(ori_ori_n382_), .B0(ori_ori_n384_), .Y(ori_ori_n385_));
  NAi41      o0357(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n386_));
  NA2        o0358(.A(ori_ori_n51_), .B(ori_ori_n114_), .Y(ori_ori_n387_));
  NO2        o0359(.A(ori_ori_n387_), .B(ori_ori_n386_), .Y(ori_ori_n388_));
  AOI220     o0360(.A0(ori_ori_n388_), .A1(b), .B0(ori_ori_n385_), .B1(ori_ori_n381_), .Y(ori_ori_n389_));
  NA4        o0361(.A(ori_ori_n389_), .B(ori_ori_n380_), .C(ori_ori_n374_), .D(ori_ori_n371_), .Y(ori_ori_n390_));
  NO4        o0362(.A(ori_ori_n390_), .B(ori_ori_n365_), .C(ori_ori_n349_), .D(ori_ori_n342_), .Y(ori_ori_n391_));
  NA4        o0363(.A(ori_ori_n391_), .B(ori_ori_n325_), .C(ori_ori_n276_), .D(ori_ori_n203_), .Y(ori10));
  NA3        o0364(.A(m), .B(k), .C(i), .Y(ori_ori_n393_));
  NO3        o0365(.A(ori_ori_n393_), .B(j), .C(ori_ori_n219_), .Y(ori_ori_n394_));
  NOi21      o0366(.An(e), .B(f), .Y(ori_ori_n395_));
  NO4        o0367(.A(ori_ori_n154_), .B(ori_ori_n395_), .C(n), .D(ori_ori_n111_), .Y(ori_ori_n396_));
  NAi31      o0368(.An(b), .B(f), .C(c), .Y(ori_ori_n397_));
  INV        o0369(.A(ori_ori_n397_), .Y(ori_ori_n398_));
  NOi32      o0370(.An(k), .Bn(h), .C(j), .Y(ori_ori_n399_));
  NA2        o0371(.A(ori_ori_n399_), .B(ori_ori_n226_), .Y(ori_ori_n400_));
  NA2        o0372(.A(ori_ori_n164_), .B(ori_ori_n400_), .Y(ori_ori_n401_));
  AOI220     o0373(.A0(ori_ori_n401_), .A1(ori_ori_n398_), .B0(ori_ori_n396_), .B1(ori_ori_n394_), .Y(ori_ori_n402_));
  AN2        o0374(.A(j), .B(h), .Y(ori_ori_n403_));
  NO3        o0375(.A(n), .B(m), .C(k), .Y(ori_ori_n404_));
  NA2        o0376(.A(ori_ori_n404_), .B(ori_ori_n403_), .Y(ori_ori_n405_));
  NO3        o0377(.A(ori_ori_n405_), .B(ori_ori_n154_), .C(ori_ori_n218_), .Y(ori_ori_n406_));
  OR2        o0378(.A(m), .B(k), .Y(ori_ori_n407_));
  NO2        o0379(.A(ori_ori_n177_), .B(ori_ori_n407_), .Y(ori_ori_n408_));
  NA4        o0380(.A(n), .B(f), .C(c), .D(ori_ori_n117_), .Y(ori_ori_n409_));
  NOi21      o0381(.An(ori_ori_n408_), .B(ori_ori_n409_), .Y(ori_ori_n410_));
  NOi32      o0382(.An(d), .Bn(a), .C(c), .Y(ori_ori_n411_));
  NA2        o0383(.A(ori_ori_n411_), .B(ori_ori_n185_), .Y(ori_ori_n412_));
  NAi21      o0384(.An(i), .B(g), .Y(ori_ori_n413_));
  NAi31      o0385(.An(k), .B(m), .C(j), .Y(ori_ori_n414_));
  NO2        o0386(.A(ori_ori_n410_), .B(ori_ori_n406_), .Y(ori_ori_n415_));
  NO2        o0387(.A(ori_ori_n409_), .B(ori_ori_n306_), .Y(ori_ori_n416_));
  NOi32      o0388(.An(f), .Bn(d), .C(c), .Y(ori_ori_n417_));
  AOI220     o0389(.A0(ori_ori_n417_), .A1(ori_ori_n317_), .B0(ori_ori_n416_), .B1(ori_ori_n220_), .Y(ori_ori_n418_));
  NA3        o0390(.A(ori_ori_n418_), .B(ori_ori_n415_), .C(ori_ori_n402_), .Y(ori_ori_n419_));
  NO2        o0391(.A(ori_ori_n59_), .B(ori_ori_n117_), .Y(ori_ori_n420_));
  NA2        o0392(.A(ori_ori_n256_), .B(ori_ori_n420_), .Y(ori_ori_n421_));
  INV        o0393(.A(e), .Y(ori_ori_n422_));
  NA2        o0394(.A(ori_ori_n46_), .B(e), .Y(ori_ori_n423_));
  OAI220     o0395(.A0(ori_ori_n423_), .A1(ori_ori_n204_), .B0(ori_ori_n208_), .B1(ori_ori_n422_), .Y(ori_ori_n424_));
  AN2        o0396(.A(g), .B(e), .Y(ori_ori_n425_));
  NA3        o0397(.A(ori_ori_n425_), .B(ori_ori_n207_), .C(i), .Y(ori_ori_n426_));
  OAI210     o0398(.A0(ori_ori_n88_), .A1(ori_ori_n422_), .B0(ori_ori_n426_), .Y(ori_ori_n427_));
  NO2        o0399(.A(ori_ori_n100_), .B(ori_ori_n422_), .Y(ori_ori_n428_));
  NO3        o0400(.A(ori_ori_n428_), .B(ori_ori_n427_), .C(ori_ori_n424_), .Y(ori_ori_n429_));
  NOi32      o0401(.An(h), .Bn(e), .C(g), .Y(ori_ori_n430_));
  NA3        o0402(.A(ori_ori_n430_), .B(ori_ori_n299_), .C(m), .Y(ori_ori_n431_));
  NOi21      o0403(.An(g), .B(h), .Y(ori_ori_n432_));
  AN3        o0404(.A(m), .B(l), .C(i), .Y(ori_ori_n433_));
  NA3        o0405(.A(ori_ori_n433_), .B(ori_ori_n432_), .C(e), .Y(ori_ori_n434_));
  AN3        o0406(.A(h), .B(g), .C(e), .Y(ori_ori_n435_));
  NA2        o0407(.A(ori_ori_n435_), .B(ori_ori_n97_), .Y(ori_ori_n436_));
  AN3        o0408(.A(ori_ori_n436_), .B(ori_ori_n434_), .C(ori_ori_n431_), .Y(ori_ori_n437_));
  AOI210     o0409(.A0(ori_ori_n437_), .A1(ori_ori_n429_), .B0(ori_ori_n421_), .Y(ori_ori_n438_));
  NA3        o0410(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(e), .Y(ori_ori_n439_));
  NO2        o0411(.A(ori_ori_n439_), .B(ori_ori_n421_), .Y(ori_ori_n440_));
  NA3        o0412(.A(ori_ori_n411_), .B(ori_ori_n185_), .C(ori_ori_n83_), .Y(ori_ori_n441_));
  NAi31      o0413(.An(b), .B(c), .C(a), .Y(ori_ori_n442_));
  NO2        o0414(.A(ori_ori_n442_), .B(n), .Y(ori_ori_n443_));
  NA2        o0415(.A(ori_ori_n51_), .B(m), .Y(ori_ori_n444_));
  NO2        o0416(.A(ori_ori_n444_), .B(ori_ori_n150_), .Y(ori_ori_n445_));
  NA2        o0417(.A(ori_ori_n445_), .B(ori_ori_n443_), .Y(ori_ori_n446_));
  INV        o0418(.A(ori_ori_n446_), .Y(ori_ori_n447_));
  NO4        o0419(.A(ori_ori_n447_), .B(ori_ori_n440_), .C(ori_ori_n438_), .D(ori_ori_n419_), .Y(ori_ori_n448_));
  NA2        o0420(.A(i), .B(g), .Y(ori_ori_n449_));
  NOi21      o0421(.An(d), .B(c), .Y(ori_ori_n450_));
  NA3        o0422(.A(i), .B(g), .C(f), .Y(ori_ori_n451_));
  OR2        o0423(.A(n), .B(m), .Y(ori_ori_n452_));
  NO2        o0424(.A(ori_ori_n452_), .B(ori_ori_n155_), .Y(ori_ori_n453_));
  NO2        o0425(.A(ori_ori_n186_), .B(ori_ori_n150_), .Y(ori_ori_n454_));
  OAI210     o0426(.A0(ori_ori_n453_), .A1(ori_ori_n179_), .B0(ori_ori_n454_), .Y(ori_ori_n455_));
  INV        o0427(.A(ori_ori_n387_), .Y(ori_ori_n456_));
  NA3        o0428(.A(ori_ori_n456_), .B(ori_ori_n375_), .C(d), .Y(ori_ori_n457_));
  NO2        o0429(.A(ori_ori_n442_), .B(ori_ori_n49_), .Y(ori_ori_n458_));
  NO3        o0430(.A(ori_ori_n66_), .B(ori_ori_n113_), .C(e), .Y(ori_ori_n459_));
  NAi21      o0431(.An(k), .B(j), .Y(ori_ori_n460_));
  NA2        o0432(.A(ori_ori_n259_), .B(ori_ori_n460_), .Y(ori_ori_n461_));
  NA3        o0433(.A(ori_ori_n461_), .B(ori_ori_n459_), .C(ori_ori_n458_), .Y(ori_ori_n462_));
  NAi21      o0434(.An(e), .B(d), .Y(ori_ori_n463_));
  INV        o0435(.A(ori_ori_n463_), .Y(ori_ori_n464_));
  NO2        o0436(.A(ori_ori_n260_), .B(ori_ori_n218_), .Y(ori_ori_n465_));
  NA3        o0437(.A(ori_ori_n465_), .B(ori_ori_n464_), .C(ori_ori_n232_), .Y(ori_ori_n466_));
  NA4        o0438(.A(ori_ori_n466_), .B(ori_ori_n462_), .C(ori_ori_n457_), .D(ori_ori_n455_), .Y(ori_ori_n467_));
  NO2        o0439(.A(ori_ori_n347_), .B(ori_ori_n218_), .Y(ori_ori_n468_));
  NA2        o0440(.A(ori_ori_n468_), .B(ori_ori_n464_), .Y(ori_ori_n469_));
  NOi31      o0441(.An(n), .B(m), .C(k), .Y(ori_ori_n470_));
  AOI220     o0442(.A0(ori_ori_n470_), .A1(ori_ori_n403_), .B0(ori_ori_n226_), .B1(ori_ori_n50_), .Y(ori_ori_n471_));
  NAi31      o0443(.An(g), .B(f), .C(c), .Y(ori_ori_n472_));
  OR3        o0444(.A(ori_ori_n472_), .B(ori_ori_n471_), .C(e), .Y(ori_ori_n473_));
  NA3        o0445(.A(ori_ori_n473_), .B(ori_ori_n469_), .C(ori_ori_n318_), .Y(ori_ori_n474_));
  NO3        o0446(.A(ori_ori_n474_), .B(ori_ori_n467_), .C(ori_ori_n274_), .Y(ori_ori_n475_));
  NOi32      o0447(.An(c), .Bn(a), .C(b), .Y(ori_ori_n476_));
  NA2        o0448(.A(ori_ori_n476_), .B(ori_ori_n114_), .Y(ori_ori_n477_));
  INV        o0449(.A(ori_ori_n283_), .Y(ori_ori_n478_));
  AN2        o0450(.A(e), .B(d), .Y(ori_ori_n479_));
  NA2        o0451(.A(ori_ori_n479_), .B(ori_ori_n478_), .Y(ori_ori_n480_));
  INV        o0452(.A(ori_ori_n150_), .Y(ori_ori_n481_));
  NO2        o0453(.A(ori_ori_n132_), .B(ori_ori_n41_), .Y(ori_ori_n482_));
  NO2        o0454(.A(ori_ori_n66_), .B(e), .Y(ori_ori_n483_));
  NA4        o0455(.A(ori_ori_n332_), .B(ori_ori_n168_), .C(ori_ori_n268_), .D(ori_ori_n120_), .Y(ori_ori_n484_));
  AOI220     o0456(.A0(ori_ori_n484_), .A1(ori_ori_n483_), .B0(ori_ori_n482_), .B1(ori_ori_n481_), .Y(ori_ori_n485_));
  AOI210     o0457(.A0(ori_ori_n485_), .A1(ori_ori_n480_), .B0(ori_ori_n477_), .Y(ori_ori_n486_));
  NO2        o0458(.A(ori_ori_n214_), .B(ori_ori_n209_), .Y(ori_ori_n487_));
  NOi21      o0459(.An(a), .B(b), .Y(ori_ori_n488_));
  NA3        o0460(.A(e), .B(d), .C(c), .Y(ori_ori_n489_));
  NAi21      o0461(.An(ori_ori_n489_), .B(ori_ori_n488_), .Y(ori_ori_n490_));
  NO2        o0462(.A(ori_ori_n441_), .B(ori_ori_n208_), .Y(ori_ori_n491_));
  NOi21      o0463(.An(ori_ori_n490_), .B(ori_ori_n491_), .Y(ori_ori_n492_));
  AOI210     o0464(.A0(ori_ori_n277_), .A1(ori_ori_n487_), .B0(ori_ori_n492_), .Y(ori_ori_n493_));
  NO4        o0465(.A(ori_ori_n191_), .B(ori_ori_n103_), .C(ori_ori_n56_), .D(b), .Y(ori_ori_n494_));
  NA2        o0466(.A(ori_ori_n398_), .B(ori_ori_n156_), .Y(ori_ori_n495_));
  OR2        o0467(.A(k), .B(j), .Y(ori_ori_n496_));
  NA2        o0468(.A(l), .B(k), .Y(ori_ori_n497_));
  NA3        o0469(.A(ori_ori_n497_), .B(ori_ori_n496_), .C(ori_ori_n226_), .Y(ori_ori_n498_));
  AOI210     o0470(.A0(ori_ori_n239_), .A1(ori_ori_n350_), .B0(ori_ori_n83_), .Y(ori_ori_n499_));
  NOi21      o0471(.An(ori_ori_n498_), .B(ori_ori_n499_), .Y(ori_ori_n500_));
  OR3        o0472(.A(ori_ori_n500_), .B(ori_ori_n146_), .C(ori_ori_n136_), .Y(ori_ori_n501_));
  NA3        o0473(.A(ori_ori_n286_), .B(ori_ori_n129_), .C(ori_ori_n127_), .Y(ori_ori_n502_));
  NO3        o0474(.A(ori_ori_n441_), .B(ori_ori_n91_), .C(ori_ori_n132_), .Y(ori_ori_n503_));
  NO3        o0475(.A(ori_ori_n503_), .B(ori_ori_n502_), .C(ori_ori_n333_), .Y(ori_ori_n504_));
  NA3        o0476(.A(ori_ori_n504_), .B(ori_ori_n501_), .C(ori_ori_n495_), .Y(ori_ori_n505_));
  NO4        o0477(.A(ori_ori_n505_), .B(ori_ori_n494_), .C(ori_ori_n493_), .D(ori_ori_n486_), .Y(ori_ori_n506_));
  INV        o0478(.A(e), .Y(ori_ori_n507_));
  NO2        o0479(.A(ori_ori_n191_), .B(ori_ori_n56_), .Y(ori_ori_n508_));
  NAi31      o0480(.An(j), .B(l), .C(i), .Y(ori_ori_n509_));
  OAI210     o0481(.A0(ori_ori_n509_), .A1(ori_ori_n133_), .B0(ori_ori_n103_), .Y(ori_ori_n510_));
  NA4        o0482(.A(ori_ori_n510_), .B(ori_ori_n508_), .C(ori_ori_n507_), .D(b), .Y(ori_ori_n511_));
  NO3        o0483(.A(ori_ori_n412_), .B(ori_ori_n358_), .C(ori_ori_n205_), .Y(ori_ori_n512_));
  NO2        o0484(.A(ori_ori_n412_), .B(ori_ori_n387_), .Y(ori_ori_n513_));
  NO4        o0485(.A(ori_ori_n513_), .B(ori_ori_n512_), .C(ori_ori_n188_), .D(ori_ori_n315_), .Y(ori_ori_n514_));
  NA3        o0486(.A(ori_ori_n514_), .B(ori_ori_n511_), .C(ori_ori_n248_), .Y(ori_ori_n515_));
  OAI210     o0487(.A0(ori_ori_n128_), .A1(ori_ori_n126_), .B0(n), .Y(ori_ori_n516_));
  NO2        o0488(.A(ori_ori_n516_), .B(ori_ori_n132_), .Y(ori_ori_n517_));
  AN2        o0489(.A(ori_ori_n517_), .B(ori_ori_n196_), .Y(ori_ori_n518_));
  XO2        o0490(.A(i), .B(h), .Y(ori_ori_n519_));
  NA3        o0491(.A(ori_ori_n519_), .B(ori_ori_n163_), .C(n), .Y(ori_ori_n520_));
  NAi41      o0492(.An(ori_ori_n307_), .B(ori_ori_n520_), .C(ori_ori_n471_), .D(ori_ori_n400_), .Y(ori_ori_n521_));
  NOi32      o0493(.An(ori_ori_n521_), .Bn(ori_ori_n483_), .C(ori_ori_n279_), .Y(ori_ori_n522_));
  NAi31      o0494(.An(c), .B(f), .C(d), .Y(ori_ori_n523_));
  AOI210     o0495(.A0(ori_ori_n287_), .A1(ori_ori_n199_), .B0(ori_ori_n523_), .Y(ori_ori_n524_));
  NOi21      o0496(.An(ori_ori_n81_), .B(ori_ori_n524_), .Y(ori_ori_n525_));
  NA2        o0497(.A(ori_ori_n233_), .B(ori_ori_n109_), .Y(ori_ori_n526_));
  AOI210     o0498(.A0(ori_ori_n526_), .A1(ori_ori_n184_), .B0(ori_ori_n523_), .Y(ori_ori_n527_));
  INV        o0499(.A(ori_ori_n527_), .Y(ori_ori_n528_));
  AO220      o0500(.A0(ori_ori_n295_), .A1(ori_ori_n271_), .B0(ori_ori_n169_), .B1(ori_ori_n67_), .Y(ori_ori_n529_));
  NA3        o0501(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n530_));
  INV        o0502(.A(ori_ori_n303_), .Y(ori_ori_n531_));
  NAi41      o0503(.An(ori_ori_n529_), .B(ori_ori_n531_), .C(ori_ori_n528_), .D(ori_ori_n525_), .Y(ori_ori_n532_));
  NO4        o0504(.A(ori_ori_n532_), .B(ori_ori_n522_), .C(ori_ori_n518_), .D(ori_ori_n515_), .Y(ori_ori_n533_));
  NA4        o0505(.A(ori_ori_n533_), .B(ori_ori_n506_), .C(ori_ori_n475_), .D(ori_ori_n448_), .Y(ori11));
  NO2        o0506(.A(ori_ori_n71_), .B(f), .Y(ori_ori_n535_));
  NA2        o0507(.A(j), .B(g), .Y(ori_ori_n536_));
  NAi31      o0508(.An(i), .B(m), .C(l), .Y(ori_ori_n537_));
  NA3        o0509(.A(m), .B(k), .C(j), .Y(ori_ori_n538_));
  OAI220     o0510(.A0(ori_ori_n538_), .A1(ori_ori_n132_), .B0(ori_ori_n537_), .B1(ori_ori_n536_), .Y(ori_ori_n539_));
  NA2        o0511(.A(ori_ori_n539_), .B(ori_ori_n535_), .Y(ori_ori_n540_));
  NOi32      o0512(.An(e), .Bn(b), .C(f), .Y(ori_ori_n541_));
  NA2        o0513(.A(ori_ori_n46_), .B(j), .Y(ori_ori_n542_));
  NO2        o0514(.A(ori_ori_n542_), .B(ori_ori_n309_), .Y(ori_ori_n543_));
  NAi31      o0515(.An(d), .B(e), .C(a), .Y(ori_ori_n544_));
  NO2        o0516(.A(ori_ori_n544_), .B(n), .Y(ori_ori_n545_));
  AOI220     o0517(.A0(ori_ori_n545_), .A1(ori_ori_n101_), .B0(ori_ori_n543_), .B1(ori_ori_n541_), .Y(ori_ori_n546_));
  NAi41      o0518(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n547_));
  AN2        o0519(.A(ori_ori_n547_), .B(ori_ori_n386_), .Y(ori_ori_n548_));
  NA2        o0520(.A(j), .B(i), .Y(ori_ori_n549_));
  NAi31      o0521(.An(n), .B(m), .C(k), .Y(ori_ori_n550_));
  NO3        o0522(.A(ori_ori_n550_), .B(ori_ori_n549_), .C(ori_ori_n113_), .Y(ori_ori_n551_));
  NO4        o0523(.A(n), .B(d), .C(ori_ori_n117_), .D(a), .Y(ori_ori_n552_));
  OR2        o0524(.A(n), .B(c), .Y(ori_ori_n553_));
  NO2        o0525(.A(ori_ori_n553_), .B(ori_ori_n152_), .Y(ori_ori_n554_));
  NO2        o0526(.A(ori_ori_n554_), .B(ori_ori_n552_), .Y(ori_ori_n555_));
  NOi32      o0527(.An(g), .Bn(f), .C(i), .Y(ori_ori_n556_));
  NA2        o0528(.A(ori_ori_n539_), .B(f), .Y(ori_ori_n557_));
  NO2        o0529(.A(ori_ori_n283_), .B(ori_ori_n49_), .Y(ori_ori_n558_));
  NO2        o0530(.A(ori_ori_n557_), .B(ori_ori_n555_), .Y(ori_ori_n559_));
  INV        o0531(.A(ori_ori_n559_), .Y(ori_ori_n560_));
  NA2        o0532(.A(ori_ori_n142_), .B(ori_ori_n34_), .Y(ori_ori_n561_));
  OAI220     o0533(.A0(ori_ori_n561_), .A1(m), .B0(ori_ori_n542_), .B1(ori_ori_n239_), .Y(ori_ori_n562_));
  NOi41      o0534(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n563_));
  NAi32      o0535(.An(e), .Bn(b), .C(c), .Y(ori_ori_n564_));
  OR2        o0536(.A(ori_ori_n564_), .B(ori_ori_n83_), .Y(ori_ori_n565_));
  AN2        o0537(.A(ori_ori_n351_), .B(ori_ori_n329_), .Y(ori_ori_n566_));
  NA2        o0538(.A(ori_ori_n566_), .B(ori_ori_n565_), .Y(ori_ori_n567_));
  OA210      o0539(.A0(ori_ori_n567_), .A1(ori_ori_n563_), .B0(ori_ori_n562_), .Y(ori_ori_n568_));
  OAI220     o0540(.A0(ori_ori_n414_), .A1(ori_ori_n413_), .B0(ori_ori_n537_), .B1(ori_ori_n536_), .Y(ori_ori_n569_));
  NAi31      o0541(.An(d), .B(c), .C(a), .Y(ori_ori_n570_));
  NO2        o0542(.A(ori_ori_n570_), .B(n), .Y(ori_ori_n571_));
  NA3        o0543(.A(ori_ori_n571_), .B(ori_ori_n569_), .C(e), .Y(ori_ori_n572_));
  INV        o0544(.A(ori_ori_n572_), .Y(ori_ori_n573_));
  NO2        o0545(.A(ori_ori_n284_), .B(n), .Y(ori_ori_n574_));
  NO2        o0546(.A(ori_ori_n443_), .B(ori_ori_n574_), .Y(ori_ori_n575_));
  NA2        o0547(.A(ori_ori_n569_), .B(f), .Y(ori_ori_n576_));
  NAi32      o0548(.An(d), .Bn(a), .C(b), .Y(ori_ori_n577_));
  NO2        o0549(.A(ori_ori_n577_), .B(ori_ori_n49_), .Y(ori_ori_n578_));
  NA2        o0550(.A(h), .B(f), .Y(ori_ori_n579_));
  NO2        o0551(.A(ori_ori_n579_), .B(ori_ori_n94_), .Y(ori_ori_n580_));
  NO3        o0552(.A(ori_ori_n180_), .B(ori_ori_n177_), .C(g), .Y(ori_ori_n581_));
  AOI220     o0553(.A0(ori_ori_n581_), .A1(ori_ori_n58_), .B0(ori_ori_n580_), .B1(ori_ori_n578_), .Y(ori_ori_n582_));
  OAI210     o0554(.A0(ori_ori_n576_), .A1(ori_ori_n575_), .B0(ori_ori_n582_), .Y(ori_ori_n583_));
  AN3        o0555(.A(j), .B(h), .C(g), .Y(ori_ori_n584_));
  NO2        o0556(.A(ori_ori_n149_), .B(c), .Y(ori_ori_n585_));
  NA3        o0557(.A(ori_ori_n585_), .B(ori_ori_n584_), .C(ori_ori_n470_), .Y(ori_ori_n586_));
  NA3        o0558(.A(f), .B(d), .C(b), .Y(ori_ori_n587_));
  NO4        o0559(.A(ori_ori_n587_), .B(ori_ori_n180_), .C(ori_ori_n177_), .D(g), .Y(ori_ori_n588_));
  NAi21      o0560(.An(ori_ori_n588_), .B(ori_ori_n586_), .Y(ori_ori_n589_));
  NO4        o0561(.A(ori_ori_n589_), .B(ori_ori_n583_), .C(ori_ori_n573_), .D(ori_ori_n568_), .Y(ori_ori_n590_));
  AN4        o0562(.A(ori_ori_n590_), .B(ori_ori_n560_), .C(ori_ori_n546_), .D(ori_ori_n540_), .Y(ori_ori_n591_));
  INV        o0563(.A(k), .Y(ori_ori_n592_));
  NA3        o0564(.A(l), .B(ori_ori_n592_), .C(i), .Y(ori_ori_n593_));
  INV        o0565(.A(ori_ori_n593_), .Y(ori_ori_n594_));
  NAi32      o0566(.An(h), .Bn(f), .C(g), .Y(ori_ori_n595_));
  NAi41      o0567(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n596_));
  OAI210     o0568(.A0(ori_ori_n544_), .A1(n), .B0(ori_ori_n596_), .Y(ori_ori_n597_));
  NA2        o0569(.A(ori_ori_n597_), .B(m), .Y(ori_ori_n598_));
  NAi31      o0570(.An(h), .B(g), .C(f), .Y(ori_ori_n599_));
  OR3        o0571(.A(ori_ori_n599_), .B(ori_ori_n284_), .C(ori_ori_n49_), .Y(ori_ori_n600_));
  NA4        o0572(.A(ori_ori_n432_), .B(ori_ori_n122_), .C(ori_ori_n114_), .D(e), .Y(ori_ori_n601_));
  AN2        o0573(.A(ori_ori_n601_), .B(ori_ori_n600_), .Y(ori_ori_n602_));
  OA210      o0574(.A0(ori_ori_n598_), .A1(ori_ori_n595_), .B0(ori_ori_n602_), .Y(ori_ori_n603_));
  NO3        o0575(.A(ori_ori_n595_), .B(ori_ori_n71_), .C(ori_ori_n72_), .Y(ori_ori_n604_));
  NO4        o0576(.A(ori_ori_n599_), .B(ori_ori_n553_), .C(ori_ori_n152_), .D(ori_ori_n72_), .Y(ori_ori_n605_));
  OR2        o0577(.A(ori_ori_n605_), .B(ori_ori_n604_), .Y(ori_ori_n606_));
  NAi21      o0578(.An(ori_ori_n606_), .B(ori_ori_n603_), .Y(ori_ori_n607_));
  NAi31      o0579(.An(f), .B(h), .C(g), .Y(ori_ori_n608_));
  NO4        o0580(.A(ori_ori_n320_), .B(ori_ori_n608_), .C(ori_ori_n71_), .D(ori_ori_n72_), .Y(ori_ori_n609_));
  NOi32      o0581(.An(b), .Bn(a), .C(c), .Y(ori_ori_n610_));
  NOi41      o0582(.An(ori_ori_n610_), .B(ori_ori_n366_), .C(ori_ori_n69_), .D(ori_ori_n118_), .Y(ori_ori_n611_));
  OR2        o0583(.A(ori_ori_n611_), .B(ori_ori_n609_), .Y(ori_ori_n612_));
  NOi32      o0584(.An(d), .Bn(a), .C(e), .Y(ori_ori_n613_));
  NA2        o0585(.A(ori_ori_n613_), .B(ori_ori_n114_), .Y(ori_ori_n614_));
  NO2        o0586(.A(n), .B(c), .Y(ori_ori_n615_));
  NA3        o0587(.A(ori_ori_n615_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n616_));
  NAi32      o0588(.An(n), .Bn(f), .C(m), .Y(ori_ori_n617_));
  NA3        o0589(.A(ori_ori_n617_), .B(ori_ori_n616_), .C(ori_ori_n614_), .Y(ori_ori_n618_));
  NOi32      o0590(.An(e), .Bn(a), .C(d), .Y(ori_ori_n619_));
  AOI210     o0591(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n619_), .Y(ori_ori_n620_));
  AOI210     o0592(.A0(ori_ori_n620_), .A1(ori_ori_n218_), .B0(ori_ori_n561_), .Y(ori_ori_n621_));
  AOI210     o0593(.A0(ori_ori_n621_), .A1(ori_ori_n618_), .B0(ori_ori_n612_), .Y(ori_ori_n622_));
  OAI210     o0594(.A0(ori_ori_n255_), .A1(ori_ori_n86_), .B0(ori_ori_n622_), .Y(ori_ori_n623_));
  AOI210     o0595(.A0(ori_ori_n607_), .A1(ori_ori_n594_), .B0(ori_ori_n623_), .Y(ori_ori_n624_));
  NO3        o0596(.A(ori_ori_n327_), .B(ori_ori_n61_), .C(n), .Y(ori_ori_n625_));
  NA3        o0597(.A(ori_ori_n523_), .B(ori_ori_n175_), .C(ori_ori_n174_), .Y(ori_ori_n626_));
  NA2        o0598(.A(ori_ori_n472_), .B(ori_ori_n236_), .Y(ori_ori_n627_));
  OR2        o0599(.A(ori_ori_n627_), .B(ori_ori_n626_), .Y(ori_ori_n628_));
  NA2        o0600(.A(ori_ori_n628_), .B(ori_ori_n625_), .Y(ori_ori_n629_));
  NO2        o0601(.A(ori_ori_n629_), .B(ori_ori_n86_), .Y(ori_ori_n630_));
  NA3        o0602(.A(ori_ori_n563_), .B(ori_ori_n353_), .C(ori_ori_n46_), .Y(ori_ori_n631_));
  NOi32      o0603(.An(e), .Bn(c), .C(f), .Y(ori_ori_n632_));
  NOi21      o0604(.An(f), .B(g), .Y(ori_ori_n633_));
  NO2        o0605(.A(ori_ori_n633_), .B(ori_ori_n216_), .Y(ori_ori_n634_));
  AOI220     o0606(.A0(ori_ori_n634_), .A1(ori_ori_n408_), .B0(ori_ori_n632_), .B1(ori_ori_n179_), .Y(ori_ori_n635_));
  NA3        o0607(.A(ori_ori_n635_), .B(ori_ori_n631_), .C(ori_ori_n182_), .Y(ori_ori_n636_));
  AOI210     o0608(.A0(ori_ori_n548_), .A1(ori_ori_n412_), .B0(ori_ori_n308_), .Y(ori_ori_n637_));
  NA2        o0609(.A(ori_ori_n637_), .B(ori_ori_n272_), .Y(ori_ori_n638_));
  NOi21      o0610(.An(j), .B(l), .Y(ori_ori_n639_));
  NAi21      o0611(.An(k), .B(h), .Y(ori_ori_n640_));
  NO2        o0612(.A(ori_ori_n640_), .B(ori_ori_n270_), .Y(ori_ori_n641_));
  NA2        o0613(.A(ori_ori_n641_), .B(ori_ori_n639_), .Y(ori_ori_n642_));
  OR2        o0614(.A(ori_ori_n642_), .B(ori_ori_n598_), .Y(ori_ori_n643_));
  NOi31      o0615(.An(m), .B(n), .C(k), .Y(ori_ori_n644_));
  NA2        o0616(.A(ori_ori_n639_), .B(ori_ori_n644_), .Y(ori_ori_n645_));
  AOI210     o0617(.A0(ori_ori_n412_), .A1(ori_ori_n386_), .B0(ori_ori_n308_), .Y(ori_ori_n646_));
  NAi21      o0618(.An(ori_ori_n645_), .B(ori_ori_n646_), .Y(ori_ori_n647_));
  NO2        o0619(.A(ori_ori_n284_), .B(ori_ori_n49_), .Y(ori_ori_n648_));
  NO2        o0620(.A(ori_ori_n320_), .B(ori_ori_n608_), .Y(ori_ori_n649_));
  NO2        o0621(.A(ori_ori_n544_), .B(ori_ori_n49_), .Y(ori_ori_n650_));
  AOI220     o0622(.A0(ori_ori_n650_), .A1(ori_ori_n649_), .B0(ori_ori_n648_), .B1(ori_ori_n580_), .Y(ori_ori_n651_));
  NA4        o0623(.A(ori_ori_n651_), .B(ori_ori_n647_), .C(ori_ori_n643_), .D(ori_ori_n638_), .Y(ori_ori_n652_));
  NA2        o0624(.A(ori_ori_n109_), .B(ori_ori_n36_), .Y(ori_ori_n653_));
  NO2        o0625(.A(k), .B(ori_ori_n219_), .Y(ori_ori_n654_));
  INV        o0626(.A(ori_ori_n375_), .Y(ori_ori_n655_));
  NO2        o0627(.A(ori_ori_n655_), .B(n), .Y(ori_ori_n656_));
  NAi31      o0628(.An(ori_ori_n653_), .B(ori_ori_n656_), .C(ori_ori_n654_), .Y(ori_ori_n657_));
  NO2        o0629(.A(ori_ori_n542_), .B(ori_ori_n180_), .Y(ori_ori_n658_));
  NA3        o0630(.A(ori_ori_n564_), .B(ori_ori_n279_), .C(ori_ori_n147_), .Y(ori_ori_n659_));
  NA2        o0631(.A(ori_ori_n519_), .B(ori_ori_n163_), .Y(ori_ori_n660_));
  NO3        o0632(.A(ori_ori_n409_), .B(ori_ori_n660_), .C(ori_ori_n86_), .Y(ori_ori_n661_));
  AOI210     o0633(.A0(ori_ori_n659_), .A1(ori_ori_n658_), .B0(ori_ori_n661_), .Y(ori_ori_n662_));
  AN3        o0634(.A(f), .B(d), .C(b), .Y(ori_ori_n663_));
  OAI210     o0635(.A0(ori_ori_n663_), .A1(ori_ori_n131_), .B0(n), .Y(ori_ori_n664_));
  NA3        o0636(.A(ori_ori_n519_), .B(ori_ori_n163_), .C(ori_ori_n219_), .Y(ori_ori_n665_));
  AOI210     o0637(.A0(ori_ori_n664_), .A1(ori_ori_n238_), .B0(ori_ori_n665_), .Y(ori_ori_n666_));
  NAi31      o0638(.An(m), .B(n), .C(k), .Y(ori_ori_n667_));
  OR2        o0639(.A(ori_ori_n136_), .B(ori_ori_n61_), .Y(ori_ori_n668_));
  OAI210     o0640(.A0(ori_ori_n668_), .A1(ori_ori_n667_), .B0(ori_ori_n257_), .Y(ori_ori_n669_));
  OAI210     o0641(.A0(ori_ori_n669_), .A1(ori_ori_n666_), .B0(j), .Y(ori_ori_n670_));
  NA3        o0642(.A(ori_ori_n670_), .B(ori_ori_n662_), .C(ori_ori_n657_), .Y(ori_ori_n671_));
  NO4        o0643(.A(ori_ori_n671_), .B(ori_ori_n652_), .C(ori_ori_n636_), .D(ori_ori_n630_), .Y(ori_ori_n672_));
  NA2        o0644(.A(ori_ori_n396_), .B(ori_ori_n166_), .Y(ori_ori_n673_));
  NAi31      o0645(.An(g), .B(h), .C(f), .Y(ori_ori_n674_));
  OR3        o0646(.A(ori_ori_n674_), .B(ori_ori_n284_), .C(n), .Y(ori_ori_n675_));
  OA210      o0647(.A0(ori_ori_n544_), .A1(n), .B0(ori_ori_n596_), .Y(ori_ori_n676_));
  NA3        o0648(.A(ori_ori_n430_), .B(ori_ori_n122_), .C(ori_ori_n83_), .Y(ori_ori_n677_));
  OAI210     o0649(.A0(ori_ori_n676_), .A1(ori_ori_n90_), .B0(ori_ori_n677_), .Y(ori_ori_n678_));
  NOi21      o0650(.An(ori_ori_n675_), .B(ori_ori_n678_), .Y(ori_ori_n679_));
  AOI210     o0651(.A0(ori_ori_n679_), .A1(ori_ori_n673_), .B0(ori_ori_n538_), .Y(ori_ori_n680_));
  NO3        o0652(.A(g), .B(ori_ori_n218_), .C(ori_ori_n56_), .Y(ori_ori_n681_));
  NAi21      o0653(.An(h), .B(j), .Y(ori_ori_n682_));
  NO2        o0654(.A(ori_ori_n526_), .B(ori_ori_n86_), .Y(ori_ori_n683_));
  OAI210     o0655(.A0(ori_ori_n683_), .A1(ori_ori_n408_), .B0(ori_ori_n681_), .Y(ori_ori_n684_));
  OR2        o0656(.A(ori_ori_n71_), .B(ori_ori_n72_), .Y(ori_ori_n685_));
  NA2        o0657(.A(ori_ori_n610_), .B(ori_ori_n355_), .Y(ori_ori_n686_));
  OA220      o0658(.A0(ori_ori_n645_), .A1(ori_ori_n686_), .B0(ori_ori_n642_), .B1(ori_ori_n685_), .Y(ori_ori_n687_));
  NA3        o0659(.A(ori_ori_n535_), .B(ori_ori_n99_), .C(ori_ori_n98_), .Y(ori_ori_n688_));
  AN2        o0660(.A(h), .B(f), .Y(ori_ori_n689_));
  NA2        o0661(.A(ori_ori_n689_), .B(ori_ori_n37_), .Y(ori_ori_n690_));
  NA2        o0662(.A(ori_ori_n99_), .B(ori_ori_n46_), .Y(ori_ori_n691_));
  OAI220     o0663(.A0(ori_ori_n691_), .A1(ori_ori_n344_), .B0(ori_ori_n690_), .B1(ori_ori_n477_), .Y(ori_ori_n692_));
  AOI210     o0664(.A0(ori_ori_n577_), .A1(ori_ori_n442_), .B0(ori_ori_n49_), .Y(ori_ori_n693_));
  OAI220     o0665(.A0(ori_ori_n599_), .A1(ori_ori_n593_), .B0(ori_ori_n337_), .B1(ori_ori_n536_), .Y(ori_ori_n694_));
  AOI210     o0666(.A0(ori_ori_n694_), .A1(ori_ori_n693_), .B0(ori_ori_n692_), .Y(ori_ori_n695_));
  NA4        o0667(.A(ori_ori_n695_), .B(ori_ori_n688_), .C(ori_ori_n687_), .D(ori_ori_n684_), .Y(ori_ori_n696_));
  NO2        o0668(.A(ori_ori_n633_), .B(ori_ori_n61_), .Y(ori_ori_n697_));
  NO2        o0669(.A(ori_ori_n697_), .B(ori_ori_n34_), .Y(ori_ori_n698_));
  NA2        o0670(.A(ori_ori_n340_), .B(ori_ori_n142_), .Y(ori_ori_n699_));
  NA2        o0671(.A(ori_ori_n133_), .B(ori_ori_n49_), .Y(ori_ori_n700_));
  AOI220     o0672(.A0(ori_ori_n700_), .A1(ori_ori_n541_), .B0(ori_ori_n375_), .B1(ori_ori_n114_), .Y(ori_ori_n701_));
  OA220      o0673(.A0(ori_ori_n701_), .A1(ori_ori_n561_), .B0(ori_ori_n373_), .B1(ori_ori_n112_), .Y(ori_ori_n702_));
  OAI210     o0674(.A0(ori_ori_n699_), .A1(ori_ori_n698_), .B0(ori_ori_n702_), .Y(ori_ori_n703_));
  NO3        o0675(.A(ori_ori_n417_), .B(ori_ori_n196_), .C(ori_ori_n195_), .Y(ori_ori_n704_));
  NA2        o0676(.A(ori_ori_n704_), .B(ori_ori_n236_), .Y(ori_ori_n705_));
  NA3        o0677(.A(ori_ori_n705_), .B(ori_ori_n261_), .C(j), .Y(ori_ori_n706_));
  NO3        o0678(.A(ori_ori_n472_), .B(ori_ori_n177_), .C(i), .Y(ori_ori_n707_));
  NA2        o0679(.A(ori_ori_n476_), .B(ori_ori_n83_), .Y(ori_ori_n708_));
  NA2        o0680(.A(ori_ori_n706_), .B(ori_ori_n415_), .Y(ori_ori_n709_));
  NO4        o0681(.A(ori_ori_n709_), .B(ori_ori_n703_), .C(ori_ori_n696_), .D(ori_ori_n680_), .Y(ori_ori_n710_));
  NA4        o0682(.A(ori_ori_n710_), .B(ori_ori_n672_), .C(ori_ori_n624_), .D(ori_ori_n591_), .Y(ori08));
  NO2        o0683(.A(k), .B(h), .Y(ori_ori_n712_));
  AO210      o0684(.A0(ori_ori_n259_), .A1(ori_ori_n460_), .B0(ori_ori_n712_), .Y(ori_ori_n713_));
  NO2        o0685(.A(ori_ori_n713_), .B(ori_ori_n306_), .Y(ori_ori_n714_));
  NA2        o0686(.A(ori_ori_n632_), .B(ori_ori_n83_), .Y(ori_ori_n715_));
  NA2        o0687(.A(ori_ori_n715_), .B(ori_ori_n472_), .Y(ori_ori_n716_));
  AOI210     o0688(.A0(ori_ori_n716_), .A1(ori_ori_n714_), .B0(ori_ori_n503_), .Y(ori_ori_n717_));
  NA2        o0689(.A(ori_ori_n83_), .B(ori_ori_n111_), .Y(ori_ori_n718_));
  NO2        o0690(.A(ori_ori_n718_), .B(ori_ori_n57_), .Y(ori_ori_n719_));
  NO4        o0691(.A(ori_ori_n393_), .B(ori_ori_n113_), .C(j), .D(ori_ori_n219_), .Y(ori_ori_n720_));
  NA2        o0692(.A(ori_ori_n587_), .B(ori_ori_n238_), .Y(ori_ori_n721_));
  AOI220     o0693(.A0(ori_ori_n721_), .A1(ori_ori_n360_), .B0(ori_ori_n720_), .B1(ori_ori_n719_), .Y(ori_ori_n722_));
  AOI210     o0694(.A0(ori_ori_n587_), .A1(ori_ori_n159_), .B0(ori_ori_n83_), .Y(ori_ori_n723_));
  NA4        o0695(.A(ori_ori_n221_), .B(ori_ori_n142_), .C(ori_ori_n45_), .D(h), .Y(ori_ori_n724_));
  AN2        o0696(.A(l), .B(k), .Y(ori_ori_n725_));
  NA4        o0697(.A(ori_ori_n725_), .B(ori_ori_n109_), .C(ori_ori_n72_), .D(ori_ori_n219_), .Y(ori_ori_n726_));
  OAI210     o0698(.A0(ori_ori_n724_), .A1(g), .B0(ori_ori_n726_), .Y(ori_ori_n727_));
  NA2        o0699(.A(ori_ori_n727_), .B(ori_ori_n723_), .Y(ori_ori_n728_));
  NA4        o0700(.A(ori_ori_n728_), .B(ori_ori_n722_), .C(ori_ori_n717_), .D(ori_ori_n362_), .Y(ori_ori_n729_));
  AN2        o0701(.A(ori_ori_n545_), .B(ori_ori_n95_), .Y(ori_ori_n730_));
  NO4        o0702(.A(ori_ori_n177_), .B(ori_ori_n407_), .C(ori_ori_n113_), .D(g), .Y(ori_ori_n731_));
  NA2        o0703(.A(ori_ori_n731_), .B(ori_ori_n721_), .Y(ori_ori_n732_));
  NO2        o0704(.A(ori_ori_n38_), .B(ori_ori_n218_), .Y(ori_ori_n733_));
  AOI220     o0705(.A0(ori_ori_n634_), .A1(ori_ori_n359_), .B0(ori_ori_n733_), .B1(ori_ori_n574_), .Y(ori_ori_n734_));
  NAi31      o0706(.An(ori_ori_n730_), .B(ori_ori_n734_), .C(ori_ori_n732_), .Y(ori_ori_n735_));
  NO2        o0707(.A(ori_ori_n548_), .B(ori_ori_n35_), .Y(ori_ori_n736_));
  OAI210     o0708(.A0(ori_ori_n564_), .A1(ori_ori_n47_), .B0(ori_ori_n668_), .Y(ori_ori_n737_));
  NO2        o0709(.A(ori_ori_n497_), .B(ori_ori_n133_), .Y(ori_ori_n738_));
  AOI210     o0710(.A0(ori_ori_n738_), .A1(ori_ori_n737_), .B0(ori_ori_n736_), .Y(ori_ori_n739_));
  NO3        o0711(.A(ori_ori_n327_), .B(ori_ori_n132_), .C(ori_ori_n41_), .Y(ori_ori_n740_));
  NAi21      o0712(.An(ori_ori_n740_), .B(ori_ori_n726_), .Y(ori_ori_n741_));
  NA2        o0713(.A(ori_ori_n713_), .B(ori_ori_n137_), .Y(ori_ori_n742_));
  AOI220     o0714(.A0(ori_ori_n742_), .A1(ori_ori_n416_), .B0(ori_ori_n741_), .B1(ori_ori_n75_), .Y(ori_ori_n743_));
  OAI210     o0715(.A0(ori_ori_n739_), .A1(ori_ori_n86_), .B0(ori_ori_n743_), .Y(ori_ori_n744_));
  NA2        o0716(.A(ori_ori_n375_), .B(ori_ori_n43_), .Y(ori_ori_n745_));
  NA3        o0717(.A(ori_ori_n705_), .B(ori_ori_n346_), .C(ori_ori_n399_), .Y(ori_ori_n746_));
  NA3        o0718(.A(m), .B(l), .C(k), .Y(ori_ori_n747_));
  AOI210     o0719(.A0(ori_ori_n677_), .A1(ori_ori_n675_), .B0(ori_ori_n747_), .Y(ori_ori_n748_));
  NA3        o0720(.A(ori_ori_n114_), .B(k), .C(ori_ori_n86_), .Y(ori_ori_n749_));
  INV        o0721(.A(ori_ori_n748_), .Y(ori_ori_n750_));
  NA3        o0722(.A(ori_ori_n750_), .B(ori_ori_n746_), .C(ori_ori_n745_), .Y(ori_ori_n751_));
  NO4        o0723(.A(ori_ori_n751_), .B(ori_ori_n744_), .C(ori_ori_n735_), .D(ori_ori_n729_), .Y(ori_ori_n752_));
  NA2        o0724(.A(ori_ori_n634_), .B(ori_ori_n408_), .Y(ori_ori_n753_));
  NOi31      o0725(.An(g), .B(h), .C(f), .Y(ori_ori_n754_));
  NA2        o0726(.A(ori_ori_n650_), .B(ori_ori_n754_), .Y(ori_ori_n755_));
  AO210      o0727(.A0(ori_ori_n755_), .A1(ori_ori_n600_), .B0(ori_ori_n549_), .Y(ori_ori_n756_));
  INV        o0728(.A(ori_ori_n513_), .Y(ori_ori_n757_));
  NA4        o0729(.A(ori_ori_n757_), .B(ori_ori_n756_), .C(ori_ori_n753_), .D(ori_ori_n258_), .Y(ori_ori_n758_));
  NA2        o0730(.A(ori_ori_n725_), .B(ori_ori_n72_), .Y(ori_ori_n759_));
  NO4        o0731(.A(ori_ori_n704_), .B(ori_ori_n177_), .C(n), .D(i), .Y(ori_ori_n760_));
  NOi21      o0732(.An(h), .B(j), .Y(ori_ori_n761_));
  NA2        o0733(.A(ori_ori_n761_), .B(f), .Y(ori_ori_n762_));
  NO2        o0734(.A(ori_ori_n762_), .B(ori_ori_n252_), .Y(ori_ori_n763_));
  NO3        o0735(.A(ori_ori_n763_), .B(ori_ori_n760_), .C(ori_ori_n707_), .Y(ori_ori_n764_));
  OAI220     o0736(.A0(ori_ori_n764_), .A1(ori_ori_n759_), .B0(ori_ori_n602_), .B1(ori_ori_n62_), .Y(ori_ori_n765_));
  AOI210     o0737(.A0(ori_ori_n758_), .A1(l), .B0(ori_ori_n765_), .Y(ori_ori_n766_));
  NO2        o0738(.A(j), .B(i), .Y(ori_ori_n767_));
  NA3        o0739(.A(ori_ori_n767_), .B(ori_ori_n79_), .C(l), .Y(ori_ori_n768_));
  NA2        o0740(.A(ori_ori_n767_), .B(ori_ori_n33_), .Y(ori_ori_n769_));
  NA2        o0741(.A(ori_ori_n435_), .B(ori_ori_n122_), .Y(ori_ori_n770_));
  OA220      o0742(.A0(ori_ori_n770_), .A1(ori_ori_n769_), .B0(ori_ori_n768_), .B1(ori_ori_n598_), .Y(ori_ori_n771_));
  NO3        o0743(.A(ori_ori_n154_), .B(ori_ori_n49_), .C(ori_ori_n111_), .Y(ori_ori_n772_));
  NO3        o0744(.A(ori_ori_n553_), .B(ori_ori_n152_), .C(ori_ori_n72_), .Y(ori_ori_n773_));
  NO3        o0745(.A(ori_ori_n497_), .B(ori_ori_n451_), .C(j), .Y(ori_ori_n774_));
  OAI210     o0746(.A0(ori_ori_n773_), .A1(ori_ori_n772_), .B0(ori_ori_n774_), .Y(ori_ori_n775_));
  OAI210     o0747(.A0(ori_ori_n755_), .A1(ori_ori_n62_), .B0(ori_ori_n775_), .Y(ori_ori_n776_));
  NA2        o0748(.A(k), .B(j), .Y(ori_ori_n777_));
  NO3        o0749(.A(ori_ori_n306_), .B(ori_ori_n777_), .C(ori_ori_n40_), .Y(ori_ori_n778_));
  AOI210     o0750(.A0(ori_ori_n541_), .A1(n), .B0(ori_ori_n563_), .Y(ori_ori_n779_));
  NA2        o0751(.A(ori_ori_n779_), .B(ori_ori_n566_), .Y(ori_ori_n780_));
  AN3        o0752(.A(ori_ori_n780_), .B(ori_ori_n778_), .C(ori_ori_n98_), .Y(ori_ori_n781_));
  NO3        o0753(.A(ori_ori_n177_), .B(ori_ori_n407_), .C(ori_ori_n113_), .Y(ori_ori_n782_));
  AOI220     o0754(.A0(ori_ori_n782_), .A1(ori_ori_n253_), .B0(ori_ori_n627_), .B1(ori_ori_n317_), .Y(ori_ori_n783_));
  INV        o0755(.A(ori_ori_n783_), .Y(ori_ori_n784_));
  NO2        o0756(.A(ori_ori_n306_), .B(ori_ori_n137_), .Y(ori_ori_n785_));
  AOI220     o0757(.A0(ori_ori_n785_), .A1(ori_ori_n634_), .B0(ori_ori_n740_), .B1(ori_ori_n723_), .Y(ori_ori_n786_));
  NO2        o0758(.A(ori_ori_n747_), .B(ori_ori_n90_), .Y(ori_ori_n787_));
  NA2        o0759(.A(ori_ori_n787_), .B(ori_ori_n597_), .Y(ori_ori_n788_));
  NO2        o0760(.A(ori_ori_n599_), .B(ori_ori_n118_), .Y(ori_ori_n789_));
  OAI210     o0761(.A0(ori_ori_n789_), .A1(ori_ori_n774_), .B0(ori_ori_n693_), .Y(ori_ori_n790_));
  NA3        o0762(.A(ori_ori_n790_), .B(ori_ori_n788_), .C(ori_ori_n786_), .Y(ori_ori_n791_));
  OR4        o0763(.A(ori_ori_n791_), .B(ori_ori_n784_), .C(ori_ori_n781_), .D(ori_ori_n776_), .Y(ori_ori_n792_));
  NA3        o0764(.A(ori_ori_n779_), .B(ori_ori_n566_), .C(ori_ori_n565_), .Y(ori_ori_n793_));
  NA4        o0765(.A(ori_ori_n793_), .B(ori_ori_n221_), .C(ori_ori_n460_), .D(ori_ori_n34_), .Y(ori_ori_n794_));
  NO4        o0766(.A(ori_ori_n497_), .B(ori_ori_n449_), .C(j), .D(f), .Y(ori_ori_n795_));
  OAI220     o0767(.A0(ori_ori_n724_), .A1(ori_ori_n715_), .B0(ori_ori_n344_), .B1(ori_ori_n38_), .Y(ori_ori_n796_));
  AOI210     o0768(.A0(ori_ori_n795_), .A1(ori_ori_n265_), .B0(ori_ori_n796_), .Y(ori_ori_n797_));
  NA3        o0769(.A(ori_ori_n556_), .B(ori_ori_n299_), .C(h), .Y(ori_ori_n798_));
  NO2        o0770(.A(ori_ori_n91_), .B(ori_ori_n47_), .Y(ori_ori_n799_));
  OAI220     o0771(.A0(ori_ori_n798_), .A1(ori_ori_n616_), .B0(ori_ori_n768_), .B1(ori_ori_n685_), .Y(ori_ori_n800_));
  AOI210     o0772(.A0(ori_ori_n799_), .A1(ori_ori_n656_), .B0(ori_ori_n800_), .Y(ori_ori_n801_));
  NA3        o0773(.A(ori_ori_n801_), .B(ori_ori_n797_), .C(ori_ori_n794_), .Y(ori_ori_n802_));
  OR2        o0774(.A(ori_ori_n787_), .B(ori_ori_n95_), .Y(ori_ori_n803_));
  AOI220     o0775(.A0(ori_ori_n803_), .A1(ori_ori_n244_), .B0(ori_ori_n774_), .B1(ori_ori_n648_), .Y(ori_ori_n804_));
  NO2        o0776(.A(ori_ori_n676_), .B(ori_ori_n72_), .Y(ori_ori_n805_));
  AOI210     o0777(.A0(ori_ori_n795_), .A1(ori_ori_n805_), .B0(ori_ori_n348_), .Y(ori_ori_n806_));
  OAI210     o0778(.A0(ori_ori_n747_), .A1(ori_ori_n674_), .B0(ori_ori_n530_), .Y(ori_ori_n807_));
  NA3        o0779(.A(ori_ori_n256_), .B(ori_ori_n59_), .C(b), .Y(ori_ori_n808_));
  AOI220     o0780(.A0(ori_ori_n615_), .A1(ori_ori_n29_), .B0(ori_ori_n476_), .B1(ori_ori_n83_), .Y(ori_ori_n809_));
  NA2        o0781(.A(ori_ori_n809_), .B(ori_ori_n808_), .Y(ori_ori_n810_));
  NA2        o0782(.A(ori_ori_n810_), .B(ori_ori_n807_), .Y(ori_ori_n811_));
  NA3        o0783(.A(ori_ori_n811_), .B(ori_ori_n806_), .C(ori_ori_n804_), .Y(ori_ori_n812_));
  NOi41      o0784(.An(ori_ori_n771_), .B(ori_ori_n812_), .C(ori_ori_n802_), .D(ori_ori_n792_), .Y(ori_ori_n813_));
  OR3        o0785(.A(ori_ori_n724_), .B(ori_ori_n238_), .C(g), .Y(ori_ori_n814_));
  NO3        o0786(.A(ori_ori_n354_), .B(ori_ori_n308_), .C(ori_ori_n113_), .Y(ori_ori_n815_));
  NA2        o0787(.A(ori_ori_n815_), .B(ori_ori_n780_), .Y(ori_ori_n816_));
  NA2        o0788(.A(ori_ori_n46_), .B(ori_ori_n56_), .Y(ori_ori_n817_));
  NO3        o0789(.A(ori_ori_n817_), .B(ori_ori_n769_), .C(ori_ori_n284_), .Y(ori_ori_n818_));
  NO3        o0790(.A(ori_ori_n536_), .B(ori_ori_n93_), .C(h), .Y(ori_ori_n819_));
  AOI210     o0791(.A0(ori_ori_n819_), .A1(ori_ori_n719_), .B0(ori_ori_n818_), .Y(ori_ori_n820_));
  NA4        o0792(.A(ori_ori_n820_), .B(ori_ori_n816_), .C(ori_ori_n814_), .D(ori_ori_n418_), .Y(ori_ori_n821_));
  OR2        o0793(.A(ori_ori_n674_), .B(ori_ori_n91_), .Y(ori_ori_n822_));
  NOi31      o0794(.An(b), .B(d), .C(a), .Y(ori_ori_n823_));
  NO2        o0795(.A(ori_ori_n823_), .B(ori_ori_n613_), .Y(ori_ori_n824_));
  NO2        o0796(.A(ori_ori_n824_), .B(n), .Y(ori_ori_n825_));
  NOi21      o0797(.An(ori_ori_n809_), .B(ori_ori_n825_), .Y(ori_ori_n826_));
  OAI220     o0798(.A0(ori_ori_n826_), .A1(ori_ori_n822_), .B0(ori_ori_n798_), .B1(ori_ori_n614_), .Y(ori_ori_n827_));
  NO2        o0799(.A(ori_ori_n564_), .B(ori_ori_n83_), .Y(ori_ori_n828_));
  NO3        o0800(.A(ori_ori_n633_), .B(ori_ori_n339_), .C(ori_ori_n118_), .Y(ori_ori_n829_));
  NOi21      o0801(.An(ori_ori_n829_), .B(ori_ori_n164_), .Y(ori_ori_n830_));
  AOI210     o0802(.A0(ori_ori_n815_), .A1(ori_ori_n828_), .B0(ori_ori_n830_), .Y(ori_ori_n831_));
  OAI210     o0803(.A0(ori_ori_n724_), .A1(ori_ori_n409_), .B0(ori_ori_n831_), .Y(ori_ori_n832_));
  NO2        o0804(.A(ori_ori_n704_), .B(n), .Y(ori_ori_n833_));
  AOI220     o0805(.A0(ori_ori_n785_), .A1(ori_ori_n681_), .B0(ori_ori_n833_), .B1(ori_ori_n714_), .Y(ori_ori_n834_));
  NO2        o0806(.A(ori_ori_n334_), .B(ori_ori_n243_), .Y(ori_ori_n835_));
  OAI210     o0807(.A0(ori_ori_n95_), .A1(ori_ori_n92_), .B0(ori_ori_n835_), .Y(ori_ori_n836_));
  NA2        o0808(.A(ori_ori_n122_), .B(ori_ori_n83_), .Y(ori_ori_n837_));
  AOI210     o0809(.A0(ori_ori_n439_), .A1(ori_ori_n431_), .B0(ori_ori_n837_), .Y(ori_ori_n838_));
  NAi21      o0810(.An(ori_ori_n838_), .B(ori_ori_n836_), .Y(ori_ori_n839_));
  OAI210     o0811(.A0(ori_ori_n605_), .A1(ori_ori_n604_), .B0(ori_ori_n376_), .Y(ori_ori_n840_));
  NAi31      o0812(.An(ori_ori_n839_), .B(ori_ori_n840_), .C(ori_ori_n834_), .Y(ori_ori_n841_));
  NO4        o0813(.A(ori_ori_n841_), .B(ori_ori_n832_), .C(ori_ori_n827_), .D(ori_ori_n821_), .Y(ori_ori_n842_));
  NA4        o0814(.A(ori_ori_n842_), .B(ori_ori_n813_), .C(ori_ori_n766_), .D(ori_ori_n752_), .Y(ori09));
  INV        o0815(.A(ori_ori_n123_), .Y(ori_ori_n844_));
  NA2        o0816(.A(f), .B(e), .Y(ori_ori_n845_));
  NO2        o0817(.A(ori_ori_n231_), .B(ori_ori_n113_), .Y(ori_ori_n846_));
  NA2        o0818(.A(ori_ori_n846_), .B(g), .Y(ori_ori_n847_));
  NA4        o0819(.A(ori_ori_n320_), .B(ori_ori_n168_), .C(ori_ori_n268_), .D(ori_ori_n120_), .Y(ori_ori_n848_));
  AOI210     o0820(.A0(ori_ori_n848_), .A1(g), .B0(ori_ori_n482_), .Y(ori_ori_n849_));
  AOI210     o0821(.A0(ori_ori_n849_), .A1(ori_ori_n847_), .B0(ori_ori_n845_), .Y(ori_ori_n850_));
  NA2        o0822(.A(ori_ori_n453_), .B(e), .Y(ori_ori_n851_));
  NO2        o0823(.A(ori_ori_n851_), .B(ori_ori_n523_), .Y(ori_ori_n852_));
  AOI210     o0824(.A0(ori_ori_n850_), .A1(ori_ori_n844_), .B0(ori_ori_n852_), .Y(ori_ori_n853_));
  NO2        o0825(.A(ori_ori_n208_), .B(ori_ori_n218_), .Y(ori_ori_n854_));
  NA3        o0826(.A(m), .B(l), .C(i), .Y(ori_ori_n855_));
  OAI220     o0827(.A0(ori_ori_n599_), .A1(ori_ori_n855_), .B0(ori_ori_n366_), .B1(ori_ori_n537_), .Y(ori_ori_n856_));
  NA4        o0828(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(g), .D(f), .Y(ori_ori_n857_));
  NAi21      o0829(.An(ori_ori_n856_), .B(ori_ori_n857_), .Y(ori_ori_n858_));
  OR2        o0830(.A(ori_ori_n858_), .B(ori_ori_n854_), .Y(ori_ori_n859_));
  NA3        o0831(.A(ori_ori_n822_), .B(ori_ori_n576_), .C(ori_ori_n530_), .Y(ori_ori_n860_));
  OA210      o0832(.A0(ori_ori_n860_), .A1(ori_ori_n859_), .B0(ori_ori_n825_), .Y(ori_ori_n861_));
  INV        o0833(.A(ori_ori_n351_), .Y(ori_ori_n862_));
  NO2        o0834(.A(ori_ori_n128_), .B(ori_ori_n126_), .Y(ori_ori_n863_));
  NOi31      o0835(.An(k), .B(m), .C(l), .Y(ori_ori_n864_));
  NO2        o0836(.A(ori_ori_n353_), .B(ori_ori_n864_), .Y(ori_ori_n865_));
  AOI210     o0837(.A0(ori_ori_n865_), .A1(ori_ori_n863_), .B0(ori_ori_n608_), .Y(ori_ori_n866_));
  NA2        o0838(.A(ori_ori_n808_), .B(ori_ori_n344_), .Y(ori_ori_n867_));
  NA2        o0839(.A(ori_ori_n355_), .B(ori_ori_n357_), .Y(ori_ori_n868_));
  OAI210     o0840(.A0(ori_ori_n208_), .A1(ori_ori_n218_), .B0(ori_ori_n868_), .Y(ori_ori_n869_));
  AOI220     o0841(.A0(ori_ori_n869_), .A1(ori_ori_n867_), .B0(ori_ori_n866_), .B1(ori_ori_n862_), .Y(ori_ori_n870_));
  NA2        o0842(.A(ori_ori_n172_), .B(ori_ori_n115_), .Y(ori_ori_n871_));
  NA3        o0843(.A(ori_ori_n871_), .B(ori_ori_n713_), .C(ori_ori_n137_), .Y(ori_ori_n872_));
  NA3        o0844(.A(ori_ori_n872_), .B(ori_ori_n193_), .C(ori_ori_n31_), .Y(ori_ori_n873_));
  NA4        o0845(.A(ori_ori_n873_), .B(ori_ori_n870_), .C(ori_ori_n635_), .D(ori_ori_n81_), .Y(ori_ori_n874_));
  NO2        o0846(.A(ori_ori_n595_), .B(ori_ori_n509_), .Y(ori_ori_n875_));
  NA2        o0847(.A(ori_ori_n875_), .B(ori_ori_n193_), .Y(ori_ori_n876_));
  NOi21      o0848(.An(f), .B(d), .Y(ori_ori_n877_));
  NA2        o0849(.A(ori_ori_n877_), .B(m), .Y(ori_ori_n878_));
  NO2        o0850(.A(ori_ori_n878_), .B(ori_ori_n52_), .Y(ori_ori_n879_));
  NOi32      o0851(.An(g), .Bn(f), .C(d), .Y(ori_ori_n880_));
  NA4        o0852(.A(ori_ori_n880_), .B(ori_ori_n615_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n881_));
  NOi21      o0853(.An(ori_ori_n321_), .B(ori_ori_n881_), .Y(ori_ori_n882_));
  AOI210     o0854(.A0(ori_ori_n879_), .A1(ori_ori_n554_), .B0(ori_ori_n882_), .Y(ori_ori_n883_));
  NA3        o0855(.A(ori_ori_n320_), .B(ori_ori_n268_), .C(ori_ori_n120_), .Y(ori_ori_n884_));
  AN2        o0856(.A(f), .B(d), .Y(ori_ori_n885_));
  NA3        o0857(.A(ori_ori_n488_), .B(ori_ori_n885_), .C(ori_ori_n83_), .Y(ori_ori_n886_));
  NO3        o0858(.A(ori_ori_n886_), .B(ori_ori_n72_), .C(ori_ori_n219_), .Y(ori_ori_n887_));
  NA2        o0859(.A(ori_ori_n884_), .B(ori_ori_n887_), .Y(ori_ori_n888_));
  NAi41      o0860(.An(ori_ori_n502_), .B(ori_ori_n888_), .C(ori_ori_n883_), .D(ori_ori_n876_), .Y(ori_ori_n889_));
  NO4        o0861(.A(ori_ori_n633_), .B(ori_ori_n133_), .C(ori_ori_n339_), .D(ori_ori_n155_), .Y(ori_ori_n890_));
  NO2        o0862(.A(ori_ori_n667_), .B(ori_ori_n339_), .Y(ori_ori_n891_));
  NO2        o0863(.A(ori_ori_n890_), .B(ori_ori_n240_), .Y(ori_ori_n892_));
  NA2        o0864(.A(ori_ori_n613_), .B(ori_ori_n83_), .Y(ori_ori_n893_));
  NO2        o0865(.A(ori_ori_n868_), .B(ori_ori_n893_), .Y(ori_ori_n894_));
  NA3        o0866(.A(ori_ori_n163_), .B(ori_ori_n109_), .C(ori_ori_n108_), .Y(ori_ori_n895_));
  OAI220     o0867(.A0(ori_ori_n886_), .A1(ori_ori_n444_), .B0(ori_ori_n351_), .B1(ori_ori_n895_), .Y(ori_ori_n896_));
  NOi41      o0868(.An(ori_ori_n229_), .B(ori_ori_n896_), .C(ori_ori_n894_), .D(ori_ori_n315_), .Y(ori_ori_n897_));
  NA2        o0869(.A(c), .B(ori_ori_n117_), .Y(ori_ori_n898_));
  NO2        o0870(.A(ori_ori_n898_), .B(ori_ori_n422_), .Y(ori_ori_n899_));
  NA3        o0871(.A(ori_ori_n899_), .B(ori_ori_n521_), .C(f), .Y(ori_ori_n900_));
  OR2        o0872(.A(ori_ori_n674_), .B(ori_ori_n550_), .Y(ori_ori_n901_));
  INV        o0873(.A(ori_ori_n901_), .Y(ori_ori_n902_));
  NA2        o0874(.A(ori_ori_n824_), .B(ori_ori_n112_), .Y(ori_ori_n903_));
  NA2        o0875(.A(ori_ori_n903_), .B(ori_ori_n902_), .Y(ori_ori_n904_));
  NA4        o0876(.A(ori_ori_n904_), .B(ori_ori_n900_), .C(ori_ori_n897_), .D(ori_ori_n892_), .Y(ori_ori_n905_));
  NO4        o0877(.A(ori_ori_n905_), .B(ori_ori_n889_), .C(ori_ori_n874_), .D(ori_ori_n861_), .Y(ori_ori_n906_));
  NA2        o0878(.A(ori_ori_n113_), .B(j), .Y(ori_ori_n907_));
  NO2        o0879(.A(ori_ori_n137_), .B(ori_ori_n133_), .Y(ori_ori_n908_));
  NO2        o0880(.A(ori_ori_n236_), .B(ori_ori_n230_), .Y(ori_ori_n909_));
  AOI220     o0881(.A0(ori_ori_n909_), .A1(ori_ori_n233_), .B0(ori_ori_n313_), .B1(ori_ori_n908_), .Y(ori_ori_n910_));
  NO2        o0882(.A(ori_ori_n444_), .B(ori_ori_n845_), .Y(ori_ori_n911_));
  NA2        o0883(.A(ori_ori_n911_), .B(ori_ori_n571_), .Y(ori_ori_n912_));
  NA2        o0884(.A(ori_ori_n912_), .B(ori_ori_n910_), .Y(ori_ori_n913_));
  NA2        o0885(.A(e), .B(d), .Y(ori_ori_n914_));
  OAI220     o0886(.A0(ori_ori_n914_), .A1(c), .B0(ori_ori_n334_), .B1(d), .Y(ori_ori_n915_));
  NA3        o0887(.A(ori_ori_n915_), .B(ori_ori_n465_), .C(ori_ori_n519_), .Y(ori_ori_n916_));
  AOI210     o0888(.A0(ori_ori_n526_), .A1(ori_ori_n184_), .B0(ori_ori_n236_), .Y(ori_ori_n917_));
  AOI210     o0889(.A0(ori_ori_n634_), .A1(ori_ori_n359_), .B0(ori_ori_n917_), .Y(ori_ori_n918_));
  INV        o0890(.A(ori_ori_n168_), .Y(ori_ori_n919_));
  NA2        o0891(.A(ori_ori_n887_), .B(ori_ori_n919_), .Y(ori_ori_n920_));
  NA3        o0892(.A(ori_ori_n171_), .B(ori_ori_n84_), .C(ori_ori_n34_), .Y(ori_ori_n921_));
  NA4        o0893(.A(ori_ori_n921_), .B(ori_ori_n920_), .C(ori_ori_n918_), .D(ori_ori_n916_), .Y(ori_ori_n922_));
  NO2        o0894(.A(ori_ori_n922_), .B(ori_ori_n913_), .Y(ori_ori_n923_));
  OR2        o0895(.A(ori_ori_n715_), .B(ori_ori_n222_), .Y(ori_ori_n924_));
  OAI220     o0896(.A0(ori_ori_n633_), .A1(ori_ori_n61_), .B0(ori_ori_n308_), .B1(j), .Y(ori_ori_n925_));
  AOI220     o0897(.A0(ori_ori_n925_), .A1(ori_ori_n891_), .B0(ori_ori_n625_), .B1(ori_ori_n632_), .Y(ori_ori_n926_));
  OAI210     o0898(.A0(ori_ori_n851_), .A1(ori_ori_n174_), .B0(ori_ori_n926_), .Y(ori_ori_n927_));
  OAI210     o0899(.A0(ori_ori_n846_), .A1(ori_ori_n919_), .B0(ori_ori_n880_), .Y(ori_ori_n928_));
  NO2        o0900(.A(ori_ori_n928_), .B(ori_ori_n616_), .Y(ori_ori_n929_));
  AOI210     o0901(.A0(ori_ori_n119_), .A1(ori_ori_n118_), .B0(ori_ori_n267_), .Y(ori_ori_n930_));
  NO2        o0902(.A(ori_ori_n930_), .B(ori_ori_n881_), .Y(ori_ori_n931_));
  AO210      o0903(.A0(ori_ori_n867_), .A1(ori_ori_n856_), .B0(ori_ori_n931_), .Y(ori_ori_n932_));
  NOi31      o0904(.An(ori_ori_n554_), .B(ori_ori_n878_), .C(ori_ori_n300_), .Y(ori_ori_n933_));
  NO4        o0905(.A(ori_ori_n933_), .B(ori_ori_n932_), .C(ori_ori_n929_), .D(ori_ori_n927_), .Y(ori_ori_n934_));
  AO220      o0906(.A0(ori_ori_n465_), .A1(ori_ori_n761_), .B0(ori_ori_n179_), .B1(f), .Y(ori_ori_n935_));
  OAI210     o0907(.A0(ori_ori_n935_), .A1(ori_ori_n468_), .B0(ori_ori_n915_), .Y(ori_ori_n936_));
  NA2        o0908(.A(ori_ori_n860_), .B(ori_ori_n719_), .Y(ori_ori_n937_));
  AN4        o0909(.A(ori_ori_n937_), .B(ori_ori_n936_), .C(ori_ori_n934_), .D(ori_ori_n924_), .Y(ori_ori_n938_));
  NA4        o0910(.A(ori_ori_n938_), .B(ori_ori_n923_), .C(ori_ori_n906_), .D(ori_ori_n853_), .Y(ori12));
  NO2        o0911(.A(ori_ori_n463_), .B(c), .Y(ori_ori_n940_));
  NO4        o0912(.A(ori_ori_n452_), .B(ori_ori_n259_), .C(ori_ori_n592_), .D(ori_ori_n219_), .Y(ori_ori_n941_));
  NA2        o0913(.A(ori_ori_n941_), .B(ori_ori_n940_), .Y(ori_ori_n942_));
  NO2        o0914(.A(ori_ori_n463_), .B(ori_ori_n117_), .Y(ori_ori_n943_));
  NO2        o0915(.A(ori_ori_n863_), .B(ori_ori_n366_), .Y(ori_ori_n944_));
  NO2        o0916(.A(ori_ori_n674_), .B(ori_ori_n393_), .Y(ori_ori_n945_));
  AOI220     o0917(.A0(ori_ori_n945_), .A1(ori_ori_n552_), .B0(ori_ori_n944_), .B1(ori_ori_n943_), .Y(ori_ori_n946_));
  NA2        o0918(.A(ori_ori_n946_), .B(ori_ori_n942_), .Y(ori_ori_n947_));
  AOI210     o0919(.A0(ori_ori_n239_), .A1(ori_ori_n350_), .B0(ori_ori_n205_), .Y(ori_ori_n948_));
  OR2        o0920(.A(ori_ori_n948_), .B(ori_ori_n941_), .Y(ori_ori_n949_));
  AOI210     o0921(.A0(ori_ori_n347_), .A1(ori_ori_n405_), .B0(ori_ori_n219_), .Y(ori_ori_n950_));
  OAI210     o0922(.A0(ori_ori_n950_), .A1(ori_ori_n949_), .B0(ori_ori_n417_), .Y(ori_ori_n951_));
  NO2        o0923(.A(ori_ori_n653_), .B(ori_ori_n270_), .Y(ori_ori_n952_));
  NO2        o0924(.A(ori_ori_n599_), .B(ori_ori_n855_), .Y(ori_ori_n953_));
  AOI220     o0925(.A0(ori_ori_n953_), .A1(ori_ori_n574_), .B0(ori_ori_n835_), .B1(ori_ori_n952_), .Y(ori_ori_n954_));
  NO2        o0926(.A(ori_ori_n154_), .B(ori_ori_n243_), .Y(ori_ori_n955_));
  NA3        o0927(.A(ori_ori_n955_), .B(ori_ori_n246_), .C(i), .Y(ori_ori_n956_));
  NA3        o0928(.A(ori_ori_n956_), .B(ori_ori_n954_), .C(ori_ori_n951_), .Y(ori_ori_n957_));
  OR2        o0929(.A(ori_ori_n335_), .B(ori_ori_n943_), .Y(ori_ori_n958_));
  NA2        o0930(.A(ori_ori_n958_), .B(ori_ori_n367_), .Y(ori_ori_n959_));
  NO3        o0931(.A(ori_ori_n133_), .B(ori_ori_n155_), .C(ori_ori_n219_), .Y(ori_ori_n960_));
  NA2        o0932(.A(ori_ori_n960_), .B(ori_ori_n541_), .Y(ori_ori_n961_));
  NA4        o0933(.A(ori_ori_n453_), .B(ori_ori_n450_), .C(ori_ori_n185_), .D(g), .Y(ori_ori_n962_));
  NA3        o0934(.A(ori_ori_n962_), .B(ori_ori_n961_), .C(ori_ori_n959_), .Y(ori_ori_n963_));
  NO3        o0935(.A(ori_ori_n679_), .B(ori_ori_n91_), .C(ori_ori_n45_), .Y(ori_ori_n964_));
  NO4        o0936(.A(ori_ori_n964_), .B(ori_ori_n963_), .C(ori_ori_n957_), .D(ori_ori_n947_), .Y(ori_ori_n965_));
  NA2        o0937(.A(ori_ori_n564_), .B(ori_ori_n147_), .Y(ori_ori_n966_));
  NOi21      o0938(.An(ori_ori_n34_), .B(ori_ori_n667_), .Y(ori_ori_n967_));
  NA2        o0939(.A(ori_ori_n967_), .B(ori_ori_n966_), .Y(ori_ori_n968_));
  OAI210     o0940(.A0(ori_ori_n257_), .A1(ori_ori_n45_), .B0(ori_ori_n968_), .Y(ori_ori_n969_));
  INV        o0941(.A(ori_ori_n331_), .Y(ori_ori_n970_));
  NO2        o0942(.A(ori_ori_n49_), .B(ori_ori_n45_), .Y(ori_ori_n971_));
  NO2        o0943(.A(ori_ori_n516_), .B(ori_ori_n308_), .Y(ori_ori_n972_));
  INV        o0944(.A(ori_ori_n972_), .Y(ori_ori_n973_));
  NO2        o0945(.A(ori_ori_n973_), .B(ori_ori_n147_), .Y(ori_ori_n974_));
  NA2        o0946(.A(ori_ori_n644_), .B(ori_ori_n376_), .Y(ori_ori_n975_));
  INV        o0947(.A(ori_ori_n380_), .Y(ori_ori_n976_));
  NO4        o0948(.A(ori_ori_n976_), .B(ori_ori_n974_), .C(ori_ori_n970_), .D(ori_ori_n969_), .Y(ori_ori_n977_));
  NA2        o0949(.A(ori_ori_n359_), .B(g), .Y(ori_ori_n978_));
  NA2        o0950(.A(ori_ori_n166_), .B(i), .Y(ori_ori_n979_));
  NA2        o0951(.A(ori_ori_n46_), .B(i), .Y(ori_ori_n980_));
  OAI220     o0952(.A0(ori_ori_n980_), .A1(ori_ori_n204_), .B0(ori_ori_n979_), .B1(ori_ori_n91_), .Y(ori_ori_n981_));
  AOI210     o0953(.A0(ori_ori_n433_), .A1(ori_ori_n37_), .B0(ori_ori_n981_), .Y(ori_ori_n982_));
  NO2        o0954(.A(ori_ori_n147_), .B(ori_ori_n83_), .Y(ori_ori_n983_));
  OR2        o0955(.A(ori_ori_n983_), .B(ori_ori_n563_), .Y(ori_ori_n984_));
  NA2        o0956(.A(ori_ori_n564_), .B(ori_ori_n397_), .Y(ori_ori_n985_));
  AOI210     o0957(.A0(ori_ori_n985_), .A1(n), .B0(ori_ori_n984_), .Y(ori_ori_n986_));
  OAI220     o0958(.A0(ori_ori_n986_), .A1(ori_ori_n978_), .B0(ori_ori_n982_), .B1(ori_ori_n344_), .Y(ori_ori_n987_));
  NO2        o0959(.A(ori_ori_n674_), .B(ori_ori_n509_), .Y(ori_ori_n988_));
  NA3        o0960(.A(ori_ori_n355_), .B(ori_ori_n639_), .C(i), .Y(ori_ori_n989_));
  OAI210     o0961(.A0(ori_ori_n451_), .A1(ori_ori_n320_), .B0(ori_ori_n989_), .Y(ori_ori_n990_));
  OAI220     o0962(.A0(ori_ori_n990_), .A1(ori_ori_n988_), .B0(ori_ori_n693_), .B1(ori_ori_n773_), .Y(ori_ori_n991_));
  NA2        o0963(.A(ori_ori_n619_), .B(ori_ori_n114_), .Y(ori_ori_n992_));
  OR3        o0964(.A(ori_ori_n320_), .B(ori_ori_n449_), .C(f), .Y(ori_ori_n993_));
  NA3        o0965(.A(ori_ori_n639_), .B(ori_ori_n79_), .C(i), .Y(ori_ori_n994_));
  OA220      o0966(.A0(ori_ori_n994_), .A1(ori_ori_n992_), .B0(ori_ori_n993_), .B1(ori_ori_n598_), .Y(ori_ori_n995_));
  NA3        o0967(.A(ori_ori_n336_), .B(ori_ori_n119_), .C(g), .Y(ori_ori_n996_));
  AOI210     o0968(.A0(ori_ori_n690_), .A1(ori_ori_n996_), .B0(m), .Y(ori_ori_n997_));
  OAI210     o0969(.A0(ori_ori_n997_), .A1(ori_ori_n944_), .B0(ori_ori_n335_), .Y(ori_ori_n998_));
  NA2        o0970(.A(ori_ori_n708_), .B(ori_ori_n893_), .Y(ori_ori_n999_));
  INV        o0971(.A(ori_ori_n857_), .Y(ori_ori_n1000_));
  NA2        o0972(.A(ori_ori_n994_), .B(ori_ori_n993_), .Y(ori_ori_n1001_));
  AOI220     o0973(.A0(ori_ori_n1001_), .A1(ori_ori_n265_), .B0(ori_ori_n1000_), .B1(ori_ori_n999_), .Y(ori_ori_n1002_));
  NA4        o0974(.A(ori_ori_n1002_), .B(ori_ori_n998_), .C(ori_ori_n995_), .D(ori_ori_n991_), .Y(ori_ori_n1003_));
  NO2        o0975(.A(ori_ori_n393_), .B(ori_ori_n90_), .Y(ori_ori_n1004_));
  OAI210     o0976(.A0(ori_ori_n1004_), .A1(ori_ori_n952_), .B0(ori_ori_n244_), .Y(ori_ori_n1005_));
  NA2        o0977(.A(ori_ori_n678_), .B(ori_ori_n87_), .Y(ori_ori_n1006_));
  NO2        o0978(.A(ori_ori_n471_), .B(ori_ori_n219_), .Y(ori_ori_n1007_));
  AOI220     o0979(.A0(ori_ori_n1007_), .A1(ori_ori_n398_), .B0(ori_ori_n958_), .B1(ori_ori_n223_), .Y(ori_ori_n1008_));
  AOI220     o0980(.A0(ori_ori_n945_), .A1(ori_ori_n955_), .B0(ori_ori_n597_), .B1(ori_ori_n89_), .Y(ori_ori_n1009_));
  NA4        o0981(.A(ori_ori_n1009_), .B(ori_ori_n1008_), .C(ori_ori_n1006_), .D(ori_ori_n1005_), .Y(ori_ori_n1010_));
  OAI210     o0982(.A0(ori_ori_n1000_), .A1(ori_ori_n953_), .B0(ori_ori_n552_), .Y(ori_ori_n1011_));
  AOI210     o0983(.A0(ori_ori_n434_), .A1(ori_ori_n426_), .B0(ori_ori_n837_), .Y(ori_ori_n1012_));
  OAI210     o0984(.A0(ori_ori_n383_), .A1(ori_ori_n382_), .B0(ori_ori_n110_), .Y(ori_ori_n1013_));
  AOI210     o0985(.A0(ori_ori_n1013_), .A1(ori_ori_n545_), .B0(ori_ori_n1012_), .Y(ori_ori_n1014_));
  NA2        o0986(.A(ori_ori_n997_), .B(ori_ori_n943_), .Y(ori_ori_n1015_));
  NO3        o0987(.A(ori_ori_n907_), .B(ori_ori_n49_), .C(ori_ori_n45_), .Y(ori_ori_n1016_));
  AOI220     o0988(.A0(ori_ori_n1016_), .A1(ori_ori_n637_), .B0(ori_ori_n658_), .B1(ori_ori_n541_), .Y(ori_ori_n1017_));
  NA4        o0989(.A(ori_ori_n1017_), .B(ori_ori_n1015_), .C(ori_ori_n1014_), .D(ori_ori_n1011_), .Y(ori_ori_n1018_));
  NO4        o0990(.A(ori_ori_n1018_), .B(ori_ori_n1010_), .C(ori_ori_n1003_), .D(ori_ori_n987_), .Y(ori_ori_n1019_));
  NAi31      o0991(.An(ori_ori_n143_), .B(ori_ori_n435_), .C(n), .Y(ori_ori_n1020_));
  NO3        o0992(.A(ori_ori_n126_), .B(ori_ori_n353_), .C(ori_ori_n864_), .Y(ori_ori_n1021_));
  NO2        o0993(.A(ori_ori_n1021_), .B(ori_ori_n1020_), .Y(ori_ori_n1022_));
  NO3        o0994(.A(ori_ori_n280_), .B(ori_ori_n143_), .C(ori_ori_n422_), .Y(ori_ori_n1023_));
  AOI210     o0995(.A0(ori_ori_n1023_), .A1(ori_ori_n510_), .B0(ori_ori_n1022_), .Y(ori_ori_n1024_));
  NA2        o0996(.A(ori_ori_n503_), .B(i), .Y(ori_ori_n1025_));
  NA2        o0997(.A(ori_ori_n1025_), .B(ori_ori_n1024_), .Y(ori_ori_n1026_));
  NA2        o0998(.A(ori_ori_n236_), .B(ori_ori_n175_), .Y(ori_ori_n1027_));
  NO3        o0999(.A(ori_ori_n317_), .B(ori_ori_n453_), .C(ori_ori_n179_), .Y(ori_ori_n1028_));
  NOi31      o1000(.An(ori_ori_n1027_), .B(ori_ori_n1028_), .C(ori_ori_n219_), .Y(ori_ori_n1029_));
  NAi21      o1001(.An(ori_ori_n564_), .B(ori_ori_n1007_), .Y(ori_ori_n1030_));
  NA2        o1002(.A(ori_ori_n494_), .B(g), .Y(ori_ori_n1031_));
  NA2        o1003(.A(ori_ori_n1031_), .B(ori_ori_n1030_), .Y(ori_ori_n1032_));
  OAI220     o1004(.A0(ori_ori_n1020_), .A1(ori_ori_n239_), .B0(ori_ori_n989_), .B1(ori_ori_n614_), .Y(ori_ori_n1033_));
  NO2        o1005(.A(ori_ori_n675_), .B(ori_ori_n393_), .Y(ori_ori_n1034_));
  NA2        o1006(.A(ori_ori_n948_), .B(ori_ori_n940_), .Y(ori_ori_n1035_));
  NO3        o1007(.A(ori_ori_n553_), .B(ori_ori_n152_), .C(ori_ori_n218_), .Y(ori_ori_n1036_));
  OAI210     o1008(.A0(ori_ori_n1036_), .A1(ori_ori_n535_), .B0(ori_ori_n394_), .Y(ori_ori_n1037_));
  OAI220     o1009(.A0(ori_ori_n945_), .A1(ori_ori_n953_), .B0(ori_ori_n554_), .B1(ori_ori_n443_), .Y(ori_ori_n1038_));
  NA4        o1010(.A(ori_ori_n1038_), .B(ori_ori_n1037_), .C(ori_ori_n1035_), .D(ori_ori_n631_), .Y(ori_ori_n1039_));
  OAI210     o1011(.A0(ori_ori_n948_), .A1(ori_ori_n941_), .B0(ori_ori_n1027_), .Y(ori_ori_n1040_));
  NA3        o1012(.A(ori_ori_n985_), .B(ori_ori_n499_), .C(ori_ori_n46_), .Y(ori_ori_n1041_));
  AOI210     o1013(.A0(ori_ori_n396_), .A1(ori_ori_n394_), .B0(ori_ori_n343_), .Y(ori_ori_n1042_));
  NA4        o1014(.A(ori_ori_n1042_), .B(ori_ori_n1041_), .C(ori_ori_n1040_), .D(ori_ori_n281_), .Y(ori_ori_n1043_));
  OR4        o1015(.A(ori_ori_n1043_), .B(ori_ori_n1039_), .C(ori_ori_n1034_), .D(ori_ori_n1033_), .Y(ori_ori_n1044_));
  NO4        o1016(.A(ori_ori_n1044_), .B(ori_ori_n1032_), .C(ori_ori_n1029_), .D(ori_ori_n1026_), .Y(ori_ori_n1045_));
  NA4        o1017(.A(ori_ori_n1045_), .B(ori_ori_n1019_), .C(ori_ori_n977_), .D(ori_ori_n965_), .Y(ori13));
  AN2        o1018(.A(c), .B(b), .Y(ori_ori_n1047_));
  NAi32      o1019(.An(d), .Bn(c), .C(e), .Y(ori_ori_n1048_));
  AN2        o1020(.A(d), .B(c), .Y(ori_ori_n1049_));
  NA2        o1021(.A(ori_ori_n1049_), .B(ori_ori_n117_), .Y(ori_ori_n1050_));
  NO3        o1022(.A(m), .B(i), .C(h), .Y(ori_ori_n1051_));
  NA3        o1023(.A(k), .B(j), .C(i), .Y(ori_ori_n1052_));
  NO3        o1024(.A(ori_ori_n1052_), .B(ori_ori_n316_), .C(ori_ori_n90_), .Y(ori_ori_n1053_));
  NOi31      o1025(.An(e), .B(d), .C(c), .Y(ori_ori_n1054_));
  NA2        o1026(.A(ori_ori_n1053_), .B(ori_ori_n1054_), .Y(ori_ori_n1055_));
  AN3        o1027(.A(g), .B(f), .C(c), .Y(ori_ori_n1056_));
  NA3        o1028(.A(l), .B(k), .C(j), .Y(ori_ori_n1057_));
  NA2        o1029(.A(i), .B(h), .Y(ori_ori_n1058_));
  NO3        o1030(.A(ori_ori_n1058_), .B(ori_ori_n1057_), .C(ori_ori_n133_), .Y(ori_ori_n1059_));
  NO3        o1031(.A(ori_ori_n144_), .B(ori_ori_n290_), .C(ori_ori_n219_), .Y(ori_ori_n1060_));
  NA3        o1032(.A(c), .B(b), .C(a), .Y(ori_ori_n1061_));
  INV        o1033(.A(ori_ori_n1055_), .Y(ori03));
  NA4        o1034(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(g), .D(ori_ori_n218_), .Y(ori_ori_n1063_));
  NA4        o1035(.A(ori_ori_n584_), .B(m), .C(ori_ori_n113_), .D(ori_ori_n218_), .Y(ori_ori_n1064_));
  NA3        o1036(.A(ori_ori_n1064_), .B(ori_ori_n384_), .C(ori_ori_n1063_), .Y(ori_ori_n1065_));
  NO2        o1037(.A(ori_ori_n1065_), .B(ori_ori_n1013_), .Y(ori_ori_n1066_));
  NOi41      o1038(.An(ori_ori_n822_), .B(ori_ori_n869_), .C(ori_ori_n858_), .D(ori_ori_n733_), .Y(ori_ori_n1067_));
  OAI220     o1039(.A0(ori_ori_n1067_), .A1(ori_ori_n708_), .B0(ori_ori_n1066_), .B1(ori_ori_n596_), .Y(ori_ori_n1068_));
  NOi31      o1040(.An(i), .B(k), .C(j), .Y(ori_ori_n1069_));
  NA4        o1041(.A(ori_ori_n1069_), .B(ori_ori_n1054_), .C(ori_ori_n355_), .D(ori_ori_n346_), .Y(ori_ori_n1070_));
  OAI210     o1042(.A0(ori_ori_n837_), .A1(ori_ori_n436_), .B0(ori_ori_n1070_), .Y(ori_ori_n1071_));
  NOi31      o1043(.An(m), .B(n), .C(f), .Y(ori_ori_n1072_));
  NA2        o1044(.A(ori_ori_n1072_), .B(ori_ori_n51_), .Y(ori_ori_n1073_));
  AN2        o1045(.A(e), .B(c), .Y(ori_ori_n1074_));
  NA2        o1046(.A(ori_ori_n1074_), .B(a), .Y(ori_ori_n1075_));
  OAI220     o1047(.A0(ori_ori_n1075_), .A1(ori_ori_n1073_), .B0(ori_ori_n901_), .B1(ori_ori_n442_), .Y(ori_ori_n1076_));
  NA2        o1048(.A(ori_ori_n519_), .B(l), .Y(ori_ori_n1077_));
  NO3        o1049(.A(ori_ori_n1076_), .B(ori_ori_n1071_), .C(ori_ori_n1012_), .Y(ori_ori_n1078_));
  NO2        o1050(.A(ori_ori_n290_), .B(a), .Y(ori_ori_n1079_));
  NO2        o1051(.A(ori_ori_n86_), .B(g), .Y(ori_ori_n1080_));
  INV        o1052(.A(ori_ori_n1078_), .Y(ori_ori_n1081_));
  NO4        o1053(.A(ori_ori_n1081_), .B(ori_ori_n1068_), .C(ori_ori_n839_), .D(ori_ori_n573_), .Y(ori_ori_n1082_));
  NA2        o1054(.A(c), .B(b), .Y(ori_ori_n1083_));
  NO2        o1055(.A(ori_ori_n718_), .B(ori_ori_n1083_), .Y(ori_ori_n1084_));
  OAI210     o1056(.A0(ori_ori_n878_), .A1(ori_ori_n849_), .B0(ori_ori_n429_), .Y(ori_ori_n1085_));
  OAI210     o1057(.A0(ori_ori_n1085_), .A1(ori_ori_n879_), .B0(ori_ori_n1084_), .Y(ori_ori_n1086_));
  NAi21      o1058(.An(ori_ori_n437_), .B(ori_ori_n1084_), .Y(ori_ori_n1087_));
  OAI210     o1059(.A0(ori_ori_n558_), .A1(ori_ori_n39_), .B0(ori_ori_n1079_), .Y(ori_ori_n1088_));
  NA2        o1060(.A(ori_ori_n1088_), .B(ori_ori_n1087_), .Y(ori_ori_n1089_));
  NA2        o1061(.A(ori_ori_n268_), .B(ori_ori_n120_), .Y(ori_ori_n1090_));
  OAI210     o1062(.A0(ori_ori_n1090_), .A1(ori_ori_n294_), .B0(g), .Y(ori_ori_n1091_));
  NAi21      o1063(.An(f), .B(d), .Y(ori_ori_n1092_));
  NO2        o1064(.A(ori_ori_n1092_), .B(ori_ori_n1061_), .Y(ori_ori_n1093_));
  INV        o1065(.A(ori_ori_n1093_), .Y(ori_ori_n1094_));
  AOI210     o1066(.A0(ori_ori_n1091_), .A1(ori_ori_n300_), .B0(ori_ori_n1094_), .Y(ori_ori_n1095_));
  AOI210     o1067(.A0(ori_ori_n1095_), .A1(ori_ori_n114_), .B0(ori_ori_n1089_), .Y(ori_ori_n1096_));
  NA2        o1068(.A(ori_ori_n482_), .B(ori_ori_n481_), .Y(ori_ori_n1097_));
  NO2        o1069(.A(ori_ori_n186_), .B(ori_ori_n243_), .Y(ori_ori_n1098_));
  NA2        o1070(.A(ori_ori_n1098_), .B(m), .Y(ori_ori_n1099_));
  NA3        o1071(.A(ori_ori_n930_), .B(ori_ori_n1077_), .C(ori_ori_n168_), .Y(ori_ori_n1100_));
  OAI210     o1072(.A0(ori_ori_n1100_), .A1(ori_ori_n321_), .B0(ori_ori_n483_), .Y(ori_ori_n1101_));
  AOI210     o1073(.A0(ori_ori_n1101_), .A1(ori_ori_n1097_), .B0(ori_ori_n1099_), .Y(ori_ori_n1102_));
  NA2        o1074(.A(ori_ori_n571_), .B(ori_ori_n424_), .Y(ori_ori_n1103_));
  NA2        o1075(.A(ori_ori_n162_), .B(ori_ori_n33_), .Y(ori_ori_n1104_));
  AOI210     o1076(.A0(ori_ori_n975_), .A1(ori_ori_n1104_), .B0(ori_ori_n219_), .Y(ori_ori_n1105_));
  OAI210     o1077(.A0(ori_ori_n1105_), .A1(ori_ori_n456_), .B0(ori_ori_n1093_), .Y(ori_ori_n1106_));
  NO2        o1078(.A(ori_ori_n387_), .B(ori_ori_n386_), .Y(ori_ori_n1107_));
  NA2        o1079(.A(ori_ori_n1098_), .B(ori_ori_n445_), .Y(ori_ori_n1108_));
  NAi41      o1080(.An(ori_ori_n1107_), .B(ori_ori_n1108_), .C(ori_ori_n1106_), .D(ori_ori_n1103_), .Y(ori_ori_n1109_));
  NO2        o1081(.A(ori_ori_n1109_), .B(ori_ori_n1102_), .Y(ori_ori_n1110_));
  NA4        o1082(.A(ori_ori_n1110_), .B(ori_ori_n1096_), .C(ori_ori_n1086_), .D(ori_ori_n1082_), .Y(ori00));
  AOI210     o1083(.A0(ori_ori_n911_), .A1(ori_ori_n955_), .B0(ori_ori_n1071_), .Y(ori_ori_n1112_));
  INV        o1084(.A(ori_ori_n730_), .Y(ori_ori_n1113_));
  NA3        o1085(.A(ori_ori_n1113_), .B(ori_ori_n1112_), .C(ori_ori_n1014_), .Y(ori_ori_n1114_));
  NA2        o1086(.A(ori_ori_n521_), .B(f), .Y(ori_ori_n1115_));
  OAI210     o1087(.A0(ori_ori_n1021_), .A1(ori_ori_n40_), .B0(ori_ori_n660_), .Y(ori_ori_n1116_));
  NA3        o1088(.A(ori_ori_n1116_), .B(ori_ori_n264_), .C(n), .Y(ori_ori_n1117_));
  AOI210     o1089(.A0(ori_ori_n1117_), .A1(ori_ori_n1115_), .B0(ori_ori_n1050_), .Y(ori_ori_n1118_));
  NO2        o1090(.A(ori_ori_n1118_), .B(ori_ori_n1114_), .Y(ori_ori_n1119_));
  NA3        o1091(.A(ori_ori_n171_), .B(ori_ori_n46_), .C(ori_ori_n45_), .Y(ori_ori_n1120_));
  NA3        o1092(.A(d), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n1121_));
  NO2        o1093(.A(ori_ori_n1121_), .B(ori_ori_n1120_), .Y(ori_ori_n1122_));
  INV        o1094(.A(ori_ori_n586_), .Y(ori_ori_n1123_));
  NO4        o1095(.A(ori_ori_n1123_), .B(ori_ori_n1122_), .C(ori_ori_n1107_), .D(ori_ori_n933_), .Y(ori_ori_n1124_));
  NO4        o1096(.A(ori_ori_n500_), .B(ori_ori_n369_), .C(ori_ori_n1083_), .D(ori_ori_n59_), .Y(ori_ori_n1125_));
  NA3        o1097(.A(ori_ori_n399_), .B(ori_ori_n226_), .C(g), .Y(ori_ori_n1126_));
  OA220      o1098(.A0(ori_ori_n1126_), .A1(ori_ori_n1121_), .B0(ori_ori_n400_), .B1(ori_ori_n136_), .Y(ori_ori_n1127_));
  NO2        o1099(.A(h), .B(g), .Y(ori_ori_n1128_));
  NA4        o1100(.A(ori_ori_n510_), .B(ori_ori_n479_), .C(ori_ori_n1128_), .D(ori_ori_n1047_), .Y(ori_ori_n1129_));
  NA2        o1101(.A(ori_ori_n960_), .B(ori_ori_n585_), .Y(ori_ori_n1130_));
  AOI220     o1102(.A0(ori_ori_n328_), .A1(ori_ori_n253_), .B0(ori_ori_n181_), .B1(ori_ori_n151_), .Y(ori_ori_n1131_));
  NA4        o1103(.A(ori_ori_n1131_), .B(ori_ori_n1130_), .C(ori_ori_n1129_), .D(ori_ori_n1127_), .Y(ori_ori_n1132_));
  NO3        o1104(.A(ori_ori_n1132_), .B(ori_ori_n1125_), .C(ori_ori_n274_), .Y(ori_ori_n1133_));
  INV        o1105(.A(ori_ori_n333_), .Y(ori_ori_n1134_));
  AOI210     o1106(.A0(ori_ori_n253_), .A1(ori_ori_n359_), .B0(ori_ori_n588_), .Y(ori_ori_n1135_));
  NA3        o1107(.A(ori_ori_n1135_), .B(ori_ori_n1134_), .C(ori_ori_n157_), .Y(ori_ori_n1136_));
  NO2        o1108(.A(ori_ori_n245_), .B(ori_ori_n185_), .Y(ori_ori_n1137_));
  NA2        o1109(.A(ori_ori_n1137_), .B(ori_ori_n443_), .Y(ori_ori_n1138_));
  NAi31      o1110(.An(ori_ori_n189_), .B(ori_ori_n875_), .C(ori_ori_n479_), .Y(ori_ori_n1139_));
  NA2        o1111(.A(ori_ori_n1139_), .B(ori_ori_n1138_), .Y(ori_ori_n1140_));
  NO3        o1112(.A(ori_ori_n1140_), .B(ori_ori_n1136_), .C(ori_ori_n529_), .Y(ori_ori_n1141_));
  AN3        o1113(.A(ori_ori_n1141_), .B(ori_ori_n1133_), .C(ori_ori_n1124_), .Y(ori_ori_n1142_));
  NA2        o1114(.A(ori_ori_n545_), .B(ori_ori_n101_), .Y(ori_ori_n1143_));
  NA3        o1115(.A(ori_ori_n1072_), .B(ori_ori_n619_), .C(ori_ori_n478_), .Y(ori_ori_n1144_));
  NA4        o1116(.A(ori_ori_n1144_), .B(ori_ori_n572_), .C(ori_ori_n1143_), .D(ori_ori_n247_), .Y(ori_ori_n1145_));
  NA2        o1117(.A(ori_ori_n1065_), .B(ori_ori_n545_), .Y(ori_ori_n1146_));
  NA4        o1118(.A(ori_ori_n663_), .B(ori_ori_n210_), .C(ori_ori_n226_), .D(ori_ori_n166_), .Y(ori_ori_n1147_));
  NA3        o1119(.A(ori_ori_n1147_), .B(ori_ori_n1146_), .C(ori_ori_n304_), .Y(ori_ori_n1148_));
  OAI210     o1120(.A0(ori_ori_n477_), .A1(ori_ori_n121_), .B0(ori_ori_n881_), .Y(ori_ori_n1149_));
  AOI220     o1121(.A0(ori_ori_n1149_), .A1(ori_ori_n1100_), .B0(ori_ori_n571_), .B1(ori_ori_n424_), .Y(ori_ori_n1150_));
  NA2        o1122(.A(n), .B(e), .Y(ori_ori_n1151_));
  NO2        o1123(.A(ori_ori_n1151_), .B(ori_ori_n149_), .Y(ori_ori_n1152_));
  NA2        o1124(.A(ori_ori_n1152_), .B(ori_ori_n282_), .Y(ori_ori_n1153_));
  OAI210     o1125(.A0(ori_ori_n370_), .A1(ori_ori_n322_), .B0(ori_ori_n458_), .Y(ori_ori_n1154_));
  NA3        o1126(.A(ori_ori_n1154_), .B(ori_ori_n1153_), .C(ori_ori_n1150_), .Y(ori_ori_n1155_));
  AOI210     o1127(.A0(ori_ori_n1152_), .A1(ori_ori_n866_), .B0(ori_ori_n838_), .Y(ori_ori_n1156_));
  AOI220     o1128(.A0(ori_ori_n967_), .A1(ori_ori_n585_), .B0(ori_ori_n663_), .B1(ori_ori_n250_), .Y(ori_ori_n1157_));
  NO2        o1129(.A(ori_ori_n68_), .B(h), .Y(ori_ori_n1158_));
  NA3        o1130(.A(ori_ori_n1157_), .B(ori_ori_n1156_), .C(ori_ori_n883_), .Y(ori_ori_n1159_));
  NO4        o1131(.A(ori_ori_n1159_), .B(ori_ori_n1155_), .C(ori_ori_n1148_), .D(ori_ori_n1145_), .Y(ori_ori_n1160_));
  NA2        o1132(.A(ori_ori_n850_), .B(ori_ori_n772_), .Y(ori_ori_n1161_));
  NA4        o1133(.A(ori_ori_n1161_), .B(ori_ori_n1160_), .C(ori_ori_n1142_), .D(ori_ori_n1119_), .Y(ori01));
  AN2        o1134(.A(ori_ori_n1037_), .B(ori_ori_n1035_), .Y(ori_ori_n1163_));
  NO3        o1135(.A(ori_ori_n818_), .B(ori_ori_n491_), .C(ori_ori_n288_), .Y(ori_ori_n1164_));
  NA2        o1136(.A(ori_ori_n410_), .B(i), .Y(ori_ori_n1165_));
  NA3        o1137(.A(ori_ori_n1165_), .B(ori_ori_n1164_), .C(ori_ori_n1163_), .Y(ori_ori_n1166_));
  NA2        o1138(.A(ori_ori_n597_), .B(ori_ori_n89_), .Y(ori_ori_n1167_));
  NA2        o1139(.A(ori_ori_n564_), .B(ori_ori_n279_), .Y(ori_ori_n1168_));
  NA2        o1140(.A(ori_ori_n972_), .B(ori_ori_n1168_), .Y(ori_ori_n1169_));
  NA4        o1141(.A(ori_ori_n1169_), .B(ori_ori_n1167_), .C(ori_ori_n926_), .D(ori_ori_n345_), .Y(ori_ori_n1170_));
  NA2        o1142(.A(ori_ori_n45_), .B(f), .Y(ori_ori_n1171_));
  NA2        o1143(.A(ori_ori_n725_), .B(ori_ori_n96_), .Y(ori_ori_n1172_));
  NO2        o1144(.A(ori_ori_n1172_), .B(ori_ori_n1171_), .Y(ori_ori_n1173_));
  OAI210     o1145(.A0(ori_ori_n798_), .A1(ori_ori_n614_), .B0(ori_ori_n1147_), .Y(ori_ori_n1174_));
  AOI210     o1146(.A0(ori_ori_n1173_), .A1(ori_ori_n648_), .B0(ori_ori_n1174_), .Y(ori_ori_n1175_));
  INV        o1147(.A(ori_ori_n119_), .Y(ori_ori_n1176_));
  OR2        o1148(.A(ori_ori_n676_), .B(ori_ori_n384_), .Y(ori_ori_n1177_));
  NAi41      o1149(.An(ori_ori_n165_), .B(ori_ori_n1177_), .C(ori_ori_n1175_), .D(ori_ori_n910_), .Y(ori_ori_n1178_));
  NO2        o1150(.A(ori_ori_n692_), .B(ori_ori_n524_), .Y(ori_ori_n1179_));
  NA4        o1151(.A(ori_ori_n725_), .B(ori_ori_n96_), .C(ori_ori_n45_), .D(ori_ori_n218_), .Y(ori_ori_n1180_));
  OA220      o1152(.A0(ori_ori_n1180_), .A1(ori_ori_n685_), .B0(ori_ori_n199_), .B1(ori_ori_n197_), .Y(ori_ori_n1181_));
  NA3        o1153(.A(ori_ori_n1181_), .B(ori_ori_n1179_), .C(ori_ori_n139_), .Y(ori_ori_n1182_));
  NO4        o1154(.A(ori_ori_n1182_), .B(ori_ori_n1178_), .C(ori_ori_n1170_), .D(ori_ori_n1166_), .Y(ori_ori_n1183_));
  INV        o1155(.A(ori_ori_n1126_), .Y(ori_ori_n1184_));
  OAI210     o1156(.A0(ori_ori_n1184_), .A1(ori_ori_n310_), .B0(ori_ori_n541_), .Y(ori_ori_n1185_));
  AOI210     o1157(.A0(ori_ori_n208_), .A1(ori_ori_n88_), .B0(ori_ori_n218_), .Y(ori_ori_n1186_));
  OAI210     o1158(.A0(ori_ori_n825_), .A1(ori_ori_n443_), .B0(ori_ori_n1186_), .Y(ori_ori_n1187_));
  AN3        o1159(.A(m), .B(l), .C(k), .Y(ori_ori_n1188_));
  OAI210     o1160(.A0(ori_ori_n372_), .A1(ori_ori_n34_), .B0(ori_ori_n1188_), .Y(ori_ori_n1189_));
  NA2        o1161(.A(ori_ori_n207_), .B(ori_ori_n34_), .Y(ori_ori_n1190_));
  AO210      o1162(.A0(ori_ori_n1190_), .A1(ori_ori_n1189_), .B0(ori_ori_n344_), .Y(ori_ori_n1191_));
  NA3        o1163(.A(ori_ori_n1191_), .B(ori_ori_n1187_), .C(ori_ori_n1185_), .Y(ori_ori_n1192_));
  AOI210     o1164(.A0(ori_ori_n606_), .A1(ori_ori_n119_), .B0(ori_ori_n612_), .Y(ori_ori_n1193_));
  OAI210     o1165(.A0(ori_ori_n1176_), .A1(ori_ori_n603_), .B0(ori_ori_n1193_), .Y(ori_ori_n1194_));
  NA2        o1166(.A(ori_ori_n287_), .B(ori_ori_n199_), .Y(ori_ori_n1195_));
  NA2        o1167(.A(ori_ori_n1195_), .B(ori_ori_n681_), .Y(ori_ori_n1196_));
  NO3        o1168(.A(ori_ori_n837_), .B(ori_ori_n208_), .C(ori_ori_n422_), .Y(ori_ori_n1197_));
  INV        o1169(.A(ori_ori_n1197_), .Y(ori_ori_n1198_));
  OAI210     o1170(.A0(ori_ori_n1173_), .A1(ori_ori_n338_), .B0(ori_ori_n693_), .Y(ori_ori_n1199_));
  NA4        o1171(.A(ori_ori_n1199_), .B(ori_ori_n1198_), .C(ori_ori_n1196_), .D(ori_ori_n801_), .Y(ori_ori_n1200_));
  NO3        o1172(.A(ori_ori_n1200_), .B(ori_ori_n1194_), .C(ori_ori_n1192_), .Y(ori_ori_n1201_));
  NA3        o1173(.A(ori_ori_n615_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1202_));
  NO2        o1174(.A(ori_ori_n1202_), .B(ori_ori_n208_), .Y(ori_ori_n1203_));
  AOI210     o1175(.A0(ori_ori_n517_), .A1(ori_ori_n58_), .B0(ori_ori_n1203_), .Y(ori_ori_n1204_));
  OR3        o1176(.A(ori_ori_n1172_), .B(ori_ori_n616_), .C(ori_ori_n1171_), .Y(ori_ori_n1205_));
  NO2        o1177(.A(ori_ori_n1180_), .B(ori_ori_n992_), .Y(ori_ori_n1206_));
  NO2        o1178(.A(ori_ori_n211_), .B(ori_ori_n112_), .Y(ori_ori_n1207_));
  NO3        o1179(.A(ori_ori_n1207_), .B(ori_ori_n1206_), .C(ori_ori_n1122_), .Y(ori_ori_n1208_));
  NA4        o1180(.A(ori_ori_n1208_), .B(ori_ori_n1205_), .C(ori_ori_n1204_), .D(ori_ori_n771_), .Y(ori_ori_n1209_));
  NO2        o1181(.A(ori_ori_n979_), .B(ori_ori_n238_), .Y(ori_ori_n1210_));
  NO2        o1182(.A(ori_ori_n980_), .B(ori_ori_n566_), .Y(ori_ori_n1211_));
  OAI210     o1183(.A0(ori_ori_n1211_), .A1(ori_ori_n1210_), .B0(ori_ori_n353_), .Y(ori_ori_n1212_));
  NA2        o1184(.A(ori_ori_n580_), .B(ori_ori_n578_), .Y(ori_ori_n1213_));
  NO3        o1185(.A(ori_ori_n78_), .B(ori_ori_n308_), .C(ori_ori_n45_), .Y(ori_ori_n1214_));
  NA2        o1186(.A(ori_ori_n1214_), .B(ori_ori_n563_), .Y(ori_ori_n1215_));
  NA3        o1187(.A(ori_ori_n1215_), .B(ori_ori_n1213_), .C(ori_ori_n687_), .Y(ori_ori_n1216_));
  OR2        o1188(.A(ori_ori_n1126_), .B(ori_ori_n1121_), .Y(ori_ori_n1217_));
  NO2        o1189(.A(ori_ori_n384_), .B(ori_ori_n71_), .Y(ori_ori_n1218_));
  INV        o1190(.A(ori_ori_n1218_), .Y(ori_ori_n1219_));
  NA2        o1191(.A(ori_ori_n1214_), .B(ori_ori_n828_), .Y(ori_ori_n1220_));
  NA4        o1192(.A(ori_ori_n1220_), .B(ori_ori_n1219_), .C(ori_ori_n1217_), .D(ori_ori_n402_), .Y(ori_ori_n1221_));
  NOi41      o1193(.An(ori_ori_n1212_), .B(ori_ori_n1221_), .C(ori_ori_n1216_), .D(ori_ori_n1209_), .Y(ori_ori_n1222_));
  NO2        o1194(.A(ori_ori_n132_), .B(ori_ori_n45_), .Y(ori_ori_n1223_));
  NO2        o1195(.A(ori_ori_n45_), .B(ori_ori_n40_), .Y(ori_ori_n1224_));
  AO220      o1196(.A0(ori_ori_n1224_), .A1(ori_ori_n634_), .B0(ori_ori_n1223_), .B1(ori_ori_n723_), .Y(ori_ori_n1225_));
  NA2        o1197(.A(ori_ori_n1225_), .B(ori_ori_n353_), .Y(ori_ori_n1226_));
  INV        o1198(.A(ori_ori_n136_), .Y(ori_ori_n1227_));
  NO3        o1199(.A(ori_ori_n1058_), .B(ori_ori_n180_), .C(ori_ori_n86_), .Y(ori_ori_n1228_));
  AOI220     o1200(.A0(ori_ori_n1228_), .A1(ori_ori_n1227_), .B0(ori_ori_n1214_), .B1(ori_ori_n983_), .Y(ori_ori_n1229_));
  NA2        o1201(.A(ori_ori_n1229_), .B(ori_ori_n1226_), .Y(ori_ori_n1230_));
  NO2        o1202(.A(ori_ori_n627_), .B(ori_ori_n626_), .Y(ori_ori_n1231_));
  NO4        o1203(.A(ori_ori_n1058_), .B(ori_ori_n1231_), .C(ori_ori_n178_), .D(ori_ori_n86_), .Y(ori_ori_n1232_));
  NO3        o1204(.A(ori_ori_n1232_), .B(ori_ori_n1230_), .C(ori_ori_n652_), .Y(ori_ori_n1233_));
  NA4        o1205(.A(ori_ori_n1233_), .B(ori_ori_n1222_), .C(ori_ori_n1201_), .D(ori_ori_n1183_), .Y(ori06));
  NO2        o1206(.A(ori_ori_n423_), .B(ori_ori_n570_), .Y(ori_ori_n1235_));
  NA2        o1207(.A(ori_ori_n275_), .B(ori_ori_n1235_), .Y(ori_ori_n1236_));
  NO2        o1208(.A(ori_ori_n230_), .B(ori_ori_n103_), .Y(ori_ori_n1237_));
  OAI210     o1209(.A0(ori_ori_n1237_), .A1(ori_ori_n1228_), .B0(ori_ori_n398_), .Y(ori_ori_n1238_));
  NO3        o1210(.A(ori_ori_n610_), .B(ori_ori_n823_), .C(ori_ori_n613_), .Y(ori_ori_n1239_));
  OR2        o1211(.A(ori_ori_n1239_), .B(ori_ori_n901_), .Y(ori_ori_n1240_));
  NA4        o1212(.A(ori_ori_n1240_), .B(ori_ori_n1238_), .C(ori_ori_n1236_), .D(ori_ori_n1212_), .Y(ori_ori_n1241_));
  NO3        o1213(.A(ori_ori_n1241_), .B(ori_ori_n1216_), .C(ori_ori_n263_), .Y(ori_ori_n1242_));
  NO2        o1214(.A(ori_ori_n308_), .B(ori_ori_n45_), .Y(ori_ori_n1243_));
  AOI210     o1215(.A0(ori_ori_n1243_), .A1(ori_ori_n984_), .B0(ori_ori_n1210_), .Y(ori_ori_n1244_));
  AOI210     o1216(.A0(ori_ori_n1243_), .A1(ori_ori_n567_), .B0(ori_ori_n1225_), .Y(ori_ori_n1245_));
  AOI210     o1217(.A0(ori_ori_n1245_), .A1(ori_ori_n1244_), .B0(ori_ori_n350_), .Y(ori_ori_n1246_));
  OAI210     o1218(.A0(ori_ori_n88_), .A1(ori_ori_n40_), .B0(ori_ori_n691_), .Y(ori_ori_n1247_));
  NA2        o1219(.A(ori_ori_n1247_), .B(ori_ori_n656_), .Y(ori_ori_n1248_));
  NO2        o1220(.A(ori_ori_n526_), .B(ori_ori_n175_), .Y(ori_ori_n1249_));
  NOi21      o1221(.An(ori_ori_n138_), .B(ori_ori_n45_), .Y(ori_ori_n1250_));
  NO2        o1222(.A(ori_ori_n620_), .B(ori_ori_n1073_), .Y(ori_ori_n1251_));
  OAI210     o1223(.A0(ori_ori_n472_), .A1(ori_ori_n254_), .B0(ori_ori_n921_), .Y(ori_ori_n1252_));
  NO4        o1224(.A(ori_ori_n1252_), .B(ori_ori_n1251_), .C(ori_ori_n1250_), .D(ori_ori_n1249_), .Y(ori_ori_n1253_));
  OR2        o1225(.A(ori_ori_n611_), .B(ori_ori_n609_), .Y(ori_ori_n1254_));
  NO2        o1226(.A(ori_ori_n383_), .B(ori_ori_n137_), .Y(ori_ori_n1255_));
  AOI210     o1227(.A0(ori_ori_n1255_), .A1(ori_ori_n597_), .B0(ori_ori_n1254_), .Y(ori_ori_n1256_));
  NA3        o1228(.A(ori_ori_n1256_), .B(ori_ori_n1253_), .C(ori_ori_n1248_), .Y(ori_ori_n1257_));
  NO2        o1229(.A(ori_ori_n762_), .B(ori_ori_n382_), .Y(ori_ori_n1258_));
  NO3        o1230(.A(ori_ori_n693_), .B(ori_ori_n773_), .C(ori_ori_n648_), .Y(ori_ori_n1259_));
  NOi21      o1231(.An(ori_ori_n1258_), .B(ori_ori_n1259_), .Y(ori_ori_n1260_));
  AN2        o1232(.A(ori_ori_n967_), .B(ori_ori_n659_), .Y(ori_ori_n1261_));
  NO4        o1233(.A(ori_ori_n1261_), .B(ori_ori_n1260_), .C(ori_ori_n1257_), .D(ori_ori_n1246_), .Y(ori_ori_n1262_));
  NO2        o1234(.A(ori_ori_n817_), .B(ori_ori_n284_), .Y(ori_ori_n1263_));
  NO2        o1235(.A(ori_ori_n749_), .B(ori_ori_n47_), .Y(ori_ori_n1264_));
  AOI220     o1236(.A0(ori_ori_n375_), .A1(ori_ori_n1264_), .B0(ori_ori_n1263_), .B1(ori_ori_n275_), .Y(ori_ori_n1265_));
  NO3        o1237(.A(ori_ori_n249_), .B(ori_ori_n103_), .C(ori_ori_n290_), .Y(ori_ori_n1266_));
  OAI220     o1238(.A0(ori_ori_n715_), .A1(ori_ori_n254_), .B0(ori_ori_n523_), .B1(ori_ori_n526_), .Y(ori_ori_n1267_));
  OAI210     o1239(.A0(l), .A1(i), .B0(k), .Y(ori_ori_n1268_));
  NO3        o1240(.A(ori_ori_n1268_), .B(ori_ori_n608_), .C(j), .Y(ori_ori_n1269_));
  NOi21      o1241(.An(ori_ori_n1269_), .B(ori_ori_n685_), .Y(ori_ori_n1270_));
  NO4        o1242(.A(ori_ori_n1270_), .B(ori_ori_n1267_), .C(ori_ori_n1266_), .D(ori_ori_n1076_), .Y(ori_ori_n1271_));
  NA3        o1243(.A(ori_ori_n809_), .B(ori_ori_n808_), .C(ori_ori_n893_), .Y(ori_ori_n1272_));
  NAi31      o1244(.An(ori_ori_n762_), .B(ori_ori_n1272_), .C(ori_ori_n207_), .Y(ori_ori_n1273_));
  NA4        o1245(.A(ori_ori_n1273_), .B(ori_ori_n1271_), .C(ori_ori_n1265_), .D(ori_ori_n1157_), .Y(ori_ori_n1274_));
  OR3        o1246(.A(ori_ori_n1239_), .B(ori_ori_n798_), .C(ori_ori_n550_), .Y(ori_ori_n1275_));
  AOI210     o1247(.A0(ori_ori_n580_), .A1(ori_ori_n458_), .B0(ori_ori_n388_), .Y(ori_ori_n1276_));
  NA2        o1248(.A(ori_ori_n1269_), .B(ori_ori_n805_), .Y(ori_ori_n1277_));
  NA3        o1249(.A(ori_ori_n1277_), .B(ori_ori_n1276_), .C(ori_ori_n1275_), .Y(ori_ori_n1278_));
  AOI220     o1250(.A0(ori_ori_n1258_), .A1(ori_ori_n772_), .B0(ori_ori_n1255_), .B1(ori_ori_n244_), .Y(ori_ori_n1279_));
  AN2        o1251(.A(ori_ori_n941_), .B(ori_ori_n940_), .Y(ori_ori_n1280_));
  NO3        o1252(.A(ori_ori_n1280_), .B(ori_ori_n513_), .C(ori_ori_n494_), .Y(ori_ori_n1281_));
  NA3        o1253(.A(ori_ori_n1281_), .B(ori_ori_n1279_), .C(ori_ori_n1220_), .Y(ori_ori_n1282_));
  NAi21      o1254(.An(j), .B(i), .Y(ori_ori_n1283_));
  NO4        o1255(.A(ori_ori_n1231_), .B(ori_ori_n1283_), .C(ori_ori_n452_), .D(ori_ori_n241_), .Y(ori_ori_n1284_));
  NO4        o1256(.A(ori_ori_n1284_), .B(ori_ori_n1282_), .C(ori_ori_n1278_), .D(ori_ori_n1274_), .Y(ori_ori_n1285_));
  NA4        o1257(.A(ori_ori_n1285_), .B(ori_ori_n1262_), .C(ori_ori_n1242_), .D(ori_ori_n1233_), .Y(ori07));
  NAi32      o1258(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1287_));
  NO3        o1259(.A(ori_ori_n1287_), .B(g), .C(f), .Y(ori_ori_n1288_));
  NAi21      o1260(.An(f), .B(c), .Y(ori_ori_n1289_));
  OR2        o1261(.A(e), .B(d), .Y(ori_ori_n1290_));
  NOi31      o1262(.An(n), .B(m), .C(b), .Y(ori_ori_n1291_));
  NOi41      o1263(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1292_));
  NO2        o1264(.A(ori_ori_n1052_), .B(ori_ori_n316_), .Y(ori_ori_n1293_));
  NA2        o1265(.A(ori_ori_n551_), .B(ori_ori_n79_), .Y(ori_ori_n1294_));
  NA2        o1266(.A(ori_ori_n1158_), .B(ori_ori_n298_), .Y(ori_ori_n1295_));
  NA2        o1267(.A(ori_ori_n1295_), .B(ori_ori_n1294_), .Y(ori_ori_n1296_));
  NO2        o1268(.A(ori_ori_n1296_), .B(ori_ori_n1288_), .Y(ori_ori_n1297_));
  NO3        o1269(.A(e), .B(d), .C(c), .Y(ori_ori_n1298_));
  NO2        o1270(.A(ori_ori_n133_), .B(ori_ori_n219_), .Y(ori_ori_n1299_));
  NA2        o1271(.A(ori_ori_n1299_), .B(ori_ori_n1298_), .Y(ori_ori_n1300_));
  INV        o1272(.A(ori_ori_n1300_), .Y(ori_ori_n1301_));
  NA3        o1273(.A(ori_ori_n712_), .B(ori_ori_n700_), .C(ori_ori_n113_), .Y(ori_ori_n1302_));
  NO2        o1274(.A(ori_ori_n1302_), .B(ori_ori_n45_), .Y(ori_ori_n1303_));
  NO2        o1275(.A(l), .B(k), .Y(ori_ori_n1304_));
  NO3        o1276(.A(ori_ori_n452_), .B(d), .C(c), .Y(ori_ori_n1305_));
  NO2        o1277(.A(ori_ori_n1303_), .B(ori_ori_n1301_), .Y(ori_ori_n1306_));
  NO2        o1278(.A(g), .B(c), .Y(ori_ori_n1307_));
  NA2        o1279(.A(ori_ori_n1307_), .B(ori_ori_n144_), .Y(ori_ori_n1308_));
  INV        o1280(.A(ori_ori_n1308_), .Y(ori_ori_n1309_));
  NA2        o1281(.A(ori_ori_n1309_), .B(ori_ori_n183_), .Y(ori_ori_n1310_));
  NO2        o1282(.A(ori_ori_n463_), .B(a), .Y(ori_ori_n1311_));
  NA2        o1283(.A(ori_ori_n1311_), .B(ori_ori_n114_), .Y(ori_ori_n1312_));
  NA2        o1284(.A(ori_ori_n140_), .B(ori_ori_n226_), .Y(ori_ori_n1313_));
  NO2        o1285(.A(ori_ori_n1313_), .B(ori_ori_n1406_), .Y(ori_ori_n1314_));
  NO2        o1286(.A(ori_ori_n769_), .B(ori_ori_n191_), .Y(ori_ori_n1315_));
  NOi31      o1287(.An(m), .B(n), .C(b), .Y(ori_ori_n1316_));
  NOi31      o1288(.An(f), .B(d), .C(c), .Y(ori_ori_n1317_));
  NA2        o1289(.A(ori_ori_n1317_), .B(ori_ori_n1316_), .Y(ori_ori_n1318_));
  INV        o1290(.A(ori_ori_n1318_), .Y(ori_ori_n1319_));
  NO3        o1291(.A(ori_ori_n1319_), .B(ori_ori_n1315_), .C(ori_ori_n1314_), .Y(ori_ori_n1320_));
  NA2        o1292(.A(ori_ori_n1056_), .B(ori_ori_n479_), .Y(ori_ori_n1321_));
  NO2        o1293(.A(ori_ori_n1321_), .B(ori_ori_n452_), .Y(ori_ori_n1322_));
  NO3        o1294(.A(ori_ori_n41_), .B(i), .C(h), .Y(ori_ori_n1323_));
  NO2        o1295(.A(ori_ori_n1051_), .B(ori_ori_n1322_), .Y(ori_ori_n1324_));
  AN4        o1296(.A(ori_ori_n1324_), .B(ori_ori_n1320_), .C(ori_ori_n1312_), .D(ori_ori_n1310_), .Y(ori_ori_n1325_));
  NA2        o1297(.A(ori_ori_n1291_), .B(ori_ori_n395_), .Y(ori_ori_n1326_));
  INV        o1298(.A(ori_ori_n1326_), .Y(ori_ori_n1327_));
  NA2        o1299(.A(ori_ori_n1305_), .B(ori_ori_n220_), .Y(ori_ori_n1328_));
  INV        o1300(.A(ori_ori_n1059_), .Y(ori_ori_n1329_));
  NAi31      o1301(.An(ori_ori_n1327_), .B(ori_ori_n1329_), .C(ori_ori_n1328_), .Y(ori_ori_n1330_));
  NO4        o1302(.A(ori_ori_n133_), .B(g), .C(f), .D(e), .Y(ori_ori_n1331_));
  NA2        o1303(.A(ori_ori_n1292_), .B(ori_ori_n1304_), .Y(ori_ori_n1332_));
  INV        o1304(.A(ori_ori_n1332_), .Y(ori_ori_n1333_));
  OR3        o1305(.A(ori_ori_n550_), .B(ori_ori_n549_), .C(ori_ori_n113_), .Y(ori_ori_n1334_));
  NA2        o1306(.A(ori_ori_n1072_), .B(ori_ori_n422_), .Y(ori_ori_n1335_));
  NO2        o1307(.A(ori_ori_n1335_), .B(ori_ori_n450_), .Y(ori_ori_n1336_));
  AO210      o1308(.A0(ori_ori_n1336_), .A1(ori_ori_n117_), .B0(ori_ori_n1333_), .Y(ori_ori_n1337_));
  NO2        o1309(.A(ori_ori_n1337_), .B(ori_ori_n1330_), .Y(ori_ori_n1338_));
  NA4        o1310(.A(ori_ori_n1338_), .B(ori_ori_n1325_), .C(ori_ori_n1306_), .D(ori_ori_n1297_), .Y(ori_ori_n1339_));
  NO2        o1311(.A(ori_ori_n1083_), .B(ori_ori_n111_), .Y(ori_ori_n1340_));
  NO2        o1312(.A(ori_ori_n407_), .B(j), .Y(ori_ori_n1341_));
  NA2        o1313(.A(ori_ori_n1323_), .B(ori_ori_n1072_), .Y(ori_ori_n1342_));
  INV        o1314(.A(ori_ori_n1342_), .Y(ori_ori_n1343_));
  NA2        o1315(.A(ori_ori_n1341_), .B(ori_ori_n162_), .Y(ori_ori_n1344_));
  INV        o1316(.A(ori_ori_n1344_), .Y(ori_ori_n1345_));
  NO2        o1317(.A(ori_ori_n1345_), .B(ori_ori_n1343_), .Y(ori_ori_n1346_));
  INV        o1318(.A(ori_ori_n49_), .Y(ori_ori_n1347_));
  NA2        o1319(.A(ori_ori_n1347_), .B(ori_ori_n1128_), .Y(ori_ori_n1348_));
  INV        o1320(.A(ori_ori_n1348_), .Y(ori_ori_n1349_));
  NO2        o1321(.A(ori_ori_n682_), .B(ori_ori_n180_), .Y(ori_ori_n1350_));
  NO2        o1322(.A(ori_ori_n1350_), .B(ori_ori_n1349_), .Y(ori_ori_n1351_));
  NO3        o1323(.A(ori_ori_n1061_), .B(ori_ori_n1290_), .C(ori_ori_n49_), .Y(ori_ori_n1352_));
  NA3        o1324(.A(ori_ori_n1340_), .B(ori_ori_n479_), .C(f), .Y(ori_ori_n1353_));
  NO2        o1325(.A(ori_ori_n1404_), .B(ori_ori_n1353_), .Y(ori_ori_n1354_));
  NO2        o1326(.A(ori_ori_n1283_), .B(ori_ori_n178_), .Y(ori_ori_n1355_));
  NOi21      o1327(.An(d), .B(f), .Y(ori_ori_n1356_));
  NO2        o1328(.A(ori_ori_n1317_), .B(ori_ori_n40_), .Y(ori_ori_n1357_));
  NA2        o1329(.A(ori_ori_n1357_), .B(ori_ori_n1355_), .Y(ori_ori_n1358_));
  INV        o1330(.A(ori_ori_n1358_), .Y(ori_ori_n1359_));
  NO2        o1331(.A(ori_ori_n1359_), .B(ori_ori_n1354_), .Y(ori_ori_n1360_));
  NA3        o1332(.A(ori_ori_n1360_), .B(ori_ori_n1351_), .C(ori_ori_n1346_), .Y(ori_ori_n1361_));
  NA2        o1333(.A(h), .B(ori_ori_n1293_), .Y(ori_ori_n1362_));
  OAI210     o1334(.A0(ori_ori_n1331_), .A1(ori_ori_n1291_), .B0(ori_ori_n898_), .Y(ori_ori_n1363_));
  NO2        o1335(.A(ori_ori_n1048_), .B(ori_ori_n133_), .Y(ori_ori_n1364_));
  NA2        o1336(.A(ori_ori_n1364_), .B(ori_ori_n633_), .Y(ori_ori_n1365_));
  NA3        o1337(.A(ori_ori_n1365_), .B(ori_ori_n1363_), .C(ori_ori_n1362_), .Y(ori_ori_n1366_));
  NA2        o1338(.A(ori_ori_n1307_), .B(ori_ori_n1356_), .Y(ori_ori_n1367_));
  NO2        o1339(.A(ori_ori_n1367_), .B(m), .Y(ori_ori_n1368_));
  NO2        o1340(.A(ori_ori_n154_), .B(ori_ori_n185_), .Y(ori_ori_n1369_));
  OAI210     o1341(.A0(ori_ori_n1369_), .A1(ori_ori_n111_), .B0(ori_ori_n1316_), .Y(ori_ori_n1370_));
  INV        o1342(.A(ori_ori_n1370_), .Y(ori_ori_n1371_));
  NO3        o1343(.A(ori_ori_n1371_), .B(ori_ori_n1368_), .C(ori_ori_n1366_), .Y(ori_ori_n1372_));
  NO2        o1344(.A(ori_ori_n1289_), .B(e), .Y(ori_ori_n1373_));
  NA2        o1345(.A(ori_ori_n1373_), .B(ori_ori_n420_), .Y(ori_ori_n1374_));
  BUFFER     o1346(.A(ori_ori_n133_), .Y(ori_ori_n1375_));
  NO2        o1347(.A(ori_ori_n1375_), .B(ori_ori_n1374_), .Y(ori_ori_n1376_));
  NO2        o1348(.A(ori_ori_n1334_), .B(ori_ori_n366_), .Y(ori_ori_n1377_));
  NO2        o1349(.A(ori_ori_n1377_), .B(ori_ori_n1376_), .Y(ori_ori_n1378_));
  NO2        o1350(.A(ori_ori_n185_), .B(c), .Y(ori_ori_n1379_));
  OAI210     o1351(.A0(ori_ori_n1379_), .A1(ori_ori_n1373_), .B0(ori_ori_n183_), .Y(ori_ori_n1380_));
  INV        o1352(.A(ori_ori_n1380_), .Y(ori_ori_n1381_));
  AOI210     o1353(.A0(j), .A1(ori_ori_n1305_), .B0(ori_ori_n1352_), .Y(ori_ori_n1382_));
  INV        o1354(.A(ori_ori_n1080_), .Y(ori_ori_n1383_));
  OAI210     o1355(.A0(ori_ori_n1383_), .A1(ori_ori_n69_), .B0(ori_ori_n1382_), .Y(ori_ori_n1384_));
  OR2        o1356(.A(h), .B(ori_ori_n549_), .Y(ori_ori_n1385_));
  NO2        o1357(.A(ori_ori_n1385_), .B(ori_ori_n178_), .Y(ori_ori_n1386_));
  NA2        o1358(.A(ori_ori_n1060_), .B(ori_ori_n226_), .Y(ori_ori_n1387_));
  NO2        o1359(.A(ori_ori_n49_), .B(l), .Y(ori_ori_n1388_));
  INV        o1360(.A(ori_ori_n496_), .Y(ori_ori_n1389_));
  NA2        o1361(.A(ori_ori_n1389_), .B(ori_ori_n1388_), .Y(ori_ori_n1390_));
  NA2        o1362(.A(ori_ori_n1390_), .B(ori_ori_n1387_), .Y(ori_ori_n1391_));
  NO4        o1363(.A(ori_ori_n1391_), .B(ori_ori_n1386_), .C(ori_ori_n1384_), .D(ori_ori_n1381_), .Y(ori_ori_n1392_));
  NA3        o1364(.A(ori_ori_n1392_), .B(ori_ori_n1378_), .C(ori_ori_n1372_), .Y(ori_ori_n1393_));
  NA3        o1365(.A(ori_ori_n971_), .B(ori_ori_n140_), .C(ori_ori_n46_), .Y(ori_ori_n1394_));
  INV        o1366(.A(ori_ori_n163_), .Y(ori_ori_n1395_));
  NOi31      o1367(.An(ori_ori_n30_), .B(ori_ori_n1395_), .C(n), .Y(ori_ori_n1396_));
  INV        o1368(.A(ori_ori_n1396_), .Y(ori_ori_n1397_));
  NO2        o1369(.A(ori_ori_n1335_), .B(d), .Y(ori_ori_n1398_));
  NA3        o1370(.A(ori_ori_n1405_), .B(ori_ori_n1397_), .C(ori_ori_n1394_), .Y(ori_ori_n1399_));
  OR4        o1371(.A(ori_ori_n1399_), .B(ori_ori_n1393_), .C(ori_ori_n1361_), .D(ori_ori_n1339_), .Y(ori04));
  INV        o1372(.A(ori_ori_n1070_), .Y(ori05));
  INV        o1373(.A(ori_ori_n114_), .Y(ori_ori_n1404_));
  INV        o1374(.A(ori_ori_n1398_), .Y(ori_ori_n1405_));
  INV        o1375(.A(h), .Y(ori_ori_n1406_));
  ZERO       o1376(.Y(ori02));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  INV        m0023(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  INV        m0025(.A(mai_mai_n53_), .Y(mai_mai_n54_));
  AOI210     m0026(.A0(mai_mai_n54_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NAi21      m0031(.An(i), .B(h), .Y(mai_mai_n60_));
  NAi31      m0032(.An(i), .B(l), .C(j), .Y(mai_mai_n61_));
  NAi41      m0033(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n62_));
  NA2        m0034(.A(g), .B(f), .Y(mai_mai_n63_));
  NO2        m0035(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n64_));
  NAi21      m0036(.An(i), .B(j), .Y(mai_mai_n65_));
  NAi32      m0037(.An(n), .Bn(k), .C(m), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi31      m0039(.An(l), .B(m), .C(k), .Y(mai_mai_n68_));
  NAi21      m0040(.An(e), .B(h), .Y(mai_mai_n69_));
  NAi41      m0041(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n70_));
  NA2        m0042(.A(mai_mai_n67_), .B(mai_mai_n64_), .Y(mai_mai_n71_));
  INV        m0043(.A(m), .Y(mai_mai_n72_));
  NOi21      m0044(.An(k), .B(l), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  AN4        m0046(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n75_));
  NOi31      m0047(.An(h), .B(g), .C(f), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  NAi32      m0049(.An(m), .Bn(k), .C(j), .Y(mai_mai_n78_));
  NOi32      m0050(.An(h), .Bn(g), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n75_), .Y(mai_mai_n80_));
  OA220      m0052(.A0(mai_mai_n80_), .A1(mai_mai_n78_), .B0(mai_mai_n77_), .B1(mai_mai_n74_), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n81_), .B(mai_mai_n71_), .Y(mai_mai_n82_));
  INV        m0054(.A(n), .Y(mai_mai_n83_));
  NOi32      m0055(.An(e), .Bn(b), .C(d), .Y(mai_mai_n84_));
  NA2        m0056(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n85_));
  INV        m0057(.A(j), .Y(mai_mai_n86_));
  AN3        m0058(.A(m), .B(k), .C(i), .Y(mai_mai_n87_));
  NA3        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(g), .Y(mai_mai_n88_));
  NAi32      m0060(.An(g), .Bn(f), .C(h), .Y(mai_mai_n89_));
  NAi31      m0061(.An(j), .B(m), .C(l), .Y(mai_mai_n90_));
  NO2        m0062(.A(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n91_));
  NA2        m0063(.A(m), .B(l), .Y(mai_mai_n92_));
  NAi31      m0064(.An(k), .B(j), .C(g), .Y(mai_mai_n93_));
  NO3        m0065(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(f), .Y(mai_mai_n94_));
  AN2        m0066(.A(j), .B(g), .Y(mai_mai_n95_));
  NOi32      m0067(.An(m), .Bn(l), .C(i), .Y(mai_mai_n96_));
  NOi21      m0068(.An(g), .B(i), .Y(mai_mai_n97_));
  NOi32      m0069(.An(m), .Bn(j), .C(k), .Y(mai_mai_n98_));
  AOI220     m0070(.A0(mai_mai_n98_), .A1(mai_mai_n97_), .B0(mai_mai_n96_), .B1(mai_mai_n95_), .Y(mai_mai_n99_));
  NO2        m0071(.A(mai_mai_n99_), .B(f), .Y(mai_mai_n100_));
  NO3        m0072(.A(mai_mai_n100_), .B(mai_mai_n94_), .C(mai_mai_n91_), .Y(mai_mai_n101_));
  NAi41      m0073(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n102_));
  AN2        m0074(.A(e), .B(b), .Y(mai_mai_n103_));
  NOi31      m0075(.An(c), .B(h), .C(f), .Y(mai_mai_n104_));
  NA2        m0076(.A(mai_mai_n104_), .B(mai_mai_n103_), .Y(mai_mai_n105_));
  NO2        m0077(.A(mai_mai_n105_), .B(mai_mai_n102_), .Y(mai_mai_n106_));
  NOi21      m0078(.An(g), .B(f), .Y(mai_mai_n107_));
  NOi21      m0079(.An(i), .B(h), .Y(mai_mai_n108_));
  NA3        m0080(.A(mai_mai_n108_), .B(mai_mai_n107_), .C(mai_mai_n36_), .Y(mai_mai_n109_));
  INV        m0081(.A(a), .Y(mai_mai_n110_));
  NA2        m0082(.A(mai_mai_n103_), .B(mai_mai_n110_), .Y(mai_mai_n111_));
  INV        m0083(.A(l), .Y(mai_mai_n112_));
  NOi21      m0084(.An(m), .B(n), .Y(mai_mai_n113_));
  AN2        m0085(.A(k), .B(h), .Y(mai_mai_n114_));
  NO2        m0086(.A(mai_mai_n109_), .B(mai_mai_n85_), .Y(mai_mai_n115_));
  INV        m0087(.A(b), .Y(mai_mai_n116_));
  NA2        m0088(.A(l), .B(j), .Y(mai_mai_n117_));
  AN2        m0089(.A(k), .B(i), .Y(mai_mai_n118_));
  NA2        m0090(.A(mai_mai_n118_), .B(mai_mai_n117_), .Y(mai_mai_n119_));
  NA2        m0091(.A(g), .B(e), .Y(mai_mai_n120_));
  NOi32      m0092(.An(c), .Bn(a), .C(d), .Y(mai_mai_n121_));
  NA2        m0093(.A(mai_mai_n121_), .B(mai_mai_n113_), .Y(mai_mai_n122_));
  NO4        m0094(.A(mai_mai_n122_), .B(mai_mai_n120_), .C(mai_mai_n119_), .D(mai_mai_n116_), .Y(mai_mai_n123_));
  NO3        m0095(.A(mai_mai_n123_), .B(mai_mai_n115_), .C(mai_mai_n106_), .Y(mai_mai_n124_));
  OAI210     m0096(.A0(mai_mai_n101_), .A1(mai_mai_n85_), .B0(mai_mai_n124_), .Y(mai_mai_n125_));
  NOi31      m0097(.An(k), .B(m), .C(j), .Y(mai_mai_n126_));
  NA3        m0098(.A(mai_mai_n126_), .B(mai_mai_n76_), .C(mai_mai_n75_), .Y(mai_mai_n127_));
  NOi31      m0099(.An(k), .B(m), .C(i), .Y(mai_mai_n128_));
  NA3        m0100(.A(mai_mai_n128_), .B(mai_mai_n79_), .C(mai_mai_n75_), .Y(mai_mai_n129_));
  NA2        m0101(.A(mai_mai_n129_), .B(mai_mai_n127_), .Y(mai_mai_n130_));
  NOi32      m0102(.An(f), .Bn(b), .C(e), .Y(mai_mai_n131_));
  NAi21      m0103(.An(g), .B(h), .Y(mai_mai_n132_));
  NAi21      m0104(.An(m), .B(n), .Y(mai_mai_n133_));
  NAi21      m0105(.An(j), .B(k), .Y(mai_mai_n134_));
  NO3        m0106(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n132_), .Y(mai_mai_n135_));
  NAi41      m0107(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n136_));
  NAi31      m0108(.An(j), .B(k), .C(h), .Y(mai_mai_n137_));
  NO3        m0109(.A(mai_mai_n137_), .B(mai_mai_n136_), .C(mai_mai_n133_), .Y(mai_mai_n138_));
  AOI210     m0110(.A0(mai_mai_n135_), .A1(mai_mai_n131_), .B0(mai_mai_n138_), .Y(mai_mai_n139_));
  NO2        m0111(.A(k), .B(j), .Y(mai_mai_n140_));
  AN2        m0112(.A(k), .B(j), .Y(mai_mai_n141_));
  NAi21      m0113(.An(c), .B(b), .Y(mai_mai_n142_));
  NA2        m0114(.A(f), .B(d), .Y(mai_mai_n143_));
  NA2        m0115(.A(h), .B(c), .Y(mai_mai_n144_));
  NAi31      m0116(.An(f), .B(e), .C(b), .Y(mai_mai_n145_));
  NA2        m0117(.A(d), .B(b), .Y(mai_mai_n146_));
  NAi21      m0118(.An(e), .B(f), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n147_), .B(mai_mai_n146_), .Y(mai_mai_n148_));
  NA2        m0120(.A(b), .B(a), .Y(mai_mai_n149_));
  NAi21      m0121(.An(e), .B(g), .Y(mai_mai_n150_));
  NAi21      m0122(.An(c), .B(d), .Y(mai_mai_n151_));
  NAi31      m0123(.An(l), .B(k), .C(h), .Y(mai_mai_n152_));
  NO2        m0124(.A(mai_mai_n133_), .B(mai_mai_n152_), .Y(mai_mai_n153_));
  NAi21      m0125(.An(mai_mai_n130_), .B(mai_mai_n139_), .Y(mai_mai_n154_));
  NAi31      m0126(.An(e), .B(f), .C(b), .Y(mai_mai_n155_));
  NOi21      m0127(.An(g), .B(d), .Y(mai_mai_n156_));
  NO2        m0128(.A(mai_mai_n156_), .B(mai_mai_n155_), .Y(mai_mai_n157_));
  NOi21      m0129(.An(h), .B(i), .Y(mai_mai_n158_));
  NOi21      m0130(.An(k), .B(m), .Y(mai_mai_n159_));
  NA3        m0131(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(n), .Y(mai_mai_n160_));
  NOi21      m0132(.An(mai_mai_n157_), .B(mai_mai_n160_), .Y(mai_mai_n161_));
  NOi21      m0133(.An(h), .B(g), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  NAi31      m0136(.An(l), .B(j), .C(h), .Y(mai_mai_n165_));
  NOi32      m0137(.An(n), .Bn(k), .C(m), .Y(mai_mai_n166_));
  NA2        m0138(.A(l), .B(i), .Y(mai_mai_n167_));
  NA2        m0139(.A(mai_mai_n167_), .B(mai_mai_n166_), .Y(mai_mai_n168_));
  NO2        m0140(.A(mai_mai_n168_), .B(mai_mai_n164_), .Y(mai_mai_n169_));
  NAi31      m0141(.An(d), .B(f), .C(c), .Y(mai_mai_n170_));
  NAi31      m0142(.An(e), .B(f), .C(c), .Y(mai_mai_n171_));
  NA2        m0143(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  NA2        m0144(.A(j), .B(h), .Y(mai_mai_n173_));
  OR3        m0145(.A(n), .B(m), .C(k), .Y(mai_mai_n174_));
  NO2        m0146(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  NAi32      m0147(.An(m), .Bn(k), .C(n), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n176_), .B(mai_mai_n173_), .Y(mai_mai_n177_));
  AOI220     m0149(.A0(mai_mai_n177_), .A1(mai_mai_n157_), .B0(mai_mai_n175_), .B1(mai_mai_n172_), .Y(mai_mai_n178_));
  NO2        m0150(.A(n), .B(m), .Y(mai_mai_n179_));
  NA2        m0151(.A(mai_mai_n179_), .B(mai_mai_n50_), .Y(mai_mai_n180_));
  NAi21      m0152(.An(f), .B(e), .Y(mai_mai_n181_));
  NA2        m0153(.A(d), .B(c), .Y(mai_mai_n182_));
  NO2        m0154(.A(mai_mai_n182_), .B(mai_mai_n181_), .Y(mai_mai_n183_));
  NOi21      m0155(.An(mai_mai_n183_), .B(mai_mai_n180_), .Y(mai_mai_n184_));
  NAi21      m0156(.An(d), .B(c), .Y(mai_mai_n185_));
  NAi31      m0157(.An(m), .B(n), .C(b), .Y(mai_mai_n186_));
  NA2        m0158(.A(k), .B(i), .Y(mai_mai_n187_));
  NAi21      m0159(.An(h), .B(f), .Y(mai_mai_n188_));
  NO2        m0160(.A(mai_mai_n188_), .B(mai_mai_n187_), .Y(mai_mai_n189_));
  NO2        m0161(.A(mai_mai_n186_), .B(mai_mai_n151_), .Y(mai_mai_n190_));
  NA2        m0162(.A(mai_mai_n190_), .B(mai_mai_n189_), .Y(mai_mai_n191_));
  NOi32      m0163(.An(f), .Bn(c), .C(d), .Y(mai_mai_n192_));
  NOi32      m0164(.An(f), .Bn(c), .C(e), .Y(mai_mai_n193_));
  NO2        m0165(.A(mai_mai_n193_), .B(mai_mai_n192_), .Y(mai_mai_n194_));
  NO3        m0166(.A(n), .B(m), .C(j), .Y(mai_mai_n195_));
  NA2        m0167(.A(mai_mai_n195_), .B(mai_mai_n114_), .Y(mai_mai_n196_));
  AO210      m0168(.A0(mai_mai_n196_), .A1(mai_mai_n180_), .B0(mai_mai_n194_), .Y(mai_mai_n197_));
  NAi41      m0169(.An(mai_mai_n184_), .B(mai_mai_n197_), .C(mai_mai_n191_), .D(mai_mai_n178_), .Y(mai_mai_n198_));
  OR4        m0170(.A(mai_mai_n198_), .B(mai_mai_n169_), .C(mai_mai_n161_), .D(mai_mai_n154_), .Y(mai_mai_n199_));
  NO4        m0171(.A(mai_mai_n199_), .B(mai_mai_n125_), .C(mai_mai_n82_), .D(mai_mai_n55_), .Y(mai_mai_n200_));
  NA3        m0172(.A(m), .B(mai_mai_n112_), .C(j), .Y(mai_mai_n201_));
  NAi31      m0173(.An(n), .B(h), .C(g), .Y(mai_mai_n202_));
  NO2        m0174(.A(mai_mai_n202_), .B(mai_mai_n201_), .Y(mai_mai_n203_));
  NOi32      m0175(.An(m), .Bn(k), .C(l), .Y(mai_mai_n204_));
  NA3        m0176(.A(mai_mai_n204_), .B(mai_mai_n86_), .C(g), .Y(mai_mai_n205_));
  NO2        m0177(.A(mai_mai_n205_), .B(n), .Y(mai_mai_n206_));
  NOi21      m0178(.An(k), .B(j), .Y(mai_mai_n207_));
  NA4        m0179(.A(mai_mai_n207_), .B(mai_mai_n113_), .C(i), .D(g), .Y(mai_mai_n208_));
  AN2        m0180(.A(i), .B(g), .Y(mai_mai_n209_));
  NA3        m0181(.A(mai_mai_n73_), .B(mai_mai_n209_), .C(mai_mai_n113_), .Y(mai_mai_n210_));
  NA2        m0182(.A(mai_mai_n210_), .B(mai_mai_n208_), .Y(mai_mai_n211_));
  NO2        m0183(.A(mai_mai_n211_), .B(mai_mai_n203_), .Y(mai_mai_n212_));
  NAi41      m0184(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n213_));
  INV        m0185(.A(mai_mai_n213_), .Y(mai_mai_n214_));
  INV        m0186(.A(f), .Y(mai_mai_n215_));
  INV        m0187(.A(g), .Y(mai_mai_n216_));
  NOi31      m0188(.An(i), .B(j), .C(h), .Y(mai_mai_n217_));
  NOi21      m0189(.An(l), .B(m), .Y(mai_mai_n218_));
  NA2        m0190(.A(mai_mai_n218_), .B(mai_mai_n217_), .Y(mai_mai_n219_));
  NO3        m0191(.A(mai_mai_n219_), .B(mai_mai_n216_), .C(mai_mai_n215_), .Y(mai_mai_n220_));
  NA2        m0192(.A(mai_mai_n220_), .B(mai_mai_n214_), .Y(mai_mai_n221_));
  OAI210     m0193(.A0(mai_mai_n212_), .A1(mai_mai_n32_), .B0(mai_mai_n221_), .Y(mai_mai_n222_));
  NOi21      m0194(.An(n), .B(m), .Y(mai_mai_n223_));
  NOi32      m0195(.An(l), .Bn(i), .C(j), .Y(mai_mai_n224_));
  NA2        m0196(.A(mai_mai_n224_), .B(mai_mai_n223_), .Y(mai_mai_n225_));
  OA220      m0197(.A0(mai_mai_n225_), .A1(mai_mai_n105_), .B0(mai_mai_n78_), .B1(mai_mai_n77_), .Y(mai_mai_n226_));
  NAi21      m0198(.An(j), .B(h), .Y(mai_mai_n227_));
  XN2        m0199(.A(i), .B(h), .Y(mai_mai_n228_));
  NA2        m0200(.A(mai_mai_n228_), .B(mai_mai_n227_), .Y(mai_mai_n229_));
  NOi31      m0201(.An(k), .B(n), .C(m), .Y(mai_mai_n230_));
  NOi31      m0202(.An(mai_mai_n230_), .B(mai_mai_n182_), .C(mai_mai_n181_), .Y(mai_mai_n231_));
  NA2        m0203(.A(mai_mai_n231_), .B(mai_mai_n229_), .Y(mai_mai_n232_));
  NAi31      m0204(.An(f), .B(e), .C(c), .Y(mai_mai_n233_));
  NO4        m0205(.A(mai_mai_n233_), .B(mai_mai_n174_), .C(mai_mai_n173_), .D(mai_mai_n59_), .Y(mai_mai_n234_));
  NA3        m0206(.A(e), .B(c), .C(b), .Y(mai_mai_n235_));
  NAi32      m0207(.An(m), .Bn(i), .C(k), .Y(mai_mai_n236_));
  INV        m0208(.A(k), .Y(mai_mai_n237_));
  INV        m0209(.A(mai_mai_n234_), .Y(mai_mai_n238_));
  NAi21      m0210(.An(n), .B(a), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n239_), .B(mai_mai_n146_), .Y(mai_mai_n240_));
  NAi41      m0212(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n241_), .B(e), .Y(mai_mai_n242_));
  NO3        m0214(.A(mai_mai_n147_), .B(mai_mai_n93_), .C(mai_mai_n92_), .Y(mai_mai_n243_));
  OAI210     m0215(.A0(mai_mai_n243_), .A1(mai_mai_n242_), .B0(mai_mai_n240_), .Y(mai_mai_n244_));
  AN4        m0216(.A(mai_mai_n244_), .B(mai_mai_n238_), .C(mai_mai_n232_), .D(mai_mai_n226_), .Y(mai_mai_n245_));
  OR2        m0217(.A(h), .B(g), .Y(mai_mai_n246_));
  NO2        m0218(.A(mai_mai_n246_), .B(mai_mai_n102_), .Y(mai_mai_n247_));
  NA2        m0219(.A(mai_mai_n247_), .B(mai_mai_n131_), .Y(mai_mai_n248_));
  NAi41      m0220(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n249_));
  NO2        m0221(.A(mai_mai_n249_), .B(mai_mai_n215_), .Y(mai_mai_n250_));
  NA2        m0222(.A(mai_mai_n159_), .B(mai_mai_n108_), .Y(mai_mai_n251_));
  NAi21      m0223(.An(mai_mai_n251_), .B(mai_mai_n250_), .Y(mai_mai_n252_));
  NO2        m0224(.A(n), .B(a), .Y(mai_mai_n253_));
  NAi31      m0225(.An(mai_mai_n241_), .B(mai_mai_n253_), .C(mai_mai_n103_), .Y(mai_mai_n254_));
  AN2        m0226(.A(mai_mai_n254_), .B(mai_mai_n252_), .Y(mai_mai_n255_));
  NAi21      m0227(.An(h), .B(i), .Y(mai_mai_n256_));
  NA2        m0228(.A(mai_mai_n179_), .B(k), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n257_), .B(mai_mai_n256_), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n258_), .B(mai_mai_n192_), .Y(mai_mai_n259_));
  NA3        m0231(.A(mai_mai_n259_), .B(mai_mai_n255_), .C(mai_mai_n248_), .Y(mai_mai_n260_));
  NOi21      m0232(.An(g), .B(e), .Y(mai_mai_n261_));
  NO2        m0233(.A(mai_mai_n70_), .B(mai_mai_n72_), .Y(mai_mai_n262_));
  NA2        m0234(.A(mai_mai_n262_), .B(mai_mai_n261_), .Y(mai_mai_n263_));
  NOi32      m0235(.An(l), .Bn(j), .C(i), .Y(mai_mai_n264_));
  AOI210     m0236(.A0(mai_mai_n73_), .A1(mai_mai_n86_), .B0(mai_mai_n264_), .Y(mai_mai_n265_));
  NO2        m0237(.A(mai_mai_n256_), .B(mai_mai_n44_), .Y(mai_mai_n266_));
  NAi21      m0238(.An(f), .B(g), .Y(mai_mai_n267_));
  NO2        m0239(.A(mai_mai_n267_), .B(mai_mai_n62_), .Y(mai_mai_n268_));
  NO2        m0240(.A(mai_mai_n66_), .B(mai_mai_n117_), .Y(mai_mai_n269_));
  AOI220     m0241(.A0(mai_mai_n269_), .A1(mai_mai_n268_), .B0(mai_mai_n266_), .B1(mai_mai_n64_), .Y(mai_mai_n270_));
  OAI210     m0242(.A0(mai_mai_n265_), .A1(mai_mai_n263_), .B0(mai_mai_n270_), .Y(mai_mai_n271_));
  NOi41      m0243(.An(mai_mai_n245_), .B(mai_mai_n271_), .C(mai_mai_n260_), .D(mai_mai_n222_), .Y(mai_mai_n272_));
  NO4        m0244(.A(mai_mai_n203_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n273_));
  NO2        m0245(.A(mai_mai_n273_), .B(mai_mai_n111_), .Y(mai_mai_n274_));
  NA3        m0246(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n275_));
  NAi21      m0247(.An(h), .B(g), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n251_), .B(mai_mai_n267_), .Y(mai_mai_n277_));
  NAi31      m0249(.An(g), .B(k), .C(h), .Y(mai_mai_n278_));
  NO3        m0250(.A(mai_mai_n133_), .B(mai_mai_n278_), .C(l), .Y(mai_mai_n279_));
  NAi31      m0251(.An(e), .B(d), .C(a), .Y(mai_mai_n280_));
  NA2        m0252(.A(mai_mai_n279_), .B(mai_mai_n131_), .Y(mai_mai_n281_));
  INV        m0253(.A(mai_mai_n281_), .Y(mai_mai_n282_));
  NA4        m0254(.A(mai_mai_n159_), .B(mai_mai_n79_), .C(mai_mai_n75_), .D(mai_mai_n117_), .Y(mai_mai_n283_));
  NA3        m0255(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(mai_mai_n83_), .Y(mai_mai_n284_));
  NO2        m0256(.A(mai_mai_n284_), .B(mai_mai_n194_), .Y(mai_mai_n285_));
  NOi21      m0257(.An(mai_mai_n283_), .B(mai_mai_n285_), .Y(mai_mai_n286_));
  NA3        m0258(.A(e), .B(c), .C(b), .Y(mai_mai_n287_));
  NAi32      m0259(.An(k), .Bn(i), .C(j), .Y(mai_mai_n288_));
  NAi21      m0260(.An(l), .B(k), .Y(mai_mai_n289_));
  NO2        m0261(.A(mai_mai_n289_), .B(mai_mai_n49_), .Y(mai_mai_n290_));
  NOi21      m0262(.An(l), .B(j), .Y(mai_mai_n291_));
  NA2        m0263(.A(mai_mai_n162_), .B(mai_mai_n291_), .Y(mai_mai_n292_));
  NAi32      m0264(.An(j), .Bn(h), .C(i), .Y(mai_mai_n293_));
  NAi21      m0265(.An(m), .B(l), .Y(mai_mai_n294_));
  NO3        m0266(.A(mai_mai_n294_), .B(mai_mai_n293_), .C(mai_mai_n83_), .Y(mai_mai_n295_));
  NA2        m0267(.A(h), .B(g), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n166_), .B(mai_mai_n45_), .Y(mai_mai_n297_));
  NO2        m0269(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n298_));
  OAI210     m0270(.A0(mai_mai_n298_), .A1(mai_mai_n295_), .B0(mai_mai_n163_), .Y(mai_mai_n299_));
  NA2        m0271(.A(mai_mai_n299_), .B(mai_mai_n286_), .Y(mai_mai_n300_));
  NO2        m0272(.A(mai_mai_n145_), .B(d), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n301_), .B(mai_mai_n53_), .Y(mai_mai_n302_));
  NO2        m0274(.A(mai_mai_n105_), .B(mai_mai_n102_), .Y(mai_mai_n303_));
  NAi32      m0275(.An(n), .Bn(m), .C(l), .Y(mai_mai_n304_));
  NO2        m0276(.A(mai_mai_n304_), .B(mai_mai_n293_), .Y(mai_mai_n305_));
  NA2        m0277(.A(mai_mai_n305_), .B(mai_mai_n183_), .Y(mai_mai_n306_));
  NAi31      m0278(.An(k), .B(l), .C(j), .Y(mai_mai_n307_));
  OAI210     m0279(.A0(mai_mai_n289_), .A1(j), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  NOi21      m0280(.An(mai_mai_n308_), .B(mai_mai_n120_), .Y(mai_mai_n309_));
  NA2        m0281(.A(mai_mai_n306_), .B(mai_mai_n302_), .Y(mai_mai_n310_));
  NO4        m0282(.A(mai_mai_n310_), .B(mai_mai_n300_), .C(mai_mai_n282_), .D(mai_mai_n274_), .Y(mai_mai_n311_));
  NA2        m0283(.A(mai_mai_n258_), .B(mai_mai_n193_), .Y(mai_mai_n312_));
  NAi21      m0284(.An(m), .B(k), .Y(mai_mai_n313_));
  NO2        m0285(.A(mai_mai_n228_), .B(mai_mai_n313_), .Y(mai_mai_n314_));
  NAi41      m0286(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n315_));
  NO2        m0287(.A(mai_mai_n315_), .B(mai_mai_n150_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n316_), .B(mai_mai_n314_), .Y(mai_mai_n317_));
  NAi31      m0289(.An(i), .B(l), .C(h), .Y(mai_mai_n318_));
  NO4        m0290(.A(mai_mai_n318_), .B(mai_mai_n150_), .C(mai_mai_n70_), .D(mai_mai_n72_), .Y(mai_mai_n319_));
  NA2        m0291(.A(e), .B(c), .Y(mai_mai_n320_));
  NO3        m0292(.A(mai_mai_n320_), .B(n), .C(d), .Y(mai_mai_n321_));
  NOi21      m0293(.An(f), .B(h), .Y(mai_mai_n322_));
  NA2        m0294(.A(mai_mai_n322_), .B(mai_mai_n118_), .Y(mai_mai_n323_));
  NO2        m0295(.A(mai_mai_n323_), .B(mai_mai_n216_), .Y(mai_mai_n324_));
  NAi31      m0296(.An(d), .B(e), .C(b), .Y(mai_mai_n325_));
  NO2        m0297(.A(mai_mai_n133_), .B(mai_mai_n325_), .Y(mai_mai_n326_));
  NA2        m0298(.A(mai_mai_n326_), .B(mai_mai_n324_), .Y(mai_mai_n327_));
  NAi41      m0299(.An(mai_mai_n319_), .B(mai_mai_n327_), .C(mai_mai_n317_), .D(mai_mai_n312_), .Y(mai_mai_n328_));
  NO4        m0300(.A(mai_mai_n315_), .B(mai_mai_n78_), .C(mai_mai_n69_), .D(mai_mai_n216_), .Y(mai_mai_n329_));
  NA2        m0301(.A(mai_mai_n253_), .B(mai_mai_n103_), .Y(mai_mai_n330_));
  OR2        m0302(.A(mai_mai_n330_), .B(mai_mai_n205_), .Y(mai_mai_n331_));
  NOi31      m0303(.An(l), .B(n), .C(m), .Y(mai_mai_n332_));
  NA2        m0304(.A(mai_mai_n332_), .B(mai_mai_n217_), .Y(mai_mai_n333_));
  NO2        m0305(.A(mai_mai_n333_), .B(mai_mai_n194_), .Y(mai_mai_n334_));
  NAi32      m0306(.An(mai_mai_n334_), .Bn(mai_mai_n329_), .C(mai_mai_n331_), .Y(mai_mai_n335_));
  NAi32      m0307(.An(m), .Bn(j), .C(k), .Y(mai_mai_n336_));
  NAi41      m0308(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n337_));
  OAI210     m0309(.A0(mai_mai_n213_), .A1(mai_mai_n336_), .B0(mai_mai_n337_), .Y(mai_mai_n338_));
  NOi31      m0310(.An(j), .B(m), .C(k), .Y(mai_mai_n339_));
  NO2        m0311(.A(mai_mai_n126_), .B(mai_mai_n339_), .Y(mai_mai_n340_));
  AN3        m0312(.A(h), .B(g), .C(f), .Y(mai_mai_n341_));
  NAi31      m0313(.An(mai_mai_n340_), .B(mai_mai_n341_), .C(mai_mai_n338_), .Y(mai_mai_n342_));
  NOi32      m0314(.An(m), .Bn(j), .C(l), .Y(mai_mai_n343_));
  NO2        m0315(.A(mai_mai_n343_), .B(mai_mai_n96_), .Y(mai_mai_n344_));
  NAi32      m0316(.An(mai_mai_n344_), .Bn(mai_mai_n202_), .C(mai_mai_n301_), .Y(mai_mai_n345_));
  NO2        m0317(.A(mai_mai_n294_), .B(mai_mai_n293_), .Y(mai_mai_n346_));
  NO2        m0318(.A(mai_mai_n219_), .B(g), .Y(mai_mai_n347_));
  NO2        m0319(.A(mai_mai_n155_), .B(mai_mai_n83_), .Y(mai_mai_n348_));
  AOI220     m0320(.A0(mai_mai_n348_), .A1(mai_mai_n347_), .B0(mai_mai_n250_), .B1(mai_mai_n346_), .Y(mai_mai_n349_));
  NA2        m0321(.A(mai_mai_n236_), .B(mai_mai_n78_), .Y(mai_mai_n350_));
  NA3        m0322(.A(mai_mai_n350_), .B(mai_mai_n341_), .C(mai_mai_n214_), .Y(mai_mai_n351_));
  NA4        m0323(.A(mai_mai_n351_), .B(mai_mai_n349_), .C(mai_mai_n345_), .D(mai_mai_n342_), .Y(mai_mai_n352_));
  NA3        m0324(.A(h), .B(g), .C(f), .Y(mai_mai_n353_));
  NO2        m0325(.A(mai_mai_n353_), .B(mai_mai_n74_), .Y(mai_mai_n354_));
  NA2        m0326(.A(mai_mai_n337_), .B(mai_mai_n213_), .Y(mai_mai_n355_));
  NA2        m0327(.A(mai_mai_n162_), .B(e), .Y(mai_mai_n356_));
  NO2        m0328(.A(mai_mai_n356_), .B(mai_mai_n41_), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n355_), .B(mai_mai_n354_), .Y(mai_mai_n358_));
  NOi32      m0330(.An(j), .Bn(g), .C(i), .Y(mai_mai_n359_));
  NA3        m0331(.A(mai_mai_n359_), .B(mai_mai_n289_), .C(mai_mai_n113_), .Y(mai_mai_n360_));
  AO210      m0332(.A0(mai_mai_n111_), .A1(mai_mai_n32_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  NOi32      m0333(.An(e), .Bn(b), .C(a), .Y(mai_mai_n362_));
  AN2        m0334(.A(l), .B(j), .Y(mai_mai_n363_));
  NO2        m0335(.A(mai_mai_n313_), .B(mai_mai_n363_), .Y(mai_mai_n364_));
  NO3        m0336(.A(mai_mai_n315_), .B(mai_mai_n69_), .C(mai_mai_n216_), .Y(mai_mai_n365_));
  NA3        m0337(.A(mai_mai_n210_), .B(mai_mai_n208_), .C(mai_mai_n35_), .Y(mai_mai_n366_));
  AOI220     m0338(.A0(mai_mai_n366_), .A1(mai_mai_n362_), .B0(mai_mai_n365_), .B1(mai_mai_n364_), .Y(mai_mai_n367_));
  NO2        m0339(.A(mai_mai_n325_), .B(n), .Y(mai_mai_n368_));
  NA2        m0340(.A(mai_mai_n209_), .B(k), .Y(mai_mai_n369_));
  NA3        m0341(.A(m), .B(mai_mai_n112_), .C(mai_mai_n215_), .Y(mai_mai_n370_));
  NA4        m0342(.A(mai_mai_n204_), .B(mai_mai_n86_), .C(g), .D(mai_mai_n215_), .Y(mai_mai_n371_));
  OAI210     m0343(.A0(mai_mai_n370_), .A1(mai_mai_n369_), .B0(mai_mai_n371_), .Y(mai_mai_n372_));
  NAi41      m0344(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n373_));
  NA2        m0345(.A(mai_mai_n51_), .B(mai_mai_n113_), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n372_), .B(mai_mai_n368_), .Y(mai_mai_n375_));
  NA4        m0347(.A(mai_mai_n375_), .B(mai_mai_n367_), .C(mai_mai_n361_), .D(mai_mai_n358_), .Y(mai_mai_n376_));
  NO4        m0348(.A(mai_mai_n376_), .B(mai_mai_n352_), .C(mai_mai_n335_), .D(mai_mai_n328_), .Y(mai_mai_n377_));
  NA4        m0349(.A(mai_mai_n377_), .B(mai_mai_n311_), .C(mai_mai_n272_), .D(mai_mai_n200_), .Y(mai10));
  NA3        m0350(.A(m), .B(k), .C(i), .Y(mai_mai_n379_));
  NO3        m0351(.A(mai_mai_n379_), .B(j), .C(mai_mai_n216_), .Y(mai_mai_n380_));
  NOi21      m0352(.An(e), .B(f), .Y(mai_mai_n381_));
  NO4        m0353(.A(mai_mai_n151_), .B(mai_mai_n381_), .C(n), .D(mai_mai_n110_), .Y(mai_mai_n382_));
  NAi31      m0354(.An(b), .B(f), .C(c), .Y(mai_mai_n383_));
  INV        m0355(.A(mai_mai_n383_), .Y(mai_mai_n384_));
  NOi32      m0356(.An(k), .Bn(h), .C(j), .Y(mai_mai_n385_));
  NA2        m0357(.A(mai_mai_n385_), .B(mai_mai_n223_), .Y(mai_mai_n386_));
  NA2        m0358(.A(mai_mai_n160_), .B(mai_mai_n386_), .Y(mai_mai_n387_));
  NA2        m0359(.A(mai_mai_n387_), .B(mai_mai_n384_), .Y(mai_mai_n388_));
  AN2        m0360(.A(j), .B(h), .Y(mai_mai_n389_));
  NO3        m0361(.A(n), .B(m), .C(k), .Y(mai_mai_n390_));
  NA2        m0362(.A(mai_mai_n390_), .B(mai_mai_n389_), .Y(mai_mai_n391_));
  NO3        m0363(.A(mai_mai_n391_), .B(mai_mai_n151_), .C(mai_mai_n215_), .Y(mai_mai_n392_));
  OR2        m0364(.A(m), .B(k), .Y(mai_mai_n393_));
  NO2        m0365(.A(mai_mai_n173_), .B(mai_mai_n393_), .Y(mai_mai_n394_));
  NA4        m0366(.A(n), .B(f), .C(c), .D(mai_mai_n116_), .Y(mai_mai_n395_));
  NOi21      m0367(.An(mai_mai_n394_), .B(mai_mai_n395_), .Y(mai_mai_n396_));
  NOi32      m0368(.An(d), .Bn(a), .C(c), .Y(mai_mai_n397_));
  NA2        m0369(.A(mai_mai_n397_), .B(mai_mai_n181_), .Y(mai_mai_n398_));
  NAi21      m0370(.An(i), .B(g), .Y(mai_mai_n399_));
  NAi31      m0371(.An(k), .B(m), .C(j), .Y(mai_mai_n400_));
  NO3        m0372(.A(mai_mai_n400_), .B(mai_mai_n399_), .C(n), .Y(mai_mai_n401_));
  NOi21      m0373(.An(mai_mai_n401_), .B(mai_mai_n398_), .Y(mai_mai_n402_));
  NO3        m0374(.A(mai_mai_n402_), .B(mai_mai_n396_), .C(mai_mai_n392_), .Y(mai_mai_n403_));
  NO2        m0375(.A(mai_mai_n395_), .B(mai_mai_n294_), .Y(mai_mai_n404_));
  NOi32      m0376(.An(f), .Bn(d), .C(c), .Y(mai_mai_n405_));
  AOI220     m0377(.A0(mai_mai_n405_), .A1(mai_mai_n305_), .B0(mai_mai_n404_), .B1(mai_mai_n217_), .Y(mai_mai_n406_));
  NA3        m0378(.A(mai_mai_n406_), .B(mai_mai_n403_), .C(mai_mai_n388_), .Y(mai_mai_n407_));
  NO2        m0379(.A(mai_mai_n59_), .B(mai_mai_n116_), .Y(mai_mai_n408_));
  NA2        m0380(.A(mai_mai_n253_), .B(mai_mai_n408_), .Y(mai_mai_n409_));
  INV        m0381(.A(e), .Y(mai_mai_n410_));
  NA2        m0382(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n411_));
  OAI220     m0383(.A0(mai_mai_n411_), .A1(mai_mai_n201_), .B0(mai_mai_n205_), .B1(mai_mai_n410_), .Y(mai_mai_n412_));
  AN2        m0384(.A(g), .B(e), .Y(mai_mai_n413_));
  NA3        m0385(.A(mai_mai_n413_), .B(mai_mai_n204_), .C(i), .Y(mai_mai_n414_));
  OAI210     m0386(.A0(mai_mai_n88_), .A1(mai_mai_n410_), .B0(mai_mai_n414_), .Y(mai_mai_n415_));
  NO2        m0387(.A(mai_mai_n99_), .B(mai_mai_n410_), .Y(mai_mai_n416_));
  NO3        m0388(.A(mai_mai_n416_), .B(mai_mai_n415_), .C(mai_mai_n412_), .Y(mai_mai_n417_));
  NOi32      m0389(.An(h), .Bn(e), .C(g), .Y(mai_mai_n418_));
  NA3        m0390(.A(mai_mai_n418_), .B(mai_mai_n291_), .C(m), .Y(mai_mai_n419_));
  NOi21      m0391(.An(g), .B(h), .Y(mai_mai_n420_));
  AN3        m0392(.A(m), .B(l), .C(i), .Y(mai_mai_n421_));
  NA3        m0393(.A(mai_mai_n421_), .B(mai_mai_n420_), .C(e), .Y(mai_mai_n422_));
  AN3        m0394(.A(h), .B(g), .C(e), .Y(mai_mai_n423_));
  NA2        m0395(.A(mai_mai_n423_), .B(mai_mai_n96_), .Y(mai_mai_n424_));
  AN3        m0396(.A(mai_mai_n424_), .B(mai_mai_n422_), .C(mai_mai_n419_), .Y(mai_mai_n425_));
  AOI210     m0397(.A0(mai_mai_n425_), .A1(mai_mai_n417_), .B0(mai_mai_n409_), .Y(mai_mai_n426_));
  NA3        m0398(.A(mai_mai_n397_), .B(mai_mai_n181_), .C(mai_mai_n83_), .Y(mai_mai_n427_));
  NAi31      m0399(.An(b), .B(c), .C(a), .Y(mai_mai_n428_));
  NO2        m0400(.A(mai_mai_n428_), .B(n), .Y(mai_mai_n429_));
  NA2        m0401(.A(mai_mai_n51_), .B(m), .Y(mai_mai_n430_));
  NO2        m0402(.A(mai_mai_n430_), .B(mai_mai_n147_), .Y(mai_mai_n431_));
  NA2        m0403(.A(mai_mai_n431_), .B(mai_mai_n429_), .Y(mai_mai_n432_));
  INV        m0404(.A(mai_mai_n432_), .Y(mai_mai_n433_));
  NO3        m0405(.A(mai_mai_n433_), .B(mai_mai_n426_), .C(mai_mai_n407_), .Y(mai_mai_n434_));
  NA2        m0406(.A(i), .B(g), .Y(mai_mai_n435_));
  NO3        m0407(.A(mai_mai_n280_), .B(mai_mai_n435_), .C(c), .Y(mai_mai_n436_));
  NOi21      m0408(.An(a), .B(n), .Y(mai_mai_n437_));
  NOi21      m0409(.An(d), .B(c), .Y(mai_mai_n438_));
  NA2        m0410(.A(mai_mai_n438_), .B(mai_mai_n437_), .Y(mai_mai_n439_));
  NA3        m0411(.A(i), .B(g), .C(f), .Y(mai_mai_n440_));
  OR2        m0412(.A(mai_mai_n440_), .B(mai_mai_n68_), .Y(mai_mai_n441_));
  NA3        m0413(.A(mai_mai_n421_), .B(mai_mai_n420_), .C(mai_mai_n181_), .Y(mai_mai_n442_));
  AOI210     m0414(.A0(mai_mai_n442_), .A1(mai_mai_n441_), .B0(mai_mai_n439_), .Y(mai_mai_n443_));
  AOI210     m0415(.A0(mai_mai_n436_), .A1(mai_mai_n290_), .B0(mai_mai_n443_), .Y(mai_mai_n444_));
  OR2        m0416(.A(n), .B(m), .Y(mai_mai_n445_));
  NO2        m0417(.A(mai_mai_n445_), .B(mai_mai_n152_), .Y(mai_mai_n446_));
  NO2        m0418(.A(mai_mai_n182_), .B(mai_mai_n147_), .Y(mai_mai_n447_));
  OAI210     m0419(.A0(mai_mai_n446_), .A1(mai_mai_n175_), .B0(mai_mai_n447_), .Y(mai_mai_n448_));
  INV        m0420(.A(mai_mai_n374_), .Y(mai_mai_n449_));
  NA3        m0421(.A(mai_mai_n449_), .B(mai_mai_n362_), .C(d), .Y(mai_mai_n450_));
  NO2        m0422(.A(mai_mai_n428_), .B(mai_mai_n49_), .Y(mai_mai_n451_));
  NO3        m0423(.A(mai_mai_n63_), .B(mai_mai_n112_), .C(e), .Y(mai_mai_n452_));
  NAi21      m0424(.An(k), .B(j), .Y(mai_mai_n453_));
  NA2        m0425(.A(mai_mai_n256_), .B(mai_mai_n453_), .Y(mai_mai_n454_));
  NA3        m0426(.A(mai_mai_n454_), .B(mai_mai_n452_), .C(mai_mai_n451_), .Y(mai_mai_n455_));
  NAi21      m0427(.An(e), .B(d), .Y(mai_mai_n456_));
  INV        m0428(.A(mai_mai_n456_), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n257_), .B(mai_mai_n215_), .Y(mai_mai_n458_));
  NA3        m0430(.A(mai_mai_n458_), .B(mai_mai_n457_), .C(mai_mai_n229_), .Y(mai_mai_n459_));
  NA4        m0431(.A(mai_mai_n459_), .B(mai_mai_n455_), .C(mai_mai_n450_), .D(mai_mai_n448_), .Y(mai_mai_n460_));
  NO2        m0432(.A(mai_mai_n333_), .B(mai_mai_n215_), .Y(mai_mai_n461_));
  NA2        m0433(.A(mai_mai_n461_), .B(mai_mai_n457_), .Y(mai_mai_n462_));
  NOi31      m0434(.An(n), .B(m), .C(k), .Y(mai_mai_n463_));
  AOI220     m0435(.A0(mai_mai_n463_), .A1(mai_mai_n389_), .B0(mai_mai_n223_), .B1(mai_mai_n50_), .Y(mai_mai_n464_));
  NAi31      m0436(.An(g), .B(f), .C(c), .Y(mai_mai_n465_));
  OR3        m0437(.A(mai_mai_n465_), .B(mai_mai_n464_), .C(e), .Y(mai_mai_n466_));
  NA3        m0438(.A(mai_mai_n466_), .B(mai_mai_n462_), .C(mai_mai_n306_), .Y(mai_mai_n467_));
  NOi41      m0439(.An(mai_mai_n444_), .B(mai_mai_n467_), .C(mai_mai_n460_), .D(mai_mai_n271_), .Y(mai_mai_n468_));
  NOi32      m0440(.An(c), .Bn(a), .C(b), .Y(mai_mai_n469_));
  NA2        m0441(.A(mai_mai_n469_), .B(mai_mai_n113_), .Y(mai_mai_n470_));
  INV        m0442(.A(mai_mai_n278_), .Y(mai_mai_n471_));
  AN2        m0443(.A(e), .B(d), .Y(mai_mai_n472_));
  NA2        m0444(.A(mai_mai_n472_), .B(mai_mai_n471_), .Y(mai_mai_n473_));
  INV        m0445(.A(mai_mai_n147_), .Y(mai_mai_n474_));
  NO2        m0446(.A(mai_mai_n132_), .B(mai_mai_n41_), .Y(mai_mai_n475_));
  NO2        m0447(.A(mai_mai_n63_), .B(e), .Y(mai_mai_n476_));
  NOi31      m0448(.An(j), .B(k), .C(i), .Y(mai_mai_n477_));
  NOi21      m0449(.An(mai_mai_n165_), .B(mai_mai_n477_), .Y(mai_mai_n478_));
  NA4        m0450(.A(mai_mai_n318_), .B(mai_mai_n478_), .C(mai_mai_n265_), .D(mai_mai_n119_), .Y(mai_mai_n479_));
  AOI220     m0451(.A0(mai_mai_n479_), .A1(mai_mai_n476_), .B0(mai_mai_n475_), .B1(mai_mai_n474_), .Y(mai_mai_n480_));
  AOI210     m0452(.A0(mai_mai_n480_), .A1(mai_mai_n473_), .B0(mai_mai_n470_), .Y(mai_mai_n481_));
  NO2        m0453(.A(mai_mai_n211_), .B(mai_mai_n206_), .Y(mai_mai_n482_));
  NOi21      m0454(.An(a), .B(b), .Y(mai_mai_n483_));
  NA3        m0455(.A(e), .B(d), .C(c), .Y(mai_mai_n484_));
  NAi21      m0456(.An(mai_mai_n484_), .B(mai_mai_n483_), .Y(mai_mai_n485_));
  NO2        m0457(.A(mai_mai_n427_), .B(mai_mai_n205_), .Y(mai_mai_n486_));
  NOi21      m0458(.An(mai_mai_n485_), .B(mai_mai_n486_), .Y(mai_mai_n487_));
  AOI210     m0459(.A0(mai_mai_n273_), .A1(mai_mai_n482_), .B0(mai_mai_n487_), .Y(mai_mai_n488_));
  NO4        m0460(.A(mai_mai_n188_), .B(mai_mai_n102_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n489_));
  NA2        m0461(.A(mai_mai_n384_), .B(mai_mai_n153_), .Y(mai_mai_n490_));
  OR2        m0462(.A(k), .B(j), .Y(mai_mai_n491_));
  NA2        m0463(.A(l), .B(k), .Y(mai_mai_n492_));
  NA3        m0464(.A(mai_mai_n492_), .B(mai_mai_n491_), .C(mai_mai_n223_), .Y(mai_mai_n493_));
  AOI210     m0465(.A0(mai_mai_n236_), .A1(mai_mai_n336_), .B0(mai_mai_n83_), .Y(mai_mai_n494_));
  NOi21      m0466(.An(mai_mai_n493_), .B(mai_mai_n494_), .Y(mai_mai_n495_));
  OR3        m0467(.A(mai_mai_n495_), .B(mai_mai_n144_), .C(mai_mai_n136_), .Y(mai_mai_n496_));
  NA3        m0468(.A(mai_mai_n283_), .B(mai_mai_n129_), .C(mai_mai_n127_), .Y(mai_mai_n497_));
  NA2        m0469(.A(mai_mai_n397_), .B(mai_mai_n113_), .Y(mai_mai_n498_));
  NO4        m0470(.A(mai_mai_n498_), .B(mai_mai_n93_), .C(mai_mai_n112_), .D(e), .Y(mai_mai_n499_));
  NO3        m0471(.A(mai_mai_n427_), .B(mai_mai_n90_), .C(mai_mai_n132_), .Y(mai_mai_n500_));
  NO4        m0472(.A(mai_mai_n500_), .B(mai_mai_n499_), .C(mai_mai_n497_), .D(mai_mai_n319_), .Y(mai_mai_n501_));
  NA3        m0473(.A(mai_mai_n501_), .B(mai_mai_n496_), .C(mai_mai_n490_), .Y(mai_mai_n502_));
  NO4        m0474(.A(mai_mai_n502_), .B(mai_mai_n489_), .C(mai_mai_n488_), .D(mai_mai_n481_), .Y(mai_mai_n503_));
  NA2        m0475(.A(mai_mai_n67_), .B(mai_mai_n64_), .Y(mai_mai_n504_));
  NOi21      m0476(.An(d), .B(e), .Y(mai_mai_n505_));
  NO2        m0477(.A(mai_mai_n188_), .B(mai_mai_n56_), .Y(mai_mai_n506_));
  NAi31      m0478(.An(j), .B(l), .C(i), .Y(mai_mai_n507_));
  OAI210     m0479(.A0(mai_mai_n507_), .A1(mai_mai_n133_), .B0(mai_mai_n102_), .Y(mai_mai_n508_));
  NA3        m0480(.A(mai_mai_n508_), .B(mai_mai_n506_), .C(mai_mai_n505_), .Y(mai_mai_n509_));
  NO3        m0481(.A(mai_mai_n398_), .B(mai_mai_n344_), .C(mai_mai_n202_), .Y(mai_mai_n510_));
  NO2        m0482(.A(mai_mai_n398_), .B(mai_mai_n374_), .Y(mai_mai_n511_));
  NO4        m0483(.A(mai_mai_n511_), .B(mai_mai_n510_), .C(mai_mai_n184_), .D(mai_mai_n303_), .Y(mai_mai_n512_));
  NA4        m0484(.A(mai_mai_n512_), .B(mai_mai_n509_), .C(mai_mai_n504_), .D(mai_mai_n245_), .Y(mai_mai_n513_));
  OAI210     m0485(.A0(mai_mai_n128_), .A1(mai_mai_n126_), .B0(n), .Y(mai_mai_n514_));
  NO2        m0486(.A(mai_mai_n514_), .B(mai_mai_n132_), .Y(mai_mai_n515_));
  OA210      m0487(.A0(mai_mai_n247_), .A1(mai_mai_n515_), .B0(mai_mai_n193_), .Y(mai_mai_n516_));
  XO2        m0488(.A(i), .B(h), .Y(mai_mai_n517_));
  NA3        m0489(.A(mai_mai_n517_), .B(mai_mai_n159_), .C(n), .Y(mai_mai_n518_));
  NAi41      m0490(.An(mai_mai_n295_), .B(mai_mai_n518_), .C(mai_mai_n464_), .D(mai_mai_n386_), .Y(mai_mai_n519_));
  NOi32      m0491(.An(mai_mai_n519_), .Bn(mai_mai_n476_), .C(mai_mai_n275_), .Y(mai_mai_n520_));
  NAi31      m0492(.An(c), .B(f), .C(d), .Y(mai_mai_n521_));
  AOI210     m0493(.A0(mai_mai_n284_), .A1(mai_mai_n196_), .B0(mai_mai_n521_), .Y(mai_mai_n522_));
  NOi21      m0494(.An(mai_mai_n81_), .B(mai_mai_n522_), .Y(mai_mai_n523_));
  NA3        m0495(.A(mai_mai_n382_), .B(mai_mai_n96_), .C(mai_mai_n95_), .Y(mai_mai_n524_));
  NA2        m0496(.A(mai_mai_n230_), .B(mai_mai_n108_), .Y(mai_mai_n525_));
  AOI210     m0497(.A0(mai_mai_n525_), .A1(mai_mai_n180_), .B0(mai_mai_n521_), .Y(mai_mai_n526_));
  AOI210     m0498(.A0(mai_mai_n360_), .A1(mai_mai_n35_), .B0(mai_mai_n485_), .Y(mai_mai_n527_));
  NOi31      m0499(.An(mai_mai_n524_), .B(mai_mai_n527_), .C(mai_mai_n526_), .Y(mai_mai_n528_));
  NA3        m0500(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n529_));
  NO2        m0501(.A(mai_mai_n529_), .B(mai_mai_n439_), .Y(mai_mai_n530_));
  INV        m0502(.A(mai_mai_n530_), .Y(mai_mai_n531_));
  NA3        m0503(.A(mai_mai_n531_), .B(mai_mai_n528_), .C(mai_mai_n523_), .Y(mai_mai_n532_));
  NO4        m0504(.A(mai_mai_n532_), .B(mai_mai_n520_), .C(mai_mai_n516_), .D(mai_mai_n513_), .Y(mai_mai_n533_));
  NA4        m0505(.A(mai_mai_n533_), .B(mai_mai_n503_), .C(mai_mai_n468_), .D(mai_mai_n434_), .Y(mai11));
  NO2        m0506(.A(mai_mai_n70_), .B(f), .Y(mai_mai_n535_));
  NA2        m0507(.A(j), .B(g), .Y(mai_mai_n536_));
  NAi31      m0508(.An(i), .B(m), .C(l), .Y(mai_mai_n537_));
  NA3        m0509(.A(m), .B(k), .C(j), .Y(mai_mai_n538_));
  OAI220     m0510(.A0(mai_mai_n538_), .A1(mai_mai_n132_), .B0(mai_mai_n537_), .B1(mai_mai_n536_), .Y(mai_mai_n539_));
  NA2        m0511(.A(mai_mai_n539_), .B(mai_mai_n535_), .Y(mai_mai_n540_));
  NOi32      m0512(.An(e), .Bn(b), .C(f), .Y(mai_mai_n541_));
  NA2        m0513(.A(mai_mai_n264_), .B(mai_mai_n113_), .Y(mai_mai_n542_));
  NA2        m0514(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n543_));
  NO2        m0515(.A(mai_mai_n543_), .B(mai_mai_n297_), .Y(mai_mai_n544_));
  NAi31      m0516(.An(d), .B(e), .C(a), .Y(mai_mai_n545_));
  NO2        m0517(.A(mai_mai_n545_), .B(n), .Y(mai_mai_n546_));
  AOI220     m0518(.A0(mai_mai_n546_), .A1(mai_mai_n100_), .B0(mai_mai_n544_), .B1(mai_mai_n541_), .Y(mai_mai_n547_));
  NAi41      m0519(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n548_));
  AN2        m0520(.A(mai_mai_n548_), .B(mai_mai_n373_), .Y(mai_mai_n549_));
  AOI210     m0521(.A0(mai_mai_n549_), .A1(mai_mai_n398_), .B0(mai_mai_n276_), .Y(mai_mai_n550_));
  NA2        m0522(.A(j), .B(i), .Y(mai_mai_n551_));
  NAi31      m0523(.An(n), .B(m), .C(k), .Y(mai_mai_n552_));
  NO3        m0524(.A(mai_mai_n552_), .B(mai_mai_n551_), .C(mai_mai_n112_), .Y(mai_mai_n553_));
  NO4        m0525(.A(n), .B(d), .C(mai_mai_n116_), .D(a), .Y(mai_mai_n554_));
  OR2        m0526(.A(n), .B(c), .Y(mai_mai_n555_));
  NO2        m0527(.A(mai_mai_n555_), .B(mai_mai_n149_), .Y(mai_mai_n556_));
  NO2        m0528(.A(mai_mai_n556_), .B(mai_mai_n554_), .Y(mai_mai_n557_));
  NOi32      m0529(.An(g), .Bn(f), .C(i), .Y(mai_mai_n558_));
  AOI220     m0530(.A0(mai_mai_n558_), .A1(mai_mai_n98_), .B0(mai_mai_n539_), .B1(f), .Y(mai_mai_n559_));
  NO2        m0531(.A(mai_mai_n278_), .B(mai_mai_n49_), .Y(mai_mai_n560_));
  NO2        m0532(.A(mai_mai_n559_), .B(mai_mai_n557_), .Y(mai_mai_n561_));
  AOI210     m0533(.A0(mai_mai_n553_), .A1(mai_mai_n550_), .B0(mai_mai_n561_), .Y(mai_mai_n562_));
  NA2        m0534(.A(mai_mai_n141_), .B(mai_mai_n34_), .Y(mai_mai_n563_));
  OAI220     m0535(.A0(mai_mai_n563_), .A1(m), .B0(mai_mai_n543_), .B1(mai_mai_n236_), .Y(mai_mai_n564_));
  NOi41      m0536(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n565_));
  NAi32      m0537(.An(e), .Bn(b), .C(c), .Y(mai_mai_n566_));
  OR2        m0538(.A(mai_mai_n566_), .B(mai_mai_n83_), .Y(mai_mai_n567_));
  AN2        m0539(.A(mai_mai_n337_), .B(mai_mai_n315_), .Y(mai_mai_n568_));
  NA2        m0540(.A(mai_mai_n568_), .B(mai_mai_n567_), .Y(mai_mai_n569_));
  OA210      m0541(.A0(mai_mai_n569_), .A1(mai_mai_n565_), .B0(mai_mai_n564_), .Y(mai_mai_n570_));
  OAI220     m0542(.A0(mai_mai_n400_), .A1(mai_mai_n399_), .B0(mai_mai_n537_), .B1(mai_mai_n536_), .Y(mai_mai_n571_));
  NO3        m0543(.A(mai_mai_n61_), .B(mai_mai_n49_), .C(mai_mai_n216_), .Y(mai_mai_n572_));
  NO2        m0544(.A(mai_mai_n233_), .B(mai_mai_n110_), .Y(mai_mai_n573_));
  OAI210     m0545(.A0(mai_mai_n572_), .A1(mai_mai_n401_), .B0(mai_mai_n573_), .Y(mai_mai_n574_));
  INV        m0546(.A(mai_mai_n574_), .Y(mai_mai_n575_));
  NO2        m0547(.A(mai_mai_n280_), .B(n), .Y(mai_mai_n576_));
  NO2        m0548(.A(mai_mai_n429_), .B(mai_mai_n576_), .Y(mai_mai_n577_));
  NA2        m0549(.A(mai_mai_n571_), .B(f), .Y(mai_mai_n578_));
  NAi32      m0550(.An(d), .Bn(a), .C(b), .Y(mai_mai_n579_));
  NO2        m0551(.A(mai_mai_n579_), .B(mai_mai_n49_), .Y(mai_mai_n580_));
  NA2        m0552(.A(h), .B(f), .Y(mai_mai_n581_));
  NO2        m0553(.A(mai_mai_n581_), .B(mai_mai_n93_), .Y(mai_mai_n582_));
  NO3        m0554(.A(mai_mai_n176_), .B(mai_mai_n173_), .C(g), .Y(mai_mai_n583_));
  AOI220     m0555(.A0(mai_mai_n583_), .A1(mai_mai_n58_), .B0(mai_mai_n582_), .B1(mai_mai_n580_), .Y(mai_mai_n584_));
  OAI210     m0556(.A0(mai_mai_n578_), .A1(mai_mai_n577_), .B0(mai_mai_n584_), .Y(mai_mai_n585_));
  AN3        m0557(.A(j), .B(h), .C(g), .Y(mai_mai_n586_));
  NO2        m0558(.A(mai_mai_n146_), .B(c), .Y(mai_mai_n587_));
  NA3        m0559(.A(mai_mai_n587_), .B(mai_mai_n586_), .C(mai_mai_n463_), .Y(mai_mai_n588_));
  NA3        m0560(.A(f), .B(d), .C(b), .Y(mai_mai_n589_));
  INV        m0561(.A(mai_mai_n588_), .Y(mai_mai_n590_));
  NO4        m0562(.A(mai_mai_n590_), .B(mai_mai_n585_), .C(mai_mai_n575_), .D(mai_mai_n570_), .Y(mai_mai_n591_));
  AN4        m0563(.A(mai_mai_n591_), .B(mai_mai_n562_), .C(mai_mai_n547_), .D(mai_mai_n540_), .Y(mai_mai_n592_));
  INV        m0564(.A(k), .Y(mai_mai_n593_));
  NA3        m0565(.A(l), .B(mai_mai_n593_), .C(i), .Y(mai_mai_n594_));
  INV        m0566(.A(mai_mai_n594_), .Y(mai_mai_n595_));
  NA4        m0567(.A(mai_mai_n397_), .B(mai_mai_n420_), .C(mai_mai_n181_), .D(mai_mai_n113_), .Y(mai_mai_n596_));
  NAi32      m0568(.An(h), .Bn(f), .C(g), .Y(mai_mai_n597_));
  NAi41      m0569(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n598_));
  OAI210     m0570(.A0(mai_mai_n545_), .A1(n), .B0(mai_mai_n598_), .Y(mai_mai_n599_));
  NA2        m0571(.A(mai_mai_n599_), .B(m), .Y(mai_mai_n600_));
  NAi31      m0572(.An(h), .B(g), .C(f), .Y(mai_mai_n601_));
  OR3        m0573(.A(mai_mai_n601_), .B(mai_mai_n280_), .C(mai_mai_n49_), .Y(mai_mai_n602_));
  OA210      m0574(.A0(mai_mai_n600_), .A1(mai_mai_n597_), .B0(mai_mai_n602_), .Y(mai_mai_n603_));
  NO4        m0575(.A(mai_mai_n601_), .B(mai_mai_n555_), .C(mai_mai_n149_), .D(mai_mai_n72_), .Y(mai_mai_n604_));
  NAi31      m0576(.An(mai_mai_n604_), .B(mai_mai_n603_), .C(mai_mai_n596_), .Y(mai_mai_n605_));
  NAi31      m0577(.An(f), .B(h), .C(g), .Y(mai_mai_n606_));
  NO4        m0578(.A(mai_mai_n307_), .B(mai_mai_n606_), .C(mai_mai_n70_), .D(mai_mai_n72_), .Y(mai_mai_n607_));
  NOi32      m0579(.An(b), .Bn(a), .C(c), .Y(mai_mai_n608_));
  NOi32      m0580(.An(d), .Bn(a), .C(e), .Y(mai_mai_n609_));
  NA2        m0581(.A(mai_mai_n609_), .B(mai_mai_n113_), .Y(mai_mai_n610_));
  NO2        m0582(.A(n), .B(c), .Y(mai_mai_n611_));
  NA3        m0583(.A(mai_mai_n611_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n612_));
  NAi32      m0584(.An(n), .Bn(f), .C(m), .Y(mai_mai_n613_));
  NA3        m0585(.A(mai_mai_n613_), .B(mai_mai_n612_), .C(mai_mai_n610_), .Y(mai_mai_n614_));
  NOi32      m0586(.An(e), .Bn(a), .C(d), .Y(mai_mai_n615_));
  AOI210     m0587(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n615_), .Y(mai_mai_n616_));
  AOI210     m0588(.A0(mai_mai_n616_), .A1(mai_mai_n215_), .B0(mai_mai_n563_), .Y(mai_mai_n617_));
  AOI210     m0589(.A0(mai_mai_n617_), .A1(mai_mai_n614_), .B0(mai_mai_n607_), .Y(mai_mai_n618_));
  OAI210     m0590(.A0(mai_mai_n252_), .A1(mai_mai_n86_), .B0(mai_mai_n618_), .Y(mai_mai_n619_));
  AOI210     m0591(.A0(mai_mai_n605_), .A1(mai_mai_n595_), .B0(mai_mai_n619_), .Y(mai_mai_n620_));
  NO3        m0592(.A(mai_mai_n313_), .B(mai_mai_n60_), .C(n), .Y(mai_mai_n621_));
  NA3        m0593(.A(mai_mai_n521_), .B(mai_mai_n171_), .C(mai_mai_n170_), .Y(mai_mai_n622_));
  NA2        m0594(.A(mai_mai_n465_), .B(mai_mai_n233_), .Y(mai_mai_n623_));
  OR2        m0595(.A(mai_mai_n623_), .B(mai_mai_n622_), .Y(mai_mai_n624_));
  NA2        m0596(.A(mai_mai_n73_), .B(mai_mai_n113_), .Y(mai_mai_n625_));
  NO2        m0597(.A(mai_mai_n625_), .B(mai_mai_n45_), .Y(mai_mai_n626_));
  AOI220     m0598(.A0(mai_mai_n626_), .A1(mai_mai_n550_), .B0(mai_mai_n624_), .B1(mai_mai_n621_), .Y(mai_mai_n627_));
  NO2        m0599(.A(mai_mai_n627_), .B(mai_mai_n86_), .Y(mai_mai_n628_));
  NA3        m0600(.A(mai_mai_n565_), .B(mai_mai_n339_), .C(mai_mai_n46_), .Y(mai_mai_n629_));
  NOi32      m0601(.An(e), .Bn(c), .C(f), .Y(mai_mai_n630_));
  NOi21      m0602(.An(f), .B(g), .Y(mai_mai_n631_));
  NO2        m0603(.A(mai_mai_n631_), .B(mai_mai_n213_), .Y(mai_mai_n632_));
  AOI220     m0604(.A0(mai_mai_n632_), .A1(mai_mai_n394_), .B0(mai_mai_n630_), .B1(mai_mai_n175_), .Y(mai_mai_n633_));
  NA3        m0605(.A(mai_mai_n633_), .B(mai_mai_n629_), .C(mai_mai_n178_), .Y(mai_mai_n634_));
  AOI210     m0606(.A0(mai_mai_n549_), .A1(mai_mai_n398_), .B0(mai_mai_n296_), .Y(mai_mai_n635_));
  NA2        m0607(.A(mai_mai_n635_), .B(mai_mai_n269_), .Y(mai_mai_n636_));
  NOi21      m0608(.An(j), .B(l), .Y(mai_mai_n637_));
  NAi21      m0609(.An(k), .B(h), .Y(mai_mai_n638_));
  NO2        m0610(.A(mai_mai_n638_), .B(mai_mai_n267_), .Y(mai_mai_n639_));
  NA2        m0611(.A(mai_mai_n639_), .B(mai_mai_n637_), .Y(mai_mai_n640_));
  OR2        m0612(.A(mai_mai_n640_), .B(mai_mai_n600_), .Y(mai_mai_n641_));
  NOi31      m0613(.An(m), .B(n), .C(k), .Y(mai_mai_n642_));
  NO2        m0614(.A(mai_mai_n280_), .B(mai_mai_n49_), .Y(mai_mai_n643_));
  NO2        m0615(.A(mai_mai_n307_), .B(mai_mai_n606_), .Y(mai_mai_n644_));
  NO2        m0616(.A(mai_mai_n545_), .B(mai_mai_n49_), .Y(mai_mai_n645_));
  AOI220     m0617(.A0(mai_mai_n645_), .A1(mai_mai_n644_), .B0(mai_mai_n643_), .B1(mai_mai_n582_), .Y(mai_mai_n646_));
  NA3        m0618(.A(mai_mai_n646_), .B(mai_mai_n641_), .C(mai_mai_n636_), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n108_), .B(mai_mai_n36_), .Y(mai_mai_n648_));
  NO2        m0620(.A(k), .B(mai_mai_n216_), .Y(mai_mai_n649_));
  INV        m0621(.A(mai_mai_n362_), .Y(mai_mai_n650_));
  NO2        m0622(.A(mai_mai_n650_), .B(n), .Y(mai_mai_n651_));
  NAi31      m0623(.An(mai_mai_n648_), .B(mai_mai_n651_), .C(mai_mai_n649_), .Y(mai_mai_n652_));
  NO2        m0624(.A(mai_mai_n543_), .B(mai_mai_n176_), .Y(mai_mai_n653_));
  NA3        m0625(.A(mai_mai_n566_), .B(mai_mai_n275_), .C(mai_mai_n145_), .Y(mai_mai_n654_));
  NA2        m0626(.A(mai_mai_n517_), .B(mai_mai_n159_), .Y(mai_mai_n655_));
  NO3        m0627(.A(mai_mai_n395_), .B(mai_mai_n655_), .C(mai_mai_n86_), .Y(mai_mai_n656_));
  AOI210     m0628(.A0(mai_mai_n654_), .A1(mai_mai_n653_), .B0(mai_mai_n656_), .Y(mai_mai_n657_));
  AN3        m0629(.A(f), .B(d), .C(b), .Y(mai_mai_n658_));
  OAI210     m0630(.A0(mai_mai_n658_), .A1(mai_mai_n131_), .B0(n), .Y(mai_mai_n659_));
  NA3        m0631(.A(mai_mai_n517_), .B(mai_mai_n159_), .C(mai_mai_n216_), .Y(mai_mai_n660_));
  AOI210     m0632(.A0(mai_mai_n659_), .A1(mai_mai_n235_), .B0(mai_mai_n660_), .Y(mai_mai_n661_));
  NAi31      m0633(.An(m), .B(n), .C(k), .Y(mai_mai_n662_));
  INV        m0634(.A(mai_mai_n254_), .Y(mai_mai_n663_));
  OAI210     m0635(.A0(mai_mai_n663_), .A1(mai_mai_n661_), .B0(j), .Y(mai_mai_n664_));
  NA3        m0636(.A(mai_mai_n664_), .B(mai_mai_n657_), .C(mai_mai_n652_), .Y(mai_mai_n665_));
  NO4        m0637(.A(mai_mai_n665_), .B(mai_mai_n647_), .C(mai_mai_n634_), .D(mai_mai_n628_), .Y(mai_mai_n666_));
  NA2        m0638(.A(mai_mai_n382_), .B(mai_mai_n162_), .Y(mai_mai_n667_));
  NAi31      m0639(.An(g), .B(h), .C(f), .Y(mai_mai_n668_));
  OA210      m0640(.A0(mai_mai_n545_), .A1(n), .B0(mai_mai_n598_), .Y(mai_mai_n669_));
  NO2        m0641(.A(mai_mai_n669_), .B(mai_mai_n89_), .Y(mai_mai_n670_));
  INV        m0642(.A(mai_mai_n670_), .Y(mai_mai_n671_));
  AOI210     m0643(.A0(mai_mai_n671_), .A1(mai_mai_n667_), .B0(mai_mai_n538_), .Y(mai_mai_n672_));
  NO3        m0644(.A(g), .B(mai_mai_n215_), .C(mai_mai_n56_), .Y(mai_mai_n673_));
  NAi21      m0645(.An(h), .B(j), .Y(mai_mai_n674_));
  NO2        m0646(.A(mai_mai_n525_), .B(mai_mai_n86_), .Y(mai_mai_n675_));
  OAI210     m0647(.A0(mai_mai_n675_), .A1(mai_mai_n394_), .B0(mai_mai_n673_), .Y(mai_mai_n676_));
  OR2        m0648(.A(mai_mai_n70_), .B(mai_mai_n72_), .Y(mai_mai_n677_));
  AN2        m0649(.A(h), .B(f), .Y(mai_mai_n678_));
  NA2        m0650(.A(mai_mai_n678_), .B(mai_mai_n37_), .Y(mai_mai_n679_));
  NA2        m0651(.A(mai_mai_n98_), .B(mai_mai_n46_), .Y(mai_mai_n680_));
  OAI220     m0652(.A0(mai_mai_n680_), .A1(mai_mai_n330_), .B0(mai_mai_n679_), .B1(mai_mai_n470_), .Y(mai_mai_n681_));
  AOI210     m0653(.A0(mai_mai_n579_), .A1(mai_mai_n428_), .B0(mai_mai_n49_), .Y(mai_mai_n682_));
  OAI220     m0654(.A0(mai_mai_n601_), .A1(mai_mai_n594_), .B0(mai_mai_n323_), .B1(mai_mai_n536_), .Y(mai_mai_n683_));
  AOI210     m0655(.A0(mai_mai_n683_), .A1(mai_mai_n682_), .B0(mai_mai_n681_), .Y(mai_mai_n684_));
  NA2        m0656(.A(mai_mai_n684_), .B(mai_mai_n676_), .Y(mai_mai_n685_));
  NO2        m0657(.A(mai_mai_n256_), .B(f), .Y(mai_mai_n686_));
  NO2        m0658(.A(mai_mai_n631_), .B(mai_mai_n60_), .Y(mai_mai_n687_));
  NO3        m0659(.A(mai_mai_n687_), .B(mai_mai_n686_), .C(mai_mai_n34_), .Y(mai_mai_n688_));
  NA2        m0660(.A(mai_mai_n326_), .B(mai_mai_n141_), .Y(mai_mai_n689_));
  NA2        m0661(.A(mai_mai_n133_), .B(mai_mai_n49_), .Y(mai_mai_n690_));
  AOI220     m0662(.A0(mai_mai_n690_), .A1(mai_mai_n541_), .B0(mai_mai_n362_), .B1(mai_mai_n113_), .Y(mai_mai_n691_));
  OA220      m0663(.A0(mai_mai_n691_), .A1(mai_mai_n563_), .B0(mai_mai_n360_), .B1(mai_mai_n111_), .Y(mai_mai_n692_));
  OAI210     m0664(.A0(mai_mai_n689_), .A1(mai_mai_n688_), .B0(mai_mai_n692_), .Y(mai_mai_n693_));
  NO3        m0665(.A(mai_mai_n405_), .B(mai_mai_n193_), .C(mai_mai_n192_), .Y(mai_mai_n694_));
  NA2        m0666(.A(mai_mai_n694_), .B(mai_mai_n233_), .Y(mai_mai_n695_));
  NA3        m0667(.A(mai_mai_n695_), .B(mai_mai_n258_), .C(j), .Y(mai_mai_n696_));
  NO3        m0668(.A(mai_mai_n465_), .B(mai_mai_n173_), .C(i), .Y(mai_mai_n697_));
  NA2        m0669(.A(mai_mai_n469_), .B(mai_mai_n83_), .Y(mai_mai_n698_));
  NO4        m0670(.A(mai_mai_n538_), .B(mai_mai_n698_), .C(mai_mai_n132_), .D(mai_mai_n215_), .Y(mai_mai_n699_));
  INV        m0671(.A(mai_mai_n699_), .Y(mai_mai_n700_));
  NA4        m0672(.A(mai_mai_n700_), .B(mai_mai_n696_), .C(mai_mai_n524_), .D(mai_mai_n403_), .Y(mai_mai_n701_));
  NO4        m0673(.A(mai_mai_n701_), .B(mai_mai_n693_), .C(mai_mai_n685_), .D(mai_mai_n672_), .Y(mai_mai_n702_));
  NA4        m0674(.A(mai_mai_n702_), .B(mai_mai_n666_), .C(mai_mai_n620_), .D(mai_mai_n592_), .Y(mai08));
  NO2        m0675(.A(k), .B(h), .Y(mai_mai_n704_));
  AO210      m0676(.A0(mai_mai_n256_), .A1(mai_mai_n453_), .B0(mai_mai_n704_), .Y(mai_mai_n705_));
  NO2        m0677(.A(mai_mai_n705_), .B(mai_mai_n294_), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n630_), .B(mai_mai_n83_), .Y(mai_mai_n707_));
  NA2        m0679(.A(mai_mai_n707_), .B(mai_mai_n465_), .Y(mai_mai_n708_));
  AOI210     m0680(.A0(mai_mai_n708_), .A1(mai_mai_n706_), .B0(mai_mai_n500_), .Y(mai_mai_n709_));
  NA2        m0681(.A(mai_mai_n83_), .B(mai_mai_n110_), .Y(mai_mai_n710_));
  NO2        m0682(.A(mai_mai_n710_), .B(mai_mai_n57_), .Y(mai_mai_n711_));
  NO4        m0683(.A(mai_mai_n379_), .B(mai_mai_n112_), .C(j), .D(mai_mai_n216_), .Y(mai_mai_n712_));
  NA2        m0684(.A(mai_mai_n589_), .B(mai_mai_n235_), .Y(mai_mai_n713_));
  AOI220     m0685(.A0(mai_mai_n713_), .A1(mai_mai_n347_), .B0(mai_mai_n712_), .B1(mai_mai_n711_), .Y(mai_mai_n714_));
  AOI210     m0686(.A0(mai_mai_n589_), .A1(mai_mai_n155_), .B0(mai_mai_n83_), .Y(mai_mai_n715_));
  NA4        m0687(.A(mai_mai_n218_), .B(mai_mai_n141_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n716_));
  AN2        m0688(.A(l), .B(k), .Y(mai_mai_n717_));
  NO2        m0689(.A(mai_mai_n716_), .B(g), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n718_), .B(mai_mai_n715_), .Y(mai_mai_n719_));
  NA4        m0691(.A(mai_mai_n719_), .B(mai_mai_n714_), .C(mai_mai_n709_), .D(mai_mai_n349_), .Y(mai_mai_n720_));
  AN2        m0692(.A(mai_mai_n546_), .B(mai_mai_n94_), .Y(mai_mai_n721_));
  NO4        m0693(.A(mai_mai_n173_), .B(mai_mai_n393_), .C(mai_mai_n112_), .D(g), .Y(mai_mai_n722_));
  AOI210     m0694(.A0(mai_mai_n722_), .A1(mai_mai_n713_), .B0(mai_mai_n530_), .Y(mai_mai_n723_));
  NO2        m0695(.A(mai_mai_n38_), .B(mai_mai_n215_), .Y(mai_mai_n724_));
  AOI220     m0696(.A0(mai_mai_n632_), .A1(mai_mai_n346_), .B0(mai_mai_n724_), .B1(mai_mai_n576_), .Y(mai_mai_n725_));
  NAi31      m0697(.An(mai_mai_n721_), .B(mai_mai_n725_), .C(mai_mai_n723_), .Y(mai_mai_n726_));
  NO3        m0698(.A(mai_mai_n313_), .B(mai_mai_n132_), .C(mai_mai_n41_), .Y(mai_mai_n727_));
  NA2        m0699(.A(mai_mai_n705_), .B(mai_mai_n137_), .Y(mai_mai_n728_));
  AOI220     m0700(.A0(mai_mai_n728_), .A1(mai_mai_n404_), .B0(mai_mai_n727_), .B1(mai_mai_n75_), .Y(mai_mai_n729_));
  INV        m0701(.A(mai_mai_n729_), .Y(mai_mai_n730_));
  NA2        m0702(.A(mai_mai_n362_), .B(mai_mai_n43_), .Y(mai_mai_n731_));
  NA3        m0703(.A(mai_mai_n695_), .B(mai_mai_n332_), .C(mai_mai_n385_), .Y(mai_mai_n732_));
  NA2        m0704(.A(mai_mai_n717_), .B(mai_mai_n223_), .Y(mai_mai_n733_));
  NO2        m0705(.A(mai_mai_n733_), .B(mai_mai_n325_), .Y(mai_mai_n734_));
  AOI210     m0706(.A0(mai_mai_n734_), .A1(mai_mai_n686_), .B0(mai_mai_n499_), .Y(mai_mai_n735_));
  NA3        m0707(.A(m), .B(l), .C(k), .Y(mai_mai_n736_));
  NO2        m0708(.A(mai_mai_n548_), .B(mai_mai_n276_), .Y(mai_mai_n737_));
  NOi21      m0709(.An(mai_mai_n737_), .B(mai_mai_n542_), .Y(mai_mai_n738_));
  NA4        m0710(.A(mai_mai_n113_), .B(l), .C(k), .D(mai_mai_n86_), .Y(mai_mai_n739_));
  NA3        m0711(.A(mai_mai_n121_), .B(mai_mai_n413_), .C(i), .Y(mai_mai_n740_));
  NO2        m0712(.A(mai_mai_n740_), .B(mai_mai_n739_), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n741_), .B(mai_mai_n738_), .Y(mai_mai_n742_));
  NA4        m0714(.A(mai_mai_n742_), .B(mai_mai_n735_), .C(mai_mai_n732_), .D(mai_mai_n731_), .Y(mai_mai_n743_));
  NO4        m0715(.A(mai_mai_n743_), .B(mai_mai_n730_), .C(mai_mai_n726_), .D(mai_mai_n720_), .Y(mai_mai_n744_));
  NA2        m0716(.A(mai_mai_n632_), .B(mai_mai_n394_), .Y(mai_mai_n745_));
  NOi31      m0717(.An(g), .B(h), .C(f), .Y(mai_mai_n746_));
  NA2        m0718(.A(mai_mai_n645_), .B(mai_mai_n746_), .Y(mai_mai_n747_));
  AO210      m0719(.A0(mai_mai_n747_), .A1(mai_mai_n602_), .B0(mai_mai_n551_), .Y(mai_mai_n748_));
  NO3        m0720(.A(mai_mai_n398_), .B(mai_mai_n536_), .C(h), .Y(mai_mai_n749_));
  AOI210     m0721(.A0(mai_mai_n749_), .A1(mai_mai_n113_), .B0(mai_mai_n511_), .Y(mai_mai_n750_));
  NA4        m0722(.A(mai_mai_n750_), .B(mai_mai_n748_), .C(mai_mai_n745_), .D(mai_mai_n255_), .Y(mai_mai_n751_));
  NA2        m0723(.A(mai_mai_n717_), .B(mai_mai_n72_), .Y(mai_mai_n752_));
  NO4        m0724(.A(mai_mai_n694_), .B(mai_mai_n173_), .C(n), .D(i), .Y(mai_mai_n753_));
  NOi21      m0725(.An(h), .B(j), .Y(mai_mai_n754_));
  NA2        m0726(.A(mai_mai_n754_), .B(f), .Y(mai_mai_n755_));
  NO2        m0727(.A(mai_mai_n755_), .B(mai_mai_n249_), .Y(mai_mai_n756_));
  NO3        m0728(.A(mai_mai_n756_), .B(mai_mai_n753_), .C(mai_mai_n697_), .Y(mai_mai_n757_));
  OAI220     m0729(.A0(mai_mai_n757_), .A1(mai_mai_n752_), .B0(mai_mai_n602_), .B1(mai_mai_n61_), .Y(mai_mai_n758_));
  AOI210     m0730(.A0(mai_mai_n751_), .A1(l), .B0(mai_mai_n758_), .Y(mai_mai_n759_));
  NO2        m0731(.A(j), .B(i), .Y(mai_mai_n760_));
  NA3        m0732(.A(mai_mai_n760_), .B(mai_mai_n79_), .C(l), .Y(mai_mai_n761_));
  NA2        m0733(.A(mai_mai_n760_), .B(mai_mai_n33_), .Y(mai_mai_n762_));
  OR2        m0734(.A(mai_mai_n761_), .B(mai_mai_n600_), .Y(mai_mai_n763_));
  NO3        m0735(.A(mai_mai_n151_), .B(mai_mai_n49_), .C(mai_mai_n110_), .Y(mai_mai_n764_));
  NO3        m0736(.A(mai_mai_n555_), .B(mai_mai_n149_), .C(mai_mai_n72_), .Y(mai_mai_n765_));
  NO3        m0737(.A(mai_mai_n492_), .B(mai_mai_n440_), .C(j), .Y(mai_mai_n766_));
  OAI210     m0738(.A0(mai_mai_n765_), .A1(mai_mai_n764_), .B0(mai_mai_n766_), .Y(mai_mai_n767_));
  OAI210     m0739(.A0(mai_mai_n747_), .A1(mai_mai_n61_), .B0(mai_mai_n767_), .Y(mai_mai_n768_));
  NA2        m0740(.A(k), .B(j), .Y(mai_mai_n769_));
  NO3        m0741(.A(mai_mai_n294_), .B(mai_mai_n769_), .C(mai_mai_n40_), .Y(mai_mai_n770_));
  AOI210     m0742(.A0(mai_mai_n541_), .A1(n), .B0(mai_mai_n565_), .Y(mai_mai_n771_));
  NA2        m0743(.A(mai_mai_n771_), .B(mai_mai_n568_), .Y(mai_mai_n772_));
  AN3        m0744(.A(mai_mai_n772_), .B(mai_mai_n770_), .C(mai_mai_n97_), .Y(mai_mai_n773_));
  NO3        m0745(.A(mai_mai_n173_), .B(mai_mai_n393_), .C(mai_mai_n112_), .Y(mai_mai_n774_));
  AOI220     m0746(.A0(mai_mai_n774_), .A1(mai_mai_n250_), .B0(mai_mai_n623_), .B1(mai_mai_n305_), .Y(mai_mai_n775_));
  NAi31      m0747(.An(mai_mai_n616_), .B(mai_mai_n91_), .C(mai_mai_n83_), .Y(mai_mai_n776_));
  NA2        m0748(.A(mai_mai_n776_), .B(mai_mai_n775_), .Y(mai_mai_n777_));
  NO2        m0749(.A(mai_mai_n294_), .B(mai_mai_n137_), .Y(mai_mai_n778_));
  AOI220     m0750(.A0(mai_mai_n778_), .A1(mai_mai_n632_), .B0(mai_mai_n727_), .B1(mai_mai_n715_), .Y(mai_mai_n779_));
  NO2        m0751(.A(mai_mai_n736_), .B(mai_mai_n89_), .Y(mai_mai_n780_));
  NA2        m0752(.A(mai_mai_n780_), .B(mai_mai_n599_), .Y(mai_mai_n781_));
  NO2        m0753(.A(mai_mai_n601_), .B(mai_mai_n117_), .Y(mai_mai_n782_));
  OAI210     m0754(.A0(mai_mai_n782_), .A1(mai_mai_n766_), .B0(mai_mai_n682_), .Y(mai_mai_n783_));
  NA3        m0755(.A(mai_mai_n783_), .B(mai_mai_n781_), .C(mai_mai_n779_), .Y(mai_mai_n784_));
  OR4        m0756(.A(mai_mai_n784_), .B(mai_mai_n777_), .C(mai_mai_n773_), .D(mai_mai_n768_), .Y(mai_mai_n785_));
  NA3        m0757(.A(mai_mai_n771_), .B(mai_mai_n568_), .C(mai_mai_n567_), .Y(mai_mai_n786_));
  NA4        m0758(.A(mai_mai_n786_), .B(mai_mai_n218_), .C(mai_mai_n453_), .D(mai_mai_n34_), .Y(mai_mai_n787_));
  OAI220     m0759(.A0(mai_mai_n716_), .A1(mai_mai_n707_), .B0(mai_mai_n330_), .B1(mai_mai_n38_), .Y(mai_mai_n788_));
  INV        m0760(.A(mai_mai_n788_), .Y(mai_mai_n789_));
  NA3        m0761(.A(mai_mai_n558_), .B(mai_mai_n291_), .C(h), .Y(mai_mai_n790_));
  NOi21      m0762(.An(mai_mai_n682_), .B(mai_mai_n790_), .Y(mai_mai_n791_));
  NO2        m0763(.A(mai_mai_n90_), .B(mai_mai_n47_), .Y(mai_mai_n792_));
  OAI220     m0764(.A0(mai_mai_n790_), .A1(mai_mai_n612_), .B0(mai_mai_n761_), .B1(mai_mai_n677_), .Y(mai_mai_n793_));
  AOI210     m0765(.A0(mai_mai_n792_), .A1(mai_mai_n651_), .B0(mai_mai_n793_), .Y(mai_mai_n794_));
  NAi41      m0766(.An(mai_mai_n791_), .B(mai_mai_n794_), .C(mai_mai_n789_), .D(mai_mai_n787_), .Y(mai_mai_n795_));
  OR2        m0767(.A(mai_mai_n780_), .B(mai_mai_n94_), .Y(mai_mai_n796_));
  AOI220     m0768(.A0(mai_mai_n796_), .A1(mai_mai_n240_), .B0(mai_mai_n766_), .B1(mai_mai_n643_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n669_), .B(mai_mai_n72_), .Y(mai_mai_n798_));
  INV        m0770(.A(mai_mai_n334_), .Y(mai_mai_n799_));
  OAI210     m0771(.A0(mai_mai_n736_), .A1(mai_mai_n668_), .B0(mai_mai_n529_), .Y(mai_mai_n800_));
  NA3        m0772(.A(mai_mai_n253_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n801_));
  AOI220     m0773(.A0(mai_mai_n611_), .A1(mai_mai_n29_), .B0(mai_mai_n469_), .B1(mai_mai_n83_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n802_), .B(mai_mai_n801_), .Y(mai_mai_n803_));
  NO2        m0775(.A(mai_mai_n790_), .B(mai_mai_n498_), .Y(mai_mai_n804_));
  AOI210     m0776(.A0(mai_mai_n803_), .A1(mai_mai_n800_), .B0(mai_mai_n804_), .Y(mai_mai_n805_));
  NA3        m0777(.A(mai_mai_n805_), .B(mai_mai_n799_), .C(mai_mai_n797_), .Y(mai_mai_n806_));
  NOi41      m0778(.An(mai_mai_n763_), .B(mai_mai_n806_), .C(mai_mai_n795_), .D(mai_mai_n785_), .Y(mai_mai_n807_));
  NO3        m0779(.A(mai_mai_n340_), .B(mai_mai_n296_), .C(mai_mai_n112_), .Y(mai_mai_n808_));
  NA2        m0780(.A(mai_mai_n808_), .B(mai_mai_n772_), .Y(mai_mai_n809_));
  NO3        m0781(.A(mai_mai_n536_), .B(mai_mai_n92_), .C(h), .Y(mai_mai_n810_));
  NA2        m0782(.A(mai_mai_n810_), .B(mai_mai_n711_), .Y(mai_mai_n811_));
  NA3        m0783(.A(mai_mai_n811_), .B(mai_mai_n809_), .C(mai_mai_n406_), .Y(mai_mai_n812_));
  OR2        m0784(.A(mai_mai_n668_), .B(mai_mai_n90_), .Y(mai_mai_n813_));
  NOi31      m0785(.An(b), .B(d), .C(a), .Y(mai_mai_n814_));
  NO2        m0786(.A(mai_mai_n814_), .B(mai_mai_n609_), .Y(mai_mai_n815_));
  NO2        m0787(.A(mai_mai_n815_), .B(n), .Y(mai_mai_n816_));
  NOi21      m0788(.An(mai_mai_n802_), .B(mai_mai_n816_), .Y(mai_mai_n817_));
  OAI220     m0789(.A0(mai_mai_n817_), .A1(mai_mai_n813_), .B0(mai_mai_n790_), .B1(mai_mai_n610_), .Y(mai_mai_n818_));
  NO2        m0790(.A(mai_mai_n566_), .B(mai_mai_n83_), .Y(mai_mai_n819_));
  NO3        m0791(.A(mai_mai_n631_), .B(mai_mai_n325_), .C(mai_mai_n117_), .Y(mai_mai_n820_));
  NOi21      m0792(.An(mai_mai_n820_), .B(mai_mai_n160_), .Y(mai_mai_n821_));
  AOI210     m0793(.A0(mai_mai_n808_), .A1(mai_mai_n819_), .B0(mai_mai_n821_), .Y(mai_mai_n822_));
  OAI210     m0794(.A0(mai_mai_n716_), .A1(mai_mai_n395_), .B0(mai_mai_n822_), .Y(mai_mai_n823_));
  NO2        m0795(.A(mai_mai_n694_), .B(n), .Y(mai_mai_n824_));
  AOI220     m0796(.A0(mai_mai_n778_), .A1(mai_mai_n673_), .B0(mai_mai_n824_), .B1(mai_mai_n706_), .Y(mai_mai_n825_));
  NO2        m0797(.A(mai_mai_n320_), .B(mai_mai_n239_), .Y(mai_mai_n826_));
  OAI210     m0798(.A0(mai_mai_n94_), .A1(mai_mai_n91_), .B0(mai_mai_n826_), .Y(mai_mai_n827_));
  NA2        m0799(.A(mai_mai_n121_), .B(mai_mai_n83_), .Y(mai_mai_n828_));
  INV        m0800(.A(mai_mai_n827_), .Y(mai_mai_n829_));
  NA2        m0801(.A(mai_mai_n734_), .B(mai_mai_n34_), .Y(mai_mai_n830_));
  NAi21      m0802(.An(mai_mai_n739_), .B(mai_mai_n436_), .Y(mai_mai_n831_));
  NO2        m0803(.A(mai_mai_n276_), .B(i), .Y(mai_mai_n832_));
  NA2        m0804(.A(mai_mai_n722_), .B(mai_mai_n348_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n604_), .B(mai_mai_n363_), .Y(mai_mai_n834_));
  AN3        m0806(.A(mai_mai_n834_), .B(mai_mai_n833_), .C(mai_mai_n831_), .Y(mai_mai_n835_));
  NAi41      m0807(.An(mai_mai_n829_), .B(mai_mai_n835_), .C(mai_mai_n830_), .D(mai_mai_n825_), .Y(mai_mai_n836_));
  NO4        m0808(.A(mai_mai_n836_), .B(mai_mai_n823_), .C(mai_mai_n818_), .D(mai_mai_n812_), .Y(mai_mai_n837_));
  NA4        m0809(.A(mai_mai_n837_), .B(mai_mai_n807_), .C(mai_mai_n759_), .D(mai_mai_n744_), .Y(mai09));
  INV        m0810(.A(mai_mai_n122_), .Y(mai_mai_n839_));
  NA2        m0811(.A(f), .B(e), .Y(mai_mai_n840_));
  NO2        m0812(.A(mai_mai_n228_), .B(mai_mai_n112_), .Y(mai_mai_n841_));
  NA2        m0813(.A(mai_mai_n841_), .B(g), .Y(mai_mai_n842_));
  NA4        m0814(.A(mai_mai_n307_), .B(mai_mai_n478_), .C(mai_mai_n265_), .D(mai_mai_n119_), .Y(mai_mai_n843_));
  AOI210     m0815(.A0(mai_mai_n843_), .A1(g), .B0(mai_mai_n475_), .Y(mai_mai_n844_));
  AOI210     m0816(.A0(mai_mai_n844_), .A1(mai_mai_n842_), .B0(mai_mai_n840_), .Y(mai_mai_n845_));
  NA2        m0817(.A(mai_mai_n446_), .B(e), .Y(mai_mai_n846_));
  NO2        m0818(.A(mai_mai_n846_), .B(mai_mai_n521_), .Y(mai_mai_n847_));
  AOI210     m0819(.A0(mai_mai_n845_), .A1(mai_mai_n839_), .B0(mai_mai_n847_), .Y(mai_mai_n848_));
  NA3        m0820(.A(m), .B(l), .C(i), .Y(mai_mai_n849_));
  OAI220     m0821(.A0(mai_mai_n601_), .A1(mai_mai_n849_), .B0(mai_mai_n353_), .B1(mai_mai_n537_), .Y(mai_mai_n850_));
  NA4        m0822(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(g), .D(f), .Y(mai_mai_n851_));
  NAi31      m0823(.An(mai_mai_n850_), .B(mai_mai_n851_), .C(mai_mai_n441_), .Y(mai_mai_n852_));
  NA3        m0824(.A(mai_mai_n813_), .B(mai_mai_n578_), .C(mai_mai_n529_), .Y(mai_mai_n853_));
  OA210      m0825(.A0(mai_mai_n853_), .A1(mai_mai_n852_), .B0(mai_mai_n816_), .Y(mai_mai_n854_));
  INV        m0826(.A(mai_mai_n337_), .Y(mai_mai_n855_));
  NO2        m0827(.A(mai_mai_n128_), .B(mai_mai_n126_), .Y(mai_mai_n856_));
  NOi31      m0828(.An(k), .B(m), .C(l), .Y(mai_mai_n857_));
  NO2        m0829(.A(mai_mai_n339_), .B(mai_mai_n857_), .Y(mai_mai_n858_));
  AOI210     m0830(.A0(mai_mai_n858_), .A1(mai_mai_n856_), .B0(mai_mai_n606_), .Y(mai_mai_n859_));
  NA2        m0831(.A(mai_mai_n801_), .B(mai_mai_n330_), .Y(mai_mai_n860_));
  NA2        m0832(.A(mai_mai_n341_), .B(mai_mai_n343_), .Y(mai_mai_n861_));
  OAI210     m0833(.A0(mai_mai_n205_), .A1(mai_mai_n215_), .B0(mai_mai_n861_), .Y(mai_mai_n862_));
  AOI220     m0834(.A0(mai_mai_n862_), .A1(mai_mai_n860_), .B0(mai_mai_n859_), .B1(mai_mai_n855_), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n167_), .B(mai_mai_n114_), .Y(mai_mai_n864_));
  NA3        m0836(.A(mai_mai_n864_), .B(mai_mai_n705_), .C(mai_mai_n137_), .Y(mai_mai_n865_));
  NA3        m0837(.A(mai_mai_n865_), .B(mai_mai_n190_), .C(mai_mai_n31_), .Y(mai_mai_n866_));
  NA4        m0838(.A(mai_mai_n866_), .B(mai_mai_n863_), .C(mai_mai_n633_), .D(mai_mai_n81_), .Y(mai_mai_n867_));
  NOi21      m0839(.An(f), .B(d), .Y(mai_mai_n868_));
  NA2        m0840(.A(mai_mai_n868_), .B(m), .Y(mai_mai_n869_));
  NO2        m0841(.A(mai_mai_n869_), .B(mai_mai_n52_), .Y(mai_mai_n870_));
  NOi32      m0842(.An(g), .Bn(f), .C(d), .Y(mai_mai_n871_));
  NA4        m0843(.A(mai_mai_n871_), .B(mai_mai_n611_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n870_), .B(mai_mai_n556_), .Y(mai_mai_n873_));
  NA3        m0845(.A(mai_mai_n307_), .B(mai_mai_n265_), .C(mai_mai_n119_), .Y(mai_mai_n874_));
  AN2        m0846(.A(f), .B(d), .Y(mai_mai_n875_));
  NA3        m0847(.A(mai_mai_n483_), .B(mai_mai_n875_), .C(mai_mai_n83_), .Y(mai_mai_n876_));
  NO3        m0848(.A(mai_mai_n876_), .B(mai_mai_n72_), .C(mai_mai_n216_), .Y(mai_mai_n877_));
  NO2        m0849(.A(mai_mai_n288_), .B(mai_mai_n56_), .Y(mai_mai_n878_));
  NA2        m0850(.A(mai_mai_n874_), .B(mai_mai_n877_), .Y(mai_mai_n879_));
  NAi31      m0851(.An(mai_mai_n497_), .B(mai_mai_n879_), .C(mai_mai_n873_), .Y(mai_mai_n880_));
  NO4        m0852(.A(mai_mai_n631_), .B(mai_mai_n133_), .C(mai_mai_n325_), .D(mai_mai_n152_), .Y(mai_mai_n881_));
  NO2        m0853(.A(mai_mai_n662_), .B(mai_mai_n325_), .Y(mai_mai_n882_));
  AN2        m0854(.A(mai_mai_n882_), .B(mai_mai_n686_), .Y(mai_mai_n883_));
  NO2        m0855(.A(mai_mai_n883_), .B(mai_mai_n881_), .Y(mai_mai_n884_));
  NA2        m0856(.A(mai_mai_n609_), .B(mai_mai_n83_), .Y(mai_mai_n885_));
  NA3        m0857(.A(mai_mai_n159_), .B(mai_mai_n108_), .C(mai_mai_n107_), .Y(mai_mai_n886_));
  OAI220     m0858(.A0(mai_mai_n876_), .A1(mai_mai_n430_), .B0(mai_mai_n337_), .B1(mai_mai_n886_), .Y(mai_mai_n887_));
  NOi31      m0859(.An(mai_mai_n226_), .B(mai_mai_n887_), .C(mai_mai_n303_), .Y(mai_mai_n888_));
  NA2        m0860(.A(c), .B(mai_mai_n116_), .Y(mai_mai_n889_));
  NO2        m0861(.A(mai_mai_n889_), .B(mai_mai_n410_), .Y(mai_mai_n890_));
  NA3        m0862(.A(mai_mai_n890_), .B(mai_mai_n519_), .C(f), .Y(mai_mai_n891_));
  OR2        m0863(.A(mai_mai_n668_), .B(mai_mai_n552_), .Y(mai_mai_n892_));
  INV        m0864(.A(mai_mai_n892_), .Y(mai_mai_n893_));
  NA2        m0865(.A(mai_mai_n815_), .B(mai_mai_n111_), .Y(mai_mai_n894_));
  NA2        m0866(.A(mai_mai_n894_), .B(mai_mai_n893_), .Y(mai_mai_n895_));
  NA4        m0867(.A(mai_mai_n895_), .B(mai_mai_n891_), .C(mai_mai_n888_), .D(mai_mai_n884_), .Y(mai_mai_n896_));
  NO4        m0868(.A(mai_mai_n896_), .B(mai_mai_n880_), .C(mai_mai_n867_), .D(mai_mai_n854_), .Y(mai_mai_n897_));
  OR2        m0869(.A(mai_mai_n876_), .B(mai_mai_n72_), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n112_), .B(j), .Y(mai_mai_n899_));
  NA2        m0871(.A(mai_mai_n841_), .B(g), .Y(mai_mai_n900_));
  AOI210     m0872(.A0(mai_mai_n900_), .A1(mai_mai_n292_), .B0(mai_mai_n898_), .Y(mai_mai_n901_));
  NO2        m0873(.A(mai_mai_n330_), .B(mai_mai_n851_), .Y(mai_mai_n902_));
  NO2        m0874(.A(mai_mai_n233_), .B(mai_mai_n227_), .Y(mai_mai_n903_));
  NA2        m0875(.A(mai_mai_n903_), .B(mai_mai_n230_), .Y(mai_mai_n904_));
  NO2        m0876(.A(mai_mai_n430_), .B(mai_mai_n840_), .Y(mai_mai_n905_));
  INV        m0877(.A(mai_mai_n904_), .Y(mai_mai_n906_));
  NA2        m0878(.A(e), .B(d), .Y(mai_mai_n907_));
  OAI220     m0879(.A0(mai_mai_n907_), .A1(c), .B0(mai_mai_n320_), .B1(d), .Y(mai_mai_n908_));
  NA3        m0880(.A(mai_mai_n908_), .B(mai_mai_n458_), .C(mai_mai_n517_), .Y(mai_mai_n909_));
  AOI210     m0881(.A0(mai_mai_n525_), .A1(mai_mai_n180_), .B0(mai_mai_n233_), .Y(mai_mai_n910_));
  AOI210     m0882(.A0(mai_mai_n632_), .A1(mai_mai_n346_), .B0(mai_mai_n910_), .Y(mai_mai_n911_));
  NA2        m0883(.A(mai_mai_n288_), .B(mai_mai_n165_), .Y(mai_mai_n912_));
  NA2        m0884(.A(mai_mai_n877_), .B(mai_mai_n912_), .Y(mai_mai_n913_));
  NA3        m0885(.A(mai_mai_n166_), .B(mai_mai_n84_), .C(mai_mai_n34_), .Y(mai_mai_n914_));
  NA4        m0886(.A(mai_mai_n914_), .B(mai_mai_n913_), .C(mai_mai_n911_), .D(mai_mai_n909_), .Y(mai_mai_n915_));
  NO4        m0887(.A(mai_mai_n915_), .B(mai_mai_n906_), .C(mai_mai_n902_), .D(mai_mai_n901_), .Y(mai_mai_n916_));
  NA2        m0888(.A(mai_mai_n855_), .B(mai_mai_n31_), .Y(mai_mai_n917_));
  AO210      m0889(.A0(mai_mai_n917_), .A1(mai_mai_n707_), .B0(mai_mai_n219_), .Y(mai_mai_n918_));
  OAI220     m0890(.A0(mai_mai_n631_), .A1(mai_mai_n60_), .B0(mai_mai_n296_), .B1(j), .Y(mai_mai_n919_));
  AOI220     m0891(.A0(mai_mai_n919_), .A1(mai_mai_n882_), .B0(mai_mai_n621_), .B1(mai_mai_n630_), .Y(mai_mai_n920_));
  OAI210     m0892(.A0(mai_mai_n846_), .A1(mai_mai_n170_), .B0(mai_mai_n920_), .Y(mai_mai_n921_));
  OAI210     m0893(.A0(mai_mai_n841_), .A1(mai_mai_n912_), .B0(mai_mai_n871_), .Y(mai_mai_n922_));
  NO2        m0894(.A(mai_mai_n922_), .B(mai_mai_n612_), .Y(mai_mai_n923_));
  AOI210     m0895(.A0(mai_mai_n118_), .A1(mai_mai_n117_), .B0(mai_mai_n264_), .Y(mai_mai_n924_));
  NO2        m0896(.A(mai_mai_n924_), .B(mai_mai_n872_), .Y(mai_mai_n925_));
  AO210      m0897(.A0(mai_mai_n860_), .A1(mai_mai_n850_), .B0(mai_mai_n925_), .Y(mai_mai_n926_));
  NO3        m0898(.A(mai_mai_n926_), .B(mai_mai_n923_), .C(mai_mai_n921_), .Y(mai_mai_n927_));
  AO220      m0899(.A0(mai_mai_n458_), .A1(mai_mai_n754_), .B0(mai_mai_n175_), .B1(f), .Y(mai_mai_n928_));
  OAI210     m0900(.A0(mai_mai_n928_), .A1(mai_mai_n461_), .B0(mai_mai_n908_), .Y(mai_mai_n929_));
  NO2        m0901(.A(mai_mai_n440_), .B(mai_mai_n68_), .Y(mai_mai_n930_));
  OAI210     m0902(.A0(mai_mai_n853_), .A1(mai_mai_n930_), .B0(mai_mai_n711_), .Y(mai_mai_n931_));
  AN4        m0903(.A(mai_mai_n931_), .B(mai_mai_n929_), .C(mai_mai_n927_), .D(mai_mai_n918_), .Y(mai_mai_n932_));
  NA4        m0904(.A(mai_mai_n932_), .B(mai_mai_n916_), .C(mai_mai_n897_), .D(mai_mai_n848_), .Y(mai12));
  NO2        m0905(.A(mai_mai_n456_), .B(c), .Y(mai_mai_n934_));
  NO4        m0906(.A(mai_mai_n445_), .B(mai_mai_n256_), .C(mai_mai_n593_), .D(mai_mai_n216_), .Y(mai_mai_n935_));
  NA2        m0907(.A(mai_mai_n935_), .B(mai_mai_n934_), .Y(mai_mai_n936_));
  NA2        m0908(.A(mai_mai_n556_), .B(mai_mai_n930_), .Y(mai_mai_n937_));
  NO2        m0909(.A(mai_mai_n456_), .B(mai_mai_n116_), .Y(mai_mai_n938_));
  NO2        m0910(.A(mai_mai_n856_), .B(mai_mai_n353_), .Y(mai_mai_n939_));
  NO2        m0911(.A(mai_mai_n668_), .B(mai_mai_n379_), .Y(mai_mai_n940_));
  AOI220     m0912(.A0(mai_mai_n940_), .A1(mai_mai_n554_), .B0(mai_mai_n939_), .B1(mai_mai_n938_), .Y(mai_mai_n941_));
  NA4        m0913(.A(mai_mai_n941_), .B(mai_mai_n937_), .C(mai_mai_n936_), .D(mai_mai_n444_), .Y(mai_mai_n942_));
  AOI210     m0914(.A0(mai_mai_n236_), .A1(mai_mai_n336_), .B0(mai_mai_n202_), .Y(mai_mai_n943_));
  OR2        m0915(.A(mai_mai_n943_), .B(mai_mai_n935_), .Y(mai_mai_n944_));
  AOI210     m0916(.A0(mai_mai_n333_), .A1(mai_mai_n391_), .B0(mai_mai_n216_), .Y(mai_mai_n945_));
  OAI210     m0917(.A0(mai_mai_n945_), .A1(mai_mai_n944_), .B0(mai_mai_n405_), .Y(mai_mai_n946_));
  NO2        m0918(.A(mai_mai_n648_), .B(mai_mai_n267_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n601_), .B(mai_mai_n849_), .Y(mai_mai_n948_));
  AOI220     m0920(.A0(mai_mai_n948_), .A1(mai_mai_n576_), .B0(mai_mai_n826_), .B1(mai_mai_n947_), .Y(mai_mai_n949_));
  NO2        m0921(.A(mai_mai_n151_), .B(mai_mai_n239_), .Y(mai_mai_n950_));
  NA2        m0922(.A(mai_mai_n949_), .B(mai_mai_n946_), .Y(mai_mai_n951_));
  OR2        m0923(.A(mai_mai_n321_), .B(mai_mai_n938_), .Y(mai_mai_n952_));
  NA2        m0924(.A(mai_mai_n952_), .B(mai_mai_n354_), .Y(mai_mai_n953_));
  NO3        m0925(.A(mai_mai_n133_), .B(mai_mai_n152_), .C(mai_mai_n216_), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n954_), .B(mai_mai_n541_), .Y(mai_mai_n955_));
  NA4        m0927(.A(mai_mai_n446_), .B(mai_mai_n438_), .C(mai_mai_n181_), .D(g), .Y(mai_mai_n956_));
  NA3        m0928(.A(mai_mai_n956_), .B(mai_mai_n955_), .C(mai_mai_n953_), .Y(mai_mai_n957_));
  NO3        m0929(.A(mai_mai_n671_), .B(mai_mai_n90_), .C(mai_mai_n45_), .Y(mai_mai_n958_));
  NO4        m0930(.A(mai_mai_n958_), .B(mai_mai_n957_), .C(mai_mai_n951_), .D(mai_mai_n942_), .Y(mai_mai_n959_));
  NO2        m0931(.A(mai_mai_n370_), .B(mai_mai_n369_), .Y(mai_mai_n960_));
  NA2        m0932(.A(mai_mai_n598_), .B(mai_mai_n70_), .Y(mai_mai_n961_));
  NA2        m0933(.A(mai_mai_n566_), .B(mai_mai_n145_), .Y(mai_mai_n962_));
  NOi21      m0934(.An(mai_mai_n34_), .B(mai_mai_n662_), .Y(mai_mai_n963_));
  AOI220     m0935(.A0(mai_mai_n963_), .A1(mai_mai_n962_), .B0(mai_mai_n961_), .B1(mai_mai_n960_), .Y(mai_mai_n964_));
  OAI210     m0936(.A0(mai_mai_n254_), .A1(mai_mai_n45_), .B0(mai_mai_n964_), .Y(mai_mai_n965_));
  NA2        m0937(.A(mai_mai_n436_), .B(mai_mai_n269_), .Y(mai_mai_n966_));
  NO3        m0938(.A(mai_mai_n828_), .B(mai_mai_n88_), .C(mai_mai_n410_), .Y(mai_mai_n967_));
  NAi31      m0939(.An(mai_mai_n967_), .B(mai_mai_n966_), .C(mai_mai_n317_), .Y(mai_mai_n968_));
  NO2        m0940(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n969_));
  NO2        m0941(.A(mai_mai_n514_), .B(mai_mai_n296_), .Y(mai_mai_n970_));
  INV        m0942(.A(mai_mai_n970_), .Y(mai_mai_n971_));
  NO2        m0943(.A(mai_mai_n971_), .B(mai_mai_n145_), .Y(mai_mai_n972_));
  NA2        m0944(.A(mai_mai_n642_), .B(mai_mai_n363_), .Y(mai_mai_n973_));
  OAI210     m0945(.A0(mai_mai_n740_), .A1(mai_mai_n973_), .B0(mai_mai_n367_), .Y(mai_mai_n974_));
  NO4        m0946(.A(mai_mai_n974_), .B(mai_mai_n972_), .C(mai_mai_n968_), .D(mai_mai_n965_), .Y(mai_mai_n975_));
  NA2        m0947(.A(mai_mai_n346_), .B(g), .Y(mai_mai_n976_));
  NA2        m0948(.A(mai_mai_n162_), .B(i), .Y(mai_mai_n977_));
  NA2        m0949(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n978_));
  OAI220     m0950(.A0(mai_mai_n978_), .A1(mai_mai_n201_), .B0(mai_mai_n977_), .B1(mai_mai_n90_), .Y(mai_mai_n979_));
  INV        m0951(.A(mai_mai_n979_), .Y(mai_mai_n980_));
  NO2        m0952(.A(mai_mai_n145_), .B(mai_mai_n83_), .Y(mai_mai_n981_));
  OR2        m0953(.A(mai_mai_n981_), .B(mai_mai_n565_), .Y(mai_mai_n982_));
  NA2        m0954(.A(mai_mai_n566_), .B(mai_mai_n383_), .Y(mai_mai_n983_));
  AOI210     m0955(.A0(mai_mai_n983_), .A1(n), .B0(mai_mai_n982_), .Y(mai_mai_n984_));
  OAI220     m0956(.A0(mai_mai_n984_), .A1(mai_mai_n976_), .B0(mai_mai_n980_), .B1(mai_mai_n330_), .Y(mai_mai_n985_));
  NO2        m0957(.A(mai_mai_n668_), .B(mai_mai_n507_), .Y(mai_mai_n986_));
  NA3        m0958(.A(mai_mai_n341_), .B(mai_mai_n637_), .C(i), .Y(mai_mai_n987_));
  OAI210     m0959(.A0(mai_mai_n440_), .A1(mai_mai_n307_), .B0(mai_mai_n987_), .Y(mai_mai_n988_));
  OAI210     m0960(.A0(mai_mai_n988_), .A1(mai_mai_n986_), .B0(mai_mai_n682_), .Y(mai_mai_n989_));
  NA2        m0961(.A(mai_mai_n615_), .B(mai_mai_n113_), .Y(mai_mai_n990_));
  OR3        m0962(.A(mai_mai_n307_), .B(mai_mai_n435_), .C(f), .Y(mai_mai_n991_));
  OR2        m0963(.A(mai_mai_n991_), .B(mai_mai_n600_), .Y(mai_mai_n992_));
  NA3        m0964(.A(mai_mai_n322_), .B(mai_mai_n118_), .C(g), .Y(mai_mai_n993_));
  AOI210     m0965(.A0(mai_mai_n679_), .A1(mai_mai_n993_), .B0(m), .Y(mai_mai_n994_));
  OAI210     m0966(.A0(mai_mai_n994_), .A1(mai_mai_n939_), .B0(mai_mai_n321_), .Y(mai_mai_n995_));
  NA2        m0967(.A(mai_mai_n698_), .B(mai_mai_n885_), .Y(mai_mai_n996_));
  NA2        m0968(.A(mai_mai_n851_), .B(mai_mai_n441_), .Y(mai_mai_n997_));
  NA2        m0969(.A(mai_mai_n224_), .B(mai_mai_n76_), .Y(mai_mai_n998_));
  NA2        m0970(.A(mai_mai_n998_), .B(mai_mai_n991_), .Y(mai_mai_n999_));
  AOI220     m0971(.A0(mai_mai_n999_), .A1(mai_mai_n262_), .B0(mai_mai_n997_), .B1(mai_mai_n996_), .Y(mai_mai_n1000_));
  NA4        m0972(.A(mai_mai_n1000_), .B(mai_mai_n995_), .C(mai_mai_n992_), .D(mai_mai_n989_), .Y(mai_mai_n1001_));
  NO2        m0973(.A(mai_mai_n379_), .B(mai_mai_n89_), .Y(mai_mai_n1002_));
  NA2        m0974(.A(mai_mai_n1002_), .B(mai_mai_n240_), .Y(mai_mai_n1003_));
  NA2        m0975(.A(mai_mai_n670_), .B(mai_mai_n87_), .Y(mai_mai_n1004_));
  NO2        m0976(.A(mai_mai_n464_), .B(mai_mai_n216_), .Y(mai_mai_n1005_));
  AOI220     m0977(.A0(mai_mai_n1005_), .A1(mai_mai_n384_), .B0(mai_mai_n952_), .B1(mai_mai_n220_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n940_), .B(mai_mai_n950_), .Y(mai_mai_n1007_));
  NA4        m0979(.A(mai_mai_n1007_), .B(mai_mai_n1006_), .C(mai_mai_n1004_), .D(mai_mai_n1003_), .Y(mai_mai_n1008_));
  OAI210     m0980(.A0(mai_mai_n997_), .A1(mai_mai_n948_), .B0(mai_mai_n554_), .Y(mai_mai_n1009_));
  OAI210     m0981(.A0(mai_mai_n370_), .A1(mai_mai_n369_), .B0(mai_mai_n109_), .Y(mai_mai_n1010_));
  NA2        m0982(.A(mai_mai_n1010_), .B(mai_mai_n546_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(mai_mai_n994_), .B(mai_mai_n938_), .Y(mai_mai_n1012_));
  NO3        m0984(.A(mai_mai_n899_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n1013_));
  AOI220     m0985(.A0(mai_mai_n1013_), .A1(mai_mai_n635_), .B0(mai_mai_n653_), .B1(mai_mai_n541_), .Y(mai_mai_n1014_));
  NA4        m0986(.A(mai_mai_n1014_), .B(mai_mai_n1012_), .C(mai_mai_n1011_), .D(mai_mai_n1009_), .Y(mai_mai_n1015_));
  NO4        m0987(.A(mai_mai_n1015_), .B(mai_mai_n1008_), .C(mai_mai_n1001_), .D(mai_mai_n985_), .Y(mai_mai_n1016_));
  NAi31      m0988(.An(mai_mai_n142_), .B(mai_mai_n423_), .C(n), .Y(mai_mai_n1017_));
  NO3        m0989(.A(mai_mai_n126_), .B(mai_mai_n339_), .C(mai_mai_n857_), .Y(mai_mai_n1018_));
  NO2        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1017_), .Y(mai_mai_n1019_));
  NO3        m0991(.A(mai_mai_n276_), .B(mai_mai_n142_), .C(mai_mai_n410_), .Y(mai_mai_n1020_));
  AOI210     m0992(.A0(mai_mai_n1020_), .A1(mai_mai_n508_), .B0(mai_mai_n1019_), .Y(mai_mai_n1021_));
  NA2        m0993(.A(mai_mai_n500_), .B(i), .Y(mai_mai_n1022_));
  NA2        m0994(.A(mai_mai_n1022_), .B(mai_mai_n1021_), .Y(mai_mai_n1023_));
  NA2        m0995(.A(mai_mai_n233_), .B(mai_mai_n171_), .Y(mai_mai_n1024_));
  NO3        m0996(.A(mai_mai_n305_), .B(mai_mai_n446_), .C(mai_mai_n175_), .Y(mai_mai_n1025_));
  NOi31      m0997(.An(mai_mai_n1024_), .B(mai_mai_n1025_), .C(mai_mai_n216_), .Y(mai_mai_n1026_));
  NAi21      m0998(.An(mai_mai_n566_), .B(mai_mai_n1005_), .Y(mai_mai_n1027_));
  NA2        m0999(.A(mai_mai_n439_), .B(mai_mai_n885_), .Y(mai_mai_n1028_));
  NO3        m1000(.A(mai_mai_n440_), .B(mai_mai_n307_), .C(mai_mai_n72_), .Y(mai_mai_n1029_));
  AOI220     m1001(.A0(mai_mai_n1029_), .A1(mai_mai_n1028_), .B0(mai_mai_n489_), .B1(g), .Y(mai_mai_n1030_));
  NA2        m1002(.A(mai_mai_n1030_), .B(mai_mai_n1027_), .Y(mai_mai_n1031_));
  NO2        m1003(.A(mai_mai_n1017_), .B(mai_mai_n236_), .Y(mai_mai_n1032_));
  NA2        m1004(.A(mai_mai_n943_), .B(mai_mai_n934_), .Y(mai_mai_n1033_));
  NO3        m1005(.A(mai_mai_n555_), .B(mai_mai_n149_), .C(mai_mai_n215_), .Y(mai_mai_n1034_));
  OAI210     m1006(.A0(mai_mai_n1034_), .A1(mai_mai_n535_), .B0(mai_mai_n380_), .Y(mai_mai_n1035_));
  OAI220     m1007(.A0(mai_mai_n940_), .A1(mai_mai_n948_), .B0(mai_mai_n556_), .B1(mai_mai_n429_), .Y(mai_mai_n1036_));
  NA4        m1008(.A(mai_mai_n1036_), .B(mai_mai_n1035_), .C(mai_mai_n1033_), .D(mai_mai_n629_), .Y(mai_mai_n1037_));
  OAI210     m1009(.A0(mai_mai_n943_), .A1(mai_mai_n935_), .B0(mai_mai_n1024_), .Y(mai_mai_n1038_));
  NA3        m1010(.A(mai_mai_n983_), .B(mai_mai_n494_), .C(mai_mai_n46_), .Y(mai_mai_n1039_));
  INV        m1011(.A(mai_mai_n329_), .Y(mai_mai_n1040_));
  NA3        m1012(.A(mai_mai_n1040_), .B(mai_mai_n1039_), .C(mai_mai_n1038_), .Y(mai_mai_n1041_));
  OR3        m1013(.A(mai_mai_n1041_), .B(mai_mai_n1037_), .C(mai_mai_n1032_), .Y(mai_mai_n1042_));
  NO4        m1014(.A(mai_mai_n1042_), .B(mai_mai_n1031_), .C(mai_mai_n1026_), .D(mai_mai_n1023_), .Y(mai_mai_n1043_));
  NA4        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1016_), .C(mai_mai_n975_), .D(mai_mai_n959_), .Y(mai13));
  INV        m1016(.A(mai_mai_n46_), .Y(mai_mai_n1045_));
  AN2        m1017(.A(c), .B(b), .Y(mai_mai_n1046_));
  NA3        m1018(.A(mai_mai_n253_), .B(mai_mai_n1046_), .C(m), .Y(mai_mai_n1047_));
  NA2        m1019(.A(mai_mai_n505_), .B(f), .Y(mai_mai_n1048_));
  NO4        m1020(.A(mai_mai_n1048_), .B(mai_mai_n1047_), .C(mai_mai_n1045_), .D(mai_mai_n594_), .Y(mai_mai_n1049_));
  NA2        m1021(.A(mai_mai_n269_), .B(mai_mai_n1046_), .Y(mai_mai_n1050_));
  NO4        m1022(.A(mai_mai_n1050_), .B(mai_mai_n1048_), .C(mai_mai_n977_), .D(a), .Y(mai_mai_n1051_));
  NAi32      m1023(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1052_));
  NA2        m1024(.A(mai_mai_n141_), .B(mai_mai_n45_), .Y(mai_mai_n1053_));
  NO4        m1025(.A(mai_mai_n1053_), .B(mai_mai_n1052_), .C(mai_mai_n601_), .D(mai_mai_n304_), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n674_), .B(mai_mai_n227_), .Y(mai_mai_n1055_));
  NA2        m1027(.A(mai_mai_n413_), .B(mai_mai_n215_), .Y(mai_mai_n1056_));
  AN2        m1028(.A(d), .B(c), .Y(mai_mai_n1057_));
  NA2        m1029(.A(mai_mai_n1057_), .B(mai_mai_n116_), .Y(mai_mai_n1058_));
  NO4        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1056_), .C(mai_mai_n176_), .D(mai_mai_n167_), .Y(mai_mai_n1059_));
  NA2        m1031(.A(mai_mai_n505_), .B(c), .Y(mai_mai_n1060_));
  NO4        m1032(.A(mai_mai_n1053_), .B(mai_mai_n597_), .C(mai_mai_n1060_), .D(mai_mai_n304_), .Y(mai_mai_n1061_));
  AO210      m1033(.A0(mai_mai_n1059_), .A1(mai_mai_n1055_), .B0(mai_mai_n1061_), .Y(mai_mai_n1062_));
  OR4        m1034(.A(mai_mai_n1062_), .B(mai_mai_n1054_), .C(mai_mai_n1051_), .D(mai_mai_n1049_), .Y(mai_mai_n1063_));
  NAi32      m1035(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1064_));
  NO2        m1036(.A(mai_mai_n1064_), .B(mai_mai_n146_), .Y(mai_mai_n1065_));
  NA2        m1037(.A(mai_mai_n1065_), .B(g), .Y(mai_mai_n1066_));
  OR3        m1038(.A(mai_mai_n227_), .B(mai_mai_n176_), .C(mai_mai_n167_), .Y(mai_mai_n1067_));
  NO2        m1039(.A(mai_mai_n1067_), .B(mai_mai_n1066_), .Y(mai_mai_n1068_));
  NO2        m1040(.A(mai_mai_n1060_), .B(mai_mai_n304_), .Y(mai_mai_n1069_));
  NO2        m1041(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1070_));
  NA2        m1042(.A(mai_mai_n639_), .B(mai_mai_n1070_), .Y(mai_mai_n1071_));
  NOi21      m1043(.An(mai_mai_n1069_), .B(mai_mai_n1071_), .Y(mai_mai_n1072_));
  NO2        m1044(.A(mai_mai_n769_), .B(mai_mai_n112_), .Y(mai_mai_n1073_));
  NOi41      m1045(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1074_));
  NA2        m1046(.A(mai_mai_n1074_), .B(mai_mai_n1073_), .Y(mai_mai_n1075_));
  NO2        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1066_), .Y(mai_mai_n1076_));
  OR3        m1048(.A(e), .B(d), .C(c), .Y(mai_mai_n1077_));
  NA3        m1049(.A(k), .B(j), .C(i), .Y(mai_mai_n1078_));
  NO3        m1050(.A(mai_mai_n1078_), .B(mai_mai_n304_), .C(mai_mai_n89_), .Y(mai_mai_n1079_));
  NOi21      m1051(.An(mai_mai_n1079_), .B(mai_mai_n1077_), .Y(mai_mai_n1080_));
  OR4        m1052(.A(mai_mai_n1080_), .B(mai_mai_n1076_), .C(mai_mai_n1072_), .D(mai_mai_n1068_), .Y(mai_mai_n1081_));
  NA3        m1053(.A(mai_mai_n472_), .B(mai_mai_n332_), .C(mai_mai_n56_), .Y(mai_mai_n1082_));
  NO2        m1054(.A(mai_mai_n1082_), .B(mai_mai_n1071_), .Y(mai_mai_n1083_));
  NO4        m1055(.A(mai_mai_n1082_), .B(mai_mai_n597_), .C(mai_mai_n453_), .D(mai_mai_n45_), .Y(mai_mai_n1084_));
  NO2        m1056(.A(f), .B(c), .Y(mai_mai_n1085_));
  NOi21      m1057(.An(mai_mai_n1085_), .B(mai_mai_n445_), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n59_), .Y(mai_mai_n1087_));
  OR2        m1059(.A(k), .B(i), .Y(mai_mai_n1088_));
  NO3        m1060(.A(mai_mai_n1088_), .B(mai_mai_n246_), .C(l), .Y(mai_mai_n1089_));
  NOi31      m1061(.An(mai_mai_n1089_), .B(mai_mai_n1087_), .C(j), .Y(mai_mai_n1090_));
  OR3        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1084_), .C(mai_mai_n1083_), .Y(mai_mai_n1091_));
  OR3        m1063(.A(mai_mai_n1091_), .B(mai_mai_n1081_), .C(mai_mai_n1063_), .Y(mai02));
  OR2        m1064(.A(l), .B(k), .Y(mai_mai_n1093_));
  OR3        m1065(.A(h), .B(g), .C(f), .Y(mai_mai_n1094_));
  OR3        m1066(.A(n), .B(m), .C(i), .Y(mai_mai_n1095_));
  NO4        m1067(.A(mai_mai_n1095_), .B(mai_mai_n1094_), .C(mai_mai_n1093_), .D(mai_mai_n1077_), .Y(mai_mai_n1096_));
  INV        m1068(.A(mai_mai_n1054_), .Y(mai_mai_n1097_));
  AN3        m1069(.A(g), .B(f), .C(c), .Y(mai_mai_n1098_));
  NA3        m1070(.A(mai_mai_n1098_), .B(mai_mai_n472_), .C(h), .Y(mai_mai_n1099_));
  OR2        m1071(.A(mai_mai_n1078_), .B(mai_mai_n304_), .Y(mai_mai_n1100_));
  OR2        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1099_), .Y(mai_mai_n1101_));
  NO3        m1073(.A(mai_mai_n1082_), .B(mai_mai_n1053_), .C(mai_mai_n597_), .Y(mai_mai_n1102_));
  NO2        m1074(.A(mai_mai_n1102_), .B(mai_mai_n1068_), .Y(mai_mai_n1103_));
  NA3        m1075(.A(l), .B(k), .C(j), .Y(mai_mai_n1104_));
  NA2        m1076(.A(i), .B(h), .Y(mai_mai_n1105_));
  NO3        m1077(.A(mai_mai_n1105_), .B(mai_mai_n1104_), .C(mai_mai_n133_), .Y(mai_mai_n1106_));
  NO3        m1078(.A(mai_mai_n143_), .B(mai_mai_n287_), .C(mai_mai_n216_), .Y(mai_mai_n1107_));
  AOI210     m1079(.A0(mai_mai_n1107_), .A1(mai_mai_n1106_), .B0(mai_mai_n1072_), .Y(mai_mai_n1108_));
  NA3        m1080(.A(c), .B(b), .C(a), .Y(mai_mai_n1109_));
  NO3        m1081(.A(mai_mai_n1109_), .B(mai_mai_n907_), .C(mai_mai_n215_), .Y(mai_mai_n1110_));
  NO4        m1082(.A(mai_mai_n1078_), .B(mai_mai_n296_), .C(mai_mai_n49_), .D(mai_mai_n112_), .Y(mai_mai_n1111_));
  AOI210     m1083(.A0(mai_mai_n1111_), .A1(mai_mai_n1110_), .B0(mai_mai_n1083_), .Y(mai_mai_n1112_));
  AN4        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1108_), .C(mai_mai_n1103_), .D(mai_mai_n1101_), .Y(mai_mai_n1113_));
  NO2        m1085(.A(mai_mai_n1058_), .B(mai_mai_n1056_), .Y(mai_mai_n1114_));
  NA2        m1086(.A(mai_mai_n1075_), .B(mai_mai_n1067_), .Y(mai_mai_n1115_));
  AOI210     m1087(.A0(mai_mai_n1115_), .A1(mai_mai_n1114_), .B0(mai_mai_n1049_), .Y(mai_mai_n1116_));
  NAi41      m1088(.An(mai_mai_n1096_), .B(mai_mai_n1116_), .C(mai_mai_n1113_), .D(mai_mai_n1097_), .Y(mai03));
  NO2        m1089(.A(mai_mai_n537_), .B(mai_mai_n606_), .Y(mai_mai_n1118_));
  NA4        m1090(.A(mai_mai_n586_), .B(m), .C(mai_mai_n112_), .D(mai_mai_n215_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n1119_), .B(mai_mai_n371_), .Y(mai_mai_n1120_));
  NO3        m1092(.A(mai_mai_n1120_), .B(mai_mai_n1118_), .C(mai_mai_n1010_), .Y(mai_mai_n1121_));
  NOi41      m1093(.An(mai_mai_n813_), .B(mai_mai_n862_), .C(mai_mai_n852_), .D(mai_mai_n724_), .Y(mai_mai_n1122_));
  OAI220     m1094(.A0(mai_mai_n1122_), .A1(mai_mai_n698_), .B0(mai_mai_n1121_), .B1(mai_mai_n598_), .Y(mai_mai_n1123_));
  NOi31      m1095(.An(m), .B(n), .C(f), .Y(mai_mai_n1124_));
  NA2        m1096(.A(mai_mai_n1124_), .B(mai_mai_n51_), .Y(mai_mai_n1125_));
  AN2        m1097(.A(e), .B(c), .Y(mai_mai_n1126_));
  NO2        m1098(.A(mai_mai_n892_), .B(mai_mai_n428_), .Y(mai_mai_n1127_));
  NA2        m1099(.A(mai_mai_n517_), .B(l), .Y(mai_mai_n1128_));
  NOi31      m1100(.An(mai_mai_n871_), .B(mai_mai_n1047_), .C(mai_mai_n1128_), .Y(mai_mai_n1129_));
  NO2        m1101(.A(mai_mai_n1129_), .B(mai_mai_n1127_), .Y(mai_mai_n1130_));
  NO2        m1102(.A(mai_mai_n287_), .B(a), .Y(mai_mai_n1131_));
  INV        m1103(.A(mai_mai_n1054_), .Y(mai_mai_n1132_));
  NO2        m1104(.A(mai_mai_n1105_), .B(mai_mai_n492_), .Y(mai_mai_n1133_));
  NO2        m1105(.A(mai_mai_n86_), .B(g), .Y(mai_mai_n1134_));
  AOI210     m1106(.A0(mai_mai_n1134_), .A1(mai_mai_n1133_), .B0(mai_mai_n1089_), .Y(mai_mai_n1135_));
  OR2        m1107(.A(mai_mai_n1135_), .B(mai_mai_n1087_), .Y(mai_mai_n1136_));
  NA3        m1108(.A(mai_mai_n1136_), .B(mai_mai_n1132_), .C(mai_mai_n1130_), .Y(mai_mai_n1137_));
  NO4        m1109(.A(mai_mai_n1137_), .B(mai_mai_n1123_), .C(mai_mai_n829_), .D(mai_mai_n575_), .Y(mai_mai_n1138_));
  NA2        m1110(.A(c), .B(b), .Y(mai_mai_n1139_));
  NO2        m1111(.A(mai_mai_n710_), .B(mai_mai_n1139_), .Y(mai_mai_n1140_));
  OAI210     m1112(.A0(mai_mai_n869_), .A1(mai_mai_n844_), .B0(mai_mai_n417_), .Y(mai_mai_n1141_));
  OAI210     m1113(.A0(mai_mai_n1141_), .A1(mai_mai_n870_), .B0(mai_mai_n1140_), .Y(mai_mai_n1142_));
  NAi21      m1114(.An(mai_mai_n425_), .B(mai_mai_n1140_), .Y(mai_mai_n1143_));
  NA3        m1115(.A(mai_mai_n429_), .B(mai_mai_n571_), .C(f), .Y(mai_mai_n1144_));
  NA2        m1116(.A(mai_mai_n560_), .B(mai_mai_n1131_), .Y(mai_mai_n1145_));
  NA3        m1117(.A(mai_mai_n1145_), .B(mai_mai_n1144_), .C(mai_mai_n1143_), .Y(mai_mai_n1146_));
  NAi21      m1118(.An(f), .B(d), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n1147_), .B(mai_mai_n1109_), .Y(mai_mai_n1148_));
  INV        m1120(.A(mai_mai_n1146_), .Y(mai_mai_n1149_));
  NO2        m1121(.A(mai_mai_n182_), .B(mai_mai_n239_), .Y(mai_mai_n1150_));
  NA2        m1122(.A(mai_mai_n1150_), .B(m), .Y(mai_mai_n1151_));
  NA3        m1123(.A(mai_mai_n924_), .B(mai_mai_n1128_), .C(mai_mai_n478_), .Y(mai_mai_n1152_));
  NA2        m1124(.A(mai_mai_n1152_), .B(mai_mai_n476_), .Y(mai_mai_n1153_));
  NO2        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1151_), .Y(mai_mai_n1154_));
  NA2        m1126(.A(mai_mai_n158_), .B(mai_mai_n33_), .Y(mai_mai_n1155_));
  AOI210     m1127(.A0(mai_mai_n973_), .A1(mai_mai_n1155_), .B0(mai_mai_n216_), .Y(mai_mai_n1156_));
  OAI210     m1128(.A0(mai_mai_n1156_), .A1(mai_mai_n449_), .B0(mai_mai_n1148_), .Y(mai_mai_n1157_));
  NO2        m1129(.A(mai_mai_n374_), .B(mai_mai_n373_), .Y(mai_mai_n1158_));
  INV        m1130(.A(mai_mai_n967_), .Y(mai_mai_n1159_));
  NAi31      m1131(.An(mai_mai_n1158_), .B(mai_mai_n1159_), .C(mai_mai_n1157_), .Y(mai_mai_n1160_));
  NO2        m1132(.A(mai_mai_n1160_), .B(mai_mai_n1154_), .Y(mai_mai_n1161_));
  NA4        m1133(.A(mai_mai_n1161_), .B(mai_mai_n1149_), .C(mai_mai_n1142_), .D(mai_mai_n1138_), .Y(mai00));
  AOI210     m1134(.A0(mai_mai_n295_), .A1(mai_mai_n216_), .B0(mai_mai_n279_), .Y(mai_mai_n1163_));
  NO2        m1135(.A(mai_mai_n1163_), .B(mai_mai_n589_), .Y(mai_mai_n1164_));
  NA2        m1136(.A(mai_mai_n905_), .B(mai_mai_n950_), .Y(mai_mai_n1165_));
  NO3        m1137(.A(mai_mai_n1102_), .B(mai_mai_n967_), .C(mai_mai_n721_), .Y(mai_mai_n1166_));
  NA3        m1138(.A(mai_mai_n1166_), .B(mai_mai_n1165_), .C(mai_mai_n1011_), .Y(mai_mai_n1167_));
  NA2        m1139(.A(mai_mai_n519_), .B(f), .Y(mai_mai_n1168_));
  OAI210     m1140(.A0(mai_mai_n1018_), .A1(mai_mai_n40_), .B0(mai_mai_n655_), .Y(mai_mai_n1169_));
  NA3        m1141(.A(mai_mai_n1169_), .B(mai_mai_n261_), .C(n), .Y(mai_mai_n1170_));
  AOI210     m1142(.A0(mai_mai_n1170_), .A1(mai_mai_n1168_), .B0(mai_mai_n1058_), .Y(mai_mai_n1171_));
  NO4        m1143(.A(mai_mai_n1171_), .B(mai_mai_n1167_), .C(mai_mai_n1164_), .D(mai_mai_n1081_), .Y(mai_mai_n1172_));
  NA3        m1144(.A(mai_mai_n166_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1173_));
  NA3        m1145(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1174_));
  NOi31      m1146(.An(n), .B(m), .C(i), .Y(mai_mai_n1175_));
  NA3        m1147(.A(mai_mai_n1175_), .B(mai_mai_n658_), .C(mai_mai_n51_), .Y(mai_mai_n1176_));
  OAI210     m1148(.A0(mai_mai_n1174_), .A1(mai_mai_n1173_), .B0(mai_mai_n1176_), .Y(mai_mai_n1177_));
  INV        m1149(.A(mai_mai_n588_), .Y(mai_mai_n1178_));
  NO2        m1150(.A(mai_mai_n1178_), .B(mai_mai_n1177_), .Y(mai_mai_n1179_));
  NO4        m1151(.A(mai_mai_n495_), .B(mai_mai_n356_), .C(mai_mai_n1139_), .D(mai_mai_n59_), .Y(mai_mai_n1180_));
  NA3        m1152(.A(mai_mai_n385_), .B(mai_mai_n223_), .C(g), .Y(mai_mai_n1181_));
  OA220      m1153(.A0(mai_mai_n1181_), .A1(mai_mai_n1174_), .B0(mai_mai_n386_), .B1(mai_mai_n136_), .Y(mai_mai_n1182_));
  NO2        m1154(.A(h), .B(g), .Y(mai_mai_n1183_));
  NA4        m1155(.A(mai_mai_n508_), .B(mai_mai_n472_), .C(mai_mai_n1183_), .D(mai_mai_n1046_), .Y(mai_mai_n1184_));
  OAI220     m1156(.A0(mai_mai_n537_), .A1(mai_mai_n606_), .B0(mai_mai_n90_), .B1(mai_mai_n89_), .Y(mai_mai_n1185_));
  AOI220     m1157(.A0(mai_mai_n1185_), .A1(mai_mai_n546_), .B0(mai_mai_n954_), .B1(mai_mai_n587_), .Y(mai_mai_n1186_));
  AOI220     m1158(.A0(mai_mai_n314_), .A1(mai_mai_n250_), .B0(mai_mai_n177_), .B1(mai_mai_n148_), .Y(mai_mai_n1187_));
  NA4        m1159(.A(mai_mai_n1187_), .B(mai_mai_n1186_), .C(mai_mai_n1184_), .D(mai_mai_n1182_), .Y(mai_mai_n1188_));
  NO3        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1180_), .C(mai_mai_n271_), .Y(mai_mai_n1189_));
  INV        m1161(.A(mai_mai_n319_), .Y(mai_mai_n1190_));
  NA2        m1162(.A(mai_mai_n250_), .B(mai_mai_n346_), .Y(mai_mai_n1191_));
  NA2        m1163(.A(mai_mai_n1191_), .B(mai_mai_n1190_), .Y(mai_mai_n1192_));
  NA3        m1164(.A(mai_mai_n179_), .B(mai_mai_n112_), .C(g), .Y(mai_mai_n1193_));
  NA3        m1165(.A(mai_mai_n472_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1194_));
  NOi31      m1166(.An(mai_mai_n878_), .B(mai_mai_n1194_), .C(mai_mai_n1193_), .Y(mai_mai_n1195_));
  NO2        m1167(.A(mai_mai_n278_), .B(mai_mai_n72_), .Y(mai_mai_n1196_));
  NO3        m1168(.A(mai_mai_n428_), .B(mai_mai_n840_), .C(n), .Y(mai_mai_n1197_));
  AOI210     m1169(.A0(mai_mai_n1197_), .A1(mai_mai_n1196_), .B0(mai_mai_n1096_), .Y(mai_mai_n1198_));
  NAi31      m1170(.An(mai_mai_n1061_), .B(mai_mai_n1198_), .C(mai_mai_n71_), .Y(mai_mai_n1199_));
  NO3        m1171(.A(mai_mai_n1199_), .B(mai_mai_n1195_), .C(mai_mai_n1192_), .Y(mai_mai_n1200_));
  AN3        m1172(.A(mai_mai_n1200_), .B(mai_mai_n1189_), .C(mai_mai_n1179_), .Y(mai_mai_n1201_));
  NA2        m1173(.A(mai_mai_n546_), .B(mai_mai_n100_), .Y(mai_mai_n1202_));
  NA3        m1174(.A(mai_mai_n1124_), .B(mai_mai_n615_), .C(mai_mai_n471_), .Y(mai_mai_n1203_));
  NA3        m1175(.A(mai_mai_n1203_), .B(mai_mai_n1202_), .C(mai_mai_n244_), .Y(mai_mai_n1204_));
  NA2        m1176(.A(mai_mai_n1120_), .B(mai_mai_n546_), .Y(mai_mai_n1205_));
  INV        m1177(.A(mai_mai_n1205_), .Y(mai_mai_n1206_));
  OAI210     m1178(.A0(mai_mai_n470_), .A1(mai_mai_n120_), .B0(mai_mai_n872_), .Y(mai_mai_n1207_));
  NA2        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1152_), .Y(mai_mai_n1208_));
  OR4        m1180(.A(mai_mai_n1058_), .B(mai_mai_n276_), .C(mai_mai_n225_), .D(e), .Y(mai_mai_n1209_));
  NO2        m1181(.A(mai_mai_n219_), .B(mai_mai_n216_), .Y(mai_mai_n1210_));
  NA2        m1182(.A(n), .B(e), .Y(mai_mai_n1211_));
  NO2        m1183(.A(mai_mai_n1211_), .B(mai_mai_n146_), .Y(mai_mai_n1212_));
  AOI220     m1184(.A0(mai_mai_n1212_), .A1(mai_mai_n277_), .B0(mai_mai_n855_), .B1(mai_mai_n1210_), .Y(mai_mai_n1213_));
  OAI210     m1185(.A0(mai_mai_n357_), .A1(mai_mai_n309_), .B0(mai_mai_n451_), .Y(mai_mai_n1214_));
  NA4        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1213_), .C(mai_mai_n1209_), .D(mai_mai_n1208_), .Y(mai_mai_n1215_));
  NA2        m1187(.A(mai_mai_n1212_), .B(mai_mai_n859_), .Y(mai_mai_n1216_));
  AOI220     m1188(.A0(mai_mai_n963_), .A1(mai_mai_n587_), .B0(mai_mai_n658_), .B1(mai_mai_n247_), .Y(mai_mai_n1217_));
  NO2        m1189(.A(mai_mai_n65_), .B(h), .Y(mai_mai_n1218_));
  NO3        m1190(.A(mai_mai_n1058_), .B(mai_mai_n1056_), .C(mai_mai_n733_), .Y(mai_mai_n1219_));
  NO2        m1191(.A(mai_mai_n1093_), .B(mai_mai_n133_), .Y(mai_mai_n1220_));
  AN2        m1192(.A(mai_mai_n1220_), .B(mai_mai_n1107_), .Y(mai_mai_n1221_));
  OAI210     m1193(.A0(mai_mai_n1221_), .A1(mai_mai_n1219_), .B0(mai_mai_n1218_), .Y(mai_mai_n1222_));
  NA4        m1194(.A(mai_mai_n1222_), .B(mai_mai_n1217_), .C(mai_mai_n1216_), .D(mai_mai_n873_), .Y(mai_mai_n1223_));
  NO4        m1195(.A(mai_mai_n1223_), .B(mai_mai_n1215_), .C(mai_mai_n1206_), .D(mai_mai_n1204_), .Y(mai_mai_n1224_));
  NA2        m1196(.A(mai_mai_n845_), .B(mai_mai_n764_), .Y(mai_mai_n1225_));
  NA4        m1197(.A(mai_mai_n1225_), .B(mai_mai_n1224_), .C(mai_mai_n1201_), .D(mai_mai_n1172_), .Y(mai01));
  AN2        m1198(.A(mai_mai_n1035_), .B(mai_mai_n1033_), .Y(mai_mai_n1227_));
  NO3        m1199(.A(mai_mai_n804_), .B(mai_mai_n486_), .C(mai_mai_n285_), .Y(mai_mai_n1228_));
  NA2        m1200(.A(mai_mai_n396_), .B(i), .Y(mai_mai_n1229_));
  NA3        m1201(.A(mai_mai_n1229_), .B(mai_mai_n1228_), .C(mai_mai_n1227_), .Y(mai_mai_n1230_));
  NA2        m1202(.A(mai_mai_n566_), .B(mai_mai_n275_), .Y(mai_mai_n1231_));
  NA2        m1203(.A(mai_mai_n970_), .B(mai_mai_n1231_), .Y(mai_mai_n1232_));
  NA3        m1204(.A(mai_mai_n1232_), .B(mai_mai_n920_), .C(mai_mai_n331_), .Y(mai_mai_n1233_));
  NA2        m1205(.A(mai_mai_n45_), .B(f), .Y(mai_mai_n1234_));
  NA2        m1206(.A(mai_mai_n717_), .B(mai_mai_n95_), .Y(mai_mai_n1235_));
  NO2        m1207(.A(mai_mai_n1235_), .B(mai_mai_n1234_), .Y(mai_mai_n1236_));
  NO2        m1208(.A(mai_mai_n790_), .B(mai_mai_n610_), .Y(mai_mai_n1237_));
  AOI210     m1209(.A0(mai_mai_n1236_), .A1(mai_mai_n643_), .B0(mai_mai_n1237_), .Y(mai_mai_n1238_));
  INV        m1210(.A(mai_mai_n118_), .Y(mai_mai_n1239_));
  OA220      m1211(.A0(mai_mai_n1239_), .A1(mai_mai_n596_), .B0(mai_mai_n669_), .B1(mai_mai_n371_), .Y(mai_mai_n1240_));
  NAi41      m1212(.An(mai_mai_n161_), .B(mai_mai_n1240_), .C(mai_mai_n1238_), .D(mai_mai_n904_), .Y(mai_mai_n1241_));
  NO3        m1213(.A(mai_mai_n791_), .B(mai_mai_n681_), .C(mai_mai_n522_), .Y(mai_mai_n1242_));
  NA4        m1214(.A(mai_mai_n717_), .B(mai_mai_n95_), .C(mai_mai_n45_), .D(mai_mai_n215_), .Y(mai_mai_n1243_));
  OA220      m1215(.A0(mai_mai_n1243_), .A1(mai_mai_n677_), .B0(mai_mai_n196_), .B1(mai_mai_n194_), .Y(mai_mai_n1244_));
  NA3        m1216(.A(mai_mai_n1244_), .B(mai_mai_n1242_), .C(mai_mai_n139_), .Y(mai_mai_n1245_));
  NO4        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1241_), .C(mai_mai_n1233_), .D(mai_mai_n1230_), .Y(mai_mai_n1246_));
  INV        m1218(.A(mai_mai_n1181_), .Y(mai_mai_n1247_));
  OAI210     m1219(.A0(mai_mai_n1247_), .A1(mai_mai_n298_), .B0(mai_mai_n541_), .Y(mai_mai_n1248_));
  NA2        m1220(.A(mai_mai_n549_), .B(mai_mai_n398_), .Y(mai_mai_n1249_));
  NOi21      m1221(.An(mai_mai_n572_), .B(mai_mai_n593_), .Y(mai_mai_n1250_));
  NA2        m1222(.A(mai_mai_n1250_), .B(mai_mai_n1249_), .Y(mai_mai_n1251_));
  AOI210     m1223(.A0(mai_mai_n205_), .A1(mai_mai_n88_), .B0(mai_mai_n215_), .Y(mai_mai_n1252_));
  OAI210     m1224(.A0(mai_mai_n816_), .A1(mai_mai_n429_), .B0(mai_mai_n1252_), .Y(mai_mai_n1253_));
  AN3        m1225(.A(m), .B(l), .C(k), .Y(mai_mai_n1254_));
  OAI210     m1226(.A0(mai_mai_n359_), .A1(mai_mai_n34_), .B0(mai_mai_n1254_), .Y(mai_mai_n1255_));
  NA2        m1227(.A(mai_mai_n204_), .B(mai_mai_n34_), .Y(mai_mai_n1256_));
  AO210      m1228(.A0(mai_mai_n1256_), .A1(mai_mai_n1255_), .B0(mai_mai_n330_), .Y(mai_mai_n1257_));
  NA4        m1229(.A(mai_mai_n1257_), .B(mai_mai_n1253_), .C(mai_mai_n1251_), .D(mai_mai_n1248_), .Y(mai_mai_n1258_));
  AOI210     m1230(.A0(mai_mai_n604_), .A1(mai_mai_n118_), .B0(mai_mai_n607_), .Y(mai_mai_n1259_));
  OAI210     m1231(.A0(mai_mai_n1239_), .A1(mai_mai_n603_), .B0(mai_mai_n1259_), .Y(mai_mai_n1260_));
  NA2        m1232(.A(mai_mai_n284_), .B(mai_mai_n196_), .Y(mai_mai_n1261_));
  NA2        m1233(.A(mai_mai_n1261_), .B(mai_mai_n673_), .Y(mai_mai_n1262_));
  INV        m1234(.A(mai_mai_n967_), .Y(mai_mai_n1263_));
  OAI210     m1235(.A0(mai_mai_n1236_), .A1(mai_mai_n324_), .B0(mai_mai_n682_), .Y(mai_mai_n1264_));
  NA4        m1236(.A(mai_mai_n1264_), .B(mai_mai_n1263_), .C(mai_mai_n1262_), .D(mai_mai_n794_), .Y(mai_mai_n1265_));
  NO3        m1237(.A(mai_mai_n1265_), .B(mai_mai_n1260_), .C(mai_mai_n1258_), .Y(mai_mai_n1266_));
  NA2        m1238(.A(mai_mai_n515_), .B(mai_mai_n58_), .Y(mai_mai_n1267_));
  OR3        m1239(.A(mai_mai_n1235_), .B(mai_mai_n612_), .C(mai_mai_n1234_), .Y(mai_mai_n1268_));
  NO2        m1240(.A(mai_mai_n1243_), .B(mai_mai_n990_), .Y(mai_mai_n1269_));
  NO2        m1241(.A(mai_mai_n208_), .B(mai_mai_n111_), .Y(mai_mai_n1270_));
  NO3        m1242(.A(mai_mai_n1270_), .B(mai_mai_n1269_), .C(mai_mai_n1177_), .Y(mai_mai_n1271_));
  NA4        m1243(.A(mai_mai_n1271_), .B(mai_mai_n1268_), .C(mai_mai_n1267_), .D(mai_mai_n763_), .Y(mai_mai_n1272_));
  NO2        m1244(.A(mai_mai_n977_), .B(mai_mai_n235_), .Y(mai_mai_n1273_));
  NO2        m1245(.A(mai_mai_n978_), .B(mai_mai_n568_), .Y(mai_mai_n1274_));
  OAI210     m1246(.A0(mai_mai_n1274_), .A1(mai_mai_n1273_), .B0(mai_mai_n339_), .Y(mai_mai_n1275_));
  NA2        m1247(.A(mai_mai_n582_), .B(mai_mai_n580_), .Y(mai_mai_n1276_));
  NO3        m1248(.A(mai_mai_n78_), .B(mai_mai_n296_), .C(mai_mai_n45_), .Y(mai_mai_n1277_));
  NA2        m1249(.A(mai_mai_n1277_), .B(mai_mai_n565_), .Y(mai_mai_n1278_));
  NA2        m1250(.A(mai_mai_n1278_), .B(mai_mai_n1276_), .Y(mai_mai_n1279_));
  OR2        m1251(.A(mai_mai_n1181_), .B(mai_mai_n1174_), .Y(mai_mai_n1280_));
  NA2        m1252(.A(mai_mai_n1277_), .B(mai_mai_n819_), .Y(mai_mai_n1281_));
  NA3        m1253(.A(mai_mai_n1281_), .B(mai_mai_n1280_), .C(mai_mai_n388_), .Y(mai_mai_n1282_));
  NOi41      m1254(.An(mai_mai_n1275_), .B(mai_mai_n1282_), .C(mai_mai_n1279_), .D(mai_mai_n1272_), .Y(mai_mai_n1283_));
  NO2        m1255(.A(mai_mai_n132_), .B(mai_mai_n45_), .Y(mai_mai_n1284_));
  NO2        m1256(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1285_));
  AO220      m1257(.A0(mai_mai_n1285_), .A1(mai_mai_n632_), .B0(mai_mai_n1284_), .B1(mai_mai_n715_), .Y(mai_mai_n1286_));
  NA2        m1258(.A(mai_mai_n1286_), .B(mai_mai_n339_), .Y(mai_mai_n1287_));
  INV        m1259(.A(mai_mai_n136_), .Y(mai_mai_n1288_));
  NO3        m1260(.A(mai_mai_n1105_), .B(mai_mai_n176_), .C(mai_mai_n86_), .Y(mai_mai_n1289_));
  AOI220     m1261(.A0(mai_mai_n1289_), .A1(mai_mai_n1288_), .B0(mai_mai_n1277_), .B1(mai_mai_n981_), .Y(mai_mai_n1290_));
  NA2        m1262(.A(mai_mai_n1290_), .B(mai_mai_n1287_), .Y(mai_mai_n1291_));
  NO2        m1263(.A(mai_mai_n623_), .B(mai_mai_n622_), .Y(mai_mai_n1292_));
  NO4        m1264(.A(mai_mai_n1105_), .B(mai_mai_n1292_), .C(mai_mai_n174_), .D(mai_mai_n86_), .Y(mai_mai_n1293_));
  NO3        m1265(.A(mai_mai_n1293_), .B(mai_mai_n1291_), .C(mai_mai_n647_), .Y(mai_mai_n1294_));
  NA4        m1266(.A(mai_mai_n1294_), .B(mai_mai_n1283_), .C(mai_mai_n1266_), .D(mai_mai_n1246_), .Y(mai06));
  NO2        m1267(.A(mai_mai_n227_), .B(mai_mai_n102_), .Y(mai_mai_n1296_));
  OAI210     m1268(.A0(mai_mai_n1296_), .A1(mai_mai_n1289_), .B0(mai_mai_n384_), .Y(mai_mai_n1297_));
  NO3        m1269(.A(mai_mai_n608_), .B(mai_mai_n814_), .C(mai_mai_n609_), .Y(mai_mai_n1298_));
  OR2        m1270(.A(mai_mai_n1298_), .B(mai_mai_n892_), .Y(mai_mai_n1299_));
  NA3        m1271(.A(mai_mai_n1299_), .B(mai_mai_n1297_), .C(mai_mai_n1275_), .Y(mai_mai_n1300_));
  NO3        m1272(.A(mai_mai_n1300_), .B(mai_mai_n1279_), .C(mai_mai_n260_), .Y(mai_mai_n1301_));
  NO2        m1273(.A(mai_mai_n296_), .B(mai_mai_n45_), .Y(mai_mai_n1302_));
  AOI210     m1274(.A0(mai_mai_n1302_), .A1(mai_mai_n982_), .B0(mai_mai_n1273_), .Y(mai_mai_n1303_));
  AOI210     m1275(.A0(mai_mai_n1302_), .A1(mai_mai_n569_), .B0(mai_mai_n1286_), .Y(mai_mai_n1304_));
  AOI210     m1276(.A0(mai_mai_n1304_), .A1(mai_mai_n1303_), .B0(mai_mai_n336_), .Y(mai_mai_n1305_));
  OAI210     m1277(.A0(mai_mai_n88_), .A1(mai_mai_n40_), .B0(mai_mai_n680_), .Y(mai_mai_n1306_));
  NA2        m1278(.A(mai_mai_n1306_), .B(mai_mai_n651_), .Y(mai_mai_n1307_));
  NO2        m1279(.A(mai_mai_n525_), .B(mai_mai_n171_), .Y(mai_mai_n1308_));
  NOi21      m1280(.An(mai_mai_n138_), .B(mai_mai_n45_), .Y(mai_mai_n1309_));
  NO2        m1281(.A(mai_mai_n616_), .B(mai_mai_n1125_), .Y(mai_mai_n1310_));
  OAI210     m1282(.A0(mai_mai_n465_), .A1(mai_mai_n251_), .B0(mai_mai_n914_), .Y(mai_mai_n1311_));
  NO4        m1283(.A(mai_mai_n1311_), .B(mai_mai_n1310_), .C(mai_mai_n1309_), .D(mai_mai_n1308_), .Y(mai_mai_n1312_));
  NO2        m1284(.A(mai_mai_n370_), .B(mai_mai_n137_), .Y(mai_mai_n1313_));
  AOI210     m1285(.A0(mai_mai_n1313_), .A1(mai_mai_n599_), .B0(mai_mai_n607_), .Y(mai_mai_n1314_));
  NA3        m1286(.A(mai_mai_n1314_), .B(mai_mai_n1312_), .C(mai_mai_n1307_), .Y(mai_mai_n1315_));
  NO2        m1287(.A(mai_mai_n755_), .B(mai_mai_n369_), .Y(mai_mai_n1316_));
  NO3        m1288(.A(mai_mai_n682_), .B(mai_mai_n765_), .C(mai_mai_n643_), .Y(mai_mai_n1317_));
  NOi21      m1289(.An(mai_mai_n1316_), .B(mai_mai_n1317_), .Y(mai_mai_n1318_));
  AN2        m1290(.A(mai_mai_n963_), .B(mai_mai_n654_), .Y(mai_mai_n1319_));
  NO4        m1291(.A(mai_mai_n1319_), .B(mai_mai_n1318_), .C(mai_mai_n1315_), .D(mai_mai_n1305_), .Y(mai_mai_n1320_));
  OAI220     m1292(.A0(mai_mai_n739_), .A1(mai_mai_n47_), .B0(mai_mai_n227_), .B1(mai_mai_n625_), .Y(mai_mai_n1321_));
  OAI210     m1293(.A0(mai_mai_n280_), .A1(c), .B0(mai_mai_n650_), .Y(mai_mai_n1322_));
  NA2        m1294(.A(mai_mai_n1322_), .B(mai_mai_n1321_), .Y(mai_mai_n1323_));
  NO3        m1295(.A(mai_mai_n246_), .B(mai_mai_n102_), .C(mai_mai_n287_), .Y(mai_mai_n1324_));
  OAI220     m1296(.A0(mai_mai_n707_), .A1(mai_mai_n251_), .B0(mai_mai_n521_), .B1(mai_mai_n525_), .Y(mai_mai_n1325_));
  OAI210     m1297(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1326_));
  NO3        m1298(.A(mai_mai_n1326_), .B(mai_mai_n606_), .C(j), .Y(mai_mai_n1327_));
  NOi21      m1299(.An(mai_mai_n1327_), .B(mai_mai_n677_), .Y(mai_mai_n1328_));
  NO4        m1300(.A(mai_mai_n1328_), .B(mai_mai_n1325_), .C(mai_mai_n1324_), .D(mai_mai_n1127_), .Y(mai_mai_n1329_));
  NA3        m1301(.A(mai_mai_n802_), .B(mai_mai_n801_), .C(mai_mai_n439_), .Y(mai_mai_n1330_));
  NAi31      m1302(.An(mai_mai_n755_), .B(mai_mai_n1330_), .C(mai_mai_n204_), .Y(mai_mai_n1331_));
  NA4        m1303(.A(mai_mai_n1331_), .B(mai_mai_n1329_), .C(mai_mai_n1323_), .D(mai_mai_n1217_), .Y(mai_mai_n1332_));
  NOi31      m1304(.An(mai_mai_n1298_), .B(mai_mai_n469_), .C(mai_mai_n397_), .Y(mai_mai_n1333_));
  OR3        m1305(.A(mai_mai_n1333_), .B(mai_mai_n790_), .C(mai_mai_n552_), .Y(mai_mai_n1334_));
  NA2        m1306(.A(mai_mai_n582_), .B(mai_mai_n451_), .Y(mai_mai_n1335_));
  NA2        m1307(.A(mai_mai_n1327_), .B(mai_mai_n798_), .Y(mai_mai_n1336_));
  NA3        m1308(.A(mai_mai_n1336_), .B(mai_mai_n1335_), .C(mai_mai_n1334_), .Y(mai_mai_n1337_));
  AN2        m1309(.A(mai_mai_n935_), .B(mai_mai_n934_), .Y(mai_mai_n1338_));
  NO4        m1310(.A(mai_mai_n1338_), .B(mai_mai_n883_), .C(mai_mai_n511_), .D(mai_mai_n489_), .Y(mai_mai_n1339_));
  NA2        m1311(.A(mai_mai_n1339_), .B(mai_mai_n1281_), .Y(mai_mai_n1340_));
  NAi21      m1312(.An(j), .B(i), .Y(mai_mai_n1341_));
  NO4        m1313(.A(mai_mai_n1292_), .B(mai_mai_n1341_), .C(mai_mai_n445_), .D(mai_mai_n237_), .Y(mai_mai_n1342_));
  NO4        m1314(.A(mai_mai_n1342_), .B(mai_mai_n1340_), .C(mai_mai_n1337_), .D(mai_mai_n1332_), .Y(mai_mai_n1343_));
  NA4        m1315(.A(mai_mai_n1343_), .B(mai_mai_n1320_), .C(mai_mai_n1301_), .D(mai_mai_n1294_), .Y(mai07));
  NOi21      m1316(.An(j), .B(k), .Y(mai_mai_n1345_));
  NA4        m1317(.A(mai_mai_n179_), .B(mai_mai_n108_), .C(mai_mai_n1345_), .D(f), .Y(mai_mai_n1346_));
  NAi32      m1318(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1347_));
  NO3        m1319(.A(mai_mai_n1347_), .B(g), .C(f), .Y(mai_mai_n1348_));
  OAI210     m1320(.A0(mai_mai_n318_), .A1(mai_mai_n491_), .B0(mai_mai_n1348_), .Y(mai_mai_n1349_));
  NAi21      m1321(.An(f), .B(c), .Y(mai_mai_n1350_));
  OR2        m1322(.A(e), .B(d), .Y(mai_mai_n1351_));
  OAI220     m1323(.A0(mai_mai_n1351_), .A1(mai_mai_n1350_), .B0(mai_mai_n638_), .B1(mai_mai_n320_), .Y(mai_mai_n1352_));
  NA3        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1070_), .C(mai_mai_n179_), .Y(mai_mai_n1353_));
  NOi31      m1325(.An(n), .B(m), .C(b), .Y(mai_mai_n1354_));
  NO3        m1326(.A(mai_mai_n133_), .B(mai_mai_n453_), .C(h), .Y(mai_mai_n1355_));
  NA3        m1327(.A(mai_mai_n1353_), .B(mai_mai_n1349_), .C(mai_mai_n1346_), .Y(mai_mai_n1356_));
  NOi41      m1328(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1357_));
  NOi21      m1329(.An(h), .B(k), .Y(mai_mai_n1358_));
  NO2        m1330(.A(k), .B(i), .Y(mai_mai_n1359_));
  NA3        m1331(.A(mai_mai_n1359_), .B(mai_mai_n903_), .C(mai_mai_n179_), .Y(mai_mai_n1360_));
  NA2        m1332(.A(mai_mai_n86_), .B(mai_mai_n45_), .Y(mai_mai_n1361_));
  NO2        m1333(.A(mai_mai_n1064_), .B(mai_mai_n445_), .Y(mai_mai_n1362_));
  NA3        m1334(.A(mai_mai_n1362_), .B(mai_mai_n1361_), .C(mai_mai_n216_), .Y(mai_mai_n1363_));
  NO2        m1335(.A(mai_mai_n1078_), .B(mai_mai_n304_), .Y(mai_mai_n1364_));
  NA2        m1336(.A(mai_mai_n553_), .B(mai_mai_n79_), .Y(mai_mai_n1365_));
  NA2        m1337(.A(mai_mai_n1218_), .B(mai_mai_n290_), .Y(mai_mai_n1366_));
  NA4        m1338(.A(mai_mai_n1366_), .B(mai_mai_n1365_), .C(mai_mai_n1363_), .D(mai_mai_n1360_), .Y(mai_mai_n1367_));
  NO2        m1339(.A(mai_mai_n1367_), .B(mai_mai_n1356_), .Y(mai_mai_n1368_));
  NO3        m1340(.A(e), .B(d), .C(c), .Y(mai_mai_n1369_));
  OAI210     m1341(.A0(mai_mai_n133_), .A1(mai_mai_n216_), .B0(mai_mai_n613_), .Y(mai_mai_n1370_));
  NA2        m1342(.A(mai_mai_n1370_), .B(mai_mai_n1369_), .Y(mai_mai_n1371_));
  NO2        m1343(.A(mai_mai_n1371_), .B(c), .Y(mai_mai_n1372_));
  OR2        m1344(.A(h), .B(f), .Y(mai_mai_n1373_));
  NO3        m1345(.A(n), .B(m), .C(i), .Y(mai_mai_n1374_));
  OAI210     m1346(.A0(mai_mai_n1126_), .A1(mai_mai_n156_), .B0(mai_mai_n1374_), .Y(mai_mai_n1375_));
  NO2        m1347(.A(mai_mai_n1375_), .B(mai_mai_n1373_), .Y(mai_mai_n1376_));
  NA3        m1348(.A(mai_mai_n704_), .B(mai_mai_n690_), .C(mai_mai_n112_), .Y(mai_mai_n1377_));
  NO2        m1349(.A(mai_mai_n1377_), .B(mai_mai_n45_), .Y(mai_mai_n1378_));
  NA2        m1350(.A(mai_mai_n1374_), .B(mai_mai_n649_), .Y(mai_mai_n1379_));
  NO2        m1351(.A(l), .B(k), .Y(mai_mai_n1380_));
  NOi41      m1352(.An(mai_mai_n558_), .B(mai_mai_n1380_), .C(mai_mai_n484_), .D(mai_mai_n445_), .Y(mai_mai_n1381_));
  NO3        m1353(.A(mai_mai_n445_), .B(d), .C(c), .Y(mai_mai_n1382_));
  NO4        m1354(.A(mai_mai_n1381_), .B(mai_mai_n1378_), .C(mai_mai_n1376_), .D(mai_mai_n1372_), .Y(mai_mai_n1383_));
  NO2        m1355(.A(mai_mai_n147_), .B(h), .Y(mai_mai_n1384_));
  NO2        m1356(.A(mai_mai_n1088_), .B(l), .Y(mai_mai_n1385_));
  NO2        m1357(.A(g), .B(c), .Y(mai_mai_n1386_));
  NA3        m1358(.A(mai_mai_n1386_), .B(mai_mai_n143_), .C(mai_mai_n187_), .Y(mai_mai_n1387_));
  NO2        m1359(.A(mai_mai_n1387_), .B(mai_mai_n1385_), .Y(mai_mai_n1388_));
  NA2        m1360(.A(mai_mai_n1388_), .B(mai_mai_n179_), .Y(mai_mai_n1389_));
  NA2        m1361(.A(mai_mai_n1358_), .B(mai_mai_n1088_), .Y(mai_mai_n1390_));
  NO2        m1362(.A(mai_mai_n456_), .B(a), .Y(mai_mai_n1391_));
  NA3        m1363(.A(mai_mai_n1391_), .B(mai_mai_n1390_), .C(mai_mai_n113_), .Y(mai_mai_n1392_));
  NO2        m1364(.A(i), .B(h), .Y(mai_mai_n1393_));
  NA2        m1365(.A(mai_mai_n1393_), .B(mai_mai_n223_), .Y(mai_mai_n1394_));
  AOI210     m1366(.A0(mai_mai_n1147_), .A1(h), .B0(mai_mai_n418_), .Y(mai_mai_n1395_));
  NA2        m1367(.A(mai_mai_n140_), .B(mai_mai_n223_), .Y(mai_mai_n1396_));
  AOI210     m1368(.A0(mai_mai_n261_), .A1(mai_mai_n116_), .B0(mai_mai_n541_), .Y(mai_mai_n1397_));
  OAI220     m1369(.A0(mai_mai_n1397_), .A1(mai_mai_n1394_), .B0(mai_mai_n1396_), .B1(mai_mai_n1395_), .Y(mai_mai_n1398_));
  NO2        m1370(.A(mai_mai_n762_), .B(mai_mai_n188_), .Y(mai_mai_n1399_));
  NOi31      m1371(.An(m), .B(n), .C(b), .Y(mai_mai_n1400_));
  NOi31      m1372(.An(f), .B(d), .C(c), .Y(mai_mai_n1401_));
  NA2        m1373(.A(mai_mai_n1401_), .B(mai_mai_n1400_), .Y(mai_mai_n1402_));
  INV        m1374(.A(mai_mai_n1402_), .Y(mai_mai_n1403_));
  NO3        m1375(.A(mai_mai_n1403_), .B(mai_mai_n1399_), .C(mai_mai_n1398_), .Y(mai_mai_n1404_));
  NA2        m1376(.A(mai_mai_n1098_), .B(mai_mai_n472_), .Y(mai_mai_n1405_));
  NO4        m1377(.A(mai_mai_n1405_), .B(mai_mai_n1073_), .C(mai_mai_n445_), .D(mai_mai_n45_), .Y(mai_mai_n1406_));
  OAI210     m1378(.A0(mai_mai_n182_), .A1(mai_mai_n536_), .B0(mai_mai_n1074_), .Y(mai_mai_n1407_));
  NO3        m1379(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1408_));
  INV        m1380(.A(mai_mai_n1407_), .Y(mai_mai_n1409_));
  NO2        m1381(.A(mai_mai_n1409_), .B(mai_mai_n1406_), .Y(mai_mai_n1410_));
  AN4        m1382(.A(mai_mai_n1410_), .B(mai_mai_n1404_), .C(mai_mai_n1392_), .D(mai_mai_n1389_), .Y(mai_mai_n1411_));
  NA2        m1383(.A(mai_mai_n1354_), .B(mai_mai_n381_), .Y(mai_mai_n1412_));
  NO2        m1384(.A(mai_mai_n1412_), .B(mai_mai_n1055_), .Y(mai_mai_n1413_));
  NA2        m1385(.A(mai_mai_n1382_), .B(mai_mai_n217_), .Y(mai_mai_n1414_));
  NO2        m1386(.A(mai_mai_n188_), .B(b), .Y(mai_mai_n1415_));
  AOI220     m1387(.A0(mai_mai_n1175_), .A1(mai_mai_n1415_), .B0(mai_mai_n1106_), .B1(mai_mai_n1405_), .Y(mai_mai_n1416_));
  NAi31      m1388(.An(mai_mai_n1413_), .B(mai_mai_n1416_), .C(mai_mai_n1414_), .Y(mai_mai_n1417_));
  NO4        m1389(.A(mai_mai_n133_), .B(g), .C(f), .D(e), .Y(mai_mai_n1418_));
  NA3        m1390(.A(mai_mai_n1359_), .B(mai_mai_n291_), .C(h), .Y(mai_mai_n1419_));
  NA2        m1391(.A(mai_mai_n195_), .B(mai_mai_n97_), .Y(mai_mai_n1420_));
  OR2        m1392(.A(e), .B(a), .Y(mai_mai_n1421_));
  NO2        m1393(.A(mai_mai_n1351_), .B(mai_mai_n1350_), .Y(mai_mai_n1422_));
  AOI210     m1394(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1422_), .Y(mai_mai_n1423_));
  NO2        m1395(.A(mai_mai_n1423_), .B(mai_mai_n1095_), .Y(mai_mai_n1424_));
  NA2        m1396(.A(mai_mai_n1357_), .B(mai_mai_n1380_), .Y(mai_mai_n1425_));
  INV        m1397(.A(mai_mai_n1425_), .Y(mai_mai_n1426_));
  OR3        m1398(.A(mai_mai_n552_), .B(mai_mai_n551_), .C(mai_mai_n112_), .Y(mai_mai_n1427_));
  NA2        m1399(.A(mai_mai_n1124_), .B(mai_mai_n410_), .Y(mai_mai_n1428_));
  OAI220     m1400(.A0(mai_mai_n1428_), .A1(mai_mai_n438_), .B0(mai_mai_n1427_), .B1(mai_mai_n296_), .Y(mai_mai_n1429_));
  AO210      m1401(.A0(mai_mai_n1429_), .A1(mai_mai_n116_), .B0(mai_mai_n1426_), .Y(mai_mai_n1430_));
  NO3        m1402(.A(mai_mai_n1430_), .B(mai_mai_n1424_), .C(mai_mai_n1417_), .Y(mai_mai_n1431_));
  NA4        m1403(.A(mai_mai_n1431_), .B(mai_mai_n1411_), .C(mai_mai_n1383_), .D(mai_mai_n1368_), .Y(mai_mai_n1432_));
  NO2        m1404(.A(mai_mai_n1139_), .B(mai_mai_n110_), .Y(mai_mai_n1433_));
  NA2        m1405(.A(mai_mai_n381_), .B(mai_mai_n56_), .Y(mai_mai_n1434_));
  AOI210     m1406(.A0(mai_mai_n1434_), .A1(mai_mai_n1064_), .B0(mai_mai_n1379_), .Y(mai_mai_n1435_));
  NA2        m1407(.A(mai_mai_n217_), .B(mai_mai_n179_), .Y(mai_mai_n1436_));
  AOI210     m1408(.A0(mai_mai_n1436_), .A1(mai_mai_n1193_), .B0(mai_mai_n1434_), .Y(mai_mai_n1437_));
  NO2        m1409(.A(mai_mai_n1099_), .B(mai_mai_n1095_), .Y(mai_mai_n1438_));
  NO3        m1410(.A(mai_mai_n1438_), .B(mai_mai_n1437_), .C(mai_mai_n1435_), .Y(mai_mai_n1439_));
  NO2        m1411(.A(mai_mai_n393_), .B(j), .Y(mai_mai_n1440_));
  NA3        m1412(.A(mai_mai_n1408_), .B(mai_mai_n1351_), .C(mai_mai_n1124_), .Y(mai_mai_n1441_));
  NAi41      m1413(.An(mai_mai_n1393_), .B(mai_mai_n1086_), .C(mai_mai_n167_), .D(mai_mai_n150_), .Y(mai_mai_n1442_));
  NA2        m1414(.A(mai_mai_n1442_), .B(mai_mai_n1441_), .Y(mai_mai_n1443_));
  NA3        m1415(.A(g), .B(mai_mai_n1440_), .C(mai_mai_n158_), .Y(mai_mai_n1444_));
  INV        m1416(.A(mai_mai_n1444_), .Y(mai_mai_n1445_));
  NO2        m1417(.A(mai_mai_n755_), .B(mai_mai_n174_), .Y(mai_mai_n1446_));
  NO3        m1418(.A(mai_mai_n1446_), .B(mai_mai_n1445_), .C(mai_mai_n1443_), .Y(mai_mai_n1447_));
  AOI210     m1419(.A0(mai_mai_n1436_), .A1(mai_mai_n1420_), .B0(mai_mai_n1064_), .Y(mai_mai_n1448_));
  OR2        m1420(.A(n), .B(i), .Y(mai_mai_n1449_));
  OAI210     m1421(.A0(mai_mai_n1449_), .A1(mai_mai_n1085_), .B0(mai_mai_n49_), .Y(mai_mai_n1450_));
  AOI220     m1422(.A0(mai_mai_n1450_), .A1(mai_mai_n1183_), .B0(mai_mai_n832_), .B1(mai_mai_n195_), .Y(mai_mai_n1451_));
  INV        m1423(.A(mai_mai_n1451_), .Y(mai_mai_n1452_));
  OAI220     m1424(.A0(mai_mai_n674_), .A1(g), .B0(mai_mai_n227_), .B1(c), .Y(mai_mai_n1453_));
  INV        m1425(.A(mai_mai_n1453_), .Y(mai_mai_n1454_));
  NO2        m1426(.A(mai_mai_n133_), .B(l), .Y(mai_mai_n1455_));
  NO2        m1427(.A(mai_mai_n227_), .B(k), .Y(mai_mai_n1456_));
  OAI210     m1428(.A0(mai_mai_n1456_), .A1(mai_mai_n1393_), .B0(mai_mai_n1455_), .Y(mai_mai_n1457_));
  OAI220     m1429(.A0(mai_mai_n1457_), .A1(mai_mai_n31_), .B0(mai_mai_n1454_), .B1(mai_mai_n176_), .Y(mai_mai_n1458_));
  NO3        m1430(.A(mai_mai_n1427_), .B(mai_mai_n472_), .C(mai_mai_n353_), .Y(mai_mai_n1459_));
  NO4        m1431(.A(mai_mai_n1459_), .B(mai_mai_n1458_), .C(mai_mai_n1452_), .D(mai_mai_n1448_), .Y(mai_mai_n1460_));
  NO3        m1432(.A(mai_mai_n1109_), .B(mai_mai_n1351_), .C(mai_mai_n49_), .Y(mai_mai_n1461_));
  NO2        m1433(.A(mai_mai_n1095_), .B(h), .Y(mai_mai_n1462_));
  NA3        m1434(.A(mai_mai_n1462_), .B(d), .C(mai_mai_n1056_), .Y(mai_mai_n1463_));
  NO2        m1435(.A(mai_mai_n1463_), .B(c), .Y(mai_mai_n1464_));
  NA3        m1436(.A(mai_mai_n1433_), .B(mai_mai_n472_), .C(f), .Y(mai_mai_n1465_));
  NA2        m1437(.A(mai_mai_n179_), .B(mai_mai_n112_), .Y(mai_mai_n1466_));
  NO2        m1438(.A(mai_mai_n1345_), .B(mai_mai_n42_), .Y(mai_mai_n1467_));
  AOI210     m1439(.A0(mai_mai_n113_), .A1(mai_mai_n40_), .B0(mai_mai_n1467_), .Y(mai_mai_n1468_));
  NO2        m1440(.A(mai_mai_n1468_), .B(mai_mai_n1465_), .Y(mai_mai_n1469_));
  NO2        m1441(.A(mai_mai_n1341_), .B(mai_mai_n174_), .Y(mai_mai_n1470_));
  NOi21      m1442(.An(d), .B(f), .Y(mai_mai_n1471_));
  NO2        m1443(.A(mai_mai_n1351_), .B(f), .Y(mai_mai_n1472_));
  NA2        m1444(.A(mai_mai_n1391_), .B(mai_mai_n1467_), .Y(mai_mai_n1473_));
  INV        m1445(.A(mai_mai_n1473_), .Y(mai_mai_n1474_));
  NO3        m1446(.A(mai_mai_n1474_), .B(mai_mai_n1469_), .C(mai_mai_n1464_), .Y(mai_mai_n1475_));
  NA4        m1447(.A(mai_mai_n1475_), .B(mai_mai_n1460_), .C(mai_mai_n1447_), .D(mai_mai_n1439_), .Y(mai_mai_n1476_));
  NO3        m1448(.A(mai_mai_n1098_), .B(mai_mai_n1085_), .C(mai_mai_n40_), .Y(mai_mai_n1477_));
  NO2        m1449(.A(mai_mai_n472_), .B(mai_mai_n296_), .Y(mai_mai_n1478_));
  OAI210     m1450(.A0(mai_mai_n1478_), .A1(mai_mai_n1477_), .B0(mai_mai_n1364_), .Y(mai_mai_n1479_));
  OAI210     m1451(.A0(mai_mai_n1418_), .A1(mai_mai_n1354_), .B0(mai_mai_n889_), .Y(mai_mai_n1480_));
  NO2        m1452(.A(mai_mai_n1052_), .B(mai_mai_n133_), .Y(mai_mai_n1481_));
  NA2        m1453(.A(mai_mai_n1481_), .B(mai_mai_n631_), .Y(mai_mai_n1482_));
  NA3        m1454(.A(mai_mai_n1482_), .B(mai_mai_n1480_), .C(mai_mai_n1479_), .Y(mai_mai_n1483_));
  NA2        m1455(.A(mai_mai_n1386_), .B(mai_mai_n1471_), .Y(mai_mai_n1484_));
  NO2        m1456(.A(mai_mai_n1484_), .B(m), .Y(mai_mai_n1485_));
  NO2        m1457(.A(mai_mai_n151_), .B(mai_mai_n181_), .Y(mai_mai_n1486_));
  OAI210     m1458(.A0(mai_mai_n1486_), .A1(mai_mai_n110_), .B0(mai_mai_n1400_), .Y(mai_mai_n1487_));
  INV        m1459(.A(mai_mai_n1487_), .Y(mai_mai_n1488_));
  NO3        m1460(.A(mai_mai_n1488_), .B(mai_mai_n1485_), .C(mai_mai_n1483_), .Y(mai_mai_n1489_));
  NO2        m1461(.A(mai_mai_n1350_), .B(e), .Y(mai_mai_n1490_));
  NA2        m1462(.A(mai_mai_n1490_), .B(mai_mai_n408_), .Y(mai_mai_n1491_));
  OAI210     m1463(.A0(mai_mai_n1472_), .A1(mai_mai_n1134_), .B0(mai_mai_n642_), .Y(mai_mai_n1492_));
  OR3        m1464(.A(mai_mai_n1456_), .B(mai_mai_n1218_), .C(mai_mai_n133_), .Y(mai_mai_n1493_));
  OAI220     m1465(.A0(mai_mai_n1493_), .A1(mai_mai_n1491_), .B0(mai_mai_n1492_), .B1(mai_mai_n447_), .Y(mai_mai_n1494_));
  NO3        m1466(.A(mai_mai_n1427_), .B(mai_mai_n353_), .C(a), .Y(mai_mai_n1495_));
  NO2        m1467(.A(mai_mai_n1495_), .B(mai_mai_n1494_), .Y(mai_mai_n1496_));
  NO2        m1468(.A(mai_mai_n181_), .B(c), .Y(mai_mai_n1497_));
  OAI210     m1469(.A0(mai_mai_n1497_), .A1(mai_mai_n1490_), .B0(mai_mai_n179_), .Y(mai_mai_n1498_));
  AOI220     m1470(.A0(mai_mai_n1498_), .A1(mai_mai_n1087_), .B0(mai_mai_n543_), .B1(mai_mai_n369_), .Y(mai_mai_n1499_));
  AOI210     m1471(.A0(i), .A1(mai_mai_n1382_), .B0(mai_mai_n1461_), .Y(mai_mai_n1500_));
  NO2        m1472(.A(mai_mai_n1421_), .B(f), .Y(mai_mai_n1501_));
  NA2        m1473(.A(mai_mai_n1134_), .B(a), .Y(mai_mai_n1502_));
  OAI220     m1474(.A0(mai_mai_n1502_), .A1(mai_mai_n66_), .B0(mai_mai_n1500_), .B1(mai_mai_n215_), .Y(mai_mai_n1503_));
  AOI210     m1475(.A0(mai_mai_n907_), .A1(mai_mai_n420_), .B0(mai_mai_n104_), .Y(mai_mai_n1504_));
  OR2        m1476(.A(mai_mai_n1504_), .B(mai_mai_n551_), .Y(mai_mai_n1505_));
  NA2        m1477(.A(mai_mai_n1501_), .B(mai_mai_n1361_), .Y(mai_mai_n1506_));
  OAI220     m1478(.A0(mai_mai_n1506_), .A1(mai_mai_n49_), .B0(mai_mai_n1505_), .B1(mai_mai_n174_), .Y(mai_mai_n1507_));
  NA4        m1479(.A(mai_mai_n1107_), .B(mai_mai_n1104_), .C(mai_mai_n223_), .D(mai_mai_n65_), .Y(mai_mai_n1508_));
  NA2        m1480(.A(mai_mai_n1355_), .B(mai_mai_n182_), .Y(mai_mai_n1509_));
  NO2        m1481(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1510_));
  OAI210     m1482(.A0(mai_mai_n1421_), .A1(mai_mai_n868_), .B0(mai_mai_n491_), .Y(mai_mai_n1511_));
  OAI210     m1483(.A0(mai_mai_n1511_), .A1(mai_mai_n1110_), .B0(mai_mai_n1510_), .Y(mai_mai_n1512_));
  NO2        m1484(.A(mai_mai_n256_), .B(g), .Y(mai_mai_n1513_));
  NO2        m1485(.A(m), .B(i), .Y(mai_mai_n1514_));
  BUFFER     m1486(.A(mai_mai_n1514_), .Y(mai_mai_n1515_));
  AOI220     m1487(.A0(mai_mai_n1515_), .A1(mai_mai_n1384_), .B0(mai_mai_n1086_), .B1(mai_mai_n1513_), .Y(mai_mai_n1516_));
  NA4        m1488(.A(mai_mai_n1516_), .B(mai_mai_n1512_), .C(mai_mai_n1509_), .D(mai_mai_n1508_), .Y(mai_mai_n1517_));
  NO4        m1489(.A(mai_mai_n1517_), .B(mai_mai_n1507_), .C(mai_mai_n1503_), .D(mai_mai_n1499_), .Y(mai_mai_n1518_));
  NA3        m1490(.A(mai_mai_n1518_), .B(mai_mai_n1496_), .C(mai_mai_n1489_), .Y(mai_mai_n1519_));
  NA3        m1491(.A(mai_mai_n969_), .B(mai_mai_n140_), .C(mai_mai_n46_), .Y(mai_mai_n1520_));
  AOI210     m1492(.A0(mai_mai_n148_), .A1(c), .B0(mai_mai_n1520_), .Y(mai_mai_n1521_));
  INV        m1493(.A(mai_mai_n185_), .Y(mai_mai_n1522_));
  NA2        m1494(.A(mai_mai_n1522_), .B(mai_mai_n1462_), .Y(mai_mai_n1523_));
  OR2        m1495(.A(mai_mai_n134_), .B(mai_mai_n1412_), .Y(mai_mai_n1524_));
  NO2        m1496(.A(mai_mai_n69_), .B(c), .Y(mai_mai_n1525_));
  NA2        m1497(.A(mai_mai_n1470_), .B(mai_mai_n1525_), .Y(mai_mai_n1526_));
  NA3        m1498(.A(mai_mai_n1526_), .B(mai_mai_n1524_), .C(mai_mai_n1523_), .Y(mai_mai_n1527_));
  NO2        m1499(.A(mai_mai_n1527_), .B(mai_mai_n1521_), .Y(mai_mai_n1528_));
  AOI210     m1500(.A0(mai_mai_n156_), .A1(mai_mai_n56_), .B0(mai_mai_n1490_), .Y(mai_mai_n1529_));
  NO2        m1501(.A(mai_mai_n1529_), .B(mai_mai_n1466_), .Y(mai_mai_n1530_));
  NOi21      m1502(.An(mai_mai_n1355_), .B(e), .Y(mai_mai_n1531_));
  NO2        m1503(.A(mai_mai_n1531_), .B(mai_mai_n1530_), .Y(mai_mai_n1532_));
  AN2        m1504(.A(mai_mai_n1107_), .B(mai_mai_n1093_), .Y(mai_mai_n1533_));
  AOI220     m1505(.A0(mai_mai_n1514_), .A1(mai_mai_n649_), .B0(mai_mai_n1070_), .B1(mai_mai_n159_), .Y(mai_mai_n1534_));
  NOi31      m1506(.An(mai_mai_n30_), .B(mai_mai_n1534_), .C(n), .Y(mai_mai_n1535_));
  AOI210     m1507(.A0(mai_mai_n1533_), .A1(mai_mai_n1175_), .B0(mai_mai_n1535_), .Y(mai_mai_n1536_));
  NO2        m1508(.A(mai_mai_n1465_), .B(mai_mai_n66_), .Y(mai_mai_n1537_));
  NA2        m1509(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1538_));
  NO2        m1510(.A(mai_mai_n1359_), .B(mai_mai_n118_), .Y(mai_mai_n1539_));
  OAI220     m1511(.A0(mai_mai_n1539_), .A1(mai_mai_n1412_), .B0(mai_mai_n1428_), .B1(mai_mai_n1538_), .Y(mai_mai_n1540_));
  NO2        m1512(.A(mai_mai_n1540_), .B(mai_mai_n1537_), .Y(mai_mai_n1541_));
  NA4        m1513(.A(mai_mai_n1541_), .B(mai_mai_n1536_), .C(mai_mai_n1532_), .D(mai_mai_n1528_), .Y(mai_mai_n1542_));
  OR4        m1514(.A(mai_mai_n1542_), .B(mai_mai_n1519_), .C(mai_mai_n1476_), .D(mai_mai_n1432_), .Y(mai04));
  NOi31      m1515(.An(mai_mai_n1418_), .B(mai_mai_n1419_), .C(mai_mai_n1058_), .Y(mai_mai_n1544_));
  NA2        m1516(.A(mai_mai_n1472_), .B(mai_mai_n832_), .Y(mai_mai_n1545_));
  NO4        m1517(.A(mai_mai_n1545_), .B(mai_mai_n1047_), .C(mai_mai_n492_), .D(j), .Y(mai_mai_n1546_));
  OR3        m1518(.A(mai_mai_n1546_), .B(mai_mai_n1544_), .C(mai_mai_n1076_), .Y(mai_mai_n1547_));
  NO2        m1519(.A(mai_mai_n1361_), .B(mai_mai_n89_), .Y(mai_mai_n1548_));
  AOI210     m1520(.A0(mai_mai_n1548_), .A1(mai_mai_n1069_), .B0(mai_mai_n1195_), .Y(mai_mai_n1549_));
  NA2        m1521(.A(mai_mai_n1549_), .B(mai_mai_n1222_), .Y(mai_mai_n1550_));
  NO4        m1522(.A(mai_mai_n1550_), .B(mai_mai_n1547_), .C(mai_mai_n1084_), .D(mai_mai_n1063_), .Y(mai_mai_n1551_));
  NA3        m1523(.A(mai_mai_n1551_), .B(mai_mai_n1136_), .C(mai_mai_n1113_), .Y(mai05));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  INV        u0023(.A(men_men_n51_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  NO2        u0026(.A(men_men_n54_), .B(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(g), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(g), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(g), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(g), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(g), .Y(men_men_n97_));
  AN2        u0069(.A(j), .B(g), .Y(men_men_n98_));
  NOi32      u0070(.An(m), .Bn(l), .C(i), .Y(men_men_n99_));
  NOi21      u0071(.An(g), .B(i), .Y(men_men_n100_));
  NOi32      u0072(.An(m), .Bn(j), .C(k), .Y(men_men_n101_));
  AOI220     u0073(.A0(men_men_n101_), .A1(men_men_n100_), .B0(men_men_n99_), .B1(men_men_n98_), .Y(men_men_n102_));
  NO2        u0074(.A(men_men_n95_), .B(men_men_n92_), .Y(men_men_n103_));
  NAi41      u0075(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n104_));
  AN2        u0076(.A(e), .B(b), .Y(men_men_n105_));
  NOi31      u0077(.An(c), .B(h), .C(f), .Y(men_men_n106_));
  NA2        u0078(.A(men_men_n106_), .B(men_men_n105_), .Y(men_men_n107_));
  NO2        u0079(.A(men_men_n107_), .B(men_men_n104_), .Y(men_men_n108_));
  NOi21      u0080(.An(g), .B(f), .Y(men_men_n109_));
  NOi21      u0081(.An(i), .B(h), .Y(men_men_n110_));
  INV        u0082(.A(a), .Y(men_men_n111_));
  NA2        u0083(.A(men_men_n105_), .B(men_men_n111_), .Y(men_men_n112_));
  INV        u0084(.A(l), .Y(men_men_n113_));
  NOi21      u0085(.An(m), .B(n), .Y(men_men_n114_));
  AN2        u0086(.A(k), .B(h), .Y(men_men_n115_));
  INV        u0087(.A(b), .Y(men_men_n116_));
  NA2        u0088(.A(l), .B(j), .Y(men_men_n117_));
  AN2        u0089(.A(k), .B(i), .Y(men_men_n118_));
  NA2        u0090(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n119_));
  NA2        u0091(.A(g), .B(e), .Y(men_men_n120_));
  NOi32      u0092(.An(c), .Bn(a), .C(d), .Y(men_men_n121_));
  NA2        u0093(.A(men_men_n121_), .B(men_men_n114_), .Y(men_men_n122_));
  NO4        u0094(.A(men_men_n122_), .B(men_men_n120_), .C(men_men_n119_), .D(men_men_n116_), .Y(men_men_n123_));
  NO2        u0095(.A(men_men_n123_), .B(men_men_n108_), .Y(men_men_n124_));
  OAI210     u0096(.A0(men_men_n103_), .A1(men_men_n88_), .B0(men_men_n124_), .Y(men_men_n125_));
  NOi31      u0097(.An(k), .B(m), .C(j), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(i), .Y(men_men_n127_));
  NOi32      u0099(.An(f), .Bn(b), .C(e), .Y(men_men_n128_));
  NAi21      u0100(.An(g), .B(h), .Y(men_men_n129_));
  NAi21      u0101(.An(m), .B(n), .Y(men_men_n130_));
  NAi21      u0102(.An(j), .B(k), .Y(men_men_n131_));
  NO3        u0103(.A(men_men_n131_), .B(men_men_n130_), .C(men_men_n129_), .Y(men_men_n132_));
  NAi41      u0104(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n133_));
  NAi31      u0105(.An(j), .B(k), .C(h), .Y(men_men_n134_));
  NA2        u0106(.A(men_men_n132_), .B(men_men_n128_), .Y(men_men_n135_));
  NO2        u0107(.A(k), .B(j), .Y(men_men_n136_));
  NO2        u0108(.A(men_men_n136_), .B(men_men_n130_), .Y(men_men_n137_));
  AN2        u0109(.A(k), .B(j), .Y(men_men_n138_));
  NAi21      u0110(.An(c), .B(b), .Y(men_men_n139_));
  NA2        u0111(.A(f), .B(d), .Y(men_men_n140_));
  NO4        u0112(.A(men_men_n140_), .B(men_men_n139_), .C(men_men_n138_), .D(men_men_n129_), .Y(men_men_n141_));
  NAi31      u0113(.An(f), .B(e), .C(b), .Y(men_men_n142_));
  NA2        u0114(.A(men_men_n141_), .B(men_men_n137_), .Y(men_men_n143_));
  NA2        u0115(.A(d), .B(b), .Y(men_men_n144_));
  NAi21      u0116(.An(e), .B(f), .Y(men_men_n145_));
  NO2        u0117(.A(men_men_n145_), .B(men_men_n144_), .Y(men_men_n146_));
  NA2        u0118(.A(b), .B(a), .Y(men_men_n147_));
  NAi21      u0119(.An(e), .B(g), .Y(men_men_n148_));
  NAi21      u0120(.An(c), .B(d), .Y(men_men_n149_));
  NAi31      u0121(.An(l), .B(k), .C(h), .Y(men_men_n150_));
  NO2        u0122(.A(men_men_n130_), .B(men_men_n150_), .Y(men_men_n151_));
  NA2        u0123(.A(men_men_n151_), .B(men_men_n146_), .Y(men_men_n152_));
  NA3        u0124(.A(men_men_n152_), .B(men_men_n143_), .C(men_men_n135_), .Y(men_men_n153_));
  NAi31      u0125(.An(e), .B(f), .C(b), .Y(men_men_n154_));
  NOi21      u0126(.An(g), .B(d), .Y(men_men_n155_));
  NO2        u0127(.A(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  NOi21      u0128(.An(h), .B(i), .Y(men_men_n157_));
  NOi21      u0129(.An(k), .B(m), .Y(men_men_n158_));
  NA3        u0130(.A(men_men_n158_), .B(men_men_n157_), .C(n), .Y(men_men_n159_));
  NOi21      u0131(.An(men_men_n156_), .B(men_men_n159_), .Y(men_men_n160_));
  NOi21      u0132(.An(h), .B(g), .Y(men_men_n161_));
  NO2        u0133(.A(men_men_n140_), .B(men_men_n139_), .Y(men_men_n162_));
  NA2        u0134(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  NAi31      u0135(.An(l), .B(j), .C(h), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n164_), .B(men_men_n49_), .Y(men_men_n165_));
  NA2        u0137(.A(men_men_n165_), .B(men_men_n67_), .Y(men_men_n166_));
  NOi32      u0138(.An(n), .Bn(k), .C(m), .Y(men_men_n167_));
  NA2        u0139(.A(l), .B(i), .Y(men_men_n168_));
  NA2        u0140(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  OAI210     u0141(.A0(men_men_n169_), .A1(men_men_n163_), .B0(men_men_n166_), .Y(men_men_n170_));
  NAi31      u0142(.An(d), .B(f), .C(c), .Y(men_men_n171_));
  NAi31      u0143(.An(e), .B(f), .C(c), .Y(men_men_n172_));
  NA2        u0144(.A(men_men_n172_), .B(men_men_n171_), .Y(men_men_n173_));
  NA2        u0145(.A(j), .B(h), .Y(men_men_n174_));
  OR3        u0146(.A(n), .B(m), .C(k), .Y(men_men_n175_));
  NO2        u0147(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  NAi32      u0148(.An(m), .Bn(k), .C(n), .Y(men_men_n177_));
  NO2        u0149(.A(men_men_n177_), .B(men_men_n174_), .Y(men_men_n178_));
  AOI220     u0150(.A0(men_men_n178_), .A1(men_men_n156_), .B0(men_men_n176_), .B1(men_men_n173_), .Y(men_men_n179_));
  NO2        u0151(.A(n), .B(m), .Y(men_men_n180_));
  NA2        u0152(.A(men_men_n180_), .B(men_men_n50_), .Y(men_men_n181_));
  NAi21      u0153(.An(f), .B(e), .Y(men_men_n182_));
  NA2        u0154(.A(d), .B(c), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  NOi21      u0156(.An(men_men_n184_), .B(men_men_n181_), .Y(men_men_n185_));
  NAi21      u0157(.An(d), .B(c), .Y(men_men_n186_));
  NAi31      u0158(.An(m), .B(n), .C(b), .Y(men_men_n187_));
  NA2        u0159(.A(k), .B(i), .Y(men_men_n188_));
  NAi21      u0160(.An(h), .B(f), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NO2        u0162(.A(men_men_n187_), .B(men_men_n149_), .Y(men_men_n191_));
  NA2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NOi32      u0164(.An(f), .Bn(c), .C(d), .Y(men_men_n193_));
  NOi32      u0165(.An(f), .Bn(c), .C(e), .Y(men_men_n194_));
  NO2        u0166(.A(men_men_n194_), .B(men_men_n193_), .Y(men_men_n195_));
  NO3        u0167(.A(n), .B(m), .C(j), .Y(men_men_n196_));
  NA2        u0168(.A(men_men_n196_), .B(men_men_n115_), .Y(men_men_n197_));
  AO210      u0169(.A0(men_men_n197_), .A1(men_men_n181_), .B0(men_men_n195_), .Y(men_men_n198_));
  NAi41      u0170(.An(men_men_n185_), .B(men_men_n198_), .C(men_men_n192_), .D(men_men_n179_), .Y(men_men_n199_));
  OR4        u0171(.A(men_men_n199_), .B(men_men_n170_), .C(men_men_n160_), .D(men_men_n153_), .Y(men_men_n200_));
  NO4        u0172(.A(men_men_n200_), .B(men_men_n125_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n201_));
  NA3        u0173(.A(m), .B(men_men_n113_), .C(j), .Y(men_men_n202_));
  NAi31      u0174(.An(n), .B(h), .C(g), .Y(men_men_n203_));
  NO2        u0175(.A(men_men_n203_), .B(men_men_n202_), .Y(men_men_n204_));
  NOi32      u0176(.An(m), .Bn(k), .C(l), .Y(men_men_n205_));
  NA3        u0177(.A(men_men_n205_), .B(men_men_n89_), .C(g), .Y(men_men_n206_));
  NO2        u0178(.A(men_men_n206_), .B(n), .Y(men_men_n207_));
  NOi21      u0179(.An(k), .B(j), .Y(men_men_n208_));
  AN2        u0180(.A(i), .B(g), .Y(men_men_n209_));
  NA3        u0181(.A(men_men_n76_), .B(men_men_n209_), .C(men_men_n114_), .Y(men_men_n210_));
  NO2        u0182(.A(men_men_n207_), .B(men_men_n204_), .Y(men_men_n211_));
  NAi41      u0183(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n212_));
  INV        u0184(.A(men_men_n212_), .Y(men_men_n213_));
  INV        u0185(.A(f), .Y(men_men_n214_));
  INV        u0186(.A(g), .Y(men_men_n215_));
  NOi31      u0187(.An(i), .B(j), .C(h), .Y(men_men_n216_));
  NOi21      u0188(.An(l), .B(m), .Y(men_men_n217_));
  NA2        u0189(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n218_));
  NO3        u0190(.A(men_men_n218_), .B(men_men_n215_), .C(men_men_n214_), .Y(men_men_n219_));
  NA2        u0191(.A(men_men_n219_), .B(men_men_n213_), .Y(men_men_n220_));
  OAI210     u0192(.A0(men_men_n211_), .A1(men_men_n32_), .B0(men_men_n220_), .Y(men_men_n221_));
  NOi21      u0193(.An(n), .B(m), .Y(men_men_n222_));
  NOi32      u0194(.An(l), .Bn(i), .C(j), .Y(men_men_n223_));
  NA2        u0195(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n224_));
  OA220      u0196(.A0(men_men_n224_), .A1(men_men_n107_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n225_));
  NAi21      u0197(.An(j), .B(h), .Y(men_men_n226_));
  XN2        u0198(.A(i), .B(h), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n228_));
  NOi31      u0200(.An(k), .B(n), .C(m), .Y(men_men_n229_));
  NOi31      u0201(.An(men_men_n229_), .B(men_men_n183_), .C(men_men_n182_), .Y(men_men_n230_));
  NA2        u0202(.A(men_men_n230_), .B(men_men_n228_), .Y(men_men_n231_));
  NAi31      u0203(.An(f), .B(e), .C(c), .Y(men_men_n232_));
  NO4        u0204(.A(men_men_n232_), .B(men_men_n175_), .C(men_men_n174_), .D(men_men_n59_), .Y(men_men_n233_));
  NA4        u0205(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n234_));
  NAi32      u0206(.An(m), .Bn(i), .C(k), .Y(men_men_n235_));
  NO3        u0207(.A(men_men_n235_), .B(men_men_n93_), .C(men_men_n234_), .Y(men_men_n236_));
  INV        u0208(.A(k), .Y(men_men_n237_));
  NO2        u0209(.A(men_men_n236_), .B(men_men_n233_), .Y(men_men_n238_));
  NAi21      u0210(.An(n), .B(a), .Y(men_men_n239_));
  NO2        u0211(.A(men_men_n239_), .B(men_men_n144_), .Y(men_men_n240_));
  NAi41      u0212(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(e), .Y(men_men_n242_));
  NO3        u0214(.A(men_men_n145_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n243_));
  OAI210     u0215(.A0(men_men_n243_), .A1(men_men_n242_), .B0(men_men_n240_), .Y(men_men_n244_));
  AN4        u0216(.A(men_men_n244_), .B(men_men_n238_), .C(men_men_n231_), .D(men_men_n225_), .Y(men_men_n245_));
  OR2        u0217(.A(h), .B(g), .Y(men_men_n246_));
  NO2        u0218(.A(men_men_n246_), .B(men_men_n104_), .Y(men_men_n247_));
  NA2        u0219(.A(men_men_n247_), .B(men_men_n128_), .Y(men_men_n248_));
  NA2        u0220(.A(men_men_n158_), .B(men_men_n110_), .Y(men_men_n249_));
  NO2        u0221(.A(n), .B(a), .Y(men_men_n250_));
  NAi31      u0222(.An(men_men_n241_), .B(men_men_n250_), .C(men_men_n105_), .Y(men_men_n251_));
  NAi21      u0223(.An(h), .B(i), .Y(men_men_n252_));
  NA2        u0224(.A(men_men_n180_), .B(k), .Y(men_men_n253_));
  NO2        u0225(.A(men_men_n253_), .B(men_men_n252_), .Y(men_men_n254_));
  NA2        u0226(.A(men_men_n254_), .B(men_men_n193_), .Y(men_men_n255_));
  NA3        u0227(.A(men_men_n255_), .B(men_men_n251_), .C(men_men_n248_), .Y(men_men_n256_));
  NOi21      u0228(.An(g), .B(e), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n258_));
  NA2        u0230(.A(men_men_n258_), .B(men_men_n257_), .Y(men_men_n259_));
  NOi32      u0231(.An(l), .Bn(j), .C(i), .Y(men_men_n260_));
  AOI210     u0232(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n260_), .Y(men_men_n261_));
  NAi21      u0233(.An(f), .B(g), .Y(men_men_n262_));
  NO2        u0234(.A(men_men_n262_), .B(men_men_n65_), .Y(men_men_n263_));
  NO2        u0235(.A(men_men_n69_), .B(men_men_n117_), .Y(men_men_n264_));
  NO2        u0236(.A(men_men_n261_), .B(men_men_n259_), .Y(men_men_n265_));
  NO3        u0237(.A(men_men_n131_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n266_));
  NOi41      u0238(.An(men_men_n245_), .B(men_men_n265_), .C(men_men_n256_), .D(men_men_n221_), .Y(men_men_n267_));
  NO4        u0239(.A(men_men_n204_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n268_));
  NO2        u0240(.A(men_men_n268_), .B(men_men_n112_), .Y(men_men_n269_));
  NA3        u0241(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n270_));
  NAi21      u0242(.An(h), .B(g), .Y(men_men_n271_));
  OR4        u0243(.A(men_men_n271_), .B(men_men_n270_), .C(men_men_n224_), .D(e), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n249_), .B(men_men_n262_), .Y(men_men_n273_));
  NAi31      u0245(.An(g), .B(k), .C(h), .Y(men_men_n274_));
  NO3        u0246(.A(men_men_n130_), .B(men_men_n274_), .C(l), .Y(men_men_n275_));
  NAi31      u0247(.An(e), .B(d), .C(a), .Y(men_men_n276_));
  NA2        u0248(.A(men_men_n275_), .B(men_men_n128_), .Y(men_men_n277_));
  NA2        u0249(.A(men_men_n277_), .B(men_men_n272_), .Y(men_men_n278_));
  NA4        u0250(.A(men_men_n158_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n117_), .Y(men_men_n279_));
  NA3        u0251(.A(men_men_n158_), .B(men_men_n157_), .C(men_men_n86_), .Y(men_men_n280_));
  NO2        u0252(.A(men_men_n280_), .B(men_men_n195_), .Y(men_men_n281_));
  NOi21      u0253(.An(men_men_n279_), .B(men_men_n281_), .Y(men_men_n282_));
  NA3        u0254(.A(e), .B(c), .C(b), .Y(men_men_n283_));
  NO2        u0255(.A(men_men_n60_), .B(men_men_n283_), .Y(men_men_n284_));
  NAi32      u0256(.An(k), .Bn(i), .C(j), .Y(men_men_n285_));
  NAi31      u0257(.An(h), .B(l), .C(i), .Y(men_men_n286_));
  NA3        u0258(.A(men_men_n286_), .B(men_men_n285_), .C(men_men_n164_), .Y(men_men_n287_));
  NOi21      u0259(.An(men_men_n287_), .B(men_men_n49_), .Y(men_men_n288_));
  OAI210     u0260(.A0(men_men_n263_), .A1(men_men_n284_), .B0(men_men_n288_), .Y(men_men_n289_));
  NAi21      u0261(.An(l), .B(k), .Y(men_men_n290_));
  NO2        u0262(.A(men_men_n290_), .B(men_men_n49_), .Y(men_men_n291_));
  NOi21      u0263(.An(l), .B(j), .Y(men_men_n292_));
  NA2        u0264(.A(men_men_n161_), .B(men_men_n292_), .Y(men_men_n293_));
  NA3        u0265(.A(men_men_n118_), .B(men_men_n117_), .C(g), .Y(men_men_n294_));
  OR3        u0266(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n295_));
  AOI210     u0267(.A0(men_men_n294_), .A1(men_men_n293_), .B0(men_men_n295_), .Y(men_men_n296_));
  INV        u0268(.A(men_men_n296_), .Y(men_men_n297_));
  NAi32      u0269(.An(j), .Bn(h), .C(i), .Y(men_men_n298_));
  NAi21      u0270(.An(m), .B(l), .Y(men_men_n299_));
  NO3        u0271(.A(men_men_n299_), .B(men_men_n298_), .C(men_men_n86_), .Y(men_men_n300_));
  NA2        u0272(.A(h), .B(g), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n300_), .B(men_men_n162_), .Y(men_men_n302_));
  NA4        u0274(.A(men_men_n302_), .B(men_men_n297_), .C(men_men_n289_), .D(men_men_n282_), .Y(men_men_n303_));
  NO2        u0275(.A(men_men_n142_), .B(d), .Y(men_men_n304_));
  NA2        u0276(.A(men_men_n304_), .B(men_men_n53_), .Y(men_men_n305_));
  NO2        u0277(.A(men_men_n107_), .B(men_men_n104_), .Y(men_men_n306_));
  NAi32      u0278(.An(n), .Bn(m), .C(l), .Y(men_men_n307_));
  NO2        u0279(.A(men_men_n307_), .B(men_men_n298_), .Y(men_men_n308_));
  NA2        u0280(.A(men_men_n308_), .B(men_men_n184_), .Y(men_men_n309_));
  NO2        u0281(.A(men_men_n122_), .B(men_men_n116_), .Y(men_men_n310_));
  NAi31      u0282(.An(k), .B(l), .C(j), .Y(men_men_n311_));
  OAI210     u0283(.A0(men_men_n290_), .A1(j), .B0(men_men_n311_), .Y(men_men_n312_));
  NOi21      u0284(.An(men_men_n312_), .B(men_men_n120_), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n313_), .B(men_men_n310_), .Y(men_men_n314_));
  NA3        u0286(.A(men_men_n314_), .B(men_men_n309_), .C(men_men_n305_), .Y(men_men_n315_));
  NO4        u0287(.A(men_men_n315_), .B(men_men_n303_), .C(men_men_n278_), .D(men_men_n269_), .Y(men_men_n316_));
  NA2        u0288(.A(men_men_n254_), .B(men_men_n194_), .Y(men_men_n317_));
  NAi21      u0289(.An(m), .B(k), .Y(men_men_n318_));
  NO2        u0290(.A(men_men_n227_), .B(men_men_n318_), .Y(men_men_n319_));
  NAi41      u0291(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n320_), .B(men_men_n148_), .Y(men_men_n321_));
  NA2        u0293(.A(men_men_n321_), .B(men_men_n319_), .Y(men_men_n322_));
  NAi31      u0294(.An(i), .B(l), .C(h), .Y(men_men_n323_));
  NA2        u0295(.A(e), .B(c), .Y(men_men_n324_));
  NO3        u0296(.A(men_men_n324_), .B(n), .C(d), .Y(men_men_n325_));
  NOi21      u0297(.An(f), .B(h), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n326_), .B(men_men_n118_), .Y(men_men_n327_));
  NO2        u0299(.A(men_men_n327_), .B(men_men_n215_), .Y(men_men_n328_));
  NAi31      u0300(.An(d), .B(e), .C(b), .Y(men_men_n329_));
  NO2        u0301(.A(men_men_n130_), .B(men_men_n329_), .Y(men_men_n330_));
  NA2        u0302(.A(men_men_n330_), .B(men_men_n328_), .Y(men_men_n331_));
  NA3        u0303(.A(men_men_n331_), .B(men_men_n322_), .C(men_men_n317_), .Y(men_men_n332_));
  NO4        u0304(.A(men_men_n320_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n215_), .Y(men_men_n333_));
  NA2        u0305(.A(men_men_n250_), .B(men_men_n105_), .Y(men_men_n334_));
  OR2        u0306(.A(men_men_n334_), .B(men_men_n206_), .Y(men_men_n335_));
  NOi31      u0307(.An(l), .B(n), .C(m), .Y(men_men_n336_));
  NA2        u0308(.A(men_men_n336_), .B(men_men_n216_), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n337_), .B(men_men_n195_), .Y(men_men_n338_));
  NAi32      u0310(.An(men_men_n338_), .Bn(men_men_n333_), .C(men_men_n335_), .Y(men_men_n339_));
  NAi32      u0311(.An(m), .Bn(j), .C(k), .Y(men_men_n340_));
  NAi41      u0312(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n341_));
  OAI210     u0313(.A0(men_men_n212_), .A1(men_men_n340_), .B0(men_men_n341_), .Y(men_men_n342_));
  NOi31      u0314(.An(j), .B(m), .C(k), .Y(men_men_n343_));
  NO2        u0315(.A(men_men_n126_), .B(men_men_n343_), .Y(men_men_n344_));
  AN3        u0316(.A(h), .B(g), .C(f), .Y(men_men_n345_));
  NAi31      u0317(.An(men_men_n344_), .B(men_men_n345_), .C(men_men_n342_), .Y(men_men_n346_));
  NOi32      u0318(.An(m), .Bn(j), .C(l), .Y(men_men_n347_));
  NO2        u0319(.A(men_men_n347_), .B(men_men_n99_), .Y(men_men_n348_));
  NAi32      u0320(.An(men_men_n348_), .Bn(men_men_n203_), .C(men_men_n304_), .Y(men_men_n349_));
  NO2        u0321(.A(men_men_n299_), .B(men_men_n298_), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n218_), .B(g), .Y(men_men_n351_));
  NO2        u0323(.A(men_men_n154_), .B(men_men_n86_), .Y(men_men_n352_));
  NA2        u0324(.A(men_men_n352_), .B(men_men_n351_), .Y(men_men_n353_));
  NA2        u0325(.A(men_men_n235_), .B(men_men_n81_), .Y(men_men_n354_));
  NA3        u0326(.A(men_men_n354_), .B(men_men_n345_), .C(men_men_n213_), .Y(men_men_n355_));
  NA4        u0327(.A(men_men_n355_), .B(men_men_n353_), .C(men_men_n349_), .D(men_men_n346_), .Y(men_men_n356_));
  NA3        u0328(.A(h), .B(g), .C(f), .Y(men_men_n357_));
  NO2        u0329(.A(men_men_n357_), .B(men_men_n77_), .Y(men_men_n358_));
  NA2        u0330(.A(men_men_n341_), .B(men_men_n212_), .Y(men_men_n359_));
  NA2        u0331(.A(men_men_n161_), .B(e), .Y(men_men_n360_));
  NO2        u0332(.A(men_men_n360_), .B(men_men_n41_), .Y(men_men_n361_));
  AOI220     u0333(.A0(men_men_n361_), .A1(men_men_n310_), .B0(men_men_n359_), .B1(men_men_n358_), .Y(men_men_n362_));
  NOi32      u0334(.An(j), .Bn(g), .C(i), .Y(men_men_n363_));
  NA3        u0335(.A(men_men_n363_), .B(men_men_n290_), .C(men_men_n114_), .Y(men_men_n364_));
  AO210      u0336(.A0(men_men_n112_), .A1(men_men_n32_), .B0(men_men_n364_), .Y(men_men_n365_));
  NOi32      u0337(.An(e), .Bn(b), .C(a), .Y(men_men_n366_));
  AN2        u0338(.A(l), .B(j), .Y(men_men_n367_));
  NO2        u0339(.A(men_men_n318_), .B(men_men_n367_), .Y(men_men_n368_));
  NO3        u0340(.A(men_men_n320_), .B(men_men_n72_), .C(men_men_n215_), .Y(men_men_n369_));
  NA2        u0341(.A(men_men_n210_), .B(men_men_n35_), .Y(men_men_n370_));
  AOI220     u0342(.A0(men_men_n370_), .A1(men_men_n366_), .B0(men_men_n369_), .B1(men_men_n368_), .Y(men_men_n371_));
  NA2        u0343(.A(men_men_n209_), .B(k), .Y(men_men_n372_));
  NA3        u0344(.A(m), .B(men_men_n113_), .C(men_men_n214_), .Y(men_men_n373_));
  NA4        u0345(.A(men_men_n205_), .B(men_men_n89_), .C(g), .D(men_men_n214_), .Y(men_men_n374_));
  NAi41      u0346(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n375_));
  NA2        u0347(.A(men_men_n51_), .B(men_men_n114_), .Y(men_men_n376_));
  NO2        u0348(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n377_));
  NA2        u0349(.A(men_men_n377_), .B(b), .Y(men_men_n378_));
  NA4        u0350(.A(men_men_n378_), .B(men_men_n371_), .C(men_men_n365_), .D(men_men_n362_), .Y(men_men_n379_));
  NO4        u0351(.A(men_men_n379_), .B(men_men_n356_), .C(men_men_n339_), .D(men_men_n332_), .Y(men_men_n380_));
  NA4        u0352(.A(men_men_n380_), .B(men_men_n316_), .C(men_men_n267_), .D(men_men_n201_), .Y(men10));
  NA3        u0353(.A(m), .B(k), .C(i), .Y(men_men_n382_));
  NO3        u0354(.A(men_men_n382_), .B(j), .C(men_men_n215_), .Y(men_men_n383_));
  NOi21      u0355(.An(e), .B(f), .Y(men_men_n384_));
  NO4        u0356(.A(men_men_n149_), .B(men_men_n384_), .C(n), .D(men_men_n111_), .Y(men_men_n385_));
  NAi31      u0357(.An(b), .B(f), .C(c), .Y(men_men_n386_));
  INV        u0358(.A(men_men_n386_), .Y(men_men_n387_));
  NOi32      u0359(.An(k), .Bn(h), .C(j), .Y(men_men_n388_));
  NA2        u0360(.A(men_men_n388_), .B(men_men_n222_), .Y(men_men_n389_));
  NA2        u0361(.A(men_men_n159_), .B(men_men_n389_), .Y(men_men_n390_));
  AOI220     u0362(.A0(men_men_n390_), .A1(men_men_n387_), .B0(men_men_n385_), .B1(men_men_n383_), .Y(men_men_n391_));
  AN2        u0363(.A(j), .B(h), .Y(men_men_n392_));
  NO3        u0364(.A(n), .B(m), .C(k), .Y(men_men_n393_));
  NA2        u0365(.A(men_men_n393_), .B(men_men_n392_), .Y(men_men_n394_));
  NO3        u0366(.A(men_men_n394_), .B(men_men_n149_), .C(men_men_n214_), .Y(men_men_n395_));
  OR2        u0367(.A(m), .B(k), .Y(men_men_n396_));
  NO2        u0368(.A(men_men_n174_), .B(men_men_n396_), .Y(men_men_n397_));
  NA4        u0369(.A(n), .B(f), .C(c), .D(men_men_n116_), .Y(men_men_n398_));
  NOi21      u0370(.An(men_men_n397_), .B(men_men_n398_), .Y(men_men_n399_));
  NOi32      u0371(.An(d), .Bn(a), .C(c), .Y(men_men_n400_));
  NA2        u0372(.A(men_men_n400_), .B(men_men_n182_), .Y(men_men_n401_));
  NAi21      u0373(.An(i), .B(g), .Y(men_men_n402_));
  NAi31      u0374(.An(k), .B(m), .C(j), .Y(men_men_n403_));
  NO3        u0375(.A(men_men_n403_), .B(men_men_n402_), .C(n), .Y(men_men_n404_));
  NOi21      u0376(.An(men_men_n404_), .B(men_men_n401_), .Y(men_men_n405_));
  NO3        u0377(.A(men_men_n405_), .B(men_men_n399_), .C(men_men_n395_), .Y(men_men_n406_));
  NO2        u0378(.A(men_men_n398_), .B(men_men_n299_), .Y(men_men_n407_));
  NOi32      u0379(.An(f), .Bn(d), .C(c), .Y(men_men_n408_));
  AOI220     u0380(.A0(men_men_n408_), .A1(men_men_n308_), .B0(men_men_n407_), .B1(men_men_n216_), .Y(men_men_n409_));
  NA3        u0381(.A(men_men_n409_), .B(men_men_n406_), .C(men_men_n391_), .Y(men_men_n410_));
  NO2        u0382(.A(men_men_n59_), .B(men_men_n116_), .Y(men_men_n411_));
  NA2        u0383(.A(men_men_n250_), .B(men_men_n411_), .Y(men_men_n412_));
  INV        u0384(.A(e), .Y(men_men_n413_));
  NA2        u0385(.A(men_men_n46_), .B(e), .Y(men_men_n414_));
  OAI220     u0386(.A0(men_men_n414_), .A1(men_men_n202_), .B0(men_men_n206_), .B1(men_men_n413_), .Y(men_men_n415_));
  AN2        u0387(.A(g), .B(e), .Y(men_men_n416_));
  NA3        u0388(.A(men_men_n416_), .B(men_men_n205_), .C(i), .Y(men_men_n417_));
  INV        u0389(.A(men_men_n417_), .Y(men_men_n418_));
  NO2        u0390(.A(men_men_n102_), .B(men_men_n413_), .Y(men_men_n419_));
  NO3        u0391(.A(men_men_n419_), .B(men_men_n418_), .C(men_men_n415_), .Y(men_men_n420_));
  NOi32      u0392(.An(h), .Bn(e), .C(g), .Y(men_men_n421_));
  NA3        u0393(.A(men_men_n421_), .B(men_men_n292_), .C(m), .Y(men_men_n422_));
  NOi21      u0394(.An(g), .B(h), .Y(men_men_n423_));
  AN3        u0395(.A(m), .B(l), .C(i), .Y(men_men_n424_));
  NA3        u0396(.A(men_men_n424_), .B(men_men_n423_), .C(e), .Y(men_men_n425_));
  AN3        u0397(.A(h), .B(g), .C(e), .Y(men_men_n426_));
  NA2        u0398(.A(men_men_n426_), .B(men_men_n99_), .Y(men_men_n427_));
  AN3        u0399(.A(men_men_n427_), .B(men_men_n425_), .C(men_men_n422_), .Y(men_men_n428_));
  AOI210     u0400(.A0(men_men_n428_), .A1(men_men_n420_), .B0(men_men_n412_), .Y(men_men_n429_));
  NA3        u0401(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n430_));
  NO2        u0402(.A(men_men_n430_), .B(men_men_n412_), .Y(men_men_n431_));
  NAi31      u0403(.An(b), .B(c), .C(a), .Y(men_men_n432_));
  NO2        u0404(.A(men_men_n432_), .B(n), .Y(men_men_n433_));
  NA2        u0405(.A(men_men_n51_), .B(m), .Y(men_men_n434_));
  NO2        u0406(.A(men_men_n434_), .B(men_men_n145_), .Y(men_men_n435_));
  NA2        u0407(.A(men_men_n435_), .B(men_men_n433_), .Y(men_men_n436_));
  INV        u0408(.A(men_men_n436_), .Y(men_men_n437_));
  NO4        u0409(.A(men_men_n437_), .B(men_men_n431_), .C(men_men_n429_), .D(men_men_n410_), .Y(men_men_n438_));
  NA2        u0410(.A(i), .B(g), .Y(men_men_n439_));
  NO3        u0411(.A(men_men_n276_), .B(men_men_n439_), .C(c), .Y(men_men_n440_));
  NOi21      u0412(.An(a), .B(n), .Y(men_men_n441_));
  NOi21      u0413(.An(d), .B(c), .Y(men_men_n442_));
  NA2        u0414(.A(men_men_n442_), .B(men_men_n441_), .Y(men_men_n443_));
  NA3        u0415(.A(i), .B(g), .C(f), .Y(men_men_n444_));
  OR2        u0416(.A(men_men_n444_), .B(men_men_n71_), .Y(men_men_n445_));
  NA3        u0417(.A(men_men_n424_), .B(men_men_n423_), .C(men_men_n182_), .Y(men_men_n446_));
  AOI210     u0418(.A0(men_men_n446_), .A1(men_men_n445_), .B0(men_men_n443_), .Y(men_men_n447_));
  AOI210     u0419(.A0(men_men_n440_), .A1(men_men_n291_), .B0(men_men_n447_), .Y(men_men_n448_));
  OR2        u0420(.A(n), .B(m), .Y(men_men_n449_));
  NO2        u0421(.A(men_men_n449_), .B(men_men_n150_), .Y(men_men_n450_));
  NO2        u0422(.A(men_men_n183_), .B(men_men_n145_), .Y(men_men_n451_));
  OAI210     u0423(.A0(men_men_n450_), .A1(men_men_n176_), .B0(men_men_n451_), .Y(men_men_n452_));
  INV        u0424(.A(men_men_n376_), .Y(men_men_n453_));
  NA3        u0425(.A(men_men_n453_), .B(men_men_n366_), .C(d), .Y(men_men_n454_));
  NO2        u0426(.A(men_men_n432_), .B(men_men_n49_), .Y(men_men_n455_));
  NAi21      u0427(.An(k), .B(j), .Y(men_men_n456_));
  NAi21      u0428(.An(e), .B(d), .Y(men_men_n457_));
  INV        u0429(.A(men_men_n457_), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n253_), .B(men_men_n214_), .Y(men_men_n459_));
  NA3        u0431(.A(men_men_n459_), .B(men_men_n458_), .C(men_men_n228_), .Y(men_men_n460_));
  NA3        u0432(.A(men_men_n460_), .B(men_men_n454_), .C(men_men_n452_), .Y(men_men_n461_));
  NO2        u0433(.A(men_men_n337_), .B(men_men_n214_), .Y(men_men_n462_));
  NA2        u0434(.A(men_men_n462_), .B(men_men_n458_), .Y(men_men_n463_));
  NOi31      u0435(.An(n), .B(m), .C(k), .Y(men_men_n464_));
  AOI220     u0436(.A0(men_men_n464_), .A1(men_men_n392_), .B0(men_men_n222_), .B1(men_men_n50_), .Y(men_men_n465_));
  NAi31      u0437(.An(g), .B(f), .C(c), .Y(men_men_n466_));
  OR3        u0438(.A(men_men_n466_), .B(men_men_n465_), .C(e), .Y(men_men_n467_));
  NA3        u0439(.A(men_men_n467_), .B(men_men_n463_), .C(men_men_n309_), .Y(men_men_n468_));
  NOi41      u0440(.An(men_men_n448_), .B(men_men_n468_), .C(men_men_n461_), .D(men_men_n265_), .Y(men_men_n469_));
  NOi32      u0441(.An(c), .Bn(a), .C(b), .Y(men_men_n470_));
  NA2        u0442(.A(men_men_n470_), .B(men_men_n114_), .Y(men_men_n471_));
  INV        u0443(.A(men_men_n274_), .Y(men_men_n472_));
  AN2        u0444(.A(e), .B(d), .Y(men_men_n473_));
  NA2        u0445(.A(men_men_n473_), .B(men_men_n472_), .Y(men_men_n474_));
  INV        u0446(.A(men_men_n145_), .Y(men_men_n475_));
  NO2        u0447(.A(men_men_n129_), .B(men_men_n41_), .Y(men_men_n476_));
  NO2        u0448(.A(men_men_n66_), .B(e), .Y(men_men_n477_));
  NOi31      u0449(.An(j), .B(k), .C(i), .Y(men_men_n478_));
  NOi21      u0450(.An(men_men_n164_), .B(men_men_n478_), .Y(men_men_n479_));
  NA4        u0451(.A(men_men_n323_), .B(men_men_n479_), .C(men_men_n261_), .D(men_men_n119_), .Y(men_men_n480_));
  AOI220     u0452(.A0(men_men_n480_), .A1(men_men_n477_), .B0(men_men_n476_), .B1(men_men_n475_), .Y(men_men_n481_));
  AOI210     u0453(.A0(men_men_n481_), .A1(men_men_n474_), .B0(men_men_n471_), .Y(men_men_n482_));
  INV        u0454(.A(men_men_n207_), .Y(men_men_n483_));
  NOi21      u0455(.An(a), .B(b), .Y(men_men_n484_));
  NA3        u0456(.A(e), .B(d), .C(c), .Y(men_men_n485_));
  NAi21      u0457(.An(men_men_n485_), .B(men_men_n484_), .Y(men_men_n486_));
  AOI210     u0458(.A0(men_men_n268_), .A1(men_men_n483_), .B0(men_men_n486_), .Y(men_men_n487_));
  NO4        u0459(.A(men_men_n189_), .B(men_men_n104_), .C(men_men_n56_), .D(b), .Y(men_men_n488_));
  NA2        u0460(.A(men_men_n387_), .B(men_men_n151_), .Y(men_men_n489_));
  OR2        u0461(.A(k), .B(j), .Y(men_men_n490_));
  NA2        u0462(.A(l), .B(k), .Y(men_men_n491_));
  NA3        u0463(.A(men_men_n491_), .B(men_men_n490_), .C(men_men_n222_), .Y(men_men_n492_));
  AOI210     u0464(.A0(men_men_n235_), .A1(men_men_n340_), .B0(men_men_n86_), .Y(men_men_n493_));
  NOi21      u0465(.An(men_men_n492_), .B(men_men_n493_), .Y(men_men_n494_));
  INV        u0466(.A(men_men_n279_), .Y(men_men_n495_));
  NA2        u0467(.A(men_men_n400_), .B(men_men_n114_), .Y(men_men_n496_));
  NO4        u0468(.A(men_men_n496_), .B(men_men_n97_), .C(men_men_n113_), .D(e), .Y(men_men_n497_));
  NO2        u0469(.A(men_men_n497_), .B(men_men_n495_), .Y(men_men_n498_));
  NA2        u0470(.A(men_men_n498_), .B(men_men_n489_), .Y(men_men_n499_));
  NO4        u0471(.A(men_men_n499_), .B(men_men_n488_), .C(men_men_n487_), .D(men_men_n482_), .Y(men_men_n500_));
  NA2        u0472(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n501_));
  NOi21      u0473(.An(d), .B(e), .Y(men_men_n502_));
  NAi31      u0474(.An(j), .B(l), .C(i), .Y(men_men_n503_));
  OAI210     u0475(.A0(men_men_n503_), .A1(men_men_n130_), .B0(men_men_n104_), .Y(men_men_n504_));
  NO3        u0476(.A(men_men_n401_), .B(men_men_n348_), .C(men_men_n203_), .Y(men_men_n505_));
  NO2        u0477(.A(men_men_n401_), .B(men_men_n376_), .Y(men_men_n506_));
  NO4        u0478(.A(men_men_n506_), .B(men_men_n505_), .C(men_men_n185_), .D(men_men_n306_), .Y(men_men_n507_));
  NA3        u0479(.A(men_men_n507_), .B(men_men_n501_), .C(men_men_n245_), .Y(men_men_n508_));
  OAI210     u0480(.A0(men_men_n127_), .A1(men_men_n126_), .B0(n), .Y(men_men_n509_));
  NO2        u0481(.A(men_men_n509_), .B(men_men_n129_), .Y(men_men_n510_));
  OR2        u0482(.A(men_men_n300_), .B(men_men_n247_), .Y(men_men_n511_));
  OA210      u0483(.A0(men_men_n511_), .A1(men_men_n510_), .B0(men_men_n194_), .Y(men_men_n512_));
  XO2        u0484(.A(i), .B(h), .Y(men_men_n513_));
  NA3        u0485(.A(men_men_n513_), .B(men_men_n158_), .C(n), .Y(men_men_n514_));
  NAi41      u0486(.An(men_men_n300_), .B(men_men_n514_), .C(men_men_n465_), .D(men_men_n389_), .Y(men_men_n515_));
  NOi32      u0487(.An(men_men_n515_), .Bn(men_men_n477_), .C(men_men_n270_), .Y(men_men_n516_));
  NAi31      u0488(.An(c), .B(f), .C(d), .Y(men_men_n517_));
  AOI210     u0489(.A0(men_men_n280_), .A1(men_men_n197_), .B0(men_men_n517_), .Y(men_men_n518_));
  NOi21      u0490(.An(men_men_n84_), .B(men_men_n518_), .Y(men_men_n519_));
  NA3        u0491(.A(men_men_n385_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n520_));
  NA2        u0492(.A(men_men_n229_), .B(men_men_n110_), .Y(men_men_n521_));
  AOI210     u0493(.A0(men_men_n521_), .A1(men_men_n181_), .B0(men_men_n517_), .Y(men_men_n522_));
  AOI210     u0494(.A0(men_men_n364_), .A1(men_men_n35_), .B0(men_men_n486_), .Y(men_men_n523_));
  NOi31      u0495(.An(men_men_n520_), .B(men_men_n523_), .C(men_men_n522_), .Y(men_men_n524_));
  AO220      u0496(.A0(men_men_n288_), .A1(men_men_n263_), .B0(men_men_n165_), .B1(men_men_n67_), .Y(men_men_n525_));
  NA3        u0497(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n526_));
  NO2        u0498(.A(men_men_n526_), .B(men_men_n443_), .Y(men_men_n527_));
  NO2        u0499(.A(men_men_n527_), .B(men_men_n296_), .Y(men_men_n528_));
  NAi41      u0500(.An(men_men_n525_), .B(men_men_n528_), .C(men_men_n524_), .D(men_men_n519_), .Y(men_men_n529_));
  NO4        u0501(.A(men_men_n529_), .B(men_men_n516_), .C(men_men_n512_), .D(men_men_n508_), .Y(men_men_n530_));
  NA4        u0502(.A(men_men_n530_), .B(men_men_n500_), .C(men_men_n469_), .D(men_men_n438_), .Y(men11));
  NO2        u0503(.A(men_men_n73_), .B(f), .Y(men_men_n532_));
  NA2        u0504(.A(j), .B(g), .Y(men_men_n533_));
  NAi31      u0505(.An(i), .B(m), .C(l), .Y(men_men_n534_));
  NA3        u0506(.A(m), .B(k), .C(j), .Y(men_men_n535_));
  OAI220     u0507(.A0(men_men_n535_), .A1(men_men_n129_), .B0(men_men_n534_), .B1(men_men_n533_), .Y(men_men_n536_));
  NA2        u0508(.A(men_men_n536_), .B(men_men_n532_), .Y(men_men_n537_));
  NOi32      u0509(.An(e), .Bn(b), .C(f), .Y(men_men_n538_));
  NA2        u0510(.A(men_men_n260_), .B(men_men_n114_), .Y(men_men_n539_));
  NA2        u0511(.A(men_men_n46_), .B(j), .Y(men_men_n540_));
  NAi31      u0512(.An(d), .B(e), .C(a), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n541_), .B(n), .Y(men_men_n542_));
  NAi41      u0514(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n543_));
  AN2        u0515(.A(men_men_n543_), .B(men_men_n375_), .Y(men_men_n544_));
  AOI210     u0516(.A0(men_men_n544_), .A1(men_men_n401_), .B0(men_men_n271_), .Y(men_men_n545_));
  NA2        u0517(.A(j), .B(i), .Y(men_men_n546_));
  NAi31      u0518(.An(n), .B(m), .C(k), .Y(men_men_n547_));
  NO3        u0519(.A(men_men_n547_), .B(men_men_n546_), .C(men_men_n113_), .Y(men_men_n548_));
  NO4        u0520(.A(n), .B(d), .C(men_men_n116_), .D(a), .Y(men_men_n549_));
  OR2        u0521(.A(n), .B(c), .Y(men_men_n550_));
  NO2        u0522(.A(men_men_n550_), .B(men_men_n147_), .Y(men_men_n551_));
  NO2        u0523(.A(men_men_n551_), .B(men_men_n549_), .Y(men_men_n552_));
  NOi32      u0524(.An(g), .Bn(f), .C(i), .Y(men_men_n553_));
  AOI220     u0525(.A0(men_men_n553_), .A1(men_men_n101_), .B0(men_men_n536_), .B1(f), .Y(men_men_n554_));
  NO2        u0526(.A(men_men_n274_), .B(men_men_n49_), .Y(men_men_n555_));
  NO2        u0527(.A(men_men_n554_), .B(men_men_n552_), .Y(men_men_n556_));
  AOI210     u0528(.A0(men_men_n548_), .A1(men_men_n545_), .B0(men_men_n556_), .Y(men_men_n557_));
  NA2        u0529(.A(men_men_n138_), .B(men_men_n34_), .Y(men_men_n558_));
  OAI220     u0530(.A0(men_men_n558_), .A1(m), .B0(men_men_n540_), .B1(men_men_n235_), .Y(men_men_n559_));
  NOi41      u0531(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n560_));
  NAi32      u0532(.An(e), .Bn(b), .C(c), .Y(men_men_n561_));
  OR2        u0533(.A(men_men_n561_), .B(men_men_n86_), .Y(men_men_n562_));
  AN2        u0534(.A(men_men_n341_), .B(men_men_n320_), .Y(men_men_n563_));
  NA2        u0535(.A(men_men_n563_), .B(men_men_n562_), .Y(men_men_n564_));
  OA210      u0536(.A0(men_men_n564_), .A1(men_men_n560_), .B0(men_men_n559_), .Y(men_men_n565_));
  OAI220     u0537(.A0(men_men_n403_), .A1(men_men_n402_), .B0(men_men_n534_), .B1(men_men_n533_), .Y(men_men_n566_));
  NAi31      u0538(.An(d), .B(c), .C(a), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n567_), .B(n), .Y(men_men_n568_));
  NA3        u0540(.A(men_men_n568_), .B(men_men_n566_), .C(e), .Y(men_men_n569_));
  NO3        u0541(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n215_), .Y(men_men_n570_));
  NO2        u0542(.A(men_men_n232_), .B(men_men_n111_), .Y(men_men_n571_));
  OAI210     u0543(.A0(men_men_n570_), .A1(men_men_n404_), .B0(men_men_n571_), .Y(men_men_n572_));
  NA2        u0544(.A(men_men_n572_), .B(men_men_n569_), .Y(men_men_n573_));
  INV        u0545(.A(men_men_n433_), .Y(men_men_n574_));
  NA2        u0546(.A(men_men_n566_), .B(f), .Y(men_men_n575_));
  NAi32      u0547(.An(d), .Bn(a), .C(b), .Y(men_men_n576_));
  NO2        u0548(.A(men_men_n576_), .B(men_men_n49_), .Y(men_men_n577_));
  NA2        u0549(.A(h), .B(f), .Y(men_men_n578_));
  NO2        u0550(.A(men_men_n578_), .B(men_men_n97_), .Y(men_men_n579_));
  NO3        u0551(.A(men_men_n177_), .B(men_men_n174_), .C(g), .Y(men_men_n580_));
  AOI220     u0552(.A0(men_men_n580_), .A1(men_men_n58_), .B0(men_men_n579_), .B1(men_men_n577_), .Y(men_men_n581_));
  OAI210     u0553(.A0(men_men_n575_), .A1(men_men_n574_), .B0(men_men_n581_), .Y(men_men_n582_));
  AN3        u0554(.A(j), .B(h), .C(g), .Y(men_men_n583_));
  NO2        u0555(.A(men_men_n144_), .B(c), .Y(men_men_n584_));
  NA3        u0556(.A(men_men_n584_), .B(men_men_n583_), .C(men_men_n464_), .Y(men_men_n585_));
  NA3        u0557(.A(f), .B(d), .C(b), .Y(men_men_n586_));
  NO4        u0558(.A(men_men_n586_), .B(men_men_n177_), .C(men_men_n174_), .D(g), .Y(men_men_n587_));
  NAi21      u0559(.An(men_men_n587_), .B(men_men_n585_), .Y(men_men_n588_));
  NO4        u0560(.A(men_men_n588_), .B(men_men_n582_), .C(men_men_n573_), .D(men_men_n565_), .Y(men_men_n589_));
  AN3        u0561(.A(men_men_n589_), .B(men_men_n557_), .C(men_men_n537_), .Y(men_men_n590_));
  INV        u0562(.A(k), .Y(men_men_n591_));
  NA3        u0563(.A(l), .B(men_men_n591_), .C(i), .Y(men_men_n592_));
  INV        u0564(.A(men_men_n592_), .Y(men_men_n593_));
  NA4        u0565(.A(men_men_n400_), .B(men_men_n423_), .C(men_men_n182_), .D(men_men_n114_), .Y(men_men_n594_));
  NAi32      u0566(.An(h), .Bn(f), .C(g), .Y(men_men_n595_));
  NAi41      u0567(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n596_));
  OAI210     u0568(.A0(men_men_n541_), .A1(n), .B0(men_men_n596_), .Y(men_men_n597_));
  NAi31      u0569(.An(h), .B(g), .C(f), .Y(men_men_n598_));
  NA4        u0570(.A(men_men_n423_), .B(men_men_n121_), .C(men_men_n114_), .D(e), .Y(men_men_n599_));
  NO3        u0571(.A(men_men_n595_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n600_));
  NAi31      u0572(.An(men_men_n600_), .B(men_men_n599_), .C(men_men_n594_), .Y(men_men_n601_));
  NAi31      u0573(.An(f), .B(h), .C(g), .Y(men_men_n602_));
  NOi32      u0574(.An(b), .Bn(a), .C(c), .Y(men_men_n603_));
  NOi41      u0575(.An(men_men_n603_), .B(men_men_n357_), .C(men_men_n69_), .D(men_men_n117_), .Y(men_men_n604_));
  NOi32      u0576(.An(d), .Bn(a), .C(e), .Y(men_men_n605_));
  NA2        u0577(.A(men_men_n605_), .B(men_men_n114_), .Y(men_men_n606_));
  NO2        u0578(.A(n), .B(c), .Y(men_men_n607_));
  NA3        u0579(.A(men_men_n607_), .B(men_men_n29_), .C(m), .Y(men_men_n608_));
  NOi32      u0580(.An(e), .Bn(a), .C(d), .Y(men_men_n609_));
  AOI210     u0581(.A0(men_men_n29_), .A1(d), .B0(men_men_n609_), .Y(men_men_n610_));
  AOI210     u0582(.A0(men_men_n601_), .A1(men_men_n593_), .B0(men_men_n604_), .Y(men_men_n611_));
  NO3        u0583(.A(men_men_n318_), .B(men_men_n61_), .C(n), .Y(men_men_n612_));
  NA3        u0584(.A(men_men_n517_), .B(men_men_n172_), .C(men_men_n171_), .Y(men_men_n613_));
  NA2        u0585(.A(men_men_n466_), .B(men_men_n232_), .Y(men_men_n614_));
  OR2        u0586(.A(men_men_n614_), .B(men_men_n613_), .Y(men_men_n615_));
  NA2        u0587(.A(men_men_n76_), .B(men_men_n114_), .Y(men_men_n616_));
  NO2        u0588(.A(men_men_n616_), .B(men_men_n45_), .Y(men_men_n617_));
  AOI220     u0589(.A0(men_men_n617_), .A1(men_men_n545_), .B0(men_men_n615_), .B1(men_men_n612_), .Y(men_men_n618_));
  NO2        u0590(.A(men_men_n618_), .B(men_men_n89_), .Y(men_men_n619_));
  NA3        u0591(.A(men_men_n560_), .B(men_men_n343_), .C(men_men_n46_), .Y(men_men_n620_));
  NOi32      u0592(.An(e), .Bn(c), .C(f), .Y(men_men_n621_));
  NOi21      u0593(.An(f), .B(g), .Y(men_men_n622_));
  NO2        u0594(.A(men_men_n622_), .B(men_men_n212_), .Y(men_men_n623_));
  AOI220     u0595(.A0(men_men_n623_), .A1(men_men_n397_), .B0(men_men_n621_), .B1(men_men_n176_), .Y(men_men_n624_));
  NA3        u0596(.A(men_men_n624_), .B(men_men_n620_), .C(men_men_n179_), .Y(men_men_n625_));
  AOI210     u0597(.A0(men_men_n544_), .A1(men_men_n401_), .B0(men_men_n301_), .Y(men_men_n626_));
  NA2        u0598(.A(men_men_n626_), .B(men_men_n264_), .Y(men_men_n627_));
  NOi21      u0599(.An(j), .B(l), .Y(men_men_n628_));
  NAi21      u0600(.An(k), .B(h), .Y(men_men_n629_));
  NO2        u0601(.A(men_men_n629_), .B(men_men_n262_), .Y(men_men_n630_));
  NA2        u0602(.A(men_men_n630_), .B(men_men_n628_), .Y(men_men_n631_));
  NOi31      u0603(.An(m), .B(n), .C(k), .Y(men_men_n632_));
  NA2        u0604(.A(men_men_n628_), .B(men_men_n632_), .Y(men_men_n633_));
  AOI210     u0605(.A0(men_men_n401_), .A1(men_men_n375_), .B0(men_men_n301_), .Y(men_men_n634_));
  NAi21      u0606(.An(men_men_n633_), .B(men_men_n634_), .Y(men_men_n635_));
  NA2        u0607(.A(men_men_n635_), .B(men_men_n627_), .Y(men_men_n636_));
  NA2        u0608(.A(men_men_n110_), .B(men_men_n36_), .Y(men_men_n637_));
  NO2        u0609(.A(k), .B(men_men_n215_), .Y(men_men_n638_));
  INV        u0610(.A(men_men_n366_), .Y(men_men_n639_));
  NO2        u0611(.A(men_men_n639_), .B(n), .Y(men_men_n640_));
  NAi31      u0612(.An(men_men_n637_), .B(men_men_n640_), .C(men_men_n638_), .Y(men_men_n641_));
  NO2        u0613(.A(men_men_n540_), .B(men_men_n177_), .Y(men_men_n642_));
  NA3        u0614(.A(men_men_n561_), .B(men_men_n270_), .C(men_men_n142_), .Y(men_men_n643_));
  NA2        u0615(.A(men_men_n513_), .B(men_men_n158_), .Y(men_men_n644_));
  NO3        u0616(.A(men_men_n398_), .B(men_men_n644_), .C(men_men_n89_), .Y(men_men_n645_));
  AOI210     u0617(.A0(men_men_n643_), .A1(men_men_n642_), .B0(men_men_n645_), .Y(men_men_n646_));
  AN3        u0618(.A(f), .B(d), .C(b), .Y(men_men_n647_));
  OAI210     u0619(.A0(men_men_n647_), .A1(men_men_n128_), .B0(n), .Y(men_men_n648_));
  NA3        u0620(.A(men_men_n513_), .B(men_men_n158_), .C(men_men_n215_), .Y(men_men_n649_));
  AOI210     u0621(.A0(men_men_n648_), .A1(men_men_n234_), .B0(men_men_n649_), .Y(men_men_n650_));
  NAi31      u0622(.An(m), .B(n), .C(k), .Y(men_men_n651_));
  OR2        u0623(.A(men_men_n133_), .B(men_men_n61_), .Y(men_men_n652_));
  OAI210     u0624(.A0(men_men_n652_), .A1(men_men_n651_), .B0(men_men_n251_), .Y(men_men_n653_));
  OAI210     u0625(.A0(men_men_n653_), .A1(men_men_n650_), .B0(j), .Y(men_men_n654_));
  NA3        u0626(.A(men_men_n654_), .B(men_men_n646_), .C(men_men_n641_), .Y(men_men_n655_));
  NO4        u0627(.A(men_men_n655_), .B(men_men_n636_), .C(men_men_n625_), .D(men_men_n619_), .Y(men_men_n656_));
  NA2        u0628(.A(men_men_n385_), .B(men_men_n161_), .Y(men_men_n657_));
  NAi31      u0629(.An(g), .B(h), .C(f), .Y(men_men_n658_));
  OR3        u0630(.A(men_men_n658_), .B(men_men_n276_), .C(n), .Y(men_men_n659_));
  OA210      u0631(.A0(men_men_n541_), .A1(n), .B0(men_men_n596_), .Y(men_men_n660_));
  NA3        u0632(.A(men_men_n421_), .B(men_men_n121_), .C(men_men_n86_), .Y(men_men_n661_));
  OAI210     u0633(.A0(men_men_n660_), .A1(men_men_n93_), .B0(men_men_n661_), .Y(men_men_n662_));
  NOi21      u0634(.An(men_men_n659_), .B(men_men_n662_), .Y(men_men_n663_));
  AOI210     u0635(.A0(men_men_n663_), .A1(men_men_n657_), .B0(men_men_n535_), .Y(men_men_n664_));
  NO3        u0636(.A(g), .B(men_men_n214_), .C(men_men_n56_), .Y(men_men_n665_));
  NAi21      u0637(.An(h), .B(j), .Y(men_men_n666_));
  NO2        u0638(.A(men_men_n521_), .B(men_men_n89_), .Y(men_men_n667_));
  OAI210     u0639(.A0(men_men_n667_), .A1(men_men_n397_), .B0(men_men_n665_), .Y(men_men_n668_));
  OR2        u0640(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n669_));
  NA2        u0641(.A(men_men_n603_), .B(men_men_n345_), .Y(men_men_n670_));
  OA220      u0642(.A0(men_men_n633_), .A1(men_men_n670_), .B0(men_men_n631_), .B1(men_men_n669_), .Y(men_men_n671_));
  NA3        u0643(.A(men_men_n532_), .B(men_men_n101_), .C(men_men_n100_), .Y(men_men_n672_));
  AN2        u0644(.A(h), .B(f), .Y(men_men_n673_));
  NA2        u0645(.A(men_men_n673_), .B(men_men_n37_), .Y(men_men_n674_));
  NA2        u0646(.A(men_men_n101_), .B(men_men_n46_), .Y(men_men_n675_));
  OAI220     u0647(.A0(men_men_n675_), .A1(men_men_n334_), .B0(men_men_n674_), .B1(men_men_n471_), .Y(men_men_n676_));
  AOI210     u0648(.A0(men_men_n576_), .A1(men_men_n432_), .B0(men_men_n49_), .Y(men_men_n677_));
  OAI220     u0649(.A0(men_men_n598_), .A1(men_men_n592_), .B0(men_men_n327_), .B1(men_men_n533_), .Y(men_men_n678_));
  AOI210     u0650(.A0(men_men_n678_), .A1(men_men_n677_), .B0(men_men_n676_), .Y(men_men_n679_));
  NA4        u0651(.A(men_men_n679_), .B(men_men_n672_), .C(men_men_n671_), .D(men_men_n668_), .Y(men_men_n680_));
  NO2        u0652(.A(men_men_n252_), .B(f), .Y(men_men_n681_));
  NO2        u0653(.A(men_men_n622_), .B(men_men_n61_), .Y(men_men_n682_));
  NO3        u0654(.A(men_men_n682_), .B(men_men_n681_), .C(men_men_n34_), .Y(men_men_n683_));
  NA2        u0655(.A(men_men_n330_), .B(men_men_n138_), .Y(men_men_n684_));
  NA2        u0656(.A(men_men_n130_), .B(men_men_n49_), .Y(men_men_n685_));
  AOI220     u0657(.A0(men_men_n685_), .A1(men_men_n538_), .B0(men_men_n366_), .B1(men_men_n114_), .Y(men_men_n686_));
  OA220      u0658(.A0(men_men_n686_), .A1(men_men_n558_), .B0(men_men_n364_), .B1(men_men_n112_), .Y(men_men_n687_));
  OAI210     u0659(.A0(men_men_n684_), .A1(men_men_n683_), .B0(men_men_n687_), .Y(men_men_n688_));
  NO3        u0660(.A(men_men_n408_), .B(men_men_n194_), .C(men_men_n193_), .Y(men_men_n689_));
  NA2        u0661(.A(men_men_n689_), .B(men_men_n232_), .Y(men_men_n690_));
  NA3        u0662(.A(men_men_n690_), .B(men_men_n254_), .C(j), .Y(men_men_n691_));
  NO3        u0663(.A(men_men_n466_), .B(men_men_n174_), .C(i), .Y(men_men_n692_));
  NA2        u0664(.A(men_men_n470_), .B(men_men_n86_), .Y(men_men_n693_));
  NO4        u0665(.A(men_men_n535_), .B(men_men_n693_), .C(men_men_n129_), .D(men_men_n214_), .Y(men_men_n694_));
  INV        u0666(.A(men_men_n694_), .Y(men_men_n695_));
  NA4        u0667(.A(men_men_n695_), .B(men_men_n691_), .C(men_men_n520_), .D(men_men_n406_), .Y(men_men_n696_));
  NO4        u0668(.A(men_men_n696_), .B(men_men_n688_), .C(men_men_n680_), .D(men_men_n664_), .Y(men_men_n697_));
  NA4        u0669(.A(men_men_n697_), .B(men_men_n656_), .C(men_men_n611_), .D(men_men_n590_), .Y(men08));
  NO2        u0670(.A(k), .B(h), .Y(men_men_n699_));
  AO210      u0671(.A0(men_men_n252_), .A1(men_men_n456_), .B0(men_men_n699_), .Y(men_men_n700_));
  NO2        u0672(.A(men_men_n700_), .B(men_men_n299_), .Y(men_men_n701_));
  NA2        u0673(.A(men_men_n621_), .B(men_men_n86_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n702_), .B(men_men_n466_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n703_), .B(men_men_n701_), .Y(men_men_n704_));
  NA2        u0676(.A(men_men_n86_), .B(men_men_n111_), .Y(men_men_n705_));
  NO2        u0677(.A(men_men_n705_), .B(men_men_n57_), .Y(men_men_n706_));
  NA2        u0678(.A(men_men_n586_), .B(men_men_n234_), .Y(men_men_n707_));
  NA2        u0679(.A(men_men_n707_), .B(men_men_n351_), .Y(men_men_n708_));
  AOI210     u0680(.A0(men_men_n586_), .A1(men_men_n154_), .B0(men_men_n86_), .Y(men_men_n709_));
  NA4        u0681(.A(men_men_n217_), .B(men_men_n138_), .C(men_men_n45_), .D(h), .Y(men_men_n710_));
  AN2        u0682(.A(l), .B(k), .Y(men_men_n711_));
  NA4        u0683(.A(men_men_n711_), .B(men_men_n110_), .C(men_men_n75_), .D(men_men_n215_), .Y(men_men_n712_));
  OAI210     u0684(.A0(men_men_n710_), .A1(g), .B0(men_men_n712_), .Y(men_men_n713_));
  NA2        u0685(.A(men_men_n713_), .B(men_men_n709_), .Y(men_men_n714_));
  NA4        u0686(.A(men_men_n714_), .B(men_men_n708_), .C(men_men_n704_), .D(men_men_n353_), .Y(men_men_n715_));
  NO4        u0687(.A(men_men_n174_), .B(men_men_n396_), .C(men_men_n113_), .D(g), .Y(men_men_n716_));
  AOI210     u0688(.A0(men_men_n716_), .A1(men_men_n707_), .B0(men_men_n527_), .Y(men_men_n717_));
  NA2        u0689(.A(men_men_n623_), .B(men_men_n350_), .Y(men_men_n718_));
  NA2        u0690(.A(men_men_n718_), .B(men_men_n717_), .Y(men_men_n719_));
  NO2        u0691(.A(men_men_n544_), .B(men_men_n35_), .Y(men_men_n720_));
  OAI210     u0692(.A0(men_men_n561_), .A1(men_men_n47_), .B0(men_men_n652_), .Y(men_men_n721_));
  NO2        u0693(.A(men_men_n491_), .B(men_men_n130_), .Y(men_men_n722_));
  AOI210     u0694(.A0(men_men_n722_), .A1(men_men_n721_), .B0(men_men_n720_), .Y(men_men_n723_));
  NO3        u0695(.A(men_men_n318_), .B(men_men_n129_), .C(men_men_n41_), .Y(men_men_n724_));
  NAi21      u0696(.An(men_men_n724_), .B(men_men_n712_), .Y(men_men_n725_));
  NA2        u0697(.A(men_men_n700_), .B(men_men_n134_), .Y(men_men_n726_));
  AOI220     u0698(.A0(men_men_n726_), .A1(men_men_n407_), .B0(men_men_n725_), .B1(men_men_n78_), .Y(men_men_n727_));
  OAI210     u0699(.A0(men_men_n723_), .A1(men_men_n89_), .B0(men_men_n727_), .Y(men_men_n728_));
  NA2        u0700(.A(men_men_n366_), .B(men_men_n43_), .Y(men_men_n729_));
  NA3        u0701(.A(men_men_n690_), .B(men_men_n336_), .C(men_men_n388_), .Y(men_men_n730_));
  NA2        u0702(.A(men_men_n711_), .B(men_men_n222_), .Y(men_men_n731_));
  NO2        u0703(.A(men_men_n731_), .B(men_men_n329_), .Y(men_men_n732_));
  AOI210     u0704(.A0(men_men_n732_), .A1(men_men_n681_), .B0(men_men_n497_), .Y(men_men_n733_));
  NA3        u0705(.A(m), .B(l), .C(k), .Y(men_men_n734_));
  AOI210     u0706(.A0(men_men_n661_), .A1(men_men_n659_), .B0(men_men_n734_), .Y(men_men_n735_));
  NO2        u0707(.A(men_men_n543_), .B(men_men_n271_), .Y(men_men_n736_));
  NOi21      u0708(.An(men_men_n736_), .B(men_men_n539_), .Y(men_men_n737_));
  NA4        u0709(.A(men_men_n114_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n738_));
  NA3        u0710(.A(men_men_n121_), .B(men_men_n416_), .C(i), .Y(men_men_n739_));
  NO2        u0711(.A(men_men_n739_), .B(men_men_n738_), .Y(men_men_n740_));
  NO3        u0712(.A(men_men_n740_), .B(men_men_n737_), .C(men_men_n735_), .Y(men_men_n741_));
  NA4        u0713(.A(men_men_n741_), .B(men_men_n733_), .C(men_men_n730_), .D(men_men_n729_), .Y(men_men_n742_));
  NO4        u0714(.A(men_men_n742_), .B(men_men_n728_), .C(men_men_n719_), .D(men_men_n715_), .Y(men_men_n743_));
  NA2        u0715(.A(men_men_n623_), .B(men_men_n397_), .Y(men_men_n744_));
  NO3        u0716(.A(men_men_n401_), .B(men_men_n533_), .C(h), .Y(men_men_n745_));
  AOI210     u0717(.A0(men_men_n745_), .A1(men_men_n114_), .B0(men_men_n506_), .Y(men_men_n746_));
  NA3        u0718(.A(men_men_n746_), .B(men_men_n744_), .C(men_men_n251_), .Y(men_men_n747_));
  NA2        u0719(.A(men_men_n711_), .B(men_men_n75_), .Y(men_men_n748_));
  NO4        u0720(.A(men_men_n689_), .B(men_men_n174_), .C(n), .D(i), .Y(men_men_n749_));
  NOi21      u0721(.An(h), .B(j), .Y(men_men_n750_));
  NA2        u0722(.A(men_men_n750_), .B(f), .Y(men_men_n751_));
  NO2        u0723(.A(men_men_n749_), .B(men_men_n692_), .Y(men_men_n752_));
  OAI220     u0724(.A0(men_men_n752_), .A1(men_men_n748_), .B0(men_men_n599_), .B1(men_men_n62_), .Y(men_men_n753_));
  AOI210     u0725(.A0(men_men_n747_), .A1(l), .B0(men_men_n753_), .Y(men_men_n754_));
  NO2        u0726(.A(j), .B(i), .Y(men_men_n755_));
  NA2        u0727(.A(men_men_n755_), .B(men_men_n33_), .Y(men_men_n756_));
  NA2        u0728(.A(men_men_n426_), .B(men_men_n121_), .Y(men_men_n757_));
  OR2        u0729(.A(men_men_n757_), .B(men_men_n756_), .Y(men_men_n758_));
  NO3        u0730(.A(men_men_n149_), .B(men_men_n49_), .C(men_men_n111_), .Y(men_men_n759_));
  NO3        u0731(.A(men_men_n550_), .B(men_men_n147_), .C(men_men_n75_), .Y(men_men_n760_));
  NO3        u0732(.A(men_men_n491_), .B(men_men_n444_), .C(j), .Y(men_men_n761_));
  NA2        u0733(.A(k), .B(j), .Y(men_men_n762_));
  NO3        u0734(.A(men_men_n299_), .B(men_men_n762_), .C(men_men_n40_), .Y(men_men_n763_));
  AOI210     u0735(.A0(men_men_n538_), .A1(n), .B0(men_men_n560_), .Y(men_men_n764_));
  NA2        u0736(.A(men_men_n764_), .B(men_men_n563_), .Y(men_men_n765_));
  AN3        u0737(.A(men_men_n765_), .B(men_men_n763_), .C(men_men_n100_), .Y(men_men_n766_));
  NA2        u0738(.A(men_men_n614_), .B(men_men_n308_), .Y(men_men_n767_));
  NAi31      u0739(.An(men_men_n610_), .B(men_men_n95_), .C(men_men_n86_), .Y(men_men_n768_));
  NA2        u0740(.A(men_men_n768_), .B(men_men_n767_), .Y(men_men_n769_));
  NO2        u0741(.A(men_men_n299_), .B(men_men_n134_), .Y(men_men_n770_));
  AOI220     u0742(.A0(men_men_n770_), .A1(men_men_n623_), .B0(men_men_n724_), .B1(men_men_n709_), .Y(men_men_n771_));
  NO2        u0743(.A(men_men_n734_), .B(men_men_n93_), .Y(men_men_n772_));
  NA2        u0744(.A(men_men_n772_), .B(men_men_n597_), .Y(men_men_n773_));
  NO2        u0745(.A(men_men_n598_), .B(men_men_n117_), .Y(men_men_n774_));
  OAI210     u0746(.A0(men_men_n774_), .A1(men_men_n761_), .B0(men_men_n677_), .Y(men_men_n775_));
  NA3        u0747(.A(men_men_n775_), .B(men_men_n773_), .C(men_men_n771_), .Y(men_men_n776_));
  OR3        u0748(.A(men_men_n776_), .B(men_men_n769_), .C(men_men_n766_), .Y(men_men_n777_));
  NA3        u0749(.A(men_men_n764_), .B(men_men_n563_), .C(men_men_n562_), .Y(men_men_n778_));
  NA4        u0750(.A(men_men_n778_), .B(men_men_n217_), .C(men_men_n456_), .D(men_men_n34_), .Y(men_men_n779_));
  NO4        u0751(.A(men_men_n491_), .B(men_men_n439_), .C(j), .D(f), .Y(men_men_n780_));
  OAI220     u0752(.A0(men_men_n710_), .A1(men_men_n702_), .B0(men_men_n334_), .B1(men_men_n38_), .Y(men_men_n781_));
  AOI210     u0753(.A0(men_men_n780_), .A1(men_men_n258_), .B0(men_men_n781_), .Y(men_men_n782_));
  NA3        u0754(.A(men_men_n553_), .B(men_men_n292_), .C(h), .Y(men_men_n783_));
  NOi21      u0755(.An(men_men_n677_), .B(men_men_n783_), .Y(men_men_n784_));
  NO2        u0756(.A(men_men_n94_), .B(men_men_n47_), .Y(men_men_n785_));
  NO2        u0757(.A(men_men_n783_), .B(men_men_n608_), .Y(men_men_n786_));
  AOI210     u0758(.A0(men_men_n785_), .A1(men_men_n640_), .B0(men_men_n786_), .Y(men_men_n787_));
  NAi41      u0759(.An(men_men_n784_), .B(men_men_n787_), .C(men_men_n782_), .D(men_men_n779_), .Y(men_men_n788_));
  BUFFER     u0760(.A(men_men_n772_), .Y(men_men_n789_));
  NA2        u0761(.A(men_men_n789_), .B(men_men_n240_), .Y(men_men_n790_));
  NO2        u0762(.A(men_men_n660_), .B(men_men_n75_), .Y(men_men_n791_));
  AOI210     u0763(.A0(men_men_n780_), .A1(men_men_n791_), .B0(men_men_n338_), .Y(men_men_n792_));
  OAI210     u0764(.A0(men_men_n734_), .A1(men_men_n658_), .B0(men_men_n526_), .Y(men_men_n793_));
  NA3        u0765(.A(men_men_n250_), .B(men_men_n59_), .C(b), .Y(men_men_n794_));
  AOI220     u0766(.A0(men_men_n607_), .A1(men_men_n29_), .B0(men_men_n470_), .B1(men_men_n86_), .Y(men_men_n795_));
  NA2        u0767(.A(men_men_n795_), .B(men_men_n794_), .Y(men_men_n796_));
  NO2        u0768(.A(men_men_n783_), .B(men_men_n496_), .Y(men_men_n797_));
  AOI210     u0769(.A0(men_men_n796_), .A1(men_men_n793_), .B0(men_men_n797_), .Y(men_men_n798_));
  NA3        u0770(.A(men_men_n798_), .B(men_men_n792_), .C(men_men_n790_), .Y(men_men_n799_));
  NOi41      u0771(.An(men_men_n758_), .B(men_men_n799_), .C(men_men_n788_), .D(men_men_n777_), .Y(men_men_n800_));
  OR3        u0772(.A(men_men_n710_), .B(men_men_n234_), .C(g), .Y(men_men_n801_));
  NO3        u0773(.A(men_men_n344_), .B(men_men_n301_), .C(men_men_n113_), .Y(men_men_n802_));
  NA2        u0774(.A(men_men_n802_), .B(men_men_n765_), .Y(men_men_n803_));
  NA2        u0775(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n804_));
  NO3        u0776(.A(men_men_n804_), .B(men_men_n756_), .C(men_men_n276_), .Y(men_men_n805_));
  NO3        u0777(.A(men_men_n533_), .B(men_men_n96_), .C(h), .Y(men_men_n806_));
  AOI210     u0778(.A0(men_men_n806_), .A1(men_men_n706_), .B0(men_men_n805_), .Y(men_men_n807_));
  NA4        u0779(.A(men_men_n807_), .B(men_men_n803_), .C(men_men_n801_), .D(men_men_n409_), .Y(men_men_n808_));
  OR2        u0780(.A(men_men_n658_), .B(men_men_n94_), .Y(men_men_n809_));
  NOi31      u0781(.An(b), .B(d), .C(a), .Y(men_men_n810_));
  NO2        u0782(.A(men_men_n810_), .B(men_men_n605_), .Y(men_men_n811_));
  NO2        u0783(.A(men_men_n811_), .B(n), .Y(men_men_n812_));
  NOi21      u0784(.An(men_men_n795_), .B(men_men_n812_), .Y(men_men_n813_));
  NO2        u0785(.A(men_men_n813_), .B(men_men_n809_), .Y(men_men_n814_));
  NO2        u0786(.A(men_men_n561_), .B(men_men_n86_), .Y(men_men_n815_));
  NA2        u0787(.A(men_men_n802_), .B(men_men_n815_), .Y(men_men_n816_));
  OAI210     u0788(.A0(men_men_n710_), .A1(men_men_n398_), .B0(men_men_n816_), .Y(men_men_n817_));
  NO2        u0789(.A(men_men_n689_), .B(n), .Y(men_men_n818_));
  AOI220     u0790(.A0(men_men_n770_), .A1(men_men_n665_), .B0(men_men_n818_), .B1(men_men_n701_), .Y(men_men_n819_));
  NA2        u0791(.A(men_men_n121_), .B(men_men_n86_), .Y(men_men_n820_));
  AOI210     u0792(.A0(men_men_n430_), .A1(men_men_n422_), .B0(men_men_n820_), .Y(men_men_n821_));
  NA2        u0793(.A(men_men_n732_), .B(men_men_n34_), .Y(men_men_n822_));
  NAi21      u0794(.An(men_men_n738_), .B(men_men_n440_), .Y(men_men_n823_));
  NO2        u0795(.A(men_men_n271_), .B(i), .Y(men_men_n824_));
  NA2        u0796(.A(men_men_n716_), .B(men_men_n352_), .Y(men_men_n825_));
  NA2        u0797(.A(men_men_n600_), .B(men_men_n367_), .Y(men_men_n826_));
  AN3        u0798(.A(men_men_n826_), .B(men_men_n825_), .C(men_men_n823_), .Y(men_men_n827_));
  NAi41      u0799(.An(men_men_n821_), .B(men_men_n827_), .C(men_men_n822_), .D(men_men_n819_), .Y(men_men_n828_));
  NO4        u0800(.A(men_men_n828_), .B(men_men_n817_), .C(men_men_n814_), .D(men_men_n808_), .Y(men_men_n829_));
  NA4        u0801(.A(men_men_n829_), .B(men_men_n800_), .C(men_men_n754_), .D(men_men_n743_), .Y(men09));
  INV        u0802(.A(men_men_n122_), .Y(men_men_n831_));
  NA2        u0803(.A(f), .B(e), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n227_), .B(men_men_n113_), .Y(men_men_n833_));
  NA2        u0805(.A(men_men_n833_), .B(g), .Y(men_men_n834_));
  NA4        u0806(.A(men_men_n311_), .B(men_men_n479_), .C(men_men_n261_), .D(men_men_n119_), .Y(men_men_n835_));
  AOI210     u0807(.A0(men_men_n835_), .A1(g), .B0(men_men_n476_), .Y(men_men_n836_));
  AOI210     u0808(.A0(men_men_n836_), .A1(men_men_n834_), .B0(men_men_n832_), .Y(men_men_n837_));
  NA2        u0809(.A(men_men_n450_), .B(e), .Y(men_men_n838_));
  NO2        u0810(.A(men_men_n838_), .B(men_men_n517_), .Y(men_men_n839_));
  AOI210     u0811(.A0(men_men_n837_), .A1(men_men_n831_), .B0(men_men_n839_), .Y(men_men_n840_));
  NO2        u0812(.A(men_men_n206_), .B(men_men_n214_), .Y(men_men_n841_));
  NA3        u0813(.A(m), .B(l), .C(i), .Y(men_men_n842_));
  OAI220     u0814(.A0(men_men_n598_), .A1(men_men_n842_), .B0(men_men_n357_), .B1(men_men_n534_), .Y(men_men_n843_));
  NA4        u0815(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(f), .Y(men_men_n844_));
  NAi31      u0816(.An(men_men_n843_), .B(men_men_n844_), .C(men_men_n445_), .Y(men_men_n845_));
  OR2        u0817(.A(men_men_n845_), .B(men_men_n841_), .Y(men_men_n846_));
  NA3        u0818(.A(men_men_n809_), .B(men_men_n575_), .C(men_men_n526_), .Y(men_men_n847_));
  OA210      u0819(.A0(men_men_n847_), .A1(men_men_n846_), .B0(men_men_n812_), .Y(men_men_n848_));
  INV        u0820(.A(men_men_n341_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n850_));
  NOi31      u0822(.An(k), .B(m), .C(l), .Y(men_men_n851_));
  NO2        u0823(.A(men_men_n343_), .B(men_men_n851_), .Y(men_men_n852_));
  AOI210     u0824(.A0(men_men_n852_), .A1(men_men_n850_), .B0(men_men_n602_), .Y(men_men_n853_));
  NA2        u0825(.A(men_men_n794_), .B(men_men_n334_), .Y(men_men_n854_));
  NA2        u0826(.A(men_men_n345_), .B(men_men_n347_), .Y(men_men_n855_));
  OAI210     u0827(.A0(men_men_n206_), .A1(men_men_n214_), .B0(men_men_n855_), .Y(men_men_n856_));
  AOI220     u0828(.A0(men_men_n856_), .A1(men_men_n854_), .B0(men_men_n853_), .B1(men_men_n849_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n168_), .B(men_men_n115_), .Y(men_men_n858_));
  NA3        u0830(.A(men_men_n858_), .B(men_men_n700_), .C(men_men_n134_), .Y(men_men_n859_));
  NA3        u0831(.A(men_men_n859_), .B(men_men_n191_), .C(men_men_n31_), .Y(men_men_n860_));
  NA4        u0832(.A(men_men_n860_), .B(men_men_n857_), .C(men_men_n624_), .D(men_men_n84_), .Y(men_men_n861_));
  NO2        u0833(.A(men_men_n595_), .B(men_men_n503_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n862_), .B(men_men_n191_), .Y(men_men_n863_));
  NOi21      u0835(.An(f), .B(d), .Y(men_men_n864_));
  NA2        u0836(.A(men_men_n864_), .B(m), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n865_), .B(men_men_n52_), .Y(men_men_n866_));
  NOi32      u0838(.An(g), .Bn(f), .C(d), .Y(men_men_n867_));
  NA4        u0839(.A(men_men_n867_), .B(men_men_n607_), .C(men_men_n29_), .D(m), .Y(men_men_n868_));
  NOi21      u0840(.An(men_men_n312_), .B(men_men_n868_), .Y(men_men_n869_));
  AOI210     u0841(.A0(men_men_n866_), .A1(men_men_n551_), .B0(men_men_n869_), .Y(men_men_n870_));
  NA3        u0842(.A(men_men_n311_), .B(men_men_n261_), .C(men_men_n119_), .Y(men_men_n871_));
  AN2        u0843(.A(f), .B(d), .Y(men_men_n872_));
  NA3        u0844(.A(men_men_n484_), .B(men_men_n872_), .C(men_men_n86_), .Y(men_men_n873_));
  NO3        u0845(.A(men_men_n873_), .B(men_men_n75_), .C(men_men_n215_), .Y(men_men_n874_));
  NO2        u0846(.A(men_men_n285_), .B(men_men_n56_), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n871_), .B(men_men_n874_), .Y(men_men_n876_));
  NAi41      u0848(.An(men_men_n495_), .B(men_men_n876_), .C(men_men_n870_), .D(men_men_n863_), .Y(men_men_n877_));
  NO4        u0849(.A(men_men_n622_), .B(men_men_n130_), .C(men_men_n329_), .D(men_men_n150_), .Y(men_men_n878_));
  NO2        u0850(.A(men_men_n651_), .B(men_men_n329_), .Y(men_men_n879_));
  AN2        u0851(.A(men_men_n879_), .B(men_men_n681_), .Y(men_men_n880_));
  NO3        u0852(.A(men_men_n880_), .B(men_men_n878_), .C(men_men_n236_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n605_), .B(men_men_n86_), .Y(men_men_n882_));
  NO2        u0854(.A(men_men_n855_), .B(men_men_n882_), .Y(men_men_n883_));
  NA3        u0855(.A(men_men_n158_), .B(men_men_n110_), .C(men_men_n109_), .Y(men_men_n884_));
  OAI220     u0856(.A0(men_men_n873_), .A1(men_men_n434_), .B0(men_men_n341_), .B1(men_men_n884_), .Y(men_men_n885_));
  NOi41      u0857(.An(men_men_n225_), .B(men_men_n885_), .C(men_men_n883_), .D(men_men_n306_), .Y(men_men_n886_));
  NA2        u0858(.A(c), .B(men_men_n116_), .Y(men_men_n887_));
  NO2        u0859(.A(men_men_n887_), .B(men_men_n413_), .Y(men_men_n888_));
  NA3        u0860(.A(men_men_n888_), .B(men_men_n515_), .C(f), .Y(men_men_n889_));
  OR2        u0861(.A(men_men_n658_), .B(men_men_n547_), .Y(men_men_n890_));
  INV        u0862(.A(men_men_n890_), .Y(men_men_n891_));
  NA2        u0863(.A(men_men_n811_), .B(men_men_n112_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n892_), .B(men_men_n891_), .Y(men_men_n893_));
  NA4        u0865(.A(men_men_n893_), .B(men_men_n889_), .C(men_men_n886_), .D(men_men_n881_), .Y(men_men_n894_));
  NO4        u0866(.A(men_men_n894_), .B(men_men_n877_), .C(men_men_n861_), .D(men_men_n848_), .Y(men_men_n895_));
  OR2        u0867(.A(men_men_n873_), .B(men_men_n75_), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n833_), .B(g), .Y(men_men_n897_));
  AOI210     u0869(.A0(men_men_n897_), .A1(men_men_n293_), .B0(men_men_n896_), .Y(men_men_n898_));
  NO2        u0870(.A(men_men_n334_), .B(men_men_n844_), .Y(men_men_n899_));
  NO2        u0871(.A(men_men_n134_), .B(men_men_n130_), .Y(men_men_n900_));
  NO2        u0872(.A(men_men_n232_), .B(men_men_n226_), .Y(men_men_n901_));
  AOI220     u0873(.A0(men_men_n901_), .A1(men_men_n229_), .B0(men_men_n304_), .B1(men_men_n900_), .Y(men_men_n902_));
  NO2        u0874(.A(men_men_n434_), .B(men_men_n832_), .Y(men_men_n903_));
  NA2        u0875(.A(men_men_n903_), .B(men_men_n568_), .Y(men_men_n904_));
  NA2        u0876(.A(men_men_n904_), .B(men_men_n902_), .Y(men_men_n905_));
  NA2        u0877(.A(e), .B(d), .Y(men_men_n906_));
  OAI220     u0878(.A0(men_men_n906_), .A1(c), .B0(men_men_n324_), .B1(d), .Y(men_men_n907_));
  NA3        u0879(.A(men_men_n907_), .B(men_men_n459_), .C(men_men_n513_), .Y(men_men_n908_));
  AOI210     u0880(.A0(men_men_n521_), .A1(men_men_n181_), .B0(men_men_n232_), .Y(men_men_n909_));
  AOI210     u0881(.A0(men_men_n623_), .A1(men_men_n350_), .B0(men_men_n909_), .Y(men_men_n910_));
  NA2        u0882(.A(men_men_n285_), .B(men_men_n164_), .Y(men_men_n911_));
  NA2        u0883(.A(men_men_n874_), .B(men_men_n911_), .Y(men_men_n912_));
  NA3        u0884(.A(men_men_n167_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n913_));
  NA4        u0885(.A(men_men_n913_), .B(men_men_n912_), .C(men_men_n910_), .D(men_men_n908_), .Y(men_men_n914_));
  NO4        u0886(.A(men_men_n914_), .B(men_men_n905_), .C(men_men_n899_), .D(men_men_n898_), .Y(men_men_n915_));
  NA2        u0887(.A(men_men_n849_), .B(men_men_n31_), .Y(men_men_n916_));
  AO210      u0888(.A0(men_men_n916_), .A1(men_men_n702_), .B0(men_men_n218_), .Y(men_men_n917_));
  OAI220     u0889(.A0(men_men_n622_), .A1(men_men_n61_), .B0(men_men_n301_), .B1(j), .Y(men_men_n918_));
  AOI220     u0890(.A0(men_men_n918_), .A1(men_men_n879_), .B0(men_men_n612_), .B1(men_men_n621_), .Y(men_men_n919_));
  OAI210     u0891(.A0(men_men_n838_), .A1(men_men_n171_), .B0(men_men_n919_), .Y(men_men_n920_));
  OAI210     u0892(.A0(men_men_n833_), .A1(men_men_n911_), .B0(men_men_n867_), .Y(men_men_n921_));
  NO2        u0893(.A(men_men_n921_), .B(men_men_n608_), .Y(men_men_n922_));
  AN2        u0894(.A(men_men_n854_), .B(men_men_n843_), .Y(men_men_n923_));
  NOi31      u0895(.An(men_men_n551_), .B(men_men_n865_), .C(men_men_n293_), .Y(men_men_n924_));
  NO4        u0896(.A(men_men_n924_), .B(men_men_n923_), .C(men_men_n922_), .D(men_men_n920_), .Y(men_men_n925_));
  AO220      u0897(.A0(men_men_n459_), .A1(men_men_n750_), .B0(men_men_n176_), .B1(f), .Y(men_men_n926_));
  OAI210     u0898(.A0(men_men_n926_), .A1(men_men_n462_), .B0(men_men_n907_), .Y(men_men_n927_));
  NO2        u0899(.A(men_men_n444_), .B(men_men_n71_), .Y(men_men_n928_));
  OAI210     u0900(.A0(men_men_n847_), .A1(men_men_n928_), .B0(men_men_n706_), .Y(men_men_n929_));
  AN4        u0901(.A(men_men_n929_), .B(men_men_n927_), .C(men_men_n925_), .D(men_men_n917_), .Y(men_men_n930_));
  NA4        u0902(.A(men_men_n930_), .B(men_men_n915_), .C(men_men_n895_), .D(men_men_n840_), .Y(men12));
  NO2        u0903(.A(men_men_n457_), .B(c), .Y(men_men_n932_));
  NO4        u0904(.A(men_men_n449_), .B(men_men_n252_), .C(men_men_n591_), .D(men_men_n215_), .Y(men_men_n933_));
  NA2        u0905(.A(men_men_n933_), .B(men_men_n932_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n551_), .B(men_men_n928_), .Y(men_men_n935_));
  NO2        u0907(.A(men_men_n457_), .B(men_men_n116_), .Y(men_men_n936_));
  NO2        u0908(.A(men_men_n850_), .B(men_men_n357_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n658_), .B(men_men_n382_), .Y(men_men_n938_));
  AOI220     u0910(.A0(men_men_n938_), .A1(men_men_n549_), .B0(men_men_n937_), .B1(men_men_n936_), .Y(men_men_n939_));
  NA4        u0911(.A(men_men_n939_), .B(men_men_n935_), .C(men_men_n934_), .D(men_men_n448_), .Y(men_men_n940_));
  AOI210     u0912(.A0(men_men_n235_), .A1(men_men_n340_), .B0(men_men_n203_), .Y(men_men_n941_));
  OR2        u0913(.A(men_men_n941_), .B(men_men_n933_), .Y(men_men_n942_));
  AOI210     u0914(.A0(men_men_n337_), .A1(men_men_n394_), .B0(men_men_n215_), .Y(men_men_n943_));
  OAI210     u0915(.A0(men_men_n943_), .A1(men_men_n942_), .B0(men_men_n408_), .Y(men_men_n944_));
  NO2        u0916(.A(men_men_n637_), .B(men_men_n262_), .Y(men_men_n945_));
  NO2        u0917(.A(men_men_n598_), .B(men_men_n842_), .Y(men_men_n946_));
  NO2        u0918(.A(men_men_n149_), .B(men_men_n239_), .Y(men_men_n947_));
  NA3        u0919(.A(men_men_n947_), .B(men_men_n242_), .C(i), .Y(men_men_n948_));
  NA2        u0920(.A(men_men_n948_), .B(men_men_n944_), .Y(men_men_n949_));
  OR2        u0921(.A(men_men_n325_), .B(men_men_n936_), .Y(men_men_n950_));
  NA2        u0922(.A(men_men_n950_), .B(men_men_n358_), .Y(men_men_n951_));
  NA4        u0923(.A(men_men_n450_), .B(men_men_n442_), .C(men_men_n182_), .D(g), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n952_), .B(men_men_n951_), .Y(men_men_n953_));
  NO3        u0925(.A(men_men_n663_), .B(men_men_n94_), .C(men_men_n45_), .Y(men_men_n954_));
  NO4        u0926(.A(men_men_n954_), .B(men_men_n953_), .C(men_men_n949_), .D(men_men_n940_), .Y(men_men_n955_));
  NO2        u0927(.A(men_men_n373_), .B(men_men_n372_), .Y(men_men_n956_));
  NA2        u0928(.A(men_men_n596_), .B(men_men_n73_), .Y(men_men_n957_));
  NA2        u0929(.A(men_men_n561_), .B(men_men_n142_), .Y(men_men_n958_));
  NOi21      u0930(.An(men_men_n34_), .B(men_men_n651_), .Y(men_men_n959_));
  AOI220     u0931(.A0(men_men_n959_), .A1(men_men_n958_), .B0(men_men_n957_), .B1(men_men_n956_), .Y(men_men_n960_));
  OAI210     u0932(.A0(men_men_n251_), .A1(men_men_n45_), .B0(men_men_n960_), .Y(men_men_n961_));
  NA2        u0933(.A(men_men_n440_), .B(men_men_n264_), .Y(men_men_n962_));
  NO3        u0934(.A(men_men_n820_), .B(men_men_n91_), .C(men_men_n413_), .Y(men_men_n963_));
  NAi31      u0935(.An(men_men_n963_), .B(men_men_n962_), .C(men_men_n322_), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n965_));
  NO2        u0937(.A(men_men_n509_), .B(men_men_n301_), .Y(men_men_n966_));
  INV        u0938(.A(men_men_n966_), .Y(men_men_n967_));
  NO2        u0939(.A(men_men_n967_), .B(men_men_n142_), .Y(men_men_n968_));
  NA2        u0940(.A(men_men_n632_), .B(men_men_n367_), .Y(men_men_n969_));
  OAI210     u0941(.A0(men_men_n739_), .A1(men_men_n969_), .B0(men_men_n371_), .Y(men_men_n970_));
  NO4        u0942(.A(men_men_n970_), .B(men_men_n968_), .C(men_men_n964_), .D(men_men_n961_), .Y(men_men_n971_));
  NA2        u0943(.A(men_men_n350_), .B(g), .Y(men_men_n972_));
  NA2        u0944(.A(men_men_n161_), .B(i), .Y(men_men_n973_));
  NA2        u0945(.A(men_men_n46_), .B(i), .Y(men_men_n974_));
  OAI220     u0946(.A0(men_men_n974_), .A1(men_men_n202_), .B0(men_men_n973_), .B1(men_men_n94_), .Y(men_men_n975_));
  AOI210     u0947(.A0(men_men_n424_), .A1(men_men_n37_), .B0(men_men_n975_), .Y(men_men_n976_));
  NO2        u0948(.A(men_men_n142_), .B(men_men_n86_), .Y(men_men_n977_));
  OR2        u0949(.A(men_men_n977_), .B(men_men_n560_), .Y(men_men_n978_));
  NA2        u0950(.A(men_men_n561_), .B(men_men_n386_), .Y(men_men_n979_));
  AOI210     u0951(.A0(men_men_n979_), .A1(n), .B0(men_men_n978_), .Y(men_men_n980_));
  OAI220     u0952(.A0(men_men_n980_), .A1(men_men_n972_), .B0(men_men_n976_), .B1(men_men_n334_), .Y(men_men_n981_));
  NO2        u0953(.A(men_men_n658_), .B(men_men_n503_), .Y(men_men_n982_));
  NA3        u0954(.A(men_men_n345_), .B(men_men_n628_), .C(i), .Y(men_men_n983_));
  OAI210     u0955(.A0(men_men_n444_), .A1(men_men_n311_), .B0(men_men_n983_), .Y(men_men_n984_));
  OAI220     u0956(.A0(men_men_n984_), .A1(men_men_n982_), .B0(men_men_n677_), .B1(men_men_n760_), .Y(men_men_n985_));
  NA2        u0957(.A(men_men_n609_), .B(men_men_n114_), .Y(men_men_n986_));
  NA3        u0958(.A(men_men_n628_), .B(men_men_n82_), .C(i), .Y(men_men_n987_));
  OR2        u0959(.A(men_men_n987_), .B(men_men_n986_), .Y(men_men_n988_));
  NA3        u0960(.A(men_men_n326_), .B(men_men_n118_), .C(g), .Y(men_men_n989_));
  AOI210     u0961(.A0(men_men_n674_), .A1(men_men_n989_), .B0(m), .Y(men_men_n990_));
  OAI210     u0962(.A0(men_men_n990_), .A1(men_men_n937_), .B0(men_men_n325_), .Y(men_men_n991_));
  NA2        u0963(.A(men_men_n693_), .B(men_men_n882_), .Y(men_men_n992_));
  INV        u0964(.A(men_men_n445_), .Y(men_men_n993_));
  NA2        u0965(.A(men_men_n223_), .B(men_men_n79_), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n994_), .B(men_men_n987_), .Y(men_men_n995_));
  AOI220     u0967(.A0(men_men_n995_), .A1(men_men_n258_), .B0(men_men_n993_), .B1(men_men_n992_), .Y(men_men_n996_));
  NA4        u0968(.A(men_men_n996_), .B(men_men_n991_), .C(men_men_n988_), .D(men_men_n985_), .Y(men_men_n997_));
  NO2        u0969(.A(men_men_n382_), .B(men_men_n93_), .Y(men_men_n998_));
  OAI210     u0970(.A0(men_men_n998_), .A1(men_men_n945_), .B0(men_men_n240_), .Y(men_men_n999_));
  NA2        u0971(.A(men_men_n662_), .B(men_men_n90_), .Y(men_men_n1000_));
  NO2        u0972(.A(men_men_n465_), .B(men_men_n215_), .Y(men_men_n1001_));
  AOI220     u0973(.A0(men_men_n1001_), .A1(men_men_n387_), .B0(men_men_n950_), .B1(men_men_n219_), .Y(men_men_n1002_));
  AOI220     u0974(.A0(men_men_n938_), .A1(men_men_n947_), .B0(men_men_n597_), .B1(men_men_n92_), .Y(men_men_n1003_));
  NA4        u0975(.A(men_men_n1003_), .B(men_men_n1002_), .C(men_men_n1000_), .D(men_men_n999_), .Y(men_men_n1004_));
  OAI210     u0976(.A0(men_men_n993_), .A1(men_men_n946_), .B0(men_men_n549_), .Y(men_men_n1005_));
  AOI210     u0977(.A0(men_men_n425_), .A1(men_men_n417_), .B0(men_men_n820_), .Y(men_men_n1006_));
  INV        u0978(.A(men_men_n1006_), .Y(men_men_n1007_));
  NA2        u0979(.A(men_men_n990_), .B(men_men_n936_), .Y(men_men_n1008_));
  NA2        u0980(.A(men_men_n642_), .B(men_men_n538_), .Y(men_men_n1009_));
  NA4        u0981(.A(men_men_n1009_), .B(men_men_n1008_), .C(men_men_n1007_), .D(men_men_n1005_), .Y(men_men_n1010_));
  NO4        u0982(.A(men_men_n1010_), .B(men_men_n1004_), .C(men_men_n997_), .D(men_men_n981_), .Y(men_men_n1011_));
  NAi31      u0983(.An(men_men_n139_), .B(men_men_n426_), .C(n), .Y(men_men_n1012_));
  NO3        u0984(.A(men_men_n126_), .B(men_men_n343_), .C(men_men_n851_), .Y(men_men_n1013_));
  NO2        u0985(.A(men_men_n1013_), .B(men_men_n1012_), .Y(men_men_n1014_));
  NO3        u0986(.A(men_men_n271_), .B(men_men_n139_), .C(men_men_n413_), .Y(men_men_n1015_));
  AOI210     u0987(.A0(men_men_n1015_), .A1(men_men_n504_), .B0(men_men_n1014_), .Y(men_men_n1016_));
  INV        u0988(.A(men_men_n1016_), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n232_), .B(men_men_n172_), .Y(men_men_n1018_));
  NO3        u0990(.A(men_men_n308_), .B(men_men_n450_), .C(men_men_n176_), .Y(men_men_n1019_));
  NOi31      u0991(.An(men_men_n1018_), .B(men_men_n1019_), .C(men_men_n215_), .Y(men_men_n1020_));
  NAi21      u0992(.An(men_men_n561_), .B(men_men_n1001_), .Y(men_men_n1021_));
  NA2        u0993(.A(men_men_n443_), .B(men_men_n882_), .Y(men_men_n1022_));
  NO3        u0994(.A(men_men_n444_), .B(men_men_n311_), .C(men_men_n75_), .Y(men_men_n1023_));
  AOI220     u0995(.A0(men_men_n1023_), .A1(men_men_n1022_), .B0(men_men_n488_), .B1(g), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n1024_), .B(men_men_n1021_), .Y(men_men_n1025_));
  NO2        u0997(.A(men_men_n983_), .B(men_men_n606_), .Y(men_men_n1026_));
  NO2        u0998(.A(men_men_n659_), .B(men_men_n382_), .Y(men_men_n1027_));
  NA2        u0999(.A(men_men_n941_), .B(men_men_n932_), .Y(men_men_n1028_));
  OAI220     u1000(.A0(men_men_n938_), .A1(men_men_n946_), .B0(men_men_n551_), .B1(men_men_n433_), .Y(men_men_n1029_));
  NA3        u1001(.A(men_men_n1029_), .B(men_men_n1028_), .C(men_men_n620_), .Y(men_men_n1030_));
  OAI210     u1002(.A0(men_men_n941_), .A1(men_men_n933_), .B0(men_men_n1018_), .Y(men_men_n1031_));
  NA3        u1003(.A(men_men_n979_), .B(men_men_n493_), .C(men_men_n46_), .Y(men_men_n1032_));
  AOI210     u1004(.A0(men_men_n385_), .A1(men_men_n383_), .B0(men_men_n333_), .Y(men_men_n1033_));
  NA4        u1005(.A(men_men_n1033_), .B(men_men_n1032_), .C(men_men_n1031_), .D(men_men_n272_), .Y(men_men_n1034_));
  OR4        u1006(.A(men_men_n1034_), .B(men_men_n1030_), .C(men_men_n1027_), .D(men_men_n1026_), .Y(men_men_n1035_));
  NO4        u1007(.A(men_men_n1035_), .B(men_men_n1025_), .C(men_men_n1020_), .D(men_men_n1017_), .Y(men_men_n1036_));
  NA4        u1008(.A(men_men_n1036_), .B(men_men_n1011_), .C(men_men_n971_), .D(men_men_n955_), .Y(men13));
  AN2        u1009(.A(c), .B(b), .Y(men_men_n1038_));
  NA3        u1010(.A(men_men_n250_), .B(men_men_n1038_), .C(m), .Y(men_men_n1039_));
  NA2        u1011(.A(men_men_n502_), .B(f), .Y(men_men_n1040_));
  NO4        u1012(.A(men_men_n1040_), .B(men_men_n1039_), .C(j), .D(men_men_n592_), .Y(men_men_n1041_));
  NA2        u1013(.A(men_men_n264_), .B(men_men_n1038_), .Y(men_men_n1042_));
  NO4        u1014(.A(men_men_n1042_), .B(men_men_n1040_), .C(men_men_n973_), .D(a), .Y(men_men_n1043_));
  NAi32      u1015(.An(d), .Bn(c), .C(e), .Y(men_men_n1044_));
  NA2        u1016(.A(men_men_n138_), .B(men_men_n45_), .Y(men_men_n1045_));
  NO4        u1017(.A(men_men_n1045_), .B(men_men_n1044_), .C(men_men_n598_), .D(men_men_n307_), .Y(men_men_n1046_));
  NA2        u1018(.A(men_men_n666_), .B(men_men_n226_), .Y(men_men_n1047_));
  NA2        u1019(.A(men_men_n416_), .B(men_men_n214_), .Y(men_men_n1048_));
  AN2        u1020(.A(d), .B(c), .Y(men_men_n1049_));
  NA2        u1021(.A(men_men_n1049_), .B(men_men_n116_), .Y(men_men_n1050_));
  NO4        u1022(.A(men_men_n1050_), .B(men_men_n1048_), .C(men_men_n177_), .D(men_men_n168_), .Y(men_men_n1051_));
  NA2        u1023(.A(men_men_n502_), .B(c), .Y(men_men_n1052_));
  NO4        u1024(.A(men_men_n1045_), .B(men_men_n595_), .C(men_men_n1052_), .D(men_men_n307_), .Y(men_men_n1053_));
  AO210      u1025(.A0(men_men_n1051_), .A1(men_men_n1047_), .B0(men_men_n1053_), .Y(men_men_n1054_));
  OR4        u1026(.A(men_men_n1054_), .B(men_men_n1046_), .C(men_men_n1043_), .D(men_men_n1041_), .Y(men_men_n1055_));
  NAi32      u1027(.An(f), .Bn(e), .C(c), .Y(men_men_n1056_));
  NO2        u1028(.A(men_men_n1056_), .B(men_men_n144_), .Y(men_men_n1057_));
  NA2        u1029(.A(men_men_n1057_), .B(g), .Y(men_men_n1058_));
  OR3        u1030(.A(men_men_n226_), .B(men_men_n177_), .C(men_men_n168_), .Y(men_men_n1059_));
  NO2        u1031(.A(men_men_n1059_), .B(men_men_n1058_), .Y(men_men_n1060_));
  NO2        u1032(.A(men_men_n1052_), .B(men_men_n307_), .Y(men_men_n1061_));
  NO2        u1033(.A(j), .B(men_men_n45_), .Y(men_men_n1062_));
  NA2        u1034(.A(men_men_n630_), .B(men_men_n1062_), .Y(men_men_n1063_));
  NOi21      u1035(.An(men_men_n1061_), .B(men_men_n1063_), .Y(men_men_n1064_));
  NO2        u1036(.A(men_men_n762_), .B(men_men_n113_), .Y(men_men_n1065_));
  NOi41      u1037(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1066_));
  NA2        u1038(.A(men_men_n1066_), .B(men_men_n1065_), .Y(men_men_n1067_));
  NO2        u1039(.A(men_men_n1067_), .B(men_men_n1058_), .Y(men_men_n1068_));
  OR3        u1040(.A(e), .B(d), .C(c), .Y(men_men_n1069_));
  NA3        u1041(.A(k), .B(j), .C(i), .Y(men_men_n1070_));
  NO3        u1042(.A(men_men_n1070_), .B(men_men_n307_), .C(men_men_n93_), .Y(men_men_n1071_));
  NOi21      u1043(.An(men_men_n1071_), .B(men_men_n1069_), .Y(men_men_n1072_));
  OR4        u1044(.A(men_men_n1072_), .B(men_men_n1068_), .C(men_men_n1064_), .D(men_men_n1060_), .Y(men_men_n1073_));
  NA3        u1045(.A(men_men_n473_), .B(men_men_n336_), .C(men_men_n56_), .Y(men_men_n1074_));
  NO2        u1046(.A(men_men_n1074_), .B(men_men_n1063_), .Y(men_men_n1075_));
  NO4        u1047(.A(men_men_n1074_), .B(men_men_n595_), .C(men_men_n456_), .D(men_men_n45_), .Y(men_men_n1076_));
  NO2        u1048(.A(f), .B(c), .Y(men_men_n1077_));
  NOi21      u1049(.An(men_men_n1077_), .B(men_men_n449_), .Y(men_men_n1078_));
  NA2        u1050(.A(men_men_n1078_), .B(men_men_n59_), .Y(men_men_n1079_));
  OR2        u1051(.A(k), .B(i), .Y(men_men_n1080_));
  NO3        u1052(.A(men_men_n1080_), .B(men_men_n246_), .C(l), .Y(men_men_n1081_));
  NOi31      u1053(.An(men_men_n1081_), .B(men_men_n1079_), .C(j), .Y(men_men_n1082_));
  OR3        u1054(.A(men_men_n1082_), .B(men_men_n1076_), .C(men_men_n1075_), .Y(men_men_n1083_));
  OR3        u1055(.A(men_men_n1083_), .B(men_men_n1073_), .C(men_men_n1055_), .Y(men02));
  OR2        u1056(.A(l), .B(k), .Y(men_men_n1085_));
  OR3        u1057(.A(h), .B(g), .C(f), .Y(men_men_n1086_));
  OR3        u1058(.A(n), .B(m), .C(i), .Y(men_men_n1087_));
  NO4        u1059(.A(men_men_n1087_), .B(men_men_n1086_), .C(men_men_n1085_), .D(men_men_n1069_), .Y(men_men_n1088_));
  NOi31      u1060(.An(e), .B(d), .C(c), .Y(men_men_n1089_));
  AOI210     u1061(.A0(men_men_n1071_), .A1(men_men_n1089_), .B0(men_men_n1046_), .Y(men_men_n1090_));
  AN3        u1062(.A(g), .B(f), .C(c), .Y(men_men_n1091_));
  NA3        u1063(.A(men_men_n1091_), .B(men_men_n473_), .C(h), .Y(men_men_n1092_));
  OR2        u1064(.A(men_men_n1070_), .B(men_men_n307_), .Y(men_men_n1093_));
  OR2        u1065(.A(men_men_n1093_), .B(men_men_n1092_), .Y(men_men_n1094_));
  NO3        u1066(.A(men_men_n1074_), .B(men_men_n1045_), .C(men_men_n595_), .Y(men_men_n1095_));
  NO2        u1067(.A(men_men_n1095_), .B(men_men_n1060_), .Y(men_men_n1096_));
  NA3        u1068(.A(l), .B(k), .C(j), .Y(men_men_n1097_));
  NA2        u1069(.A(i), .B(h), .Y(men_men_n1098_));
  NO3        u1070(.A(men_men_n1098_), .B(men_men_n1097_), .C(men_men_n130_), .Y(men_men_n1099_));
  NO3        u1071(.A(men_men_n140_), .B(men_men_n283_), .C(men_men_n215_), .Y(men_men_n1100_));
  AOI210     u1072(.A0(men_men_n1100_), .A1(men_men_n1099_), .B0(men_men_n1064_), .Y(men_men_n1101_));
  NA3        u1073(.A(c), .B(b), .C(a), .Y(men_men_n1102_));
  NO3        u1074(.A(men_men_n1102_), .B(men_men_n906_), .C(men_men_n214_), .Y(men_men_n1103_));
  NO4        u1075(.A(men_men_n1070_), .B(men_men_n301_), .C(men_men_n49_), .D(men_men_n113_), .Y(men_men_n1104_));
  AOI210     u1076(.A0(men_men_n1104_), .A1(men_men_n1103_), .B0(men_men_n1075_), .Y(men_men_n1105_));
  AN4        u1077(.A(men_men_n1105_), .B(men_men_n1101_), .C(men_men_n1096_), .D(men_men_n1094_), .Y(men_men_n1106_));
  NO2        u1078(.A(men_men_n1050_), .B(men_men_n1048_), .Y(men_men_n1107_));
  NA2        u1079(.A(men_men_n1067_), .B(men_men_n1059_), .Y(men_men_n1108_));
  AOI210     u1080(.A0(men_men_n1108_), .A1(men_men_n1107_), .B0(men_men_n1041_), .Y(men_men_n1109_));
  NAi41      u1081(.An(men_men_n1088_), .B(men_men_n1109_), .C(men_men_n1106_), .D(men_men_n1090_), .Y(men03));
  NO2        u1082(.A(men_men_n534_), .B(men_men_n602_), .Y(men_men_n1111_));
  NA4        u1083(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(men_men_n214_), .Y(men_men_n1112_));
  NA4        u1084(.A(men_men_n583_), .B(m), .C(men_men_n113_), .D(men_men_n214_), .Y(men_men_n1113_));
  NA3        u1085(.A(men_men_n1113_), .B(men_men_n374_), .C(men_men_n1112_), .Y(men_men_n1114_));
  NO2        u1086(.A(men_men_n1114_), .B(men_men_n1111_), .Y(men_men_n1115_));
  NOi31      u1087(.An(men_men_n809_), .B(men_men_n856_), .C(men_men_n845_), .Y(men_men_n1116_));
  OAI220     u1088(.A0(men_men_n1116_), .A1(men_men_n693_), .B0(men_men_n1115_), .B1(men_men_n596_), .Y(men_men_n1117_));
  NOi31      u1089(.An(i), .B(k), .C(j), .Y(men_men_n1118_));
  NA4        u1090(.A(men_men_n1118_), .B(men_men_n1089_), .C(men_men_n345_), .D(men_men_n336_), .Y(men_men_n1119_));
  OAI210     u1091(.A0(men_men_n820_), .A1(men_men_n427_), .B0(men_men_n1119_), .Y(men_men_n1120_));
  NOi31      u1092(.An(m), .B(n), .C(f), .Y(men_men_n1121_));
  NA2        u1093(.A(men_men_n1121_), .B(men_men_n51_), .Y(men_men_n1122_));
  AN2        u1094(.A(e), .B(c), .Y(men_men_n1123_));
  NA2        u1095(.A(men_men_n1123_), .B(a), .Y(men_men_n1124_));
  OAI220     u1096(.A0(men_men_n1124_), .A1(men_men_n1122_), .B0(men_men_n890_), .B1(men_men_n432_), .Y(men_men_n1125_));
  NA2        u1097(.A(men_men_n513_), .B(l), .Y(men_men_n1126_));
  NOi31      u1098(.An(men_men_n867_), .B(men_men_n1039_), .C(men_men_n1126_), .Y(men_men_n1127_));
  NO4        u1099(.A(men_men_n1127_), .B(men_men_n1125_), .C(men_men_n1120_), .D(men_men_n1006_), .Y(men_men_n1128_));
  NO2        u1100(.A(men_men_n283_), .B(a), .Y(men_men_n1129_));
  INV        u1101(.A(men_men_n1046_), .Y(men_men_n1130_));
  NO2        u1102(.A(men_men_n1098_), .B(men_men_n491_), .Y(men_men_n1131_));
  NO2        u1103(.A(men_men_n89_), .B(g), .Y(men_men_n1132_));
  AOI210     u1104(.A0(men_men_n1132_), .A1(men_men_n1131_), .B0(men_men_n1081_), .Y(men_men_n1133_));
  OR2        u1105(.A(men_men_n1133_), .B(men_men_n1079_), .Y(men_men_n1134_));
  NA3        u1106(.A(men_men_n1134_), .B(men_men_n1130_), .C(men_men_n1128_), .Y(men_men_n1135_));
  NO4        u1107(.A(men_men_n1135_), .B(men_men_n1117_), .C(men_men_n821_), .D(men_men_n573_), .Y(men_men_n1136_));
  NA2        u1108(.A(c), .B(b), .Y(men_men_n1137_));
  NO2        u1109(.A(men_men_n705_), .B(men_men_n1137_), .Y(men_men_n1138_));
  OAI210     u1110(.A0(men_men_n865_), .A1(men_men_n836_), .B0(men_men_n420_), .Y(men_men_n1139_));
  OAI210     u1111(.A0(men_men_n1139_), .A1(men_men_n866_), .B0(men_men_n1138_), .Y(men_men_n1140_));
  NAi21      u1112(.An(men_men_n428_), .B(men_men_n1138_), .Y(men_men_n1141_));
  NA3        u1113(.A(men_men_n433_), .B(men_men_n566_), .C(f), .Y(men_men_n1142_));
  OAI210     u1114(.A0(men_men_n555_), .A1(men_men_n39_), .B0(men_men_n1129_), .Y(men_men_n1143_));
  NA3        u1115(.A(men_men_n1143_), .B(men_men_n1142_), .C(men_men_n1141_), .Y(men_men_n1144_));
  NA2        u1116(.A(men_men_n261_), .B(men_men_n119_), .Y(men_men_n1145_));
  OAI210     u1117(.A0(men_men_n1145_), .A1(men_men_n287_), .B0(g), .Y(men_men_n1146_));
  NAi21      u1118(.An(f), .B(d), .Y(men_men_n1147_));
  NO2        u1119(.A(men_men_n1147_), .B(men_men_n1102_), .Y(men_men_n1148_));
  INV        u1120(.A(men_men_n1148_), .Y(men_men_n1149_));
  AOI210     u1121(.A0(men_men_n1146_), .A1(men_men_n293_), .B0(men_men_n1149_), .Y(men_men_n1150_));
  AOI210     u1122(.A0(men_men_n1150_), .A1(men_men_n114_), .B0(men_men_n1144_), .Y(men_men_n1151_));
  NA2        u1123(.A(men_men_n476_), .B(men_men_n475_), .Y(men_men_n1152_));
  NO2        u1124(.A(men_men_n183_), .B(men_men_n239_), .Y(men_men_n1153_));
  NA2        u1125(.A(men_men_n1153_), .B(m), .Y(men_men_n1154_));
  NA2        u1126(.A(men_men_n1126_), .B(men_men_n479_), .Y(men_men_n1155_));
  OAI210     u1127(.A0(men_men_n1155_), .A1(men_men_n312_), .B0(men_men_n477_), .Y(men_men_n1156_));
  AOI210     u1128(.A0(men_men_n1156_), .A1(men_men_n1152_), .B0(men_men_n1154_), .Y(men_men_n1157_));
  NA2        u1129(.A(men_men_n568_), .B(men_men_n415_), .Y(men_men_n1158_));
  NA2        u1130(.A(men_men_n453_), .B(men_men_n1148_), .Y(men_men_n1159_));
  NO2        u1131(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n1160_));
  AOI210     u1132(.A0(men_men_n1153_), .A1(men_men_n435_), .B0(men_men_n963_), .Y(men_men_n1161_));
  NAi41      u1133(.An(men_men_n1160_), .B(men_men_n1161_), .C(men_men_n1159_), .D(men_men_n1158_), .Y(men_men_n1162_));
  NO2        u1134(.A(men_men_n1162_), .B(men_men_n1157_), .Y(men_men_n1163_));
  NA4        u1135(.A(men_men_n1163_), .B(men_men_n1151_), .C(men_men_n1140_), .D(men_men_n1136_), .Y(men00));
  AOI210     u1136(.A0(men_men_n300_), .A1(men_men_n215_), .B0(men_men_n275_), .Y(men_men_n1165_));
  NO2        u1137(.A(men_men_n1165_), .B(men_men_n586_), .Y(men_men_n1166_));
  AOI210     u1138(.A0(men_men_n903_), .A1(men_men_n947_), .B0(men_men_n1120_), .Y(men_men_n1167_));
  NO2        u1139(.A(men_men_n1095_), .B(men_men_n963_), .Y(men_men_n1168_));
  NA3        u1140(.A(men_men_n1168_), .B(men_men_n1167_), .C(men_men_n1007_), .Y(men_men_n1169_));
  NA2        u1141(.A(men_men_n515_), .B(f), .Y(men_men_n1170_));
  OAI210     u1142(.A0(men_men_n1013_), .A1(men_men_n40_), .B0(men_men_n644_), .Y(men_men_n1171_));
  NA3        u1143(.A(men_men_n1171_), .B(men_men_n257_), .C(n), .Y(men_men_n1172_));
  AOI210     u1144(.A0(men_men_n1172_), .A1(men_men_n1170_), .B0(men_men_n1050_), .Y(men_men_n1173_));
  NO4        u1145(.A(men_men_n1173_), .B(men_men_n1169_), .C(men_men_n1166_), .D(men_men_n1073_), .Y(men_men_n1174_));
  NA3        u1146(.A(men_men_n167_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1175_));
  NA3        u1147(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1176_));
  NOi31      u1148(.An(n), .B(m), .C(i), .Y(men_men_n1177_));
  NA3        u1149(.A(men_men_n1177_), .B(men_men_n647_), .C(men_men_n51_), .Y(men_men_n1178_));
  OAI210     u1150(.A0(men_men_n1176_), .A1(men_men_n1175_), .B0(men_men_n1178_), .Y(men_men_n1179_));
  INV        u1151(.A(men_men_n585_), .Y(men_men_n1180_));
  NO4        u1152(.A(men_men_n1180_), .B(men_men_n1179_), .C(men_men_n1160_), .D(men_men_n924_), .Y(men_men_n1181_));
  NO4        u1153(.A(men_men_n494_), .B(men_men_n360_), .C(men_men_n1137_), .D(men_men_n59_), .Y(men_men_n1182_));
  NA3        u1154(.A(men_men_n388_), .B(men_men_n222_), .C(g), .Y(men_men_n1183_));
  OR2        u1155(.A(men_men_n1183_), .B(men_men_n1176_), .Y(men_men_n1184_));
  NO2        u1156(.A(h), .B(g), .Y(men_men_n1185_));
  NA4        u1157(.A(men_men_n504_), .B(men_men_n473_), .C(men_men_n1185_), .D(men_men_n1038_), .Y(men_men_n1186_));
  OAI220     u1158(.A0(men_men_n534_), .A1(men_men_n602_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1187_));
  NA2        u1159(.A(men_men_n1187_), .B(men_men_n542_), .Y(men_men_n1188_));
  NA3        u1160(.A(men_men_n1188_), .B(men_men_n1186_), .C(men_men_n1184_), .Y(men_men_n1189_));
  NO3        u1161(.A(men_men_n1189_), .B(men_men_n1182_), .C(men_men_n265_), .Y(men_men_n1190_));
  INV        u1162(.A(men_men_n587_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n1191_), .B(men_men_n152_), .Y(men_men_n1192_));
  NO2        u1164(.A(men_men_n241_), .B(men_men_n182_), .Y(men_men_n1193_));
  NA2        u1165(.A(men_men_n1193_), .B(men_men_n433_), .Y(men_men_n1194_));
  NA3        u1166(.A(men_men_n180_), .B(men_men_n113_), .C(g), .Y(men_men_n1195_));
  NA3        u1167(.A(men_men_n473_), .B(men_men_n40_), .C(f), .Y(men_men_n1196_));
  NOi31      u1168(.An(men_men_n875_), .B(men_men_n1196_), .C(men_men_n1195_), .Y(men_men_n1197_));
  NAi31      u1169(.An(men_men_n187_), .B(men_men_n862_), .C(men_men_n473_), .Y(men_men_n1198_));
  NAi31      u1170(.An(men_men_n1197_), .B(men_men_n1198_), .C(men_men_n1194_), .Y(men_men_n1199_));
  NO2        u1171(.A(men_men_n274_), .B(men_men_n75_), .Y(men_men_n1200_));
  NO3        u1172(.A(men_men_n432_), .B(men_men_n832_), .C(n), .Y(men_men_n1201_));
  AOI210     u1173(.A0(men_men_n1201_), .A1(men_men_n1200_), .B0(men_men_n1088_), .Y(men_men_n1202_));
  NAi31      u1174(.An(men_men_n1053_), .B(men_men_n1202_), .C(men_men_n74_), .Y(men_men_n1203_));
  NO4        u1175(.A(men_men_n1203_), .B(men_men_n1199_), .C(men_men_n1192_), .D(men_men_n525_), .Y(men_men_n1204_));
  AN3        u1176(.A(men_men_n1204_), .B(men_men_n1190_), .C(men_men_n1181_), .Y(men_men_n1205_));
  NA3        u1177(.A(men_men_n1121_), .B(men_men_n609_), .C(men_men_n472_), .Y(men_men_n1206_));
  NA3        u1178(.A(men_men_n1206_), .B(men_men_n569_), .C(men_men_n244_), .Y(men_men_n1207_));
  NA2        u1179(.A(men_men_n1114_), .B(men_men_n542_), .Y(men_men_n1208_));
  NA4        u1180(.A(men_men_n647_), .B(men_men_n208_), .C(men_men_n222_), .D(men_men_n161_), .Y(men_men_n1209_));
  NA3        u1181(.A(men_men_n1209_), .B(men_men_n1208_), .C(men_men_n297_), .Y(men_men_n1210_));
  OAI210     u1182(.A0(men_men_n471_), .A1(men_men_n120_), .B0(men_men_n868_), .Y(men_men_n1211_));
  AOI220     u1183(.A0(men_men_n1211_), .A1(men_men_n1155_), .B0(men_men_n568_), .B1(men_men_n415_), .Y(men_men_n1212_));
  OR4        u1184(.A(men_men_n1050_), .B(men_men_n271_), .C(men_men_n224_), .D(e), .Y(men_men_n1213_));
  NO2        u1185(.A(men_men_n218_), .B(men_men_n215_), .Y(men_men_n1214_));
  NA2        u1186(.A(n), .B(e), .Y(men_men_n1215_));
  NO2        u1187(.A(men_men_n1215_), .B(men_men_n144_), .Y(men_men_n1216_));
  AOI220     u1188(.A0(men_men_n1216_), .A1(men_men_n273_), .B0(men_men_n849_), .B1(men_men_n1214_), .Y(men_men_n1217_));
  OAI210     u1189(.A0(men_men_n361_), .A1(men_men_n313_), .B0(men_men_n455_), .Y(men_men_n1218_));
  NA4        u1190(.A(men_men_n1218_), .B(men_men_n1217_), .C(men_men_n1213_), .D(men_men_n1212_), .Y(men_men_n1219_));
  AOI210     u1191(.A0(men_men_n1216_), .A1(men_men_n853_), .B0(men_men_n821_), .Y(men_men_n1220_));
  AOI220     u1192(.A0(men_men_n959_), .A1(men_men_n584_), .B0(men_men_n647_), .B1(men_men_n247_), .Y(men_men_n1221_));
  NO2        u1193(.A(men_men_n68_), .B(h), .Y(men_men_n1222_));
  NO3        u1194(.A(men_men_n1050_), .B(men_men_n1048_), .C(men_men_n731_), .Y(men_men_n1223_));
  NO2        u1195(.A(men_men_n1085_), .B(men_men_n130_), .Y(men_men_n1224_));
  AN2        u1196(.A(men_men_n1224_), .B(men_men_n1100_), .Y(men_men_n1225_));
  OAI210     u1197(.A0(men_men_n1225_), .A1(men_men_n1223_), .B0(men_men_n1222_), .Y(men_men_n1226_));
  NA4        u1198(.A(men_men_n1226_), .B(men_men_n1221_), .C(men_men_n1220_), .D(men_men_n870_), .Y(men_men_n1227_));
  NO4        u1199(.A(men_men_n1227_), .B(men_men_n1219_), .C(men_men_n1210_), .D(men_men_n1207_), .Y(men_men_n1228_));
  NA2        u1200(.A(men_men_n837_), .B(men_men_n759_), .Y(men_men_n1229_));
  NA4        u1201(.A(men_men_n1229_), .B(men_men_n1228_), .C(men_men_n1205_), .D(men_men_n1174_), .Y(men01));
  NO3        u1202(.A(men_men_n805_), .B(men_men_n797_), .C(men_men_n281_), .Y(men_men_n1231_));
  NA2        u1203(.A(men_men_n399_), .B(i), .Y(men_men_n1232_));
  NA3        u1204(.A(men_men_n1232_), .B(men_men_n1231_), .C(men_men_n1028_), .Y(men_men_n1233_));
  NA2        u1205(.A(men_men_n597_), .B(men_men_n92_), .Y(men_men_n1234_));
  NA2        u1206(.A(men_men_n561_), .B(men_men_n270_), .Y(men_men_n1235_));
  NA2        u1207(.A(men_men_n966_), .B(men_men_n1235_), .Y(men_men_n1236_));
  NA4        u1208(.A(men_men_n1236_), .B(men_men_n1234_), .C(men_men_n919_), .D(men_men_n335_), .Y(men_men_n1237_));
  NA2        u1209(.A(men_men_n45_), .B(f), .Y(men_men_n1238_));
  NA2        u1210(.A(men_men_n711_), .B(men_men_n98_), .Y(men_men_n1239_));
  NO2        u1211(.A(men_men_n1239_), .B(men_men_n1238_), .Y(men_men_n1240_));
  INV        u1212(.A(men_men_n118_), .Y(men_men_n1241_));
  OA220      u1213(.A0(men_men_n1241_), .A1(men_men_n594_), .B0(men_men_n660_), .B1(men_men_n374_), .Y(men_men_n1242_));
  NAi41      u1214(.An(men_men_n160_), .B(men_men_n1242_), .C(men_men_n1209_), .D(men_men_n902_), .Y(men_men_n1243_));
  NO3        u1215(.A(men_men_n784_), .B(men_men_n676_), .C(men_men_n518_), .Y(men_men_n1244_));
  OR2        u1216(.A(men_men_n197_), .B(men_men_n195_), .Y(men_men_n1245_));
  NA3        u1217(.A(men_men_n1245_), .B(men_men_n1244_), .C(men_men_n135_), .Y(men_men_n1246_));
  NO4        u1218(.A(men_men_n1246_), .B(men_men_n1243_), .C(men_men_n1237_), .D(men_men_n1233_), .Y(men_men_n1247_));
  INV        u1219(.A(men_men_n1183_), .Y(men_men_n1248_));
  NA2        u1220(.A(men_men_n1248_), .B(men_men_n538_), .Y(men_men_n1249_));
  NA2        u1221(.A(men_men_n544_), .B(men_men_n401_), .Y(men_men_n1250_));
  NOi21      u1222(.An(men_men_n570_), .B(men_men_n591_), .Y(men_men_n1251_));
  NA2        u1223(.A(men_men_n1251_), .B(men_men_n1250_), .Y(men_men_n1252_));
  AOI210     u1224(.A0(men_men_n206_), .A1(men_men_n91_), .B0(men_men_n214_), .Y(men_men_n1253_));
  OAI210     u1225(.A0(men_men_n812_), .A1(men_men_n433_), .B0(men_men_n1253_), .Y(men_men_n1254_));
  AN3        u1226(.A(m), .B(l), .C(k), .Y(men_men_n1255_));
  OAI210     u1227(.A0(men_men_n363_), .A1(men_men_n34_), .B0(men_men_n1255_), .Y(men_men_n1256_));
  NA2        u1228(.A(men_men_n205_), .B(men_men_n34_), .Y(men_men_n1257_));
  AO210      u1229(.A0(men_men_n1257_), .A1(men_men_n1256_), .B0(men_men_n334_), .Y(men_men_n1258_));
  NA4        u1230(.A(men_men_n1258_), .B(men_men_n1254_), .C(men_men_n1252_), .D(men_men_n1249_), .Y(men_men_n1259_));
  AOI210     u1231(.A0(men_men_n600_), .A1(men_men_n118_), .B0(men_men_n604_), .Y(men_men_n1260_));
  OAI210     u1232(.A0(men_men_n1241_), .A1(men_men_n599_), .B0(men_men_n1260_), .Y(men_men_n1261_));
  NA2        u1233(.A(men_men_n280_), .B(men_men_n197_), .Y(men_men_n1262_));
  NA2        u1234(.A(men_men_n1262_), .B(men_men_n665_), .Y(men_men_n1263_));
  NO3        u1235(.A(men_men_n820_), .B(men_men_n206_), .C(men_men_n413_), .Y(men_men_n1264_));
  NO2        u1236(.A(men_men_n1264_), .B(men_men_n963_), .Y(men_men_n1265_));
  OAI210     u1237(.A0(men_men_n1240_), .A1(men_men_n328_), .B0(men_men_n677_), .Y(men_men_n1266_));
  NA4        u1238(.A(men_men_n1266_), .B(men_men_n1265_), .C(men_men_n1263_), .D(men_men_n787_), .Y(men_men_n1267_));
  NO3        u1239(.A(men_men_n1267_), .B(men_men_n1261_), .C(men_men_n1259_), .Y(men_men_n1268_));
  NA3        u1240(.A(men_men_n607_), .B(men_men_n29_), .C(f), .Y(men_men_n1269_));
  NO2        u1241(.A(men_men_n1269_), .B(men_men_n206_), .Y(men_men_n1270_));
  AOI210     u1242(.A0(men_men_n510_), .A1(men_men_n58_), .B0(men_men_n1270_), .Y(men_men_n1271_));
  INV        u1243(.A(men_men_n1179_), .Y(men_men_n1272_));
  NA3        u1244(.A(men_men_n1272_), .B(men_men_n1271_), .C(men_men_n758_), .Y(men_men_n1273_));
  NO2        u1245(.A(men_men_n973_), .B(men_men_n234_), .Y(men_men_n1274_));
  NO2        u1246(.A(men_men_n974_), .B(men_men_n563_), .Y(men_men_n1275_));
  OAI210     u1247(.A0(men_men_n1275_), .A1(men_men_n1274_), .B0(men_men_n343_), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n579_), .B(men_men_n577_), .Y(men_men_n1277_));
  NO3        u1249(.A(men_men_n81_), .B(men_men_n301_), .C(men_men_n45_), .Y(men_men_n1278_));
  NA2        u1250(.A(men_men_n1278_), .B(men_men_n560_), .Y(men_men_n1279_));
  NA3        u1251(.A(men_men_n1279_), .B(men_men_n1277_), .C(men_men_n671_), .Y(men_men_n1280_));
  OR2        u1252(.A(men_men_n1183_), .B(men_men_n1176_), .Y(men_men_n1281_));
  NO2        u1253(.A(men_men_n374_), .B(men_men_n73_), .Y(men_men_n1282_));
  INV        u1254(.A(men_men_n1282_), .Y(men_men_n1283_));
  NA2        u1255(.A(men_men_n1278_), .B(men_men_n815_), .Y(men_men_n1284_));
  NA4        u1256(.A(men_men_n1284_), .B(men_men_n1283_), .C(men_men_n1281_), .D(men_men_n391_), .Y(men_men_n1285_));
  NOi41      u1257(.An(men_men_n1276_), .B(men_men_n1285_), .C(men_men_n1280_), .D(men_men_n1273_), .Y(men_men_n1286_));
  NO2        u1258(.A(men_men_n129_), .B(men_men_n45_), .Y(men_men_n1287_));
  NO2        u1259(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1288_));
  AO220      u1260(.A0(men_men_n1288_), .A1(men_men_n623_), .B0(men_men_n1287_), .B1(men_men_n709_), .Y(men_men_n1289_));
  NA2        u1261(.A(men_men_n1289_), .B(men_men_n343_), .Y(men_men_n1290_));
  NO3        u1262(.A(men_men_n1098_), .B(men_men_n177_), .C(men_men_n89_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n1278_), .B(men_men_n977_), .Y(men_men_n1292_));
  NA2        u1264(.A(men_men_n1292_), .B(men_men_n1290_), .Y(men_men_n1293_));
  NO2        u1265(.A(men_men_n614_), .B(men_men_n613_), .Y(men_men_n1294_));
  NO4        u1266(.A(men_men_n1098_), .B(men_men_n1294_), .C(men_men_n175_), .D(men_men_n89_), .Y(men_men_n1295_));
  NO3        u1267(.A(men_men_n1295_), .B(men_men_n1293_), .C(men_men_n636_), .Y(men_men_n1296_));
  NA4        u1268(.A(men_men_n1296_), .B(men_men_n1286_), .C(men_men_n1268_), .D(men_men_n1247_), .Y(men06));
  NO2        u1269(.A(men_men_n414_), .B(men_men_n567_), .Y(men_men_n1298_));
  INV        u1270(.A(men_men_n738_), .Y(men_men_n1299_));
  OAI210     u1271(.A0(men_men_n1299_), .A1(men_men_n266_), .B0(men_men_n1298_), .Y(men_men_n1300_));
  NO2        u1272(.A(men_men_n226_), .B(men_men_n104_), .Y(men_men_n1301_));
  OAI210     u1273(.A0(men_men_n1301_), .A1(men_men_n1291_), .B0(men_men_n387_), .Y(men_men_n1302_));
  NO3        u1274(.A(men_men_n603_), .B(men_men_n810_), .C(men_men_n605_), .Y(men_men_n1303_));
  OR2        u1275(.A(men_men_n1303_), .B(men_men_n890_), .Y(men_men_n1304_));
  NA4        u1276(.A(men_men_n1304_), .B(men_men_n1302_), .C(men_men_n1300_), .D(men_men_n1276_), .Y(men_men_n1305_));
  NO3        u1277(.A(men_men_n1305_), .B(men_men_n1280_), .C(men_men_n256_), .Y(men_men_n1306_));
  NO2        u1278(.A(men_men_n301_), .B(men_men_n45_), .Y(men_men_n1307_));
  AOI210     u1279(.A0(men_men_n1307_), .A1(men_men_n978_), .B0(men_men_n1274_), .Y(men_men_n1308_));
  AOI210     u1280(.A0(men_men_n1307_), .A1(men_men_n564_), .B0(men_men_n1289_), .Y(men_men_n1309_));
  AOI210     u1281(.A0(men_men_n1309_), .A1(men_men_n1308_), .B0(men_men_n340_), .Y(men_men_n1310_));
  INV        u1282(.A(men_men_n675_), .Y(men_men_n1311_));
  NA2        u1283(.A(men_men_n1311_), .B(men_men_n640_), .Y(men_men_n1312_));
  NO2        u1284(.A(men_men_n521_), .B(men_men_n172_), .Y(men_men_n1313_));
  NO2        u1285(.A(men_men_n610_), .B(men_men_n1122_), .Y(men_men_n1314_));
  OAI210     u1286(.A0(men_men_n466_), .A1(men_men_n249_), .B0(men_men_n913_), .Y(men_men_n1315_));
  NO3        u1287(.A(men_men_n1315_), .B(men_men_n1314_), .C(men_men_n1313_), .Y(men_men_n1316_));
  NO2        u1288(.A(men_men_n373_), .B(men_men_n134_), .Y(men_men_n1317_));
  AOI210     u1289(.A0(men_men_n1317_), .A1(men_men_n597_), .B0(men_men_n604_), .Y(men_men_n1318_));
  NA3        u1290(.A(men_men_n1318_), .B(men_men_n1316_), .C(men_men_n1312_), .Y(men_men_n1319_));
  NO2        u1291(.A(men_men_n751_), .B(men_men_n372_), .Y(men_men_n1320_));
  AN2        u1292(.A(men_men_n959_), .B(men_men_n643_), .Y(men_men_n1321_));
  NO3        u1293(.A(men_men_n1321_), .B(men_men_n1319_), .C(men_men_n1310_), .Y(men_men_n1322_));
  NO2        u1294(.A(men_men_n804_), .B(men_men_n276_), .Y(men_men_n1323_));
  OAI220     u1295(.A0(men_men_n738_), .A1(men_men_n47_), .B0(men_men_n226_), .B1(men_men_n616_), .Y(men_men_n1324_));
  AOI220     u1296(.A0(men_men_n366_), .A1(men_men_n1324_), .B0(men_men_n1323_), .B1(men_men_n266_), .Y(men_men_n1325_));
  NO3        u1297(.A(men_men_n246_), .B(men_men_n104_), .C(men_men_n283_), .Y(men_men_n1326_));
  OAI220     u1298(.A0(men_men_n702_), .A1(men_men_n249_), .B0(men_men_n517_), .B1(men_men_n521_), .Y(men_men_n1327_));
  NO3        u1299(.A(men_men_n1327_), .B(men_men_n1326_), .C(men_men_n1125_), .Y(men_men_n1328_));
  NA4        u1300(.A(men_men_n795_), .B(men_men_n794_), .C(men_men_n443_), .D(men_men_n882_), .Y(men_men_n1329_));
  NAi31      u1301(.An(men_men_n751_), .B(men_men_n1329_), .C(men_men_n205_), .Y(men_men_n1330_));
  NA4        u1302(.A(men_men_n1330_), .B(men_men_n1328_), .C(men_men_n1325_), .D(men_men_n1221_), .Y(men_men_n1331_));
  NOi31      u1303(.An(men_men_n1303_), .B(men_men_n470_), .C(men_men_n400_), .Y(men_men_n1332_));
  OR3        u1304(.A(men_men_n1332_), .B(men_men_n783_), .C(men_men_n547_), .Y(men_men_n1333_));
  OR3        u1305(.A(men_men_n375_), .B(men_men_n226_), .C(men_men_n616_), .Y(men_men_n1334_));
  AOI210     u1306(.A0(men_men_n579_), .A1(men_men_n455_), .B0(men_men_n377_), .Y(men_men_n1335_));
  NA3        u1307(.A(men_men_n1335_), .B(men_men_n1334_), .C(men_men_n1333_), .Y(men_men_n1336_));
  AOI220     u1308(.A0(men_men_n1320_), .A1(men_men_n759_), .B0(men_men_n1317_), .B1(men_men_n240_), .Y(men_men_n1337_));
  AN2        u1309(.A(men_men_n933_), .B(men_men_n932_), .Y(men_men_n1338_));
  NO4        u1310(.A(men_men_n1338_), .B(men_men_n880_), .C(men_men_n506_), .D(men_men_n488_), .Y(men_men_n1339_));
  NA3        u1311(.A(men_men_n1339_), .B(men_men_n1337_), .C(men_men_n1284_), .Y(men_men_n1340_));
  NAi21      u1312(.An(j), .B(i), .Y(men_men_n1341_));
  NO4        u1313(.A(men_men_n1294_), .B(men_men_n1341_), .C(men_men_n449_), .D(men_men_n237_), .Y(men_men_n1342_));
  NO4        u1314(.A(men_men_n1342_), .B(men_men_n1340_), .C(men_men_n1336_), .D(men_men_n1331_), .Y(men_men_n1343_));
  NA4        u1315(.A(men_men_n1343_), .B(men_men_n1322_), .C(men_men_n1306_), .D(men_men_n1296_), .Y(men07));
  NOi21      u1316(.An(j), .B(k), .Y(men_men_n1345_));
  NA4        u1317(.A(men_men_n180_), .B(men_men_n110_), .C(men_men_n1345_), .D(f), .Y(men_men_n1346_));
  NAi32      u1318(.An(m), .Bn(b), .C(n), .Y(men_men_n1347_));
  NO3        u1319(.A(men_men_n1347_), .B(g), .C(f), .Y(men_men_n1348_));
  OAI210     u1320(.A0(men_men_n323_), .A1(men_men_n490_), .B0(men_men_n1348_), .Y(men_men_n1349_));
  NAi21      u1321(.An(f), .B(c), .Y(men_men_n1350_));
  OR2        u1322(.A(e), .B(d), .Y(men_men_n1351_));
  OAI220     u1323(.A0(men_men_n1351_), .A1(men_men_n1350_), .B0(men_men_n629_), .B1(men_men_n324_), .Y(men_men_n1352_));
  NA3        u1324(.A(men_men_n1352_), .B(men_men_n1062_), .C(men_men_n180_), .Y(men_men_n1353_));
  NOi31      u1325(.An(n), .B(m), .C(b), .Y(men_men_n1354_));
  NO3        u1326(.A(men_men_n130_), .B(men_men_n456_), .C(h), .Y(men_men_n1355_));
  NA3        u1327(.A(men_men_n1353_), .B(men_men_n1349_), .C(men_men_n1346_), .Y(men_men_n1356_));
  NOi41      u1328(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1357_));
  NA3        u1329(.A(men_men_n1357_), .B(men_men_n872_), .C(men_men_n416_), .Y(men_men_n1358_));
  NO2        u1330(.A(men_men_n1358_), .B(men_men_n56_), .Y(men_men_n1359_));
  NA2        u1331(.A(men_men_n1100_), .B(men_men_n222_), .Y(men_men_n1360_));
  NO2        u1332(.A(men_men_n1360_), .B(men_men_n61_), .Y(men_men_n1361_));
  NO2        u1333(.A(k), .B(i), .Y(men_men_n1362_));
  NA3        u1334(.A(men_men_n1362_), .B(men_men_n901_), .C(men_men_n180_), .Y(men_men_n1363_));
  NA2        u1335(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1364_));
  NO2        u1336(.A(men_men_n1056_), .B(men_men_n449_), .Y(men_men_n1365_));
  NA3        u1337(.A(men_men_n1365_), .B(men_men_n1364_), .C(men_men_n215_), .Y(men_men_n1366_));
  NO2        u1338(.A(men_men_n1070_), .B(men_men_n307_), .Y(men_men_n1367_));
  NA2        u1339(.A(men_men_n548_), .B(men_men_n82_), .Y(men_men_n1368_));
  NA2        u1340(.A(men_men_n1222_), .B(men_men_n291_), .Y(men_men_n1369_));
  NA4        u1341(.A(men_men_n1369_), .B(men_men_n1368_), .C(men_men_n1366_), .D(men_men_n1363_), .Y(men_men_n1370_));
  NO4        u1342(.A(men_men_n1370_), .B(men_men_n1361_), .C(men_men_n1359_), .D(men_men_n1356_), .Y(men_men_n1371_));
  NO3        u1343(.A(e), .B(d), .C(c), .Y(men_men_n1372_));
  NO2        u1344(.A(men_men_n130_), .B(men_men_n215_), .Y(men_men_n1373_));
  NA2        u1345(.A(men_men_n1373_), .B(men_men_n1372_), .Y(men_men_n1374_));
  NO2        u1346(.A(men_men_n1374_), .B(c), .Y(men_men_n1375_));
  OR2        u1347(.A(h), .B(f), .Y(men_men_n1376_));
  NO3        u1348(.A(n), .B(m), .C(i), .Y(men_men_n1377_));
  OAI210     u1349(.A0(men_men_n1123_), .A1(men_men_n155_), .B0(men_men_n1377_), .Y(men_men_n1378_));
  NO2        u1350(.A(i), .B(g), .Y(men_men_n1379_));
  OR3        u1351(.A(men_men_n1379_), .B(men_men_n1347_), .C(men_men_n72_), .Y(men_men_n1380_));
  OAI220     u1352(.A0(men_men_n1380_), .A1(men_men_n490_), .B0(men_men_n1378_), .B1(men_men_n1376_), .Y(men_men_n1381_));
  NA3        u1353(.A(men_men_n699_), .B(men_men_n685_), .C(men_men_n113_), .Y(men_men_n1382_));
  NA3        u1354(.A(men_men_n1354_), .B(men_men_n1065_), .C(men_men_n673_), .Y(men_men_n1383_));
  AOI210     u1355(.A0(men_men_n1383_), .A1(men_men_n1382_), .B0(men_men_n45_), .Y(men_men_n1384_));
  NA2        u1356(.A(men_men_n1377_), .B(men_men_n638_), .Y(men_men_n1385_));
  NO2        u1357(.A(l), .B(k), .Y(men_men_n1386_));
  NOi41      u1358(.An(men_men_n553_), .B(men_men_n1386_), .C(men_men_n485_), .D(men_men_n449_), .Y(men_men_n1387_));
  NO3        u1359(.A(men_men_n449_), .B(d), .C(c), .Y(men_men_n1388_));
  NO4        u1360(.A(men_men_n1387_), .B(men_men_n1384_), .C(men_men_n1381_), .D(men_men_n1375_), .Y(men_men_n1389_));
  NO2        u1361(.A(men_men_n145_), .B(h), .Y(men_men_n1390_));
  NO2        u1362(.A(men_men_n1080_), .B(l), .Y(men_men_n1391_));
  NO2        u1363(.A(g), .B(c), .Y(men_men_n1392_));
  NA3        u1364(.A(men_men_n1392_), .B(men_men_n140_), .C(men_men_n188_), .Y(men_men_n1393_));
  NO2        u1365(.A(men_men_n1393_), .B(men_men_n1391_), .Y(men_men_n1394_));
  NA2        u1366(.A(men_men_n1394_), .B(men_men_n180_), .Y(men_men_n1395_));
  NO2        u1367(.A(men_men_n457_), .B(a), .Y(men_men_n1396_));
  NA3        u1368(.A(men_men_n1396_), .B(k), .C(men_men_n114_), .Y(men_men_n1397_));
  NO2        u1369(.A(i), .B(h), .Y(men_men_n1398_));
  AOI210     u1370(.A0(men_men_n1147_), .A1(h), .B0(men_men_n421_), .Y(men_men_n1399_));
  NA2        u1371(.A(men_men_n136_), .B(men_men_n222_), .Y(men_men_n1400_));
  NO2        u1372(.A(men_men_n1400_), .B(men_men_n1399_), .Y(men_men_n1401_));
  NO2        u1373(.A(men_men_n756_), .B(men_men_n189_), .Y(men_men_n1402_));
  NOi31      u1374(.An(m), .B(n), .C(b), .Y(men_men_n1403_));
  NOi31      u1375(.An(f), .B(d), .C(c), .Y(men_men_n1404_));
  NA2        u1376(.A(men_men_n1404_), .B(men_men_n1403_), .Y(men_men_n1405_));
  INV        u1377(.A(men_men_n1405_), .Y(men_men_n1406_));
  NO3        u1378(.A(men_men_n1406_), .B(men_men_n1402_), .C(men_men_n1401_), .Y(men_men_n1407_));
  NA2        u1379(.A(men_men_n1091_), .B(men_men_n473_), .Y(men_men_n1408_));
  NO4        u1380(.A(men_men_n1408_), .B(men_men_n1065_), .C(men_men_n449_), .D(men_men_n45_), .Y(men_men_n1409_));
  OAI210     u1381(.A0(men_men_n183_), .A1(men_men_n533_), .B0(men_men_n1066_), .Y(men_men_n1410_));
  NO3        u1382(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1411_));
  INV        u1383(.A(men_men_n1410_), .Y(men_men_n1412_));
  NO2        u1384(.A(men_men_n1412_), .B(men_men_n1409_), .Y(men_men_n1413_));
  AN4        u1385(.A(men_men_n1413_), .B(men_men_n1407_), .C(men_men_n1397_), .D(men_men_n1395_), .Y(men_men_n1414_));
  NA2        u1386(.A(men_men_n1354_), .B(men_men_n384_), .Y(men_men_n1415_));
  NO2        u1387(.A(men_men_n1415_), .B(men_men_n1047_), .Y(men_men_n1416_));
  NA2        u1388(.A(men_men_n1388_), .B(men_men_n216_), .Y(men_men_n1417_));
  NO2        u1389(.A(men_men_n189_), .B(b), .Y(men_men_n1418_));
  AOI220     u1390(.A0(men_men_n1177_), .A1(men_men_n1418_), .B0(men_men_n1099_), .B1(men_men_n1408_), .Y(men_men_n1419_));
  NO2        u1391(.A(i), .B(men_men_n214_), .Y(men_men_n1420_));
  NA4        u1392(.A(men_men_n1153_), .B(men_men_n1420_), .C(men_men_n105_), .D(m), .Y(men_men_n1421_));
  NAi41      u1393(.An(men_men_n1416_), .B(men_men_n1421_), .C(men_men_n1419_), .D(men_men_n1417_), .Y(men_men_n1422_));
  NO4        u1394(.A(men_men_n130_), .B(g), .C(f), .D(e), .Y(men_men_n1423_));
  NA3        u1395(.A(men_men_n1362_), .B(men_men_n292_), .C(h), .Y(men_men_n1424_));
  NA2        u1396(.A(men_men_n196_), .B(men_men_n100_), .Y(men_men_n1425_));
  OR2        u1397(.A(e), .B(a), .Y(men_men_n1426_));
  NO2        u1398(.A(men_men_n1351_), .B(men_men_n1350_), .Y(men_men_n1427_));
  AOI210     u1399(.A0(men_men_n30_), .A1(h), .B0(men_men_n1427_), .Y(men_men_n1428_));
  NO2        u1400(.A(men_men_n1428_), .B(men_men_n1087_), .Y(men_men_n1429_));
  NOi41      u1401(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1430_));
  NA2        u1402(.A(men_men_n1430_), .B(men_men_n114_), .Y(men_men_n1431_));
  NA2        u1403(.A(men_men_n1357_), .B(men_men_n1386_), .Y(men_men_n1432_));
  NA2        u1404(.A(men_men_n1432_), .B(men_men_n1431_), .Y(men_men_n1433_));
  NA2        u1405(.A(men_men_n1121_), .B(men_men_n413_), .Y(men_men_n1434_));
  NO2        u1406(.A(men_men_n1434_), .B(men_men_n442_), .Y(men_men_n1435_));
  AO210      u1407(.A0(men_men_n1435_), .A1(men_men_n116_), .B0(men_men_n1433_), .Y(men_men_n1436_));
  NO3        u1408(.A(men_men_n1436_), .B(men_men_n1429_), .C(men_men_n1422_), .Y(men_men_n1437_));
  NA4        u1409(.A(men_men_n1437_), .B(men_men_n1414_), .C(men_men_n1389_), .D(men_men_n1371_), .Y(men_men_n1438_));
  NA2        u1410(.A(men_men_n384_), .B(men_men_n56_), .Y(men_men_n1439_));
  AOI210     u1411(.A0(men_men_n1439_), .A1(men_men_n1056_), .B0(men_men_n1385_), .Y(men_men_n1440_));
  NA2        u1412(.A(men_men_n216_), .B(men_men_n180_), .Y(men_men_n1441_));
  AOI210     u1413(.A0(men_men_n1441_), .A1(men_men_n1195_), .B0(men_men_n1439_), .Y(men_men_n1442_));
  NO2        u1414(.A(men_men_n1092_), .B(men_men_n1087_), .Y(men_men_n1443_));
  NO3        u1415(.A(men_men_n1443_), .B(men_men_n1442_), .C(men_men_n1440_), .Y(men_men_n1444_));
  NO2        u1416(.A(men_men_n396_), .B(j), .Y(men_men_n1445_));
  NA3        u1417(.A(men_men_n1411_), .B(men_men_n1351_), .C(men_men_n1121_), .Y(men_men_n1446_));
  NAi41      u1418(.An(men_men_n1398_), .B(men_men_n1078_), .C(men_men_n168_), .D(men_men_n148_), .Y(men_men_n1447_));
  NA2        u1419(.A(men_men_n1447_), .B(men_men_n1446_), .Y(men_men_n1448_));
  NA3        u1420(.A(g), .B(men_men_n1445_), .C(men_men_n157_), .Y(men_men_n1449_));
  INV        u1421(.A(men_men_n1449_), .Y(men_men_n1450_));
  NO3        u1422(.A(men_men_n751_), .B(men_men_n175_), .C(men_men_n416_), .Y(men_men_n1451_));
  NO3        u1423(.A(men_men_n1451_), .B(men_men_n1450_), .C(men_men_n1448_), .Y(men_men_n1452_));
  NO3        u1424(.A(men_men_n1087_), .B(men_men_n591_), .C(g), .Y(men_men_n1453_));
  NOi21      u1425(.An(men_men_n1441_), .B(men_men_n1453_), .Y(men_men_n1454_));
  AOI210     u1426(.A0(men_men_n1454_), .A1(men_men_n1425_), .B0(men_men_n1056_), .Y(men_men_n1455_));
  OR2        u1427(.A(n), .B(i), .Y(men_men_n1456_));
  OAI210     u1428(.A0(men_men_n1456_), .A1(men_men_n1077_), .B0(men_men_n49_), .Y(men_men_n1457_));
  AOI220     u1429(.A0(men_men_n1457_), .A1(men_men_n1185_), .B0(men_men_n824_), .B1(men_men_n196_), .Y(men_men_n1458_));
  INV        u1430(.A(men_men_n1458_), .Y(men_men_n1459_));
  NA2        u1431(.A(men_men_n1418_), .B(men_men_n41_), .Y(men_men_n1460_));
  NO2        u1432(.A(men_men_n130_), .B(l), .Y(men_men_n1461_));
  NO2        u1433(.A(men_men_n226_), .B(k), .Y(men_men_n1462_));
  OAI210     u1434(.A0(men_men_n1462_), .A1(men_men_n1398_), .B0(men_men_n1461_), .Y(men_men_n1463_));
  OAI220     u1435(.A0(men_men_n1463_), .A1(men_men_n31_), .B0(men_men_n1460_), .B1(men_men_n177_), .Y(men_men_n1464_));
  NO3        u1436(.A(men_men_n1464_), .B(men_men_n1459_), .C(men_men_n1455_), .Y(men_men_n1465_));
  INV        u1437(.A(men_men_n49_), .Y(men_men_n1466_));
  NO3        u1438(.A(men_men_n1102_), .B(men_men_n1351_), .C(men_men_n49_), .Y(men_men_n1467_));
  NA2        u1439(.A(men_men_n1103_), .B(men_men_n1466_), .Y(men_men_n1468_));
  NO2        u1440(.A(men_men_n1087_), .B(h), .Y(men_men_n1469_));
  NA3        u1441(.A(men_men_n1469_), .B(d), .C(men_men_n1048_), .Y(men_men_n1470_));
  OAI220     u1442(.A0(men_men_n1470_), .A1(c), .B0(men_men_n1468_), .B1(j), .Y(men_men_n1471_));
  NA2        u1443(.A(men_men_n180_), .B(men_men_n113_), .Y(men_men_n1472_));
  AOI210     u1444(.A0(men_men_n533_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1473_));
  NA2        u1445(.A(men_men_n1473_), .B(men_men_n1396_), .Y(men_men_n1474_));
  NO2        u1446(.A(men_men_n1341_), .B(men_men_n175_), .Y(men_men_n1475_));
  NOi21      u1447(.An(d), .B(f), .Y(men_men_n1476_));
  NO3        u1448(.A(men_men_n1404_), .B(men_men_n1476_), .C(men_men_n40_), .Y(men_men_n1477_));
  NA2        u1449(.A(men_men_n1477_), .B(men_men_n1475_), .Y(men_men_n1478_));
  NO2        u1450(.A(men_men_n1351_), .B(f), .Y(men_men_n1479_));
  NO2        u1451(.A(men_men_n301_), .B(c), .Y(men_men_n1480_));
  NA2        u1452(.A(men_men_n1480_), .B(men_men_n548_), .Y(men_men_n1481_));
  NA3        u1453(.A(men_men_n1481_), .B(men_men_n1478_), .C(men_men_n1474_), .Y(men_men_n1482_));
  NO2        u1454(.A(men_men_n1482_), .B(men_men_n1471_), .Y(men_men_n1483_));
  NA4        u1455(.A(men_men_n1483_), .B(men_men_n1465_), .C(men_men_n1452_), .D(men_men_n1444_), .Y(men_men_n1484_));
  NO3        u1456(.A(men_men_n1091_), .B(men_men_n1077_), .C(men_men_n40_), .Y(men_men_n1485_));
  NO2        u1457(.A(men_men_n473_), .B(men_men_n301_), .Y(men_men_n1486_));
  OAI210     u1458(.A0(men_men_n1486_), .A1(men_men_n1485_), .B0(men_men_n1367_), .Y(men_men_n1487_));
  OAI210     u1459(.A0(men_men_n1423_), .A1(men_men_n1354_), .B0(men_men_n887_), .Y(men_men_n1488_));
  NO2        u1460(.A(men_men_n1044_), .B(men_men_n130_), .Y(men_men_n1489_));
  NA2        u1461(.A(men_men_n1489_), .B(men_men_n622_), .Y(men_men_n1490_));
  NA3        u1462(.A(men_men_n1490_), .B(men_men_n1488_), .C(men_men_n1487_), .Y(men_men_n1491_));
  NA2        u1463(.A(men_men_n1392_), .B(men_men_n1476_), .Y(men_men_n1492_));
  NO2        u1464(.A(men_men_n1492_), .B(m), .Y(men_men_n1493_));
  NA3        u1465(.A(men_men_n1100_), .B(men_men_n110_), .C(men_men_n222_), .Y(men_men_n1494_));
  NO2        u1466(.A(men_men_n149_), .B(men_men_n182_), .Y(men_men_n1495_));
  OAI210     u1467(.A0(men_men_n1495_), .A1(men_men_n111_), .B0(men_men_n1403_), .Y(men_men_n1496_));
  NA2        u1468(.A(men_men_n1496_), .B(men_men_n1494_), .Y(men_men_n1497_));
  NO3        u1469(.A(men_men_n1497_), .B(men_men_n1493_), .C(men_men_n1491_), .Y(men_men_n1498_));
  NO2        u1470(.A(men_men_n1350_), .B(e), .Y(men_men_n1499_));
  NA2        u1471(.A(men_men_n1499_), .B(men_men_n411_), .Y(men_men_n1500_));
  OAI210     u1472(.A0(men_men_n1479_), .A1(men_men_n1132_), .B0(men_men_n632_), .Y(men_men_n1501_));
  OR3        u1473(.A(men_men_n1462_), .B(men_men_n1222_), .C(men_men_n130_), .Y(men_men_n1502_));
  OAI220     u1474(.A0(men_men_n1502_), .A1(men_men_n1500_), .B0(men_men_n1501_), .B1(men_men_n451_), .Y(men_men_n1503_));
  INV        u1475(.A(men_men_n1503_), .Y(men_men_n1504_));
  NO2        u1476(.A(men_men_n182_), .B(c), .Y(men_men_n1505_));
  OAI210     u1477(.A0(men_men_n1505_), .A1(men_men_n1499_), .B0(men_men_n180_), .Y(men_men_n1506_));
  AOI220     u1478(.A0(men_men_n1506_), .A1(men_men_n1079_), .B0(men_men_n540_), .B1(men_men_n372_), .Y(men_men_n1507_));
  NA2        u1479(.A(men_men_n546_), .B(g), .Y(men_men_n1508_));
  AOI210     u1480(.A0(men_men_n1508_), .A1(men_men_n1388_), .B0(men_men_n1467_), .Y(men_men_n1509_));
  NA2        u1481(.A(men_men_n1132_), .B(a), .Y(men_men_n1510_));
  OAI220     u1482(.A0(men_men_n1510_), .A1(men_men_n69_), .B0(men_men_n1509_), .B1(men_men_n214_), .Y(men_men_n1511_));
  AOI210     u1483(.A0(men_men_n906_), .A1(men_men_n423_), .B0(men_men_n106_), .Y(men_men_n1512_));
  OR2        u1484(.A(men_men_n1512_), .B(men_men_n546_), .Y(men_men_n1513_));
  NO2        u1485(.A(men_men_n1513_), .B(men_men_n175_), .Y(men_men_n1514_));
  NA4        u1486(.A(men_men_n1100_), .B(men_men_n1097_), .C(men_men_n222_), .D(men_men_n68_), .Y(men_men_n1515_));
  NA2        u1487(.A(men_men_n1355_), .B(men_men_n183_), .Y(men_men_n1516_));
  NO2        u1488(.A(men_men_n49_), .B(l), .Y(men_men_n1517_));
  OAI210     u1489(.A0(men_men_n1426_), .A1(men_men_n864_), .B0(men_men_n490_), .Y(men_men_n1518_));
  OAI210     u1490(.A0(men_men_n1518_), .A1(men_men_n1103_), .B0(men_men_n1517_), .Y(men_men_n1519_));
  NO2        u1491(.A(men_men_n252_), .B(g), .Y(men_men_n1520_));
  NO2        u1492(.A(m), .B(i), .Y(men_men_n1521_));
  BUFFER     u1493(.A(men_men_n1521_), .Y(men_men_n1522_));
  AOI220     u1494(.A0(men_men_n1522_), .A1(men_men_n1390_), .B0(men_men_n1078_), .B1(men_men_n1520_), .Y(men_men_n1523_));
  NA4        u1495(.A(men_men_n1523_), .B(men_men_n1519_), .C(men_men_n1516_), .D(men_men_n1515_), .Y(men_men_n1524_));
  NO4        u1496(.A(men_men_n1524_), .B(men_men_n1514_), .C(men_men_n1511_), .D(men_men_n1507_), .Y(men_men_n1525_));
  NA3        u1497(.A(men_men_n1525_), .B(men_men_n1504_), .C(men_men_n1498_), .Y(men_men_n1526_));
  NA3        u1498(.A(men_men_n965_), .B(men_men_n136_), .C(men_men_n46_), .Y(men_men_n1527_));
  AOI210     u1499(.A0(men_men_n146_), .A1(c), .B0(men_men_n1527_), .Y(men_men_n1528_));
  INV        u1500(.A(men_men_n186_), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n1529_), .B(men_men_n1469_), .Y(men_men_n1530_));
  OR2        u1502(.A(men_men_n131_), .B(men_men_n1415_), .Y(men_men_n1531_));
  NO2        u1503(.A(men_men_n72_), .B(c), .Y(men_men_n1532_));
  NO4        u1504(.A(men_men_n1376_), .B(men_men_n187_), .C(men_men_n456_), .D(men_men_n45_), .Y(men_men_n1533_));
  AOI210     u1505(.A0(men_men_n1475_), .A1(men_men_n1532_), .B0(men_men_n1533_), .Y(men_men_n1534_));
  NA3        u1506(.A(men_men_n1534_), .B(men_men_n1531_), .C(men_men_n1530_), .Y(men_men_n1535_));
  NO2        u1507(.A(men_men_n1535_), .B(men_men_n1528_), .Y(men_men_n1536_));
  NO4        u1508(.A(men_men_n226_), .B(men_men_n187_), .C(men_men_n257_), .D(k), .Y(men_men_n1537_));
  AOI210     u1509(.A0(men_men_n155_), .A1(men_men_n56_), .B0(men_men_n1499_), .Y(men_men_n1538_));
  NO2        u1510(.A(men_men_n1538_), .B(men_men_n1472_), .Y(men_men_n1539_));
  NO2        u1511(.A(men_men_n1527_), .B(men_men_n111_), .Y(men_men_n1540_));
  NOi21      u1512(.An(men_men_n1355_), .B(e), .Y(men_men_n1541_));
  NO4        u1513(.A(men_men_n1541_), .B(men_men_n1540_), .C(men_men_n1539_), .D(men_men_n1537_), .Y(men_men_n1542_));
  AN2        u1514(.A(men_men_n1100_), .B(men_men_n1085_), .Y(men_men_n1543_));
  AOI220     u1515(.A0(men_men_n1521_), .A1(men_men_n638_), .B0(men_men_n1062_), .B1(men_men_n158_), .Y(men_men_n1544_));
  NOi31      u1516(.An(men_men_n30_), .B(men_men_n1544_), .C(n), .Y(men_men_n1545_));
  AOI210     u1517(.A0(men_men_n1543_), .A1(men_men_n1177_), .B0(men_men_n1545_), .Y(men_men_n1546_));
  NA2        u1518(.A(men_men_n59_), .B(a), .Y(men_men_n1547_));
  NO2        u1519(.A(men_men_n1362_), .B(men_men_n118_), .Y(men_men_n1548_));
  OAI220     u1520(.A0(men_men_n1548_), .A1(men_men_n1415_), .B0(men_men_n1434_), .B1(men_men_n1547_), .Y(men_men_n1549_));
  INV        u1521(.A(men_men_n1549_), .Y(men_men_n1550_));
  NA4        u1522(.A(men_men_n1550_), .B(men_men_n1546_), .C(men_men_n1542_), .D(men_men_n1536_), .Y(men_men_n1551_));
  OR4        u1523(.A(men_men_n1551_), .B(men_men_n1526_), .C(men_men_n1484_), .D(men_men_n1438_), .Y(men04));
  NOi31      u1524(.An(men_men_n1423_), .B(men_men_n1424_), .C(men_men_n1050_), .Y(men_men_n1553_));
  NA2        u1525(.A(men_men_n1479_), .B(men_men_n824_), .Y(men_men_n1554_));
  NO4        u1526(.A(men_men_n1554_), .B(men_men_n1039_), .C(men_men_n491_), .D(j), .Y(men_men_n1555_));
  OR3        u1527(.A(men_men_n1555_), .B(men_men_n1553_), .C(men_men_n1068_), .Y(men_men_n1556_));
  NO3        u1528(.A(men_men_n1364_), .B(men_men_n93_), .C(k), .Y(men_men_n1557_));
  AOI210     u1529(.A0(men_men_n1557_), .A1(men_men_n1061_), .B0(men_men_n1197_), .Y(men_men_n1558_));
  NA2        u1530(.A(men_men_n1558_), .B(men_men_n1226_), .Y(men_men_n1559_));
  NO4        u1531(.A(men_men_n1559_), .B(men_men_n1556_), .C(men_men_n1076_), .D(men_men_n1055_), .Y(men_men_n1560_));
  NA4        u1532(.A(men_men_n1560_), .B(men_men_n1134_), .C(men_men_n1119_), .D(men_men_n1106_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule