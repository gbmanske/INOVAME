//Benchmark atmr_intb_466_0.125

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n302_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n329_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n345_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO2        o027(.A(ori_ori_n49_), .B(x11), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x07), .Y(ori_ori_n54_));
  OAI210     o032(.A0(ori_ori_n54_), .A1(ori_ori_n50_), .B0(ori_ori_n47_), .Y(ori_ori_n55_));
  NOi21      o033(.An(x01), .B(x09), .Y(ori_ori_n56_));
  INV        o034(.A(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n51_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(x09), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o038(.A(x07), .Y(ori_ori_n61_));
  AOI220     o039(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n61_), .Y(ori_ori_n62_));
  INV        o040(.A(ori_ori_n59_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n64_), .B(ori_ori_n24_), .Y(ori_ori_n65_));
  OAI220     o043(.A0(ori_ori_n65_), .A1(ori_ori_n63_), .B0(ori_ori_n62_), .B1(ori_ori_n60_), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n61_), .B(ori_ori_n48_), .Y(ori_ori_n67_));
  OAI210     o045(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n67_), .Y(ori_ori_n68_));
  AOI220     o046(.A0(ori_ori_n68_), .A1(ori_ori_n59_), .B0(ori_ori_n66_), .B1(ori_ori_n31_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(ori_ori_n69_), .A1(ori_ori_n55_), .B0(x05), .Y(ori_ori_n70_));
  INV        o048(.A(x10), .Y(ori_ori_n71_));
  NA2        o049(.A(x09), .B(x05), .Y(ori_ori_n72_));
  NA2        o050(.A(x10), .B(x06), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n61_), .B(ori_ori_n41_), .Y(ori_ori_n74_));
  NA2        o052(.A(x07), .B(x03), .Y(ori_ori_n75_));
  NOi31      o053(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n76_));
  INV        o054(.A(x07), .Y(ori_ori_n77_));
  NO2        o055(.A(ori_ori_n77_), .B(ori_ori_n24_), .Y(ori_ori_n78_));
  NO2        o056(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n79_), .B(ori_ori_n36_), .Y(ori_ori_n80_));
  OAI210     o058(.A0(ori_ori_n79_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n81_));
  AOI210     o059(.A0(ori_ori_n80_), .A1(ori_ori_n48_), .B0(ori_ori_n81_), .Y(ori_ori_n82_));
  NO2        o060(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n83_));
  NO2        o061(.A(x08), .B(x01), .Y(ori_ori_n84_));
  OAI210     o062(.A0(ori_ori_n84_), .A1(ori_ori_n83_), .B0(ori_ori_n35_), .Y(ori_ori_n85_));
  NO3        o063(.A(ori_ori_n85_), .B(ori_ori_n82_), .C(ori_ori_n78_), .Y(ori_ori_n86_));
  AN2        o064(.A(ori_ori_n86_), .B(ori_ori_n75_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n85_), .Y(ori_ori_n88_));
  NA2        o066(.A(x11), .B(x00), .Y(ori_ori_n89_));
  NO2        o067(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n90_));
  NOi21      o068(.An(ori_ori_n89_), .B(ori_ori_n90_), .Y(ori_ori_n91_));
  NOi21      o069(.An(x01), .B(x10), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n29_), .B(ori_ori_n57_), .Y(ori_ori_n93_));
  NO3        o071(.A(ori_ori_n93_), .B(ori_ori_n92_), .C(x06), .Y(ori_ori_n94_));
  NA2        o072(.A(ori_ori_n94_), .B(ori_ori_n27_), .Y(ori_ori_n95_));
  OAI210     o073(.A0(ori_ori_n352_), .A1(x07), .B0(ori_ori_n95_), .Y(ori_ori_n96_));
  NO3        o074(.A(ori_ori_n96_), .B(ori_ori_n87_), .C(ori_ori_n70_), .Y(ori01));
  INV        o075(.A(x12), .Y(ori_ori_n98_));
  INV        o076(.A(x13), .Y(ori_ori_n99_));
  NO2        o077(.A(x10), .B(x01), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  NO2        o080(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n103_));
  INV        o081(.A(x13), .Y(ori_ori_n104_));
  NA2        o082(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n105_));
  NO2        o083(.A(ori_ori_n105_), .B(x05), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n35_), .B(ori_ori_n57_), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n108_));
  NA2        o086(.A(x10), .B(ori_ori_n57_), .Y(ori_ori_n109_));
  NA2        o087(.A(ori_ori_n109_), .B(ori_ori_n108_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n112_));
  NA3        o090(.A(ori_ori_n112_), .B(ori_ori_n111_), .C(x13), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n114_));
  NOi31      o092(.An(ori_ori_n113_), .B(ori_ori_n114_), .C(ori_ori_n110_), .Y(ori_ori_n115_));
  NO3        o093(.A(ori_ori_n115_), .B(x06), .C(x03), .Y(ori_ori_n116_));
  INV        o094(.A(ori_ori_n116_), .Y(ori_ori_n117_));
  NA2        o095(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n118_));
  OAI210     o096(.A0(ori_ori_n84_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n119_));
  NO2        o097(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n121_));
  NO2        o099(.A(x09), .B(x05), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n122_), .B(ori_ori_n47_), .Y(ori_ori_n123_));
  AOI210     o101(.A0(ori_ori_n123_), .A1(ori_ori_n102_), .B0(ori_ori_n49_), .Y(ori_ori_n124_));
  NA2        o102(.A(x09), .B(x00), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n103_), .B(ori_ori_n125_), .Y(ori_ori_n126_));
  INV        o104(.A(ori_ori_n124_), .Y(ori_ori_n127_));
  NO2        o105(.A(x03), .B(x02), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n85_), .B(ori_ori_n99_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n129_), .B(ori_ori_n128_), .Y(ori_ori_n130_));
  OA210      o108(.A0(ori_ori_n127_), .A1(x11), .B0(ori_ori_n130_), .Y(ori_ori_n131_));
  OAI210     o109(.A0(ori_ori_n117_), .A1(ori_ori_n23_), .B0(ori_ori_n131_), .Y(ori_ori_n132_));
  NAi21      o110(.An(x06), .B(x10), .Y(ori_ori_n133_));
  NOi21      o111(.An(x01), .B(x13), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n134_), .B(ori_ori_n133_), .Y(ori_ori_n135_));
  NO2        o113(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n99_), .B(x01), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n137_), .B(x08), .Y(ori_ori_n138_));
  OAI210     o116(.A0(x05), .A1(ori_ori_n138_), .B0(ori_ori_n51_), .Y(ori_ori_n139_));
  AOI210     o117(.A0(ori_ori_n139_), .A1(ori_ori_n136_), .B0(ori_ori_n48_), .Y(ori_ori_n140_));
  AOI210     o118(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n141_));
  NA2        o119(.A(ori_ori_n140_), .B(ori_ori_n141_), .Y(ori_ori_n142_));
  NA2        o120(.A(x10), .B(x05), .Y(ori_ori_n143_));
  NO2        o121(.A(x09), .B(x01), .Y(ori_ori_n144_));
  INV        o122(.A(ori_ori_n25_), .Y(ori_ori_n145_));
  NAi21      o123(.An(x13), .B(x00), .Y(ori_ori_n146_));
  AN2        o124(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n93_), .B(x06), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n146_), .B(ori_ori_n36_), .Y(ori_ori_n149_));
  INV        o127(.A(ori_ori_n149_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n148_), .B(ori_ori_n147_), .Y(ori_ori_n151_));
  NA2        o129(.A(ori_ori_n151_), .B(ori_ori_n145_), .Y(ori_ori_n152_));
  NOi21      o130(.An(x09), .B(x00), .Y(ori_ori_n153_));
  NO3        o131(.A(ori_ori_n83_), .B(ori_ori_n153_), .C(ori_ori_n47_), .Y(ori_ori_n154_));
  NA2        o132(.A(ori_ori_n154_), .B(ori_ori_n109_), .Y(ori_ori_n155_));
  NA2        o133(.A(x10), .B(x08), .Y(ori_ori_n156_));
  INV        o134(.A(ori_ori_n156_), .Y(ori_ori_n157_));
  NA2        o135(.A(x06), .B(x05), .Y(ori_ori_n158_));
  OAI210     o136(.A0(ori_ori_n158_), .A1(ori_ori_n35_), .B0(ori_ori_n98_), .Y(ori_ori_n159_));
  AOI210     o137(.A0(ori_ori_n157_), .A1(ori_ori_n58_), .B0(ori_ori_n159_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(ori_ori_n155_), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n99_), .B(x12), .Y(ori_ori_n162_));
  AOI210     o140(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n162_), .Y(ori_ori_n163_));
  NO2        o141(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n164_));
  NA2        o142(.A(ori_ori_n164_), .B(x02), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n163_), .B(ori_ori_n161_), .Y(ori_ori_n166_));
  NA3        o144(.A(ori_ori_n166_), .B(ori_ori_n152_), .C(ori_ori_n142_), .Y(ori_ori_n167_));
  AOI210     o145(.A0(ori_ori_n132_), .A1(ori_ori_n98_), .B0(ori_ori_n167_), .Y(ori_ori_n168_));
  NA2        o146(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n169_));
  NA2        o147(.A(ori_ori_n169_), .B(ori_ori_n119_), .Y(ori_ori_n170_));
  AOI210     o148(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n171_), .B(ori_ori_n170_), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n172_), .B(x12), .Y(ori_ori_n173_));
  INV        o151(.A(ori_ori_n76_), .Y(ori_ori_n174_));
  NO2        o152(.A(x05), .B(ori_ori_n51_), .Y(ori_ori_n175_));
  OAI210     o153(.A0(ori_ori_n175_), .A1(ori_ori_n135_), .B0(ori_ori_n57_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(ori_ori_n174_), .Y(ori_ori_n177_));
  NO2        o155(.A(ori_ori_n92_), .B(x06), .Y(ori_ori_n178_));
  AOI210     o156(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n179_));
  NO3        o157(.A(ori_ori_n179_), .B(ori_ori_n178_), .C(ori_ori_n41_), .Y(ori_ori_n180_));
  INV        o158(.A(ori_ori_n121_), .Y(ori_ori_n181_));
  OAI210     o159(.A0(ori_ori_n181_), .A1(ori_ori_n180_), .B0(x02), .Y(ori_ori_n182_));
  AOI210     o160(.A0(ori_ori_n182_), .A1(ori_ori_n177_), .B0(ori_ori_n23_), .Y(ori_ori_n183_));
  OAI210     o161(.A0(ori_ori_n173_), .A1(ori_ori_n57_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  INV        o162(.A(ori_ori_n121_), .Y(ori_ori_n185_));
  NO2        o163(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n186_));
  OAI210     o164(.A0(ori_ori_n79_), .A1(ori_ori_n36_), .B0(x04), .Y(ori_ori_n187_));
  NO2        o165(.A(ori_ori_n99_), .B(x03), .Y(ori_ori_n188_));
  AOI220     o166(.A0(ori_ori_n188_), .A1(ori_ori_n187_), .B0(ori_ori_n76_), .B1(ori_ori_n186_), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n190_));
  INV        o168(.A(ori_ori_n133_), .Y(ori_ori_n191_));
  NOi21      o169(.An(x13), .B(x04), .Y(ori_ori_n192_));
  NO3        o170(.A(ori_ori_n192_), .B(ori_ori_n76_), .C(ori_ori_n153_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n193_), .B(x05), .Y(ori_ori_n194_));
  AOI220     o172(.A0(ori_ori_n194_), .A1(ori_ori_n190_), .B0(ori_ori_n191_), .B1(ori_ori_n57_), .Y(ori_ori_n195_));
  OAI210     o173(.A0(ori_ori_n189_), .A1(ori_ori_n185_), .B0(ori_ori_n195_), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n90_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n197_), .B(x12), .Y(ori_ori_n198_));
  NA2        o176(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n199_));
  NO2        o177(.A(x06), .B(x00), .Y(ori_ori_n200_));
  NA2        o178(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n201_), .B(x03), .Y(ori_ori_n202_));
  BUFFER     o180(.A(ori_ori_n202_), .Y(ori_ori_n203_));
  NA2        o181(.A(x13), .B(ori_ori_n98_), .Y(ori_ori_n204_));
  NA3        o182(.A(ori_ori_n204_), .B(ori_ori_n159_), .C(ori_ori_n91_), .Y(ori_ori_n205_));
  OAI210     o183(.A0(ori_ori_n203_), .A1(ori_ori_n199_), .B0(ori_ori_n205_), .Y(ori_ori_n206_));
  AOI210     o184(.A0(ori_ori_n198_), .A1(ori_ori_n196_), .B0(ori_ori_n206_), .Y(ori_ori_n207_));
  AOI210     o185(.A0(ori_ori_n207_), .A1(ori_ori_n184_), .B0(x07), .Y(ori_ori_n208_));
  NA2        o186(.A(ori_ori_n72_), .B(ori_ori_n29_), .Y(ori_ori_n209_));
  NOi31      o187(.An(ori_ori_n118_), .B(ori_ori_n192_), .C(ori_ori_n153_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n210_), .B(ori_ori_n209_), .Y(ori_ori_n211_));
  NO2        o189(.A(x08), .B(x05), .Y(ori_ori_n212_));
  OAI210     o190(.A0(ori_ori_n76_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n213_));
  INV        o191(.A(ori_ori_n213_), .Y(ori_ori_n214_));
  NO2        o192(.A(x12), .B(x02), .Y(ori_ori_n215_));
  INV        o193(.A(ori_ori_n215_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n216_), .B(ori_ori_n197_), .Y(ori_ori_n217_));
  OA210      o195(.A0(ori_ori_n214_), .A1(ori_ori_n211_), .B0(ori_ori_n217_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n219_));
  NO2        o197(.A(ori_ori_n219_), .B(x01), .Y(ori_ori_n220_));
  INV        o198(.A(ori_ori_n220_), .Y(ori_ori_n221_));
  AOI210     o199(.A0(ori_ori_n221_), .A1(ori_ori_n113_), .B0(ori_ori_n29_), .Y(ori_ori_n222_));
  NA2        o200(.A(ori_ori_n99_), .B(x04), .Y(ori_ori_n223_));
  NO2        o201(.A(x02), .B(ori_ori_n104_), .Y(ori_ori_n224_));
  NO3        o202(.A(ori_ori_n89_), .B(x12), .C(x03), .Y(ori_ori_n225_));
  OAI210     o203(.A0(ori_ori_n224_), .A1(ori_ori_n222_), .B0(ori_ori_n225_), .Y(ori_ori_n226_));
  NOi21      o204(.An(ori_ori_n209_), .B(ori_ori_n178_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n227_), .B(ori_ori_n228_), .Y(ori_ori_n229_));
  NO2        o207(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n230_));
  NO3        o208(.A(ori_ori_n230_), .B(ori_ori_n179_), .C(ori_ori_n148_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n199_), .B(ori_ori_n28_), .Y(ori_ori_n232_));
  OAI210     o210(.A0(ori_ori_n231_), .A1(ori_ori_n185_), .B0(ori_ori_n232_), .Y(ori_ori_n233_));
  NA3        o211(.A(ori_ori_n233_), .B(ori_ori_n229_), .C(ori_ori_n226_), .Y(ori_ori_n234_));
  NO3        o212(.A(ori_ori_n234_), .B(ori_ori_n218_), .C(ori_ori_n208_), .Y(ori_ori_n235_));
  OAI210     o213(.A0(ori_ori_n168_), .A1(ori_ori_n61_), .B0(ori_ori_n235_), .Y(ori02));
  NO2        o214(.A(ori_ori_n99_), .B(ori_ori_n35_), .Y(ori_ori_n237_));
  NA3        o215(.A(ori_ori_n237_), .B(ori_ori_n157_), .C(ori_ori_n56_), .Y(ori_ori_n238_));
  INV        o216(.A(ori_ori_n143_), .Y(ori_ori_n239_));
  AOI220     o217(.A0(x09), .A1(ori_ori_n239_), .B0(ori_ori_n129_), .B1(ori_ori_n128_), .Y(ori_ori_n240_));
  AOI210     o218(.A0(ori_ori_n240_), .A1(ori_ori_n238_), .B0(ori_ori_n48_), .Y(ori_ori_n241_));
  NO2        o219(.A(x05), .B(x02), .Y(ori_ori_n242_));
  OAI210     o220(.A0(ori_ori_n170_), .A1(ori_ori_n153_), .B0(ori_ori_n242_), .Y(ori_ori_n243_));
  AOI220     o221(.A0(ori_ori_n212_), .A1(ori_ori_n58_), .B0(ori_ori_n56_), .B1(ori_ori_n36_), .Y(ori_ori_n244_));
  NOi21      o222(.An(ori_ori_n237_), .B(ori_ori_n244_), .Y(ori_ori_n245_));
  AOI210     o223(.A0(ori_ori_n192_), .A1(ori_ori_n79_), .B0(ori_ori_n245_), .Y(ori_ori_n246_));
  AOI210     o224(.A0(ori_ori_n246_), .A1(ori_ori_n243_), .B0(ori_ori_n121_), .Y(ori_ori_n247_));
  NAi21      o225(.An(ori_ori_n194_), .B(ori_ori_n189_), .Y(ori_ori_n248_));
  NO2        o226(.A(ori_ori_n201_), .B(ori_ori_n47_), .Y(ori_ori_n249_));
  NA2        o227(.A(ori_ori_n249_), .B(ori_ori_n248_), .Y(ori_ori_n250_));
  AN2        o228(.A(ori_ori_n188_), .B(ori_ori_n187_), .Y(ori_ori_n251_));
  NA2        o229(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n252_));
  OAI210     o230(.A0(ori_ori_n354_), .A1(ori_ori_n251_), .B0(ori_ori_n93_), .Y(ori_ori_n253_));
  INV        o231(.A(ori_ori_n128_), .Y(ori_ori_n254_));
  NO2        o232(.A(ori_ori_n254_), .B(ori_ori_n110_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n255_), .B(x13), .Y(ori_ori_n256_));
  NA3        o234(.A(ori_ori_n256_), .B(ori_ori_n253_), .C(ori_ori_n250_), .Y(ori_ori_n257_));
  NO3        o235(.A(ori_ori_n257_), .B(ori_ori_n247_), .C(ori_ori_n241_), .Y(ori_ori_n258_));
  NA2        o236(.A(ori_ori_n120_), .B(x03), .Y(ori_ori_n259_));
  OAI210     o237(.A0(ori_ori_n35_), .A1(ori_ori_n230_), .B0(ori_ori_n259_), .Y(ori_ori_n260_));
  NA2        o238(.A(ori_ori_n260_), .B(ori_ori_n100_), .Y(ori_ori_n261_));
  OAI220     o239(.A0(ori_ori_n223_), .A1(x09), .B0(ori_ori_n111_), .B1(ori_ori_n28_), .Y(ori_ori_n262_));
  NA2        o240(.A(ori_ori_n262_), .B(ori_ori_n101_), .Y(ori_ori_n263_));
  NA2        o241(.A(ori_ori_n223_), .B(ori_ori_n98_), .Y(ori_ori_n264_));
  NA3        o242(.A(x12), .B(ori_ori_n264_), .C(ori_ori_n110_), .Y(ori_ori_n265_));
  NA4        o243(.A(ori_ori_n265_), .B(ori_ori_n263_), .C(ori_ori_n261_), .D(ori_ori_n48_), .Y(ori_ori_n266_));
  INV        o244(.A(ori_ori_n164_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n138_), .B(ori_ori_n40_), .Y(ori_ori_n268_));
  NA2        o246(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n269_));
  OAI220     o247(.A0(ori_ori_n269_), .A1(ori_ori_n268_), .B0(ori_ori_n267_), .B1(ori_ori_n59_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n270_), .B(x02), .Y(ori_ori_n271_));
  NO3        o249(.A(ori_ori_n162_), .B(ori_ori_n136_), .C(ori_ori_n52_), .Y(ori_ori_n272_));
  OAI210     o250(.A0(ori_ori_n125_), .A1(ori_ori_n36_), .B0(ori_ori_n98_), .Y(ori_ori_n273_));
  OAI210     o251(.A0(ori_ori_n273_), .A1(ori_ori_n154_), .B0(ori_ori_n272_), .Y(ori_ori_n274_));
  NA3        o252(.A(ori_ori_n274_), .B(ori_ori_n271_), .C(x06), .Y(ori_ori_n275_));
  NA2        o253(.A(x09), .B(x03), .Y(ori_ori_n276_));
  OAI220     o254(.A0(ori_ori_n276_), .A1(ori_ori_n109_), .B0(ori_ori_n169_), .B1(ori_ori_n64_), .Y(ori_ori_n277_));
  NO2        o255(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n278_));
  NO3        o256(.A(ori_ori_n103_), .B(ori_ori_n109_), .C(ori_ori_n38_), .Y(ori_ori_n279_));
  AOI210     o257(.A0(ori_ori_n272_), .A1(ori_ori_n278_), .B0(ori_ori_n279_), .Y(ori_ori_n280_));
  AO220      o258(.A0(ori_ori_n353_), .A1(x04), .B0(ori_ori_n277_), .B1(x05), .Y(ori_ori_n281_));
  AOI210     o259(.A0(ori_ori_n275_), .A1(ori_ori_n266_), .B0(ori_ori_n281_), .Y(ori_ori_n282_));
  OAI210     o260(.A0(ori_ori_n258_), .A1(x12), .B0(ori_ori_n282_), .Y(ori03));
  OR2        o261(.A(ori_ori_n42_), .B(ori_ori_n186_), .Y(ori_ori_n284_));
  AOI210     o262(.A0(ori_ori_n129_), .A1(ori_ori_n98_), .B0(ori_ori_n284_), .Y(ori_ori_n285_));
  NA2        o263(.A(ori_ori_n162_), .B(ori_ori_n128_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n286_), .B(ori_ori_n165_), .Y(ori_ori_n287_));
  OAI210     o265(.A0(ori_ori_n287_), .A1(ori_ori_n285_), .B0(x05), .Y(ori_ori_n288_));
  NA2        o266(.A(ori_ori_n284_), .B(x05), .Y(ori_ori_n289_));
  AOI210     o267(.A0(ori_ori_n119_), .A1(ori_ori_n174_), .B0(ori_ori_n289_), .Y(ori_ori_n290_));
  AOI210     o268(.A0(ori_ori_n188_), .A1(ori_ori_n80_), .B0(ori_ori_n106_), .Y(ori_ori_n291_));
  OAI220     o269(.A0(ori_ori_n291_), .A1(ori_ori_n59_), .B0(ori_ori_n252_), .B1(ori_ori_n244_), .Y(ori_ori_n292_));
  OAI210     o270(.A0(ori_ori_n292_), .A1(ori_ori_n290_), .B0(ori_ori_n98_), .Y(ori_ori_n293_));
  AOI210     o271(.A0(ori_ori_n123_), .A1(ori_ori_n60_), .B0(ori_ori_n38_), .Y(ori_ori_n294_));
  NO2        o272(.A(ori_ori_n144_), .B(ori_ori_n114_), .Y(ori_ori_n295_));
  OAI220     o273(.A0(ori_ori_n295_), .A1(ori_ori_n37_), .B0(ori_ori_n126_), .B1(x13), .Y(ori_ori_n296_));
  OAI210     o274(.A0(ori_ori_n296_), .A1(ori_ori_n294_), .B0(x04), .Y(ori_ori_n297_));
  AOI210     o275(.A0(ori_ori_n150_), .A1(ori_ori_n98_), .B0(ori_ori_n123_), .Y(ori_ori_n298_));
  OA210      o276(.A0(ori_ori_n138_), .A1(x12), .B0(ori_ori_n114_), .Y(ori_ori_n299_));
  NO2        o277(.A(ori_ori_n299_), .B(ori_ori_n298_), .Y(ori_ori_n300_));
  NA4        o278(.A(ori_ori_n300_), .B(ori_ori_n297_), .C(ori_ori_n293_), .D(ori_ori_n288_), .Y(ori04));
  NO2        o279(.A(ori_ori_n88_), .B(ori_ori_n39_), .Y(ori_ori_n302_));
  XO2        o280(.A(ori_ori_n302_), .B(ori_ori_n204_), .Y(ori05));
  NA3        o281(.A(ori_ori_n121_), .B(ori_ori_n111_), .C(ori_ori_n31_), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n191_), .B(ori_ori_n57_), .Y(ori_ori_n305_));
  AOI210     o283(.A0(ori_ori_n305_), .A1(ori_ori_n304_), .B0(ori_ori_n24_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n306_), .B(ori_ori_n98_), .Y(ori_ori_n307_));
  NA2        o285(.A(ori_ori_n209_), .B(x03), .Y(ori_ori_n308_));
  OAI210     o286(.A0(ori_ori_n26_), .A1(ori_ori_n98_), .B0(x07), .Y(ori_ori_n309_));
  INV        o287(.A(ori_ori_n309_), .Y(ori_ori_n310_));
  AOI210     o288(.A0(ori_ori_n81_), .A1(ori_ori_n31_), .B0(ori_ori_n52_), .Y(ori_ori_n311_));
  NO3        o289(.A(ori_ori_n311_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n312_));
  NA2        o290(.A(ori_ori_n71_), .B(x02), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n313_), .B(ori_ori_n308_), .Y(ori_ori_n314_));
  OR2        o292(.A(ori_ori_n314_), .B(ori_ori_n199_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n200_), .B(ori_ori_n197_), .Y(ori_ori_n316_));
  NA2        o294(.A(ori_ori_n316_), .B(ori_ori_n315_), .Y(ori_ori_n317_));
  OAI210     o295(.A0(ori_ori_n317_), .A1(ori_ori_n312_), .B0(ori_ori_n98_), .Y(ori_ori_n318_));
  NA2        o296(.A(ori_ori_n33_), .B(ori_ori_n98_), .Y(ori_ori_n319_));
  AOI210     o297(.A0(ori_ori_n319_), .A1(ori_ori_n90_), .B0(x07), .Y(ori_ori_n320_));
  AOI220     o298(.A0(ori_ori_n320_), .A1(ori_ori_n318_), .B0(ori_ori_n310_), .B1(ori_ori_n307_), .Y(ori_ori_n321_));
  NOi21      o299(.An(ori_ori_n259_), .B(ori_ori_n114_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n322_), .B(ori_ori_n216_), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n323_), .B(x08), .Y(ori_ori_n324_));
  NO2        o302(.A(x05), .B(x03), .Y(ori_ori_n325_));
  NO2        o303(.A(x13), .B(x12), .Y(ori_ori_n326_));
  NO2        o304(.A(ori_ori_n111_), .B(ori_ori_n28_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n327_), .B(ori_ori_n220_), .Y(ori_ori_n328_));
  OR3        o306(.A(ori_ori_n328_), .B(x12), .C(x03), .Y(ori_ori_n329_));
  NA3        o307(.A(ori_ori_n267_), .B(ori_ori_n107_), .C(x12), .Y(ori_ori_n330_));
  AO210      o308(.A0(ori_ori_n267_), .A1(ori_ori_n107_), .B0(ori_ori_n204_), .Y(ori_ori_n331_));
  NA4        o309(.A(ori_ori_n331_), .B(ori_ori_n330_), .C(ori_ori_n329_), .D(x08), .Y(ori_ori_n332_));
  AOI210     o310(.A0(ori_ori_n326_), .A1(ori_ori_n325_), .B0(ori_ori_n332_), .Y(ori_ori_n333_));
  NO2        o311(.A(ori_ori_n324_), .B(ori_ori_n333_), .Y(ori_ori_n334_));
  NO2        o312(.A(ori_ori_n122_), .B(ori_ori_n43_), .Y(ori_ori_n335_));
  NA2        o313(.A(ori_ori_n335_), .B(ori_ori_n149_), .Y(ori_ori_n336_));
  NA3        o314(.A(ori_ori_n328_), .B(ori_ori_n322_), .C(ori_ori_n264_), .Y(ori_ori_n337_));
  INV        o315(.A(x14), .Y(ori_ori_n338_));
  NO3        o316(.A(ori_ori_n137_), .B(ori_ori_n74_), .C(ori_ori_n57_), .Y(ori_ori_n339_));
  NO2        o317(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n340_));
  NA3        o318(.A(ori_ori_n340_), .B(ori_ori_n337_), .C(ori_ori_n336_), .Y(ori_ori_n341_));
  NA2        o319(.A(ori_ori_n319_), .B(ori_ori_n61_), .Y(ori_ori_n342_));
  NOi21      o320(.An(ori_ori_n223_), .B(ori_ori_n126_), .Y(ori_ori_n343_));
  NO3        o321(.A(ori_ori_n108_), .B(ori_ori_n24_), .C(x06), .Y(ori_ori_n344_));
  AOI210     o322(.A0(ori_ori_n228_), .A1(ori_ori_n191_), .B0(ori_ori_n344_), .Y(ori_ori_n345_));
  OAI210     o323(.A0(ori_ori_n44_), .A1(x04), .B0(ori_ori_n345_), .Y(ori_ori_n346_));
  OAI210     o324(.A0(ori_ori_n346_), .A1(ori_ori_n343_), .B0(ori_ori_n98_), .Y(ori_ori_n347_));
  OAI210     o325(.A0(ori_ori_n342_), .A1(ori_ori_n89_), .B0(ori_ori_n347_), .Y(ori_ori_n348_));
  NO4        o326(.A(ori_ori_n348_), .B(ori_ori_n341_), .C(ori_ori_n334_), .D(ori_ori_n321_), .Y(ori06));
  INV        o327(.A(ori_ori_n91_), .Y(ori_ori_n352_));
  INV        o328(.A(ori_ori_n280_), .Y(ori_ori_n353_));
  INV        o329(.A(ori_ori_n123_), .Y(ori_ori_n354_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  NOi21      m029(.An(x01), .B(x09), .Y(mai_mai_n52_));
  INV        m030(.A(x00), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n50_), .B(mai_mai_n53_), .Y(mai_mai_n54_));
  NO2        m032(.A(mai_mai_n54_), .B(mai_mai_n52_), .Y(mai_mai_n55_));
  NA2        m033(.A(x09), .B(mai_mai_n53_), .Y(mai_mai_n56_));
  INV        m034(.A(x07), .Y(mai_mai_n57_));
  AOI210     m035(.A0(x11), .A1(mai_mai_n48_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  INV        m036(.A(mai_mai_n55_), .Y(mai_mai_n59_));
  OAI220     m037(.A0(x02), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .B1(mai_mai_n56_), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n60_), .B(mai_mai_n31_), .Y(mai_mai_n61_));
  NO2        m039(.A(mai_mai_n61_), .B(x05), .Y(mai_mai_n62_));
  NO2        m040(.A(mai_mai_n57_), .B(mai_mai_n23_), .Y(mai_mai_n63_));
  NA2        m041(.A(x09), .B(x05), .Y(mai_mai_n64_));
  NA2        m042(.A(x10), .B(x06), .Y(mai_mai_n65_));
  NA3        m043(.A(mai_mai_n65_), .B(mai_mai_n64_), .C(mai_mai_n28_), .Y(mai_mai_n66_));
  NO2        m044(.A(mai_mai_n57_), .B(mai_mai_n41_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n66_), .A1(mai_mai_n63_), .B0(x03), .Y(mai_mai_n68_));
  NOi31      m046(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n69_));
  INV        m047(.A(mai_mai_n24_), .Y(mai_mai_n70_));
  NO2        m048(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n71_));
  OAI210     m049(.A0(mai_mai_n71_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n72_));
  INV        m050(.A(mai_mai_n72_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n74_));
  NO2        m052(.A(x08), .B(x01), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n75_), .A1(mai_mai_n74_), .B0(mai_mai_n35_), .Y(mai_mai_n76_));
  NA2        m054(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n77_));
  NO3        m055(.A(mai_mai_n76_), .B(mai_mai_n73_), .C(mai_mai_n70_), .Y(mai_mai_n78_));
  AN2        m056(.A(mai_mai_n78_), .B(mai_mai_n68_), .Y(mai_mai_n79_));
  INV        m057(.A(mai_mai_n76_), .Y(mai_mai_n80_));
  NO2        m058(.A(x06), .B(x05), .Y(mai_mai_n81_));
  NA2        m059(.A(x11), .B(x00), .Y(mai_mai_n82_));
  NO2        m060(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n83_));
  NOi21      m061(.An(mai_mai_n82_), .B(mai_mai_n83_), .Y(mai_mai_n84_));
  AOI210     m062(.A0(mai_mai_n81_), .A1(mai_mai_n80_), .B0(mai_mai_n84_), .Y(mai_mai_n85_));
  NOi21      m063(.An(x01), .B(x10), .Y(mai_mai_n86_));
  NO2        m064(.A(mai_mai_n29_), .B(mai_mai_n53_), .Y(mai_mai_n87_));
  NO3        m065(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(x06), .Y(mai_mai_n88_));
  NA2        m066(.A(mai_mai_n88_), .B(mai_mai_n27_), .Y(mai_mai_n89_));
  OAI210     m067(.A0(mai_mai_n85_), .A1(x07), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NO3        m068(.A(mai_mai_n90_), .B(mai_mai_n79_), .C(mai_mai_n62_), .Y(mai01));
  INV        m069(.A(x12), .Y(mai_mai_n92_));
  INV        m070(.A(x13), .Y(mai_mai_n93_));
  NA2        m071(.A(x08), .B(x04), .Y(mai_mai_n94_));
  NA2        m072(.A(mai_mai_n86_), .B(mai_mai_n28_), .Y(mai_mai_n95_));
  NO2        m073(.A(mai_mai_n95_), .B(mai_mai_n64_), .Y(mai_mai_n96_));
  NO2        m074(.A(x10), .B(x01), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n98_));
  NO2        m076(.A(mai_mai_n98_), .B(mai_mai_n97_), .Y(mai_mai_n99_));
  NA2        m077(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n36_), .Y(mai_mai_n101_));
  AOI210     m079(.A0(mai_mai_n101_), .A1(mai_mai_n99_), .B0(mai_mai_n96_), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(mai_mai_n93_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n52_), .B(x05), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n105_));
  NA3        m083(.A(x13), .B(mai_mai_n105_), .C(x06), .Y(mai_mai_n106_));
  INV        m084(.A(mai_mai_n106_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n75_), .B(x13), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n392_), .B(x05), .Y(mai_mai_n109_));
  NA2        m087(.A(mai_mai_n35_), .B(mai_mai_n53_), .Y(mai_mai_n110_));
  AOI210     m088(.A0(mai_mai_n35_), .A1(x08), .B0(mai_mai_n104_), .Y(mai_mai_n111_));
  AOI210     m089(.A0(mai_mai_n111_), .A1(mai_mai_n108_), .B0(mai_mai_n65_), .Y(mai_mai_n112_));
  NA2        m090(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n113_));
  NA2        m091(.A(x10), .B(mai_mai_n53_), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n114_), .B(mai_mai_n113_), .Y(mai_mai_n115_));
  NA2        m093(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n117_));
  NO3        m095(.A(x00), .B(x06), .C(x03), .Y(mai_mai_n118_));
  NO4        m096(.A(mai_mai_n118_), .B(mai_mai_n112_), .C(mai_mai_n107_), .D(mai_mai_n103_), .Y(mai_mai_n119_));
  NA2        m097(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n120_));
  OAI210     m098(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n121_), .B(mai_mai_n120_), .Y(mai_mai_n122_));
  NO2        m100(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n124_));
  AOI210     m102(.A0(mai_mai_n124_), .A1(mai_mai_n49_), .B0(mai_mai_n123_), .Y(mai_mai_n125_));
  AN2        m103(.A(mai_mai_n125_), .B(mai_mai_n122_), .Y(mai_mai_n126_));
  NO2        m104(.A(x09), .B(x05), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(mai_mai_n47_), .Y(mai_mai_n128_));
  NO2        m106(.A(mai_mai_n99_), .B(mai_mai_n49_), .Y(mai_mai_n129_));
  NA2        m107(.A(x09), .B(x00), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n104_), .B(mai_mai_n130_), .Y(mai_mai_n131_));
  INV        m109(.A(mai_mai_n69_), .Y(mai_mai_n132_));
  AOI210     m110(.A0(mai_mai_n132_), .A1(mai_mai_n131_), .B0(mai_mai_n124_), .Y(mai_mai_n133_));
  NO3        m111(.A(mai_mai_n133_), .B(mai_mai_n129_), .C(mai_mai_n126_), .Y(mai_mai_n134_));
  NO2        m112(.A(x03), .B(x02), .Y(mai_mai_n135_));
  NA2        m113(.A(mai_mai_n76_), .B(mai_mai_n93_), .Y(mai_mai_n136_));
  OAI210     m114(.A0(mai_mai_n136_), .A1(mai_mai_n104_), .B0(mai_mai_n135_), .Y(mai_mai_n137_));
  OA210      m115(.A0(mai_mai_n134_), .A1(x11), .B0(mai_mai_n137_), .Y(mai_mai_n138_));
  OAI210     m116(.A0(mai_mai_n119_), .A1(mai_mai_n23_), .B0(mai_mai_n138_), .Y(mai_mai_n139_));
  NA2        m117(.A(mai_mai_n99_), .B(mai_mai_n40_), .Y(mai_mai_n140_));
  NAi21      m118(.An(x06), .B(x10), .Y(mai_mai_n141_));
  NOi21      m119(.An(x01), .B(x13), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n142_), .B(mai_mai_n141_), .Y(mai_mai_n143_));
  BUFFER     m121(.A(mai_mai_n143_), .Y(mai_mai_n144_));
  AOI210     m122(.A0(mai_mai_n144_), .A1(mai_mai_n140_), .B0(mai_mai_n41_), .Y(mai_mai_n145_));
  NO2        m123(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n93_), .B(x01), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n147_), .B(x08), .Y(mai_mai_n148_));
  NO2        m126(.A(mai_mai_n146_), .B(mai_mai_n48_), .Y(mai_mai_n149_));
  AOI210     m127(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n150_));
  OAI210     m128(.A0(mai_mai_n149_), .A1(mai_mai_n145_), .B0(mai_mai_n150_), .Y(mai_mai_n151_));
  NA2        m129(.A(x04), .B(x02), .Y(mai_mai_n152_));
  NA2        m130(.A(x10), .B(x05), .Y(mai_mai_n153_));
  NA2        m131(.A(x09), .B(x06), .Y(mai_mai_n154_));
  NO2        m132(.A(x09), .B(x01), .Y(mai_mai_n155_));
  NO3        m133(.A(mai_mai_n155_), .B(mai_mai_n97_), .C(mai_mai_n31_), .Y(mai_mai_n156_));
  INV        m134(.A(mai_mai_n156_), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n104_), .B(x08), .Y(mai_mai_n158_));
  OAI210     m136(.A0(mai_mai_n390_), .A1(x11), .B0(mai_mai_n157_), .Y(mai_mai_n159_));
  NAi21      m137(.An(mai_mai_n152_), .B(mai_mai_n159_), .Y(mai_mai_n160_));
  INV        m138(.A(mai_mai_n25_), .Y(mai_mai_n161_));
  NAi21      m139(.An(x13), .B(x00), .Y(mai_mai_n162_));
  AOI210     m140(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  AOI220     m141(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n164_));
  OAI210     m142(.A0(mai_mai_n153_), .A1(mai_mai_n35_), .B0(mai_mai_n164_), .Y(mai_mai_n165_));
  AN2        m143(.A(mai_mai_n165_), .B(mai_mai_n163_), .Y(mai_mai_n166_));
  BUFFER     m144(.A(mai_mai_n64_), .Y(mai_mai_n167_));
  NO2        m145(.A(mai_mai_n87_), .B(x06), .Y(mai_mai_n168_));
  NO2        m146(.A(mai_mai_n162_), .B(mai_mai_n36_), .Y(mai_mai_n169_));
  INV        m147(.A(mai_mai_n169_), .Y(mai_mai_n170_));
  OAI220     m148(.A0(mai_mai_n170_), .A1(mai_mai_n154_), .B0(mai_mai_n168_), .B1(mai_mai_n167_), .Y(mai_mai_n171_));
  OAI210     m149(.A0(mai_mai_n171_), .A1(mai_mai_n166_), .B0(mai_mai_n161_), .Y(mai_mai_n172_));
  NOi21      m150(.An(x09), .B(x00), .Y(mai_mai_n173_));
  NO3        m151(.A(mai_mai_n74_), .B(mai_mai_n173_), .C(mai_mai_n47_), .Y(mai_mai_n174_));
  INV        m152(.A(mai_mai_n174_), .Y(mai_mai_n175_));
  NA2        m153(.A(x06), .B(x05), .Y(mai_mai_n176_));
  NA2        m154(.A(mai_mai_n92_), .B(mai_mai_n175_), .Y(mai_mai_n177_));
  NO2        m155(.A(mai_mai_n93_), .B(x12), .Y(mai_mai_n178_));
  AOI210     m156(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n178_), .Y(mai_mai_n179_));
  INV        m157(.A(mai_mai_n86_), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n181_));
  NA2        m159(.A(mai_mai_n181_), .B(x02), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n182_), .B(mai_mai_n180_), .Y(mai_mai_n183_));
  AOI210     m161(.A0(mai_mai_n179_), .A1(mai_mai_n177_), .B0(mai_mai_n183_), .Y(mai_mai_n184_));
  NA4        m162(.A(mai_mai_n184_), .B(mai_mai_n172_), .C(mai_mai_n160_), .D(mai_mai_n151_), .Y(mai_mai_n185_));
  AOI210     m163(.A0(mai_mai_n139_), .A1(mai_mai_n92_), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  INV        m164(.A(mai_mai_n66_), .Y(mai_mai_n187_));
  NA2        m165(.A(mai_mai_n187_), .B(mai_mai_n122_), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n113_), .B(x06), .Y(mai_mai_n189_));
  INV        m167(.A(mai_mai_n189_), .Y(mai_mai_n190_));
  AOI210     m168(.A0(mai_mai_n190_), .A1(mai_mai_n188_), .B0(x12), .Y(mai_mai_n191_));
  INV        m169(.A(mai_mai_n69_), .Y(mai_mai_n192_));
  NA2        m170(.A(mai_mai_n143_), .B(mai_mai_n53_), .Y(mai_mai_n193_));
  NA2        m171(.A(mai_mai_n193_), .B(mai_mai_n192_), .Y(mai_mai_n194_));
  AOI210     m172(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n50_), .Y(mai_mai_n195_));
  NA4        m173(.A(mai_mai_n141_), .B(mai_mai_n52_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n196_));
  NA2        m174(.A(mai_mai_n196_), .B(mai_mai_n124_), .Y(mai_mai_n197_));
  NA2        m175(.A(mai_mai_n197_), .B(x02), .Y(mai_mai_n198_));
  AOI210     m176(.A0(mai_mai_n198_), .A1(mai_mai_n194_), .B0(mai_mai_n23_), .Y(mai_mai_n199_));
  OAI210     m177(.A0(mai_mai_n191_), .A1(mai_mai_n53_), .B0(mai_mai_n199_), .Y(mai_mai_n200_));
  INV        m178(.A(mai_mai_n124_), .Y(mai_mai_n201_));
  NO2        m179(.A(mai_mai_n50_), .B(x03), .Y(mai_mai_n202_));
  NA2        m180(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n203_));
  NOi21      m181(.An(x13), .B(x04), .Y(mai_mai_n204_));
  NO3        m182(.A(mai_mai_n204_), .B(mai_mai_n69_), .C(mai_mai_n173_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n205_), .B(x05), .Y(mai_mai_n206_));
  NA2        m184(.A(mai_mai_n206_), .B(mai_mai_n203_), .Y(mai_mai_n207_));
  INV        m185(.A(mai_mai_n207_), .Y(mai_mai_n208_));
  INV        m186(.A(mai_mai_n83_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n209_), .B(x12), .Y(mai_mai_n210_));
  NA2        m188(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n212_));
  OAI210     m190(.A0(mai_mai_n212_), .A1(mai_mai_n165_), .B0(mai_mai_n163_), .Y(mai_mai_n213_));
  AOI210     m191(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n214_));
  NO2        m192(.A(x06), .B(x00), .Y(mai_mai_n215_));
  NO3        m193(.A(mai_mai_n215_), .B(mai_mai_n214_), .C(mai_mai_n41_), .Y(mai_mai_n216_));
  OAI210     m194(.A0(mai_mai_n94_), .A1(mai_mai_n130_), .B0(mai_mai_n65_), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  NA2        m196(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n219_));
  NA2        m197(.A(mai_mai_n219_), .B(x03), .Y(mai_mai_n220_));
  OA210      m198(.A0(mai_mai_n220_), .A1(mai_mai_n218_), .B0(mai_mai_n213_), .Y(mai_mai_n221_));
  NA2        m199(.A(x13), .B(mai_mai_n92_), .Y(mai_mai_n222_));
  NA3        m200(.A(mai_mai_n222_), .B(x12), .C(mai_mai_n84_), .Y(mai_mai_n223_));
  OAI210     m201(.A0(mai_mai_n221_), .A1(mai_mai_n211_), .B0(mai_mai_n223_), .Y(mai_mai_n224_));
  AOI210     m202(.A0(mai_mai_n210_), .A1(mai_mai_n208_), .B0(mai_mai_n224_), .Y(mai_mai_n225_));
  AOI210     m203(.A0(mai_mai_n225_), .A1(mai_mai_n200_), .B0(x07), .Y(mai_mai_n226_));
  NA2        m204(.A(mai_mai_n64_), .B(mai_mai_n29_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n204_), .B(mai_mai_n173_), .Y(mai_mai_n228_));
  AOI210     m206(.A0(mai_mai_n228_), .A1(mai_mai_n132_), .B0(mai_mai_n227_), .Y(mai_mai_n229_));
  NO2        m207(.A(mai_mai_n93_), .B(x06), .Y(mai_mai_n230_));
  INV        m208(.A(mai_mai_n230_), .Y(mai_mai_n231_));
  NO2        m209(.A(x08), .B(x05), .Y(mai_mai_n232_));
  NO2        m210(.A(mai_mai_n232_), .B(mai_mai_n214_), .Y(mai_mai_n233_));
  NO2        m211(.A(mai_mai_n233_), .B(mai_mai_n231_), .Y(mai_mai_n234_));
  NO2        m212(.A(x12), .B(x02), .Y(mai_mai_n235_));
  INV        m213(.A(mai_mai_n235_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n236_), .B(mai_mai_n209_), .Y(mai_mai_n237_));
  OA210      m215(.A0(mai_mai_n234_), .A1(mai_mai_n229_), .B0(mai_mai_n237_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n239_));
  NO2        m217(.A(mai_mai_n239_), .B(x01), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n93_), .B(x04), .Y(mai_mai_n241_));
  NO3        m219(.A(mai_mai_n82_), .B(x12), .C(x03), .Y(mai_mai_n242_));
  OAI210     m220(.A0(mai_mai_n230_), .A1(mai_mai_n75_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  AOI210     m221(.A0(mai_mai_n180_), .A1(mai_mai_n176_), .B0(mai_mai_n94_), .Y(mai_mai_n244_));
  NO2        m222(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n244_), .B(mai_mai_n245_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n54_), .B(x05), .Y(mai_mai_n247_));
  NO3        m225(.A(mai_mai_n247_), .B(mai_mai_n195_), .C(mai_mai_n168_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n211_), .B(mai_mai_n28_), .Y(mai_mai_n249_));
  OAI210     m227(.A0(mai_mai_n248_), .A1(mai_mai_n201_), .B0(mai_mai_n249_), .Y(mai_mai_n250_));
  NA3        m228(.A(mai_mai_n250_), .B(mai_mai_n246_), .C(mai_mai_n243_), .Y(mai_mai_n251_));
  NO3        m229(.A(mai_mai_n251_), .B(mai_mai_n238_), .C(mai_mai_n226_), .Y(mai_mai_n252_));
  OAI210     m230(.A0(mai_mai_n186_), .A1(mai_mai_n57_), .B0(mai_mai_n252_), .Y(mai02));
  AOI210     m231(.A0(mai_mai_n120_), .A1(mai_mai_n76_), .B0(mai_mai_n116_), .Y(mai_mai_n254_));
  NOi21      m232(.An(mai_mai_n205_), .B(mai_mai_n155_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n255_), .B(mai_mai_n32_), .Y(mai_mai_n256_));
  OAI210     m234(.A0(mai_mai_n256_), .A1(mai_mai_n254_), .B0(mai_mai_n153_), .Y(mai_mai_n257_));
  INV        m235(.A(mai_mai_n153_), .Y(mai_mai_n258_));
  AOI210     m236(.A0(mai_mai_n105_), .A1(mai_mai_n77_), .B0(mai_mai_n195_), .Y(mai_mai_n259_));
  NO2        m237(.A(mai_mai_n259_), .B(mai_mai_n93_), .Y(mai_mai_n260_));
  AOI220     m238(.A0(mai_mai_n260_), .A1(mai_mai_n258_), .B0(mai_mai_n136_), .B1(mai_mai_n135_), .Y(mai_mai_n261_));
  AOI210     m239(.A0(mai_mai_n261_), .A1(mai_mai_n257_), .B0(mai_mai_n48_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n219_), .B(mai_mai_n47_), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n263_), .B(mai_mai_n206_), .Y(mai_mai_n264_));
  OAI210     m242(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n265_));
  OA210      m243(.A0(mai_mai_n391_), .A1(x08), .B0(mai_mai_n128_), .Y(mai_mai_n266_));
  AOI210     m244(.A0(mai_mai_n266_), .A1(mai_mai_n121_), .B0(mai_mai_n265_), .Y(mai_mai_n267_));
  NA2        m245(.A(mai_mai_n267_), .B(mai_mai_n87_), .Y(mai_mai_n268_));
  NA3        m246(.A(mai_mai_n87_), .B(mai_mai_n75_), .C(mai_mai_n202_), .Y(mai_mai_n269_));
  NA3        m247(.A(mai_mai_n86_), .B(mai_mai_n74_), .C(mai_mai_n42_), .Y(mai_mai_n270_));
  AOI210     m248(.A0(mai_mai_n270_), .A1(mai_mai_n269_), .B0(x04), .Y(mai_mai_n271_));
  INV        m249(.A(mai_mai_n135_), .Y(mai_mai_n272_));
  OAI220     m250(.A0(mai_mai_n233_), .A1(mai_mai_n95_), .B0(mai_mai_n272_), .B1(mai_mai_n115_), .Y(mai_mai_n273_));
  AOI210     m251(.A0(mai_mai_n273_), .A1(x13), .B0(mai_mai_n271_), .Y(mai_mai_n274_));
  NA3        m252(.A(mai_mai_n274_), .B(mai_mai_n268_), .C(mai_mai_n264_), .Y(mai_mai_n275_));
  NO2        m253(.A(mai_mai_n275_), .B(mai_mai_n262_), .Y(mai_mai_n276_));
  NA2        m254(.A(mai_mai_n123_), .B(x03), .Y(mai_mai_n277_));
  OAI210     m255(.A0(mai_mai_n162_), .A1(mai_mai_n247_), .B0(mai_mai_n277_), .Y(mai_mai_n278_));
  NA2        m256(.A(mai_mai_n278_), .B(mai_mai_n97_), .Y(mai_mai_n279_));
  NA2        m257(.A(mai_mai_n158_), .B(mai_mai_n98_), .Y(mai_mai_n280_));
  NA2        m258(.A(mai_mai_n241_), .B(mai_mai_n92_), .Y(mai_mai_n281_));
  NA2        m259(.A(mai_mai_n92_), .B(mai_mai_n41_), .Y(mai_mai_n282_));
  NA3        m260(.A(mai_mai_n282_), .B(mai_mai_n281_), .C(mai_mai_n115_), .Y(mai_mai_n283_));
  NA4        m261(.A(mai_mai_n283_), .B(mai_mai_n280_), .C(mai_mai_n279_), .D(mai_mai_n48_), .Y(mai_mai_n284_));
  INV        m262(.A(mai_mai_n181_), .Y(mai_mai_n285_));
  NO2        m263(.A(mai_mai_n148_), .B(mai_mai_n40_), .Y(mai_mai_n286_));
  NA2        m264(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n287_));
  OAI220     m265(.A0(mai_mai_n287_), .A1(mai_mai_n286_), .B0(mai_mai_n285_), .B1(mai_mai_n55_), .Y(mai_mai_n288_));
  NA2        m266(.A(mai_mai_n288_), .B(x02), .Y(mai_mai_n289_));
  INV        m267(.A(mai_mai_n212_), .Y(mai_mai_n290_));
  NA2        m268(.A(mai_mai_n178_), .B(x04), .Y(mai_mai_n291_));
  NO2        m269(.A(mai_mai_n291_), .B(mai_mai_n290_), .Y(mai_mai_n292_));
  NO3        m270(.A(mai_mai_n164_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n293_));
  OAI210     m271(.A0(mai_mai_n293_), .A1(mai_mai_n292_), .B0(mai_mai_n87_), .Y(mai_mai_n294_));
  NO3        m272(.A(mai_mai_n178_), .B(mai_mai_n146_), .C(mai_mai_n51_), .Y(mai_mai_n295_));
  OAI210     m273(.A0(mai_mai_n130_), .A1(mai_mai_n36_), .B0(mai_mai_n92_), .Y(mai_mai_n296_));
  OAI210     m274(.A0(mai_mai_n296_), .A1(mai_mai_n174_), .B0(mai_mai_n295_), .Y(mai_mai_n297_));
  NA4        m275(.A(mai_mai_n297_), .B(mai_mai_n294_), .C(mai_mai_n289_), .D(x06), .Y(mai_mai_n298_));
  OAI220     m276(.A0(mai_mai_n147_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n299_));
  NO3        m277(.A(mai_mai_n247_), .B(mai_mai_n113_), .C(x08), .Y(mai_mai_n300_));
  AOI210     m278(.A0(mai_mai_n299_), .A1(mai_mai_n201_), .B0(mai_mai_n300_), .Y(mai_mai_n301_));
  NO2        m279(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n302_));
  NO3        m280(.A(mai_mai_n104_), .B(mai_mai_n114_), .C(mai_mai_n38_), .Y(mai_mai_n303_));
  AOI210     m281(.A0(mai_mai_n295_), .A1(mai_mai_n302_), .B0(mai_mai_n303_), .Y(mai_mai_n304_));
  OAI210     m282(.A0(mai_mai_n301_), .A1(mai_mai_n28_), .B0(mai_mai_n304_), .Y(mai_mai_n305_));
  AN2        m283(.A(mai_mai_n305_), .B(x04), .Y(mai_mai_n306_));
  AOI210     m284(.A0(mai_mai_n298_), .A1(mai_mai_n284_), .B0(mai_mai_n306_), .Y(mai_mai_n307_));
  OAI210     m285(.A0(mai_mai_n276_), .A1(x12), .B0(mai_mai_n307_), .Y(mai03));
  OR2        m286(.A(mai_mai_n42_), .B(mai_mai_n202_), .Y(mai_mai_n309_));
  AOI210     m287(.A0(mai_mai_n136_), .A1(mai_mai_n92_), .B0(mai_mai_n309_), .Y(mai_mai_n310_));
  AO210      m288(.A0(mai_mai_n290_), .A1(mai_mai_n77_), .B0(mai_mai_n291_), .Y(mai_mai_n311_));
  NA2        m289(.A(mai_mai_n178_), .B(mai_mai_n135_), .Y(mai_mai_n312_));
  NA3        m290(.A(mai_mai_n312_), .B(mai_mai_n311_), .C(mai_mai_n182_), .Y(mai_mai_n313_));
  OAI210     m291(.A0(mai_mai_n313_), .A1(mai_mai_n310_), .B0(x05), .Y(mai_mai_n314_));
  NA2        m292(.A(mai_mai_n309_), .B(x05), .Y(mai_mai_n315_));
  AOI210     m293(.A0(mai_mai_n121_), .A1(mai_mai_n192_), .B0(mai_mai_n315_), .Y(mai_mai_n316_));
  INV        m294(.A(mai_mai_n109_), .Y(mai_mai_n317_));
  NO2        m295(.A(mai_mai_n317_), .B(mai_mai_n55_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(mai_mai_n318_), .A1(mai_mai_n316_), .B0(mai_mai_n92_), .Y(mai_mai_n319_));
  AOI210     m297(.A0(mai_mai_n128_), .A1(mai_mai_n56_), .B0(mai_mai_n38_), .Y(mai_mai_n320_));
  NO2        m298(.A(mai_mai_n155_), .B(mai_mai_n117_), .Y(mai_mai_n321_));
  OAI220     m299(.A0(mai_mai_n321_), .A1(mai_mai_n37_), .B0(mai_mai_n131_), .B1(x13), .Y(mai_mai_n322_));
  OAI210     m300(.A0(mai_mai_n322_), .A1(mai_mai_n320_), .B0(x04), .Y(mai_mai_n323_));
  NO3        m301(.A(mai_mai_n282_), .B(mai_mai_n76_), .C(mai_mai_n55_), .Y(mai_mai_n324_));
  AOI210     m302(.A0(mai_mai_n170_), .A1(mai_mai_n92_), .B0(mai_mai_n128_), .Y(mai_mai_n325_));
  OA210      m303(.A0(mai_mai_n148_), .A1(x12), .B0(mai_mai_n117_), .Y(mai_mai_n326_));
  NO3        m304(.A(mai_mai_n326_), .B(mai_mai_n325_), .C(mai_mai_n324_), .Y(mai_mai_n327_));
  NA4        m305(.A(mai_mai_n327_), .B(mai_mai_n323_), .C(mai_mai_n319_), .D(mai_mai_n314_), .Y(mai04));
  NO2        m306(.A(mai_mai_n80_), .B(mai_mai_n39_), .Y(mai_mai_n329_));
  XO2        m307(.A(mai_mai_n329_), .B(mai_mai_n222_), .Y(mai05));
  NO2        m308(.A(mai_mai_n51_), .B(mai_mai_n189_), .Y(mai_mai_n331_));
  AOI210     m309(.A0(mai_mai_n331_), .A1(mai_mai_n265_), .B0(mai_mai_n25_), .Y(mai_mai_n332_));
  NO2        m310(.A(x06), .B(mai_mai_n24_), .Y(mai_mai_n333_));
  OAI210     m311(.A0(mai_mai_n333_), .A1(mai_mai_n332_), .B0(mai_mai_n92_), .Y(mai_mai_n334_));
  NA2        m312(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n336_));
  NA2        m314(.A(mai_mai_n227_), .B(x03), .Y(mai_mai_n337_));
  OAI220     m315(.A0(mai_mai_n337_), .A1(mai_mai_n336_), .B0(mai_mai_n335_), .B1(mai_mai_n72_), .Y(mai_mai_n338_));
  OAI210     m316(.A0(mai_mai_n26_), .A1(mai_mai_n92_), .B0(x07), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n338_), .A1(x06), .B0(mai_mai_n339_), .Y(mai_mai_n340_));
  OR2        m318(.A(mai_mai_n93_), .B(mai_mai_n211_), .Y(mai_mai_n341_));
  NA2        m319(.A(mai_mai_n142_), .B(x05), .Y(mai_mai_n342_));
  NA3        m320(.A(mai_mai_n342_), .B(mai_mai_n215_), .C(mai_mai_n209_), .Y(mai_mai_n343_));
  NO2        m321(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n344_));
  OAI210     m322(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n345_));
  OR3        m323(.A(mai_mai_n345_), .B(mai_mai_n344_), .C(mai_mai_n44_), .Y(mai_mai_n346_));
  NA3        m324(.A(mai_mai_n346_), .B(mai_mai_n343_), .C(mai_mai_n341_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n347_), .B(mai_mai_n92_), .Y(mai_mai_n348_));
  NA2        m326(.A(mai_mai_n33_), .B(mai_mai_n92_), .Y(mai_mai_n349_));
  AOI210     m327(.A0(mai_mai_n349_), .A1(mai_mai_n83_), .B0(x07), .Y(mai_mai_n350_));
  AOI220     m328(.A0(mai_mai_n350_), .A1(mai_mai_n348_), .B0(mai_mai_n340_), .B1(mai_mai_n334_), .Y(mai_mai_n351_));
  NA3        m329(.A(mai_mai_n23_), .B(mai_mai_n57_), .C(mai_mai_n48_), .Y(mai_mai_n352_));
  AO210      m330(.A0(mai_mai_n352_), .A1(mai_mai_n239_), .B0(mai_mai_n236_), .Y(mai_mai_n353_));
  NO2        m331(.A(mai_mai_n67_), .B(mai_mai_n123_), .Y(mai_mai_n354_));
  OR2        m332(.A(mai_mai_n354_), .B(x03), .Y(mai_mai_n355_));
  NA2        m333(.A(mai_mai_n302_), .B(mai_mai_n57_), .Y(mai_mai_n356_));
  NO3        m334(.A(mai_mai_n302_), .B(mai_mai_n127_), .C(mai_mai_n28_), .Y(mai_mai_n357_));
  AOI220     m335(.A0(mai_mai_n357_), .A1(mai_mai_n355_), .B0(mai_mai_n353_), .B1(mai_mai_n47_), .Y(mai_mai_n358_));
  NA2        m336(.A(mai_mai_n358_), .B(mai_mai_n93_), .Y(mai_mai_n359_));
  AOI210     m337(.A0(mai_mai_n291_), .A1(mai_mai_n100_), .B0(mai_mai_n235_), .Y(mai_mai_n360_));
  NOi21      m338(.An(mai_mai_n277_), .B(mai_mai_n117_), .Y(mai_mai_n361_));
  NO2        m339(.A(mai_mai_n361_), .B(mai_mai_n236_), .Y(mai_mai_n362_));
  OAI210     m340(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n363_));
  AOI210     m341(.A0(mai_mai_n222_), .A1(mai_mai_n47_), .B0(mai_mai_n363_), .Y(mai_mai_n364_));
  NO4        m342(.A(mai_mai_n364_), .B(mai_mai_n362_), .C(mai_mai_n360_), .D(x08), .Y(mai_mai_n365_));
  NO2        m343(.A(mai_mai_n116_), .B(mai_mai_n28_), .Y(mai_mai_n366_));
  NO2        m344(.A(mai_mai_n366_), .B(mai_mai_n240_), .Y(mai_mai_n367_));
  NA3        m345(.A(mai_mai_n285_), .B(mai_mai_n110_), .C(x12), .Y(mai_mai_n368_));
  NA2        m346(.A(mai_mai_n368_), .B(x08), .Y(mai_mai_n369_));
  INV        m347(.A(mai_mai_n369_), .Y(mai_mai_n370_));
  AOI210     m348(.A0(mai_mai_n365_), .A1(mai_mai_n359_), .B0(mai_mai_n370_), .Y(mai_mai_n371_));
  OAI210     m349(.A0(mai_mai_n356_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n372_));
  OAI220     m350(.A0(mai_mai_n153_), .A1(mai_mai_n336_), .B0(mai_mai_n127_), .B1(mai_mai_n43_), .Y(mai_mai_n373_));
  OAI210     m351(.A0(mai_mai_n373_), .A1(mai_mai_n372_), .B0(mai_mai_n169_), .Y(mai_mai_n374_));
  NA3        m352(.A(mai_mai_n367_), .B(mai_mai_n361_), .C(mai_mai_n281_), .Y(mai_mai_n375_));
  INV        m353(.A(x14), .Y(mai_mai_n376_));
  NO3        m354(.A(mai_mai_n277_), .B(mai_mai_n95_), .C(x11), .Y(mai_mai_n377_));
  NO2        m355(.A(mai_mai_n147_), .B(mai_mai_n53_), .Y(mai_mai_n378_));
  NO3        m356(.A(mai_mai_n352_), .B(mai_mai_n282_), .C(mai_mai_n162_), .Y(mai_mai_n379_));
  NO4        m357(.A(mai_mai_n379_), .B(mai_mai_n378_), .C(mai_mai_n377_), .D(mai_mai_n376_), .Y(mai_mai_n380_));
  NA3        m358(.A(mai_mai_n380_), .B(mai_mai_n375_), .C(mai_mai_n374_), .Y(mai_mai_n381_));
  AOI220     m359(.A0(mai_mai_n349_), .A1(mai_mai_n57_), .B0(mai_mai_n366_), .B1(mai_mai_n146_), .Y(mai_mai_n382_));
  NOi21      m360(.An(mai_mai_n241_), .B(mai_mai_n131_), .Y(mai_mai_n383_));
  NO2        m361(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n384_));
  OAI210     m362(.A0(mai_mai_n384_), .A1(mai_mai_n383_), .B0(mai_mai_n92_), .Y(mai_mai_n385_));
  OAI210     m363(.A0(mai_mai_n382_), .A1(mai_mai_n82_), .B0(mai_mai_n385_), .Y(mai_mai_n386_));
  NO4        m364(.A(mai_mai_n386_), .B(mai_mai_n381_), .C(mai_mai_n371_), .D(mai_mai_n351_), .Y(mai06));
  INV        m365(.A(x01), .Y(mai_mai_n390_));
  INV        m366(.A(x13), .Y(mai_mai_n391_));
  INV        m367(.A(x13), .Y(mai_mai_n392_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  INV        u030(.A(men_men_n52_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  INV        u039(.A(men_men_n59_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  NO2        u042(.A(men_men_n64_), .B(men_men_n62_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n30_), .A1(x11), .B0(men_men_n66_), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n59_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  NA2        u048(.A(x09), .B(x05), .Y(men_men_n71_));
  NA2        u049(.A(x10), .B(x06), .Y(men_men_n72_));
  NA2        u050(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n73_));
  OAI210     u051(.A0(men_men_n73_), .A1(x11), .B0(x03), .Y(men_men_n74_));
  NOi31      u052(.An(x08), .B(x04), .C(x00), .Y(men_men_n75_));
  NO2        u053(.A(x10), .B(x09), .Y(men_men_n76_));
  NO2        u054(.A(men_men_n411_), .B(men_men_n24_), .Y(men_men_n77_));
  NO2        u055(.A(x09), .B(men_men_n41_), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n78_), .B(men_men_n36_), .Y(men_men_n79_));
  OAI210     u057(.A0(men_men_n78_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n80_));
  NO2        u058(.A(men_men_n48_), .B(men_men_n80_), .Y(men_men_n81_));
  NO2        u059(.A(men_men_n36_), .B(x00), .Y(men_men_n82_));
  NO2        u060(.A(x08), .B(x01), .Y(men_men_n83_));
  OAI210     u061(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n35_), .Y(men_men_n84_));
  NO3        u062(.A(men_men_n84_), .B(men_men_n81_), .C(men_men_n77_), .Y(men_men_n85_));
  AN2        u063(.A(men_men_n85_), .B(men_men_n74_), .Y(men_men_n86_));
  INV        u064(.A(men_men_n84_), .Y(men_men_n87_));
  NO2        u065(.A(x06), .B(x05), .Y(men_men_n88_));
  NA2        u066(.A(x11), .B(x00), .Y(men_men_n89_));
  NO2        u067(.A(x11), .B(men_men_n47_), .Y(men_men_n90_));
  NOi21      u068(.An(men_men_n89_), .B(men_men_n90_), .Y(men_men_n91_));
  NOi21      u069(.An(x01), .B(x10), .Y(men_men_n92_));
  NO2        u070(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n93_));
  NO3        u071(.A(men_men_n93_), .B(men_men_n92_), .C(x06), .Y(men_men_n94_));
  NA2        u072(.A(men_men_n94_), .B(men_men_n27_), .Y(men_men_n95_));
  OAI210     u073(.A0(men_men_n413_), .A1(x07), .B0(men_men_n95_), .Y(men_men_n96_));
  NO3        u074(.A(men_men_n96_), .B(men_men_n86_), .C(men_men_n69_), .Y(men01));
  INV        u075(.A(x12), .Y(men_men_n98_));
  INV        u076(.A(x13), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n88_), .B(x01), .Y(men_men_n100_));
  NA2        u078(.A(men_men_n100_), .B(men_men_n70_), .Y(men_men_n101_));
  NA2        u079(.A(x08), .B(x04), .Y(men_men_n102_));
  NO2        u080(.A(men_men_n102_), .B(men_men_n57_), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n103_), .B(men_men_n101_), .Y(men_men_n104_));
  NA2        u082(.A(men_men_n92_), .B(men_men_n28_), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n105_), .B(men_men_n71_), .Y(men_men_n106_));
  NO2        u084(.A(x10), .B(x01), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n29_), .B(x00), .Y(men_men_n108_));
  NO2        u086(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NA2        u087(.A(x04), .B(men_men_n28_), .Y(men_men_n110_));
  NO3        u088(.A(men_men_n110_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n111_), .B(men_men_n106_), .Y(men_men_n112_));
  AOI210     u090(.A0(men_men_n112_), .A1(men_men_n104_), .B0(men_men_n99_), .Y(men_men_n113_));
  NO2        u091(.A(men_men_n56_), .B(x05), .Y(men_men_n114_));
  NOi21      u092(.An(men_men_n114_), .B(men_men_n58_), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n99_), .B(men_men_n36_), .Y(men_men_n116_));
  NA3        u094(.A(men_men_n116_), .B(men_men_n415_), .C(x06), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n117_), .B(men_men_n115_), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n83_), .B(x13), .Y(men_men_n119_));
  NA2        u097(.A(x09), .B(men_men_n35_), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n120_), .B(men_men_n119_), .Y(men_men_n121_));
  NA2        u099(.A(x13), .B(men_men_n35_), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n122_), .B(x05), .Y(men_men_n123_));
  NO2        u101(.A(men_men_n123_), .B(men_men_n121_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n125_));
  AOI210     u103(.A0(men_men_n57_), .A1(men_men_n79_), .B0(men_men_n115_), .Y(men_men_n126_));
  AOI210     u104(.A0(men_men_n126_), .A1(men_men_n124_), .B0(men_men_n72_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n128_));
  NA2        u106(.A(x10), .B(men_men_n57_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n129_), .B(men_men_n128_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n51_), .B(x05), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n36_), .B(x04), .Y(men_men_n132_));
  NA3        u110(.A(men_men_n132_), .B(men_men_n131_), .C(x13), .Y(men_men_n133_));
  NO3        u111(.A(men_men_n125_), .B(men_men_n78_), .C(men_men_n36_), .Y(men_men_n134_));
  NO2        u112(.A(men_men_n60_), .B(x05), .Y(men_men_n135_));
  NOi31      u113(.An(men_men_n133_), .B(men_men_n134_), .C(men_men_n130_), .Y(men_men_n136_));
  NO3        u114(.A(men_men_n136_), .B(x06), .C(x03), .Y(men_men_n137_));
  NO4        u115(.A(men_men_n137_), .B(men_men_n127_), .C(men_men_n118_), .D(men_men_n113_), .Y(men_men_n138_));
  NA2        u116(.A(x13), .B(men_men_n36_), .Y(men_men_n139_));
  OAI210     u117(.A0(men_men_n83_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n140_));
  NA2        u118(.A(men_men_n140_), .B(men_men_n139_), .Y(men_men_n141_));
  OA210      u119(.A0(x00), .A1(men_men_n76_), .B0(x04), .Y(men_men_n142_));
  NO2        u120(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n29_), .B(x06), .Y(men_men_n144_));
  AOI210     u122(.A0(men_men_n144_), .A1(men_men_n49_), .B0(men_men_n143_), .Y(men_men_n145_));
  OA210      u123(.A0(men_men_n145_), .A1(men_men_n142_), .B0(men_men_n141_), .Y(men_men_n146_));
  NO2        u124(.A(x09), .B(x05), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n147_), .B(men_men_n47_), .Y(men_men_n148_));
  AOI210     u126(.A0(men_men_n148_), .A1(men_men_n109_), .B0(men_men_n49_), .Y(men_men_n149_));
  NA2        u127(.A(x09), .B(x00), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n114_), .B(men_men_n150_), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n75_), .B(men_men_n51_), .Y(men_men_n152_));
  AOI210     u130(.A0(men_men_n152_), .A1(men_men_n151_), .B0(men_men_n144_), .Y(men_men_n153_));
  NO3        u131(.A(men_men_n153_), .B(men_men_n149_), .C(men_men_n146_), .Y(men_men_n154_));
  NO2        u132(.A(x03), .B(x02), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n84_), .B(men_men_n99_), .Y(men_men_n156_));
  OAI210     u134(.A0(men_men_n156_), .A1(men_men_n115_), .B0(men_men_n155_), .Y(men_men_n157_));
  OA210      u135(.A0(men_men_n154_), .A1(x11), .B0(men_men_n157_), .Y(men_men_n158_));
  OAI210     u136(.A0(men_men_n138_), .A1(men_men_n23_), .B0(men_men_n158_), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n109_), .B(men_men_n40_), .Y(men_men_n160_));
  NAi21      u138(.An(x06), .B(x10), .Y(men_men_n161_));
  NOi21      u139(.An(x01), .B(x13), .Y(men_men_n162_));
  NA2        u140(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  OR2        u141(.A(men_men_n163_), .B(x08), .Y(men_men_n164_));
  AOI210     u142(.A0(men_men_n164_), .A1(men_men_n160_), .B0(men_men_n41_), .Y(men_men_n165_));
  NO2        u143(.A(men_men_n29_), .B(x03), .Y(men_men_n166_));
  NA2        u144(.A(men_men_n99_), .B(x01), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n167_), .B(x08), .Y(men_men_n168_));
  OAI210     u146(.A0(x05), .A1(men_men_n168_), .B0(men_men_n51_), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n169_), .A1(men_men_n166_), .B0(men_men_n48_), .Y(men_men_n170_));
  AOI210     u148(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n170_), .A1(men_men_n165_), .B0(men_men_n171_), .Y(men_men_n172_));
  NA2        u150(.A(x04), .B(x02), .Y(men_men_n173_));
  NA2        u151(.A(x10), .B(x05), .Y(men_men_n174_));
  NA2        u152(.A(x03), .B(x00), .Y(men_men_n175_));
  NO2        u153(.A(men_men_n114_), .B(x08), .Y(men_men_n176_));
  NA3        u154(.A(men_men_n162_), .B(men_men_n161_), .C(men_men_n51_), .Y(men_men_n177_));
  NA2        u155(.A(men_men_n92_), .B(x05), .Y(men_men_n178_));
  OAI210     u156(.A0(men_men_n178_), .A1(men_men_n116_), .B0(men_men_n177_), .Y(men_men_n179_));
  AOI210     u157(.A0(men_men_n176_), .A1(x06), .B0(men_men_n179_), .Y(men_men_n180_));
  OAI210     u158(.A0(men_men_n180_), .A1(x11), .B0(men_men_n175_), .Y(men_men_n181_));
  NAi21      u159(.An(men_men_n173_), .B(men_men_n181_), .Y(men_men_n182_));
  INV        u160(.A(men_men_n25_), .Y(men_men_n183_));
  NAi21      u161(.An(x13), .B(x00), .Y(men_men_n184_));
  AOI210     u162(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n184_), .Y(men_men_n185_));
  AOI220     u163(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n186_));
  OAI210     u164(.A0(men_men_n174_), .A1(men_men_n35_), .B0(men_men_n186_), .Y(men_men_n187_));
  NO2        u165(.A(men_men_n184_), .B(men_men_n36_), .Y(men_men_n188_));
  INV        u166(.A(men_men_n72_), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n189_), .A1(men_men_n185_), .B0(men_men_n183_), .Y(men_men_n190_));
  INV        u168(.A(x00), .Y(men_men_n191_));
  NA2        u169(.A(x06), .B(x05), .Y(men_men_n192_));
  OAI210     u170(.A0(men_men_n192_), .A1(men_men_n35_), .B0(men_men_n98_), .Y(men_men_n193_));
  AOI210     u171(.A0(x10), .A1(men_men_n58_), .B0(men_men_n193_), .Y(men_men_n194_));
  NO2        u172(.A(men_men_n99_), .B(x12), .Y(men_men_n195_));
  AOI210     u173(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n195_), .Y(men_men_n196_));
  NA2        u174(.A(men_men_n92_), .B(men_men_n51_), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n198_));
  NA2        u176(.A(men_men_n198_), .B(x02), .Y(men_men_n199_));
  NO2        u177(.A(men_men_n199_), .B(men_men_n197_), .Y(men_men_n200_));
  AOI210     u178(.A0(men_men_n196_), .A1(men_men_n416_), .B0(men_men_n200_), .Y(men_men_n201_));
  NA4        u179(.A(men_men_n201_), .B(men_men_n190_), .C(men_men_n182_), .D(men_men_n172_), .Y(men_men_n202_));
  AOI210     u180(.A0(men_men_n159_), .A1(men_men_n98_), .B0(men_men_n202_), .Y(men_men_n203_));
  NA2        u181(.A(men_men_n28_), .B(men_men_n141_), .Y(men_men_n204_));
  NA2        u182(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n205_));
  NA2        u183(.A(men_men_n205_), .B(men_men_n140_), .Y(men_men_n206_));
  AOI210     u184(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n207_));
  NO2        u185(.A(men_men_n128_), .B(x06), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n207_), .A1(men_men_n206_), .B0(men_men_n208_), .Y(men_men_n209_));
  AOI210     u187(.A0(men_men_n209_), .A1(men_men_n204_), .B0(x12), .Y(men_men_n210_));
  INV        u188(.A(men_men_n75_), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n92_), .B(x06), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n212_), .B(men_men_n41_), .Y(men_men_n213_));
  OAI210     u191(.A0(men_men_n56_), .A1(men_men_n213_), .B0(x02), .Y(men_men_n214_));
  AOI210     u192(.A0(men_men_n214_), .A1(men_men_n57_), .B0(men_men_n23_), .Y(men_men_n215_));
  OAI210     u193(.A0(men_men_n210_), .A1(men_men_n57_), .B0(men_men_n215_), .Y(men_men_n216_));
  INV        u194(.A(men_men_n144_), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n51_), .B(x03), .Y(men_men_n218_));
  OAI210     u196(.A0(men_men_n78_), .A1(men_men_n36_), .B0(men_men_n120_), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n99_), .B(x03), .Y(men_men_n220_));
  AOI220     u198(.A0(men_men_n220_), .A1(men_men_n219_), .B0(men_men_n75_), .B1(men_men_n218_), .Y(men_men_n221_));
  INV        u199(.A(men_men_n161_), .Y(men_men_n222_));
  NA2        u200(.A(men_men_n222_), .B(men_men_n57_), .Y(men_men_n223_));
  NA2        u201(.A(men_men_n221_), .B(men_men_n223_), .Y(men_men_n224_));
  INV        u202(.A(men_men_n90_), .Y(men_men_n225_));
  NO2        u203(.A(men_men_n225_), .B(x12), .Y(men_men_n226_));
  NA2        u204(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n228_));
  OAI210     u206(.A0(men_men_n228_), .A1(men_men_n187_), .B0(men_men_n185_), .Y(men_men_n229_));
  OAI210     u207(.A0(men_men_n102_), .A1(men_men_n150_), .B0(men_men_n72_), .Y(men_men_n230_));
  INV        u208(.A(men_men_n230_), .Y(men_men_n231_));
  INV        u209(.A(x03), .Y(men_men_n232_));
  OA210      u210(.A0(men_men_n232_), .A1(men_men_n231_), .B0(men_men_n229_), .Y(men_men_n233_));
  NA2        u211(.A(x13), .B(men_men_n98_), .Y(men_men_n234_));
  NA3        u212(.A(men_men_n234_), .B(men_men_n193_), .C(men_men_n91_), .Y(men_men_n235_));
  OAI210     u213(.A0(men_men_n233_), .A1(men_men_n227_), .B0(men_men_n235_), .Y(men_men_n236_));
  AOI210     u214(.A0(men_men_n226_), .A1(men_men_n224_), .B0(men_men_n236_), .Y(men_men_n237_));
  AOI210     u215(.A0(men_men_n237_), .A1(men_men_n216_), .B0(x07), .Y(men_men_n238_));
  NA2        u216(.A(men_men_n71_), .B(men_men_n29_), .Y(men_men_n239_));
  NA2        u217(.A(men_men_n139_), .B(men_men_n152_), .Y(men_men_n240_));
  NO2        u218(.A(men_men_n99_), .B(x06), .Y(men_men_n241_));
  INV        u219(.A(men_men_n241_), .Y(men_men_n242_));
  NO2        u220(.A(x08), .B(x05), .Y(men_men_n243_));
  NA2        u221(.A(x13), .B(men_men_n31_), .Y(men_men_n244_));
  NA2        u222(.A(men_men_n242_), .B(men_men_n244_), .Y(men_men_n245_));
  NO2        u223(.A(x12), .B(x02), .Y(men_men_n246_));
  INV        u224(.A(men_men_n246_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n247_), .B(men_men_n225_), .Y(men_men_n248_));
  OA210      u226(.A0(men_men_n245_), .A1(men_men_n240_), .B0(men_men_n248_), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n250_));
  NO2        u228(.A(men_men_n250_), .B(x01), .Y(men_men_n251_));
  NOi21      u229(.An(men_men_n83_), .B(men_men_n120_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n252_), .B(men_men_n251_), .Y(men_men_n253_));
  AOI210     u231(.A0(men_men_n253_), .A1(men_men_n133_), .B0(men_men_n29_), .Y(men_men_n254_));
  NA2        u232(.A(men_men_n241_), .B(men_men_n219_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n99_), .B(x04), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n256_), .B(men_men_n28_), .Y(men_men_n257_));
  OAI210     u235(.A0(men_men_n257_), .A1(men_men_n119_), .B0(men_men_n255_), .Y(men_men_n258_));
  NO3        u236(.A(men_men_n89_), .B(x12), .C(x03), .Y(men_men_n259_));
  OAI210     u237(.A0(men_men_n258_), .A1(men_men_n254_), .B0(men_men_n259_), .Y(men_men_n260_));
  AOI210     u238(.A0(men_men_n197_), .A1(men_men_n192_), .B0(men_men_n102_), .Y(men_men_n261_));
  NOi21      u239(.An(men_men_n239_), .B(men_men_n212_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n25_), .B(x00), .Y(men_men_n263_));
  OAI210     u241(.A0(men_men_n262_), .A1(men_men_n261_), .B0(men_men_n263_), .Y(men_men_n264_));
  NA2        u242(.A(men_men_n264_), .B(men_men_n260_), .Y(men_men_n265_));
  NO3        u243(.A(men_men_n265_), .B(men_men_n249_), .C(men_men_n238_), .Y(men_men_n266_));
  OAI210     u244(.A0(men_men_n203_), .A1(men_men_n61_), .B0(men_men_n266_), .Y(men02));
  AOI210     u245(.A0(men_men_n139_), .A1(men_men_n84_), .B0(men_men_n131_), .Y(men_men_n268_));
  NA2        u246(.A(x13), .B(men_men_n56_), .Y(men_men_n269_));
  NA2        u247(.A(men_men_n32_), .B(men_men_n269_), .Y(men_men_n270_));
  OAI210     u248(.A0(men_men_n270_), .A1(men_men_n268_), .B0(men_men_n174_), .Y(men_men_n271_));
  INV        u249(.A(men_men_n174_), .Y(men_men_n272_));
  OAI220     u250(.A0(x02), .A1(men_men_n99_), .B0(men_men_n84_), .B1(men_men_n51_), .Y(men_men_n273_));
  AOI220     u251(.A0(men_men_n273_), .A1(men_men_n272_), .B0(men_men_n156_), .B1(men_men_n155_), .Y(men_men_n274_));
  AOI210     u252(.A0(men_men_n274_), .A1(men_men_n271_), .B0(men_men_n48_), .Y(men_men_n275_));
  NO2        u253(.A(x05), .B(x02), .Y(men_men_n276_));
  OAI210     u254(.A0(men_men_n206_), .A1(men_men_n191_), .B0(men_men_n276_), .Y(men_men_n277_));
  AOI220     u255(.A0(men_men_n243_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n278_));
  NOi21      u256(.An(x13), .B(men_men_n278_), .Y(men_men_n279_));
  AOI210     u257(.A0(x13), .A1(men_men_n78_), .B0(men_men_n279_), .Y(men_men_n280_));
  AOI210     u258(.A0(men_men_n280_), .A1(men_men_n277_), .B0(men_men_n144_), .Y(men_men_n281_));
  INV        u259(.A(men_men_n221_), .Y(men_men_n282_));
  NO2        u260(.A(x10), .B(men_men_n47_), .Y(men_men_n283_));
  NA2        u261(.A(men_men_n283_), .B(men_men_n282_), .Y(men_men_n284_));
  AN2        u262(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n285_));
  OAI210     u263(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n286_));
  NA2        u264(.A(x13), .B(men_men_n28_), .Y(men_men_n287_));
  AOI210     u265(.A0(men_men_n287_), .A1(men_men_n140_), .B0(men_men_n286_), .Y(men_men_n288_));
  OAI210     u266(.A0(men_men_n288_), .A1(men_men_n285_), .B0(men_men_n93_), .Y(men_men_n289_));
  NA3        u267(.A(men_men_n93_), .B(men_men_n83_), .C(men_men_n218_), .Y(men_men_n290_));
  NA3        u268(.A(men_men_n92_), .B(men_men_n82_), .C(men_men_n42_), .Y(men_men_n291_));
  AOI210     u269(.A0(men_men_n291_), .A1(men_men_n290_), .B0(x04), .Y(men_men_n292_));
  INV        u270(.A(men_men_n105_), .Y(men_men_n293_));
  AOI210     u271(.A0(men_men_n293_), .A1(x13), .B0(men_men_n292_), .Y(men_men_n294_));
  NA3        u272(.A(men_men_n294_), .B(men_men_n289_), .C(men_men_n284_), .Y(men_men_n295_));
  NO3        u273(.A(men_men_n295_), .B(men_men_n281_), .C(men_men_n275_), .Y(men_men_n296_));
  NA2        u274(.A(men_men_n143_), .B(x03), .Y(men_men_n297_));
  INV        u275(.A(men_men_n184_), .Y(men_men_n298_));
  AOI220     u276(.A0(x08), .A1(men_men_n298_), .B0(men_men_n198_), .B1(x08), .Y(men_men_n299_));
  NA2        u277(.A(men_men_n299_), .B(men_men_n297_), .Y(men_men_n300_));
  NA2        u278(.A(men_men_n300_), .B(men_men_n107_), .Y(men_men_n301_));
  NA2        u279(.A(men_men_n173_), .B(men_men_n167_), .Y(men_men_n302_));
  AN2        u280(.A(men_men_n302_), .B(men_men_n176_), .Y(men_men_n303_));
  INV        u281(.A(men_men_n56_), .Y(men_men_n304_));
  OAI220     u282(.A0(men_men_n256_), .A1(men_men_n304_), .B0(men_men_n131_), .B1(men_men_n28_), .Y(men_men_n305_));
  OAI210     u283(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n108_), .Y(men_men_n306_));
  NA2        u284(.A(men_men_n256_), .B(men_men_n98_), .Y(men_men_n307_));
  NA2        u285(.A(men_men_n98_), .B(men_men_n41_), .Y(men_men_n308_));
  NA3        u286(.A(men_men_n308_), .B(men_men_n307_), .C(men_men_n130_), .Y(men_men_n309_));
  NA4        u287(.A(men_men_n309_), .B(men_men_n306_), .C(men_men_n301_), .D(men_men_n48_), .Y(men_men_n310_));
  INV        u288(.A(men_men_n198_), .Y(men_men_n311_));
  NO2        u289(.A(men_men_n414_), .B(men_men_n31_), .Y(men_men_n312_));
  NA2        u290(.A(men_men_n312_), .B(x02), .Y(men_men_n313_));
  INV        u291(.A(men_men_n228_), .Y(men_men_n314_));
  NA2        u292(.A(men_men_n195_), .B(x04), .Y(men_men_n315_));
  NO2        u293(.A(men_men_n315_), .B(men_men_n314_), .Y(men_men_n316_));
  NO3        u294(.A(men_men_n186_), .B(x13), .C(men_men_n31_), .Y(men_men_n317_));
  OAI210     u295(.A0(men_men_n317_), .A1(men_men_n316_), .B0(men_men_n93_), .Y(men_men_n318_));
  NO3        u296(.A(men_men_n195_), .B(men_men_n166_), .C(men_men_n52_), .Y(men_men_n319_));
  OAI210     u297(.A0(x12), .A1(x01), .B0(men_men_n319_), .Y(men_men_n320_));
  NA4        u298(.A(men_men_n320_), .B(men_men_n318_), .C(men_men_n313_), .D(x06), .Y(men_men_n321_));
  NA2        u299(.A(x09), .B(x03), .Y(men_men_n322_));
  OAI220     u300(.A0(men_men_n322_), .A1(men_men_n129_), .B0(men_men_n205_), .B1(men_men_n63_), .Y(men_men_n323_));
  NO2        u301(.A(men_men_n128_), .B(x08), .Y(men_men_n324_));
  AOI210     u302(.A0(x01), .A1(men_men_n217_), .B0(men_men_n324_), .Y(men_men_n325_));
  NO2        u303(.A(men_men_n325_), .B(men_men_n28_), .Y(men_men_n326_));
  AO220      u304(.A0(men_men_n326_), .A1(x04), .B0(men_men_n323_), .B1(x05), .Y(men_men_n327_));
  AOI210     u305(.A0(men_men_n321_), .A1(men_men_n310_), .B0(men_men_n327_), .Y(men_men_n328_));
  OAI210     u306(.A0(men_men_n296_), .A1(x12), .B0(men_men_n328_), .Y(men03));
  OR2        u307(.A(men_men_n42_), .B(men_men_n218_), .Y(men_men_n330_));
  AOI210     u308(.A0(men_men_n156_), .A1(men_men_n98_), .B0(men_men_n330_), .Y(men_men_n331_));
  OAI210     u309(.A0(men_men_n417_), .A1(men_men_n331_), .B0(x05), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n330_), .B(x05), .Y(men_men_n333_));
  AOI210     u311(.A0(men_men_n140_), .A1(men_men_n211_), .B0(men_men_n333_), .Y(men_men_n334_));
  AOI210     u312(.A0(men_men_n220_), .A1(men_men_n79_), .B0(men_men_n123_), .Y(men_men_n335_));
  OAI220     u313(.A0(men_men_n335_), .A1(men_men_n59_), .B0(men_men_n287_), .B1(men_men_n278_), .Y(men_men_n336_));
  OAI210     u314(.A0(men_men_n336_), .A1(men_men_n334_), .B0(men_men_n98_), .Y(men_men_n337_));
  NO2        u315(.A(men_men_n151_), .B(x13), .Y(men_men_n338_));
  NA2        u316(.A(men_men_n338_), .B(x04), .Y(men_men_n339_));
  NO3        u317(.A(men_men_n308_), .B(men_men_n84_), .C(men_men_n59_), .Y(men_men_n340_));
  NO2        u318(.A(men_men_n98_), .B(men_men_n148_), .Y(men_men_n341_));
  OA210      u319(.A0(men_men_n168_), .A1(x12), .B0(men_men_n135_), .Y(men_men_n342_));
  NO3        u320(.A(men_men_n342_), .B(men_men_n341_), .C(men_men_n340_), .Y(men_men_n343_));
  NA4        u321(.A(men_men_n343_), .B(men_men_n339_), .C(men_men_n337_), .D(men_men_n332_), .Y(men04));
  NO2        u322(.A(men_men_n87_), .B(men_men_n39_), .Y(men_men_n345_));
  XO2        u323(.A(men_men_n345_), .B(men_men_n234_), .Y(men05));
  AOI210     u324(.A0(men_men_n71_), .A1(men_men_n52_), .B0(men_men_n208_), .Y(men_men_n347_));
  AOI210     u325(.A0(men_men_n347_), .A1(men_men_n286_), .B0(men_men_n25_), .Y(men_men_n348_));
  NAi31      u326(.An(men_men_n76_), .B(men_men_n131_), .C(men_men_n31_), .Y(men_men_n349_));
  AOI210     u327(.A0(men_men_n412_), .A1(men_men_n349_), .B0(men_men_n24_), .Y(men_men_n350_));
  OAI210     u328(.A0(men_men_n350_), .A1(men_men_n348_), .B0(men_men_n98_), .Y(men_men_n351_));
  NA2        u329(.A(x11), .B(men_men_n31_), .Y(men_men_n352_));
  NA2        u330(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n353_));
  NA2        u331(.A(men_men_n239_), .B(x03), .Y(men_men_n354_));
  OAI220     u332(.A0(men_men_n354_), .A1(men_men_n353_), .B0(men_men_n352_), .B1(men_men_n80_), .Y(men_men_n355_));
  OAI210     u333(.A0(men_men_n26_), .A1(men_men_n98_), .B0(x07), .Y(men_men_n356_));
  AOI210     u334(.A0(men_men_n355_), .A1(x06), .B0(men_men_n356_), .Y(men_men_n357_));
  AOI220     u335(.A0(men_men_n80_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n358_));
  NO3        u336(.A(men_men_n358_), .B(men_men_n23_), .C(x00), .Y(men_men_n359_));
  NA2        u337(.A(men_men_n70_), .B(x02), .Y(men_men_n360_));
  AOI210     u338(.A0(men_men_n360_), .A1(men_men_n354_), .B0(men_men_n241_), .Y(men_men_n361_));
  OR2        u339(.A(men_men_n361_), .B(men_men_n227_), .Y(men_men_n362_));
  NO2        u340(.A(men_men_n23_), .B(x10), .Y(men_men_n363_));
  OAI210     u341(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n364_));
  OR3        u342(.A(men_men_n364_), .B(men_men_n363_), .C(men_men_n44_), .Y(men_men_n365_));
  NA2        u343(.A(men_men_n365_), .B(men_men_n362_), .Y(men_men_n366_));
  OAI210     u344(.A0(men_men_n366_), .A1(men_men_n359_), .B0(men_men_n98_), .Y(men_men_n367_));
  AOI210     u345(.A0(x12), .A1(men_men_n90_), .B0(x07), .Y(men_men_n368_));
  AOI220     u346(.A0(men_men_n368_), .A1(men_men_n367_), .B0(men_men_n357_), .B1(men_men_n351_), .Y(men_men_n369_));
  BUFFER     u347(.A(men_men_n247_), .Y(men_men_n370_));
  AOI210     u348(.A0(men_men_n363_), .A1(x07), .B0(men_men_n143_), .Y(men_men_n371_));
  OR2        u349(.A(men_men_n371_), .B(x03), .Y(men_men_n372_));
  NO2        u350(.A(x07), .B(x11), .Y(men_men_n373_));
  NO3        u351(.A(men_men_n373_), .B(men_men_n147_), .C(men_men_n28_), .Y(men_men_n374_));
  AOI220     u352(.A0(men_men_n374_), .A1(men_men_n372_), .B0(men_men_n370_), .B1(men_men_n47_), .Y(men_men_n375_));
  NA2        u353(.A(men_men_n375_), .B(men_men_n99_), .Y(men_men_n376_));
  AOI210     u354(.A0(men_men_n315_), .A1(men_men_n110_), .B0(men_men_n246_), .Y(men_men_n377_));
  NOi21      u355(.An(men_men_n297_), .B(men_men_n135_), .Y(men_men_n378_));
  OAI210     u356(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n234_), .A1(men_men_n47_), .B0(men_men_n379_), .Y(men_men_n380_));
  NO3        u358(.A(men_men_n380_), .B(men_men_n377_), .C(x08), .Y(men_men_n381_));
  NO2        u359(.A(men_men_n352_), .B(men_men_n66_), .Y(men_men_n382_));
  NO2        u360(.A(men_men_n131_), .B(men_men_n28_), .Y(men_men_n383_));
  NO2        u361(.A(men_men_n383_), .B(men_men_n251_), .Y(men_men_n384_));
  OR3        u362(.A(men_men_n384_), .B(x12), .C(x03), .Y(men_men_n385_));
  NA3        u363(.A(men_men_n311_), .B(men_men_n125_), .C(x12), .Y(men_men_n386_));
  AO210      u364(.A0(men_men_n311_), .A1(men_men_n125_), .B0(men_men_n234_), .Y(men_men_n387_));
  NA4        u365(.A(men_men_n387_), .B(men_men_n386_), .C(men_men_n385_), .D(x08), .Y(men_men_n388_));
  NO2        u366(.A(men_men_n382_), .B(men_men_n388_), .Y(men_men_n389_));
  AOI210     u367(.A0(men_men_n381_), .A1(men_men_n376_), .B0(men_men_n389_), .Y(men_men_n390_));
  OAI210     u368(.A0(x07), .A1(men_men_n23_), .B0(x03), .Y(men_men_n391_));
  INV        u369(.A(x07), .Y(men_men_n392_));
  NO2        u370(.A(men_men_n392_), .B(men_men_n353_), .Y(men_men_n393_));
  OAI210     u371(.A0(men_men_n393_), .A1(men_men_n391_), .B0(men_men_n188_), .Y(men_men_n394_));
  NA3        u372(.A(men_men_n384_), .B(men_men_n378_), .C(men_men_n307_), .Y(men_men_n395_));
  INV        u373(.A(x14), .Y(men_men_n396_));
  NO3        u374(.A(men_men_n297_), .B(men_men_n105_), .C(x11), .Y(men_men_n397_));
  NO3        u375(.A(x07), .B(men_men_n308_), .C(men_men_n184_), .Y(men_men_n398_));
  NO3        u376(.A(men_men_n398_), .B(men_men_n397_), .C(men_men_n396_), .Y(men_men_n399_));
  NA3        u377(.A(men_men_n399_), .B(men_men_n395_), .C(men_men_n394_), .Y(men_men_n400_));
  AOI220     u378(.A0(x12), .A1(men_men_n61_), .B0(men_men_n383_), .B1(men_men_n166_), .Y(men_men_n401_));
  INV        u379(.A(men_men_n151_), .Y(men_men_n402_));
  NO3        u380(.A(men_men_n128_), .B(men_men_n24_), .C(x06), .Y(men_men_n403_));
  AOI210     u381(.A0(men_men_n263_), .A1(men_men_n222_), .B0(men_men_n403_), .Y(men_men_n404_));
  OAI210     u382(.A0(men_men_n44_), .A1(x04), .B0(men_men_n404_), .Y(men_men_n405_));
  OAI210     u383(.A0(men_men_n405_), .A1(men_men_n402_), .B0(men_men_n98_), .Y(men_men_n406_));
  OAI210     u384(.A0(men_men_n401_), .A1(men_men_n89_), .B0(men_men_n406_), .Y(men_men_n407_));
  NO4        u385(.A(men_men_n407_), .B(men_men_n400_), .C(men_men_n390_), .D(men_men_n369_), .Y(men06));
  INV        u386(.A(x07), .Y(men_men_n411_));
  INV        u387(.A(men_men_n88_), .Y(men_men_n412_));
  INV        u388(.A(men_men_n91_), .Y(men_men_n413_));
  INV        u389(.A(x05), .Y(men_men_n414_));
  INV        u390(.A(x02), .Y(men_men_n415_));
  INV        u391(.A(men_men_n194_), .Y(men_men_n416_));
  INV        u392(.A(men_men_n315_), .Y(men_men_n417_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule