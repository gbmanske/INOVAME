// Benchmark "top" written by ABC on Thu Jun 20 14:00:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n97_, new_new_n98_, new_new_n100_,
    new_new_n101_, new_new_n102_, new_new_n103_, new_new_n104_,
    new_new_n105_, new_new_n106_, new_new_n107_, new_new_n108_,
    new_new_n109_, new_new_n110_, new_new_n111_, new_new_n112_,
    new_new_n113_, new_new_n114_, new_new_n115_, new_new_n116_,
    new_new_n117_, new_new_n118_, new_new_n119_, new_new_n120_,
    new_new_n121_, new_new_n122_, new_new_n123_, new_new_n124_,
    new_new_n125_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n395_, new_new_n396_, new_new_n397_,
    new_new_n398_, new_new_n399_, new_new_n400_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n406_, new_new_n407_, new_new_n408_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n489_, new_new_n490_,
    new_new_n491_, new_new_n492_, new_new_n493_, new_new_n494_,
    new_new_n495_, new_new_n496_, new_new_n497_, new_new_n498_,
    new_new_n499_, new_new_n500_, new_new_n501_, new_new_n502_,
    new_new_n503_, new_new_n504_, new_new_n505_, new_new_n506_,
    new_new_n507_, new_new_n508_, new_new_n509_, new_new_n510_,
    new_new_n511_, new_new_n512_, new_new_n513_, new_new_n514_,
    new_new_n515_, new_new_n516_, new_new_n517_, new_new_n518_,
    new_new_n519_, new_new_n520_, new_new_n521_, new_new_n522_,
    new_new_n523_, new_new_n524_, new_new_n525_, new_new_n526_,
    new_new_n527_, new_new_n528_, new_new_n529_, new_new_n530_,
    new_new_n531_, new_new_n532_, new_new_n533_, new_new_n534_,
    new_new_n536_, new_new_n537_, new_new_n538_, new_new_n539_,
    new_new_n540_, new_new_n541_, new_new_n542_, new_new_n543_,
    new_new_n544_, new_new_n545_, new_new_n546_, new_new_n547_,
    new_new_n548_, new_new_n549_, new_new_n550_, new_new_n551_,
    new_new_n552_, new_new_n553_, new_new_n554_, new_new_n555_,
    new_new_n556_, new_new_n557_, new_new_n558_, new_new_n559_,
    new_new_n560_, new_new_n561_, new_new_n562_, new_new_n563_,
    new_new_n564_, new_new_n565_, new_new_n566_, new_new_n567_,
    new_new_n568_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n653_, new_new_n654_, new_new_n655_, new_new_n656_,
    new_new_n657_, new_new_n658_, new_new_n659_, new_new_n660_,
    new_new_n661_, new_new_n662_, new_new_n663_, new_new_n664_,
    new_new_n665_, new_new_n666_, new_new_n667_, new_new_n668_,
    new_new_n669_, new_new_n670_, new_new_n671_, new_new_n672_,
    new_new_n673_, new_new_n674_, new_new_n675_, new_new_n676_,
    new_new_n677_, new_new_n678_, new_new_n679_, new_new_n680_,
    new_new_n681_, new_new_n682_, new_new_n683_, new_new_n684_,
    new_new_n685_, new_new_n686_, new_new_n687_, new_new_n688_,
    new_new_n689_, new_new_n690_, new_new_n691_, new_new_n692_,
    new_new_n693_, new_new_n694_, new_new_n695_, new_new_n696_,
    new_new_n697_, new_new_n698_, new_new_n699_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n703_, new_new_n704_,
    new_new_n705_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NAi31      g018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(zz01));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  NA2        g027(.A(i_0_), .B(i_2_), .Y(new_new_n50_));
  NA2        g028(.A(i_7_), .B(i_9_), .Y(new_new_n51_));
  NO2        g029(.A(new_new_n51_), .B(new_new_n50_), .Y(new_new_n52_));
  NA3        g030(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n53_));
  NO2        g031(.A(i_1_), .B(i_6_), .Y(new_new_n54_));
  NA2        g032(.A(i_8_), .B(i_7_), .Y(new_new_n55_));
  INV        g033(.A(i_1_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n49_), .B(i_2_), .Y(new_new_n57_));
  AOI210     g035(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n58_));
  NA2        g036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NO2        g037(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n60_));
  INV        g038(.A(i_0_), .Y(new_new_n61_));
  NAi21      g039(.An(i_5_), .B(i_10_), .Y(new_new_n62_));
  NA2        g040(.A(i_5_), .B(i_9_), .Y(new_new_n63_));
  AOI210     g041(.A0(new_new_n63_), .A1(new_new_n62_), .B0(new_new_n61_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(new_new_n60_), .Y(new_new_n65_));
  NA2        g043(.A(i_12_), .B(i_5_), .Y(new_new_n66_));
  NA2        g044(.A(i_2_), .B(i_8_), .Y(new_new_n67_));
  NO2        g045(.A(i_3_), .B(i_9_), .Y(new_new_n68_));
  NO2        g046(.A(i_3_), .B(i_7_), .Y(new_new_n69_));
  INV        g047(.A(i_6_), .Y(new_new_n70_));
  INV        g048(.A(i_11_), .Y(new_new_n71_));
  NO2        g049(.A(i_2_), .B(i_7_), .Y(new_new_n72_));
  NAi21      g050(.An(i_6_), .B(i_10_), .Y(new_new_n73_));
  NA2        g051(.A(i_6_), .B(i_9_), .Y(new_new_n74_));
  NA2        g052(.A(i_2_), .B(i_6_), .Y(new_new_n75_));
  AN3        g053(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n76_));
  NAi21      g054(.An(i_6_), .B(i_11_), .Y(new_new_n77_));
  NA2        g055(.A(new_new_n76_), .B(new_new_n32_), .Y(new_new_n78_));
  INV        g056(.A(i_7_), .Y(new_new_n79_));
  NO2        g057(.A(i_0_), .B(i_5_), .Y(new_new_n80_));
  NA2        g058(.A(i_12_), .B(i_3_), .Y(new_new_n81_));
  NAi21      g059(.An(i_7_), .B(i_11_), .Y(new_new_n82_));
  AN2        g060(.A(i_2_), .B(i_10_), .Y(new_new_n83_));
  NO2        g061(.A(new_new_n83_), .B(i_7_), .Y(new_new_n84_));
  NA2        g062(.A(i_12_), .B(i_7_), .Y(new_new_n85_));
  NO2        g063(.A(new_new_n56_), .B(new_new_n26_), .Y(new_new_n86_));
  NA2        g064(.A(i_11_), .B(i_12_), .Y(new_new_n87_));
  NA2        g065(.A(new_new_n87_), .B(new_new_n78_), .Y(new_new_n88_));
  NA2        g066(.A(new_new_n79_), .B(new_new_n37_), .Y(new_new_n89_));
  NA2        g067(.A(i_7_), .B(new_new_n25_), .Y(new_new_n90_));
  NA2        g068(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n91_));
  NO2        g069(.A(new_new_n91_), .B(new_new_n45_), .Y(new_new_n92_));
  NA2        g070(.A(new_new_n74_), .B(new_new_n73_), .Y(new_new_n93_));
  NO2        g071(.A(i_1_), .B(new_new_n70_), .Y(new_new_n94_));
  NO2        g072(.A(i_6_), .B(i_5_), .Y(new_new_n95_));
  NA2        g073(.A(new_new_n750_), .B(new_new_n745_), .Y(zz02));
  NO2        g074(.A(new_new_n56_), .B(new_new_n37_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n752_), .B(new_new_n97_), .Y(new_new_n98_));
  NA4        g076(.A(new_new_n98_), .B(new_new_n65_), .C(new_new_n57_), .D(new_new_n30_), .Y(zz00));
  AN2        g077(.A(i_8_), .B(i_7_), .Y(new_new_n100_));
  NA2        g078(.A(new_new_n100_), .B(i_6_), .Y(new_new_n101_));
  NO2        g079(.A(i_12_), .B(i_13_), .Y(new_new_n102_));
  NAi21      g080(.An(i_5_), .B(i_11_), .Y(new_new_n103_));
  NOi21      g081(.An(new_new_n102_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g082(.A(i_0_), .B(i_1_), .Y(new_new_n105_));
  NA2        g083(.A(i_2_), .B(i_3_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(i_4_), .Y(new_new_n107_));
  NA3        g085(.A(new_new_n107_), .B(new_new_n105_), .C(new_new_n104_), .Y(new_new_n108_));
  AN2        g086(.A(new_new_n102_), .B(new_new_n68_), .Y(new_new_n109_));
  NA2        g087(.A(i_1_), .B(i_5_), .Y(new_new_n110_));
  NA2        g088(.A(i_2_), .B(new_new_n36_), .Y(new_new_n111_));
  NO3        g089(.A(new_new_n111_), .B(new_new_n110_), .C(i_13_), .Y(new_new_n112_));
  OR2        g090(.A(i_0_), .B(i_1_), .Y(new_new_n113_));
  NO3        g091(.A(new_new_n113_), .B(new_new_n66_), .C(i_13_), .Y(new_new_n114_));
  NAi32      g092(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n115_));
  NAi21      g093(.An(new_new_n115_), .B(new_new_n114_), .Y(new_new_n116_));
  NOi21      g094(.An(i_4_), .B(i_10_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(new_new_n39_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n118_), .B(new_new_n116_), .Y(new_new_n119_));
  NO2        g097(.A(new_new_n119_), .B(new_new_n112_), .Y(new_new_n120_));
  AOI210     g098(.A0(new_new_n120_), .A1(new_new_n108_), .B0(new_new_n101_), .Y(new_new_n121_));
  NOi21      g099(.An(i_4_), .B(i_9_), .Y(new_new_n122_));
  NOi21      g100(.An(i_11_), .B(i_13_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n122_), .Y(new_new_n124_));
  BUFFER     g102(.A(new_new_n124_), .Y(new_new_n125_));
  NO2        g103(.A(i_4_), .B(i_5_), .Y(new_new_n126_));
  NAi21      g104(.An(i_12_), .B(i_11_), .Y(new_new_n127_));
  NO2        g105(.A(new_new_n127_), .B(i_13_), .Y(new_new_n128_));
  NA3        g106(.A(new_new_n128_), .B(new_new_n126_), .C(new_new_n68_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n129_), .B(new_new_n125_), .Y(new_new_n130_));
  NO2        g108(.A(new_new_n61_), .B(new_new_n56_), .Y(new_new_n131_));
  NAi31      g109(.An(new_new_n741_), .B(new_new_n109_), .C(i_11_), .Y(new_new_n132_));
  NA2        g110(.A(i_3_), .B(i_5_), .Y(new_new_n133_));
  AOI210     g111(.A0(new_new_n124_), .A1(new_new_n132_), .B0(new_new_n56_), .Y(new_new_n134_));
  NO2        g112(.A(new_new_n61_), .B(i_5_), .Y(new_new_n135_));
  NO2        g113(.A(i_13_), .B(i_10_), .Y(new_new_n136_));
  NA3        g114(.A(new_new_n136_), .B(new_new_n135_), .C(new_new_n43_), .Y(new_new_n137_));
  NO2        g115(.A(i_2_), .B(i_1_), .Y(new_new_n138_));
  NAi21      g116(.An(i_4_), .B(i_12_), .Y(new_new_n139_));
  NO4        g117(.A(new_new_n139_), .B(i_2_), .C(new_new_n137_), .D(new_new_n25_), .Y(new_new_n140_));
  NO3        g118(.A(new_new_n140_), .B(new_new_n134_), .C(new_new_n130_), .Y(new_new_n141_));
  INV        g119(.A(i_8_), .Y(new_new_n142_));
  NO3        g120(.A(i_3_), .B(new_new_n70_), .C(new_new_n47_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(i_7_), .Y(new_new_n144_));
  NA2        g122(.A(new_new_n39_), .B(new_new_n43_), .Y(new_new_n145_));
  NO3        g123(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n146_));
  OAI210     g124(.A0(new_new_n76_), .A1(i_12_), .B0(new_new_n146_), .Y(new_new_n147_));
  AOI210     g125(.A0(new_new_n147_), .A1(new_new_n145_), .B0(new_new_n144_), .Y(new_new_n148_));
  NO3        g126(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n149_));
  NA2        g127(.A(new_new_n149_), .B(new_new_n39_), .Y(new_new_n150_));
  NO2        g128(.A(i_13_), .B(i_9_), .Y(new_new_n151_));
  NAi21      g129(.An(i_12_), .B(i_3_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n43_), .B(i_5_), .Y(new_new_n153_));
  NO2        g131(.A(new_new_n54_), .B(new_new_n150_), .Y(new_new_n154_));
  AOI210     g132(.A0(new_new_n154_), .A1(i_7_), .B0(new_new_n148_), .Y(new_new_n155_));
  OAI210     g133(.A0(new_new_n155_), .A1(i_4_), .B0(new_new_n141_), .Y(new_new_n156_));
  NA3        g134(.A(i_13_), .B(new_new_n142_), .C(i_10_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n157_), .B(i_12_), .Y(new_new_n158_));
  NA2        g136(.A(i_0_), .B(i_5_), .Y(new_new_n159_));
  NAi31      g137(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n45_), .B(new_new_n56_), .Y(new_new_n161_));
  INV        g139(.A(i_13_), .Y(new_new_n162_));
  NO2        g140(.A(i_12_), .B(new_new_n162_), .Y(new_new_n163_));
  NA2        g141(.A(new_new_n163_), .B(new_new_n143_), .Y(new_new_n164_));
  INV        g142(.A(new_new_n164_), .Y(new_new_n165_));
  AOI210     g143(.A0(new_new_n165_), .A1(new_new_n100_), .B0(new_new_n158_), .Y(new_new_n166_));
  NO2        g144(.A(i_12_), .B(new_new_n37_), .Y(new_new_n167_));
  NO2        g145(.A(new_new_n133_), .B(i_4_), .Y(new_new_n168_));
  NA2        g146(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n169_));
  OR2        g147(.A(i_8_), .B(i_7_), .Y(new_new_n170_));
  INV        g148(.A(i_12_), .Y(new_new_n171_));
  NO3        g149(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n172_));
  NA2        g150(.A(i_2_), .B(i_1_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n170_), .B(new_new_n169_), .Y(new_new_n174_));
  NO3        g152(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n175_));
  NAi21      g153(.An(i_4_), .B(i_3_), .Y(new_new_n176_));
  NO2        g154(.A(i_0_), .B(i_6_), .Y(new_new_n177_));
  NOi41      g155(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n178_));
  NA2        g156(.A(new_new_n178_), .B(new_new_n177_), .Y(new_new_n179_));
  AOI220     g157(.A0(new_new_n178_), .A1(new_new_n39_), .B0(new_new_n174_), .B1(new_new_n151_), .Y(new_new_n180_));
  NO2        g158(.A(i_11_), .B(new_new_n162_), .Y(new_new_n181_));
  NOi21      g159(.An(i_1_), .B(i_6_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n171_), .B(i_9_), .Y(new_new_n183_));
  NO2        g161(.A(i_12_), .B(i_3_), .Y(new_new_n184_));
  NA2        g162(.A(i_3_), .B(i_9_), .Y(new_new_n185_));
  NAi21      g163(.An(i_7_), .B(i_10_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n186_), .B(new_new_n185_), .Y(new_new_n187_));
  NA3        g165(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n188_));
  INV        g166(.A(new_new_n101_), .Y(new_new_n189_));
  NA2        g167(.A(new_new_n171_), .B(i_13_), .Y(new_new_n190_));
  NO2        g168(.A(new_new_n190_), .B(new_new_n63_), .Y(new_new_n191_));
  AOI220     g169(.A0(new_new_n191_), .A1(new_new_n189_), .B0(i_9_), .B1(new_new_n181_), .Y(new_new_n192_));
  NO2        g170(.A(new_new_n170_), .B(new_new_n37_), .Y(new_new_n193_));
  NA2        g171(.A(i_12_), .B(i_6_), .Y(new_new_n194_));
  OR2        g172(.A(i_13_), .B(i_9_), .Y(new_new_n195_));
  NO3        g173(.A(new_new_n195_), .B(new_new_n194_), .C(new_new_n47_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n176_), .B(i_2_), .Y(new_new_n197_));
  NA3        g175(.A(new_new_n197_), .B(new_new_n196_), .C(new_new_n43_), .Y(new_new_n198_));
  NA2        g176(.A(new_new_n181_), .B(i_9_), .Y(new_new_n199_));
  OAI210     g177(.A0(new_new_n56_), .A1(new_new_n199_), .B0(new_new_n198_), .Y(new_new_n200_));
  NO3        g178(.A(i_11_), .B(new_new_n162_), .C(new_new_n25_), .Y(new_new_n201_));
  INV        g179(.A(new_new_n201_), .Y(new_new_n202_));
  NA3        g180(.A(i_6_), .B(new_new_n193_), .C(new_new_n163_), .Y(new_new_n203_));
  AOI210     g181(.A0(new_new_n203_), .A1(new_new_n202_), .B0(new_new_n45_), .Y(new_new_n204_));
  AOI210     g182(.A0(new_new_n200_), .A1(new_new_n193_), .B0(new_new_n204_), .Y(new_new_n205_));
  NA4        g183(.A(new_new_n205_), .B(new_new_n192_), .C(new_new_n180_), .D(new_new_n166_), .Y(new_new_n206_));
  NO3        g184(.A(i_12_), .B(new_new_n162_), .C(new_new_n37_), .Y(new_new_n207_));
  INV        g185(.A(new_new_n207_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n173_), .B(i_0_), .Y(new_new_n209_));
  NO2        g187(.A(i_3_), .B(i_10_), .Y(new_new_n210_));
  NA3        g188(.A(new_new_n210_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n211_));
  AN2        g189(.A(i_3_), .B(i_10_), .Y(new_new_n212_));
  NO2        g190(.A(i_5_), .B(new_new_n37_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n45_), .B(new_new_n26_), .Y(new_new_n214_));
  OAI220     g192(.A0(new_new_n211_), .A1(i_6_), .B0(i_3_), .B1(new_new_n208_), .Y(new_new_n215_));
  NO4        g193(.A(new_new_n215_), .B(new_new_n206_), .C(new_new_n156_), .D(new_new_n121_), .Y(new_new_n216_));
  NO3        g194(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n217_));
  NO2        g195(.A(i_2_), .B(i_3_), .Y(new_new_n218_));
  NO2        g196(.A(i_12_), .B(i_10_), .Y(new_new_n219_));
  NOi21      g197(.An(i_5_), .B(i_0_), .Y(new_new_n220_));
  NA3        g198(.A(new_new_n36_), .B(new_new_n70_), .C(i_8_), .Y(new_new_n221_));
  NO2        g199(.A(i_6_), .B(i_8_), .Y(new_new_n222_));
  NO2        g200(.A(i_1_), .B(i_7_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n75_), .B(new_new_n142_), .Y(new_new_n224_));
  AOI210     g202(.A0(new_new_n54_), .A1(i_3_), .B0(new_new_n118_), .Y(new_new_n225_));
  AOI210     g203(.A0(i_12_), .A1(new_new_n217_), .B0(new_new_n225_), .Y(new_new_n226_));
  NOi32      g204(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n227_));
  INV        g205(.A(new_new_n227_), .Y(new_new_n228_));
  NAi21      g206(.An(i_1_), .B(i_5_), .Y(new_new_n229_));
  OAI210     g207(.A0(i_9_), .A1(new_new_n115_), .B0(new_new_n179_), .Y(new_new_n230_));
  NAi41      g208(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n231_));
  OAI220     g209(.A0(new_new_n231_), .A1(new_new_n229_), .B0(new_new_n160_), .B1(new_new_n115_), .Y(new_new_n232_));
  AOI210     g210(.A0(new_new_n231_), .A1(new_new_n115_), .B0(new_new_n113_), .Y(new_new_n233_));
  NOi32      g211(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n234_), .B(new_new_n45_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n235_), .B(i_0_), .Y(new_new_n236_));
  OR3        g214(.A(new_new_n236_), .B(new_new_n233_), .C(new_new_n232_), .Y(new_new_n237_));
  NAi21      g215(.An(i_3_), .B(i_4_), .Y(new_new_n238_));
  NO2        g216(.A(new_new_n238_), .B(i_9_), .Y(new_new_n239_));
  INV        g217(.A(new_new_n239_), .Y(new_new_n240_));
  NA2        g218(.A(i_2_), .B(i_7_), .Y(new_new_n241_));
  NO2        g219(.A(new_new_n238_), .B(i_10_), .Y(new_new_n242_));
  NA3        g220(.A(new_new_n242_), .B(new_new_n241_), .C(new_new_n177_), .Y(new_new_n243_));
  AOI210     g221(.A0(new_new_n243_), .A1(new_new_n240_), .B0(new_new_n135_), .Y(new_new_n244_));
  AOI210     g222(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n245_));
  INV        g223(.A(new_new_n242_), .Y(new_new_n246_));
  AOI220     g224(.A0(new_new_n242_), .A1(new_new_n223_), .B0(new_new_n172_), .B1(new_new_n138_), .Y(new_new_n247_));
  AOI210     g225(.A0(new_new_n247_), .A1(new_new_n246_), .B0(i_5_), .Y(new_new_n248_));
  NO4        g226(.A(new_new_n248_), .B(new_new_n244_), .C(new_new_n237_), .D(new_new_n230_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n249_), .B(new_new_n228_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n55_), .B(new_new_n25_), .Y(new_new_n251_));
  AN2        g229(.A(i_12_), .B(i_5_), .Y(new_new_n252_));
  NO2        g230(.A(i_4_), .B(new_new_n26_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n253_), .B(new_new_n252_), .Y(new_new_n254_));
  NO2        g232(.A(i_11_), .B(new_new_n254_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n176_), .B(i_5_), .Y(new_new_n256_));
  NO2        g234(.A(i_5_), .B(i_10_), .Y(new_new_n257_));
  NO2        g235(.A(i_11_), .B(new_new_n176_), .Y(new_new_n258_));
  OAI210     g236(.A0(new_new_n258_), .A1(new_new_n255_), .B0(new_new_n251_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n108_), .B(new_new_n70_), .Y(new_new_n261_));
  OAI210     g239(.A0(new_new_n261_), .A1(new_new_n255_), .B0(new_new_n260_), .Y(new_new_n262_));
  NO3        g240(.A(new_new_n70_), .B(new_new_n47_), .C(i_9_), .Y(new_new_n263_));
  NO2        g241(.A(i_11_), .B(i_12_), .Y(new_new_n264_));
  NO2        g242(.A(i_10_), .B(i_11_), .Y(new_new_n265_));
  NAi21      g243(.An(i_13_), .B(i_0_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n266_), .B(new_new_n173_), .Y(new_new_n267_));
  OAI210     g245(.A0(new_new_n740_), .A1(new_new_n265_), .B0(new_new_n267_), .Y(new_new_n268_));
  NA3        g246(.A(new_new_n268_), .B(new_new_n262_), .C(new_new_n259_), .Y(new_new_n269_));
  NO2        g247(.A(i_0_), .B(i_11_), .Y(new_new_n270_));
  AN2        g248(.A(i_1_), .B(i_6_), .Y(new_new_n271_));
  NOi21      g249(.An(i_2_), .B(i_12_), .Y(new_new_n272_));
  NA2        g250(.A(new_new_n100_), .B(i_9_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n273_), .B(i_4_), .Y(new_new_n274_));
  NA2        g252(.A(new_new_n272_), .B(new_new_n274_), .Y(new_new_n275_));
  OR2        g253(.A(i_13_), .B(i_10_), .Y(new_new_n276_));
  NO3        g254(.A(new_new_n276_), .B(new_new_n87_), .C(i_9_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n124_), .B(new_new_n89_), .Y(new_new_n278_));
  BUFFER     g256(.A(new_new_n157_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n79_), .B(new_new_n25_), .Y(new_new_n280_));
  NA2        g258(.A(new_new_n207_), .B(new_new_n280_), .Y(new_new_n281_));
  NA2        g259(.A(i_5_), .B(i_1_), .Y(new_new_n282_));
  OAI220     g260(.A0(new_new_n282_), .A1(new_new_n279_), .B0(new_new_n281_), .B1(new_new_n80_), .Y(new_new_n283_));
  INV        g261(.A(new_new_n283_), .Y(new_new_n284_));
  AOI210     g262(.A0(new_new_n284_), .A1(new_new_n275_), .B0(new_new_n26_), .Y(new_new_n285_));
  NO4        g263(.A(new_new_n748_), .B(new_new_n285_), .C(new_new_n269_), .D(new_new_n250_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n61_), .B(i_13_), .Y(new_new_n287_));
  NO2        g265(.A(i_10_), .B(i_9_), .Y(new_new_n288_));
  NO2        g266(.A(i_12_), .B(i_3_), .Y(new_new_n289_));
  NO2        g267(.A(i_4_), .B(new_new_n150_), .Y(new_new_n290_));
  NO3        g268(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n291_));
  NA2        g269(.A(new_new_n194_), .B(new_new_n77_), .Y(new_new_n292_));
  NA2        g270(.A(new_new_n292_), .B(new_new_n291_), .Y(new_new_n293_));
  NA2        g271(.A(i_8_), .B(i_9_), .Y(new_new_n294_));
  INV        g272(.A(new_new_n207_), .Y(new_new_n295_));
  OAI220     g273(.A0(new_new_n295_), .A1(new_new_n294_), .B0(new_new_n293_), .B1(new_new_n214_), .Y(new_new_n296_));
  NA2        g274(.A(new_new_n181_), .B(new_new_n213_), .Y(new_new_n297_));
  NO3        g275(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n298_));
  AOI210     g276(.A0(new_new_n184_), .A1(new_new_n138_), .B0(new_new_n298_), .Y(new_new_n299_));
  NA3        g277(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n300_));
  NA4        g278(.A(new_new_n103_), .B(new_new_n86_), .C(new_new_n66_), .D(new_new_n23_), .Y(new_new_n301_));
  OAI220     g279(.A0(new_new_n301_), .A1(new_new_n300_), .B0(new_new_n299_), .B1(new_new_n297_), .Y(new_new_n302_));
  NO3        g280(.A(new_new_n302_), .B(new_new_n296_), .C(new_new_n290_), .Y(new_new_n303_));
  OR2        g281(.A(i_8_), .B(new_new_n169_), .Y(new_new_n304_));
  NA2        g282(.A(new_new_n76_), .B(i_13_), .Y(new_new_n305_));
  NA2        g283(.A(i_3_), .B(new_new_n251_), .Y(new_new_n306_));
  NO2        g284(.A(i_2_), .B(i_13_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n306_), .B(new_new_n305_), .Y(new_new_n308_));
  NO3        g286(.A(i_4_), .B(new_new_n47_), .C(i_8_), .Y(new_new_n309_));
  NO2        g287(.A(i_6_), .B(i_7_), .Y(new_new_n310_));
  NO2        g288(.A(i_11_), .B(i_1_), .Y(new_new_n311_));
  OR2        g289(.A(i_11_), .B(i_8_), .Y(new_new_n312_));
  NOi21      g290(.An(i_2_), .B(i_7_), .Y(new_new_n313_));
  NAi31      g291(.An(new_new_n312_), .B(new_new_n313_), .C(i_0_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n276_), .B(new_new_n314_), .Y(new_new_n315_));
  NO2        g293(.A(i_6_), .B(i_10_), .Y(new_new_n316_));
  NA3        g294(.A(new_new_n178_), .B(new_new_n123_), .C(new_new_n95_), .Y(new_new_n317_));
  NO2        g295(.A(new_new_n113_), .B(i_3_), .Y(new_new_n318_));
  NAi31      g296(.An(i_11_), .B(new_new_n318_), .C(new_new_n163_), .Y(new_new_n319_));
  NA3        g297(.A(new_new_n260_), .B(new_new_n131_), .C(new_new_n107_), .Y(new_new_n320_));
  NA3        g298(.A(new_new_n320_), .B(new_new_n319_), .C(new_new_n317_), .Y(new_new_n321_));
  NO4        g299(.A(new_new_n321_), .B(new_new_n217_), .C(new_new_n315_), .D(new_new_n308_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n291_), .B(new_new_n252_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n298_), .B(new_new_n257_), .Y(new_new_n324_));
  INV        g302(.A(new_new_n323_), .Y(new_new_n325_));
  NAi21      g303(.An(new_new_n157_), .B(new_new_n264_), .Y(new_new_n326_));
  NA3        g304(.A(i_6_), .B(i_3_), .C(new_new_n100_), .Y(new_new_n327_));
  OAI220     g305(.A0(new_new_n38_), .A1(new_new_n327_), .B0(i_1_), .B1(new_new_n326_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n27_), .B(i_10_), .Y(new_new_n329_));
  NA2        g307(.A(new_new_n217_), .B(new_new_n172_), .Y(new_new_n330_));
  OAI210     g308(.A0(new_new_n329_), .A1(new_new_n305_), .B0(new_new_n330_), .Y(new_new_n331_));
  NO3        g309(.A(new_new_n331_), .B(new_new_n328_), .C(new_new_n325_), .Y(new_new_n332_));
  NA4        g310(.A(new_new_n332_), .B(new_new_n322_), .C(new_new_n304_), .D(new_new_n303_), .Y(new_new_n333_));
  NA3        g311(.A(new_new_n212_), .B(new_new_n128_), .C(new_new_n126_), .Y(new_new_n334_));
  OAI210     g312(.A0(new_new_n211_), .A1(new_new_n741_), .B0(new_new_n334_), .Y(new_new_n335_));
  INV        g313(.A(new_new_n335_), .Y(new_new_n336_));
  NA2        g314(.A(new_new_n252_), .B(new_new_n162_), .Y(new_new_n337_));
  NA2        g315(.A(new_new_n227_), .B(new_new_n61_), .Y(new_new_n338_));
  NA2        g316(.A(i_6_), .B(new_new_n234_), .Y(new_new_n339_));
  AO210      g317(.A0(new_new_n338_), .A1(new_new_n337_), .B0(new_new_n339_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n36_), .B(i_8_), .Y(new_new_n341_));
  NAi31      g319(.An(new_new_n338_), .B(new_new_n316_), .C(new_new_n45_), .Y(new_new_n342_));
  INV        g320(.A(new_new_n277_), .Y(new_new_n343_));
  NA3        g321(.A(new_new_n343_), .B(new_new_n342_), .C(new_new_n340_), .Y(new_new_n344_));
  INV        g322(.A(new_new_n344_), .Y(new_new_n345_));
  NO2        g323(.A(i_7_), .B(new_new_n145_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n133_), .B(new_new_n70_), .Y(new_new_n347_));
  AOI210     g325(.A0(new_new_n347_), .A1(new_new_n346_), .B0(new_new_n278_), .Y(new_new_n348_));
  NA3        g326(.A(new_new_n348_), .B(new_new_n345_), .C(new_new_n336_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n276_), .B(new_new_n38_), .Y(new_new_n350_));
  NA2        g328(.A(new_new_n350_), .B(new_new_n253_), .Y(new_new_n351_));
  NO2        g329(.A(i_8_), .B(i_7_), .Y(new_new_n352_));
  INV        g330(.A(new_new_n161_), .Y(new_new_n353_));
  NA2        g331(.A(new_new_n43_), .B(i_10_), .Y(new_new_n354_));
  NO2        g332(.A(new_new_n354_), .B(i_6_), .Y(new_new_n355_));
  NA3        g333(.A(new_new_n355_), .B(new_new_n739_), .C(new_new_n352_), .Y(new_new_n356_));
  OAI210     g334(.A0(new_new_n133_), .A1(new_new_n190_), .B0(new_new_n305_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n357_), .B(new_new_n193_), .Y(new_new_n358_));
  NOi31      g336(.An(new_new_n209_), .B(new_new_n211_), .C(new_new_n741_), .Y(new_new_n359_));
  NA3        g337(.A(new_new_n212_), .B(new_new_n126_), .C(new_new_n76_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n113_), .B(i_5_), .Y(new_new_n361_));
  NA2        g339(.A(new_new_n361_), .B(new_new_n218_), .Y(new_new_n362_));
  NA2        g340(.A(new_new_n362_), .B(new_new_n360_), .Y(new_new_n363_));
  OAI210     g341(.A0(new_new_n363_), .A1(new_new_n359_), .B0(new_new_n298_), .Y(new_new_n364_));
  NA4        g342(.A(new_new_n364_), .B(new_new_n358_), .C(new_new_n356_), .D(new_new_n351_), .Y(new_new_n365_));
  NA2        g343(.A(new_new_n207_), .B(new_new_n69_), .Y(new_new_n366_));
  AOI210     g344(.A0(i_11_), .A1(new_new_n67_), .B0(new_new_n366_), .Y(new_new_n367_));
  NA2        g345(.A(i_0_), .B(new_new_n47_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n201_), .B(new_new_n367_), .Y(new_new_n369_));
  NO4        g347(.A(new_new_n182_), .B(new_new_n41_), .C(i_2_), .D(new_new_n47_), .Y(new_new_n370_));
  NO3        g348(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n371_));
  OA210      g349(.A0(new_new_n371_), .A1(new_new_n370_), .B0(new_new_n227_), .Y(new_new_n372_));
  NO2        g350(.A(new_new_n276_), .B(i_1_), .Y(new_new_n373_));
  NOi31      g351(.An(new_new_n373_), .B(new_new_n292_), .C(new_new_n61_), .Y(new_new_n374_));
  AN4        g352(.A(new_new_n374_), .B(new_new_n274_), .C(i_3_), .D(i_2_), .Y(new_new_n375_));
  INV        g353(.A(new_new_n129_), .Y(new_new_n376_));
  NO3        g354(.A(new_new_n376_), .B(new_new_n375_), .C(new_new_n372_), .Y(new_new_n377_));
  NO2        g355(.A(new_new_n70_), .B(new_new_n25_), .Y(new_new_n378_));
  AOI220     g356(.A0(new_new_n207_), .A1(new_new_n378_), .B0(new_new_n201_), .B1(i_6_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n214_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n85_), .B(new_new_n23_), .Y(new_new_n381_));
  NA2        g359(.A(new_new_n124_), .B(new_new_n132_), .Y(new_new_n382_));
  NOi21      g360(.An(new_new_n104_), .B(new_new_n221_), .Y(new_new_n383_));
  NO3        g361(.A(new_new_n383_), .B(new_new_n382_), .C(new_new_n380_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n338_), .B(new_new_n247_), .Y(new_new_n385_));
  NA2        g363(.A(i_6_), .B(new_new_n201_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n207_), .B(new_new_n159_), .Y(new_new_n387_));
  AOI210     g365(.A0(new_new_n387_), .A1(new_new_n386_), .B0(i_3_), .Y(new_new_n388_));
  NO3        g366(.A(i_4_), .B(i_8_), .C(new_new_n211_), .Y(new_new_n389_));
  INV        g367(.A(new_new_n326_), .Y(new_new_n390_));
  NO4        g368(.A(new_new_n390_), .B(new_new_n389_), .C(new_new_n388_), .D(new_new_n385_), .Y(new_new_n391_));
  NA4        g369(.A(new_new_n391_), .B(new_new_n384_), .C(new_new_n377_), .D(new_new_n369_), .Y(new_new_n392_));
  NO4        g370(.A(new_new_n392_), .B(new_new_n365_), .C(new_new_n349_), .D(new_new_n333_), .Y(new_new_n393_));
  NA4        g371(.A(new_new_n393_), .B(new_new_n286_), .C(new_new_n226_), .D(new_new_n216_), .Y(zz07));
  NA2        g372(.A(new_new_n316_), .B(new_new_n69_), .Y(new_new_n395_));
  NA2        g373(.A(i_11_), .B(new_new_n142_), .Y(new_new_n396_));
  NO2        g374(.A(i_13_), .B(new_new_n395_), .Y(new_new_n397_));
  NA3        g375(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n171_), .B(i_4_), .Y(new_new_n399_));
  NA2        g377(.A(new_new_n399_), .B(i_8_), .Y(new_new_n400_));
  NA2        g378(.A(i_2_), .B(new_new_n70_), .Y(new_new_n401_));
  INV        g379(.A(new_new_n149_), .Y(new_new_n402_));
  NO2        g380(.A(i_7_), .B(new_new_n37_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n402_), .B(i_13_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n404_), .B(new_new_n397_), .Y(new_new_n405_));
  OR2        g383(.A(i_6_), .B(i_10_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n406_), .B(new_new_n23_), .Y(new_new_n407_));
  OR3        g385(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n408_));
  INV        g386(.A(new_new_n146_), .Y(new_new_n409_));
  OA220      g387(.A0(new_new_n408_), .A1(i_3_), .B0(i_10_), .B1(new_new_n195_), .Y(new_new_n410_));
  AOI210     g388(.A0(new_new_n410_), .A1(new_new_n405_), .B0(new_new_n56_), .Y(new_new_n411_));
  NOi21      g389(.An(i_11_), .B(i_7_), .Y(new_new_n412_));
  AO210      g390(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n413_), .B(new_new_n412_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n71_), .B(new_new_n56_), .Y(new_new_n415_));
  AO210      g393(.A0(new_new_n415_), .A1(new_new_n247_), .B0(new_new_n40_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n163_), .B(new_new_n56_), .Y(new_new_n417_));
  OR2        g395(.A(new_new_n152_), .B(new_new_n82_), .Y(new_new_n418_));
  NO2        g396(.A(new_new_n56_), .B(i_9_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n417_), .B(new_new_n416_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n420_), .B(i_6_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n171_), .B(new_new_n70_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n422_), .B(i_11_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n343_), .B(new_new_n293_), .Y(new_new_n424_));
  NO3        g402(.A(i_12_), .B(i_13_), .C(new_new_n70_), .Y(new_new_n425_));
  NA2        g403(.A(new_new_n425_), .B(new_new_n419_), .Y(new_new_n426_));
  NO3        g404(.A(new_new_n406_), .B(new_new_n170_), .C(new_new_n23_), .Y(new_new_n427_));
  AOI210     g405(.A0(i_1_), .A1(new_new_n187_), .B0(new_new_n427_), .Y(new_new_n428_));
  OAI210     g406(.A0(new_new_n428_), .A1(new_new_n43_), .B0(new_new_n426_), .Y(new_new_n429_));
  NA3        g407(.A(new_new_n352_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n430_));
  INV        g408(.A(i_2_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n97_), .B(i_9_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n432_), .B(new_new_n431_), .Y(new_new_n433_));
  NA3        g411(.A(new_new_n419_), .B(new_new_n218_), .C(i_6_), .Y(new_new_n434_));
  NO2        g412(.A(new_new_n434_), .B(new_new_n23_), .Y(new_new_n435_));
  AOI210     g413(.A0(new_new_n311_), .A1(new_new_n280_), .B0(new_new_n175_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n401_), .Y(new_new_n437_));
  NO2        g415(.A(i_11_), .B(new_new_n37_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n438_), .B(new_new_n24_), .Y(new_new_n439_));
  OR3        g417(.A(new_new_n437_), .B(new_new_n435_), .C(new_new_n433_), .Y(new_new_n440_));
  NO3        g418(.A(new_new_n440_), .B(new_new_n429_), .C(new_new_n424_), .Y(new_new_n441_));
  NO2        g419(.A(new_new_n171_), .B(new_new_n79_), .Y(new_new_n442_));
  NO2        g420(.A(new_new_n442_), .B(new_new_n412_), .Y(new_new_n443_));
  NO2        g421(.A(new_new_n757_), .B(new_new_n408_), .Y(new_new_n444_));
  NO2        g422(.A(i_9_), .B(new_new_n70_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n444_), .B(new_new_n45_), .Y(new_new_n446_));
  NA2        g424(.A(i_3_), .B(new_new_n142_), .Y(new_new_n447_));
  NA2        g425(.A(i_1_), .B(i_3_), .Y(new_new_n448_));
  NA3        g426(.A(new_new_n446_), .B(new_new_n441_), .C(new_new_n421_), .Y(new_new_n449_));
  AN2        g427(.A(new_new_n178_), .B(new_new_n70_), .Y(new_new_n450_));
  NA2        g428(.A(i_6_), .B(new_new_n239_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n316_), .B(new_new_n45_), .Y(new_new_n452_));
  NA2        g430(.A(i_6_), .B(new_new_n25_), .Y(new_new_n453_));
  NA3        g431(.A(new_new_n117_), .B(new_new_n69_), .C(new_new_n70_), .Y(new_new_n454_));
  NA4        g432(.A(new_new_n454_), .B(new_new_n453_), .C(new_new_n452_), .D(new_new_n451_), .Y(new_new_n455_));
  OAI210     g433(.A0(new_new_n455_), .A1(new_new_n450_), .B0(i_1_), .Y(new_new_n456_));
  AOI210     g434(.A0(new_new_n194_), .A1(new_new_n77_), .B0(i_1_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n238_), .B(i_2_), .Y(new_new_n458_));
  NA2        g436(.A(new_new_n458_), .B(new_new_n457_), .Y(new_new_n459_));
  OAI210     g437(.A0(new_new_n434_), .A1(i_12_), .B0(new_new_n459_), .Y(new_new_n460_));
  INV        g438(.A(new_new_n460_), .Y(new_new_n461_));
  AOI210     g439(.A0(new_new_n461_), .A1(new_new_n456_), .B0(i_13_), .Y(new_new_n462_));
  NA2        g440(.A(new_new_n307_), .B(new_new_n117_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n463_), .B(new_new_n43_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n51_), .B(i_12_), .Y(new_new_n465_));
  AOI210     g443(.A0(new_new_n178_), .A1(new_new_n94_), .B0(new_new_n445_), .Y(new_new_n466_));
  OAI220     g444(.A0(new_new_n466_), .A1(new_new_n40_), .B0(new_new_n736_), .B1(new_new_n75_), .Y(new_new_n467_));
  AOI210     g445(.A0(new_new_n464_), .A1(new_new_n222_), .B0(new_new_n467_), .Y(new_new_n468_));
  NOi31      g446(.An(new_new_n753_), .B(new_new_n395_), .C(new_new_n43_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n93_), .B(i_13_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n470_), .B(new_new_n457_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n59_), .B(new_new_n79_), .Y(new_new_n472_));
  NO3        g450(.A(new_new_n313_), .B(new_new_n171_), .C(new_new_n70_), .Y(new_new_n473_));
  NO2        g451(.A(new_new_n473_), .B(new_new_n472_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n474_), .B(new_new_n409_), .Y(new_new_n475_));
  NO3        g453(.A(new_new_n475_), .B(new_new_n471_), .C(new_new_n469_), .Y(new_new_n476_));
  NA3        g454(.A(new_new_n272_), .B(new_new_n403_), .C(new_new_n77_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n423_), .B(i_13_), .Y(new_new_n478_));
  NAi21      g456(.An(i_11_), .B(i_12_), .Y(new_new_n479_));
  NOi41      g457(.An(new_new_n84_), .B(new_new_n479_), .C(i_13_), .D(new_new_n70_), .Y(new_new_n480_));
  AOI210     g458(.A0(new_new_n755_), .A1(new_new_n217_), .B0(new_new_n480_), .Y(new_new_n481_));
  NA3        g459(.A(new_new_n481_), .B(new_new_n478_), .C(new_new_n477_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n482_), .B(new_new_n56_), .Y(new_new_n483_));
  NO2        g461(.A(i_2_), .B(i_12_), .Y(new_new_n484_));
  NO2        g462(.A(i_3_), .B(i_2_), .Y(new_new_n485_));
  NA3        g463(.A(new_new_n756_), .B(new_new_n44_), .C(new_new_n162_), .Y(new_new_n486_));
  NA4        g464(.A(new_new_n486_), .B(new_new_n483_), .C(new_new_n476_), .D(new_new_n468_), .Y(new_new_n487_));
  OR4        g465(.A(new_new_n487_), .B(new_new_n462_), .C(new_new_n449_), .D(new_new_n411_), .Y(zz05));
  AOI210     g466(.A0(new_new_n443_), .A1(new_new_n197_), .B0(new_new_n278_), .Y(new_new_n489_));
  AO210      g467(.A0(new_new_n24_), .A1(i_10_), .B0(new_new_n181_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n490_), .B(new_new_n484_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n400_), .B(i_11_), .Y(new_new_n492_));
  OAI210     g470(.A0(new_new_n403_), .A1(new_new_n72_), .B0(new_new_n492_), .Y(new_new_n493_));
  NA4        g471(.A(new_new_n493_), .B(new_new_n491_), .C(new_new_n489_), .D(new_new_n343_), .Y(new_new_n494_));
  NO3        g472(.A(i_11_), .B(new_new_n171_), .C(i_13_), .Y(new_new_n495_));
  NO2        g473(.A(new_new_n90_), .B(new_new_n23_), .Y(new_new_n496_));
  NA2        g474(.A(i_12_), .B(i_8_), .Y(new_new_n497_));
  OAI210     g475(.A0(new_new_n45_), .A1(i_3_), .B0(new_new_n497_), .Y(new_new_n498_));
  INV        g476(.A(new_new_n288_), .Y(new_new_n499_));
  AOI220     g477(.A0(new_new_n218_), .A1(new_new_n381_), .B0(new_new_n498_), .B1(new_new_n496_), .Y(new_new_n500_));
  INV        g478(.A(new_new_n500_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n501_), .B(new_new_n494_), .Y(new_new_n502_));
  INV        g480(.A(new_new_n123_), .Y(new_new_n503_));
  INV        g481(.A(new_new_n178_), .Y(new_new_n504_));
  OAI210     g482(.A0(new_new_n458_), .A1(new_new_n289_), .B0(new_new_n84_), .Y(new_new_n505_));
  AOI210     g483(.A0(new_new_n505_), .A1(new_new_n504_), .B0(new_new_n503_), .Y(new_new_n506_));
  NO2        g484(.A(new_new_n294_), .B(new_new_n26_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(new_new_n280_), .Y(new_new_n508_));
  NA2        g486(.A(new_new_n508_), .B(i_2_), .Y(new_new_n509_));
  INV        g487(.A(new_new_n509_), .Y(new_new_n510_));
  AOI210     g488(.A0(new_new_n754_), .A1(new_new_n510_), .B0(new_new_n506_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n139_), .B(new_new_n91_), .Y(new_new_n512_));
  OAI210     g490(.A0(new_new_n512_), .A1(new_new_n496_), .B0(i_2_), .Y(new_new_n513_));
  INV        g491(.A(new_new_n124_), .Y(new_new_n514_));
  NO3        g492(.A(new_new_n413_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n515_));
  AOI210     g493(.A0(new_new_n514_), .A1(new_new_n72_), .B0(new_new_n515_), .Y(new_new_n516_));
  AOI210     g494(.A0(new_new_n516_), .A1(new_new_n513_), .B0(new_new_n142_), .Y(new_new_n517_));
  OA210      g495(.A0(new_new_n414_), .A1(new_new_n92_), .B0(i_13_), .Y(new_new_n518_));
  INV        g496(.A(new_new_n146_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n109_), .B(new_new_n396_), .Y(new_new_n520_));
  AOI210     g498(.A0(new_new_n520_), .A1(new_new_n519_), .B0(new_new_n241_), .Y(new_new_n521_));
  AOI210     g499(.A0(new_new_n152_), .A1(new_new_n106_), .B0(new_new_n341_), .Y(new_new_n522_));
  OAI210     g500(.A0(new_new_n522_), .A1(new_new_n163_), .B0(new_new_n280_), .Y(new_new_n523_));
  NO2        g501(.A(i_2_), .B(new_new_n43_), .Y(new_new_n524_));
  NA3        g502(.A(new_new_n212_), .B(new_new_n90_), .C(new_new_n41_), .Y(new_new_n525_));
  OAI210     g503(.A0(new_new_n525_), .A1(new_new_n524_), .B0(new_new_n523_), .Y(new_new_n526_));
  NO4        g504(.A(new_new_n526_), .B(new_new_n521_), .C(new_new_n518_), .D(new_new_n517_), .Y(new_new_n527_));
  INV        g505(.A(new_new_n381_), .Y(new_new_n528_));
  NA2        g506(.A(new_new_n495_), .B(i_7_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n529_), .B(new_new_n528_), .Y(new_new_n530_));
  NO2        g508(.A(i_2_), .B(i_12_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n531_), .B(new_new_n92_), .Y(new_new_n532_));
  NO2        g510(.A(new_new_n532_), .B(new_new_n396_), .Y(new_new_n533_));
  AOI220     g511(.A0(new_new_n533_), .A1(new_new_n36_), .B0(new_new_n530_), .B1(new_new_n45_), .Y(new_new_n534_));
  NA4        g512(.A(new_new_n534_), .B(new_new_n527_), .C(new_new_n511_), .D(new_new_n502_), .Y(zz06));
  OAI210     g513(.A0(new_new_n25_), .A1(new_new_n742_), .B0(new_new_n485_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n160_), .B(i_11_), .Y(new_new_n537_));
  NO2        g515(.A(i_11_), .B(i_9_), .Y(new_new_n538_));
  OR2        g516(.A(new_new_n536_), .B(i_12_), .Y(new_new_n539_));
  NA2        g517(.A(new_new_n242_), .B(new_new_n223_), .Y(new_new_n540_));
  NA4        g518(.A(new_new_n415_), .B(new_new_n312_), .C(i_12_), .D(new_new_n540_), .Y(new_new_n541_));
  AOI220     g519(.A0(new_new_n143_), .A1(new_new_n538_), .B0(new_new_n541_), .B1(new_new_n61_), .Y(new_new_n542_));
  INV        g520(.A(new_new_n219_), .Y(new_new_n543_));
  AOI210     g521(.A0(new_new_n90_), .A1(i_5_), .B0(new_new_n543_), .Y(new_new_n544_));
  NA2        g522(.A(new_new_n737_), .B(new_new_n531_), .Y(new_new_n545_));
  AOI210     g523(.A0(new_new_n545_), .A1(new_new_n339_), .B0(new_new_n135_), .Y(new_new_n546_));
  INV        g524(.A(i_11_), .Y(new_new_n547_));
  NA3        g525(.A(new_new_n547_), .B(new_new_n310_), .C(new_new_n257_), .Y(new_new_n548_));
  NAi32      g526(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n549_));
  AOI210     g527(.A0(i_11_), .A1(i_11_), .B0(new_new_n549_), .Y(new_new_n550_));
  NA2        g528(.A(i_4_), .B(new_new_n371_), .Y(new_new_n551_));
  NAi31      g529(.An(new_new_n550_), .B(new_new_n551_), .C(new_new_n548_), .Y(new_new_n552_));
  OR3        g530(.A(new_new_n552_), .B(new_new_n546_), .C(new_new_n544_), .Y(new_new_n553_));
  NA3        g531(.A(new_new_n749_), .B(new_new_n184_), .C(i_7_), .Y(new_new_n554_));
  OR2        g532(.A(new_new_n414_), .B(new_new_n289_), .Y(new_new_n555_));
  NA2        g533(.A(new_new_n555_), .B(new_new_n105_), .Y(new_new_n556_));
  AO210      g534(.A0(new_new_n324_), .A1(new_new_n499_), .B0(new_new_n36_), .Y(new_new_n557_));
  NA3        g535(.A(new_new_n557_), .B(new_new_n556_), .C(new_new_n554_), .Y(new_new_n558_));
  AOI210     g536(.A0(new_new_n738_), .A1(new_new_n371_), .B0(new_new_n537_), .Y(new_new_n559_));
  NA3        g537(.A(new_new_n241_), .B(new_new_n172_), .C(new_new_n105_), .Y(new_new_n560_));
  OAI210     g538(.A0(new_new_n263_), .A1(new_new_n149_), .B0(new_new_n58_), .Y(new_new_n561_));
  NA4        g539(.A(new_new_n561_), .B(new_new_n560_), .C(new_new_n559_), .D(new_new_n402_), .Y(new_new_n562_));
  AO210      g540(.A0(new_new_n341_), .A1(new_new_n45_), .B0(new_new_n71_), .Y(new_new_n563_));
  NA3        g541(.A(new_new_n563_), .B(new_new_n316_), .C(new_new_n159_), .Y(new_new_n564_));
  AOI210     g542(.A0(new_new_n289_), .A1(new_new_n288_), .B0(new_new_n370_), .Y(new_new_n565_));
  NA3        g543(.A(new_new_n744_), .B(new_new_n219_), .C(i_7_), .Y(new_new_n566_));
  NA4        g544(.A(new_new_n566_), .B(new_new_n743_), .C(new_new_n565_), .D(new_new_n564_), .Y(new_new_n567_));
  NO4        g545(.A(new_new_n567_), .B(new_new_n562_), .C(new_new_n558_), .D(new_new_n553_), .Y(new_new_n568_));
  NA4        g546(.A(new_new_n568_), .B(new_new_n542_), .C(new_new_n539_), .D(new_new_n249_), .Y(zz03));
  NA2        g547(.A(i_12_), .B(i_10_), .Y(new_new_n570_));
  NA2        g548(.A(i_6_), .B(i_7_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n571_), .B(i_0_), .Y(new_new_n572_));
  NO2        g550(.A(i_11_), .B(new_new_n171_), .Y(new_new_n573_));
  OAI210     g551(.A0(new_new_n572_), .A1(new_new_n209_), .B0(new_new_n573_), .Y(new_new_n574_));
  NA3        g552(.A(new_new_n560_), .B(new_new_n402_), .C(new_new_n240_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n575_), .B(new_new_n39_), .Y(new_new_n576_));
  NO3        g554(.A(new_new_n418_), .B(new_new_n294_), .C(new_new_n94_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n272_), .B(new_new_n44_), .Y(new_new_n578_));
  NO2        g556(.A(new_new_n52_), .B(new_new_n577_), .Y(new_new_n579_));
  AOI210     g557(.A0(new_new_n579_), .A1(new_new_n576_), .B0(new_new_n47_), .Y(new_new_n580_));
  NO3        g558(.A(new_new_n245_), .B(new_new_n38_), .C(i_0_), .Y(new_new_n581_));
  INV        g559(.A(new_new_n581_), .Y(new_new_n582_));
  NA2        g560(.A(new_new_n753_), .B(new_new_n746_), .Y(new_new_n583_));
  NA2        g561(.A(i_0_), .B(i_5_), .Y(new_new_n584_));
  OAI220     g562(.A0(new_new_n584_), .A1(new_new_n583_), .B0(new_new_n582_), .B1(new_new_n56_), .Y(new_new_n585_));
  NOi21      g563(.An(i_5_), .B(i_9_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n586_), .B(new_new_n287_), .Y(new_new_n587_));
  NO3        g565(.A(new_new_n273_), .B(new_new_n194_), .C(new_new_n61_), .Y(new_new_n588_));
  NO2        g566(.A(new_new_n127_), .B(new_new_n106_), .Y(new_new_n589_));
  AOI210     g567(.A0(new_new_n589_), .A1(new_new_n177_), .B0(new_new_n588_), .Y(new_new_n590_));
  OAI220     g568(.A0(new_new_n590_), .A1(new_new_n741_), .B0(i_12_), .B1(new_new_n587_), .Y(new_new_n591_));
  NO4        g569(.A(new_new_n591_), .B(new_new_n585_), .C(new_new_n580_), .D(new_new_n751_), .Y(new_new_n592_));
  INV        g570(.A(new_new_n217_), .Y(new_new_n593_));
  OAI220     g571(.A0(new_new_n118_), .A1(i_0_), .B0(new_new_n593_), .B1(i_10_), .Y(new_new_n594_));
  INV        g572(.A(new_new_n594_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n378_), .B(i_0_), .Y(new_new_n596_));
  NO3        g574(.A(new_new_n596_), .B(new_new_n254_), .C(new_new_n72_), .Y(new_new_n597_));
  NO4        g575(.A(i_5_), .B(i_12_), .C(new_new_n276_), .D(new_new_n271_), .Y(new_new_n598_));
  AOI210     g576(.A0(new_new_n598_), .A1(i_11_), .B0(new_new_n597_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n495_), .B(new_new_n220_), .Y(new_new_n600_));
  OAI220     g578(.A0(i_6_), .A1(new_new_n600_), .B0(new_new_n439_), .B1(new_new_n353_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n183_), .B(new_new_n110_), .Y(new_new_n602_));
  NO4        g580(.A(new_new_n85_), .B(new_new_n54_), .C(new_new_n447_), .D(i_5_), .Y(new_new_n603_));
  AO220      g581(.A0(new_new_n603_), .A1(new_new_n43_), .B0(new_new_n602_), .B1(i_6_), .Y(new_new_n604_));
  NO2        g582(.A(i_3_), .B(new_new_n600_), .Y(new_new_n605_));
  NO3        g583(.A(new_new_n605_), .B(new_new_n604_), .C(new_new_n601_), .Y(new_new_n606_));
  NA3        g584(.A(new_new_n606_), .B(new_new_n599_), .C(new_new_n595_), .Y(new_new_n607_));
  NA2        g585(.A(i_11_), .B(i_9_), .Y(new_new_n608_));
  NO3        g586(.A(i_12_), .B(new_new_n608_), .C(new_new_n401_), .Y(new_new_n609_));
  AO220      g587(.A0(new_new_n609_), .A1(i_10_), .B0(new_new_n196_), .B1(new_new_n71_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n608_), .B(new_new_n61_), .Y(new_new_n611_));
  NO2        g589(.A(new_new_n127_), .B(i_0_), .Y(new_new_n612_));
  NA2        g590(.A(new_new_n310_), .B(new_new_n168_), .Y(new_new_n613_));
  OAI220     g591(.A0(i_12_), .A1(new_new_n587_), .B0(new_new_n613_), .B1(new_new_n127_), .Y(new_new_n614_));
  NO3        g592(.A(new_new_n614_), .B(new_new_n114_), .C(new_new_n610_), .Y(new_new_n615_));
  NA2        g593(.A(new_new_n438_), .B(i_1_), .Y(new_new_n616_));
  NO2        g594(.A(i_6_), .B(new_new_n616_), .Y(new_new_n617_));
  NA2        g595(.A(new_new_n123_), .B(new_new_n80_), .Y(new_new_n618_));
  NOi21      g596(.An(new_new_n138_), .B(new_new_n618_), .Y(new_new_n619_));
  NO2        g597(.A(i_0_), .B(new_new_n578_), .Y(new_new_n620_));
  NO3        g598(.A(new_new_n620_), .B(new_new_n619_), .C(new_new_n617_), .Y(new_new_n621_));
  NOi21      g599(.An(i_7_), .B(new_new_n479_), .Y(new_new_n622_));
  NA3        g600(.A(new_new_n622_), .B(new_new_n253_), .C(i_6_), .Y(new_new_n623_));
  OA210      g601(.A0(new_new_n618_), .A1(new_new_n339_), .B0(new_new_n623_), .Y(new_new_n624_));
  NO3        g602(.A(new_new_n266_), .B(new_new_n231_), .C(new_new_n229_), .Y(new_new_n625_));
  INV        g603(.A(new_new_n188_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n479_), .B(new_new_n185_), .Y(new_new_n627_));
  AOI210     g605(.A0(new_new_n627_), .A1(new_new_n626_), .B0(new_new_n625_), .Y(new_new_n628_));
  NA4        g606(.A(new_new_n628_), .B(new_new_n624_), .C(new_new_n621_), .D(new_new_n615_), .Y(new_new_n629_));
  AN2        g607(.A(new_new_n220_), .B(new_new_n589_), .Y(new_new_n630_));
  NA2        g608(.A(new_new_n630_), .B(i_10_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n570_), .B(new_new_n218_), .Y(new_new_n632_));
  OA210      g610(.A0(new_new_n310_), .A1(new_new_n161_), .B0(new_new_n309_), .Y(new_new_n633_));
  OAI210     g611(.A0(new_new_n633_), .A1(new_new_n632_), .B0(new_new_n611_), .Y(new_new_n634_));
  NA3        g612(.A(new_new_n309_), .B(new_new_n272_), .C(new_new_n44_), .Y(new_new_n635_));
  OAI210     g613(.A0(new_new_n118_), .A1(i_7_), .B0(new_new_n635_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n611_), .B(new_new_n212_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n137_), .B(new_new_n637_), .Y(new_new_n638_));
  AOI220     g616(.A0(new_new_n638_), .A1(new_new_n310_), .B0(new_new_n636_), .B1(new_new_n61_), .Y(new_new_n639_));
  NA3        g617(.A(i_5_), .B(new_new_n251_), .C(new_new_n422_), .Y(new_new_n640_));
  NA2        g618(.A(new_new_n75_), .B(new_new_n43_), .Y(new_new_n641_));
  NO2        g619(.A(new_new_n63_), .B(new_new_n497_), .Y(new_new_n642_));
  NA2        g620(.A(new_new_n642_), .B(new_new_n641_), .Y(new_new_n643_));
  AOI210     g621(.A0(new_new_n643_), .A1(new_new_n640_), .B0(new_new_n46_), .Y(new_new_n644_));
  NAi21      g622(.An(i_9_), .B(i_5_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n266_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n398_), .B(new_new_n81_), .Y(new_new_n647_));
  AOI220     g625(.A0(new_new_n647_), .A1(i_0_), .B0(new_new_n646_), .B1(new_new_n414_), .Y(new_new_n648_));
  OAI220     g626(.A0(new_new_n648_), .A1(new_new_n70_), .B0(i_0_), .B1(new_new_n124_), .Y(new_new_n649_));
  NO3        g627(.A(new_new_n649_), .B(new_new_n644_), .C(new_new_n344_), .Y(new_new_n650_));
  NA4        g628(.A(new_new_n650_), .B(new_new_n639_), .C(new_new_n634_), .D(new_new_n631_), .Y(new_new_n651_));
  NO3        g629(.A(new_new_n651_), .B(new_new_n629_), .C(new_new_n607_), .Y(new_new_n652_));
  INV        g630(.A(new_new_n479_), .Y(new_new_n653_));
  NO3        g631(.A(new_new_n81_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n654_));
  AO220      g632(.A0(new_new_n654_), .A1(new_new_n43_), .B0(new_new_n653_), .B1(new_new_n126_), .Y(new_new_n655_));
  AOI210     g633(.A0(i_12_), .A1(new_new_n451_), .B0(new_new_n618_), .Y(new_new_n656_));
  AOI210     g634(.A0(new_new_n655_), .A1(new_new_n224_), .B0(new_new_n656_), .Y(new_new_n657_));
  NA3        g635(.A(new_new_n104_), .B(new_new_n746_), .C(new_new_n61_), .Y(new_new_n658_));
  NO2        g636(.A(new_new_n551_), .B(new_new_n266_), .Y(new_new_n659_));
  NA2        g637(.A(new_new_n573_), .B(i_9_), .Y(new_new_n660_));
  AOI210     g638(.A0(i_0_), .A1(new_new_n327_), .B0(new_new_n660_), .Y(new_new_n661_));
  OAI210     g639(.A0(new_new_n177_), .A1(i_9_), .B0(new_new_n167_), .Y(new_new_n662_));
  NO2        g640(.A(new_new_n662_), .B(new_new_n110_), .Y(new_new_n663_));
  NO3        g641(.A(new_new_n663_), .B(new_new_n661_), .C(new_new_n659_), .Y(new_new_n664_));
  NA3        g642(.A(new_new_n664_), .B(new_new_n658_), .C(new_new_n657_), .Y(new_new_n665_));
  NA2        g643(.A(new_new_n220_), .B(new_new_n241_), .Y(new_new_n666_));
  AOI210     g644(.A0(new_new_n211_), .A1(new_new_n118_), .B0(new_new_n666_), .Y(new_new_n667_));
  INV        g645(.A(new_new_n667_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n374_), .B(new_new_n63_), .Y(new_new_n669_));
  NO3        g647(.A(new_new_n153_), .B(new_new_n252_), .C(i_0_), .Y(new_new_n670_));
  OAI210     g648(.A0(new_new_n670_), .A1(new_new_n64_), .B0(i_13_), .Y(new_new_n671_));
  INV        g649(.A(new_new_n159_), .Y(new_new_n672_));
  NO2        g650(.A(i_12_), .B(new_new_n409_), .Y(new_new_n673_));
  NA3        g651(.A(new_new_n673_), .B(i_7_), .C(new_new_n672_), .Y(new_new_n674_));
  NA4        g652(.A(new_new_n674_), .B(new_new_n671_), .C(new_new_n669_), .D(new_new_n668_), .Y(new_new_n675_));
  NO2        g653(.A(new_new_n176_), .B(new_new_n75_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n676_), .B(new_new_n653_), .Y(new_new_n677_));
  NA2        g655(.A(new_new_n749_), .B(new_new_n128_), .Y(new_new_n678_));
  OA220      g656(.A0(new_new_n678_), .A1(i_0_), .B0(new_new_n677_), .B1(i_5_), .Y(new_new_n679_));
  AOI210     g657(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n127_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n680_), .B(new_new_n633_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n407_), .B(new_new_n135_), .Y(new_new_n682_));
  NA2        g660(.A(new_new_n682_), .B(new_new_n360_), .Y(new_new_n683_));
  NO3        g661(.A(new_new_n578_), .B(new_new_n51_), .C(new_new_n47_), .Y(new_new_n684_));
  NA2        g662(.A(new_new_n323_), .B(new_new_n317_), .Y(new_new_n685_));
  NO3        g663(.A(new_new_n685_), .B(new_new_n684_), .C(new_new_n683_), .Y(new_new_n686_));
  NA3        g664(.A(new_new_n257_), .B(new_new_n123_), .C(new_new_n122_), .Y(new_new_n687_));
  INV        g665(.A(new_new_n687_), .Y(new_new_n688_));
  NOi31      g666(.An(new_new_n256_), .B(i_11_), .C(new_new_n173_), .Y(new_new_n689_));
  NO3        g667(.A(new_new_n608_), .B(new_new_n159_), .C(new_new_n139_), .Y(new_new_n690_));
  NO3        g668(.A(new_new_n690_), .B(new_new_n689_), .C(new_new_n688_), .Y(new_new_n691_));
  NA4        g669(.A(new_new_n691_), .B(new_new_n686_), .C(new_new_n681_), .D(new_new_n679_), .Y(new_new_n692_));
  NO3        g670(.A(new_new_n408_), .B(new_new_n368_), .C(i_7_), .Y(new_new_n693_));
  NA3        g671(.A(new_new_n573_), .B(new_new_n83_), .C(new_new_n90_), .Y(new_new_n694_));
  INV        g672(.A(new_new_n694_), .Y(new_new_n695_));
  AOI210     g673(.A0(new_new_n695_), .A1(i_6_), .B0(new_new_n693_), .Y(new_new_n696_));
  NAi21      g674(.An(new_new_n175_), .B(new_new_n176_), .Y(new_new_n697_));
  NO3        g675(.A(new_new_n173_), .B(i_0_), .C(i_12_), .Y(new_new_n698_));
  AOI220     g676(.A0(new_new_n698_), .A1(new_new_n697_), .B0(new_new_n257_), .B1(new_new_n128_), .Y(new_new_n699_));
  NO3        g677(.A(i_12_), .B(new_new_n430_), .C(new_new_n94_), .Y(new_new_n700_));
  NA2        g678(.A(new_new_n700_), .B(new_new_n159_), .Y(new_new_n701_));
  NA2        g679(.A(new_new_n307_), .B(new_new_n612_), .Y(new_new_n702_));
  NA4        g680(.A(new_new_n702_), .B(new_new_n701_), .C(new_new_n699_), .D(new_new_n696_), .Y(new_new_n703_));
  NO4        g681(.A(new_new_n703_), .B(new_new_n692_), .C(new_new_n675_), .D(new_new_n665_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n747_), .B(new_new_n151_), .Y(new_new_n705_));
  NO2        g683(.A(new_new_n300_), .B(new_new_n194_), .Y(new_new_n706_));
  NO2        g684(.A(new_new_n706_), .B(new_new_n598_), .Y(new_new_n707_));
  INV        g685(.A(new_new_n707_), .Y(new_new_n708_));
  AOI210     g686(.A0(new_new_n136_), .A1(new_new_n47_), .B0(new_new_n708_), .Y(new_new_n709_));
  AOI210     g687(.A0(new_new_n709_), .A1(new_new_n705_), .B0(new_new_n61_), .Y(new_new_n710_));
  NO2        g688(.A(new_new_n371_), .B(new_new_n248_), .Y(new_new_n711_));
  NO2        g689(.A(new_new_n711_), .B(new_new_n503_), .Y(new_new_n712_));
  INV        g690(.A(new_new_n622_), .Y(new_new_n713_));
  NO2        g691(.A(new_new_n713_), .B(new_new_n448_), .Y(new_new_n714_));
  INV        g692(.A(new_new_n53_), .Y(new_new_n715_));
  NA2        g693(.A(new_new_n715_), .B(new_new_n64_), .Y(new_new_n716_));
  NO2        g694(.A(new_new_n716_), .B(new_new_n171_), .Y(new_new_n717_));
  NO2        g695(.A(new_new_n717_), .B(new_new_n714_), .Y(new_new_n718_));
  OAI210     g696(.A0(new_new_n196_), .A1(new_new_n114_), .B0(new_new_n72_), .Y(new_new_n719_));
  NA3        g697(.A(new_new_n507_), .B(new_new_n209_), .C(new_new_n66_), .Y(new_new_n720_));
  AOI210     g698(.A0(new_new_n720_), .A1(new_new_n719_), .B0(i_11_), .Y(new_new_n721_));
  INV        g699(.A(new_new_n151_), .Y(new_new_n722_));
  NA2        g700(.A(i_0_), .B(i_5_), .Y(new_new_n723_));
  AOI210     g701(.A0(new_new_n722_), .A1(new_new_n519_), .B0(new_new_n723_), .Y(new_new_n724_));
  NO3        g702(.A(new_new_n55_), .B(new_new_n54_), .C(i_4_), .Y(new_new_n725_));
  OAI210     g703(.A0(new_new_n626_), .A1(new_new_n213_), .B0(new_new_n725_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n726_), .B(new_new_n479_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n550_), .B(new_new_n232_), .Y(new_new_n728_));
  NO2        g706(.A(new_new_n728_), .B(new_new_n40_), .Y(new_new_n729_));
  NO4        g707(.A(new_new_n729_), .B(new_new_n727_), .C(new_new_n724_), .D(new_new_n721_), .Y(new_new_n730_));
  OAI210     g708(.A0(new_new_n718_), .A1(i_4_), .B0(new_new_n730_), .Y(new_new_n731_));
  NO3        g709(.A(new_new_n731_), .B(new_new_n712_), .C(new_new_n710_), .Y(new_new_n732_));
  NA4        g710(.A(new_new_n732_), .B(new_new_n704_), .C(new_new_n652_), .D(new_new_n592_), .Y(zz04));
  INV        g711(.A(new_new_n465_), .Y(new_new_n736_));
  INV        g712(.A(i_9_), .Y(new_new_n737_));
  INV        g713(.A(i_11_), .Y(new_new_n738_));
  INV        g714(.A(new_new_n176_), .Y(new_new_n739_));
  INV        g715(.A(new_new_n160_), .Y(new_new_n740_));
  INV        g716(.A(i_5_), .Y(new_new_n741_));
  INV        g717(.A(i_9_), .Y(new_new_n742_));
  INV        g718(.A(new_new_n270_), .Y(new_new_n743_));
  INV        g719(.A(i_5_), .Y(new_new_n744_));
  INV        g720(.A(new_new_n64_), .Y(new_new_n745_));
  INV        g721(.A(i_9_), .Y(new_new_n746_));
  INV        g722(.A(i_10_), .Y(new_new_n747_));
  INV        g723(.A(new_new_n199_), .Y(new_new_n748_));
  INV        g724(.A(i_9_), .Y(new_new_n749_));
  INV        g725(.A(new_new_n88_), .Y(new_new_n750_));
  INV        g726(.A(new_new_n574_), .Y(new_new_n751_));
  INV        g727(.A(i_6_), .Y(new_new_n752_));
  INV        g728(.A(i_13_), .Y(new_new_n753_));
  INV        g729(.A(new_new_n276_), .Y(new_new_n754_));
  INV        g730(.A(i_6_), .Y(new_new_n755_));
  INV        g731(.A(i_1_), .Y(new_new_n756_));
  INV        g732(.A(i_1_), .Y(new_new_n757_));
endmodule


