//Benchmark atmr_9sym_175_0.0313

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n169_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  NA2        o002(.A(i_4_), .B(ori_ori_n12_), .Y(ori_ori_n13_));
  INV        o003(.A(i_5_), .Y(ori_ori_n14_));
  NOi21      o004(.An(i_3_), .B(i_7_), .Y(ori_ori_n15_));
  NA3        o005(.A(ori_ori_n15_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n16_));
  INV        o006(.A(i_0_), .Y(ori_ori_n17_));
  NOi21      o007(.An(i_1_), .B(i_3_), .Y(ori_ori_n18_));
  NA3        o008(.A(ori_ori_n18_), .B(ori_ori_n17_), .C(i_2_), .Y(ori_ori_n19_));
  AOI210     o009(.A0(ori_ori_n19_), .A1(ori_ori_n16_), .B0(ori_ori_n13_), .Y(ori_ori_n20_));
  INV        o010(.A(i_4_), .Y(ori_ori_n21_));
  NA2        o011(.A(i_0_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  INV        o012(.A(i_7_), .Y(ori_ori_n23_));
  NA3        o013(.A(i_6_), .B(i_5_), .C(ori_ori_n23_), .Y(ori_ori_n24_));
  NOi21      o014(.An(i_8_), .B(i_6_), .Y(ori_ori_n25_));
  NOi21      o015(.An(i_1_), .B(i_8_), .Y(ori_ori_n26_));
  AOI220     o016(.A0(ori_ori_n26_), .A1(i_2_), .B0(ori_ori_n25_), .B1(i_5_), .Y(ori_ori_n27_));
  AOI210     o017(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n22_), .Y(ori_ori_n28_));
  AOI210     o018(.A0(ori_ori_n28_), .A1(ori_ori_n11_), .B0(ori_ori_n20_), .Y(ori_ori_n29_));
  NO2        o019(.A(i_2_), .B(i_4_), .Y(ori_ori_n30_));
  INV        o020(.A(i_2_), .Y(ori_ori_n31_));
  NOi21      o021(.An(i_6_), .B(i_8_), .Y(ori_ori_n32_));
  NOi21      o022(.An(i_7_), .B(i_1_), .Y(ori_ori_n33_));
  NOi21      o023(.An(i_5_), .B(i_6_), .Y(ori_ori_n34_));
  AOI220     o024(.A0(ori_ori_n34_), .A1(ori_ori_n33_), .B0(ori_ori_n32_), .B1(i_5_), .Y(ori_ori_n35_));
  NO3        o025(.A(ori_ori_n35_), .B(ori_ori_n31_), .C(i_4_), .Y(ori_ori_n36_));
  NOi21      o026(.An(i_0_), .B(i_4_), .Y(ori_ori_n37_));
  XO2        o027(.A(i_1_), .B(i_3_), .Y(ori_ori_n38_));
  NOi21      o028(.An(i_7_), .B(i_5_), .Y(ori_ori_n39_));
  AN3        o029(.A(ori_ori_n39_), .B(ori_ori_n38_), .C(ori_ori_n37_), .Y(ori_ori_n40_));
  INV        o030(.A(i_1_), .Y(ori_ori_n41_));
  NOi21      o031(.An(i_3_), .B(i_0_), .Y(ori_ori_n42_));
  NA2        o032(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NO2        o033(.A(ori_ori_n169_), .B(ori_ori_n43_), .Y(ori_ori_n44_));
  NO3        o034(.A(ori_ori_n44_), .B(ori_ori_n40_), .C(ori_ori_n36_), .Y(ori_ori_n45_));
  NA2        o035(.A(i_1_), .B(ori_ori_n11_), .Y(ori_ori_n46_));
  NOi21      o036(.An(i_4_), .B(i_0_), .Y(ori_ori_n47_));
  NO2        o037(.A(ori_ori_n25_), .B(ori_ori_n15_), .Y(ori_ori_n48_));
  NA2        o038(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n49_));
  NOi21      o039(.An(i_2_), .B(i_8_), .Y(ori_ori_n50_));
  NO3        o040(.A(ori_ori_n50_), .B(ori_ori_n47_), .C(ori_ori_n37_), .Y(ori_ori_n51_));
  NO3        o041(.A(ori_ori_n51_), .B(ori_ori_n49_), .C(ori_ori_n48_), .Y(ori_ori_n52_));
  INV        o042(.A(ori_ori_n52_), .Y(ori_ori_n53_));
  NOi31      o043(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n54_));
  NA2        o044(.A(ori_ori_n54_), .B(i_0_), .Y(ori_ori_n55_));
  NOi21      o045(.An(i_4_), .B(i_3_), .Y(ori_ori_n56_));
  NOi21      o046(.An(i_1_), .B(i_4_), .Y(ori_ori_n57_));
  OAI210     o047(.A0(ori_ori_n57_), .A1(ori_ori_n56_), .B0(ori_ori_n50_), .Y(ori_ori_n58_));
  NA2        o048(.A(ori_ori_n58_), .B(ori_ori_n55_), .Y(ori_ori_n59_));
  AN2        o049(.A(i_8_), .B(i_7_), .Y(ori_ori_n60_));
  INV        o050(.A(ori_ori_n60_), .Y(ori_ori_n61_));
  NOi21      o051(.An(i_8_), .B(i_7_), .Y(ori_ori_n62_));
  NO2        o052(.A(ori_ori_n61_), .B(ori_ori_n49_), .Y(ori_ori_n63_));
  AOI220     o053(.A0(ori_ori_n63_), .A1(ori_ori_n31_), .B0(ori_ori_n59_), .B1(ori_ori_n34_), .Y(ori_ori_n64_));
  NA4        o054(.A(ori_ori_n64_), .B(ori_ori_n53_), .C(ori_ori_n45_), .D(ori_ori_n29_), .Y(ori_ori_n65_));
  NA2        o055(.A(i_8_), .B(i_7_), .Y(ori_ori_n66_));
  NO3        o056(.A(ori_ori_n66_), .B(ori_ori_n13_), .C(i_1_), .Y(ori_ori_n67_));
  NA2        o057(.A(i_8_), .B(ori_ori_n23_), .Y(ori_ori_n68_));
  AOI220     o058(.A0(ori_ori_n42_), .A1(i_1_), .B0(ori_ori_n38_), .B1(i_2_), .Y(ori_ori_n69_));
  NOi21      o059(.An(i_1_), .B(i_2_), .Y(ori_ori_n70_));
  NO2        o060(.A(ori_ori_n69_), .B(ori_ori_n68_), .Y(ori_ori_n71_));
  OAI210     o061(.A0(ori_ori_n71_), .A1(ori_ori_n67_), .B0(ori_ori_n14_), .Y(ori_ori_n72_));
  NA3        o062(.A(ori_ori_n62_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n73_));
  NA3        o063(.A(ori_ori_n26_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n74_));
  NA2        o064(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  NOi32      o065(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(ori_ori_n76_));
  NA2        o066(.A(ori_ori_n76_), .B(i_3_), .Y(ori_ori_n77_));
  NA3        o067(.A(ori_ori_n18_), .B(i_2_), .C(i_6_), .Y(ori_ori_n78_));
  NA2        o068(.A(ori_ori_n78_), .B(ori_ori_n77_), .Y(ori_ori_n79_));
  NO2        o069(.A(i_0_), .B(i_4_), .Y(ori_ori_n80_));
  AOI220     o070(.A0(ori_ori_n80_), .A1(ori_ori_n79_), .B0(ori_ori_n75_), .B1(ori_ori_n56_), .Y(ori_ori_n81_));
  NA2        o071(.A(ori_ori_n81_), .B(ori_ori_n72_), .Y(ori_ori_n82_));
  INV        o072(.A(i_6_), .Y(ori_ori_n83_));
  NO2        o073(.A(ori_ori_n83_), .B(i_0_), .Y(ori_ori_n84_));
  NOi21      o074(.An(i_7_), .B(i_8_), .Y(ori_ori_n85_));
  NOi21      o075(.An(i_6_), .B(i_5_), .Y(ori_ori_n86_));
  AOI210     o076(.A0(ori_ori_n85_), .A1(ori_ori_n12_), .B0(ori_ori_n86_), .Y(ori_ori_n87_));
  NO2        o077(.A(ori_ori_n87_), .B(ori_ori_n11_), .Y(ori_ori_n88_));
  OAI210     o078(.A0(ori_ori_n88_), .A1(ori_ori_n84_), .B0(ori_ori_n70_), .Y(ori_ori_n89_));
  NA3        o079(.A(ori_ori_n25_), .B(i_2_), .C(ori_ori_n14_), .Y(ori_ori_n90_));
  AOI210     o080(.A0(ori_ori_n22_), .A1(ori_ori_n46_), .B0(ori_ori_n90_), .Y(ori_ori_n91_));
  AOI220     o081(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n18_), .B1(ori_ori_n31_), .Y(ori_ori_n92_));
  NA3        o082(.A(ori_ori_n21_), .B(i_5_), .C(i_7_), .Y(ori_ori_n93_));
  NA2        o083(.A(i_4_), .B(i_5_), .Y(ori_ori_n94_));
  NA3        o084(.A(ori_ori_n66_), .B(ori_ori_n18_), .C(ori_ori_n17_), .Y(ori_ori_n95_));
  OAI220     o085(.A0(ori_ori_n95_), .A1(ori_ori_n94_), .B0(ori_ori_n93_), .B1(ori_ori_n92_), .Y(ori_ori_n96_));
  NO2        o086(.A(ori_ori_n96_), .B(ori_ori_n91_), .Y(ori_ori_n97_));
  NA2        o087(.A(ori_ori_n41_), .B(i_6_), .Y(ori_ori_n98_));
  NOi21      o088(.An(i_2_), .B(i_1_), .Y(ori_ori_n99_));
  AN3        o089(.A(ori_ori_n85_), .B(ori_ori_n99_), .C(ori_ori_n47_), .Y(ori_ori_n100_));
  NAi21      o090(.An(i_6_), .B(i_0_), .Y(ori_ori_n101_));
  NA3        o091(.A(ori_ori_n57_), .B(i_5_), .C(ori_ori_n23_), .Y(ori_ori_n102_));
  NOi21      o092(.An(i_4_), .B(i_6_), .Y(ori_ori_n103_));
  NOi21      o093(.An(i_5_), .B(i_3_), .Y(ori_ori_n104_));
  NA3        o094(.A(ori_ori_n104_), .B(ori_ori_n70_), .C(ori_ori_n103_), .Y(ori_ori_n105_));
  OAI210     o095(.A0(ori_ori_n102_), .A1(ori_ori_n101_), .B0(ori_ori_n105_), .Y(ori_ori_n106_));
  NA2        o096(.A(ori_ori_n70_), .B(ori_ori_n32_), .Y(ori_ori_n107_));
  NO2        o097(.A(ori_ori_n106_), .B(ori_ori_n100_), .Y(ori_ori_n108_));
  BUFFER     o098(.A(i_6_), .Y(ori_ori_n109_));
  AOI210     o099(.A0(ori_ori_n109_), .A1(i_7_), .B0(i_5_), .Y(ori_ori_n110_));
  NOi31      o100(.An(ori_ori_n47_), .B(ori_ori_n110_), .C(i_2_), .Y(ori_ori_n111_));
  NA2        o101(.A(ori_ori_n62_), .B(ori_ori_n12_), .Y(ori_ori_n112_));
  NA2        o102(.A(ori_ori_n32_), .B(ori_ori_n14_), .Y(ori_ori_n113_));
  NOi21      o103(.An(i_3_), .B(i_1_), .Y(ori_ori_n114_));
  NA2        o104(.A(ori_ori_n114_), .B(i_4_), .Y(ori_ori_n115_));
  AOI210     o105(.A0(ori_ori_n113_), .A1(ori_ori_n112_), .B0(ori_ori_n115_), .Y(ori_ori_n116_));
  AOI220     o106(.A0(ori_ori_n85_), .A1(ori_ori_n14_), .B0(ori_ori_n103_), .B1(ori_ori_n23_), .Y(ori_ori_n117_));
  NOi31      o107(.An(ori_ori_n42_), .B(ori_ori_n117_), .C(ori_ori_n31_), .Y(ori_ori_n118_));
  NO3        o108(.A(ori_ori_n118_), .B(ori_ori_n116_), .C(ori_ori_n111_), .Y(ori_ori_n119_));
  NA4        o109(.A(ori_ori_n119_), .B(ori_ori_n108_), .C(ori_ori_n97_), .D(ori_ori_n89_), .Y(ori_ori_n120_));
  NA2        o110(.A(ori_ori_n50_), .B(ori_ori_n15_), .Y(ori_ori_n121_));
  NOi31      o111(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n122_));
  NOi31      o112(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n123_));
  OAI210     o113(.A0(ori_ori_n123_), .A1(ori_ori_n122_), .B0(i_7_), .Y(ori_ori_n124_));
  NA3        o114(.A(ori_ori_n32_), .B(i_2_), .C(ori_ori_n14_), .Y(ori_ori_n125_));
  NA4        o115(.A(ori_ori_n125_), .B(ori_ori_n124_), .C(ori_ori_n121_), .D(ori_ori_n107_), .Y(ori_ori_n126_));
  NA2        o116(.A(ori_ori_n126_), .B(ori_ori_n37_), .Y(ori_ori_n127_));
  NA3        o117(.A(ori_ori_n60_), .B(ori_ori_n99_), .C(ori_ori_n17_), .Y(ori_ori_n128_));
  NAi31      o118(.An(ori_ori_n101_), .B(ori_ori_n85_), .C(ori_ori_n99_), .Y(ori_ori_n129_));
  NA3        o119(.A(ori_ori_n62_), .B(ori_ori_n54_), .C(i_6_), .Y(ori_ori_n130_));
  NA3        o120(.A(ori_ori_n130_), .B(ori_ori_n129_), .C(ori_ori_n128_), .Y(ori_ori_n131_));
  NOi21      o121(.An(i_0_), .B(i_2_), .Y(ori_ori_n132_));
  NA3        o122(.A(ori_ori_n132_), .B(ori_ori_n33_), .C(ori_ori_n103_), .Y(ori_ori_n133_));
  NA3        o123(.A(ori_ori_n47_), .B(ori_ori_n39_), .C(ori_ori_n18_), .Y(ori_ori_n134_));
  NOi32      o124(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n135_));
  NA2        o125(.A(ori_ori_n135_), .B(ori_ori_n122_), .Y(ori_ori_n136_));
  NA3        o126(.A(ori_ori_n132_), .B(ori_ori_n56_), .C(ori_ori_n32_), .Y(ori_ori_n137_));
  NA4        o127(.A(ori_ori_n137_), .B(ori_ori_n136_), .C(ori_ori_n134_), .D(ori_ori_n133_), .Y(ori_ori_n138_));
  NA4        o128(.A(ori_ori_n54_), .B(i_6_), .C(ori_ori_n14_), .D(i_7_), .Y(ori_ori_n139_));
  NA4        o129(.A(ori_ori_n57_), .B(ori_ori_n34_), .C(ori_ori_n17_), .D(i_8_), .Y(ori_ori_n140_));
  NA2        o130(.A(ori_ori_n140_), .B(ori_ori_n139_), .Y(ori_ori_n141_));
  NO3        o131(.A(ori_ori_n141_), .B(ori_ori_n138_), .C(ori_ori_n131_), .Y(ori_ori_n142_));
  NOi21      o132(.An(i_5_), .B(i_2_), .Y(ori_ori_n143_));
  AOI220     o133(.A0(ori_ori_n143_), .A1(ori_ori_n85_), .B0(ori_ori_n60_), .B1(ori_ori_n30_), .Y(ori_ori_n144_));
  NO2        o134(.A(ori_ori_n144_), .B(ori_ori_n98_), .Y(ori_ori_n145_));
  NO3        o135(.A(i_2_), .B(ori_ori_n11_), .C(ori_ori_n14_), .Y(ori_ori_n146_));
  NA2        o136(.A(i_2_), .B(i_4_), .Y(ori_ori_n147_));
  AOI210     o137(.A0(ori_ori_n101_), .A1(ori_ori_n83_), .B0(ori_ori_n147_), .Y(ori_ori_n148_));
  NO2        o138(.A(i_8_), .B(i_7_), .Y(ori_ori_n149_));
  OA210      o139(.A0(ori_ori_n148_), .A1(ori_ori_n146_), .B0(ori_ori_n149_), .Y(ori_ori_n150_));
  NA3        o140(.A(ori_ori_n114_), .B(i_5_), .C(ori_ori_n23_), .Y(ori_ori_n151_));
  NO2        o141(.A(ori_ori_n151_), .B(i_4_), .Y(ori_ori_n152_));
  NO3        o142(.A(ori_ori_n152_), .B(ori_ori_n150_), .C(ori_ori_n145_), .Y(ori_ori_n153_));
  NA2        o143(.A(ori_ori_n85_), .B(ori_ori_n12_), .Y(ori_ori_n154_));
  NA3        o144(.A(i_2_), .B(i_1_), .C(ori_ori_n14_), .Y(ori_ori_n155_));
  NA2        o145(.A(ori_ori_n47_), .B(i_3_), .Y(ori_ori_n156_));
  AOI210     o146(.A0(ori_ori_n156_), .A1(ori_ori_n155_), .B0(ori_ori_n154_), .Y(ori_ori_n157_));
  NA2        o147(.A(ori_ori_n132_), .B(ori_ori_n62_), .Y(ori_ori_n158_));
  INV        o148(.A(ori_ori_n158_), .Y(ori_ori_n159_));
  NA4        o149(.A(ori_ori_n104_), .B(ori_ori_n60_), .C(ori_ori_n41_), .D(ori_ori_n21_), .Y(ori_ori_n160_));
  NOi31      o150(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n161_));
  OAI210     o151(.A0(ori_ori_n135_), .A1(ori_ori_n76_), .B0(ori_ori_n161_), .Y(ori_ori_n162_));
  NA2        o152(.A(ori_ori_n162_), .B(ori_ori_n160_), .Y(ori_ori_n163_));
  NO3        o153(.A(ori_ori_n163_), .B(ori_ori_n159_), .C(ori_ori_n157_), .Y(ori_ori_n164_));
  NA4        o154(.A(ori_ori_n164_), .B(ori_ori_n153_), .C(ori_ori_n142_), .D(ori_ori_n127_), .Y(ori_ori_n165_));
  OR4        o155(.A(ori_ori_n165_), .B(ori_ori_n120_), .C(ori_ori_n82_), .D(ori_ori_n65_), .Y(ori00));
  INV        o156(.A(i_6_), .Y(ori_ori_n169_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NA3        m013(.A(i_6_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_8_), .B(i_6_), .Y(mai_mai_n25_));
  NOi21      m015(.An(i_1_), .B(i_8_), .Y(mai_mai_n26_));
  AOI220     m016(.A0(mai_mai_n26_), .A1(i_2_), .B0(mai_mai_n25_), .B1(i_5_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n22_), .Y(mai_mai_n28_));
  AOI210     m018(.A0(mai_mai_n28_), .A1(mai_mai_n11_), .B0(mai_mai_n20_), .Y(mai_mai_n29_));
  NA2        m019(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n30_));
  NA2        m020(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n31_));
  NO2        m021(.A(i_2_), .B(i_4_), .Y(mai_mai_n32_));
  NA3        m022(.A(mai_mai_n32_), .B(i_6_), .C(i_8_), .Y(mai_mai_n33_));
  AOI210     m023(.A0(mai_mai_n31_), .A1(mai_mai_n30_), .B0(mai_mai_n33_), .Y(mai_mai_n34_));
  INV        m024(.A(i_2_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_5_), .B(i_0_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_6_), .B(i_8_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_5_), .B(i_6_), .Y(mai_mai_n38_));
  NA2        m028(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n39_));
  NO2        m029(.A(mai_mai_n39_), .B(mai_mai_n35_), .Y(mai_mai_n40_));
  NOi21      m030(.An(i_0_), .B(i_4_), .Y(mai_mai_n41_));
  XO2        m031(.A(i_1_), .B(i_3_), .Y(mai_mai_n42_));
  NOi21      m032(.An(i_7_), .B(i_5_), .Y(mai_mai_n43_));
  AN3        m033(.A(mai_mai_n43_), .B(mai_mai_n42_), .C(mai_mai_n41_), .Y(mai_mai_n44_));
  INV        m034(.A(i_1_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_3_), .B(i_0_), .Y(mai_mai_n46_));
  NA2        m036(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m037(.A(mai_mai_n24_), .B(mai_mai_n47_), .Y(mai_mai_n48_));
  NO4        m038(.A(mai_mai_n48_), .B(mai_mai_n44_), .C(mai_mai_n40_), .D(mai_mai_n34_), .Y(mai_mai_n49_));
  INV        m039(.A(i_8_), .Y(mai_mai_n50_));
  NA2        m040(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n51_));
  NO4        m041(.A(mai_mai_n51_), .B(mai_mai_n30_), .C(i_2_), .D(mai_mai_n50_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_4_), .B(i_0_), .Y(mai_mai_n53_));
  AOI210     m043(.A0(mai_mai_n53_), .A1(mai_mai_n25_), .B0(mai_mai_n15_), .Y(mai_mai_n54_));
  NA2        m044(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n55_));
  NOi21      m045(.An(i_2_), .B(i_8_), .Y(mai_mai_n56_));
  NO3        m046(.A(mai_mai_n56_), .B(mai_mai_n53_), .C(mai_mai_n41_), .Y(mai_mai_n57_));
  NO3        m047(.A(mai_mai_n57_), .B(mai_mai_n55_), .C(mai_mai_n54_), .Y(mai_mai_n58_));
  NO2        m048(.A(mai_mai_n58_), .B(mai_mai_n52_), .Y(mai_mai_n59_));
  NOi31      m049(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n60_));
  NOi21      m050(.An(i_4_), .B(i_3_), .Y(mai_mai_n61_));
  NOi21      m051(.An(i_1_), .B(i_4_), .Y(mai_mai_n62_));
  AN2        m052(.A(i_8_), .B(i_7_), .Y(mai_mai_n63_));
  NA2        m053(.A(mai_mai_n63_), .B(mai_mai_n12_), .Y(mai_mai_n64_));
  NOi21      m054(.An(i_8_), .B(i_7_), .Y(mai_mai_n65_));
  NA3        m055(.A(mai_mai_n65_), .B(mai_mai_n61_), .C(i_6_), .Y(mai_mai_n66_));
  OAI210     m056(.A0(mai_mai_n64_), .A1(mai_mai_n55_), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  AOI220     m057(.A0(mai_mai_n67_), .A1(mai_mai_n35_), .B0(mai_mai_n56_), .B1(mai_mai_n38_), .Y(mai_mai_n68_));
  NA4        m058(.A(mai_mai_n68_), .B(mai_mai_n59_), .C(mai_mai_n49_), .D(mai_mai_n29_), .Y(mai_mai_n69_));
  INV        m059(.A(i_7_), .Y(mai_mai_n70_));
  NO3        m060(.A(mai_mai_n70_), .B(mai_mai_n13_), .C(i_1_), .Y(mai_mai_n71_));
  NA2        m061(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n72_));
  NA2        m062(.A(mai_mai_n42_), .B(i_2_), .Y(mai_mai_n73_));
  NOi21      m063(.An(i_1_), .B(i_2_), .Y(mai_mai_n74_));
  NA3        m064(.A(mai_mai_n74_), .B(mai_mai_n53_), .C(i_6_), .Y(mai_mai_n75_));
  OAI210     m065(.A0(mai_mai_n73_), .A1(mai_mai_n72_), .B0(mai_mai_n75_), .Y(mai_mai_n76_));
  OAI210     m066(.A0(mai_mai_n76_), .A1(mai_mai_n71_), .B0(mai_mai_n14_), .Y(mai_mai_n77_));
  NA3        m067(.A(mai_mai_n65_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n78_));
  NA3        m068(.A(mai_mai_n26_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n79_));
  NA2        m069(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  NOi32      m070(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n81_));
  NA2        m071(.A(mai_mai_n81_), .B(i_3_), .Y(mai_mai_n82_));
  NA3        m072(.A(mai_mai_n18_), .B(i_2_), .C(i_6_), .Y(mai_mai_n83_));
  NA2        m073(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n84_));
  INV        m074(.A(i_0_), .Y(mai_mai_n85_));
  AOI220     m075(.A0(mai_mai_n85_), .A1(mai_mai_n84_), .B0(mai_mai_n80_), .B1(mai_mai_n61_), .Y(mai_mai_n86_));
  NA2        m076(.A(mai_mai_n86_), .B(mai_mai_n77_), .Y(mai_mai_n87_));
  NAi21      m077(.An(i_3_), .B(i_6_), .Y(mai_mai_n88_));
  NO3        m078(.A(mai_mai_n88_), .B(i_0_), .C(mai_mai_n50_), .Y(mai_mai_n89_));
  NA2        m079(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n90_));
  NOi21      m080(.An(i_7_), .B(i_8_), .Y(mai_mai_n91_));
  NOi31      m081(.An(i_6_), .B(i_5_), .C(i_7_), .Y(mai_mai_n92_));
  AOI210     m082(.A0(mai_mai_n91_), .A1(mai_mai_n12_), .B0(mai_mai_n92_), .Y(mai_mai_n93_));
  OAI210     m083(.A0(mai_mai_n93_), .A1(mai_mai_n11_), .B0(mai_mai_n90_), .Y(mai_mai_n94_));
  OAI210     m084(.A0(mai_mai_n94_), .A1(mai_mai_n89_), .B0(mai_mai_n74_), .Y(mai_mai_n95_));
  NA3        m085(.A(mai_mai_n25_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n96_));
  AOI210     m086(.A0(mai_mai_n22_), .A1(mai_mai_n51_), .B0(mai_mai_n96_), .Y(mai_mai_n97_));
  AOI220     m087(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n18_), .B1(mai_mai_n35_), .Y(mai_mai_n98_));
  NA3        m088(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n99_));
  NO2        m089(.A(mai_mai_n99_), .B(mai_mai_n98_), .Y(mai_mai_n100_));
  NO2        m090(.A(mai_mai_n100_), .B(mai_mai_n97_), .Y(mai_mai_n101_));
  NA3        m091(.A(mai_mai_n65_), .B(mai_mai_n35_), .C(i_3_), .Y(mai_mai_n102_));
  NA2        m092(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n103_));
  AOI210     m093(.A0(mai_mai_n103_), .A1(mai_mai_n22_), .B0(mai_mai_n102_), .Y(mai_mai_n104_));
  NAi21      m094(.An(i_6_), .B(i_0_), .Y(mai_mai_n105_));
  NA3        m095(.A(mai_mai_n62_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n106_));
  NOi21      m096(.An(i_4_), .B(i_6_), .Y(mai_mai_n107_));
  NOi21      m097(.An(i_5_), .B(i_3_), .Y(mai_mai_n108_));
  NA3        m098(.A(mai_mai_n108_), .B(mai_mai_n74_), .C(mai_mai_n107_), .Y(mai_mai_n109_));
  OAI210     m099(.A0(mai_mai_n106_), .A1(mai_mai_n105_), .B0(mai_mai_n109_), .Y(mai_mai_n110_));
  NA2        m100(.A(mai_mai_n74_), .B(mai_mai_n37_), .Y(mai_mai_n111_));
  NOi21      m101(.An(mai_mai_n43_), .B(mai_mai_n111_), .Y(mai_mai_n112_));
  NO3        m102(.A(mai_mai_n112_), .B(mai_mai_n110_), .C(mai_mai_n104_), .Y(mai_mai_n113_));
  NOi21      m103(.An(i_6_), .B(i_1_), .Y(mai_mai_n114_));
  AOI220     m104(.A0(mai_mai_n114_), .A1(i_7_), .B0(mai_mai_n25_), .B1(i_5_), .Y(mai_mai_n115_));
  NOi31      m105(.An(mai_mai_n53_), .B(mai_mai_n115_), .C(i_2_), .Y(mai_mai_n116_));
  NA2        m106(.A(mai_mai_n65_), .B(mai_mai_n12_), .Y(mai_mai_n117_));
  NA2        m107(.A(mai_mai_n37_), .B(mai_mai_n14_), .Y(mai_mai_n118_));
  NOi21      m108(.An(i_3_), .B(i_1_), .Y(mai_mai_n119_));
  NA2        m109(.A(mai_mai_n119_), .B(i_4_), .Y(mai_mai_n120_));
  AOI210     m110(.A0(mai_mai_n118_), .A1(mai_mai_n117_), .B0(mai_mai_n120_), .Y(mai_mai_n121_));
  NOi31      m111(.An(mai_mai_n46_), .B(i_5_), .C(mai_mai_n35_), .Y(mai_mai_n122_));
  NO3        m112(.A(mai_mai_n122_), .B(mai_mai_n121_), .C(mai_mai_n116_), .Y(mai_mai_n123_));
  NA4        m113(.A(mai_mai_n123_), .B(mai_mai_n113_), .C(mai_mai_n101_), .D(mai_mai_n95_), .Y(mai_mai_n124_));
  NA2        m114(.A(mai_mai_n56_), .B(mai_mai_n15_), .Y(mai_mai_n125_));
  NOi31      m115(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n126_));
  NOi31      m116(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n127_));
  OAI210     m117(.A0(mai_mai_n127_), .A1(mai_mai_n126_), .B0(i_7_), .Y(mai_mai_n128_));
  NA3        m118(.A(mai_mai_n37_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n129_));
  NA4        m119(.A(mai_mai_n129_), .B(mai_mai_n128_), .C(mai_mai_n125_), .D(mai_mai_n111_), .Y(mai_mai_n130_));
  NA2        m120(.A(mai_mai_n130_), .B(mai_mai_n41_), .Y(mai_mai_n131_));
  NO2        m121(.A(mai_mai_n78_), .B(mai_mai_n31_), .Y(mai_mai_n132_));
  NA4        m122(.A(mai_mai_n63_), .B(i_2_), .C(mai_mai_n17_), .D(mai_mai_n12_), .Y(mai_mai_n133_));
  NA3        m123(.A(mai_mai_n65_), .B(mai_mai_n60_), .C(i_6_), .Y(mai_mai_n134_));
  NA2        m124(.A(mai_mai_n134_), .B(mai_mai_n133_), .Y(mai_mai_n135_));
  NOi21      m125(.An(i_0_), .B(i_2_), .Y(mai_mai_n136_));
  NOi32      m126(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(mai_mai_n137_));
  NA2        m127(.A(mai_mai_n137_), .B(mai_mai_n126_), .Y(mai_mai_n138_));
  NA3        m128(.A(mai_mai_n136_), .B(mai_mai_n61_), .C(mai_mai_n37_), .Y(mai_mai_n139_));
  NA2        m129(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n140_));
  NA4        m130(.A(mai_mai_n60_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n141_));
  NA4        m131(.A(mai_mai_n62_), .B(mai_mai_n38_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n142_));
  NA4        m132(.A(mai_mai_n62_), .B(mai_mai_n46_), .C(i_5_), .D(mai_mai_n23_), .Y(mai_mai_n143_));
  NA3        m133(.A(mai_mai_n143_), .B(mai_mai_n142_), .C(mai_mai_n141_), .Y(mai_mai_n144_));
  NO4        m134(.A(mai_mai_n144_), .B(mai_mai_n140_), .C(mai_mai_n135_), .D(mai_mai_n132_), .Y(mai_mai_n145_));
  NOi21      m135(.An(i_5_), .B(i_2_), .Y(mai_mai_n146_));
  AOI220     m136(.A0(mai_mai_n146_), .A1(mai_mai_n91_), .B0(mai_mai_n63_), .B1(mai_mai_n32_), .Y(mai_mai_n147_));
  AOI210     m137(.A0(mai_mai_n147_), .A1(mai_mai_n125_), .B0(mai_mai_n103_), .Y(mai_mai_n148_));
  NO4        m138(.A(i_2_), .B(mai_mai_n21_), .C(mai_mai_n11_), .D(mai_mai_n14_), .Y(mai_mai_n149_));
  NA2        m139(.A(i_2_), .B(i_4_), .Y(mai_mai_n150_));
  AOI210     m140(.A0(mai_mai_n105_), .A1(mai_mai_n88_), .B0(mai_mai_n150_), .Y(mai_mai_n151_));
  NO2        m141(.A(i_8_), .B(i_7_), .Y(mai_mai_n152_));
  OA210      m142(.A0(mai_mai_n151_), .A1(mai_mai_n149_), .B0(mai_mai_n152_), .Y(mai_mai_n153_));
  NA3        m143(.A(mai_mai_n119_), .B(i_0_), .C(mai_mai_n23_), .Y(mai_mai_n154_));
  NO2        m144(.A(mai_mai_n154_), .B(i_4_), .Y(mai_mai_n155_));
  NO3        m145(.A(mai_mai_n155_), .B(mai_mai_n153_), .C(mai_mai_n148_), .Y(mai_mai_n156_));
  NA2        m146(.A(mai_mai_n91_), .B(mai_mai_n12_), .Y(mai_mai_n157_));
  NA3        m147(.A(i_2_), .B(i_1_), .C(mai_mai_n14_), .Y(mai_mai_n158_));
  INV        m148(.A(mai_mai_n53_), .Y(mai_mai_n159_));
  AOI210     m149(.A0(mai_mai_n159_), .A1(mai_mai_n158_), .B0(mai_mai_n157_), .Y(mai_mai_n160_));
  NA3        m150(.A(mai_mai_n136_), .B(mai_mai_n65_), .C(mai_mai_n107_), .Y(mai_mai_n161_));
  OAI210     m151(.A0(mai_mai_n102_), .A1(mai_mai_n31_), .B0(mai_mai_n161_), .Y(mai_mai_n162_));
  NA3        m152(.A(mai_mai_n108_), .B(mai_mai_n63_), .C(mai_mai_n45_), .Y(mai_mai_n163_));
  NOi31      m153(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n164_));
  OAI210     m154(.A0(mai_mai_n137_), .A1(mai_mai_n81_), .B0(mai_mai_n164_), .Y(mai_mai_n165_));
  NA2        m155(.A(mai_mai_n165_), .B(mai_mai_n163_), .Y(mai_mai_n166_));
  NO3        m156(.A(mai_mai_n166_), .B(mai_mai_n162_), .C(mai_mai_n160_), .Y(mai_mai_n167_));
  NA4        m157(.A(mai_mai_n167_), .B(mai_mai_n156_), .C(mai_mai_n145_), .D(mai_mai_n131_), .Y(mai_mai_n168_));
  OR4        m158(.A(mai_mai_n168_), .B(mai_mai_n124_), .C(mai_mai_n87_), .D(mai_mai_n69_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  INV        u002(.A(i_5_), .Y(men_men_n13_));
  NOi21      u003(.An(i_3_), .B(i_7_), .Y(men_men_n14_));
  INV        u004(.A(i_0_), .Y(men_men_n15_));
  NOi21      u005(.An(i_1_), .B(i_3_), .Y(men_men_n16_));
  INV        u006(.A(i_4_), .Y(men_men_n17_));
  NA2        u007(.A(i_0_), .B(men_men_n17_), .Y(men_men_n18_));
  INV        u008(.A(i_7_), .Y(men_men_n19_));
  NA3        u009(.A(i_6_), .B(i_5_), .C(men_men_n19_), .Y(men_men_n20_));
  NOi21      u010(.An(i_8_), .B(i_6_), .Y(men_men_n21_));
  NOi21      u011(.An(i_1_), .B(i_8_), .Y(men_men_n22_));
  AOI220     u012(.A0(men_men_n22_), .A1(i_2_), .B0(men_men_n21_), .B1(i_5_), .Y(men_men_n23_));
  AOI210     u013(.A0(men_men_n23_), .A1(men_men_n20_), .B0(men_men_n18_), .Y(men_men_n24_));
  NA2        u014(.A(men_men_n24_), .B(men_men_n11_), .Y(men_men_n25_));
  NA2        u015(.A(i_0_), .B(men_men_n13_), .Y(men_men_n26_));
  NA2        u016(.A(men_men_n15_), .B(i_5_), .Y(men_men_n27_));
  NO2        u017(.A(i_2_), .B(i_4_), .Y(men_men_n28_));
  NA3        u018(.A(men_men_n28_), .B(i_6_), .C(i_8_), .Y(men_men_n29_));
  AOI210     u019(.A0(men_men_n27_), .A1(men_men_n26_), .B0(men_men_n29_), .Y(men_men_n30_));
  INV        u020(.A(i_2_), .Y(men_men_n31_));
  NOi21      u021(.An(i_5_), .B(i_0_), .Y(men_men_n32_));
  NOi21      u022(.An(i_6_), .B(i_8_), .Y(men_men_n33_));
  NOi21      u023(.An(i_7_), .B(i_1_), .Y(men_men_n34_));
  NOi21      u024(.An(i_5_), .B(i_6_), .Y(men_men_n35_));
  AOI220     u025(.A0(men_men_n35_), .A1(men_men_n34_), .B0(men_men_n33_), .B1(men_men_n32_), .Y(men_men_n36_));
  NO3        u026(.A(men_men_n36_), .B(men_men_n31_), .C(i_4_), .Y(men_men_n37_));
  NOi21      u027(.An(i_0_), .B(i_4_), .Y(men_men_n38_));
  XO2        u028(.A(i_1_), .B(i_3_), .Y(men_men_n39_));
  NOi21      u029(.An(i_7_), .B(i_5_), .Y(men_men_n40_));
  AN3        u030(.A(men_men_n40_), .B(men_men_n39_), .C(men_men_n38_), .Y(men_men_n41_));
  INV        u031(.A(i_1_), .Y(men_men_n42_));
  NOi21      u032(.An(i_3_), .B(i_0_), .Y(men_men_n43_));
  NA2        u033(.A(men_men_n43_), .B(men_men_n42_), .Y(men_men_n44_));
  NA3        u034(.A(i_6_), .B(men_men_n13_), .C(i_7_), .Y(men_men_n45_));
  AOI210     u035(.A0(men_men_n45_), .A1(men_men_n20_), .B0(men_men_n44_), .Y(men_men_n46_));
  NO4        u036(.A(men_men_n46_), .B(men_men_n41_), .C(men_men_n37_), .D(men_men_n30_), .Y(men_men_n47_));
  INV        u037(.A(i_8_), .Y(men_men_n48_));
  NA2        u038(.A(i_1_), .B(men_men_n11_), .Y(men_men_n49_));
  NO4        u039(.A(men_men_n49_), .B(men_men_n26_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n50_));
  NOi21      u040(.An(i_4_), .B(i_0_), .Y(men_men_n51_));
  AOI210     u041(.A0(men_men_n51_), .A1(men_men_n21_), .B0(men_men_n14_), .Y(men_men_n52_));
  NA2        u042(.A(i_1_), .B(men_men_n13_), .Y(men_men_n53_));
  NOi21      u043(.An(i_2_), .B(i_8_), .Y(men_men_n54_));
  NO2        u044(.A(men_men_n53_), .B(men_men_n52_), .Y(men_men_n55_));
  NO2        u045(.A(men_men_n55_), .B(men_men_n50_), .Y(men_men_n56_));
  NOi31      u046(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n57_));
  NA2        u047(.A(men_men_n57_), .B(i_0_), .Y(men_men_n58_));
  NOi21      u048(.An(i_4_), .B(i_3_), .Y(men_men_n59_));
  NOi21      u049(.An(i_1_), .B(i_4_), .Y(men_men_n60_));
  OAI210     u050(.A0(men_men_n60_), .A1(men_men_n59_), .B0(men_men_n54_), .Y(men_men_n61_));
  NA2        u051(.A(men_men_n61_), .B(men_men_n58_), .Y(men_men_n62_));
  AN2        u052(.A(i_8_), .B(i_7_), .Y(men_men_n63_));
  NA2        u053(.A(men_men_n63_), .B(men_men_n12_), .Y(men_men_n64_));
  NOi21      u054(.An(i_8_), .B(i_7_), .Y(men_men_n65_));
  NA3        u055(.A(men_men_n65_), .B(men_men_n59_), .C(i_6_), .Y(men_men_n66_));
  NA2        u056(.A(men_men_n64_), .B(men_men_n66_), .Y(men_men_n67_));
  AOI220     u057(.A0(men_men_n67_), .A1(men_men_n31_), .B0(men_men_n62_), .B1(men_men_n35_), .Y(men_men_n68_));
  NA4        u058(.A(men_men_n68_), .B(men_men_n56_), .C(men_men_n47_), .D(men_men_n25_), .Y(men_men_n69_));
  NA2        u059(.A(i_8_), .B(i_7_), .Y(men_men_n70_));
  NA2        u060(.A(i_8_), .B(men_men_n19_), .Y(men_men_n71_));
  NA2        u061(.A(men_men_n39_), .B(i_2_), .Y(men_men_n72_));
  NOi21      u062(.An(i_1_), .B(i_2_), .Y(men_men_n73_));
  NA3        u063(.A(men_men_n73_), .B(men_men_n51_), .C(i_6_), .Y(men_men_n74_));
  OAI210     u064(.A0(men_men_n72_), .A1(men_men_n71_), .B0(men_men_n74_), .Y(men_men_n75_));
  NA2        u065(.A(men_men_n75_), .B(men_men_n13_), .Y(men_men_n76_));
  NA3        u066(.A(men_men_n65_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n77_));
  NA3        u067(.A(men_men_n22_), .B(i_0_), .C(men_men_n13_), .Y(men_men_n78_));
  NA2        u068(.A(men_men_n78_), .B(men_men_n77_), .Y(men_men_n79_));
  NOi32      u069(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n80_));
  NA2        u070(.A(men_men_n80_), .B(i_3_), .Y(men_men_n81_));
  NA3        u071(.A(men_men_n16_), .B(i_2_), .C(i_6_), .Y(men_men_n82_));
  NA2        u072(.A(men_men_n82_), .B(men_men_n81_), .Y(men_men_n83_));
  NO2        u073(.A(i_0_), .B(i_4_), .Y(men_men_n84_));
  AOI220     u074(.A0(men_men_n84_), .A1(men_men_n83_), .B0(men_men_n79_), .B1(men_men_n59_), .Y(men_men_n85_));
  NA2        u075(.A(men_men_n85_), .B(men_men_n76_), .Y(men_men_n86_));
  NAi21      u076(.An(i_3_), .B(i_6_), .Y(men_men_n87_));
  NO3        u077(.A(men_men_n87_), .B(i_0_), .C(men_men_n48_), .Y(men_men_n88_));
  NA2        u078(.A(men_men_n33_), .B(men_men_n32_), .Y(men_men_n89_));
  NOi21      u079(.An(i_7_), .B(i_8_), .Y(men_men_n90_));
  OAI210     u080(.A0(i_6_), .A1(men_men_n11_), .B0(men_men_n89_), .Y(men_men_n91_));
  OAI210     u081(.A0(men_men_n91_), .A1(men_men_n88_), .B0(men_men_n73_), .Y(men_men_n92_));
  NA3        u082(.A(men_men_n21_), .B(i_2_), .C(men_men_n13_), .Y(men_men_n93_));
  AOI210     u083(.A0(men_men_n18_), .A1(men_men_n49_), .B0(men_men_n93_), .Y(men_men_n94_));
  AOI220     u084(.A0(men_men_n43_), .A1(men_men_n42_), .B0(men_men_n16_), .B1(men_men_n31_), .Y(men_men_n95_));
  NA3        u085(.A(men_men_n17_), .B(i_5_), .C(i_7_), .Y(men_men_n96_));
  NA2        u086(.A(i_4_), .B(i_5_), .Y(men_men_n97_));
  NA3        u087(.A(men_men_n70_), .B(men_men_n16_), .C(men_men_n15_), .Y(men_men_n98_));
  OAI220     u088(.A0(men_men_n98_), .A1(men_men_n97_), .B0(men_men_n96_), .B1(men_men_n95_), .Y(men_men_n99_));
  NO2        u089(.A(men_men_n99_), .B(men_men_n94_), .Y(men_men_n100_));
  NA3        u090(.A(men_men_n65_), .B(men_men_n31_), .C(i_3_), .Y(men_men_n101_));
  NA2        u091(.A(men_men_n42_), .B(i_6_), .Y(men_men_n102_));
  AOI210     u092(.A0(men_men_n102_), .A1(men_men_n18_), .B0(men_men_n101_), .Y(men_men_n103_));
  NAi21      u093(.An(i_6_), .B(i_0_), .Y(men_men_n104_));
  NA3        u094(.A(men_men_n60_), .B(i_5_), .C(men_men_n19_), .Y(men_men_n105_));
  NOi21      u095(.An(i_4_), .B(i_6_), .Y(men_men_n106_));
  NOi21      u096(.An(i_5_), .B(i_3_), .Y(men_men_n107_));
  NA3        u097(.A(men_men_n107_), .B(men_men_n73_), .C(men_men_n106_), .Y(men_men_n108_));
  OAI210     u098(.A0(men_men_n105_), .A1(men_men_n104_), .B0(men_men_n108_), .Y(men_men_n109_));
  NA2        u099(.A(men_men_n73_), .B(men_men_n33_), .Y(men_men_n110_));
  NOi21      u100(.An(men_men_n40_), .B(men_men_n110_), .Y(men_men_n111_));
  NO3        u101(.A(men_men_n111_), .B(men_men_n109_), .C(men_men_n103_), .Y(men_men_n112_));
  NOi21      u102(.An(i_6_), .B(i_1_), .Y(men_men_n113_));
  AOI220     u103(.A0(men_men_n113_), .A1(i_7_), .B0(men_men_n21_), .B1(i_5_), .Y(men_men_n114_));
  NOi31      u104(.An(men_men_n51_), .B(men_men_n114_), .C(i_2_), .Y(men_men_n115_));
  NOi21      u105(.An(i_3_), .B(i_1_), .Y(men_men_n116_));
  NA2        u106(.A(men_men_n116_), .B(i_4_), .Y(men_men_n117_));
  AOI210     u107(.A0(i_8_), .A1(i_6_), .B0(men_men_n117_), .Y(men_men_n118_));
  NA2        u108(.A(men_men_n90_), .B(men_men_n13_), .Y(men_men_n119_));
  NOi31      u109(.An(men_men_n43_), .B(men_men_n119_), .C(men_men_n31_), .Y(men_men_n120_));
  NO3        u110(.A(men_men_n120_), .B(men_men_n118_), .C(men_men_n115_), .Y(men_men_n121_));
  NA4        u111(.A(men_men_n121_), .B(men_men_n112_), .C(men_men_n100_), .D(men_men_n92_), .Y(men_men_n122_));
  NA2        u112(.A(men_men_n54_), .B(men_men_n14_), .Y(men_men_n123_));
  NOi31      u113(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n124_));
  NA2        u114(.A(men_men_n124_), .B(i_7_), .Y(men_men_n125_));
  NA2        u115(.A(men_men_n33_), .B(men_men_n13_), .Y(men_men_n126_));
  NA4        u116(.A(men_men_n126_), .B(men_men_n125_), .C(men_men_n123_), .D(men_men_n110_), .Y(men_men_n127_));
  NA2        u117(.A(men_men_n127_), .B(men_men_n38_), .Y(men_men_n128_));
  NA2        u118(.A(men_men_n59_), .B(men_men_n34_), .Y(men_men_n129_));
  AOI210     u119(.A0(men_men_n129_), .A1(men_men_n77_), .B0(men_men_n27_), .Y(men_men_n130_));
  NA3        u120(.A(men_men_n65_), .B(men_men_n57_), .C(i_6_), .Y(men_men_n131_));
  INV        u121(.A(men_men_n131_), .Y(men_men_n132_));
  NA3        u122(.A(men_men_n51_), .B(men_men_n40_), .C(men_men_n16_), .Y(men_men_n133_));
  NA2        u123(.A(men_men_n59_), .B(men_men_n33_), .Y(men_men_n134_));
  NA2        u124(.A(men_men_n134_), .B(men_men_n133_), .Y(men_men_n135_));
  NA3        u125(.A(men_men_n57_), .B(men_men_n13_), .C(i_7_), .Y(men_men_n136_));
  NA4        u126(.A(men_men_n60_), .B(men_men_n35_), .C(men_men_n15_), .D(i_8_), .Y(men_men_n137_));
  NA4        u127(.A(men_men_n60_), .B(men_men_n43_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n138_));
  NA3        u128(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n139_));
  NO4        u129(.A(men_men_n139_), .B(men_men_n135_), .C(men_men_n132_), .D(men_men_n130_), .Y(men_men_n140_));
  BUFFER     u130(.A(i_5_), .Y(men_men_n141_));
  AOI220     u131(.A0(men_men_n141_), .A1(men_men_n90_), .B0(men_men_n63_), .B1(men_men_n28_), .Y(men_men_n142_));
  AOI210     u132(.A0(men_men_n142_), .A1(men_men_n123_), .B0(men_men_n102_), .Y(men_men_n143_));
  NA2        u133(.A(i_2_), .B(i_4_), .Y(men_men_n144_));
  NO2        u134(.A(men_men_n104_), .B(men_men_n144_), .Y(men_men_n145_));
  NO2        u135(.A(i_8_), .B(i_7_), .Y(men_men_n146_));
  AN2        u136(.A(men_men_n145_), .B(men_men_n146_), .Y(men_men_n147_));
  NA4        u137(.A(men_men_n116_), .B(i_0_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n148_));
  NO2        u138(.A(men_men_n148_), .B(i_4_), .Y(men_men_n149_));
  NO3        u139(.A(men_men_n149_), .B(men_men_n147_), .C(men_men_n143_), .Y(men_men_n150_));
  NA2        u140(.A(men_men_n90_), .B(men_men_n12_), .Y(men_men_n151_));
  NA2        u141(.A(i_2_), .B(men_men_n13_), .Y(men_men_n152_));
  NA2        u142(.A(men_men_n51_), .B(i_3_), .Y(men_men_n153_));
  AOI210     u143(.A0(men_men_n153_), .A1(men_men_n152_), .B0(men_men_n151_), .Y(men_men_n154_));
  NO2        u144(.A(men_men_n101_), .B(men_men_n27_), .Y(men_men_n155_));
  NA4        u145(.A(men_men_n107_), .B(men_men_n63_), .C(men_men_n42_), .D(men_men_n17_), .Y(men_men_n156_));
  NA3        u146(.A(men_men_n54_), .B(men_men_n32_), .C(men_men_n14_), .Y(men_men_n157_));
  NOi31      u147(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n158_));
  NA2        u148(.A(i_4_), .B(men_men_n158_), .Y(men_men_n159_));
  NA3        u149(.A(men_men_n159_), .B(men_men_n157_), .C(men_men_n156_), .Y(men_men_n160_));
  NO3        u150(.A(men_men_n160_), .B(men_men_n155_), .C(men_men_n154_), .Y(men_men_n161_));
  NA4        u151(.A(men_men_n161_), .B(men_men_n150_), .C(men_men_n140_), .D(men_men_n128_), .Y(men_men_n162_));
  OR4        u152(.A(men_men_n162_), .B(men_men_n122_), .C(men_men_n86_), .D(men_men_n69_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule