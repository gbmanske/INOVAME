library verilog;
use verilog.vl_types.all;
entity ContDe1_1always_vlg_vec_tst is
end ContDe1_1always_vlg_vec_tst;
