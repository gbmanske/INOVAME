//Benchmark atmr_max1024_476_0.0625

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n448_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(x8), .B(x7), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n61_));
  INV        o045(.A(x9), .Y(ori_ori_n62_));
  NO2        o046(.A(x7), .B(x6), .Y(ori_ori_n63_));
  NO2        o047(.A(ori_ori_n61_), .B(x5), .Y(ori_ori_n64_));
  NO2        o048(.A(x8), .B(x2), .Y(ori_ori_n65_));
  INV        o049(.A(ori_ori_n65_), .Y(ori_ori_n66_));
  NO2        o050(.A(ori_ori_n66_), .B(x1), .Y(ori_ori_n67_));
  AN2        o051(.A(ori_ori_n67_), .B(ori_ori_n63_), .Y(ori_ori_n68_));
  OAI210     o052(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n69_), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n70_), .B(ori_ori_n68_), .Y(ori_ori_n71_));
  NA2        o055(.A(ori_ori_n71_), .B(x4), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n73_));
  OAI210     o057(.A0(ori_ori_n73_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n74_));
  NA2        o058(.A(x5), .B(x3), .Y(ori_ori_n75_));
  NO2        o059(.A(x8), .B(x6), .Y(ori_ori_n76_));
  NO4        o060(.A(ori_ori_n76_), .B(ori_ori_n75_), .C(ori_ori_n63_), .D(ori_ori_n54_), .Y(ori_ori_n77_));
  NAi21      o061(.An(x4), .B(x3), .Y(ori_ori_n78_));
  INV        o062(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NO2        o063(.A(ori_ori_n79_), .B(ori_ori_n22_), .Y(ori_ori_n80_));
  NO2        o064(.A(x4), .B(x2), .Y(ori_ori_n81_));
  NO2        o065(.A(ori_ori_n81_), .B(x3), .Y(ori_ori_n82_));
  NO3        o066(.A(ori_ori_n82_), .B(ori_ori_n80_), .C(ori_ori_n18_), .Y(ori_ori_n83_));
  NO3        o067(.A(ori_ori_n83_), .B(ori_ori_n77_), .C(ori_ori_n74_), .Y(ori_ori_n84_));
  NA2        o068(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n85_));
  NO2        o069(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n86_));
  INV        o070(.A(x8), .Y(ori_ori_n87_));
  NA2        o071(.A(x2), .B(x1), .Y(ori_ori_n88_));
  INV        o072(.A(ori_ori_n86_), .Y(ori_ori_n89_));
  NO2        o073(.A(ori_ori_n89_), .B(ori_ori_n26_), .Y(ori_ori_n90_));
  AOI210     o074(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n91_));
  OAI210     o075(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n92_));
  NO3        o076(.A(ori_ori_n92_), .B(ori_ori_n91_), .C(ori_ori_n90_), .Y(ori_ori_n93_));
  NA2        o077(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n94_));
  NO2        o078(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n95_));
  OAI210     o079(.A0(ori_ori_n95_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n96_));
  AOI210     o080(.A0(ori_ori_n94_), .A1(ori_ori_n52_), .B0(ori_ori_n96_), .Y(ori_ori_n97_));
  NO2        o081(.A(x3), .B(x2), .Y(ori_ori_n98_));
  NA3        o082(.A(ori_ori_n98_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n99_));
  INV        o083(.A(ori_ori_n99_), .Y(ori_ori_n100_));
  NA2        o084(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n101_));
  OAI210     o085(.A0(ori_ori_n101_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n102_));
  NO4        o086(.A(ori_ori_n102_), .B(ori_ori_n100_), .C(ori_ori_n97_), .D(ori_ori_n93_), .Y(ori_ori_n103_));
  AO210      o087(.A0(ori_ori_n84_), .A1(ori_ori_n72_), .B0(ori_ori_n103_), .Y(ori02));
  NO2        o088(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n105_));
  NO2        o089(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n106_));
  NA2        o090(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n107_));
  NAi21      o091(.An(x2), .B(x8), .Y(ori_ori_n108_));
  NO2        o092(.A(x4), .B(x1), .Y(ori_ori_n109_));
  NA2        o093(.A(ori_ori_n109_), .B(x2), .Y(ori_ori_n110_));
  NOi21      o094(.An(x0), .B(x1), .Y(ori_ori_n111_));
  NO3        o095(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n112_));
  NOi21      o096(.An(x0), .B(x4), .Y(ori_ori_n113_));
  AOI220     o097(.A0(x7), .A1(ori_ori_n113_), .B0(ori_ori_n112_), .B1(ori_ori_n111_), .Y(ori_ori_n114_));
  AOI210     o098(.A0(ori_ori_n114_), .A1(ori_ori_n110_), .B0(ori_ori_n75_), .Y(ori_ori_n115_));
  NO2        o099(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n116_));
  NA2        o100(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n117_));
  AOI210     o101(.A0(ori_ori_n117_), .A1(ori_ori_n101_), .B0(ori_ori_n107_), .Y(ori_ori_n118_));
  OAI210     o102(.A0(ori_ori_n118_), .A1(ori_ori_n35_), .B0(ori_ori_n116_), .Y(ori_ori_n119_));
  NAi21      o103(.An(x0), .B(x4), .Y(ori_ori_n120_));
  NO2        o104(.A(ori_ori_n120_), .B(x1), .Y(ori_ori_n121_));
  NO2        o105(.A(x7), .B(x0), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n81_), .B(ori_ori_n95_), .Y(ori_ori_n123_));
  NO2        o107(.A(ori_ori_n123_), .B(x3), .Y(ori_ori_n124_));
  OAI210     o108(.A0(ori_ori_n122_), .A1(ori_ori_n121_), .B0(ori_ori_n124_), .Y(ori_ori_n125_));
  NO2        o109(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n126_));
  NA2        o110(.A(x5), .B(x0), .Y(ori_ori_n127_));
  NO2        o111(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n128_));
  NA3        o112(.A(ori_ori_n128_), .B(ori_ori_n127_), .C(ori_ori_n126_), .Y(ori_ori_n129_));
  NA4        o113(.A(ori_ori_n129_), .B(ori_ori_n125_), .C(ori_ori_n119_), .D(ori_ori_n36_), .Y(ori_ori_n130_));
  NO2        o114(.A(ori_ori_n130_), .B(ori_ori_n115_), .Y(ori_ori_n131_));
  NO3        o115(.A(ori_ori_n75_), .B(ori_ori_n73_), .C(ori_ori_n24_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n133_));
  NA2        o117(.A(x7), .B(x3), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n94_), .B(x5), .Y(ori_ori_n135_));
  NO2        o119(.A(x9), .B(x7), .Y(ori_ori_n136_));
  NOi21      o120(.An(x8), .B(x0), .Y(ori_ori_n137_));
  NO2        o121(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n138_));
  INV        o122(.A(x7), .Y(ori_ori_n139_));
  NA2        o123(.A(ori_ori_n139_), .B(ori_ori_n18_), .Y(ori_ori_n140_));
  AOI220     o124(.A0(ori_ori_n140_), .A1(ori_ori_n138_), .B0(ori_ori_n105_), .B1(ori_ori_n38_), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n142_));
  NO2        o126(.A(ori_ori_n142_), .B(ori_ori_n113_), .Y(ori_ori_n143_));
  NO2        o127(.A(ori_ori_n143_), .B(ori_ori_n141_), .Y(ori_ori_n144_));
  INV        o128(.A(ori_ori_n144_), .Y(ori_ori_n145_));
  OAI210     o129(.A0(ori_ori_n134_), .A1(ori_ori_n50_), .B0(ori_ori_n145_), .Y(ori_ori_n146_));
  NA2        o130(.A(x5), .B(x1), .Y(ori_ori_n147_));
  INV        o131(.A(ori_ori_n147_), .Y(ori_ori_n148_));
  AOI210     o132(.A0(ori_ori_n148_), .A1(ori_ori_n113_), .B0(ori_ori_n36_), .Y(ori_ori_n149_));
  NAi21      o133(.An(x2), .B(x7), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n150_), .B(ori_ori_n48_), .Y(ori_ori_n151_));
  NA2        o135(.A(ori_ori_n151_), .B(ori_ori_n64_), .Y(ori_ori_n152_));
  NAi31      o136(.An(ori_ori_n75_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n153_));
  NA3        o137(.A(ori_ori_n153_), .B(ori_ori_n152_), .C(ori_ori_n149_), .Y(ori_ori_n154_));
  NO3        o138(.A(ori_ori_n154_), .B(ori_ori_n146_), .C(ori_ori_n132_), .Y(ori_ori_n155_));
  NO2        o139(.A(ori_ori_n155_), .B(ori_ori_n131_), .Y(ori_ori_n156_));
  NO2        o140(.A(ori_ori_n127_), .B(ori_ori_n123_), .Y(ori_ori_n157_));
  NA2        o141(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n158_));
  NA2        o142(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n159_));
  NA3        o143(.A(ori_ori_n159_), .B(ori_ori_n158_), .C(ori_ori_n24_), .Y(ori_ori_n160_));
  AN2        o144(.A(ori_ori_n160_), .B(ori_ori_n128_), .Y(ori_ori_n161_));
  NA2        o145(.A(x8), .B(x0), .Y(ori_ori_n162_));
  NO2        o146(.A(ori_ori_n139_), .B(ori_ori_n25_), .Y(ori_ori_n163_));
  NA2        o147(.A(x2), .B(x0), .Y(ori_ori_n164_));
  NA2        o148(.A(x4), .B(x1), .Y(ori_ori_n165_));
  NAi21      o149(.An(ori_ori_n109_), .B(ori_ori_n165_), .Y(ori_ori_n166_));
  NOi31      o150(.An(ori_ori_n166_), .B(ori_ori_n142_), .C(ori_ori_n164_), .Y(ori_ori_n167_));
  NO3        o151(.A(ori_ori_n167_), .B(ori_ori_n161_), .C(ori_ori_n157_), .Y(ori_ori_n168_));
  NO2        o152(.A(ori_ori_n168_), .B(ori_ori_n43_), .Y(ori_ori_n169_));
  NO2        o153(.A(ori_ori_n160_), .B(ori_ori_n73_), .Y(ori_ori_n170_));
  INV        o154(.A(ori_ori_n116_), .Y(ori_ori_n171_));
  NO2        o155(.A(ori_ori_n101_), .B(ori_ori_n17_), .Y(ori_ori_n172_));
  AOI210     o156(.A0(ori_ori_n35_), .A1(ori_ori_n87_), .B0(ori_ori_n172_), .Y(ori_ori_n173_));
  NO3        o157(.A(ori_ori_n173_), .B(ori_ori_n171_), .C(x7), .Y(ori_ori_n174_));
  NA3        o158(.A(ori_ori_n166_), .B(ori_ori_n171_), .C(ori_ori_n42_), .Y(ori_ori_n175_));
  OAI210     o159(.A0(ori_ori_n159_), .A1(ori_ori_n123_), .B0(ori_ori_n175_), .Y(ori_ori_n176_));
  NO3        o160(.A(ori_ori_n176_), .B(ori_ori_n174_), .C(ori_ori_n170_), .Y(ori_ori_n177_));
  NO2        o161(.A(ori_ori_n177_), .B(x3), .Y(ori_ori_n178_));
  NO3        o162(.A(ori_ori_n178_), .B(ori_ori_n169_), .C(ori_ori_n156_), .Y(ori03));
  NO2        o163(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n180_));
  NO2        o164(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n181_));
  NO2        o165(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n182_));
  NO2        o166(.A(ori_ori_n75_), .B(x6), .Y(ori_ori_n183_));
  NA2        o167(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n184_));
  NO2        o168(.A(ori_ori_n184_), .B(x4), .Y(ori_ori_n185_));
  NO2        o169(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n186_));
  NA2        o170(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n187_));
  NO2        o171(.A(ori_ori_n187_), .B(ori_ori_n184_), .Y(ori_ori_n188_));
  NA2        o172(.A(x9), .B(ori_ori_n54_), .Y(ori_ori_n189_));
  NA2        o173(.A(ori_ori_n189_), .B(x4), .Y(ori_ori_n190_));
  NA2        o174(.A(ori_ori_n184_), .B(ori_ori_n78_), .Y(ori_ori_n191_));
  AOI210     o175(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n164_), .Y(ori_ori_n192_));
  AOI220     o176(.A0(ori_ori_n192_), .A1(ori_ori_n191_), .B0(ori_ori_n190_), .B1(ori_ori_n188_), .Y(ori_ori_n193_));
  NO3        o177(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n194_));
  NO2        o178(.A(x5), .B(x1), .Y(ori_ori_n195_));
  NO2        o179(.A(ori_ori_n187_), .B(ori_ori_n158_), .Y(ori_ori_n196_));
  NO3        o180(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n197_));
  NO2        o181(.A(ori_ori_n197_), .B(ori_ori_n196_), .Y(ori_ori_n198_));
  INV        o182(.A(ori_ori_n198_), .Y(ori_ori_n199_));
  AOI220     o183(.A0(ori_ori_n199_), .A1(ori_ori_n48_), .B0(ori_ori_n194_), .B1(ori_ori_n116_), .Y(ori_ori_n200_));
  NA2        o184(.A(ori_ori_n200_), .B(ori_ori_n193_), .Y(ori_ori_n201_));
  NO2        o185(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n202_));
  NA2        o186(.A(ori_ori_n202_), .B(ori_ori_n19_), .Y(ori_ori_n203_));
  NO2        o187(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n204_));
  NO2        o188(.A(ori_ori_n204_), .B(x6), .Y(ori_ori_n205_));
  NOi21      o189(.An(ori_ori_n81_), .B(ori_ori_n205_), .Y(ori_ori_n206_));
  NA2        o190(.A(ori_ori_n62_), .B(ori_ori_n87_), .Y(ori_ori_n207_));
  NA3        o191(.A(ori_ori_n207_), .B(ori_ori_n204_), .C(x6), .Y(ori_ori_n208_));
  AOI210     o192(.A0(ori_ori_n208_), .A1(ori_ori_n206_), .B0(ori_ori_n139_), .Y(ori_ori_n209_));
  AO210      o193(.A0(ori_ori_n209_), .A1(ori_ori_n203_), .B0(ori_ori_n163_), .Y(ori_ori_n210_));
  NA2        o194(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n211_));
  OAI210     o195(.A0(ori_ori_n211_), .A1(ori_ori_n25_), .B0(ori_ori_n159_), .Y(ori_ori_n212_));
  NO3        o196(.A(ori_ori_n165_), .B(ori_ori_n62_), .C(x6), .Y(ori_ori_n213_));
  AOI220     o197(.A0(ori_ori_n213_), .A1(ori_ori_n212_), .B0(ori_ori_n128_), .B1(ori_ori_n86_), .Y(ori_ori_n214_));
  NA2        o198(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n215_));
  NO2        o199(.A(ori_ori_n215_), .B(ori_ori_n75_), .Y(ori_ori_n216_));
  INV        o200(.A(x6), .Y(ori_ori_n217_));
  NO2        o201(.A(ori_ori_n147_), .B(ori_ori_n43_), .Y(ori_ori_n218_));
  OAI210     o202(.A0(ori_ori_n218_), .A1(ori_ori_n196_), .B0(ori_ori_n217_), .Y(ori_ori_n219_));
  NA2        o203(.A(ori_ori_n181_), .B(ori_ori_n121_), .Y(ori_ori_n220_));
  NA3        o204(.A(ori_ori_n187_), .B(ori_ori_n116_), .C(x6), .Y(ori_ori_n221_));
  OAI210     o205(.A0(ori_ori_n87_), .A1(ori_ori_n36_), .B0(ori_ori_n64_), .Y(ori_ori_n222_));
  NA4        o206(.A(ori_ori_n222_), .B(ori_ori_n221_), .C(ori_ori_n220_), .D(ori_ori_n219_), .Y(ori_ori_n223_));
  OAI210     o207(.A0(ori_ori_n223_), .A1(ori_ori_n216_), .B0(x2), .Y(ori_ori_n224_));
  NA3        o208(.A(ori_ori_n224_), .B(ori_ori_n214_), .C(ori_ori_n210_), .Y(ori_ori_n225_));
  AOI210     o209(.A0(ori_ori_n201_), .A1(x8), .B0(ori_ori_n225_), .Y(ori_ori_n226_));
  NO2        o210(.A(ori_ori_n87_), .B(x3), .Y(ori_ori_n227_));
  NA2        o211(.A(ori_ori_n227_), .B(ori_ori_n185_), .Y(ori_ori_n228_));
  NO3        o212(.A(ori_ori_n85_), .B(ori_ori_n76_), .C(ori_ori_n25_), .Y(ori_ori_n229_));
  AOI210     o213(.A0(ori_ori_n205_), .A1(ori_ori_n142_), .B0(ori_ori_n229_), .Y(ori_ori_n230_));
  AOI210     o214(.A0(ori_ori_n230_), .A1(ori_ori_n228_), .B0(x2), .Y(ori_ori_n231_));
  NO2        o215(.A(x4), .B(ori_ori_n54_), .Y(ori_ori_n232_));
  AOI220     o216(.A0(ori_ori_n185_), .A1(ori_ori_n172_), .B0(ori_ori_n232_), .B1(ori_ori_n64_), .Y(ori_ori_n233_));
  NA2        o217(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n234_));
  NA3        o218(.A(ori_ori_n25_), .B(x3), .C(x2), .Y(ori_ori_n235_));
  AOI210     o219(.A0(ori_ori_n235_), .A1(ori_ori_n127_), .B0(ori_ori_n234_), .Y(ori_ori_n236_));
  NA2        o220(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n237_));
  NO2        o221(.A(ori_ori_n237_), .B(ori_ori_n25_), .Y(ori_ori_n238_));
  OAI210     o222(.A0(ori_ori_n238_), .A1(ori_ori_n236_), .B0(ori_ori_n109_), .Y(ori_ori_n239_));
  NA2        o223(.A(ori_ori_n187_), .B(x6), .Y(ori_ori_n240_));
  NO2        o224(.A(ori_ori_n187_), .B(x6), .Y(ori_ori_n241_));
  INV        o225(.A(ori_ori_n241_), .Y(ori_ori_n242_));
  NA3        o226(.A(ori_ori_n242_), .B(ori_ori_n240_), .C(ori_ori_n133_), .Y(ori_ori_n243_));
  NA4        o227(.A(ori_ori_n243_), .B(ori_ori_n239_), .C(ori_ori_n233_), .D(ori_ori_n139_), .Y(ori_ori_n244_));
  NA2        o228(.A(ori_ori_n181_), .B(ori_ori_n204_), .Y(ori_ori_n245_));
  NO2        o229(.A(x9), .B(x6), .Y(ori_ori_n246_));
  NO2        o230(.A(ori_ori_n127_), .B(ori_ori_n18_), .Y(ori_ori_n247_));
  NAi21      o231(.An(ori_ori_n247_), .B(ori_ori_n235_), .Y(ori_ori_n248_));
  NAi21      o232(.An(x1), .B(x4), .Y(ori_ori_n249_));
  AOI210     o233(.A0(x3), .A1(x2), .B0(ori_ori_n48_), .Y(ori_ori_n250_));
  OAI210     o234(.A0(ori_ori_n127_), .A1(x3), .B0(ori_ori_n250_), .Y(ori_ori_n251_));
  AOI220     o235(.A0(ori_ori_n251_), .A1(ori_ori_n249_), .B0(ori_ori_n248_), .B1(ori_ori_n246_), .Y(ori_ori_n252_));
  NA2        o236(.A(ori_ori_n252_), .B(ori_ori_n245_), .Y(ori_ori_n253_));
  NA2        o237(.A(ori_ori_n62_), .B(x2), .Y(ori_ori_n254_));
  NO2        o238(.A(ori_ori_n254_), .B(ori_ori_n245_), .Y(ori_ori_n255_));
  NA2        o239(.A(x6), .B(x2), .Y(ori_ori_n256_));
  OAI210     o240(.A0(x4), .A1(ori_ori_n255_), .B0(ori_ori_n253_), .Y(ori_ori_n257_));
  NO2        o241(.A(x3), .B(ori_ori_n184_), .Y(ori_ori_n258_));
  OR2        o242(.A(ori_ori_n258_), .B(ori_ori_n183_), .Y(ori_ori_n259_));
  NA2        o243(.A(x4), .B(x0), .Y(ori_ori_n260_));
  NA2        o244(.A(ori_ori_n259_), .B(ori_ori_n42_), .Y(ori_ori_n261_));
  AOI210     o245(.A0(ori_ori_n261_), .A1(ori_ori_n257_), .B0(x8), .Y(ori_ori_n262_));
  INV        o246(.A(ori_ori_n234_), .Y(ori_ori_n263_));
  NA2        o247(.A(ori_ori_n247_), .B(ori_ori_n263_), .Y(ori_ori_n264_));
  INV        o248(.A(ori_ori_n162_), .Y(ori_ori_n265_));
  OAI210     o249(.A0(ori_ori_n265_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n266_));
  AOI210     o250(.A0(ori_ori_n266_), .A1(ori_ori_n264_), .B0(ori_ori_n211_), .Y(ori_ori_n267_));
  NO4        o251(.A(ori_ori_n267_), .B(ori_ori_n262_), .C(ori_ori_n244_), .D(ori_ori_n231_), .Y(ori_ori_n268_));
  INV        o252(.A(x1), .Y(ori_ori_n269_));
  OAI210     o253(.A0(x1), .A1(ori_ori_n241_), .B0(x2), .Y(ori_ori_n270_));
  OAI210     o254(.A0(ori_ori_n265_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n271_));
  AOI210     o255(.A0(ori_ori_n271_), .A1(ori_ori_n270_), .B0(ori_ori_n171_), .Y(ori_ori_n272_));
  NOi21      o256(.An(ori_ori_n256_), .B(ori_ori_n17_), .Y(ori_ori_n273_));
  NA3        o257(.A(ori_ori_n273_), .B(ori_ori_n195_), .C(ori_ori_n40_), .Y(ori_ori_n274_));
  AOI210     o258(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n275_));
  NA3        o259(.A(ori_ori_n275_), .B(ori_ori_n148_), .C(ori_ori_n32_), .Y(ori_ori_n276_));
  NA2        o260(.A(x3), .B(x2), .Y(ori_ori_n277_));
  AOI220     o261(.A0(ori_ori_n277_), .A1(ori_ori_n211_), .B0(ori_ori_n276_), .B1(ori_ori_n274_), .Y(ori_ori_n278_));
  NAi21      o262(.An(x4), .B(x0), .Y(ori_ori_n279_));
  NO3        o263(.A(ori_ori_n279_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n280_));
  OAI210     o264(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n280_), .Y(ori_ori_n281_));
  OAI220     o265(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n282_));
  NO2        o266(.A(x9), .B(x8), .Y(ori_ori_n283_));
  NA3        o267(.A(ori_ori_n283_), .B(ori_ori_n36_), .C(ori_ori_n54_), .Y(ori_ori_n284_));
  OAI210     o268(.A0(ori_ori_n275_), .A1(ori_ori_n273_), .B0(ori_ori_n284_), .Y(ori_ori_n285_));
  AOI220     o269(.A0(ori_ori_n285_), .A1(ori_ori_n79_), .B0(ori_ori_n282_), .B1(ori_ori_n31_), .Y(ori_ori_n286_));
  AOI210     o270(.A0(ori_ori_n286_), .A1(ori_ori_n281_), .B0(ori_ori_n25_), .Y(ori_ori_n287_));
  NO2        o271(.A(ori_ori_n275_), .B(ori_ori_n273_), .Y(ori_ori_n288_));
  INV        o272(.A(ori_ori_n196_), .Y(ori_ori_n289_));
  NA2        o273(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n290_));
  OR2        o274(.A(ori_ori_n290_), .B(ori_ori_n260_), .Y(ori_ori_n291_));
  OAI220     o275(.A0(ori_ori_n291_), .A1(ori_ori_n147_), .B0(ori_ori_n215_), .B1(ori_ori_n289_), .Y(ori_ori_n292_));
  AO210      o276(.A0(ori_ori_n288_), .A1(ori_ori_n135_), .B0(ori_ori_n292_), .Y(ori_ori_n293_));
  NO4        o277(.A(ori_ori_n293_), .B(ori_ori_n287_), .C(ori_ori_n278_), .D(ori_ori_n272_), .Y(ori_ori_n294_));
  OAI210     o278(.A0(ori_ori_n268_), .A1(ori_ori_n226_), .B0(ori_ori_n294_), .Y(ori04));
  NO2        o279(.A(x2), .B(x1), .Y(ori_ori_n296_));
  OAI210     o280(.A0(ori_ori_n237_), .A1(ori_ori_n296_), .B0(ori_ori_n36_), .Y(ori_ori_n297_));
  NO2        o281(.A(ori_ori_n296_), .B(ori_ori_n279_), .Y(ori_ori_n298_));
  OAI210     o282(.A0(ori_ori_n54_), .A1(ori_ori_n298_), .B0(ori_ori_n227_), .Y(ori_ori_n299_));
  NO2        o283(.A(ori_ori_n254_), .B(ori_ori_n85_), .Y(ori_ori_n300_));
  NO2        o284(.A(ori_ori_n300_), .B(ori_ori_n36_), .Y(ori_ori_n301_));
  NO2        o285(.A(ori_ori_n277_), .B(ori_ori_n186_), .Y(ori_ori_n302_));
  NA2        o286(.A(x9), .B(x0), .Y(ori_ori_n303_));
  AOI210     o287(.A0(ori_ori_n85_), .A1(ori_ori_n73_), .B0(ori_ori_n303_), .Y(ori_ori_n304_));
  OAI210     o288(.A0(ori_ori_n304_), .A1(ori_ori_n302_), .B0(ori_ori_n87_), .Y(ori_ori_n305_));
  NA3        o289(.A(ori_ori_n305_), .B(ori_ori_n301_), .C(ori_ori_n299_), .Y(ori_ori_n306_));
  NA2        o290(.A(ori_ori_n306_), .B(ori_ori_n297_), .Y(ori_ori_n307_));
  OAI210     o291(.A0(x0), .A1(ori_ori_n101_), .B0(ori_ori_n162_), .Y(ori_ori_n308_));
  NA3        o292(.A(ori_ori_n308_), .B(x6), .C(x3), .Y(ori_ori_n309_));
  AOI210     o293(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n310_));
  NO2        o294(.A(ori_ori_n310_), .B(ori_ori_n290_), .Y(ori_ori_n311_));
  INV        o295(.A(ori_ori_n311_), .Y(ori_ori_n312_));
  NA2        o296(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n313_));
  OAI210     o297(.A0(ori_ori_n101_), .A1(ori_ori_n17_), .B0(ori_ori_n313_), .Y(ori_ori_n314_));
  AOI220     o298(.A0(ori_ori_n314_), .A1(ori_ori_n76_), .B0(ori_ori_n300_), .B1(ori_ori_n87_), .Y(ori_ori_n315_));
  NA3        o299(.A(ori_ori_n315_), .B(ori_ori_n312_), .C(ori_ori_n309_), .Y(ori_ori_n316_));
  OAI210     o300(.A0(ori_ori_n106_), .A1(x3), .B0(ori_ori_n280_), .Y(ori_ori_n317_));
  NA2        o301(.A(ori_ori_n194_), .B(ori_ori_n81_), .Y(ori_ori_n318_));
  NA3        o302(.A(ori_ori_n318_), .B(ori_ori_n317_), .C(ori_ori_n139_), .Y(ori_ori_n319_));
  AOI210     o303(.A0(ori_ori_n316_), .A1(x4), .B0(ori_ori_n319_), .Y(ori_ori_n320_));
  NA3        o304(.A(ori_ori_n298_), .B(ori_ori_n189_), .C(ori_ori_n87_), .Y(ori_ori_n321_));
  NOi21      o305(.An(x4), .B(x0), .Y(ori_ori_n322_));
  XO2        o306(.A(x4), .B(x0), .Y(ori_ori_n323_));
  INV        o307(.A(ori_ori_n249_), .Y(ori_ori_n324_));
  AOI220     o308(.A0(ori_ori_n324_), .A1(x8), .B0(ori_ori_n322_), .B1(ori_ori_n88_), .Y(ori_ori_n325_));
  AOI210     o309(.A0(ori_ori_n325_), .A1(ori_ori_n321_), .B0(x3), .Y(ori_ori_n326_));
  INV        o310(.A(ori_ori_n88_), .Y(ori_ori_n327_));
  NO2        o311(.A(ori_ori_n87_), .B(x4), .Y(ori_ori_n328_));
  AOI220     o312(.A0(ori_ori_n328_), .A1(ori_ori_n44_), .B0(ori_ori_n113_), .B1(ori_ori_n327_), .Y(ori_ori_n329_));
  NO2        o313(.A(ori_ori_n323_), .B(x2), .Y(ori_ori_n330_));
  NO3        o314(.A(ori_ori_n207_), .B(ori_ori_n28_), .C(ori_ori_n24_), .Y(ori_ori_n331_));
  NO2        o315(.A(ori_ori_n331_), .B(ori_ori_n330_), .Y(ori_ori_n332_));
  NA4        o316(.A(ori_ori_n332_), .B(ori_ori_n329_), .C(ori_ori_n203_), .D(x6), .Y(ori_ori_n333_));
  NO2        o317(.A(ori_ori_n164_), .B(ori_ori_n87_), .Y(ori_ori_n334_));
  NO2        o318(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n335_));
  OR2        o319(.A(ori_ori_n328_), .B(ori_ori_n335_), .Y(ori_ori_n336_));
  NO2        o320(.A(ori_ori_n137_), .B(ori_ori_n101_), .Y(ori_ori_n337_));
  AOI220     o321(.A0(ori_ori_n337_), .A1(ori_ori_n336_), .B0(ori_ori_n334_), .B1(ori_ori_n61_), .Y(ori_ori_n338_));
  NO2        o322(.A(ori_ori_n137_), .B(ori_ori_n78_), .Y(ori_ori_n339_));
  NO2        o323(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n340_));
  NOi21      o324(.An(ori_ori_n109_), .B(ori_ori_n27_), .Y(ori_ori_n341_));
  AOI210     o325(.A0(ori_ori_n340_), .A1(ori_ori_n339_), .B0(ori_ori_n341_), .Y(ori_ori_n342_));
  OAI210     o326(.A0(ori_ori_n338_), .A1(ori_ori_n62_), .B0(ori_ori_n342_), .Y(ori_ori_n343_));
  OAI220     o327(.A0(ori_ori_n343_), .A1(x6), .B0(ori_ori_n333_), .B1(ori_ori_n326_), .Y(ori_ori_n344_));
  OAI210     o328(.A0(x6), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n345_));
  OAI210     o329(.A0(ori_ori_n345_), .A1(ori_ori_n87_), .B0(ori_ori_n291_), .Y(ori_ori_n346_));
  AOI210     o330(.A0(ori_ori_n346_), .A1(ori_ori_n18_), .B0(ori_ori_n139_), .Y(ori_ori_n347_));
  AO220      o331(.A0(ori_ori_n347_), .A1(ori_ori_n344_), .B0(ori_ori_n320_), .B1(ori_ori_n307_), .Y(ori_ori_n348_));
  NA2        o332(.A(ori_ori_n340_), .B(x6), .Y(ori_ori_n349_));
  AOI210     o333(.A0(x6), .A1(x1), .B0(ori_ori_n138_), .Y(ori_ori_n350_));
  NA2        o334(.A(ori_ori_n328_), .B(x0), .Y(ori_ori_n351_));
  NA2        o335(.A(ori_ori_n81_), .B(x6), .Y(ori_ori_n352_));
  OAI210     o336(.A0(ori_ori_n351_), .A1(ori_ori_n350_), .B0(ori_ori_n352_), .Y(ori_ori_n353_));
  AOI220     o337(.A0(ori_ori_n353_), .A1(ori_ori_n349_), .B0(ori_ori_n197_), .B1(ori_ori_n49_), .Y(ori_ori_n354_));
  NA2        o338(.A(ori_ori_n354_), .B(ori_ori_n348_), .Y(ori_ori_n355_));
  AOI210     o339(.A0(ori_ori_n182_), .A1(x8), .B0(ori_ori_n106_), .Y(ori_ori_n356_));
  NA2        o340(.A(ori_ori_n356_), .B(ori_ori_n313_), .Y(ori_ori_n357_));
  NA3        o341(.A(ori_ori_n357_), .B(ori_ori_n180_), .C(ori_ori_n139_), .Y(ori_ori_n358_));
  NA3        o342(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n359_));
  NA2        o343(.A(ori_ori_n202_), .B(x0), .Y(ori_ori_n360_));
  OAI220     o344(.A0(ori_ori_n360_), .A1(ori_ori_n189_), .B0(ori_ori_n359_), .B1(ori_ori_n327_), .Y(ori_ori_n361_));
  INV        o345(.A(ori_ori_n361_), .Y(ori_ori_n362_));
  AOI210     o346(.A0(ori_ori_n362_), .A1(ori_ori_n358_), .B0(ori_ori_n25_), .Y(ori_ori_n363_));
  OAI210     o347(.A0(ori_ori_n180_), .A1(ori_ori_n65_), .B0(ori_ori_n186_), .Y(ori_ori_n364_));
  NA3        o348(.A(ori_ori_n182_), .B(ori_ori_n204_), .C(x8), .Y(ori_ori_n365_));
  AOI210     o349(.A0(ori_ori_n365_), .A1(ori_ori_n364_), .B0(ori_ori_n25_), .Y(ori_ori_n366_));
  AOI210     o350(.A0(ori_ori_n108_), .A1(x0), .B0(ori_ori_n42_), .Y(ori_ori_n367_));
  NOi31      o351(.An(ori_ori_n367_), .B(ori_ori_n335_), .C(ori_ori_n165_), .Y(ori_ori_n368_));
  OAI210     o352(.A0(ori_ori_n368_), .A1(ori_ori_n366_), .B0(ori_ori_n136_), .Y(ori_ori_n369_));
  NAi31      o353(.An(ori_ori_n50_), .B(ori_ori_n269_), .C(ori_ori_n163_), .Y(ori_ori_n370_));
  NA2        o354(.A(ori_ori_n370_), .B(ori_ori_n369_), .Y(ori_ori_n371_));
  OAI210     o355(.A0(ori_ori_n371_), .A1(ori_ori_n363_), .B0(x6), .Y(ori_ori_n372_));
  NO2        o356(.A(x0), .B(ori_ori_n32_), .Y(ori_ori_n373_));
  NA2        o357(.A(ori_ori_n180_), .B(ori_ori_n139_), .Y(ori_ori_n374_));
  AOI210     o358(.A0(x7), .A1(ori_ori_n232_), .B0(x1), .Y(ori_ori_n375_));
  OAI210     o359(.A0(ori_ori_n374_), .A1(x8), .B0(ori_ori_n375_), .Y(ori_ori_n376_));
  NAi31      o360(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n377_));
  OAI210     o361(.A0(ori_ori_n377_), .A1(x4), .B0(ori_ori_n150_), .Y(ori_ori_n378_));
  NA3        o362(.A(ori_ori_n378_), .B(ori_ori_n134_), .C(x9), .Y(ori_ori_n379_));
  NO4        o363(.A(x8), .B(ori_ori_n279_), .C(x9), .D(x2), .Y(ori_ori_n380_));
  NOi21      o364(.An(ori_ori_n112_), .B(ori_ori_n164_), .Y(ori_ori_n381_));
  NO3        o365(.A(ori_ori_n381_), .B(ori_ori_n380_), .C(ori_ori_n18_), .Y(ori_ori_n382_));
  NA2        o366(.A(ori_ori_n339_), .B(ori_ori_n139_), .Y(ori_ori_n383_));
  NA4        o367(.A(ori_ori_n383_), .B(ori_ori_n382_), .C(ori_ori_n379_), .D(ori_ori_n50_), .Y(ori_ori_n384_));
  OAI210     o368(.A0(ori_ori_n376_), .A1(ori_ori_n373_), .B0(ori_ori_n384_), .Y(ori_ori_n385_));
  AOI210     o369(.A0(ori_ori_n38_), .A1(x9), .B0(ori_ori_n120_), .Y(ori_ori_n386_));
  NO3        o370(.A(ori_ori_n386_), .B(ori_ori_n112_), .C(ori_ori_n43_), .Y(ori_ori_n387_));
  NOi31      o371(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n388_));
  AOI220     o372(.A0(ori_ori_n388_), .A1(ori_ori_n322_), .B0(ori_ori_n113_), .B1(x3), .Y(ori_ori_n389_));
  AOI210     o373(.A0(ori_ori_n249_), .A1(ori_ori_n60_), .B0(ori_ori_n111_), .Y(ori_ori_n390_));
  OAI210     o374(.A0(ori_ori_n390_), .A1(x3), .B0(ori_ori_n389_), .Y(ori_ori_n391_));
  NO3        o375(.A(ori_ori_n391_), .B(ori_ori_n387_), .C(x2), .Y(ori_ori_n392_));
  OAI220     o376(.A0(ori_ori_n323_), .A1(ori_ori_n283_), .B0(ori_ori_n279_), .B1(ori_ori_n43_), .Y(ori_ori_n393_));
  NA2        o377(.A(ori_ori_n393_), .B(ori_ori_n139_), .Y(ori_ori_n394_));
  NO2        o378(.A(ori_ori_n394_), .B(ori_ori_n54_), .Y(ori_ori_n395_));
  NO2        o379(.A(ori_ori_n395_), .B(ori_ori_n392_), .Y(ori_ori_n396_));
  AOI210     o380(.A0(ori_ori_n396_), .A1(ori_ori_n385_), .B0(ori_ori_n25_), .Y(ori_ori_n397_));
  NA4        o381(.A(ori_ori_n31_), .B(ori_ori_n87_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n398_));
  NO3        o382(.A(ori_ori_n62_), .B(x4), .C(x1), .Y(ori_ori_n399_));
  NO3        o383(.A(ori_ori_n65_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n400_));
  AOI220     o384(.A0(ori_ori_n400_), .A1(ori_ori_n250_), .B0(ori_ori_n399_), .B1(ori_ori_n367_), .Y(ori_ori_n401_));
  NO2        o385(.A(ori_ori_n401_), .B(ori_ori_n98_), .Y(ori_ori_n402_));
  NO3        o386(.A(ori_ori_n254_), .B(ori_ori_n162_), .C(ori_ori_n40_), .Y(ori_ori_n403_));
  OAI210     o387(.A0(ori_ori_n403_), .A1(ori_ori_n402_), .B0(x7), .Y(ori_ori_n404_));
  NA2        o388(.A(ori_ori_n207_), .B(x7), .Y(ori_ori_n405_));
  NA3        o389(.A(ori_ori_n405_), .B(ori_ori_n138_), .C(ori_ori_n121_), .Y(ori_ori_n406_));
  NA3        o390(.A(ori_ori_n406_), .B(ori_ori_n404_), .C(ori_ori_n398_), .Y(ori_ori_n407_));
  OAI210     o391(.A0(ori_ori_n407_), .A1(ori_ori_n397_), .B0(ori_ori_n36_), .Y(ori_ori_n408_));
  INV        o392(.A(ori_ori_n186_), .Y(ori_ori_n409_));
  NO4        o393(.A(ori_ori_n409_), .B(ori_ori_n75_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n410_));
  NA2        o394(.A(ori_ori_n237_), .B(ori_ori_n21_), .Y(ori_ori_n411_));
  NO2        o395(.A(ori_ori_n147_), .B(ori_ori_n122_), .Y(ori_ori_n412_));
  NA2        o396(.A(ori_ori_n412_), .B(ori_ori_n411_), .Y(ori_ori_n413_));
  AOI210     o397(.A0(ori_ori_n413_), .A1(ori_ori_n153_), .B0(ori_ori_n28_), .Y(ori_ori_n414_));
  AOI220     o398(.A0(ori_ori_n335_), .A1(ori_ori_n87_), .B0(ori_ori_n137_), .B1(ori_ori_n182_), .Y(ori_ori_n415_));
  NA3        o399(.A(ori_ori_n415_), .B(ori_ori_n377_), .C(ori_ori_n85_), .Y(ori_ori_n416_));
  NA2        o400(.A(ori_ori_n416_), .B(ori_ori_n163_), .Y(ori_ori_n417_));
  OAI220     o401(.A0(x3), .A1(ori_ori_n66_), .B0(ori_ori_n147_), .B1(ori_ori_n43_), .Y(ori_ori_n418_));
  NA2        o402(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n419_));
  OAI210     o403(.A0(ori_ori_n136_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n420_));
  NO3        o404(.A(ori_ori_n388_), .B(x3), .C(ori_ori_n54_), .Y(ori_ori_n421_));
  NA2        o405(.A(ori_ori_n421_), .B(ori_ori_n420_), .Y(ori_ori_n422_));
  OAI210     o406(.A0(ori_ori_n140_), .A1(ori_ori_n419_), .B0(ori_ori_n422_), .Y(ori_ori_n423_));
  AOI220     o407(.A0(ori_ori_n423_), .A1(x0), .B0(ori_ori_n418_), .B1(ori_ori_n122_), .Y(ori_ori_n424_));
  AOI210     o408(.A0(ori_ori_n424_), .A1(ori_ori_n417_), .B0(ori_ori_n215_), .Y(ori_ori_n425_));
  NO3        o409(.A(ori_ori_n425_), .B(ori_ori_n414_), .C(ori_ori_n410_), .Y(ori_ori_n426_));
  NA3        o410(.A(ori_ori_n426_), .B(ori_ori_n408_), .C(ori_ori_n372_), .Y(ori_ori_n427_));
  AOI210     o411(.A0(ori_ori_n355_), .A1(ori_ori_n25_), .B0(ori_ori_n427_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  INV        m012(.A(mai_mai_n24_), .Y(mai_mai_n29_));
  NO2        m013(.A(x4), .B(x3), .Y(mai_mai_n30_));
  INV        m014(.A(mai_mai_n30_), .Y(mai_mai_n31_));
  OA210      m015(.A0(mai_mai_n31_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n32_));
  NOi31      m016(.An(mai_mai_n23_), .B(mai_mai_n32_), .C(mai_mai_n29_), .Y(mai00));
  NO2        m017(.A(x1), .B(x0), .Y(mai_mai_n34_));
  INV        m018(.A(x6), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n35_), .B(mai_mai_n25_), .Y(mai_mai_n36_));
  NA2        m020(.A(x4), .B(x3), .Y(mai_mai_n37_));
  NO2        m021(.A(mai_mai_n23_), .B(mai_mai_n37_), .Y(mai_mai_n38_));
  NO2        m022(.A(x2), .B(x0), .Y(mai_mai_n39_));
  INV        m023(.A(x3), .Y(mai_mai_n40_));
  NO2        m024(.A(mai_mai_n40_), .B(mai_mai_n18_), .Y(mai_mai_n41_));
  INV        m025(.A(mai_mai_n41_), .Y(mai_mai_n42_));
  NO2        m026(.A(mai_mai_n36_), .B(x4), .Y(mai_mai_n43_));
  OAI210     m027(.A0(mai_mai_n43_), .A1(mai_mai_n42_), .B0(mai_mai_n39_), .Y(mai_mai_n44_));
  INV        m028(.A(x4), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n45_), .B(mai_mai_n17_), .Y(mai_mai_n46_));
  NA2        m030(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n47_));
  OAI210     m031(.A0(mai_mai_n47_), .A1(mai_mai_n20_), .B0(mai_mai_n44_), .Y(mai_mai_n48_));
  AOI210     m032(.A0(mai_mai_n22_), .A1(mai_mai_n19_), .B0(mai_mai_n34_), .Y(mai_mai_n49_));
  INV        m033(.A(x2), .Y(mai_mai_n50_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n17_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n40_), .B(mai_mai_n18_), .Y(mai_mai_n52_));
  NA2        m036(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  OAI210     m037(.A0(mai_mai_n49_), .A1(mai_mai_n31_), .B0(mai_mai_n53_), .Y(mai_mai_n54_));
  NO3        m038(.A(mai_mai_n54_), .B(mai_mai_n48_), .C(mai_mai_n38_), .Y(mai01));
  NA2        m039(.A(x8), .B(x7), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n40_), .B(x1), .Y(mai_mai_n57_));
  INV        m041(.A(x9), .Y(mai_mai_n58_));
  NO2        m042(.A(mai_mai_n58_), .B(mai_mai_n35_), .Y(mai_mai_n59_));
  INV        m043(.A(mai_mai_n59_), .Y(mai_mai_n60_));
  NO3        m044(.A(mai_mai_n60_), .B(mai_mai_n57_), .C(mai_mai_n56_), .Y(mai_mai_n61_));
  NO2        m045(.A(x7), .B(x6), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n63_));
  NO2        m047(.A(x8), .B(x2), .Y(mai_mai_n64_));
  INV        m048(.A(mai_mai_n64_), .Y(mai_mai_n65_));
  NO2        m049(.A(mai_mai_n65_), .B(x1), .Y(mai_mai_n66_));
  OA210      m050(.A0(mai_mai_n66_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .Y(mai_mai_n67_));
  OAI210     m051(.A0(mai_mai_n41_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n68_));
  OAI210     m052(.A0(mai_mai_n52_), .A1(mai_mai_n20_), .B0(mai_mai_n68_), .Y(mai_mai_n69_));
  NAi31      m053(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n70_));
  OAI220     m054(.A0(mai_mai_n70_), .A1(mai_mai_n40_), .B0(mai_mai_n69_), .B1(mai_mai_n67_), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n71_), .A1(mai_mai_n61_), .B0(x4), .Y(mai_mai_n72_));
  NA2        m056(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n73_));
  OAI210     m057(.A0(mai_mai_n73_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n74_));
  NA2        m058(.A(x5), .B(x3), .Y(mai_mai_n75_));
  NO2        m059(.A(x8), .B(x6), .Y(mai_mai_n76_));
  NO4        m060(.A(mai_mai_n76_), .B(mai_mai_n75_), .C(mai_mai_n62_), .D(mai_mai_n50_), .Y(mai_mai_n77_));
  NAi21      m061(.An(x4), .B(x3), .Y(mai_mai_n78_));
  INV        m062(.A(mai_mai_n78_), .Y(mai_mai_n79_));
  NO2        m063(.A(mai_mai_n79_), .B(mai_mai_n22_), .Y(mai_mai_n80_));
  NO2        m064(.A(x4), .B(x2), .Y(mai_mai_n81_));
  NO2        m065(.A(mai_mai_n81_), .B(x3), .Y(mai_mai_n82_));
  NO3        m066(.A(mai_mai_n82_), .B(mai_mai_n80_), .C(mai_mai_n18_), .Y(mai_mai_n83_));
  NO3        m067(.A(mai_mai_n83_), .B(mai_mai_n77_), .C(mai_mai_n74_), .Y(mai_mai_n84_));
  NO4        m068(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n40_), .D(x1), .Y(mai_mai_n85_));
  NA2        m069(.A(mai_mai_n58_), .B(mai_mai_n45_), .Y(mai_mai_n86_));
  INV        m070(.A(mai_mai_n86_), .Y(mai_mai_n87_));
  OAI210     m071(.A0(mai_mai_n85_), .A1(mai_mai_n63_), .B0(mai_mai_n87_), .Y(mai_mai_n88_));
  NA2        m072(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n89_), .B(mai_mai_n25_), .Y(mai_mai_n90_));
  INV        m074(.A(x8), .Y(mai_mai_n91_));
  NA2        m075(.A(x2), .B(x1), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n91_), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n90_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n26_), .Y(mai_mai_n95_));
  AOI210     m079(.A0(mai_mai_n52_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n96_));
  OAI210     m080(.A0(mai_mai_n42_), .A1(mai_mai_n36_), .B0(mai_mai_n45_), .Y(mai_mai_n97_));
  NO3        m081(.A(mai_mai_n97_), .B(mai_mai_n96_), .C(mai_mai_n95_), .Y(mai_mai_n98_));
  NA2        m082(.A(x4), .B(mai_mai_n40_), .Y(mai_mai_n99_));
  NO2        m083(.A(mai_mai_n45_), .B(mai_mai_n50_), .Y(mai_mai_n100_));
  NO2        m084(.A(mai_mai_n99_), .B(x1), .Y(mai_mai_n101_));
  NO2        m085(.A(x3), .B(x2), .Y(mai_mai_n102_));
  NA3        m086(.A(mai_mai_n102_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n103_));
  AOI210     m087(.A0(x8), .A1(x6), .B0(mai_mai_n103_), .Y(mai_mai_n104_));
  NA2        m088(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n105_));
  OAI210     m089(.A0(mai_mai_n105_), .A1(mai_mai_n37_), .B0(mai_mai_n17_), .Y(mai_mai_n106_));
  NO4        m090(.A(mai_mai_n106_), .B(mai_mai_n104_), .C(mai_mai_n101_), .D(mai_mai_n98_), .Y(mai_mai_n107_));
  AO220      m091(.A0(mai_mai_n107_), .A1(mai_mai_n88_), .B0(mai_mai_n84_), .B1(mai_mai_n72_), .Y(mai02));
  NO2        m092(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n109_));
  NO2        m093(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n110_));
  NA2        m094(.A(mai_mai_n50_), .B(mai_mai_n17_), .Y(mai_mai_n111_));
  NA2        m095(.A(mai_mai_n40_), .B(x0), .Y(mai_mai_n112_));
  OAI210     m096(.A0(mai_mai_n86_), .A1(mai_mai_n111_), .B0(mai_mai_n112_), .Y(mai_mai_n113_));
  AOI220     m097(.A0(mai_mai_n113_), .A1(mai_mai_n110_), .B0(mai_mai_n109_), .B1(x4), .Y(mai_mai_n114_));
  NO3        m098(.A(mai_mai_n114_), .B(x7), .C(x5), .Y(mai_mai_n115_));
  NA2        m099(.A(x9), .B(x2), .Y(mai_mai_n116_));
  OR2        m100(.A(x8), .B(x0), .Y(mai_mai_n117_));
  INV        m101(.A(mai_mai_n117_), .Y(mai_mai_n118_));
  NAi21      m102(.An(x2), .B(x8), .Y(mai_mai_n119_));
  INV        m103(.A(mai_mai_n119_), .Y(mai_mai_n120_));
  NO2        m104(.A(mai_mai_n120_), .B(mai_mai_n118_), .Y(mai_mai_n121_));
  NO2        m105(.A(x4), .B(x1), .Y(mai_mai_n122_));
  NA3        m106(.A(mai_mai_n122_), .B(mai_mai_n121_), .C(mai_mai_n56_), .Y(mai_mai_n123_));
  NOi21      m107(.An(x0), .B(x1), .Y(mai_mai_n124_));
  NOi21      m108(.An(x0), .B(x4), .Y(mai_mai_n125_));
  NO2        m109(.A(x8), .B(mai_mai_n58_), .Y(mai_mai_n126_));
  NA2        m110(.A(mai_mai_n126_), .B(mai_mai_n125_), .Y(mai_mai_n127_));
  AOI210     m111(.A0(mai_mai_n127_), .A1(mai_mai_n123_), .B0(mai_mai_n75_), .Y(mai_mai_n128_));
  NO2        m112(.A(x5), .B(mai_mai_n45_), .Y(mai_mai_n129_));
  NA2        m113(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n130_));
  AOI210     m114(.A0(mai_mai_n130_), .A1(mai_mai_n105_), .B0(mai_mai_n112_), .Y(mai_mai_n131_));
  OAI210     m115(.A0(mai_mai_n131_), .A1(mai_mai_n34_), .B0(mai_mai_n129_), .Y(mai_mai_n132_));
  NAi21      m116(.An(x0), .B(x4), .Y(mai_mai_n133_));
  NO2        m117(.A(x7), .B(x0), .Y(mai_mai_n134_));
  NO2        m118(.A(mai_mai_n81_), .B(mai_mai_n100_), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n135_), .B(x3), .Y(mai_mai_n136_));
  NA2        m120(.A(mai_mai_n134_), .B(mai_mai_n136_), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n21_), .B(mai_mai_n40_), .Y(mai_mai_n138_));
  NA2        m122(.A(x5), .B(x0), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n140_));
  NA3        m124(.A(mai_mai_n140_), .B(mai_mai_n139_), .C(mai_mai_n138_), .Y(mai_mai_n141_));
  NA4        m125(.A(mai_mai_n141_), .B(mai_mai_n137_), .C(mai_mai_n132_), .D(mai_mai_n35_), .Y(mai_mai_n142_));
  NO3        m126(.A(mai_mai_n142_), .B(mai_mai_n128_), .C(mai_mai_n115_), .Y(mai_mai_n143_));
  NO3        m127(.A(mai_mai_n75_), .B(mai_mai_n73_), .C(mai_mai_n24_), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n145_));
  AOI220     m129(.A0(mai_mai_n124_), .A1(mai_mai_n145_), .B0(mai_mai_n63_), .B1(mai_mai_n17_), .Y(mai_mai_n146_));
  NO3        m130(.A(mai_mai_n146_), .B(mai_mai_n56_), .C(mai_mai_n58_), .Y(mai_mai_n147_));
  NA2        m131(.A(x7), .B(x3), .Y(mai_mai_n148_));
  NO2        m132(.A(mai_mai_n99_), .B(x5), .Y(mai_mai_n149_));
  NO2        m133(.A(x9), .B(x7), .Y(mai_mai_n150_));
  NOi21      m134(.An(x8), .B(x0), .Y(mai_mai_n151_));
  OA210      m135(.A0(mai_mai_n150_), .A1(x1), .B0(mai_mai_n151_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n40_), .B(x2), .Y(mai_mai_n153_));
  INV        m137(.A(x7), .Y(mai_mai_n154_));
  NA2        m138(.A(mai_mai_n154_), .B(mai_mai_n18_), .Y(mai_mai_n155_));
  NA2        m139(.A(mai_mai_n155_), .B(mai_mai_n153_), .Y(mai_mai_n156_));
  NO2        m140(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n157_));
  NO2        m141(.A(mai_mai_n157_), .B(mai_mai_n125_), .Y(mai_mai_n158_));
  NO2        m142(.A(mai_mai_n158_), .B(mai_mai_n156_), .Y(mai_mai_n159_));
  AOI210     m143(.A0(mai_mai_n152_), .A1(mai_mai_n149_), .B0(mai_mai_n159_), .Y(mai_mai_n160_));
  OAI210     m144(.A0(mai_mai_n148_), .A1(mai_mai_n47_), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  NA2        m145(.A(x5), .B(x1), .Y(mai_mai_n162_));
  INV        m146(.A(mai_mai_n162_), .Y(mai_mai_n163_));
  AOI210     m147(.A0(mai_mai_n163_), .A1(mai_mai_n125_), .B0(mai_mai_n35_), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n58_), .B(mai_mai_n91_), .Y(mai_mai_n165_));
  NAi21      m149(.An(x2), .B(x7), .Y(mai_mai_n166_));
  NO3        m150(.A(mai_mai_n166_), .B(mai_mai_n165_), .C(mai_mai_n45_), .Y(mai_mai_n167_));
  NA2        m151(.A(mai_mai_n167_), .B(mai_mai_n63_), .Y(mai_mai_n168_));
  NA2        m152(.A(mai_mai_n168_), .B(mai_mai_n164_), .Y(mai_mai_n169_));
  NO4        m153(.A(mai_mai_n169_), .B(mai_mai_n161_), .C(mai_mai_n147_), .D(mai_mai_n144_), .Y(mai_mai_n170_));
  NO2        m154(.A(mai_mai_n170_), .B(mai_mai_n143_), .Y(mai_mai_n171_));
  NO2        m155(.A(mai_mai_n139_), .B(mai_mai_n135_), .Y(mai_mai_n172_));
  NA2        m156(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n173_));
  NA2        m157(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n174_));
  NA3        m158(.A(mai_mai_n174_), .B(mai_mai_n173_), .C(mai_mai_n24_), .Y(mai_mai_n175_));
  AN2        m159(.A(mai_mai_n175_), .B(mai_mai_n140_), .Y(mai_mai_n176_));
  NA2        m160(.A(x8), .B(x0), .Y(mai_mai_n177_));
  NO2        m161(.A(mai_mai_n154_), .B(mai_mai_n25_), .Y(mai_mai_n178_));
  NO2        m162(.A(mai_mai_n124_), .B(x4), .Y(mai_mai_n179_));
  NA2        m163(.A(mai_mai_n179_), .B(mai_mai_n178_), .Y(mai_mai_n180_));
  AOI210     m164(.A0(mai_mai_n177_), .A1(mai_mai_n130_), .B0(mai_mai_n180_), .Y(mai_mai_n181_));
  NA2        m165(.A(x2), .B(x0), .Y(mai_mai_n182_));
  NA2        m166(.A(x4), .B(x1), .Y(mai_mai_n183_));
  NAi21      m167(.An(mai_mai_n122_), .B(mai_mai_n183_), .Y(mai_mai_n184_));
  NOi31      m168(.An(mai_mai_n184_), .B(mai_mai_n157_), .C(mai_mai_n182_), .Y(mai_mai_n185_));
  NO4        m169(.A(mai_mai_n185_), .B(mai_mai_n181_), .C(mai_mai_n176_), .D(mai_mai_n172_), .Y(mai_mai_n186_));
  NO2        m170(.A(mai_mai_n186_), .B(mai_mai_n40_), .Y(mai_mai_n187_));
  NO2        m171(.A(mai_mai_n175_), .B(mai_mai_n73_), .Y(mai_mai_n188_));
  INV        m172(.A(mai_mai_n129_), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n105_), .B(mai_mai_n17_), .Y(mai_mai_n190_));
  AOI210     m174(.A0(mai_mai_n34_), .A1(mai_mai_n91_), .B0(mai_mai_n190_), .Y(mai_mai_n191_));
  NO3        m175(.A(mai_mai_n191_), .B(mai_mai_n189_), .C(x7), .Y(mai_mai_n192_));
  NA3        m176(.A(mai_mai_n184_), .B(mai_mai_n189_), .C(mai_mai_n39_), .Y(mai_mai_n193_));
  OAI210     m177(.A0(mai_mai_n174_), .A1(mai_mai_n135_), .B0(mai_mai_n193_), .Y(mai_mai_n194_));
  NO3        m178(.A(mai_mai_n194_), .B(mai_mai_n192_), .C(mai_mai_n188_), .Y(mai_mai_n195_));
  NO2        m179(.A(mai_mai_n195_), .B(x3), .Y(mai_mai_n196_));
  NO3        m180(.A(mai_mai_n196_), .B(mai_mai_n187_), .C(mai_mai_n171_), .Y(mai03));
  NO2        m181(.A(mai_mai_n45_), .B(x3), .Y(mai_mai_n198_));
  NO2        m182(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n199_));
  INV        m183(.A(mai_mai_n199_), .Y(mai_mai_n200_));
  NO2        m184(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n201_));
  OAI210     m185(.A0(mai_mai_n201_), .A1(mai_mai_n25_), .B0(mai_mai_n59_), .Y(mai_mai_n202_));
  OAI220     m186(.A0(mai_mai_n202_), .A1(mai_mai_n17_), .B0(mai_mai_n200_), .B1(mai_mai_n105_), .Y(mai_mai_n203_));
  NA2        m187(.A(mai_mai_n203_), .B(mai_mai_n198_), .Y(mai_mai_n204_));
  NO2        m188(.A(mai_mai_n75_), .B(x6), .Y(mai_mai_n205_));
  NA2        m189(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n206_));
  NO2        m190(.A(mai_mai_n206_), .B(x4), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n208_));
  AO220      m192(.A0(mai_mai_n208_), .A1(mai_mai_n207_), .B0(mai_mai_n205_), .B1(mai_mai_n51_), .Y(mai_mai_n209_));
  NA2        m193(.A(mai_mai_n209_), .B(mai_mai_n58_), .Y(mai_mai_n210_));
  NA2        m194(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n211_));
  NO2        m195(.A(mai_mai_n211_), .B(mai_mai_n206_), .Y(mai_mai_n212_));
  NA2        m196(.A(x9), .B(mai_mai_n50_), .Y(mai_mai_n213_));
  NA2        m197(.A(x9), .B(mai_mai_n212_), .Y(mai_mai_n214_));
  NO3        m198(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n215_));
  NO2        m199(.A(x5), .B(x1), .Y(mai_mai_n216_));
  AOI220     m200(.A0(mai_mai_n216_), .A1(mai_mai_n17_), .B0(mai_mai_n102_), .B1(x5), .Y(mai_mai_n217_));
  NO2        m201(.A(mai_mai_n211_), .B(mai_mai_n173_), .Y(mai_mai_n218_));
  NO3        m202(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n219_));
  NO2        m203(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n220_));
  OAI210     m204(.A0(mai_mai_n217_), .A1(mai_mai_n60_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  AOI220     m205(.A0(mai_mai_n221_), .A1(mai_mai_n45_), .B0(mai_mai_n215_), .B1(mai_mai_n129_), .Y(mai_mai_n222_));
  NA4        m206(.A(mai_mai_n222_), .B(mai_mai_n214_), .C(mai_mai_n210_), .D(mai_mai_n204_), .Y(mai_mai_n223_));
  NO2        m207(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n224_));
  NA2        m208(.A(mai_mai_n224_), .B(mai_mai_n19_), .Y(mai_mai_n225_));
  NO2        m209(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n226_));
  NO2        m210(.A(mai_mai_n226_), .B(x6), .Y(mai_mai_n227_));
  NOi21      m211(.An(mai_mai_n81_), .B(mai_mai_n227_), .Y(mai_mai_n228_));
  NA2        m212(.A(mai_mai_n58_), .B(mai_mai_n91_), .Y(mai_mai_n229_));
  NA3        m213(.A(mai_mai_n229_), .B(mai_mai_n226_), .C(x6), .Y(mai_mai_n230_));
  AOI210     m214(.A0(mai_mai_n230_), .A1(mai_mai_n228_), .B0(mai_mai_n154_), .Y(mai_mai_n231_));
  AO210      m215(.A0(mai_mai_n231_), .A1(mai_mai_n225_), .B0(mai_mai_n178_), .Y(mai_mai_n232_));
  NA2        m216(.A(mai_mai_n40_), .B(mai_mai_n50_), .Y(mai_mai_n233_));
  NA2        m217(.A(mai_mai_n140_), .B(mai_mai_n90_), .Y(mai_mai_n234_));
  NA2        m218(.A(x6), .B(mai_mai_n45_), .Y(mai_mai_n235_));
  OAI210     m219(.A0(mai_mai_n118_), .A1(mai_mai_n76_), .B0(x4), .Y(mai_mai_n236_));
  AOI210     m220(.A0(mai_mai_n236_), .A1(mai_mai_n235_), .B0(mai_mai_n75_), .Y(mai_mai_n237_));
  NO2        m221(.A(mai_mai_n58_), .B(x6), .Y(mai_mai_n238_));
  NO2        m222(.A(mai_mai_n162_), .B(mai_mai_n40_), .Y(mai_mai_n239_));
  OAI210     m223(.A0(mai_mai_n239_), .A1(mai_mai_n218_), .B0(mai_mai_n238_), .Y(mai_mai_n240_));
  NA3        m224(.A(mai_mai_n211_), .B(mai_mai_n129_), .C(x6), .Y(mai_mai_n241_));
  OAI210     m225(.A0(mai_mai_n91_), .A1(mai_mai_n35_), .B0(mai_mai_n63_), .Y(mai_mai_n242_));
  NA3        m226(.A(mai_mai_n242_), .B(mai_mai_n241_), .C(mai_mai_n240_), .Y(mai_mai_n243_));
  OAI210     m227(.A0(mai_mai_n243_), .A1(mai_mai_n237_), .B0(x2), .Y(mai_mai_n244_));
  NA3        m228(.A(mai_mai_n244_), .B(mai_mai_n234_), .C(mai_mai_n232_), .Y(mai_mai_n245_));
  AOI210     m229(.A0(mai_mai_n223_), .A1(x8), .B0(mai_mai_n245_), .Y(mai_mai_n246_));
  NO2        m230(.A(mai_mai_n91_), .B(x3), .Y(mai_mai_n247_));
  NA2        m231(.A(mai_mai_n247_), .B(mai_mai_n207_), .Y(mai_mai_n248_));
  NO2        m232(.A(mai_mai_n89_), .B(mai_mai_n25_), .Y(mai_mai_n249_));
  AOI210     m233(.A0(mai_mai_n227_), .A1(mai_mai_n157_), .B0(mai_mai_n249_), .Y(mai_mai_n250_));
  AOI210     m234(.A0(mai_mai_n250_), .A1(mai_mai_n248_), .B0(x2), .Y(mai_mai_n251_));
  NO2        m235(.A(x4), .B(mai_mai_n50_), .Y(mai_mai_n252_));
  AOI220     m236(.A0(mai_mai_n207_), .A1(mai_mai_n190_), .B0(mai_mai_n252_), .B1(mai_mai_n63_), .Y(mai_mai_n253_));
  NA2        m237(.A(mai_mai_n58_), .B(x6), .Y(mai_mai_n254_));
  NA2        m238(.A(mai_mai_n40_), .B(mai_mai_n17_), .Y(mai_mai_n255_));
  NO2        m239(.A(mai_mai_n255_), .B(mai_mai_n25_), .Y(mai_mai_n256_));
  NA2        m240(.A(mai_mai_n256_), .B(mai_mai_n122_), .Y(mai_mai_n257_));
  NA2        m241(.A(mai_mai_n211_), .B(x6), .Y(mai_mai_n258_));
  NO2        m242(.A(mai_mai_n211_), .B(x6), .Y(mai_mai_n259_));
  NAi21      m243(.An(mai_mai_n165_), .B(mai_mai_n259_), .Y(mai_mai_n260_));
  NA3        m244(.A(mai_mai_n260_), .B(mai_mai_n258_), .C(mai_mai_n145_), .Y(mai_mai_n261_));
  NA4        m245(.A(mai_mai_n261_), .B(mai_mai_n257_), .C(mai_mai_n253_), .D(mai_mai_n154_), .Y(mai_mai_n262_));
  NO2        m246(.A(mai_mai_n139_), .B(mai_mai_n18_), .Y(mai_mai_n263_));
  NAi21      m247(.An(x1), .B(x4), .Y(mai_mai_n264_));
  AOI210     m248(.A0(x3), .A1(x2), .B0(mai_mai_n45_), .Y(mai_mai_n265_));
  OAI210     m249(.A0(mai_mai_n139_), .A1(x3), .B0(mai_mai_n265_), .Y(mai_mai_n266_));
  NA2        m250(.A(mai_mai_n266_), .B(mai_mai_n264_), .Y(mai_mai_n267_));
  INV        m251(.A(mai_mai_n267_), .Y(mai_mai_n268_));
  NA2        m252(.A(mai_mai_n58_), .B(x2), .Y(mai_mai_n269_));
  NO3        m253(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n270_));
  NA2        m254(.A(mai_mai_n105_), .B(mai_mai_n25_), .Y(mai_mai_n271_));
  NA2        m255(.A(x6), .B(x2), .Y(mai_mai_n272_));
  NO2        m256(.A(mai_mai_n272_), .B(mai_mai_n173_), .Y(mai_mai_n273_));
  AOI210     m257(.A0(mai_mai_n271_), .A1(mai_mai_n270_), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  OAI220     m258(.A0(mai_mai_n274_), .A1(mai_mai_n40_), .B0(mai_mai_n179_), .B1(mai_mai_n43_), .Y(mai_mai_n275_));
  NA2        m259(.A(mai_mai_n275_), .B(mai_mai_n268_), .Y(mai_mai_n276_));
  NA2        m260(.A(x9), .B(mai_mai_n40_), .Y(mai_mai_n277_));
  NO2        m261(.A(mai_mai_n277_), .B(mai_mai_n206_), .Y(mai_mai_n278_));
  OR3        m262(.A(mai_mai_n278_), .B(mai_mai_n205_), .C(mai_mai_n149_), .Y(mai_mai_n279_));
  NA2        m263(.A(x4), .B(x0), .Y(mai_mai_n280_));
  NA2        m264(.A(mai_mai_n279_), .B(mai_mai_n39_), .Y(mai_mai_n281_));
  AOI210     m265(.A0(mai_mai_n281_), .A1(mai_mai_n276_), .B0(x8), .Y(mai_mai_n282_));
  INV        m266(.A(mai_mai_n254_), .Y(mai_mai_n283_));
  OAI210     m267(.A0(mai_mai_n263_), .A1(mai_mai_n216_), .B0(mai_mai_n283_), .Y(mai_mai_n284_));
  INV        m268(.A(mai_mai_n177_), .Y(mai_mai_n285_));
  OAI210     m269(.A0(mai_mai_n285_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n286_));
  AOI210     m270(.A0(mai_mai_n286_), .A1(mai_mai_n284_), .B0(mai_mai_n233_), .Y(mai_mai_n287_));
  NO4        m271(.A(mai_mai_n287_), .B(mai_mai_n282_), .C(mai_mai_n262_), .D(mai_mai_n251_), .Y(mai_mai_n288_));
  NO2        m272(.A(mai_mai_n165_), .B(x1), .Y(mai_mai_n289_));
  NO3        m273(.A(mai_mai_n289_), .B(x3), .C(mai_mai_n35_), .Y(mai_mai_n290_));
  OAI210     m274(.A0(mai_mai_n290_), .A1(mai_mai_n259_), .B0(x2), .Y(mai_mai_n291_));
  OAI210     m275(.A0(mai_mai_n285_), .A1(x6), .B0(mai_mai_n41_), .Y(mai_mai_n292_));
  AOI210     m276(.A0(mai_mai_n292_), .A1(mai_mai_n291_), .B0(mai_mai_n189_), .Y(mai_mai_n293_));
  NOi21      m277(.An(mai_mai_n272_), .B(mai_mai_n17_), .Y(mai_mai_n294_));
  NA3        m278(.A(mai_mai_n294_), .B(mai_mai_n216_), .C(mai_mai_n37_), .Y(mai_mai_n295_));
  AOI210     m279(.A0(mai_mai_n35_), .A1(mai_mai_n50_), .B0(x0), .Y(mai_mai_n296_));
  NA3        m280(.A(mai_mai_n296_), .B(mai_mai_n163_), .C(mai_mai_n31_), .Y(mai_mai_n297_));
  NA2        m281(.A(x3), .B(x2), .Y(mai_mai_n298_));
  AOI220     m282(.A0(mai_mai_n298_), .A1(mai_mai_n233_), .B0(mai_mai_n297_), .B1(mai_mai_n295_), .Y(mai_mai_n299_));
  NAi21      m283(.An(x4), .B(x0), .Y(mai_mai_n300_));
  NO3        m284(.A(mai_mai_n300_), .B(mai_mai_n41_), .C(x2), .Y(mai_mai_n301_));
  OAI210     m285(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n301_), .Y(mai_mai_n302_));
  OAI220     m286(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n303_));
  NO2        m287(.A(mai_mai_n296_), .B(mai_mai_n294_), .Y(mai_mai_n304_));
  AOI220     m288(.A0(mai_mai_n304_), .A1(mai_mai_n79_), .B0(mai_mai_n303_), .B1(mai_mai_n30_), .Y(mai_mai_n305_));
  AOI210     m289(.A0(mai_mai_n305_), .A1(mai_mai_n302_), .B0(mai_mai_n25_), .Y(mai_mai_n306_));
  NA3        m290(.A(mai_mai_n35_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n307_));
  OAI210     m291(.A0(mai_mai_n296_), .A1(mai_mai_n294_), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  INV        m292(.A(mai_mai_n218_), .Y(mai_mai_n309_));
  NA2        m293(.A(mai_mai_n35_), .B(mai_mai_n40_), .Y(mai_mai_n310_));
  OR2        m294(.A(mai_mai_n310_), .B(mai_mai_n280_), .Y(mai_mai_n311_));
  OAI220     m295(.A0(mai_mai_n311_), .A1(mai_mai_n162_), .B0(mai_mai_n235_), .B1(mai_mai_n309_), .Y(mai_mai_n312_));
  AO210      m296(.A0(mai_mai_n308_), .A1(mai_mai_n149_), .B0(mai_mai_n312_), .Y(mai_mai_n313_));
  NO4        m297(.A(mai_mai_n313_), .B(mai_mai_n306_), .C(mai_mai_n299_), .D(mai_mai_n293_), .Y(mai_mai_n314_));
  OAI210     m298(.A0(mai_mai_n288_), .A1(mai_mai_n246_), .B0(mai_mai_n314_), .Y(mai04));
  OAI210     m299(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n316_));
  NA3        m300(.A(mai_mai_n316_), .B(mai_mai_n270_), .C(mai_mai_n82_), .Y(mai_mai_n317_));
  NO2        m301(.A(x2), .B(x1), .Y(mai_mai_n318_));
  OAI210     m302(.A0(mai_mai_n255_), .A1(mai_mai_n318_), .B0(mai_mai_n35_), .Y(mai_mai_n319_));
  NO2        m303(.A(mai_mai_n318_), .B(mai_mai_n300_), .Y(mai_mai_n320_));
  AOI210     m304(.A0(mai_mai_n58_), .A1(x4), .B0(mai_mai_n111_), .Y(mai_mai_n321_));
  OAI210     m305(.A0(mai_mai_n321_), .A1(mai_mai_n320_), .B0(mai_mai_n247_), .Y(mai_mai_n322_));
  NO2        m306(.A(mai_mai_n298_), .B(mai_mai_n208_), .Y(mai_mai_n323_));
  NA2        m307(.A(x9), .B(x0), .Y(mai_mai_n324_));
  AOI210     m308(.A0(mai_mai_n89_), .A1(mai_mai_n73_), .B0(mai_mai_n324_), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n325_), .A1(mai_mai_n323_), .B0(mai_mai_n91_), .Y(mai_mai_n326_));
  NA3        m310(.A(mai_mai_n326_), .B(x6), .C(mai_mai_n322_), .Y(mai_mai_n327_));
  NA2        m311(.A(mai_mai_n327_), .B(mai_mai_n319_), .Y(mai_mai_n328_));
  NO2        m312(.A(mai_mai_n213_), .B(mai_mai_n112_), .Y(mai_mai_n329_));
  NO3        m313(.A(mai_mai_n254_), .B(mai_mai_n119_), .C(mai_mai_n18_), .Y(mai_mai_n330_));
  NO2        m314(.A(mai_mai_n330_), .B(mai_mai_n329_), .Y(mai_mai_n331_));
  OAI210     m315(.A0(mai_mai_n117_), .A1(mai_mai_n105_), .B0(mai_mai_n177_), .Y(mai_mai_n332_));
  NA3        m316(.A(mai_mai_n332_), .B(x6), .C(x3), .Y(mai_mai_n333_));
  NOi21      m317(.An(mai_mai_n151_), .B(mai_mai_n130_), .Y(mai_mai_n334_));
  AOI210     m318(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n335_));
  OAI220     m319(.A0(mai_mai_n335_), .A1(mai_mai_n310_), .B0(mai_mai_n269_), .B1(mai_mai_n307_), .Y(mai_mai_n336_));
  AOI210     m320(.A0(mai_mai_n334_), .A1(mai_mai_n59_), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  NA2        m321(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n338_));
  OAI210     m322(.A0(mai_mai_n105_), .A1(mai_mai_n17_), .B0(mai_mai_n338_), .Y(mai_mai_n339_));
  NA2        m323(.A(mai_mai_n339_), .B(mai_mai_n76_), .Y(mai_mai_n340_));
  NA4        m324(.A(mai_mai_n340_), .B(mai_mai_n337_), .C(mai_mai_n333_), .D(mai_mai_n331_), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n110_), .A1(x3), .B0(mai_mai_n301_), .Y(mai_mai_n342_));
  NA3        m326(.A(mai_mai_n229_), .B(mai_mai_n215_), .C(mai_mai_n81_), .Y(mai_mai_n343_));
  NA3        m327(.A(mai_mai_n343_), .B(mai_mai_n342_), .C(mai_mai_n154_), .Y(mai_mai_n344_));
  AOI210     m328(.A0(mai_mai_n341_), .A1(x4), .B0(mai_mai_n344_), .Y(mai_mai_n345_));
  NA3        m329(.A(mai_mai_n320_), .B(mai_mai_n213_), .C(mai_mai_n91_), .Y(mai_mai_n346_));
  NOi21      m330(.An(x4), .B(x0), .Y(mai_mai_n347_));
  XO2        m331(.A(x4), .B(x0), .Y(mai_mai_n348_));
  OAI210     m332(.A0(mai_mai_n348_), .A1(mai_mai_n116_), .B0(mai_mai_n264_), .Y(mai_mai_n349_));
  AOI220     m333(.A0(mai_mai_n349_), .A1(x8), .B0(mai_mai_n347_), .B1(mai_mai_n92_), .Y(mai_mai_n350_));
  AOI210     m334(.A0(mai_mai_n350_), .A1(mai_mai_n346_), .B0(x3), .Y(mai_mai_n351_));
  INV        m335(.A(mai_mai_n92_), .Y(mai_mai_n352_));
  NO2        m336(.A(mai_mai_n91_), .B(x4), .Y(mai_mai_n353_));
  AOI220     m337(.A0(mai_mai_n353_), .A1(mai_mai_n41_), .B0(mai_mai_n125_), .B1(mai_mai_n352_), .Y(mai_mai_n354_));
  NO3        m338(.A(mai_mai_n348_), .B(mai_mai_n165_), .C(x2), .Y(mai_mai_n355_));
  INV        m339(.A(mai_mai_n355_), .Y(mai_mai_n356_));
  NA4        m340(.A(mai_mai_n356_), .B(mai_mai_n354_), .C(mai_mai_n225_), .D(x6), .Y(mai_mai_n357_));
  OAI220     m341(.A0(mai_mai_n300_), .A1(mai_mai_n89_), .B0(mai_mai_n182_), .B1(mai_mai_n91_), .Y(mai_mai_n358_));
  NA2        m342(.A(mai_mai_n358_), .B(mai_mai_n57_), .Y(mai_mai_n359_));
  NO2        m343(.A(mai_mai_n151_), .B(mai_mai_n78_), .Y(mai_mai_n360_));
  NO2        m344(.A(mai_mai_n34_), .B(x2), .Y(mai_mai_n361_));
  NOi21      m345(.An(mai_mai_n122_), .B(mai_mai_n27_), .Y(mai_mai_n362_));
  AOI210     m346(.A0(mai_mai_n361_), .A1(mai_mai_n360_), .B0(mai_mai_n362_), .Y(mai_mai_n363_));
  OAI210     m347(.A0(mai_mai_n359_), .A1(mai_mai_n58_), .B0(mai_mai_n363_), .Y(mai_mai_n364_));
  OAI220     m348(.A0(mai_mai_n364_), .A1(x6), .B0(mai_mai_n357_), .B1(mai_mai_n351_), .Y(mai_mai_n365_));
  OAI210     m349(.A0(mai_mai_n59_), .A1(mai_mai_n45_), .B0(mai_mai_n39_), .Y(mai_mai_n366_));
  OAI210     m350(.A0(mai_mai_n366_), .A1(mai_mai_n91_), .B0(mai_mai_n311_), .Y(mai_mai_n367_));
  AOI210     m351(.A0(mai_mai_n367_), .A1(mai_mai_n18_), .B0(mai_mai_n154_), .Y(mai_mai_n368_));
  AO220      m352(.A0(mai_mai_n368_), .A1(mai_mai_n365_), .B0(mai_mai_n345_), .B1(mai_mai_n328_), .Y(mai_mai_n369_));
  NA2        m353(.A(mai_mai_n81_), .B(x6), .Y(mai_mai_n370_));
  INV        m354(.A(mai_mai_n370_), .Y(mai_mai_n371_));
  AOI220     m355(.A0(mai_mai_n371_), .A1(mai_mai_n34_), .B0(mai_mai_n219_), .B1(mai_mai_n46_), .Y(mai_mai_n372_));
  NA3        m356(.A(mai_mai_n372_), .B(mai_mai_n369_), .C(mai_mai_n317_), .Y(mai_mai_n373_));
  AOI210     m357(.A0(mai_mai_n201_), .A1(x8), .B0(mai_mai_n110_), .Y(mai_mai_n374_));
  NA2        m358(.A(mai_mai_n374_), .B(mai_mai_n338_), .Y(mai_mai_n375_));
  NA3        m359(.A(mai_mai_n375_), .B(mai_mai_n198_), .C(mai_mai_n154_), .Y(mai_mai_n376_));
  OAI210     m360(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n233_), .Y(mai_mai_n377_));
  AO220      m361(.A0(mai_mai_n377_), .A1(mai_mai_n150_), .B0(mai_mai_n109_), .B1(x4), .Y(mai_mai_n378_));
  NA3        m362(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n379_));
  NO2        m363(.A(mai_mai_n379_), .B(mai_mai_n352_), .Y(mai_mai_n380_));
  AOI210     m364(.A0(mai_mai_n378_), .A1(mai_mai_n118_), .B0(mai_mai_n380_), .Y(mai_mai_n381_));
  AOI210     m365(.A0(mai_mai_n381_), .A1(mai_mai_n376_), .B0(mai_mai_n25_), .Y(mai_mai_n382_));
  NA3        m366(.A(mai_mai_n120_), .B(mai_mai_n224_), .C(x0), .Y(mai_mai_n383_));
  AOI210     m367(.A0(mai_mai_n119_), .A1(mai_mai_n117_), .B0(mai_mai_n39_), .Y(mai_mai_n384_));
  NOi31      m368(.An(mai_mai_n384_), .B(x3), .C(mai_mai_n183_), .Y(mai_mai_n385_));
  NA2        m369(.A(mai_mai_n385_), .B(mai_mai_n150_), .Y(mai_mai_n386_));
  NA2        m370(.A(mai_mai_n386_), .B(mai_mai_n383_), .Y(mai_mai_n387_));
  OAI210     m371(.A0(mai_mai_n387_), .A1(mai_mai_n382_), .B0(x6), .Y(mai_mai_n388_));
  OAI210     m372(.A0(mai_mai_n165_), .A1(mai_mai_n45_), .B0(mai_mai_n134_), .Y(mai_mai_n389_));
  AOI210     m373(.A0(mai_mai_n37_), .A1(mai_mai_n31_), .B0(mai_mai_n389_), .Y(mai_mai_n390_));
  NO2        m374(.A(mai_mai_n154_), .B(x0), .Y(mai_mai_n391_));
  AOI220     m375(.A0(mai_mai_n391_), .A1(mai_mai_n224_), .B0(mai_mai_n198_), .B1(mai_mai_n154_), .Y(mai_mai_n392_));
  AOI210     m376(.A0(mai_mai_n126_), .A1(mai_mai_n252_), .B0(x1), .Y(mai_mai_n393_));
  OAI210     m377(.A0(mai_mai_n392_), .A1(x8), .B0(mai_mai_n393_), .Y(mai_mai_n394_));
  NAi31      m378(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n395_));
  OAI210     m379(.A0(mai_mai_n395_), .A1(x4), .B0(mai_mai_n166_), .Y(mai_mai_n396_));
  NA3        m380(.A(mai_mai_n396_), .B(mai_mai_n148_), .C(x9), .Y(mai_mai_n397_));
  NO3        m381(.A(x9), .B(mai_mai_n154_), .C(x0), .Y(mai_mai_n398_));
  AOI220     m382(.A0(mai_mai_n398_), .A1(mai_mai_n247_), .B0(mai_mai_n360_), .B1(mai_mai_n154_), .Y(mai_mai_n399_));
  NA4        m383(.A(mai_mai_n399_), .B(x1), .C(mai_mai_n397_), .D(mai_mai_n47_), .Y(mai_mai_n400_));
  OAI210     m384(.A0(mai_mai_n394_), .A1(mai_mai_n390_), .B0(mai_mai_n400_), .Y(mai_mai_n401_));
  NOi31      m385(.An(mai_mai_n391_), .B(mai_mai_n31_), .C(x8), .Y(mai_mai_n402_));
  INV        m386(.A(mai_mai_n133_), .Y(mai_mai_n403_));
  NO2        m387(.A(mai_mai_n403_), .B(mai_mai_n40_), .Y(mai_mai_n404_));
  NOi31      m388(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n405_));
  NA2        m389(.A(mai_mai_n405_), .B(mai_mai_n347_), .Y(mai_mai_n406_));
  AOI210     m390(.A0(mai_mai_n264_), .A1(mai_mai_n56_), .B0(mai_mai_n124_), .Y(mai_mai_n407_));
  OAI210     m391(.A0(mai_mai_n407_), .A1(x3), .B0(mai_mai_n406_), .Y(mai_mai_n408_));
  NO3        m392(.A(mai_mai_n408_), .B(mai_mai_n404_), .C(x2), .Y(mai_mai_n409_));
  OAI210     m393(.A0(mai_mai_n300_), .A1(mai_mai_n40_), .B0(mai_mai_n348_), .Y(mai_mai_n410_));
  AOI210     m394(.A0(x9), .A1(mai_mai_n45_), .B0(mai_mai_n379_), .Y(mai_mai_n411_));
  AOI220     m395(.A0(mai_mai_n411_), .A1(mai_mai_n91_), .B0(mai_mai_n410_), .B1(mai_mai_n154_), .Y(mai_mai_n412_));
  NO2        m396(.A(mai_mai_n412_), .B(mai_mai_n50_), .Y(mai_mai_n413_));
  NO3        m397(.A(mai_mai_n413_), .B(mai_mai_n409_), .C(mai_mai_n402_), .Y(mai_mai_n414_));
  AOI210     m398(.A0(mai_mai_n414_), .A1(mai_mai_n401_), .B0(mai_mai_n25_), .Y(mai_mai_n415_));
  NO3        m399(.A(mai_mai_n58_), .B(x4), .C(x1), .Y(mai_mai_n416_));
  NO3        m400(.A(mai_mai_n64_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n417_));
  AOI220     m401(.A0(mai_mai_n417_), .A1(mai_mai_n265_), .B0(mai_mai_n416_), .B1(mai_mai_n384_), .Y(mai_mai_n418_));
  NO2        m402(.A(mai_mai_n418_), .B(mai_mai_n102_), .Y(mai_mai_n419_));
  NO3        m403(.A(mai_mai_n269_), .B(mai_mai_n177_), .C(mai_mai_n37_), .Y(mai_mai_n420_));
  OAI210     m404(.A0(mai_mai_n420_), .A1(mai_mai_n419_), .B0(x7), .Y(mai_mai_n421_));
  INV        m405(.A(mai_mai_n421_), .Y(mai_mai_n422_));
  OAI210     m406(.A0(mai_mai_n422_), .A1(mai_mai_n415_), .B0(mai_mai_n35_), .Y(mai_mai_n423_));
  NO2        m407(.A(mai_mai_n398_), .B(mai_mai_n208_), .Y(mai_mai_n424_));
  NO4        m408(.A(mai_mai_n424_), .B(mai_mai_n75_), .C(x4), .D(mai_mai_n50_), .Y(mai_mai_n425_));
  NA2        m409(.A(mai_mai_n395_), .B(mai_mai_n89_), .Y(mai_mai_n426_));
  NA2        m410(.A(mai_mai_n426_), .B(mai_mai_n178_), .Y(mai_mai_n427_));
  OAI220     m411(.A0(mai_mai_n277_), .A1(mai_mai_n65_), .B0(mai_mai_n162_), .B1(mai_mai_n40_), .Y(mai_mai_n428_));
  NA2        m412(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n429_));
  AOI210     m413(.A0(mai_mai_n166_), .A1(mai_mai_n27_), .B0(mai_mai_n70_), .Y(mai_mai_n430_));
  OAI210     m414(.A0(mai_mai_n150_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n431_));
  NO3        m415(.A(mai_mai_n405_), .B(x3), .C(mai_mai_n50_), .Y(mai_mai_n432_));
  AOI210     m416(.A0(mai_mai_n432_), .A1(mai_mai_n431_), .B0(mai_mai_n430_), .Y(mai_mai_n433_));
  OAI210     m417(.A0(mai_mai_n155_), .A1(mai_mai_n429_), .B0(mai_mai_n433_), .Y(mai_mai_n434_));
  AOI220     m418(.A0(mai_mai_n434_), .A1(x0), .B0(mai_mai_n428_), .B1(mai_mai_n134_), .Y(mai_mai_n435_));
  AOI210     m419(.A0(mai_mai_n435_), .A1(mai_mai_n427_), .B0(mai_mai_n235_), .Y(mai_mai_n436_));
  NA2        m420(.A(x9), .B(x5), .Y(mai_mai_n437_));
  NO4        m421(.A(mai_mai_n105_), .B(mai_mai_n437_), .C(mai_mai_n56_), .D(mai_mai_n31_), .Y(mai_mai_n438_));
  NO3        m422(.A(mai_mai_n438_), .B(mai_mai_n436_), .C(mai_mai_n425_), .Y(mai_mai_n439_));
  NA3        m423(.A(mai_mai_n439_), .B(mai_mai_n423_), .C(mai_mai_n388_), .Y(mai_mai_n440_));
  AOI210     m424(.A0(mai_mai_n373_), .A1(mai_mai_n25_), .B0(mai_mai_n440_), .Y(mai05));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  INV        u005(.A(men_men_n19_), .Y(men_men_n22_));
  NA2        u006(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n23_));
  INV        u007(.A(x5), .Y(men_men_n24_));
  NA2        u008(.A(x7), .B(x6), .Y(men_men_n25_));
  NA2        u009(.A(x8), .B(x3), .Y(men_men_n26_));
  NA2        u010(.A(x4), .B(x2), .Y(men_men_n27_));
  NO4        u011(.A(men_men_n27_), .B(men_men_n26_), .C(men_men_n25_), .D(men_men_n24_), .Y(men_men_n28_));
  NO2        u012(.A(men_men_n28_), .B(men_men_n23_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  NOi21      u015(.An(men_men_n22_), .B(men_men_n29_), .Y(men00));
  NO2        u016(.A(x1), .B(x0), .Y(men_men_n33_));
  INV        u017(.A(x6), .Y(men_men_n34_));
  NO2        u018(.A(men_men_n34_), .B(men_men_n24_), .Y(men_men_n35_));
  AN2        u019(.A(x8), .B(x7), .Y(men_men_n36_));
  NA3        u020(.A(men_men_n36_), .B(men_men_n35_), .C(men_men_n33_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n22_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n35_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n50_), .B(men_men_n33_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  OAI210     u039(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n55_), .Y(men_men_n56_));
  NO3        u040(.A(men_men_n56_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u041(.A(x8), .B(x7), .Y(men_men_n58_));
  NA2        u042(.A(men_men_n41_), .B(x1), .Y(men_men_n59_));
  INV        u043(.A(x9), .Y(men_men_n60_));
  NO2        u044(.A(men_men_n60_), .B(men_men_n34_), .Y(men_men_n61_));
  INV        u045(.A(men_men_n61_), .Y(men_men_n62_));
  NO3        u046(.A(men_men_n62_), .B(men_men_n59_), .C(men_men_n58_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n59_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  AN2        u050(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n67_));
  OAI210     u051(.A0(men_men_n42_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n68_));
  OAI210     u052(.A0(men_men_n54_), .A1(men_men_n20_), .B0(men_men_n68_), .Y(men_men_n69_));
  NAi31      u053(.An(x1), .B(x9), .C(x5), .Y(men_men_n70_));
  NO2        u054(.A(men_men_n69_), .B(men_men_n67_), .Y(men_men_n71_));
  OAI210     u055(.A0(men_men_n71_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n72_));
  NA2        u056(.A(men_men_n46_), .B(x2), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n74_));
  NA2        u058(.A(x5), .B(x3), .Y(men_men_n75_));
  NO2        u059(.A(x8), .B(x6), .Y(men_men_n76_));
  NO4        u060(.A(men_men_n76_), .B(men_men_n75_), .C(men_men_n64_), .D(men_men_n52_), .Y(men_men_n77_));
  NAi21      u061(.An(x4), .B(x3), .Y(men_men_n78_));
  INV        u062(.A(men_men_n78_), .Y(men_men_n79_));
  NO2        u063(.A(x4), .B(x2), .Y(men_men_n80_));
  NO2        u064(.A(men_men_n80_), .B(x3), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n78_), .B(men_men_n18_), .Y(men_men_n82_));
  NO3        u066(.A(men_men_n82_), .B(men_men_n77_), .C(men_men_n74_), .Y(men_men_n83_));
  NO4        u067(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n84_));
  NA2        u068(.A(men_men_n60_), .B(men_men_n46_), .Y(men_men_n85_));
  INV        u069(.A(men_men_n85_), .Y(men_men_n86_));
  OAI210     u070(.A0(men_men_n84_), .A1(men_men_n65_), .B0(men_men_n86_), .Y(men_men_n87_));
  NA2        u071(.A(x3), .B(men_men_n18_), .Y(men_men_n88_));
  NO2        u072(.A(men_men_n88_), .B(men_men_n24_), .Y(men_men_n89_));
  INV        u073(.A(x8), .Y(men_men_n90_));
  NA2        u074(.A(x2), .B(x1), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n89_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n25_), .Y(men_men_n94_));
  AOI210     u078(.A0(men_men_n54_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n95_));
  OAI210     u079(.A0(men_men_n43_), .A1(men_men_n35_), .B0(men_men_n46_), .Y(men_men_n96_));
  NO3        u080(.A(men_men_n96_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n97_));
  NA2        u081(.A(x4), .B(men_men_n41_), .Y(men_men_n98_));
  NO2        u082(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n99_));
  OAI210     u083(.A0(men_men_n99_), .A1(men_men_n41_), .B0(men_men_n18_), .Y(men_men_n100_));
  AOI210     u084(.A0(men_men_n98_), .A1(men_men_n50_), .B0(men_men_n100_), .Y(men_men_n101_));
  NO2        u085(.A(x3), .B(x2), .Y(men_men_n102_));
  NA3        u086(.A(men_men_n102_), .B(men_men_n25_), .C(men_men_n24_), .Y(men_men_n103_));
  AOI210     u087(.A0(x8), .A1(x6), .B0(men_men_n103_), .Y(men_men_n104_));
  NA2        u088(.A(men_men_n52_), .B(x1), .Y(men_men_n105_));
  OAI210     u089(.A0(men_men_n105_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n106_));
  NO4        u090(.A(men_men_n106_), .B(men_men_n104_), .C(men_men_n101_), .D(men_men_n97_), .Y(men_men_n107_));
  AO220      u091(.A0(men_men_n107_), .A1(men_men_n87_), .B0(men_men_n83_), .B1(men_men_n72_), .Y(men02));
  NO2        u092(.A(x3), .B(men_men_n52_), .Y(men_men_n109_));
  NO2        u093(.A(x8), .B(men_men_n18_), .Y(men_men_n110_));
  NA2        u094(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n111_));
  NA2        u095(.A(men_men_n41_), .B(x0), .Y(men_men_n112_));
  OAI210     u096(.A0(men_men_n85_), .A1(men_men_n111_), .B0(men_men_n112_), .Y(men_men_n113_));
  AOI220     u097(.A0(men_men_n113_), .A1(men_men_n110_), .B0(men_men_n109_), .B1(x4), .Y(men_men_n114_));
  NO3        u098(.A(men_men_n114_), .B(x7), .C(x5), .Y(men_men_n115_));
  NA2        u099(.A(x9), .B(x2), .Y(men_men_n116_));
  OR2        u100(.A(x8), .B(x0), .Y(men_men_n117_));
  INV        u101(.A(men_men_n117_), .Y(men_men_n118_));
  INV        u102(.A(x2), .Y(men_men_n119_));
  OAI220     u103(.A0(men_men_n119_), .A1(men_men_n118_), .B0(men_men_n116_), .B1(x7), .Y(men_men_n120_));
  NO2        u104(.A(x4), .B(x1), .Y(men_men_n121_));
  NA3        u105(.A(men_men_n121_), .B(men_men_n120_), .C(men_men_n58_), .Y(men_men_n122_));
  NOi21      u106(.An(x0), .B(x1), .Y(men_men_n123_));
  NO3        u107(.A(x9), .B(x8), .C(x7), .Y(men_men_n124_));
  NOi21      u108(.An(x0), .B(x4), .Y(men_men_n125_));
  NAi21      u109(.An(x8), .B(x7), .Y(men_men_n126_));
  NA2        u110(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n127_));
  AOI210     u111(.A0(men_men_n127_), .A1(men_men_n122_), .B0(men_men_n75_), .Y(men_men_n128_));
  NO2        u112(.A(x5), .B(men_men_n46_), .Y(men_men_n129_));
  NA2        u113(.A(x2), .B(men_men_n18_), .Y(men_men_n130_));
  AOI210     u114(.A0(men_men_n130_), .A1(men_men_n105_), .B0(men_men_n112_), .Y(men_men_n131_));
  OAI210     u115(.A0(men_men_n131_), .A1(men_men_n33_), .B0(men_men_n129_), .Y(men_men_n132_));
  NAi21      u116(.An(x0), .B(x4), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n133_), .B(x1), .Y(men_men_n134_));
  NO2        u118(.A(x7), .B(x0), .Y(men_men_n135_));
  NO2        u119(.A(men_men_n80_), .B(men_men_n99_), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n136_), .B(x3), .Y(men_men_n137_));
  OAI210     u121(.A0(men_men_n135_), .A1(men_men_n134_), .B0(men_men_n137_), .Y(men_men_n138_));
  NA2        u122(.A(x5), .B(x0), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n46_), .B(x2), .Y(men_men_n140_));
  NA3        u124(.A(men_men_n138_), .B(men_men_n132_), .C(men_men_n34_), .Y(men_men_n141_));
  NO3        u125(.A(men_men_n141_), .B(men_men_n128_), .C(men_men_n115_), .Y(men_men_n142_));
  NO3        u126(.A(men_men_n75_), .B(men_men_n73_), .C(men_men_n23_), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n27_), .B(men_men_n24_), .Y(men_men_n144_));
  AOI220     u128(.A0(men_men_n123_), .A1(men_men_n144_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n145_));
  NO3        u129(.A(men_men_n145_), .B(men_men_n58_), .C(men_men_n60_), .Y(men_men_n146_));
  NA2        u130(.A(x7), .B(x3), .Y(men_men_n147_));
  NO2        u131(.A(men_men_n98_), .B(x5), .Y(men_men_n148_));
  NO2        u132(.A(x9), .B(x7), .Y(men_men_n149_));
  NOi21      u133(.An(x8), .B(x0), .Y(men_men_n150_));
  NO2        u134(.A(men_men_n41_), .B(x2), .Y(men_men_n151_));
  INV        u135(.A(x7), .Y(men_men_n152_));
  NA2        u136(.A(men_men_n152_), .B(men_men_n18_), .Y(men_men_n153_));
  AOI220     u137(.A0(men_men_n153_), .A1(men_men_n151_), .B0(men_men_n109_), .B1(men_men_n36_), .Y(men_men_n154_));
  NO2        u138(.A(men_men_n24_), .B(x4), .Y(men_men_n155_));
  NO2        u139(.A(men_men_n155_), .B(men_men_n125_), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n156_), .B(men_men_n154_), .Y(men_men_n157_));
  AOI210     u141(.A0(men_men_n150_), .A1(men_men_n148_), .B0(men_men_n157_), .Y(men_men_n158_));
  OAI210     u142(.A0(men_men_n147_), .A1(men_men_n48_), .B0(men_men_n158_), .Y(men_men_n159_));
  NA2        u143(.A(x5), .B(x1), .Y(men_men_n160_));
  INV        u144(.A(men_men_n160_), .Y(men_men_n161_));
  AOI210     u145(.A0(men_men_n161_), .A1(men_men_n125_), .B0(men_men_n34_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n60_), .B(men_men_n90_), .Y(men_men_n163_));
  NAi21      u147(.An(x2), .B(x7), .Y(men_men_n164_));
  NO3        u148(.A(men_men_n164_), .B(men_men_n163_), .C(men_men_n46_), .Y(men_men_n165_));
  NA2        u149(.A(men_men_n165_), .B(men_men_n65_), .Y(men_men_n166_));
  NAi31      u150(.An(men_men_n75_), .B(men_men_n36_), .C(men_men_n33_), .Y(men_men_n167_));
  NA3        u151(.A(men_men_n167_), .B(men_men_n166_), .C(men_men_n162_), .Y(men_men_n168_));
  NO4        u152(.A(men_men_n168_), .B(men_men_n159_), .C(men_men_n146_), .D(men_men_n143_), .Y(men_men_n169_));
  NO2        u153(.A(men_men_n169_), .B(men_men_n142_), .Y(men_men_n170_));
  NO2        u154(.A(men_men_n139_), .B(men_men_n136_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n24_), .B(men_men_n18_), .Y(men_men_n172_));
  NA2        u156(.A(men_men_n24_), .B(men_men_n17_), .Y(men_men_n173_));
  NA3        u157(.A(men_men_n173_), .B(men_men_n172_), .C(men_men_n23_), .Y(men_men_n174_));
  AN2        u158(.A(men_men_n174_), .B(men_men_n140_), .Y(men_men_n175_));
  NA2        u159(.A(x8), .B(x0), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n152_), .B(men_men_n24_), .Y(men_men_n177_));
  NO2        u161(.A(men_men_n123_), .B(x4), .Y(men_men_n178_));
  NA2        u162(.A(men_men_n178_), .B(men_men_n177_), .Y(men_men_n179_));
  AOI210     u163(.A0(men_men_n176_), .A1(men_men_n130_), .B0(men_men_n179_), .Y(men_men_n180_));
  NA2        u164(.A(x2), .B(x0), .Y(men_men_n181_));
  NA2        u165(.A(x4), .B(x1), .Y(men_men_n182_));
  NAi21      u166(.An(men_men_n121_), .B(men_men_n182_), .Y(men_men_n183_));
  NOi31      u167(.An(men_men_n183_), .B(men_men_n155_), .C(men_men_n181_), .Y(men_men_n184_));
  NO4        u168(.A(men_men_n184_), .B(men_men_n180_), .C(men_men_n175_), .D(men_men_n171_), .Y(men_men_n185_));
  NO2        u169(.A(men_men_n185_), .B(men_men_n41_), .Y(men_men_n186_));
  NO2        u170(.A(men_men_n174_), .B(men_men_n73_), .Y(men_men_n187_));
  INV        u171(.A(men_men_n129_), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n105_), .B(men_men_n17_), .Y(men_men_n189_));
  AOI210     u173(.A0(men_men_n33_), .A1(men_men_n90_), .B0(men_men_n189_), .Y(men_men_n190_));
  NO3        u174(.A(men_men_n190_), .B(men_men_n188_), .C(x7), .Y(men_men_n191_));
  NA3        u175(.A(men_men_n183_), .B(men_men_n188_), .C(men_men_n40_), .Y(men_men_n192_));
  OAI210     u176(.A0(men_men_n173_), .A1(men_men_n136_), .B0(men_men_n192_), .Y(men_men_n193_));
  NO3        u177(.A(men_men_n193_), .B(men_men_n191_), .C(men_men_n187_), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n194_), .B(x3), .Y(men_men_n195_));
  NO3        u179(.A(men_men_n195_), .B(men_men_n186_), .C(men_men_n170_), .Y(men03));
  NO2        u180(.A(men_men_n46_), .B(x3), .Y(men_men_n197_));
  NO2        u181(.A(x6), .B(men_men_n24_), .Y(men_men_n198_));
  INV        u182(.A(men_men_n198_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n52_), .B(x1), .Y(men_men_n200_));
  OAI210     u184(.A0(men_men_n200_), .A1(men_men_n24_), .B0(men_men_n61_), .Y(men_men_n201_));
  OAI220     u185(.A0(men_men_n201_), .A1(men_men_n17_), .B0(men_men_n199_), .B1(men_men_n105_), .Y(men_men_n202_));
  NA2        u186(.A(men_men_n202_), .B(men_men_n197_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n75_), .B(x6), .Y(men_men_n204_));
  NA2        u188(.A(x6), .B(men_men_n24_), .Y(men_men_n205_));
  NO2        u189(.A(men_men_n205_), .B(x4), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n18_), .B(x0), .Y(men_men_n207_));
  AO220      u191(.A0(men_men_n207_), .A1(men_men_n206_), .B0(men_men_n204_), .B1(men_men_n53_), .Y(men_men_n208_));
  INV        u192(.A(men_men_n208_), .Y(men_men_n209_));
  NA2        u193(.A(x3), .B(men_men_n17_), .Y(men_men_n210_));
  INV        u194(.A(men_men_n205_), .Y(men_men_n211_));
  AOI210     u195(.A0(men_men_n24_), .A1(x3), .B0(men_men_n181_), .Y(men_men_n212_));
  NA2        u196(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n213_));
  NO2        u197(.A(x5), .B(x1), .Y(men_men_n214_));
  AOI220     u198(.A0(men_men_n214_), .A1(men_men_n17_), .B0(men_men_n102_), .B1(x5), .Y(men_men_n215_));
  NO2        u199(.A(men_men_n210_), .B(men_men_n172_), .Y(men_men_n216_));
  INV        u200(.A(men_men_n216_), .Y(men_men_n217_));
  OAI210     u201(.A0(men_men_n215_), .A1(men_men_n62_), .B0(men_men_n217_), .Y(men_men_n218_));
  NA2        u202(.A(men_men_n218_), .B(men_men_n46_), .Y(men_men_n219_));
  NA4        u203(.A(men_men_n219_), .B(men_men_n213_), .C(men_men_n209_), .D(men_men_n203_), .Y(men_men_n220_));
  NO2        u204(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n221_));
  NA2        u205(.A(men_men_n221_), .B(men_men_n19_), .Y(men_men_n222_));
  NO2        u206(.A(x3), .B(men_men_n17_), .Y(men_men_n223_));
  NO2        u207(.A(men_men_n223_), .B(x6), .Y(men_men_n224_));
  NOi21      u208(.An(men_men_n80_), .B(men_men_n224_), .Y(men_men_n225_));
  NA2        u209(.A(men_men_n60_), .B(men_men_n90_), .Y(men_men_n226_));
  NA2        u210(.A(men_men_n223_), .B(x6), .Y(men_men_n227_));
  AOI210     u211(.A0(men_men_n227_), .A1(men_men_n225_), .B0(men_men_n152_), .Y(men_men_n228_));
  OR2        u212(.A(men_men_n228_), .B(men_men_n177_), .Y(men_men_n229_));
  NA2        u213(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n230_));
  OAI210     u214(.A0(men_men_n230_), .A1(men_men_n24_), .B0(men_men_n173_), .Y(men_men_n231_));
  NO3        u215(.A(men_men_n182_), .B(men_men_n60_), .C(x6), .Y(men_men_n232_));
  AOI220     u216(.A0(men_men_n232_), .A1(men_men_n231_), .B0(men_men_n140_), .B1(men_men_n89_), .Y(men_men_n233_));
  NA2        u217(.A(x6), .B(men_men_n46_), .Y(men_men_n234_));
  OAI210     u218(.A0(men_men_n118_), .A1(men_men_n76_), .B0(x4), .Y(men_men_n235_));
  AOI210     u219(.A0(men_men_n235_), .A1(men_men_n234_), .B0(men_men_n75_), .Y(men_men_n236_));
  NA2        u220(.A(men_men_n198_), .B(men_men_n134_), .Y(men_men_n237_));
  NA3        u221(.A(men_men_n210_), .B(men_men_n129_), .C(x6), .Y(men_men_n238_));
  OAI210     u222(.A0(men_men_n90_), .A1(men_men_n34_), .B0(men_men_n65_), .Y(men_men_n239_));
  NA3        u223(.A(men_men_n239_), .B(men_men_n238_), .C(men_men_n237_), .Y(men_men_n240_));
  OAI210     u224(.A0(men_men_n240_), .A1(men_men_n236_), .B0(x2), .Y(men_men_n241_));
  NA3        u225(.A(men_men_n241_), .B(men_men_n233_), .C(men_men_n229_), .Y(men_men_n242_));
  AOI210     u226(.A0(men_men_n220_), .A1(x8), .B0(men_men_n242_), .Y(men_men_n243_));
  NO2        u227(.A(men_men_n90_), .B(x3), .Y(men_men_n244_));
  NA2        u228(.A(men_men_n244_), .B(men_men_n206_), .Y(men_men_n245_));
  NO3        u229(.A(men_men_n88_), .B(men_men_n76_), .C(men_men_n24_), .Y(men_men_n246_));
  AOI210     u230(.A0(men_men_n224_), .A1(men_men_n155_), .B0(men_men_n246_), .Y(men_men_n247_));
  AOI210     u231(.A0(men_men_n247_), .A1(men_men_n245_), .B0(x2), .Y(men_men_n248_));
  NO2        u232(.A(x4), .B(men_men_n52_), .Y(men_men_n249_));
  AOI220     u233(.A0(men_men_n206_), .A1(men_men_n189_), .B0(men_men_n249_), .B1(men_men_n65_), .Y(men_men_n250_));
  NA2        u234(.A(men_men_n60_), .B(x6), .Y(men_men_n251_));
  NA3        u235(.A(men_men_n24_), .B(x3), .C(x2), .Y(men_men_n252_));
  AOI210     u236(.A0(men_men_n252_), .A1(men_men_n139_), .B0(men_men_n251_), .Y(men_men_n253_));
  NA2        u237(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n254_));
  NO2        u238(.A(men_men_n254_), .B(men_men_n24_), .Y(men_men_n255_));
  OAI210     u239(.A0(men_men_n255_), .A1(men_men_n253_), .B0(men_men_n121_), .Y(men_men_n256_));
  NA2        u240(.A(men_men_n210_), .B(x6), .Y(men_men_n257_));
  NO2        u241(.A(men_men_n210_), .B(x6), .Y(men_men_n258_));
  NAi21      u242(.An(men_men_n163_), .B(men_men_n258_), .Y(men_men_n259_));
  NA3        u243(.A(men_men_n259_), .B(men_men_n257_), .C(men_men_n144_), .Y(men_men_n260_));
  NA4        u244(.A(men_men_n260_), .B(men_men_n256_), .C(men_men_n250_), .D(men_men_n152_), .Y(men_men_n261_));
  NA2        u245(.A(men_men_n198_), .B(men_men_n223_), .Y(men_men_n262_));
  NO2        u246(.A(x9), .B(x6), .Y(men_men_n263_));
  NO2        u247(.A(men_men_n139_), .B(men_men_n18_), .Y(men_men_n264_));
  NAi21      u248(.An(men_men_n264_), .B(men_men_n252_), .Y(men_men_n265_));
  NAi21      u249(.An(x1), .B(x4), .Y(men_men_n266_));
  OAI210     u250(.A0(men_men_n139_), .A1(x3), .B0(x4), .Y(men_men_n267_));
  AOI220     u251(.A0(men_men_n267_), .A1(men_men_n266_), .B0(men_men_n265_), .B1(men_men_n263_), .Y(men_men_n268_));
  NA2        u252(.A(men_men_n268_), .B(men_men_n262_), .Y(men_men_n269_));
  NA2        u253(.A(men_men_n60_), .B(x2), .Y(men_men_n270_));
  NO2        u254(.A(men_men_n270_), .B(men_men_n262_), .Y(men_men_n271_));
  NO3        u255(.A(x9), .B(x6), .C(x0), .Y(men_men_n272_));
  NA2        u256(.A(men_men_n105_), .B(men_men_n24_), .Y(men_men_n273_));
  NA2        u257(.A(x6), .B(x2), .Y(men_men_n274_));
  NO2        u258(.A(men_men_n274_), .B(men_men_n172_), .Y(men_men_n275_));
  AOI210     u259(.A0(men_men_n273_), .A1(men_men_n272_), .B0(men_men_n275_), .Y(men_men_n276_));
  OAI220     u260(.A0(men_men_n276_), .A1(men_men_n41_), .B0(men_men_n178_), .B1(men_men_n44_), .Y(men_men_n277_));
  OAI210     u261(.A0(men_men_n277_), .A1(men_men_n271_), .B0(men_men_n269_), .Y(men_men_n278_));
  NA2        u262(.A(x4), .B(x0), .Y(men_men_n279_));
  NO3        u263(.A(men_men_n70_), .B(men_men_n279_), .C(x6), .Y(men_men_n280_));
  AOI210     u264(.A0(men_men_n204_), .A1(men_men_n40_), .B0(men_men_n280_), .Y(men_men_n281_));
  AOI210     u265(.A0(men_men_n281_), .A1(men_men_n278_), .B0(x8), .Y(men_men_n282_));
  NA2        u266(.A(men_men_n214_), .B(x6), .Y(men_men_n283_));
  OAI210     u267(.A0(x0), .A1(x4), .B0(men_men_n20_), .Y(men_men_n284_));
  AOI210     u268(.A0(men_men_n284_), .A1(men_men_n283_), .B0(men_men_n230_), .Y(men_men_n285_));
  NO4        u269(.A(men_men_n285_), .B(men_men_n282_), .C(men_men_n261_), .D(men_men_n248_), .Y(men_men_n286_));
  NO2        u270(.A(men_men_n163_), .B(x1), .Y(men_men_n287_));
  NO3        u271(.A(men_men_n287_), .B(x3), .C(men_men_n34_), .Y(men_men_n288_));
  OAI210     u272(.A0(men_men_n288_), .A1(men_men_n258_), .B0(x2), .Y(men_men_n289_));
  OAI210     u273(.A0(x0), .A1(x6), .B0(men_men_n42_), .Y(men_men_n290_));
  AOI210     u274(.A0(men_men_n290_), .A1(men_men_n289_), .B0(men_men_n188_), .Y(men_men_n291_));
  NOi21      u275(.An(men_men_n274_), .B(men_men_n17_), .Y(men_men_n292_));
  NA3        u276(.A(men_men_n292_), .B(men_men_n214_), .C(men_men_n38_), .Y(men_men_n293_));
  AOI210     u277(.A0(men_men_n34_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n294_));
  NA3        u278(.A(men_men_n294_), .B(men_men_n161_), .C(men_men_n31_), .Y(men_men_n295_));
  NA2        u279(.A(x3), .B(x2), .Y(men_men_n296_));
  AOI220     u280(.A0(men_men_n296_), .A1(men_men_n230_), .B0(men_men_n295_), .B1(men_men_n293_), .Y(men_men_n297_));
  NAi21      u281(.An(x4), .B(x0), .Y(men_men_n298_));
  NO3        u282(.A(men_men_n298_), .B(men_men_n42_), .C(x2), .Y(men_men_n299_));
  OAI210     u283(.A0(x6), .A1(men_men_n18_), .B0(men_men_n299_), .Y(men_men_n300_));
  OAI220     u284(.A0(men_men_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n301_));
  NO2        u285(.A(x9), .B(x8), .Y(men_men_n302_));
  NA3        u286(.A(men_men_n302_), .B(men_men_n34_), .C(men_men_n52_), .Y(men_men_n303_));
  OAI210     u287(.A0(men_men_n294_), .A1(men_men_n292_), .B0(men_men_n303_), .Y(men_men_n304_));
  AOI220     u288(.A0(men_men_n304_), .A1(men_men_n79_), .B0(men_men_n301_), .B1(men_men_n30_), .Y(men_men_n305_));
  AOI210     u289(.A0(men_men_n305_), .A1(men_men_n300_), .B0(men_men_n24_), .Y(men_men_n306_));
  NA3        u290(.A(men_men_n34_), .B(x1), .C(men_men_n17_), .Y(men_men_n307_));
  OAI210     u291(.A0(men_men_n294_), .A1(men_men_n292_), .B0(men_men_n307_), .Y(men_men_n308_));
  INV        u292(.A(men_men_n216_), .Y(men_men_n309_));
  NA2        u293(.A(men_men_n34_), .B(men_men_n41_), .Y(men_men_n310_));
  OR2        u294(.A(men_men_n310_), .B(men_men_n279_), .Y(men_men_n311_));
  OAI220     u295(.A0(men_men_n311_), .A1(men_men_n160_), .B0(men_men_n234_), .B1(men_men_n309_), .Y(men_men_n312_));
  AO210      u296(.A0(men_men_n308_), .A1(men_men_n148_), .B0(men_men_n312_), .Y(men_men_n313_));
  NO4        u297(.A(men_men_n313_), .B(men_men_n306_), .C(men_men_n297_), .D(men_men_n291_), .Y(men_men_n314_));
  OAI210     u298(.A0(men_men_n286_), .A1(men_men_n243_), .B0(men_men_n314_), .Y(men04));
  OAI210     u299(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n316_));
  NA3        u300(.A(men_men_n316_), .B(men_men_n272_), .C(men_men_n81_), .Y(men_men_n317_));
  NO2        u301(.A(x2), .B(x1), .Y(men_men_n318_));
  OAI210     u302(.A0(men_men_n254_), .A1(men_men_n318_), .B0(men_men_n34_), .Y(men_men_n319_));
  NO2        u303(.A(men_men_n318_), .B(men_men_n298_), .Y(men_men_n320_));
  AOI210     u304(.A0(men_men_n60_), .A1(x4), .B0(men_men_n111_), .Y(men_men_n321_));
  OAI210     u305(.A0(men_men_n321_), .A1(men_men_n320_), .B0(men_men_n244_), .Y(men_men_n322_));
  NO2        u306(.A(men_men_n270_), .B(men_men_n88_), .Y(men_men_n323_));
  NO2        u307(.A(men_men_n323_), .B(men_men_n34_), .Y(men_men_n324_));
  NO2        u308(.A(men_men_n296_), .B(men_men_n207_), .Y(men_men_n325_));
  NA2        u309(.A(men_men_n325_), .B(men_men_n90_), .Y(men_men_n326_));
  NA3        u310(.A(men_men_n326_), .B(men_men_n324_), .C(men_men_n322_), .Y(men_men_n327_));
  NA2        u311(.A(men_men_n327_), .B(men_men_n319_), .Y(men_men_n328_));
  NO2        u312(.A(x2), .B(men_men_n112_), .Y(men_men_n329_));
  NO3        u313(.A(men_men_n251_), .B(x2), .C(men_men_n18_), .Y(men_men_n330_));
  NO2        u314(.A(men_men_n330_), .B(men_men_n329_), .Y(men_men_n331_));
  NA3        u315(.A(men_men_n448_), .B(x6), .C(x3), .Y(men_men_n332_));
  NOi21      u316(.An(men_men_n150_), .B(men_men_n130_), .Y(men_men_n333_));
  AOI210     u317(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n334_));
  OAI220     u318(.A0(men_men_n334_), .A1(men_men_n310_), .B0(men_men_n270_), .B1(men_men_n307_), .Y(men_men_n335_));
  AOI210     u319(.A0(men_men_n333_), .A1(men_men_n61_), .B0(men_men_n335_), .Y(men_men_n336_));
  NA2        u320(.A(men_men_n323_), .B(men_men_n90_), .Y(men_men_n337_));
  NA4        u321(.A(men_men_n337_), .B(men_men_n336_), .C(men_men_n332_), .D(men_men_n331_), .Y(men_men_n338_));
  OAI210     u322(.A0(men_men_n110_), .A1(x3), .B0(men_men_n299_), .Y(men_men_n339_));
  NA2        u323(.A(men_men_n339_), .B(men_men_n152_), .Y(men_men_n340_));
  AOI210     u324(.A0(men_men_n338_), .A1(x4), .B0(men_men_n340_), .Y(men_men_n341_));
  NOi21      u325(.An(x4), .B(x0), .Y(men_men_n342_));
  XO2        u326(.A(x4), .B(x0), .Y(men_men_n343_));
  OAI210     u327(.A0(men_men_n343_), .A1(men_men_n116_), .B0(men_men_n266_), .Y(men_men_n344_));
  AOI220     u328(.A0(men_men_n344_), .A1(x8), .B0(men_men_n342_), .B1(men_men_n91_), .Y(men_men_n345_));
  NO2        u329(.A(men_men_n345_), .B(x3), .Y(men_men_n346_));
  INV        u330(.A(men_men_n91_), .Y(men_men_n347_));
  NO2        u331(.A(men_men_n90_), .B(x4), .Y(men_men_n348_));
  AOI220     u332(.A0(men_men_n348_), .A1(men_men_n42_), .B0(men_men_n125_), .B1(men_men_n347_), .Y(men_men_n349_));
  NO3        u333(.A(men_men_n343_), .B(men_men_n163_), .C(x2), .Y(men_men_n350_));
  NO3        u334(.A(men_men_n226_), .B(men_men_n27_), .C(men_men_n23_), .Y(men_men_n351_));
  NO2        u335(.A(men_men_n351_), .B(men_men_n350_), .Y(men_men_n352_));
  NA4        u336(.A(men_men_n352_), .B(men_men_n349_), .C(men_men_n222_), .D(x6), .Y(men_men_n353_));
  OAI220     u337(.A0(men_men_n298_), .A1(men_men_n88_), .B0(men_men_n181_), .B1(men_men_n90_), .Y(men_men_n354_));
  NO2        u338(.A(men_men_n41_), .B(x0), .Y(men_men_n355_));
  OR2        u339(.A(men_men_n348_), .B(men_men_n355_), .Y(men_men_n356_));
  NO2        u340(.A(men_men_n150_), .B(men_men_n105_), .Y(men_men_n357_));
  AOI220     u341(.A0(men_men_n357_), .A1(men_men_n356_), .B0(men_men_n354_), .B1(men_men_n59_), .Y(men_men_n358_));
  NO2        u342(.A(men_men_n150_), .B(men_men_n78_), .Y(men_men_n359_));
  NO2        u343(.A(men_men_n33_), .B(x2), .Y(men_men_n360_));
  NOi21      u344(.An(men_men_n121_), .B(men_men_n26_), .Y(men_men_n361_));
  AOI210     u345(.A0(men_men_n360_), .A1(men_men_n359_), .B0(men_men_n361_), .Y(men_men_n362_));
  OAI210     u346(.A0(men_men_n358_), .A1(men_men_n60_), .B0(men_men_n362_), .Y(men_men_n363_));
  OAI220     u347(.A0(men_men_n363_), .A1(x6), .B0(men_men_n353_), .B1(men_men_n346_), .Y(men_men_n364_));
  INV        u348(.A(men_men_n311_), .Y(men_men_n365_));
  AOI210     u349(.A0(men_men_n365_), .A1(men_men_n18_), .B0(men_men_n152_), .Y(men_men_n366_));
  AO220      u350(.A0(men_men_n366_), .A1(men_men_n364_), .B0(men_men_n341_), .B1(men_men_n328_), .Y(men_men_n367_));
  NA2        u351(.A(men_men_n360_), .B(x6), .Y(men_men_n368_));
  AOI210     u352(.A0(x6), .A1(x1), .B0(men_men_n151_), .Y(men_men_n369_));
  NA2        u353(.A(men_men_n348_), .B(x0), .Y(men_men_n370_));
  NA2        u354(.A(men_men_n80_), .B(x6), .Y(men_men_n371_));
  OAI210     u355(.A0(men_men_n370_), .A1(men_men_n369_), .B0(men_men_n371_), .Y(men_men_n372_));
  NA2        u356(.A(men_men_n372_), .B(men_men_n368_), .Y(men_men_n373_));
  NA3        u357(.A(men_men_n373_), .B(men_men_n367_), .C(men_men_n317_), .Y(men_men_n374_));
  AOI210     u358(.A0(men_men_n200_), .A1(x8), .B0(men_men_n110_), .Y(men_men_n375_));
  INV        u359(.A(men_men_n375_), .Y(men_men_n376_));
  NA3        u360(.A(men_men_n376_), .B(men_men_n197_), .C(men_men_n152_), .Y(men_men_n377_));
  OAI210     u361(.A0(men_men_n27_), .A1(x1), .B0(men_men_n230_), .Y(men_men_n378_));
  AO220      u362(.A0(men_men_n378_), .A1(men_men_n149_), .B0(men_men_n109_), .B1(x4), .Y(men_men_n379_));
  NA3        u363(.A(x7), .B(x3), .C(x0), .Y(men_men_n380_));
  NA2        u364(.A(men_men_n221_), .B(x0), .Y(men_men_n381_));
  OAI220     u365(.A0(men_men_n381_), .A1(x2), .B0(men_men_n380_), .B1(men_men_n347_), .Y(men_men_n382_));
  AOI210     u366(.A0(men_men_n379_), .A1(men_men_n118_), .B0(men_men_n382_), .Y(men_men_n383_));
  AOI210     u367(.A0(men_men_n383_), .A1(men_men_n377_), .B0(men_men_n24_), .Y(men_men_n384_));
  OAI210     u368(.A0(men_men_n197_), .A1(men_men_n66_), .B0(men_men_n207_), .Y(men_men_n385_));
  NA3        u369(.A(men_men_n200_), .B(men_men_n223_), .C(x8), .Y(men_men_n386_));
  AOI210     u370(.A0(men_men_n386_), .A1(men_men_n385_), .B0(men_men_n24_), .Y(men_men_n387_));
  NA2        u371(.A(men_men_n387_), .B(men_men_n149_), .Y(men_men_n388_));
  NAi31      u372(.An(men_men_n48_), .B(men_men_n287_), .C(men_men_n177_), .Y(men_men_n389_));
  NA2        u373(.A(men_men_n389_), .B(men_men_n388_), .Y(men_men_n390_));
  OAI210     u374(.A0(men_men_n390_), .A1(men_men_n384_), .B0(x6), .Y(men_men_n391_));
  OAI210     u375(.A0(men_men_n163_), .A1(men_men_n46_), .B0(men_men_n135_), .Y(men_men_n392_));
  NA2        u376(.A(men_men_n53_), .B(men_men_n36_), .Y(men_men_n393_));
  AOI220     u377(.A0(men_men_n393_), .A1(men_men_n392_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n394_));
  NO2        u378(.A(men_men_n152_), .B(x0), .Y(men_men_n395_));
  AOI220     u379(.A0(men_men_n395_), .A1(men_men_n221_), .B0(men_men_n197_), .B1(men_men_n152_), .Y(men_men_n396_));
  INV        u380(.A(x1), .Y(men_men_n397_));
  OAI210     u381(.A0(men_men_n396_), .A1(x8), .B0(men_men_n397_), .Y(men_men_n398_));
  NO4        u382(.A(men_men_n126_), .B(men_men_n298_), .C(x9), .D(x2), .Y(men_men_n399_));
  NOi21      u383(.An(men_men_n124_), .B(men_men_n181_), .Y(men_men_n400_));
  NO3        u384(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n18_), .Y(men_men_n401_));
  NO3        u385(.A(x9), .B(men_men_n152_), .C(x0), .Y(men_men_n402_));
  AOI220     u386(.A0(men_men_n402_), .A1(men_men_n244_), .B0(men_men_n359_), .B1(men_men_n152_), .Y(men_men_n403_));
  NA3        u387(.A(men_men_n403_), .B(men_men_n401_), .C(men_men_n48_), .Y(men_men_n404_));
  OAI210     u388(.A0(men_men_n398_), .A1(men_men_n394_), .B0(men_men_n404_), .Y(men_men_n405_));
  NOi31      u389(.An(men_men_n395_), .B(men_men_n31_), .C(x8), .Y(men_men_n406_));
  AOI210     u390(.A0(men_men_n36_), .A1(x9), .B0(men_men_n133_), .Y(men_men_n407_));
  NO3        u391(.A(men_men_n407_), .B(men_men_n124_), .C(men_men_n41_), .Y(men_men_n408_));
  AOI210     u392(.A0(men_men_n266_), .A1(men_men_n58_), .B0(men_men_n123_), .Y(men_men_n409_));
  NO2        u393(.A(men_men_n409_), .B(x3), .Y(men_men_n410_));
  NO3        u394(.A(men_men_n410_), .B(men_men_n408_), .C(x2), .Y(men_men_n411_));
  OAI220     u395(.A0(men_men_n343_), .A1(men_men_n302_), .B0(men_men_n298_), .B1(men_men_n41_), .Y(men_men_n412_));
  INV        u396(.A(men_men_n380_), .Y(men_men_n413_));
  AOI220     u397(.A0(men_men_n413_), .A1(men_men_n90_), .B0(men_men_n412_), .B1(men_men_n152_), .Y(men_men_n414_));
  NO2        u398(.A(men_men_n414_), .B(men_men_n52_), .Y(men_men_n415_));
  NO3        u399(.A(men_men_n415_), .B(men_men_n411_), .C(men_men_n406_), .Y(men_men_n416_));
  AOI210     u400(.A0(men_men_n416_), .A1(men_men_n405_), .B0(men_men_n24_), .Y(men_men_n417_));
  NA4        u401(.A(men_men_n30_), .B(men_men_n90_), .C(x2), .D(men_men_n17_), .Y(men_men_n418_));
  NA2        u402(.A(men_men_n226_), .B(x7), .Y(men_men_n419_));
  NA3        u403(.A(men_men_n419_), .B(men_men_n151_), .C(men_men_n134_), .Y(men_men_n420_));
  NA2        u404(.A(men_men_n420_), .B(men_men_n418_), .Y(men_men_n421_));
  OAI210     u405(.A0(men_men_n421_), .A1(men_men_n417_), .B0(men_men_n34_), .Y(men_men_n422_));
  NO2        u406(.A(men_men_n402_), .B(men_men_n207_), .Y(men_men_n423_));
  NO4        u407(.A(men_men_n423_), .B(men_men_n75_), .C(x4), .D(men_men_n52_), .Y(men_men_n424_));
  NA2        u408(.A(men_men_n254_), .B(men_men_n21_), .Y(men_men_n425_));
  NO2        u409(.A(men_men_n160_), .B(men_men_n135_), .Y(men_men_n426_));
  NA2        u410(.A(men_men_n426_), .B(men_men_n425_), .Y(men_men_n427_));
  AOI210     u411(.A0(men_men_n427_), .A1(men_men_n167_), .B0(men_men_n27_), .Y(men_men_n428_));
  AOI220     u412(.A0(men_men_n355_), .A1(men_men_n90_), .B0(men_men_n150_), .B1(men_men_n200_), .Y(men_men_n429_));
  NA2        u413(.A(men_men_n429_), .B(men_men_n88_), .Y(men_men_n430_));
  NA2        u414(.A(men_men_n430_), .B(men_men_n177_), .Y(men_men_n431_));
  NO2        u415(.A(men_men_n160_), .B(men_men_n41_), .Y(men_men_n432_));
  NA2        u416(.A(x3), .B(men_men_n52_), .Y(men_men_n433_));
  AOI210     u417(.A0(men_men_n164_), .A1(men_men_n26_), .B0(men_men_n70_), .Y(men_men_n434_));
  OAI210     u418(.A0(men_men_n149_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n435_));
  NO2        u419(.A(x3), .B(men_men_n52_), .Y(men_men_n436_));
  AOI210     u420(.A0(men_men_n436_), .A1(men_men_n435_), .B0(men_men_n434_), .Y(men_men_n437_));
  OAI210     u421(.A0(men_men_n153_), .A1(men_men_n433_), .B0(men_men_n437_), .Y(men_men_n438_));
  AOI220     u422(.A0(men_men_n438_), .A1(x0), .B0(men_men_n432_), .B1(men_men_n135_), .Y(men_men_n439_));
  AOI210     u423(.A0(men_men_n439_), .A1(men_men_n431_), .B0(men_men_n234_), .Y(men_men_n440_));
  INV        u424(.A(x5), .Y(men_men_n441_));
  NO4        u425(.A(men_men_n105_), .B(men_men_n441_), .C(men_men_n58_), .D(men_men_n31_), .Y(men_men_n442_));
  NO4        u426(.A(men_men_n442_), .B(men_men_n440_), .C(men_men_n428_), .D(men_men_n424_), .Y(men_men_n443_));
  NA3        u427(.A(men_men_n443_), .B(men_men_n422_), .C(men_men_n391_), .Y(men_men_n444_));
  AOI210     u428(.A0(men_men_n374_), .A1(men_men_n24_), .B0(men_men_n444_), .Y(men05));
  INV        u429(.A(men_men_n176_), .Y(men_men_n448_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule