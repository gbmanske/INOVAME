// Benchmark "top" written by ABC on Thu Jun 20 14:00:11 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n125_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n997_, new_new_n998_, new_new_n999_,
    new_new_n1000_, new_new_n1001_, new_new_n1002_, new_new_n1003_,
    new_new_n1004_, new_new_n1005_, new_new_n1006_, new_new_n1007_,
    new_new_n1008_, new_new_n1009_, new_new_n1010_, new_new_n1011_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NO2        g018(.A(new_new_n36_), .B(i_3_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(men1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NO2        g031(.A(i_1_), .B(i_6_), .Y(new_new_n54_));
  NA2        g032(.A(i_8_), .B(i_7_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_12_), .Y(new_new_n56_));
  INV        g034(.A(i_1_), .Y(new_new_n57_));
  NA2        g035(.A(new_new_n57_), .B(i_6_), .Y(new_new_n58_));
  INV        g036(.A(new_new_n31_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(new_new_n56_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n50_), .B(i_2_), .Y(new_new_n61_));
  AOI210     g039(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_6_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(new_new_n25_), .Y(new_new_n64_));
  INV        g042(.A(i_0_), .Y(new_new_n65_));
  NAi21      g043(.An(i_5_), .B(i_10_), .Y(new_new_n66_));
  NA2        g044(.A(i_5_), .B(i_9_), .Y(new_new_n67_));
  AOI210     g045(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n65_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n64_), .Y(new_new_n69_));
  NA2        g047(.A(new_new_n61_), .B(new_new_n69_), .Y(new_new_n70_));
  OAI210     g048(.A0(new_new_n70_), .A1(new_new_n60_), .B0(i_0_), .Y(new_new_n71_));
  NA2        g049(.A(i_12_), .B(i_5_), .Y(new_new_n72_));
  NA2        g050(.A(i_2_), .B(i_8_), .Y(new_new_n73_));
  NO2        g051(.A(i_3_), .B(i_9_), .Y(new_new_n74_));
  NO2        g052(.A(i_3_), .B(i_7_), .Y(new_new_n75_));
  NO3        g053(.A(new_new_n75_), .B(new_new_n74_), .C(new_new_n57_), .Y(new_new_n76_));
  INV        g054(.A(i_6_), .Y(new_new_n77_));
  OR4        g055(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n78_));
  INV        g056(.A(new_new_n78_), .Y(new_new_n79_));
  NO2        g057(.A(i_2_), .B(i_7_), .Y(new_new_n80_));
  OAI210     g058(.A0(new_new_n76_), .A1(i_8_), .B0(new_new_n78_), .Y(new_new_n81_));
  NAi21      g059(.An(i_6_), .B(i_10_), .Y(new_new_n82_));
  NA2        g060(.A(i_6_), .B(i_9_), .Y(new_new_n83_));
  AOI210     g061(.A0(new_new_n83_), .A1(new_new_n82_), .B0(new_new_n57_), .Y(new_new_n84_));
  NA2        g062(.A(i_2_), .B(i_6_), .Y(new_new_n85_));
  NO3        g063(.A(new_new_n85_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n86_));
  NO2        g064(.A(new_new_n86_), .B(new_new_n84_), .Y(new_new_n87_));
  AOI210     g065(.A0(new_new_n87_), .A1(new_new_n81_), .B0(new_new_n72_), .Y(new_new_n88_));
  AN3        g066(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n89_));
  NAi21      g067(.An(i_6_), .B(i_11_), .Y(new_new_n90_));
  NO2        g068(.A(i_5_), .B(i_8_), .Y(new_new_n91_));
  NOi21      g069(.An(new_new_n91_), .B(new_new_n90_), .Y(new_new_n92_));
  AOI210     g070(.A0(new_new_n89_), .A1(new_new_n32_), .B0(new_new_n92_), .Y(new_new_n93_));
  INV        g071(.A(i_7_), .Y(new_new_n94_));
  NO2        g072(.A(i_0_), .B(i_5_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n95_), .B(new_new_n77_), .Y(new_new_n96_));
  NA2        g074(.A(i_12_), .B(i_3_), .Y(new_new_n97_));
  INV        g075(.A(new_new_n97_), .Y(new_new_n98_));
  NAi21      g076(.An(i_7_), .B(i_11_), .Y(new_new_n99_));
  NO3        g077(.A(new_new_n99_), .B(new_new_n82_), .C(new_new_n51_), .Y(new_new_n100_));
  AN2        g078(.A(i_2_), .B(i_10_), .Y(new_new_n101_));
  OR2        g079(.A(new_new_n72_), .B(new_new_n54_), .Y(new_new_n102_));
  NO2        g080(.A(i_8_), .B(new_new_n94_), .Y(new_new_n103_));
  NO3        g081(.A(new_new_n103_), .B(new_new_n102_), .C(new_new_n1008_), .Y(new_new_n104_));
  NA2        g082(.A(i_12_), .B(i_7_), .Y(new_new_n105_));
  NA2        g083(.A(i_11_), .B(i_12_), .Y(new_new_n106_));
  INV        g084(.A(new_new_n104_), .Y(new_new_n107_));
  NA3        g085(.A(new_new_n107_), .B(new_new_n97_), .C(new_new_n93_), .Y(new_new_n108_));
  NOi21      g086(.An(i_1_), .B(i_5_), .Y(new_new_n109_));
  NA2        g087(.A(new_new_n109_), .B(i_11_), .Y(new_new_n110_));
  NA2        g088(.A(new_new_n94_), .B(new_new_n37_), .Y(new_new_n111_));
  NA2        g089(.A(i_7_), .B(new_new_n25_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n112_), .B(new_new_n111_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n83_), .B(new_new_n82_), .Y(new_new_n114_));
  NAi21      g092(.An(i_3_), .B(i_8_), .Y(new_new_n115_));
  INV        g093(.A(new_new_n115_), .Y(new_new_n116_));
  NOi31      g094(.An(new_new_n116_), .B(new_new_n114_), .C(i_10_), .Y(new_new_n117_));
  NO2        g095(.A(i_1_), .B(new_new_n77_), .Y(new_new_n118_));
  NO2        g096(.A(i_6_), .B(i_5_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(i_3_), .Y(new_new_n120_));
  AO210      g098(.A0(new_new_n120_), .A1(new_new_n47_), .B0(new_new_n118_), .Y(new_new_n121_));
  OAI220     g099(.A0(new_new_n121_), .A1(new_new_n99_), .B0(new_new_n117_), .B1(new_new_n110_), .Y(new_new_n122_));
  NO3        g100(.A(new_new_n122_), .B(new_new_n108_), .C(new_new_n88_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n71_), .Y(men2));
  NO2        g102(.A(new_new_n57_), .B(new_new_n37_), .Y(new_new_n125_));
  NA3        g103(.A(new_new_n69_), .B(new_new_n61_), .C(new_new_n30_), .Y(men0));
  AN2        g104(.A(i_8_), .B(i_7_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(i_6_), .Y(new_new_n128_));
  NO2        g106(.A(i_12_), .B(i_13_), .Y(new_new_n129_));
  NAi21      g107(.An(i_5_), .B(i_11_), .Y(new_new_n130_));
  NOi21      g108(.An(new_new_n129_), .B(new_new_n130_), .Y(new_new_n131_));
  NO2        g109(.A(i_0_), .B(i_1_), .Y(new_new_n132_));
  NA2        g110(.A(i_2_), .B(i_3_), .Y(new_new_n133_));
  NO2        g111(.A(new_new_n133_), .B(i_4_), .Y(new_new_n134_));
  NA3        g112(.A(new_new_n134_), .B(new_new_n132_), .C(new_new_n131_), .Y(new_new_n135_));
  OR2        g113(.A(new_new_n135_), .B(new_new_n25_), .Y(new_new_n136_));
  AN2        g114(.A(new_new_n129_), .B(new_new_n74_), .Y(new_new_n137_));
  NO2        g115(.A(new_new_n137_), .B(new_new_n27_), .Y(new_new_n138_));
  NA2        g116(.A(i_1_), .B(i_5_), .Y(new_new_n139_));
  NO2        g117(.A(new_new_n65_), .B(new_new_n46_), .Y(new_new_n140_));
  NA2        g118(.A(new_new_n140_), .B(new_new_n36_), .Y(new_new_n141_));
  NO3        g119(.A(new_new_n141_), .B(new_new_n139_), .C(new_new_n138_), .Y(new_new_n142_));
  OR2        g120(.A(i_0_), .B(i_1_), .Y(new_new_n143_));
  NO3        g121(.A(new_new_n143_), .B(new_new_n72_), .C(i_13_), .Y(new_new_n144_));
  NAi32      g122(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n145_));
  NAi21      g123(.An(new_new_n145_), .B(new_new_n144_), .Y(new_new_n146_));
  NOi21      g124(.An(i_4_), .B(i_10_), .Y(new_new_n147_));
  NA2        g125(.A(new_new_n147_), .B(new_new_n39_), .Y(new_new_n148_));
  NO2        g126(.A(i_3_), .B(i_5_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n65_), .B(i_2_), .C(i_1_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n1011_), .B(new_new_n142_), .Y(new_new_n151_));
  AOI210     g129(.A0(new_new_n151_), .A1(new_new_n136_), .B0(new_new_n128_), .Y(new_new_n152_));
  NA3        g130(.A(new_new_n65_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n153_));
  NOi21      g131(.An(i_4_), .B(i_9_), .Y(new_new_n154_));
  NOi21      g132(.An(i_11_), .B(i_13_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n154_), .Y(new_new_n156_));
  NO2        g134(.A(i_4_), .B(i_5_), .Y(new_new_n157_));
  NAi21      g135(.An(i_12_), .B(i_11_), .Y(new_new_n158_));
  NO2        g136(.A(new_new_n158_), .B(i_13_), .Y(new_new_n159_));
  NA3        g137(.A(new_new_n159_), .B(new_new_n157_), .C(new_new_n74_), .Y(new_new_n160_));
  AOI210     g138(.A0(new_new_n160_), .A1(new_new_n156_), .B0(new_new_n153_), .Y(new_new_n161_));
  NO2        g139(.A(new_new_n65_), .B(new_new_n57_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n36_), .B(i_5_), .Y(new_new_n163_));
  NAi31      g141(.An(new_new_n163_), .B(new_new_n137_), .C(i_11_), .Y(new_new_n164_));
  NA2        g142(.A(i_3_), .B(i_5_), .Y(new_new_n165_));
  OR2        g143(.A(new_new_n165_), .B(new_new_n156_), .Y(new_new_n166_));
  AOI210     g144(.A0(new_new_n166_), .A1(new_new_n164_), .B0(i_2_), .Y(new_new_n167_));
  NO2        g145(.A(new_new_n65_), .B(i_5_), .Y(new_new_n168_));
  NO2        g146(.A(i_13_), .B(i_10_), .Y(new_new_n169_));
  NA3        g147(.A(new_new_n169_), .B(new_new_n168_), .C(new_new_n44_), .Y(new_new_n170_));
  NO2        g148(.A(i_2_), .B(i_1_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n171_), .B(i_3_), .Y(new_new_n172_));
  NAi21      g150(.An(i_4_), .B(i_12_), .Y(new_new_n173_));
  NO4        g151(.A(new_new_n173_), .B(new_new_n172_), .C(new_new_n170_), .D(new_new_n25_), .Y(new_new_n174_));
  NO3        g152(.A(new_new_n174_), .B(new_new_n167_), .C(new_new_n161_), .Y(new_new_n175_));
  INV        g153(.A(i_8_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n176_), .B(i_7_), .Y(new_new_n177_));
  NA2        g155(.A(new_new_n177_), .B(i_6_), .Y(new_new_n178_));
  NO3        g156(.A(i_3_), .B(new_new_n77_), .C(new_new_n48_), .Y(new_new_n179_));
  NA2        g157(.A(new_new_n179_), .B(new_new_n103_), .Y(new_new_n180_));
  NO3        g158(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n181_));
  NA3        g159(.A(new_new_n181_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n182_));
  NO3        g160(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n183_));
  OAI210     g161(.A0(new_new_n89_), .A1(i_12_), .B0(new_new_n183_), .Y(new_new_n184_));
  AOI210     g162(.A0(new_new_n184_), .A1(new_new_n182_), .B0(new_new_n180_), .Y(new_new_n185_));
  NO2        g163(.A(i_3_), .B(i_8_), .Y(new_new_n186_));
  NO3        g164(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n187_));
  NA3        g165(.A(new_new_n187_), .B(new_new_n186_), .C(new_new_n39_), .Y(new_new_n188_));
  NO2        g166(.A(i_13_), .B(i_9_), .Y(new_new_n189_));
  NAi21      g167(.An(i_12_), .B(i_3_), .Y(new_new_n190_));
  NO3        g168(.A(i_0_), .B(i_2_), .C(new_new_n57_), .Y(new_new_n191_));
  NA2        g169(.A(new_new_n191_), .B(i_10_), .Y(new_new_n192_));
  OAI220     g170(.A0(new_new_n192_), .A1(new_new_n190_), .B0(new_new_n95_), .B1(new_new_n188_), .Y(new_new_n193_));
  AOI210     g171(.A0(new_new_n193_), .A1(i_7_), .B0(new_new_n185_), .Y(new_new_n194_));
  OAI220     g172(.A0(new_new_n194_), .A1(i_4_), .B0(new_new_n178_), .B1(new_new_n175_), .Y(new_new_n195_));
  NAi21      g173(.An(i_12_), .B(i_7_), .Y(new_new_n196_));
  NA3        g174(.A(i_13_), .B(new_new_n176_), .C(i_10_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n197_), .B(new_new_n196_), .Y(new_new_n198_));
  NA2        g176(.A(i_0_), .B(i_5_), .Y(new_new_n199_));
  NA2        g177(.A(new_new_n199_), .B(new_new_n96_), .Y(new_new_n200_));
  OAI220     g178(.A0(new_new_n200_), .A1(new_new_n172_), .B0(i_2_), .B1(new_new_n120_), .Y(new_new_n201_));
  NAi31      g179(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n202_));
  NO2        g180(.A(new_new_n36_), .B(i_13_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n46_), .B(new_new_n57_), .Y(new_new_n204_));
  NA3        g182(.A(new_new_n204_), .B(i_3_), .C(new_new_n203_), .Y(new_new_n205_));
  INV        g183(.A(i_13_), .Y(new_new_n206_));
  NO2        g184(.A(i_12_), .B(new_new_n206_), .Y(new_new_n207_));
  NA3        g185(.A(new_new_n207_), .B(new_new_n181_), .C(new_new_n179_), .Y(new_new_n208_));
  OAI210     g186(.A0(new_new_n205_), .A1(new_new_n202_), .B0(new_new_n208_), .Y(new_new_n209_));
  AOI220     g187(.A0(new_new_n209_), .A1(new_new_n127_), .B0(new_new_n201_), .B1(new_new_n198_), .Y(new_new_n210_));
  NO2        g188(.A(i_12_), .B(new_new_n37_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n165_), .B(i_4_), .Y(new_new_n212_));
  NA2        g190(.A(new_new_n212_), .B(new_new_n211_), .Y(new_new_n213_));
  OR2        g191(.A(i_8_), .B(i_7_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n214_), .B(new_new_n77_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n51_), .B(i_1_), .Y(new_new_n216_));
  NA2        g194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  INV        g195(.A(i_12_), .Y(new_new_n218_));
  NO3        g196(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n219_));
  NA2        g197(.A(i_2_), .B(i_1_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n217_), .B(new_new_n213_), .Y(new_new_n221_));
  NO3        g199(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n222_));
  NAi21      g200(.An(i_4_), .B(i_3_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n223_), .B(new_new_n67_), .Y(new_new_n224_));
  NO2        g202(.A(i_0_), .B(i_6_), .Y(new_new_n225_));
  NOi41      g203(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n226_));
  NA2        g204(.A(new_new_n226_), .B(new_new_n225_), .Y(new_new_n227_));
  NA2        g205(.A(new_new_n221_), .B(new_new_n189_), .Y(new_new_n228_));
  NO2        g206(.A(i_11_), .B(new_new_n206_), .Y(new_new_n229_));
  NOi21      g207(.An(i_1_), .B(i_6_), .Y(new_new_n230_));
  NAi21      g208(.An(i_3_), .B(i_7_), .Y(new_new_n231_));
  NA2        g209(.A(new_new_n218_), .B(i_9_), .Y(new_new_n232_));
  OR4        g210(.A(new_new_n232_), .B(new_new_n231_), .C(new_new_n230_), .D(new_new_n168_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n234_));
  NO2        g212(.A(i_12_), .B(i_3_), .Y(new_new_n235_));
  NA2        g213(.A(i_3_), .B(i_9_), .Y(new_new_n236_));
  NAi21      g214(.An(i_7_), .B(i_10_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  NA3        g216(.A(new_new_n238_), .B(new_new_n1010_), .C(new_new_n58_), .Y(new_new_n239_));
  NA2        g217(.A(new_new_n239_), .B(new_new_n233_), .Y(new_new_n240_));
  NA3        g218(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n218_), .B(i_13_), .Y(new_new_n242_));
  NO2        g220(.A(new_new_n242_), .B(new_new_n67_), .Y(new_new_n243_));
  AOI220     g221(.A0(new_new_n243_), .A1(new_new_n127_), .B0(new_new_n240_), .B1(new_new_n229_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n214_), .B(new_new_n37_), .Y(new_new_n245_));
  NA2        g223(.A(i_12_), .B(i_6_), .Y(new_new_n246_));
  NO3        g224(.A(i_9_), .B(new_new_n246_), .C(new_new_n48_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n223_), .B(i_2_), .Y(new_new_n248_));
  NA3        g226(.A(new_new_n248_), .B(new_new_n247_), .C(new_new_n44_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n229_), .B(i_9_), .Y(new_new_n250_));
  OAI210     g228(.A0(new_new_n65_), .A1(new_new_n250_), .B0(new_new_n249_), .Y(new_new_n251_));
  NO3        g229(.A(i_11_), .B(new_new_n206_), .C(new_new_n25_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n231_), .B(i_8_), .Y(new_new_n253_));
  NO2        g231(.A(i_6_), .B(new_new_n48_), .Y(new_new_n254_));
  NA3        g232(.A(new_new_n254_), .B(new_new_n253_), .C(new_new_n252_), .Y(new_new_n255_));
  NO3        g233(.A(new_new_n26_), .B(new_new_n77_), .C(i_5_), .Y(new_new_n256_));
  NA3        g234(.A(new_new_n256_), .B(new_new_n245_), .C(new_new_n207_), .Y(new_new_n257_));
  AOI210     g235(.A0(new_new_n257_), .A1(new_new_n255_), .B0(new_new_n46_), .Y(new_new_n258_));
  AOI210     g236(.A0(new_new_n251_), .A1(new_new_n245_), .B0(new_new_n258_), .Y(new_new_n259_));
  NA4        g237(.A(new_new_n259_), .B(new_new_n244_), .C(new_new_n228_), .D(new_new_n210_), .Y(new_new_n260_));
  NO3        g238(.A(i_12_), .B(new_new_n206_), .C(new_new_n37_), .Y(new_new_n261_));
  INV        g239(.A(new_new_n261_), .Y(new_new_n262_));
  INV        g240(.A(i_8_), .Y(new_new_n263_));
  NOi21      g241(.An(new_new_n149_), .B(new_new_n77_), .Y(new_new_n264_));
  NO3        g242(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n265_));
  AOI220     g243(.A0(new_new_n265_), .A1(new_new_n179_), .B0(new_new_n264_), .B1(new_new_n216_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n266_), .B(new_new_n263_), .Y(new_new_n267_));
  NO2        g245(.A(new_new_n220_), .B(i_0_), .Y(new_new_n268_));
  AOI220     g246(.A0(new_new_n268_), .A1(new_new_n177_), .B0(i_1_), .B1(new_new_n127_), .Y(new_new_n269_));
  NA2        g247(.A(new_new_n254_), .B(new_new_n26_), .Y(new_new_n270_));
  NO2        g248(.A(new_new_n270_), .B(new_new_n269_), .Y(new_new_n271_));
  NA2        g249(.A(i_0_), .B(i_1_), .Y(new_new_n272_));
  NO2        g250(.A(new_new_n272_), .B(i_2_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n55_), .B(i_6_), .Y(new_new_n274_));
  NA3        g252(.A(new_new_n274_), .B(new_new_n273_), .C(new_new_n149_), .Y(new_new_n275_));
  OAI210     g253(.A0(i_3_), .A1(new_new_n128_), .B0(new_new_n275_), .Y(new_new_n276_));
  NO3        g254(.A(new_new_n276_), .B(new_new_n271_), .C(new_new_n267_), .Y(new_new_n277_));
  NO2        g255(.A(i_3_), .B(i_10_), .Y(new_new_n278_));
  NA3        g256(.A(new_new_n278_), .B(new_new_n39_), .C(new_new_n44_), .Y(new_new_n279_));
  NO2        g257(.A(i_2_), .B(new_new_n94_), .Y(new_new_n280_));
  NA2        g258(.A(i_1_), .B(new_new_n36_), .Y(new_new_n281_));
  NOi21      g259(.An(new_new_n199_), .B(new_new_n95_), .Y(new_new_n282_));
  NA3        g260(.A(new_new_n282_), .B(i_1_), .C(new_new_n280_), .Y(new_new_n283_));
  AN2        g261(.A(i_3_), .B(i_10_), .Y(new_new_n284_));
  NA4        g262(.A(new_new_n284_), .B(new_new_n181_), .C(new_new_n159_), .D(new_new_n157_), .Y(new_new_n285_));
  NO2        g263(.A(i_5_), .B(new_new_n37_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n287_));
  OR2        g265(.A(new_new_n283_), .B(new_new_n279_), .Y(new_new_n288_));
  OAI220     g266(.A0(new_new_n288_), .A1(i_6_), .B0(new_new_n277_), .B1(new_new_n262_), .Y(new_new_n289_));
  NO4        g267(.A(new_new_n289_), .B(new_new_n260_), .C(new_new_n195_), .D(new_new_n152_), .Y(new_new_n290_));
  NO3        g268(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n55_), .B(new_new_n77_), .Y(new_new_n292_));
  NA2        g270(.A(new_new_n268_), .B(new_new_n292_), .Y(new_new_n293_));
  NO3        g271(.A(i_6_), .B(new_new_n176_), .C(i_7_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n294_), .B(new_new_n181_), .Y(new_new_n295_));
  AOI210     g273(.A0(new_new_n295_), .A1(new_new_n293_), .B0(i_5_), .Y(new_new_n296_));
  NO2        g274(.A(i_2_), .B(i_3_), .Y(new_new_n297_));
  OR2        g275(.A(i_0_), .B(i_5_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n199_), .B(new_new_n298_), .Y(new_new_n299_));
  NA4        g277(.A(new_new_n299_), .B(new_new_n215_), .C(new_new_n297_), .D(i_1_), .Y(new_new_n300_));
  NA3        g278(.A(new_new_n268_), .B(new_new_n264_), .C(new_new_n103_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n143_), .B(new_new_n46_), .Y(new_new_n302_));
  NA3        g280(.A(new_new_n302_), .B(i_7_), .C(new_new_n149_), .Y(new_new_n303_));
  NA3        g281(.A(new_new_n303_), .B(new_new_n301_), .C(new_new_n300_), .Y(new_new_n304_));
  OAI210     g282(.A0(new_new_n304_), .A1(new_new_n296_), .B0(i_4_), .Y(new_new_n305_));
  NO2        g283(.A(i_12_), .B(i_10_), .Y(new_new_n306_));
  NOi21      g284(.An(i_5_), .B(i_0_), .Y(new_new_n307_));
  AOI210     g285(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n94_), .Y(new_new_n308_));
  NO3        g286(.A(new_new_n308_), .B(new_new_n281_), .C(new_new_n115_), .Y(new_new_n309_));
  NA4        g287(.A(new_new_n75_), .B(new_new_n36_), .C(new_new_n77_), .D(i_8_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n309_), .B(new_new_n306_), .Y(new_new_n311_));
  NO2        g289(.A(i_6_), .B(i_8_), .Y(new_new_n312_));
  NOi21      g290(.An(i_0_), .B(i_2_), .Y(new_new_n313_));
  AN2        g291(.A(new_new_n313_), .B(new_new_n312_), .Y(new_new_n314_));
  NO2        g292(.A(i_1_), .B(i_7_), .Y(new_new_n315_));
  NA3        g293(.A(new_new_n312_), .B(new_new_n41_), .C(i_5_), .Y(new_new_n316_));
  NA3        g294(.A(new_new_n316_), .B(new_new_n311_), .C(new_new_n305_), .Y(new_new_n317_));
  INV        g295(.A(i_8_), .Y(new_new_n318_));
  NOi21      g296(.An(new_new_n139_), .B(new_new_n96_), .Y(new_new_n319_));
  NA2        g297(.A(new_new_n318_), .B(i_3_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n272_), .B(new_new_n73_), .Y(new_new_n321_));
  NA2        g299(.A(new_new_n321_), .B(new_new_n119_), .Y(new_new_n322_));
  NO2        g300(.A(new_new_n85_), .B(new_new_n176_), .Y(new_new_n323_));
  NA3        g301(.A(new_new_n282_), .B(new_new_n323_), .C(new_new_n57_), .Y(new_new_n324_));
  AOI210     g302(.A0(new_new_n324_), .A1(new_new_n322_), .B0(i_3_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n176_), .B(i_9_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n326_), .B(i_1_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n325_), .B(new_new_n271_), .Y(new_new_n328_));
  AOI210     g306(.A0(new_new_n328_), .A1(new_new_n320_), .B0(new_new_n148_), .Y(new_new_n329_));
  AOI210     g307(.A0(new_new_n317_), .A1(new_new_n291_), .B0(new_new_n329_), .Y(new_new_n330_));
  NOi32      g308(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n331_));
  INV        g309(.A(new_new_n331_), .Y(new_new_n332_));
  NAi21      g310(.An(i_1_), .B(i_5_), .Y(new_new_n333_));
  NA2        g311(.A(new_new_n333_), .B(i_0_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(new_new_n25_), .Y(new_new_n335_));
  OAI210     g313(.A0(new_new_n335_), .A1(new_new_n145_), .B0(new_new_n227_), .Y(new_new_n336_));
  NAi41      g314(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n337_));
  OAI220     g315(.A0(new_new_n337_), .A1(new_new_n333_), .B0(new_new_n202_), .B1(new_new_n145_), .Y(new_new_n338_));
  AOI210     g316(.A0(new_new_n337_), .A1(new_new_n145_), .B0(new_new_n143_), .Y(new_new_n339_));
  NOi32      g317(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n340_), .B(new_new_n46_), .Y(new_new_n341_));
  NO2        g319(.A(new_new_n341_), .B(i_0_), .Y(new_new_n342_));
  OR3        g320(.A(new_new_n342_), .B(new_new_n339_), .C(new_new_n338_), .Y(new_new_n343_));
  NO2        g321(.A(i_1_), .B(new_new_n94_), .Y(new_new_n344_));
  NAi21      g322(.An(i_3_), .B(i_4_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n345_), .B(i_9_), .Y(new_new_n346_));
  AN2        g324(.A(i_6_), .B(i_7_), .Y(new_new_n347_));
  OAI210     g325(.A0(new_new_n347_), .A1(new_new_n344_), .B0(new_new_n346_), .Y(new_new_n348_));
  NA2        g326(.A(i_2_), .B(i_7_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n345_), .B(i_10_), .Y(new_new_n350_));
  NA3        g328(.A(new_new_n350_), .B(new_new_n349_), .C(new_new_n225_), .Y(new_new_n351_));
  AOI210     g329(.A0(new_new_n351_), .A1(new_new_n348_), .B0(new_new_n168_), .Y(new_new_n352_));
  AOI220     g330(.A0(new_new_n350_), .A1(new_new_n315_), .B0(new_new_n219_), .B1(new_new_n171_), .Y(new_new_n353_));
  NO3        g331(.A(new_new_n352_), .B(new_new_n343_), .C(new_new_n336_), .Y(new_new_n354_));
  NO2        g332(.A(new_new_n354_), .B(new_new_n332_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n55_), .B(new_new_n25_), .Y(new_new_n356_));
  AN2        g334(.A(i_12_), .B(i_5_), .Y(new_new_n357_));
  NO2        g335(.A(i_4_), .B(new_new_n26_), .Y(new_new_n358_));
  NO2        g336(.A(i_11_), .B(i_6_), .Y(new_new_n359_));
  NA3        g337(.A(new_new_n359_), .B(new_new_n302_), .C(new_new_n206_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n360_), .B(new_new_n1007_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n223_), .B(i_5_), .Y(new_new_n362_));
  NO2        g340(.A(i_5_), .B(i_10_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n129_), .B(new_new_n45_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n364_), .B(new_new_n223_), .Y(new_new_n365_));
  OAI210     g343(.A0(new_new_n365_), .A1(new_new_n361_), .B0(new_new_n356_), .Y(new_new_n366_));
  NO2        g344(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n367_));
  INV        g345(.A(new_new_n135_), .Y(new_new_n368_));
  OAI210     g346(.A0(new_new_n368_), .A1(new_new_n361_), .B0(new_new_n367_), .Y(new_new_n369_));
  NO3        g347(.A(new_new_n77_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n370_));
  NO2        g348(.A(i_3_), .B(new_new_n94_), .Y(new_new_n371_));
  NO2        g349(.A(i_11_), .B(i_12_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n363_), .B(new_new_n218_), .Y(new_new_n373_));
  NA3        g351(.A(new_new_n103_), .B(new_new_n41_), .C(i_11_), .Y(new_new_n374_));
  OAI220     g352(.A0(new_new_n374_), .A1(new_new_n202_), .B0(new_new_n373_), .B1(new_new_n310_), .Y(new_new_n375_));
  NAi21      g353(.An(i_13_), .B(i_0_), .Y(new_new_n376_));
  INV        g354(.A(new_new_n375_), .Y(new_new_n377_));
  NA3        g355(.A(new_new_n377_), .B(new_new_n369_), .C(new_new_n366_), .Y(new_new_n378_));
  NO3        g356(.A(i_1_), .B(i_12_), .C(new_new_n77_), .Y(new_new_n379_));
  NO2        g357(.A(i_0_), .B(i_11_), .Y(new_new_n380_));
  INV        g358(.A(i_5_), .Y(new_new_n381_));
  NOi21      g359(.An(i_2_), .B(i_12_), .Y(new_new_n382_));
  NO2        g360(.A(i_12_), .B(new_new_n381_), .Y(new_new_n383_));
  NA2        g361(.A(new_new_n127_), .B(i_9_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n384_), .B(i_4_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n383_), .B(new_new_n385_), .Y(new_new_n386_));
  NAi21      g364(.An(i_9_), .B(i_4_), .Y(new_new_n387_));
  OR2        g365(.A(i_13_), .B(i_10_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n156_), .B(new_new_n111_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n94_), .B(new_new_n25_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n261_), .B(new_new_n390_), .Y(new_new_n391_));
  INV        g369(.A(new_new_n191_), .Y(new_new_n392_));
  OAI220     g370(.A0(new_new_n392_), .A1(new_new_n196_), .B0(new_new_n391_), .B1(new_new_n319_), .Y(new_new_n393_));
  INV        g371(.A(new_new_n393_), .Y(new_new_n394_));
  AOI210     g372(.A0(new_new_n394_), .A1(new_new_n386_), .B0(new_new_n26_), .Y(new_new_n395_));
  NA2        g373(.A(new_new_n301_), .B(new_new_n300_), .Y(new_new_n396_));
  AOI220     g374(.A0(new_new_n274_), .A1(new_new_n265_), .B0(new_new_n268_), .B1(new_new_n292_), .Y(new_new_n397_));
  NO2        g375(.A(new_new_n165_), .B(new_new_n77_), .Y(new_new_n398_));
  AOI220     g376(.A0(new_new_n398_), .A1(new_new_n273_), .B0(new_new_n256_), .B1(new_new_n191_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(new_new_n263_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n400_), .B(new_new_n396_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n179_), .B(new_new_n89_), .Y(new_new_n402_));
  NA3        g380(.A(new_new_n302_), .B(new_new_n149_), .C(new_new_n77_), .Y(new_new_n403_));
  AOI210     g381(.A0(new_new_n403_), .A1(new_new_n402_), .B0(i_8_), .Y(new_new_n404_));
  NA3        g382(.A(new_new_n1010_), .B(new_new_n58_), .C(i_2_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n274_), .B(new_new_n216_), .Y(new_new_n406_));
  OAI220     g384(.A0(new_new_n406_), .A1(new_new_n165_), .B0(new_new_n405_), .B1(new_new_n1004_), .Y(new_new_n407_));
  NO2        g385(.A(i_3_), .B(new_new_n48_), .Y(new_new_n408_));
  NA3        g386(.A(new_new_n315_), .B(new_new_n314_), .C(new_new_n408_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n294_), .B(new_new_n299_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n410_), .B(new_new_n409_), .Y(new_new_n411_));
  NO3        g389(.A(new_new_n411_), .B(new_new_n407_), .C(new_new_n404_), .Y(new_new_n412_));
  AOI210     g390(.A0(new_new_n412_), .A1(new_new_n401_), .B0(new_new_n250_), .Y(new_new_n413_));
  NO4        g391(.A(new_new_n413_), .B(new_new_n395_), .C(new_new_n378_), .D(new_new_n355_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n57_), .B(i_4_), .Y(new_new_n415_));
  NO2        g393(.A(new_new_n65_), .B(i_13_), .Y(new_new_n416_));
  NA3        g394(.A(new_new_n416_), .B(new_new_n415_), .C(i_2_), .Y(new_new_n417_));
  NO2        g395(.A(i_10_), .B(i_9_), .Y(new_new_n418_));
  NAi21      g396(.An(i_12_), .B(i_8_), .Y(new_new_n419_));
  NO2        g397(.A(new_new_n419_), .B(i_3_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n420_), .B(new_new_n418_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n1002_), .B(new_new_n96_), .Y(new_new_n422_));
  OAI220     g400(.A0(new_new_n422_), .A1(new_new_n188_), .B0(new_new_n421_), .B1(new_new_n417_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n287_), .B(i_0_), .Y(new_new_n424_));
  NO3        g402(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n425_));
  NA2        g403(.A(new_new_n246_), .B(new_new_n90_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n426_), .B(new_new_n425_), .Y(new_new_n427_));
  NA2        g405(.A(i_8_), .B(i_9_), .Y(new_new_n428_));
  NO2        g406(.A(new_new_n427_), .B(new_new_n424_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n229_), .B(new_new_n286_), .Y(new_new_n430_));
  NO3        g408(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n431_));
  AOI210     g409(.A0(new_new_n235_), .A1(new_new_n171_), .B0(new_new_n431_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n432_), .B(new_new_n430_), .Y(new_new_n433_));
  NO3        g411(.A(new_new_n433_), .B(new_new_n429_), .C(new_new_n423_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n273_), .B(new_new_n99_), .Y(new_new_n435_));
  OA220      g413(.A0(new_new_n327_), .A1(new_new_n148_), .B0(new_new_n435_), .B1(new_new_n213_), .Y(new_new_n436_));
  NA2        g414(.A(new_new_n89_), .B(i_13_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n398_), .B(new_new_n356_), .Y(new_new_n438_));
  NO2        g416(.A(i_2_), .B(i_13_), .Y(new_new_n439_));
  NA3        g417(.A(new_new_n439_), .B(new_new_n147_), .C(new_new_n92_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n438_), .B(new_new_n437_), .Y(new_new_n441_));
  NO3        g419(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n442_));
  NO2        g420(.A(i_6_), .B(i_7_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n443_), .B(new_new_n442_), .Y(new_new_n444_));
  OR2        g422(.A(i_11_), .B(i_8_), .Y(new_new_n445_));
  NOi21      g423(.An(i_2_), .B(i_7_), .Y(new_new_n446_));
  NAi31      g424(.An(new_new_n445_), .B(new_new_n446_), .C(new_new_n999_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n388_), .B(i_6_), .Y(new_new_n448_));
  NA3        g426(.A(new_new_n448_), .B(new_new_n415_), .C(new_new_n67_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n449_), .B(new_new_n447_), .Y(new_new_n450_));
  NO2        g428(.A(i_3_), .B(new_new_n176_), .Y(new_new_n451_));
  NO2        g429(.A(i_6_), .B(i_10_), .Y(new_new_n452_));
  NA4        g430(.A(new_new_n452_), .B(new_new_n291_), .C(new_new_n451_), .D(new_new_n218_), .Y(new_new_n453_));
  NO2        g431(.A(new_new_n453_), .B(new_new_n141_), .Y(new_new_n454_));
  NA3        g432(.A(new_new_n226_), .B(new_new_n155_), .C(new_new_n119_), .Y(new_new_n455_));
  NO2        g433(.A(new_new_n143_), .B(i_3_), .Y(new_new_n456_));
  NA3        g434(.A(new_new_n367_), .B(new_new_n162_), .C(new_new_n134_), .Y(new_new_n457_));
  NA2        g435(.A(new_new_n457_), .B(new_new_n455_), .Y(new_new_n458_));
  NO4        g436(.A(new_new_n458_), .B(new_new_n454_), .C(new_new_n450_), .D(new_new_n441_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n425_), .B(new_new_n357_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n431_), .B(new_new_n363_), .Y(new_new_n461_));
  NO2        g439(.A(new_new_n461_), .B(new_new_n205_), .Y(new_new_n462_));
  NAi21      g440(.An(new_new_n197_), .B(new_new_n372_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n26_), .B(i_5_), .Y(new_new_n464_));
  NA3        g442(.A(new_new_n1001_), .B(new_new_n464_), .C(new_new_n127_), .Y(new_new_n465_));
  NO2        g443(.A(new_new_n38_), .B(new_new_n465_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n27_), .B(i_10_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n291_), .B(new_new_n219_), .Y(new_new_n468_));
  OAI220     g446(.A0(new_new_n468_), .A1(new_new_n405_), .B0(new_new_n467_), .B1(new_new_n437_), .Y(new_new_n469_));
  NA4        g447(.A(new_new_n284_), .B(new_new_n204_), .C(new_new_n65_), .D(new_new_n218_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n470_), .B(new_new_n444_), .Y(new_new_n471_));
  NO4        g449(.A(new_new_n471_), .B(new_new_n469_), .C(new_new_n466_), .D(new_new_n462_), .Y(new_new_n472_));
  NA4        g450(.A(new_new_n472_), .B(new_new_n459_), .C(new_new_n436_), .D(new_new_n434_), .Y(new_new_n473_));
  NA3        g451(.A(new_new_n284_), .B(new_new_n159_), .C(new_new_n157_), .Y(new_new_n474_));
  OAI210     g452(.A0(new_new_n279_), .A1(new_new_n163_), .B0(new_new_n474_), .Y(new_new_n475_));
  AN2        g453(.A(new_new_n265_), .B(new_new_n215_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n476_), .B(new_new_n475_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n291_), .B(new_new_n150_), .Y(new_new_n478_));
  OAI210     g456(.A0(new_new_n478_), .A1(new_new_n213_), .B0(new_new_n285_), .Y(new_new_n479_));
  INV        g457(.A(new_new_n479_), .Y(new_new_n480_));
  NA4        g458(.A(new_new_n416_), .B(new_new_n415_), .C(new_new_n186_), .D(i_2_), .Y(new_new_n481_));
  INV        g459(.A(new_new_n481_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n357_), .B(new_new_n206_), .Y(new_new_n483_));
  NA2        g461(.A(new_new_n331_), .B(new_new_n65_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n347_), .B(new_new_n340_), .Y(new_new_n485_));
  AO210      g463(.A0(new_new_n484_), .A1(new_new_n483_), .B0(new_new_n485_), .Y(new_new_n486_));
  NO2        g464(.A(new_new_n36_), .B(i_8_), .Y(new_new_n487_));
  INV        g465(.A(new_new_n486_), .Y(new_new_n488_));
  AOI210     g466(.A0(new_new_n482_), .A1(new_new_n187_), .B0(new_new_n488_), .Y(new_new_n489_));
  OAI210     g467(.A0(i_8_), .A1(new_new_n57_), .B0(new_new_n121_), .Y(new_new_n490_));
  AOI210     g468(.A0(new_new_n177_), .A1(i_9_), .B0(new_new_n245_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n491_), .B(new_new_n182_), .Y(new_new_n492_));
  AOI220     g470(.A0(i_6_), .A1(new_new_n492_), .B0(new_new_n490_), .B1(new_new_n389_), .Y(new_new_n493_));
  NA4        g471(.A(new_new_n493_), .B(new_new_n489_), .C(new_new_n480_), .D(new_new_n477_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n362_), .B(new_new_n273_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n153_), .B(new_new_n495_), .Y(new_new_n496_));
  NO2        g474(.A(i_12_), .B(new_new_n176_), .Y(new_new_n497_));
  NA2        g475(.A(new_new_n497_), .B(new_new_n206_), .Y(new_new_n498_));
  NO3        g476(.A(i_6_), .B(new_new_n498_), .C(new_new_n435_), .Y(new_new_n499_));
  NOi21      g477(.An(new_new_n294_), .B(new_new_n38_), .Y(new_new_n500_));
  OAI210     g478(.A0(new_new_n500_), .A1(new_new_n499_), .B0(new_new_n496_), .Y(new_new_n501_));
  NO2        g479(.A(i_8_), .B(i_7_), .Y(new_new_n502_));
  OAI210     g480(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n503_), .B(new_new_n204_), .Y(new_new_n504_));
  AOI220     g482(.A0(new_new_n302_), .A1(new_new_n39_), .B0(new_new_n216_), .B1(new_new_n189_), .Y(new_new_n505_));
  OAI220     g483(.A0(new_new_n505_), .A1(new_new_n165_), .B0(new_new_n504_), .B1(new_new_n223_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n44_), .B(i_10_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(i_6_), .Y(new_new_n508_));
  NA3        g486(.A(new_new_n508_), .B(new_new_n506_), .C(new_new_n502_), .Y(new_new_n509_));
  AOI220     g487(.A0(new_new_n398_), .A1(new_new_n302_), .B0(i_2_), .B1(new_new_n225_), .Y(new_new_n510_));
  OAI220     g488(.A0(new_new_n510_), .A1(new_new_n242_), .B0(new_new_n437_), .B1(new_new_n120_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n511_), .B(new_new_n245_), .Y(new_new_n512_));
  NOi21      g490(.An(new_new_n268_), .B(new_new_n279_), .Y(new_new_n513_));
  NA3        g491(.A(new_new_n284_), .B(new_new_n157_), .C(new_new_n89_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n203_), .B(new_new_n44_), .Y(new_new_n515_));
  NO2        g493(.A(new_new_n143_), .B(i_5_), .Y(new_new_n516_));
  NA2        g494(.A(new_new_n516_), .B(new_new_n297_), .Y(new_new_n517_));
  OAI210     g495(.A0(new_new_n517_), .A1(new_new_n515_), .B0(new_new_n514_), .Y(new_new_n518_));
  OAI210     g496(.A0(new_new_n518_), .A1(new_new_n513_), .B0(new_new_n431_), .Y(new_new_n519_));
  NA4        g497(.A(new_new_n519_), .B(new_new_n512_), .C(new_new_n509_), .D(new_new_n501_), .Y(new_new_n520_));
  NA3        g498(.A(new_new_n199_), .B(new_new_n63_), .C(new_new_n44_), .Y(new_new_n521_));
  NA2        g499(.A(new_new_n261_), .B(new_new_n75_), .Y(new_new_n522_));
  AOI210     g500(.A0(new_new_n521_), .A1(new_new_n322_), .B0(new_new_n522_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n274_), .B(new_new_n265_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n524_), .B(new_new_n156_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n204_), .B(i_3_), .Y(new_new_n526_));
  NA2        g504(.A(new_new_n418_), .B(new_new_n203_), .Y(new_new_n527_));
  NO2        g505(.A(new_new_n526_), .B(new_new_n527_), .Y(new_new_n528_));
  NA2        g506(.A(i_0_), .B(new_new_n48_), .Y(new_new_n529_));
  NA3        g507(.A(new_new_n497_), .B(new_new_n252_), .C(new_new_n529_), .Y(new_new_n530_));
  NO2        g508(.A(i_2_), .B(new_new_n530_), .Y(new_new_n531_));
  NO4        g509(.A(new_new_n531_), .B(new_new_n528_), .C(new_new_n525_), .D(new_new_n523_), .Y(new_new_n532_));
  NO4        g510(.A(new_new_n230_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n533_));
  NO3        g511(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n214_), .B(new_new_n36_), .Y(new_new_n535_));
  AN2        g513(.A(new_new_n535_), .B(new_new_n534_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n388_), .B(i_1_), .Y(new_new_n537_));
  NOi31      g515(.An(new_new_n537_), .B(new_new_n426_), .C(new_new_n65_), .Y(new_new_n538_));
  AN4        g516(.A(new_new_n538_), .B(new_new_n385_), .C(new_new_n464_), .D(i_2_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n397_), .B(new_new_n160_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n540_), .B(new_new_n539_), .Y(new_new_n541_));
  NOi21      g519(.An(i_10_), .B(i_6_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n77_), .B(new_new_n25_), .Y(new_new_n543_));
  NA2        g521(.A(new_new_n261_), .B(new_new_n543_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n544_), .B(new_new_n424_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n105_), .B(new_new_n23_), .Y(new_new_n546_));
  NA2        g524(.A(new_new_n294_), .B(new_new_n150_), .Y(new_new_n547_));
  AOI220     g525(.A0(new_new_n547_), .A1(new_new_n406_), .B0(new_new_n166_), .B1(new_new_n164_), .Y(new_new_n548_));
  NOi21      g526(.An(new_new_n131_), .B(new_new_n310_), .Y(new_new_n549_));
  NO3        g527(.A(new_new_n549_), .B(new_new_n548_), .C(new_new_n545_), .Y(new_new_n550_));
  NO2        g528(.A(new_new_n484_), .B(new_new_n353_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n297_), .Y(new_new_n552_));
  NO2        g530(.A(i_12_), .B(new_new_n77_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n553_), .B(new_new_n252_), .Y(new_new_n554_));
  NA3        g532(.A(new_new_n359_), .B(new_new_n261_), .C(new_new_n199_), .Y(new_new_n555_));
  AOI210     g533(.A0(new_new_n555_), .A1(new_new_n554_), .B0(new_new_n552_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n157_), .B(i_0_), .Y(new_new_n557_));
  NO3        g535(.A(new_new_n557_), .B(i_8_), .C(new_new_n279_), .Y(new_new_n558_));
  OR2        g536(.A(i_2_), .B(i_5_), .Y(new_new_n559_));
  AOI210     g537(.A0(new_new_n349_), .A1(new_new_n225_), .B0(new_new_n181_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n560_), .B(new_new_n463_), .Y(new_new_n561_));
  NO4        g539(.A(new_new_n561_), .B(new_new_n558_), .C(new_new_n556_), .D(new_new_n551_), .Y(new_new_n562_));
  NA4        g540(.A(new_new_n562_), .B(new_new_n550_), .C(new_new_n541_), .D(new_new_n532_), .Y(new_new_n563_));
  NO4        g541(.A(new_new_n563_), .B(new_new_n520_), .C(new_new_n494_), .D(new_new_n473_), .Y(new_new_n564_));
  NA4        g542(.A(new_new_n564_), .B(new_new_n414_), .C(new_new_n330_), .D(new_new_n290_), .Y(men7));
  NO2        g543(.A(new_new_n99_), .B(new_new_n82_), .Y(new_new_n566_));
  NA2        g544(.A(new_new_n358_), .B(new_new_n566_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n452_), .B(new_new_n75_), .Y(new_new_n568_));
  NA2        g546(.A(new_new_n129_), .B(i_8_), .Y(new_new_n569_));
  OAI210     g547(.A0(new_new_n569_), .A1(new_new_n568_), .B0(new_new_n567_), .Y(new_new_n570_));
  NA3        g548(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n218_), .B(i_4_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n572_), .B(i_8_), .Y(new_new_n573_));
  NA2        g551(.A(i_2_), .B(new_new_n77_), .Y(new_new_n574_));
  OAI210     g552(.A0(new_new_n80_), .A1(new_new_n186_), .B0(new_new_n187_), .Y(new_new_n575_));
  NO2        g553(.A(i_7_), .B(new_new_n37_), .Y(new_new_n576_));
  NA2        g554(.A(i_4_), .B(i_8_), .Y(new_new_n577_));
  AOI210     g555(.A0(new_new_n577_), .A1(new_new_n284_), .B0(new_new_n576_), .Y(new_new_n578_));
  OAI220     g556(.A0(new_new_n578_), .A1(new_new_n574_), .B0(new_new_n575_), .B1(i_13_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n579_), .B(new_new_n570_), .Y(new_new_n580_));
  OR2        g558(.A(i_6_), .B(i_10_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n581_), .B(new_new_n23_), .Y(new_new_n582_));
  OR3        g560(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n583_));
  NO3        g561(.A(new_new_n583_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n584_));
  INV        g562(.A(new_new_n183_), .Y(new_new_n585_));
  INV        g563(.A(new_new_n584_), .Y(new_new_n586_));
  OR2        g564(.A(new_new_n586_), .B(new_new_n552_), .Y(new_new_n587_));
  AOI210     g565(.A0(new_new_n587_), .A1(new_new_n580_), .B0(new_new_n57_), .Y(new_new_n588_));
  NOi21      g566(.An(i_11_), .B(i_7_), .Y(new_new_n589_));
  AO210      g567(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n590_), .B(new_new_n589_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(new_new_n189_), .Y(new_new_n592_));
  NA3        g570(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n593_));
  NAi31      g571(.An(new_new_n593_), .B(new_new_n196_), .C(i_11_), .Y(new_new_n594_));
  AOI210     g572(.A0(new_new_n594_), .A1(new_new_n592_), .B0(new_new_n57_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n596_));
  AO210      g574(.A0(new_new_n596_), .A1(new_new_n353_), .B0(new_new_n40_), .Y(new_new_n597_));
  NO3        g575(.A(new_new_n237_), .B(new_new_n190_), .C(i_8_), .Y(new_new_n598_));
  OAI210     g576(.A0(new_new_n598_), .A1(new_new_n207_), .B0(new_new_n57_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n382_), .B(new_new_n31_), .Y(new_new_n600_));
  OR2        g578(.A(new_new_n190_), .B(new_new_n99_), .Y(new_new_n601_));
  NA2        g579(.A(new_new_n601_), .B(new_new_n600_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n57_), .B(i_9_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n603_), .B(i_4_), .Y(new_new_n604_));
  NA2        g582(.A(new_new_n604_), .B(new_new_n602_), .Y(new_new_n605_));
  NO2        g583(.A(i_1_), .B(i_12_), .Y(new_new_n606_));
  NA3        g584(.A(new_new_n606_), .B(new_new_n101_), .C(new_new_n24_), .Y(new_new_n607_));
  NA4        g585(.A(new_new_n607_), .B(new_new_n605_), .C(new_new_n599_), .D(new_new_n597_), .Y(new_new_n608_));
  OAI210     g586(.A0(new_new_n608_), .A1(new_new_n595_), .B0(i_6_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n593_), .B(new_new_n99_), .Y(new_new_n610_));
  NA2        g588(.A(new_new_n610_), .B(new_new_n553_), .Y(new_new_n611_));
  NO2        g589(.A(i_6_), .B(i_11_), .Y(new_new_n612_));
  NA2        g590(.A(new_new_n611_), .B(new_new_n427_), .Y(new_new_n613_));
  NO4        g591(.A(new_new_n196_), .B(new_new_n115_), .C(i_13_), .D(new_new_n77_), .Y(new_new_n614_));
  NA2        g592(.A(new_new_n614_), .B(new_new_n603_), .Y(new_new_n615_));
  NO3        g593(.A(new_new_n581_), .B(new_new_n214_), .C(new_new_n23_), .Y(new_new_n616_));
  AOI210     g594(.A0(i_1_), .A1(new_new_n238_), .B0(new_new_n616_), .Y(new_new_n617_));
  OAI210     g595(.A0(new_new_n617_), .A1(new_new_n44_), .B0(new_new_n615_), .Y(new_new_n618_));
  NA3        g596(.A(new_new_n502_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n619_));
  NA2        g597(.A(new_new_n125_), .B(i_9_), .Y(new_new_n620_));
  NA3        g598(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n621_));
  NO2        g599(.A(new_new_n46_), .B(i_1_), .Y(new_new_n622_));
  NA3        g600(.A(new_new_n622_), .B(new_new_n246_), .C(new_new_n44_), .Y(new_new_n623_));
  OAI220     g601(.A0(new_new_n623_), .A1(new_new_n621_), .B0(new_new_n620_), .B1(new_new_n997_), .Y(new_new_n624_));
  NA3        g602(.A(new_new_n603_), .B(new_new_n297_), .C(i_6_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n23_), .Y(new_new_n626_));
  NO2        g604(.A(i_11_), .B(new_new_n37_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n627_), .B(new_new_n24_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n628_), .B(new_new_n46_), .Y(new_new_n629_));
  OR3        g607(.A(new_new_n629_), .B(new_new_n626_), .C(new_new_n624_), .Y(new_new_n630_));
  NO3        g608(.A(new_new_n630_), .B(new_new_n618_), .C(new_new_n613_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n218_), .B(new_new_n94_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n632_), .B(new_new_n589_), .Y(new_new_n633_));
  NA2        g611(.A(new_new_n633_), .B(i_1_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n634_), .B(new_new_n583_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n387_), .B(new_new_n77_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n635_), .B(new_new_n46_), .Y(new_new_n637_));
  NA2        g615(.A(i_3_), .B(new_new_n176_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n638_), .B(new_new_n105_), .Y(new_new_n639_));
  AN2        g617(.A(new_new_n639_), .B(new_new_n508_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n214_), .B(new_new_n44_), .Y(new_new_n641_));
  NO2        g619(.A(new_new_n106_), .B(new_new_n37_), .Y(new_new_n642_));
  NA2        g620(.A(i_1_), .B(i_3_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n428_), .B(new_new_n85_), .Y(new_new_n644_));
  AOI210     g622(.A0(new_new_n641_), .A1(new_new_n542_), .B0(new_new_n644_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n643_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n646_), .B(new_new_n640_), .Y(new_new_n647_));
  NA4        g625(.A(new_new_n647_), .B(new_new_n637_), .C(new_new_n631_), .D(new_new_n609_), .Y(new_new_n648_));
  NO3        g626(.A(new_new_n445_), .B(i_3_), .C(i_7_), .Y(new_new_n649_));
  NOi21      g627(.An(new_new_n649_), .B(i_10_), .Y(new_new_n650_));
  AN2        g628(.A(new_new_n650_), .B(new_new_n77_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n347_), .B(new_new_n346_), .Y(new_new_n652_));
  NO3        g630(.A(new_new_n446_), .B(new_new_n577_), .C(new_new_n77_), .Y(new_new_n653_));
  NA2        g631(.A(new_new_n653_), .B(new_new_n25_), .Y(new_new_n654_));
  NA2        g632(.A(new_new_n147_), .B(new_new_n77_), .Y(new_new_n655_));
  NA3        g633(.A(new_new_n655_), .B(new_new_n654_), .C(new_new_n652_), .Y(new_new_n656_));
  OAI210     g634(.A0(new_new_n656_), .A1(new_new_n651_), .B0(i_1_), .Y(new_new_n657_));
  NO2        g635(.A(new_new_n625_), .B(new_new_n419_), .Y(new_new_n658_));
  INV        g636(.A(new_new_n658_), .Y(new_new_n659_));
  AOI210     g637(.A0(new_new_n659_), .A1(new_new_n657_), .B0(i_13_), .Y(new_new_n660_));
  OR2        g638(.A(i_11_), .B(i_7_), .Y(new_new_n661_));
  NA3        g639(.A(new_new_n661_), .B(new_new_n98_), .C(new_new_n125_), .Y(new_new_n662_));
  AOI220     g640(.A0(new_new_n439_), .A1(new_new_n147_), .B0(new_new_n1002_), .B1(new_new_n125_), .Y(new_new_n663_));
  OAI210     g641(.A0(new_new_n663_), .A1(new_new_n44_), .B0(new_new_n662_), .Y(new_new_n664_));
  AOI220     g642(.A0(i_7_), .A1(new_new_n636_), .B0(new_new_n226_), .B1(new_new_n118_), .Y(new_new_n665_));
  OAI220     g643(.A0(new_new_n665_), .A1(new_new_n40_), .B0(new_new_n52_), .B1(new_new_n85_), .Y(new_new_n666_));
  AOI210     g644(.A0(new_new_n664_), .A1(new_new_n312_), .B0(new_new_n666_), .Y(new_new_n667_));
  AOI220     g645(.A0(i_12_), .A1(new_new_n64_), .B0(new_new_n359_), .B1(new_new_n622_), .Y(new_new_n668_));
  NO2        g646(.A(new_new_n668_), .B(new_new_n223_), .Y(new_new_n669_));
  AOI210     g647(.A0(new_new_n419_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n114_), .B(i_13_), .Y(new_new_n671_));
  NO2        g649(.A(new_new_n621_), .B(new_new_n105_), .Y(new_new_n672_));
  INV        g650(.A(new_new_n672_), .Y(new_new_n673_));
  OAI220     g651(.A0(new_new_n673_), .A1(new_new_n63_), .B0(new_new_n671_), .B1(new_new_n1006_), .Y(new_new_n674_));
  NO3        g652(.A(new_new_n63_), .B(new_new_n32_), .C(new_new_n94_), .Y(new_new_n675_));
  NA2        g653(.A(new_new_n26_), .B(new_new_n176_), .Y(new_new_n676_));
  INV        g654(.A(new_new_n675_), .Y(new_new_n677_));
  AOI210     g655(.A0(new_new_n359_), .A1(new_new_n622_), .B0(new_new_n84_), .Y(new_new_n678_));
  OAI220     g656(.A0(new_new_n678_), .A1(new_new_n573_), .B0(new_new_n677_), .B1(new_new_n585_), .Y(new_new_n679_));
  NO3        g657(.A(new_new_n679_), .B(new_new_n674_), .C(new_new_n669_), .Y(new_new_n680_));
  NA3        g658(.A(new_new_n382_), .B(new_new_n576_), .C(new_new_n90_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n612_), .B(i_13_), .Y(new_new_n682_));
  INV        g660(.A(new_new_n676_), .Y(new_new_n683_));
  NAi21      g661(.An(i_11_), .B(i_12_), .Y(new_new_n684_));
  NO3        g662(.A(new_new_n684_), .B(i_13_), .C(new_new_n77_), .Y(new_new_n685_));
  NO3        g663(.A(new_new_n446_), .B(new_new_n553_), .C(new_new_n577_), .Y(new_new_n686_));
  AOI220     g664(.A0(new_new_n686_), .A1(new_new_n291_), .B0(new_new_n685_), .B1(new_new_n683_), .Y(new_new_n687_));
  NA3        g665(.A(new_new_n687_), .B(new_new_n682_), .C(new_new_n681_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n688_), .B(new_new_n57_), .Y(new_new_n689_));
  NO2        g667(.A(i_2_), .B(i_12_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n344_), .B(new_new_n690_), .Y(new_new_n691_));
  NA2        g669(.A(i_8_), .B(new_new_n25_), .Y(new_new_n692_));
  NO2        g670(.A(new_new_n692_), .B(new_new_n358_), .Y(new_new_n693_));
  OAI210     g671(.A0(new_new_n693_), .A1(new_new_n346_), .B0(new_new_n344_), .Y(new_new_n694_));
  NO2        g672(.A(new_new_n115_), .B(i_2_), .Y(new_new_n695_));
  NA2        g673(.A(new_new_n695_), .B(new_new_n606_), .Y(new_new_n696_));
  NA3        g674(.A(new_new_n696_), .B(new_new_n694_), .C(new_new_n691_), .Y(new_new_n697_));
  NA3        g675(.A(new_new_n697_), .B(new_new_n45_), .C(new_new_n206_), .Y(new_new_n698_));
  NA4        g676(.A(new_new_n698_), .B(new_new_n689_), .C(new_new_n680_), .D(new_new_n667_), .Y(new_new_n699_));
  OR4        g677(.A(new_new_n699_), .B(new_new_n660_), .C(new_new_n648_), .D(new_new_n588_), .Y(men5));
  AOI210     g678(.A0(new_new_n633_), .A1(new_new_n248_), .B0(new_new_n389_), .Y(new_new_n701_));
  NA3        g679(.A(new_new_n24_), .B(new_new_n690_), .C(new_new_n99_), .Y(new_new_n702_));
  NA2        g680(.A(new_new_n702_), .B(new_new_n701_), .Y(new_new_n703_));
  NO3        g681(.A(i_11_), .B(new_new_n218_), .C(i_13_), .Y(new_new_n704_));
  NO2        g682(.A(new_new_n112_), .B(new_new_n23_), .Y(new_new_n705_));
  NA2        g683(.A(i_12_), .B(i_8_), .Y(new_new_n706_));
  OAI210     g684(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n706_), .Y(new_new_n707_));
  INV        g685(.A(new_new_n418_), .Y(new_new_n708_));
  AOI220     g686(.A0(new_new_n297_), .A1(new_new_n546_), .B0(new_new_n707_), .B1(new_new_n705_), .Y(new_new_n709_));
  INV        g687(.A(new_new_n709_), .Y(new_new_n710_));
  NO2        g688(.A(new_new_n710_), .B(new_new_n703_), .Y(new_new_n711_));
  INV        g689(.A(new_new_n155_), .Y(new_new_n712_));
  NO2        g690(.A(new_new_n428_), .B(new_new_n26_), .Y(new_new_n713_));
  NO2        g691(.A(new_new_n713_), .B(new_new_n390_), .Y(new_new_n714_));
  NA2        g692(.A(new_new_n714_), .B(i_2_), .Y(new_new_n715_));
  INV        g693(.A(new_new_n715_), .Y(new_new_n716_));
  AOI210     g694(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n388_), .Y(new_new_n717_));
  AOI210     g695(.A0(new_new_n717_), .A1(new_new_n716_), .B0(new_new_n226_), .Y(new_new_n718_));
  NO2        g696(.A(new_new_n173_), .B(new_new_n113_), .Y(new_new_n719_));
  OAI210     g697(.A0(new_new_n719_), .A1(new_new_n705_), .B0(i_2_), .Y(new_new_n720_));
  NO3        g698(.A(new_new_n590_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n721_));
  AOI210     g699(.A0(new_new_n155_), .A1(new_new_n80_), .B0(new_new_n721_), .Y(new_new_n722_));
  AOI210     g700(.A0(new_new_n722_), .A1(new_new_n720_), .B0(new_new_n176_), .Y(new_new_n723_));
  NA2        g701(.A(new_new_n183_), .B(new_new_n186_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n137_), .B(i_8_), .Y(new_new_n725_));
  AOI210     g703(.A0(new_new_n725_), .A1(new_new_n724_), .B0(new_new_n349_), .Y(new_new_n726_));
  NA2        g704(.A(new_new_n190_), .B(new_new_n133_), .Y(new_new_n727_));
  NA2        g705(.A(new_new_n727_), .B(new_new_n390_), .Y(new_new_n728_));
  NA3        g706(.A(new_new_n284_), .B(new_new_n112_), .C(new_new_n42_), .Y(new_new_n729_));
  OAI210     g707(.A0(new_new_n729_), .A1(new_new_n46_), .B0(new_new_n728_), .Y(new_new_n730_));
  NO3        g708(.A(new_new_n730_), .B(new_new_n726_), .C(new_new_n723_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n546_), .B(new_new_n28_), .Y(new_new_n732_));
  NA2        g710(.A(new_new_n704_), .B(new_new_n253_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n733_), .B(new_new_n732_), .Y(new_new_n734_));
  INV        g712(.A(new_new_n734_), .Y(new_new_n735_));
  NA4        g713(.A(new_new_n735_), .B(new_new_n731_), .C(new_new_n718_), .D(new_new_n711_), .Y(men6));
  NA2        g714(.A(new_new_n25_), .B(new_new_n695_), .Y(new_new_n737_));
  NA4        g715(.A(new_new_n363_), .B(new_new_n451_), .C(new_new_n63_), .D(new_new_n94_), .Y(new_new_n738_));
  INV        g716(.A(new_new_n738_), .Y(new_new_n739_));
  NO2        g717(.A(new_new_n202_), .B(i_2_), .Y(new_new_n740_));
  NO2        g718(.A(i_11_), .B(i_9_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n739_), .B(new_new_n307_), .Y(new_new_n742_));
  AO210      g720(.A0(new_new_n742_), .A1(new_new_n737_), .B0(i_12_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n350_), .B(new_new_n315_), .Y(new_new_n744_));
  NA2        g722(.A(new_new_n553_), .B(new_new_n57_), .Y(new_new_n745_));
  NA2        g723(.A(new_new_n650_), .B(new_new_n63_), .Y(new_new_n746_));
  NA4        g724(.A(new_new_n596_), .B(new_new_n746_), .C(new_new_n745_), .D(new_new_n744_), .Y(new_new_n747_));
  INV        g725(.A(new_new_n180_), .Y(new_new_n748_));
  AOI220     g726(.A0(new_new_n748_), .A1(new_new_n741_), .B0(new_new_n747_), .B1(new_new_n65_), .Y(new_new_n749_));
  INV        g727(.A(new_new_n306_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n67_), .B(new_new_n118_), .Y(new_new_n751_));
  INV        g729(.A(new_new_n112_), .Y(new_new_n752_));
  NA2        g730(.A(new_new_n752_), .B(new_new_n46_), .Y(new_new_n753_));
  AOI210     g731(.A0(new_new_n753_), .A1(new_new_n751_), .B0(new_new_n750_), .Y(new_new_n754_));
  INV        g732(.A(new_new_n485_), .Y(new_new_n755_));
  NO2        g733(.A(new_new_n32_), .B(i_11_), .Y(new_new_n756_));
  NA3        g734(.A(new_new_n756_), .B(new_new_n443_), .C(new_new_n363_), .Y(new_new_n757_));
  OAI210     g735(.A0(new_new_n649_), .A1(new_new_n535_), .B0(new_new_n534_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n758_), .B(new_new_n757_), .Y(new_new_n759_));
  OR3        g737(.A(new_new_n759_), .B(new_new_n755_), .C(new_new_n754_), .Y(new_new_n760_));
  NA3        g738(.A(new_new_n326_), .B(new_new_n235_), .C(i_7_), .Y(new_new_n761_));
  NA2        g739(.A(new_new_n420_), .B(new_new_n132_), .Y(new_new_n762_));
  AO210      g740(.A0(new_new_n461_), .A1(new_new_n708_), .B0(new_new_n36_), .Y(new_new_n763_));
  NA3        g741(.A(new_new_n763_), .B(new_new_n762_), .C(new_new_n761_), .Y(new_new_n764_));
  OAI210     g742(.A0(i_6_), .A1(i_11_), .B0(new_new_n78_), .Y(new_new_n765_));
  AOI220     g743(.A0(new_new_n765_), .A1(new_new_n534_), .B0(new_new_n740_), .B1(new_new_n1009_), .Y(new_new_n766_));
  NA3        g744(.A(new_new_n349_), .B(new_new_n219_), .C(new_new_n132_), .Y(new_new_n767_));
  OAI210     g745(.A0(new_new_n370_), .A1(new_new_n187_), .B0(new_new_n62_), .Y(new_new_n768_));
  NA4        g746(.A(new_new_n768_), .B(new_new_n767_), .C(new_new_n766_), .D(new_new_n575_), .Y(new_new_n769_));
  AO210      g747(.A0(new_new_n487_), .A1(new_new_n46_), .B0(new_new_n79_), .Y(new_new_n770_));
  NA3        g748(.A(new_new_n770_), .B(new_new_n452_), .C(new_new_n199_), .Y(new_new_n771_));
  INV        g749(.A(new_new_n533_), .Y(new_new_n772_));
  NO2        g750(.A(new_new_n581_), .B(i_2_), .Y(new_new_n773_));
  OAI210     g751(.A0(new_new_n773_), .A1(new_new_n102_), .B0(new_new_n380_), .Y(new_new_n774_));
  INV        g752(.A(new_new_n559_), .Y(new_new_n775_));
  NA3        g753(.A(new_new_n775_), .B(new_new_n306_), .C(i_7_), .Y(new_new_n776_));
  NA4        g754(.A(new_new_n776_), .B(new_new_n774_), .C(new_new_n772_), .D(new_new_n771_), .Y(new_new_n777_));
  NO4        g755(.A(new_new_n777_), .B(new_new_n769_), .C(new_new_n764_), .D(new_new_n760_), .Y(new_new_n778_));
  NA4        g756(.A(new_new_n778_), .B(new_new_n749_), .C(new_new_n743_), .D(new_new_n354_), .Y(men3));
  NA2        g757(.A(i_12_), .B(i_10_), .Y(new_new_n780_));
  NA2        g758(.A(i_6_), .B(i_7_), .Y(new_new_n781_));
  NO2        g759(.A(new_new_n781_), .B(i_0_), .Y(new_new_n782_));
  NO2        g760(.A(i_11_), .B(new_new_n218_), .Y(new_new_n783_));
  NA2        g761(.A(new_new_n268_), .B(new_new_n783_), .Y(new_new_n784_));
  NO2        g762(.A(new_new_n784_), .B(new_new_n176_), .Y(new_new_n785_));
  NO3        g763(.A(new_new_n424_), .B(new_new_n82_), .C(new_new_n44_), .Y(new_new_n786_));
  OA210      g764(.A0(new_new_n786_), .A1(new_new_n785_), .B0(new_new_n157_), .Y(new_new_n787_));
  NA3        g765(.A(new_new_n767_), .B(new_new_n575_), .C(new_new_n348_), .Y(new_new_n788_));
  NA2        g766(.A(new_new_n788_), .B(new_new_n39_), .Y(new_new_n789_));
  NO3        g767(.A(new_new_n601_), .B(new_new_n428_), .C(new_new_n118_), .Y(new_new_n790_));
  NA2        g768(.A(new_new_n382_), .B(new_new_n45_), .Y(new_new_n791_));
  AN2        g769(.A(new_new_n426_), .B(new_new_n53_), .Y(new_new_n792_));
  NO2        g770(.A(new_new_n792_), .B(new_new_n790_), .Y(new_new_n793_));
  AOI210     g771(.A0(new_new_n793_), .A1(new_new_n789_), .B0(new_new_n48_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n670_), .B(new_new_n1003_), .Y(new_new_n795_));
  NA2        g773(.A(new_new_n313_), .B(new_new_n408_), .Y(new_new_n796_));
  NO2        g774(.A(new_new_n796_), .B(new_new_n795_), .Y(new_new_n797_));
  NOi21      g775(.An(i_5_), .B(i_9_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n798_), .B(new_new_n416_), .Y(new_new_n799_));
  INV        g777(.A(new_new_n653_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n800_), .B(new_new_n799_), .Y(new_new_n801_));
  NO4        g779(.A(new_new_n801_), .B(new_new_n797_), .C(new_new_n794_), .D(new_new_n787_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n168_), .B(new_new_n24_), .Y(new_new_n803_));
  NO2        g781(.A(new_new_n642_), .B(new_new_n566_), .Y(new_new_n804_));
  NO2        g782(.A(new_new_n804_), .B(new_new_n803_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n291_), .B(new_new_n116_), .Y(new_new_n806_));
  NAi21      g784(.An(new_new_n148_), .B(new_new_n408_), .Y(new_new_n807_));
  NO2        g785(.A(new_new_n806_), .B(new_new_n373_), .Y(new_new_n808_));
  NO2        g786(.A(new_new_n808_), .B(new_new_n805_), .Y(new_new_n809_));
  NO2        g787(.A(new_new_n363_), .B(new_new_n272_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n810_), .B(new_new_n672_), .Y(new_new_n811_));
  NA2        g789(.A(new_new_n543_), .B(i_0_), .Y(new_new_n812_));
  NO3        g790(.A(new_new_n812_), .B(new_new_n1007_), .C(new_new_n80_), .Y(new_new_n813_));
  NO4        g791(.A(new_new_n559_), .B(new_new_n196_), .C(new_new_n388_), .D(i_6_), .Y(new_new_n814_));
  INV        g792(.A(new_new_n813_), .Y(new_new_n815_));
  AN2        g793(.A(new_new_n89_), .B(new_new_n224_), .Y(new_new_n816_));
  NA2        g794(.A(new_new_n704_), .B(new_new_n307_), .Y(new_new_n817_));
  AOI210     g795(.A0(new_new_n452_), .A1(new_new_n80_), .B0(new_new_n54_), .Y(new_new_n818_));
  OAI220     g796(.A0(new_new_n818_), .A1(new_new_n817_), .B0(new_new_n628_), .B1(new_new_n504_), .Y(new_new_n819_));
  NA2        g797(.A(i_0_), .B(i_10_), .Y(new_new_n820_));
  NO4        g798(.A(new_new_n105_), .B(new_new_n54_), .C(new_new_n638_), .D(i_5_), .Y(new_new_n821_));
  AN2        g799(.A(new_new_n821_), .B(i_10_), .Y(new_new_n822_));
  AOI220     g800(.A0(new_new_n313_), .A1(new_new_n91_), .B0(new_new_n168_), .B1(new_new_n75_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n537_), .B(i_4_), .Y(new_new_n824_));
  NA2        g802(.A(new_new_n171_), .B(new_new_n186_), .Y(new_new_n825_));
  OAI220     g803(.A0(new_new_n825_), .A1(new_new_n817_), .B0(new_new_n824_), .B1(new_new_n823_), .Y(new_new_n826_));
  NO4        g804(.A(new_new_n826_), .B(new_new_n822_), .C(new_new_n819_), .D(new_new_n816_), .Y(new_new_n827_));
  NA4        g805(.A(new_new_n827_), .B(new_new_n815_), .C(new_new_n811_), .D(new_new_n809_), .Y(new_new_n828_));
  NO2        g806(.A(new_new_n95_), .B(new_new_n37_), .Y(new_new_n829_));
  NA2        g807(.A(i_11_), .B(i_9_), .Y(new_new_n830_));
  NO3        g808(.A(i_12_), .B(new_new_n830_), .C(new_new_n574_), .Y(new_new_n831_));
  AN2        g809(.A(new_new_n831_), .B(new_new_n829_), .Y(new_new_n832_));
  NO2        g810(.A(new_new_n48_), .B(i_7_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n367_), .B(new_new_n162_), .Y(new_new_n834_));
  NA2        g812(.A(new_new_n834_), .B(new_new_n146_), .Y(new_new_n835_));
  NO2        g813(.A(new_new_n830_), .B(new_new_n65_), .Y(new_new_n836_));
  NO2        g814(.A(new_new_n158_), .B(i_0_), .Y(new_new_n837_));
  INV        g815(.A(new_new_n837_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n443_), .B(new_new_n212_), .Y(new_new_n839_));
  AOI210     g817(.A0(new_new_n347_), .A1(new_new_n41_), .B0(new_new_n379_), .Y(new_new_n840_));
  OAI220     g818(.A0(new_new_n840_), .A1(new_new_n799_), .B0(new_new_n839_), .B1(new_new_n838_), .Y(new_new_n841_));
  NO3        g819(.A(new_new_n841_), .B(new_new_n835_), .C(new_new_n832_), .Y(new_new_n842_));
  NA2        g820(.A(new_new_n627_), .B(new_new_n109_), .Y(new_new_n843_));
  NO2        g821(.A(i_6_), .B(new_new_n843_), .Y(new_new_n844_));
  AOI210     g822(.A0(new_new_n419_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n845_));
  NA2        g823(.A(new_new_n155_), .B(new_new_n95_), .Y(new_new_n846_));
  NOi32      g824(.An(new_new_n845_), .Bn(new_new_n171_), .C(new_new_n846_), .Y(new_new_n847_));
  NO2        g825(.A(new_new_n1000_), .B(new_new_n791_), .Y(new_new_n848_));
  NO3        g826(.A(new_new_n848_), .B(new_new_n847_), .C(new_new_n844_), .Y(new_new_n849_));
  NOi21      g827(.An(i_7_), .B(i_5_), .Y(new_new_n850_));
  NOi31      g828(.An(new_new_n850_), .B(i_0_), .C(new_new_n684_), .Y(new_new_n851_));
  NA3        g829(.A(new_new_n851_), .B(new_new_n358_), .C(i_6_), .Y(new_new_n852_));
  OA210      g830(.A0(new_new_n846_), .A1(new_new_n485_), .B0(new_new_n852_), .Y(new_new_n853_));
  NO3        g831(.A(new_new_n376_), .B(new_new_n337_), .C(new_new_n333_), .Y(new_new_n854_));
  INV        g832(.A(new_new_n298_), .Y(new_new_n855_));
  INV        g833(.A(new_new_n854_), .Y(new_new_n856_));
  NA4        g834(.A(new_new_n856_), .B(new_new_n853_), .C(new_new_n849_), .D(new_new_n842_), .Y(new_new_n857_));
  NO2        g835(.A(new_new_n803_), .B(new_new_n220_), .Y(new_new_n858_));
  AN2        g836(.A(new_new_n312_), .B(new_new_n307_), .Y(new_new_n859_));
  NA2        g837(.A(new_new_n858_), .B(i_10_), .Y(new_new_n860_));
  NO2        g838(.A(new_new_n780_), .B(new_new_n297_), .Y(new_new_n861_));
  OA210      g839(.A0(new_new_n443_), .A1(new_new_n204_), .B0(new_new_n442_), .Y(new_new_n862_));
  NA2        g840(.A(new_new_n861_), .B(new_new_n836_), .Y(new_new_n863_));
  NO2        g841(.A(new_new_n807_), .B(i_6_), .Y(new_new_n864_));
  NO2        g842(.A(new_new_n235_), .B(new_new_n46_), .Y(new_new_n865_));
  NA2        g843(.A(new_new_n836_), .B(new_new_n284_), .Y(new_new_n866_));
  OAI210     g844(.A0(new_new_n865_), .A1(new_new_n170_), .B0(new_new_n866_), .Y(new_new_n867_));
  AOI220     g845(.A0(new_new_n867_), .A1(new_new_n443_), .B0(new_new_n864_), .B1(new_new_n65_), .Y(new_new_n868_));
  NO2        g846(.A(new_new_n67_), .B(new_new_n706_), .Y(new_new_n869_));
  AOI220     g847(.A0(new_new_n869_), .A1(i_11_), .B0(new_new_n157_), .B1(new_new_n566_), .Y(new_new_n870_));
  NO2        g848(.A(new_new_n870_), .B(new_new_n47_), .Y(new_new_n871_));
  NO3        g849(.A(new_new_n559_), .B(i_0_), .C(new_new_n24_), .Y(new_new_n872_));
  AOI210     g850(.A0(i_7_), .A1(new_new_n516_), .B0(new_new_n872_), .Y(new_new_n873_));
  NAi21      g851(.An(i_9_), .B(i_5_), .Y(new_new_n874_));
  NO2        g852(.A(new_new_n874_), .B(new_new_n376_), .Y(new_new_n875_));
  NO2        g853(.A(new_new_n571_), .B(new_new_n97_), .Y(new_new_n876_));
  AOI220     g854(.A0(new_new_n876_), .A1(i_0_), .B0(new_new_n875_), .B1(new_new_n591_), .Y(new_new_n877_));
  OAI220     g855(.A0(new_new_n877_), .A1(new_new_n77_), .B0(new_new_n873_), .B1(new_new_n156_), .Y(new_new_n878_));
  NO3        g856(.A(new_new_n878_), .B(new_new_n871_), .C(new_new_n488_), .Y(new_new_n879_));
  NA4        g857(.A(new_new_n879_), .B(new_new_n868_), .C(new_new_n863_), .D(new_new_n860_), .Y(new_new_n880_));
  NO3        g858(.A(new_new_n880_), .B(new_new_n857_), .C(new_new_n828_), .Y(new_new_n881_));
  NO2        g859(.A(i_0_), .B(new_new_n684_), .Y(new_new_n882_));
  NA2        g860(.A(new_new_n65_), .B(new_new_n44_), .Y(new_new_n883_));
  NO3        g861(.A(new_new_n97_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n884_));
  AO220      g862(.A0(new_new_n884_), .A1(new_new_n65_), .B0(new_new_n882_), .B1(new_new_n157_), .Y(new_new_n885_));
  AOI210     g863(.A0(new_new_n745_), .A1(new_new_n652_), .B0(new_new_n846_), .Y(new_new_n886_));
  AOI210     g864(.A0(new_new_n885_), .A1(new_new_n323_), .B0(new_new_n886_), .Y(new_new_n887_));
  NA2        g865(.A(new_new_n695_), .B(new_new_n131_), .Y(new_new_n888_));
  NO2        g866(.A(new_new_n758_), .B(new_new_n376_), .Y(new_new_n889_));
  NA3        g867(.A(new_new_n782_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n890_));
  NA2        g868(.A(new_new_n783_), .B(i_9_), .Y(new_new_n891_));
  AOI210     g869(.A0(new_new_n890_), .A1(new_new_n465_), .B0(new_new_n891_), .Y(new_new_n892_));
  OAI210     g870(.A0(new_new_n225_), .A1(i_9_), .B0(new_new_n211_), .Y(new_new_n893_));
  AOI210     g871(.A0(new_new_n893_), .A1(new_new_n812_), .B0(new_new_n139_), .Y(new_new_n894_));
  NO3        g872(.A(new_new_n894_), .B(new_new_n892_), .C(new_new_n889_), .Y(new_new_n895_));
  NA3        g873(.A(new_new_n895_), .B(new_new_n888_), .C(new_new_n887_), .Y(new_new_n896_));
  INV        g874(.A(new_new_n859_), .Y(new_new_n897_));
  AOI210     g875(.A0(new_new_n279_), .A1(new_new_n148_), .B0(new_new_n897_), .Y(new_new_n898_));
  NA3        g876(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n899_));
  NA2        g877(.A(new_new_n833_), .B(new_new_n456_), .Y(new_new_n900_));
  AOI210     g878(.A0(new_new_n899_), .A1(new_new_n148_), .B0(new_new_n900_), .Y(new_new_n901_));
  NO2        g879(.A(new_new_n901_), .B(new_new_n898_), .Y(new_new_n902_));
  NO3        g880(.A(new_new_n820_), .B(new_new_n798_), .C(new_new_n173_), .Y(new_new_n903_));
  AOI220     g881(.A0(new_new_n903_), .A1(i_11_), .B0(new_new_n538_), .B1(new_new_n67_), .Y(new_new_n904_));
  NA2        g882(.A(new_new_n68_), .B(i_13_), .Y(new_new_n905_));
  INV        g883(.A(new_new_n199_), .Y(new_new_n906_));
  OAI220     g884(.A0(new_new_n498_), .A1(new_new_n1005_), .B0(i_12_), .B1(new_new_n585_), .Y(new_new_n907_));
  NA3        g885(.A(new_new_n907_), .B(new_new_n371_), .C(new_new_n906_), .Y(new_new_n908_));
  NA4        g886(.A(new_new_n908_), .B(new_new_n905_), .C(new_new_n904_), .D(new_new_n902_), .Y(new_new_n909_));
  NO2        g887(.A(new_new_n223_), .B(new_new_n85_), .Y(new_new_n910_));
  AOI210     g888(.A0(new_new_n910_), .A1(new_new_n882_), .B0(new_new_n100_), .Y(new_new_n911_));
  AOI220     g889(.A0(new_new_n850_), .A1(new_new_n456_), .B0(new_new_n782_), .B1(new_new_n149_), .Y(new_new_n912_));
  NA2        g890(.A(new_new_n326_), .B(new_new_n159_), .Y(new_new_n913_));
  OA220      g891(.A0(new_new_n913_), .A1(new_new_n912_), .B0(new_new_n911_), .B1(i_5_), .Y(new_new_n914_));
  AOI210     g892(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n158_), .Y(new_new_n915_));
  NA2        g893(.A(new_new_n915_), .B(new_new_n862_), .Y(new_new_n916_));
  NA3        g894(.A(new_new_n582_), .B(new_new_n168_), .C(new_new_n75_), .Y(new_new_n917_));
  NA2        g895(.A(new_new_n917_), .B(new_new_n514_), .Y(new_new_n918_));
  NA3        g896(.A(new_new_n460_), .B(new_new_n455_), .C(new_new_n440_), .Y(new_new_n919_));
  NO2        g897(.A(new_new_n919_), .B(new_new_n918_), .Y(new_new_n920_));
  NA3        g898(.A(new_new_n363_), .B(new_new_n155_), .C(new_new_n154_), .Y(new_new_n921_));
  NA3        g899(.A(new_new_n833_), .B(new_new_n268_), .C(new_new_n211_), .Y(new_new_n922_));
  NA2        g900(.A(new_new_n922_), .B(new_new_n921_), .Y(new_new_n923_));
  NA3        g901(.A(new_new_n363_), .B(new_new_n314_), .C(new_new_n203_), .Y(new_new_n924_));
  INV        g902(.A(new_new_n924_), .Y(new_new_n925_));
  NOi31      g903(.An(new_new_n362_), .B(new_new_n883_), .C(new_new_n220_), .Y(new_new_n926_));
  NO3        g904(.A(new_new_n926_), .B(new_new_n925_), .C(new_new_n923_), .Y(new_new_n927_));
  NA4        g905(.A(new_new_n927_), .B(new_new_n920_), .C(new_new_n916_), .D(new_new_n914_), .Y(new_new_n928_));
  INV        g906(.A(new_new_n584_), .Y(new_new_n929_));
  NO3        g907(.A(new_new_n929_), .B(new_new_n529_), .C(i_3_), .Y(new_new_n930_));
  NO2        g908(.A(new_new_n77_), .B(i_5_), .Y(new_new_n931_));
  NA3        g909(.A(new_new_n783_), .B(new_new_n101_), .C(new_new_n112_), .Y(new_new_n932_));
  INV        g910(.A(new_new_n932_), .Y(new_new_n933_));
  AOI210     g911(.A0(new_new_n933_), .A1(new_new_n931_), .B0(new_new_n930_), .Y(new_new_n934_));
  NA3        g912(.A(new_new_n284_), .B(i_5_), .C(new_new_n176_), .Y(new_new_n935_));
  NO3        g913(.A(new_new_n220_), .B(i_0_), .C(i_12_), .Y(new_new_n936_));
  AOI220     g914(.A0(new_new_n936_), .A1(new_new_n222_), .B0(new_new_n739_), .B1(new_new_n159_), .Y(new_new_n937_));
  AN2        g915(.A(new_new_n820_), .B(new_new_n139_), .Y(new_new_n938_));
  NO4        g916(.A(new_new_n938_), .B(i_12_), .C(new_new_n619_), .D(new_new_n118_), .Y(new_new_n939_));
  NA2        g917(.A(new_new_n939_), .B(new_new_n199_), .Y(new_new_n940_));
  NA3        g918(.A(new_new_n91_), .B(new_new_n542_), .C(i_11_), .Y(new_new_n941_));
  NO2        g919(.A(new_new_n941_), .B(new_new_n141_), .Y(new_new_n942_));
  NA2        g920(.A(new_new_n850_), .B(new_new_n439_), .Y(new_new_n943_));
  INV        g921(.A(new_new_n58_), .Y(new_new_n944_));
  OAI210     g922(.A0(new_new_n944_), .A1(new_new_n935_), .B0(new_new_n943_), .Y(new_new_n945_));
  AOI210     g923(.A0(new_new_n945_), .A1(new_new_n837_), .B0(new_new_n942_), .Y(new_new_n946_));
  NA4        g924(.A(new_new_n946_), .B(new_new_n940_), .C(new_new_n937_), .D(new_new_n934_), .Y(new_new_n947_));
  NO4        g925(.A(new_new_n947_), .B(new_new_n928_), .C(new_new_n909_), .D(new_new_n896_), .Y(new_new_n948_));
  NA2        g926(.A(new_new_n756_), .B(new_new_n37_), .Y(new_new_n949_));
  NA3        g927(.A(new_new_n845_), .B(new_new_n344_), .C(i_5_), .Y(new_new_n950_));
  NA2        g928(.A(new_new_n950_), .B(new_new_n949_), .Y(new_new_n951_));
  NA2        g929(.A(new_new_n951_), .B(new_new_n189_), .Y(new_new_n952_));
  AN2        g930(.A(new_new_n661_), .B(new_new_n345_), .Y(new_new_n953_));
  NA2        g931(.A(new_new_n169_), .B(new_new_n171_), .Y(new_new_n954_));
  AO210      g932(.A0(new_new_n953_), .A1(new_new_n33_), .B0(new_new_n954_), .Y(new_new_n955_));
  OAI210     g933(.A0(new_new_n584_), .A1(new_new_n582_), .B0(new_new_n297_), .Y(new_new_n956_));
  NAi31      g934(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n957_));
  NO2        g935(.A(new_new_n62_), .B(new_new_n957_), .Y(new_new_n958_));
  NO2        g936(.A(new_new_n958_), .B(new_new_n616_), .Y(new_new_n959_));
  NA3        g937(.A(new_new_n959_), .B(new_new_n956_), .C(new_new_n955_), .Y(new_new_n960_));
  NO4        g938(.A(new_new_n214_), .B(new_new_n130_), .C(new_new_n643_), .D(new_new_n37_), .Y(new_new_n961_));
  NO2        g939(.A(new_new_n961_), .B(new_new_n814_), .Y(new_new_n962_));
  OAI210     g940(.A0(new_new_n941_), .A1(new_new_n133_), .B0(new_new_n962_), .Y(new_new_n963_));
  AOI210     g941(.A0(new_new_n960_), .A1(new_new_n48_), .B0(new_new_n963_), .Y(new_new_n964_));
  AOI210     g942(.A0(new_new_n964_), .A1(new_new_n952_), .B0(new_new_n65_), .Y(new_new_n965_));
  NO2        g943(.A(new_new_n998_), .B(new_new_n712_), .Y(new_new_n966_));
  OAI210     g944(.A0(new_new_n72_), .A1(new_new_n52_), .B0(new_new_n99_), .Y(new_new_n967_));
  NA2        g945(.A(new_new_n967_), .B(new_new_n68_), .Y(new_new_n968_));
  AOI210     g946(.A0(new_new_n915_), .A1(new_new_n833_), .B0(new_new_n851_), .Y(new_new_n969_));
  AOI210     g947(.A0(new_new_n969_), .A1(new_new_n968_), .B0(new_new_n643_), .Y(new_new_n970_));
  INV        g948(.A(new_new_n241_), .Y(new_new_n971_));
  AOI220     g949(.A0(new_new_n971_), .A1(new_new_n68_), .B0(new_new_n321_), .B1(new_new_n234_), .Y(new_new_n972_));
  NO2        g950(.A(new_new_n972_), .B(new_new_n218_), .Y(new_new_n973_));
  NA3        g951(.A(new_new_n89_), .B(new_new_n286_), .C(new_new_n31_), .Y(new_new_n974_));
  INV        g952(.A(new_new_n974_), .Y(new_new_n975_));
  NO3        g953(.A(new_new_n975_), .B(new_new_n973_), .C(new_new_n970_), .Y(new_new_n976_));
  OAI210     g954(.A0(new_new_n247_), .A1(new_new_n144_), .B0(new_new_n80_), .Y(new_new_n977_));
  NA3        g955(.A(new_new_n713_), .B(new_new_n268_), .C(new_new_n72_), .Y(new_new_n978_));
  AOI210     g956(.A0(new_new_n978_), .A1(new_new_n977_), .B0(i_11_), .Y(new_new_n979_));
  NA2        g957(.A(new_new_n577_), .B(new_new_n196_), .Y(new_new_n980_));
  NA2        g958(.A(new_new_n980_), .B(new_new_n189_), .Y(new_new_n981_));
  NA2        g959(.A(new_new_n150_), .B(i_5_), .Y(new_new_n982_));
  AOI210     g960(.A0(new_new_n981_), .A1(new_new_n724_), .B0(new_new_n982_), .Y(new_new_n983_));
  NO3        g961(.A(new_new_n55_), .B(new_new_n54_), .C(i_4_), .Y(new_new_n984_));
  OAI210     g962(.A0(new_new_n855_), .A1(new_new_n286_), .B0(new_new_n984_), .Y(new_new_n985_));
  NO2        g963(.A(new_new_n985_), .B(new_new_n684_), .Y(new_new_n986_));
  NO4        g964(.A(new_new_n874_), .B(new_new_n445_), .C(new_new_n231_), .D(new_new_n230_), .Y(new_new_n987_));
  NO2        g965(.A(new_new_n987_), .B(new_new_n533_), .Y(new_new_n988_));
  INV        g966(.A(new_new_n338_), .Y(new_new_n989_));
  AOI210     g967(.A0(new_new_n989_), .A1(new_new_n988_), .B0(new_new_n40_), .Y(new_new_n990_));
  NO4        g968(.A(new_new_n990_), .B(new_new_n986_), .C(new_new_n983_), .D(new_new_n979_), .Y(new_new_n991_));
  OAI210     g969(.A0(new_new_n976_), .A1(i_4_), .B0(new_new_n991_), .Y(new_new_n992_));
  NO3        g970(.A(new_new_n992_), .B(new_new_n966_), .C(new_new_n965_), .Y(new_new_n993_));
  NA4        g971(.A(new_new_n993_), .B(new_new_n948_), .C(new_new_n881_), .D(new_new_n802_), .Y(men4));
  INV        g972(.A(i_2_), .Y(new_new_n997_));
  INV        g973(.A(new_new_n536_), .Y(new_new_n998_));
  INV        g974(.A(i_3_), .Y(new_new_n999_));
  INV        g975(.A(new_new_n307_), .Y(new_new_n1000_));
  INV        g976(.A(i_0_), .Y(new_new_n1001_));
  INV        g977(.A(i_4_), .Y(new_new_n1002_));
  INV        g978(.A(i_9_), .Y(new_new_n1003_));
  INV        g979(.A(i_10_), .Y(new_new_n1004_));
  INV        g980(.A(i_6_), .Y(new_new_n1005_));
  INV        g981(.A(i_1_), .Y(new_new_n1006_));
  INV        g982(.A(new_new_n357_), .Y(new_new_n1007_));
  INV        g983(.A(i_10_), .Y(new_new_n1008_));
  INV        g984(.A(i_7_), .Y(new_new_n1009_));
  INV        g985(.A(i_5_), .Y(new_new_n1010_));
  INV        g986(.A(new_new_n145_), .Y(new_new_n1011_));
endmodule


