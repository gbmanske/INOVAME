//Benchmark atmr_max1024_476_0.5

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  INV        o003(.A(ori_ori_n19_), .Y(ori_ori_n20_));
  NA2        o004(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n21_));
  INV        o005(.A(x5), .Y(ori_ori_n22_));
  NA2        o006(.A(x8), .B(x3), .Y(ori_ori_n23_));
  NA2        o007(.A(x4), .B(x2), .Y(ori_ori_n24_));
  INV        o008(.A(ori_ori_n21_), .Y(ori_ori_n25_));
  NO2        o009(.A(x4), .B(x3), .Y(ori_ori_n26_));
  INV        o010(.A(ori_ori_n26_), .Y(ori_ori_n27_));
  NOi21      o011(.An(ori_ori_n20_), .B(ori_ori_n25_), .Y(ori00));
  NO2        o012(.A(x1), .B(x0), .Y(ori_ori_n29_));
  INV        o013(.A(x6), .Y(ori_ori_n30_));
  NA2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  NO2        o015(.A(ori_ori_n20_), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NO2        o016(.A(x2), .B(x0), .Y(ori_ori_n33_));
  INV        o017(.A(x3), .Y(ori_ori_n34_));
  NO2        o018(.A(ori_ori_n34_), .B(ori_ori_n18_), .Y(ori_ori_n35_));
  INV        o019(.A(ori_ori_n35_), .Y(ori_ori_n36_));
  INV        o020(.A(ori_ori_n33_), .Y(ori_ori_n37_));
  INV        o021(.A(x4), .Y(ori_ori_n38_));
  NO2        o022(.A(ori_ori_n38_), .B(ori_ori_n17_), .Y(ori_ori_n39_));
  NA2        o023(.A(ori_ori_n39_), .B(x2), .Y(ori_ori_n40_));
  NA2        o024(.A(ori_ori_n40_), .B(ori_ori_n37_), .Y(ori_ori_n41_));
  INV        o025(.A(ori_ori_n29_), .Y(ori_ori_n42_));
  INV        o026(.A(x2), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n44_));
  NA2        o028(.A(ori_ori_n34_), .B(ori_ori_n18_), .Y(ori_ori_n45_));
  NA2        o029(.A(ori_ori_n45_), .B(ori_ori_n44_), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n42_), .A1(ori_ori_n27_), .B0(ori_ori_n46_), .Y(ori_ori_n47_));
  NO3        o031(.A(ori_ori_n47_), .B(ori_ori_n41_), .C(ori_ori_n32_), .Y(ori01));
  NA2        o032(.A(ori_ori_n34_), .B(x1), .Y(ori_ori_n49_));
  INV        o033(.A(x9), .Y(ori_ori_n50_));
  NO2        o034(.A(ori_ori_n49_), .B(x5), .Y(ori_ori_n51_));
  OAI210     o035(.A0(ori_ori_n35_), .A1(ori_ori_n22_), .B0(ori_ori_n43_), .Y(ori_ori_n52_));
  NA2        o036(.A(ori_ori_n45_), .B(ori_ori_n52_), .Y(ori_ori_n53_));
  INV        o037(.A(ori_ori_n53_), .Y(ori_ori_n54_));
  NA2        o038(.A(ori_ori_n54_), .B(x4), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n38_), .B(x2), .Y(ori_ori_n56_));
  OAI210     o040(.A0(ori_ori_n56_), .A1(ori_ori_n45_), .B0(x0), .Y(ori_ori_n57_));
  NA2        o041(.A(x5), .B(x3), .Y(ori_ori_n58_));
  NO2        o042(.A(x8), .B(x6), .Y(ori_ori_n59_));
  NAi21      o043(.An(x4), .B(x3), .Y(ori_ori_n60_));
  INV        o044(.A(ori_ori_n60_), .Y(ori_ori_n61_));
  NO2        o045(.A(x4), .B(x2), .Y(ori_ori_n62_));
  NO2        o046(.A(ori_ori_n60_), .B(ori_ori_n18_), .Y(ori_ori_n63_));
  NO2        o047(.A(ori_ori_n63_), .B(ori_ori_n57_), .Y(ori_ori_n64_));
  NA2        o048(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n65_));
  INV        o049(.A(x8), .Y(ori_ori_n66_));
  NA2        o050(.A(x2), .B(x1), .Y(ori_ori_n67_));
  AOI210     o051(.A0(ori_ori_n45_), .A1(ori_ori_n22_), .B0(ori_ori_n43_), .Y(ori_ori_n68_));
  NA2        o052(.A(ori_ori_n36_), .B(ori_ori_n38_), .Y(ori_ori_n69_));
  NO2        o053(.A(ori_ori_n69_), .B(ori_ori_n68_), .Y(ori_ori_n70_));
  NA2        o054(.A(x4), .B(ori_ori_n34_), .Y(ori_ori_n71_));
  NO2        o055(.A(ori_ori_n38_), .B(ori_ori_n43_), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n73_));
  OAI210     o057(.A0(ori_ori_n73_), .A1(ori_ori_n31_), .B0(ori_ori_n17_), .Y(ori_ori_n74_));
  NO2        o058(.A(ori_ori_n74_), .B(ori_ori_n70_), .Y(ori_ori_n75_));
  AO210      o059(.A0(ori_ori_n64_), .A1(ori_ori_n55_), .B0(ori_ori_n75_), .Y(ori02));
  OR2        o060(.A(x8), .B(x0), .Y(ori_ori_n77_));
  INV        o061(.A(ori_ori_n77_), .Y(ori_ori_n78_));
  NO2        o062(.A(x4), .B(x1), .Y(ori_ori_n79_));
  NA2        o063(.A(ori_ori_n79_), .B(x2), .Y(ori_ori_n80_));
  NOi21      o064(.An(x0), .B(x4), .Y(ori_ori_n81_));
  NO2        o065(.A(ori_ori_n80_), .B(ori_ori_n58_), .Y(ori_ori_n82_));
  NO2        o066(.A(x5), .B(ori_ori_n38_), .Y(ori_ori_n83_));
  NAi21      o067(.An(x0), .B(x4), .Y(ori_ori_n84_));
  NO2        o068(.A(ori_ori_n84_), .B(x1), .Y(ori_ori_n85_));
  NO2        o069(.A(x7), .B(x0), .Y(ori_ori_n86_));
  NO2        o070(.A(ori_ori_n62_), .B(ori_ori_n72_), .Y(ori_ori_n87_));
  NO2        o071(.A(ori_ori_n87_), .B(x3), .Y(ori_ori_n88_));
  OAI210     o072(.A0(ori_ori_n86_), .A1(ori_ori_n85_), .B0(ori_ori_n88_), .Y(ori_ori_n89_));
  NA2        o073(.A(x5), .B(x0), .Y(ori_ori_n90_));
  NO2        o074(.A(ori_ori_n38_), .B(x2), .Y(ori_ori_n91_));
  NA2        o075(.A(ori_ori_n89_), .B(ori_ori_n30_), .Y(ori_ori_n92_));
  NO2        o076(.A(ori_ori_n92_), .B(ori_ori_n82_), .Y(ori_ori_n93_));
  NO3        o077(.A(ori_ori_n58_), .B(ori_ori_n56_), .C(ori_ori_n21_), .Y(ori_ori_n94_));
  NO2        o078(.A(ori_ori_n24_), .B(ori_ori_n22_), .Y(ori_ori_n95_));
  NA2        o079(.A(x7), .B(x3), .Y(ori_ori_n96_));
  NO2        o080(.A(ori_ori_n71_), .B(x5), .Y(ori_ori_n97_));
  BUFFER     o081(.A(x8), .Y(ori_ori_n98_));
  NO2        o082(.A(ori_ori_n34_), .B(x2), .Y(ori_ori_n99_));
  INV        o083(.A(x7), .Y(ori_ori_n100_));
  NA2        o084(.A(ori_ori_n100_), .B(ori_ori_n18_), .Y(ori_ori_n101_));
  NA2        o085(.A(x5), .B(x1), .Y(ori_ori_n102_));
  INV        o086(.A(ori_ori_n102_), .Y(ori_ori_n103_));
  AOI210     o087(.A0(ori_ori_n103_), .A1(ori_ori_n81_), .B0(ori_ori_n30_), .Y(ori_ori_n104_));
  NAi21      o088(.An(x2), .B(x7), .Y(ori_ori_n105_));
  NO2        o089(.A(ori_ori_n105_), .B(ori_ori_n38_), .Y(ori_ori_n106_));
  NA2        o090(.A(ori_ori_n286_), .B(ori_ori_n104_), .Y(ori_ori_n107_));
  NO2        o091(.A(ori_ori_n107_), .B(ori_ori_n94_), .Y(ori_ori_n108_));
  NO2        o092(.A(ori_ori_n108_), .B(ori_ori_n93_), .Y(ori_ori_n109_));
  NO2        o093(.A(ori_ori_n90_), .B(ori_ori_n87_), .Y(ori_ori_n110_));
  NA2        o094(.A(ori_ori_n22_), .B(ori_ori_n18_), .Y(ori_ori_n111_));
  NA2        o095(.A(ori_ori_n22_), .B(ori_ori_n17_), .Y(ori_ori_n112_));
  NA3        o096(.A(ori_ori_n112_), .B(ori_ori_n111_), .C(ori_ori_n21_), .Y(ori_ori_n113_));
  AN2        o097(.A(ori_ori_n113_), .B(ori_ori_n91_), .Y(ori_ori_n114_));
  NA2        o098(.A(x8), .B(x0), .Y(ori_ori_n115_));
  NO2        o099(.A(ori_ori_n100_), .B(ori_ori_n22_), .Y(ori_ori_n116_));
  NO2        o100(.A(ori_ori_n115_), .B(ori_ori_n22_), .Y(ori_ori_n117_));
  NA2        o101(.A(x4), .B(x1), .Y(ori_ori_n118_));
  NO3        o102(.A(ori_ori_n117_), .B(ori_ori_n114_), .C(ori_ori_n110_), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n119_), .B(ori_ori_n34_), .Y(ori_ori_n120_));
  NO2        o104(.A(ori_ori_n113_), .B(ori_ori_n56_), .Y(ori_ori_n121_));
  INV        o105(.A(ori_ori_n83_), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n73_), .B(ori_ori_n17_), .Y(ori_ori_n123_));
  NO2        o107(.A(ori_ori_n29_), .B(ori_ori_n123_), .Y(ori_ori_n124_));
  NO3        o108(.A(ori_ori_n124_), .B(ori_ori_n122_), .C(x7), .Y(ori_ori_n125_));
  NO2        o109(.A(ori_ori_n112_), .B(ori_ori_n87_), .Y(ori_ori_n126_));
  NO3        o110(.A(ori_ori_n126_), .B(ori_ori_n125_), .C(ori_ori_n121_), .Y(ori_ori_n127_));
  NO2        o111(.A(ori_ori_n127_), .B(x3), .Y(ori_ori_n128_));
  NO3        o112(.A(ori_ori_n128_), .B(ori_ori_n120_), .C(ori_ori_n109_), .Y(ori03));
  NO2        o113(.A(ori_ori_n38_), .B(x3), .Y(ori_ori_n130_));
  NO2        o114(.A(ori_ori_n58_), .B(x6), .Y(ori_ori_n131_));
  AN2        o115(.A(ori_ori_n131_), .B(ori_ori_n44_), .Y(ori_ori_n132_));
  INV        o116(.A(ori_ori_n132_), .Y(ori_ori_n133_));
  NA2        o117(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n134_));
  NO3        o118(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n135_));
  NO2        o119(.A(ori_ori_n134_), .B(ori_ori_n111_), .Y(ori_ori_n136_));
  NO3        o120(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n137_));
  NO2        o121(.A(ori_ori_n137_), .B(ori_ori_n136_), .Y(ori_ori_n138_));
  INV        o122(.A(ori_ori_n138_), .Y(ori_ori_n139_));
  NA2        o123(.A(ori_ori_n139_), .B(ori_ori_n38_), .Y(ori_ori_n140_));
  NA2        o124(.A(ori_ori_n140_), .B(ori_ori_n133_), .Y(ori_ori_n141_));
  NO2        o125(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n142_));
  NO2        o126(.A(ori_ori_n142_), .B(x6), .Y(ori_ori_n143_));
  NOi21      o127(.An(ori_ori_n62_), .B(ori_ori_n143_), .Y(ori_ori_n144_));
  NA2        o128(.A(ori_ori_n50_), .B(ori_ori_n66_), .Y(ori_ori_n145_));
  NA3        o129(.A(ori_ori_n145_), .B(ori_ori_n142_), .C(x6), .Y(ori_ori_n146_));
  AOI210     o130(.A0(ori_ori_n146_), .A1(ori_ori_n144_), .B0(ori_ori_n100_), .Y(ori_ori_n147_));
  OR2        o131(.A(ori_ori_n147_), .B(ori_ori_n116_), .Y(ori_ori_n148_));
  NA2        o132(.A(ori_ori_n34_), .B(ori_ori_n43_), .Y(ori_ori_n149_));
  OAI210     o133(.A0(ori_ori_n149_), .A1(ori_ori_n22_), .B0(ori_ori_n112_), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n118_), .B(x6), .Y(ori_ori_n151_));
  NA2        o135(.A(ori_ori_n151_), .B(ori_ori_n150_), .Y(ori_ori_n152_));
  NA2        o136(.A(x6), .B(ori_ori_n38_), .Y(ori_ori_n153_));
  OAI210     o137(.A0(ori_ori_n78_), .A1(ori_ori_n59_), .B0(x4), .Y(ori_ori_n154_));
  AOI210     o138(.A0(ori_ori_n154_), .A1(ori_ori_n153_), .B0(ori_ori_n58_), .Y(ori_ori_n155_));
  NA2        o139(.A(x5), .B(ori_ori_n85_), .Y(ori_ori_n156_));
  NA3        o140(.A(ori_ori_n134_), .B(ori_ori_n83_), .C(x6), .Y(ori_ori_n157_));
  INV        o141(.A(ori_ori_n51_), .Y(ori_ori_n158_));
  NA3        o142(.A(ori_ori_n158_), .B(ori_ori_n157_), .C(ori_ori_n156_), .Y(ori_ori_n159_));
  OAI210     o143(.A0(ori_ori_n159_), .A1(ori_ori_n155_), .B0(x2), .Y(ori_ori_n160_));
  NA3        o144(.A(ori_ori_n160_), .B(ori_ori_n152_), .C(ori_ori_n148_), .Y(ori_ori_n161_));
  AOI210     o145(.A0(ori_ori_n141_), .A1(x8), .B0(ori_ori_n161_), .Y(ori_ori_n162_));
  NO2        o146(.A(ori_ori_n66_), .B(x3), .Y(ori_ori_n163_));
  NA2        o147(.A(ori_ori_n163_), .B(x6), .Y(ori_ori_n164_));
  NO2        o148(.A(ori_ori_n65_), .B(ori_ori_n22_), .Y(ori_ori_n165_));
  AOI210     o149(.A0(ori_ori_n143_), .A1(x5), .B0(ori_ori_n165_), .Y(ori_ori_n166_));
  AOI210     o150(.A0(ori_ori_n166_), .A1(ori_ori_n164_), .B0(x2), .Y(ori_ori_n167_));
  AOI220     o151(.A0(x6), .A1(ori_ori_n123_), .B0(x2), .B1(ori_ori_n51_), .Y(ori_ori_n168_));
  NA2        o152(.A(ori_ori_n134_), .B(x6), .Y(ori_ori_n169_));
  NO2        o153(.A(ori_ori_n134_), .B(x6), .Y(ori_ori_n170_));
  INV        o154(.A(ori_ori_n170_), .Y(ori_ori_n171_));
  NA3        o155(.A(ori_ori_n171_), .B(ori_ori_n169_), .C(ori_ori_n95_), .Y(ori_ori_n172_));
  NA3        o156(.A(ori_ori_n172_), .B(ori_ori_n168_), .C(ori_ori_n100_), .Y(ori_ori_n173_));
  AOI210     o157(.A0(x3), .A1(x2), .B0(ori_ori_n38_), .Y(ori_ori_n174_));
  NA2        o158(.A(ori_ori_n131_), .B(ori_ori_n33_), .Y(ori_ori_n175_));
  NO2        o159(.A(ori_ori_n175_), .B(x8), .Y(ori_ori_n176_));
  NO3        o160(.A(ori_ori_n176_), .B(ori_ori_n173_), .C(ori_ori_n167_), .Y(ori_ori_n177_));
  NA2        o161(.A(ori_ori_n170_), .B(x2), .Y(ori_ori_n178_));
  OAI210     o162(.A0(x0), .A1(x6), .B0(ori_ori_n35_), .Y(ori_ori_n179_));
  AOI210     o163(.A0(ori_ori_n179_), .A1(ori_ori_n178_), .B0(ori_ori_n122_), .Y(ori_ori_n180_));
  AOI210     o164(.A0(ori_ori_n30_), .A1(ori_ori_n43_), .B0(x0), .Y(ori_ori_n181_));
  NA3        o165(.A(ori_ori_n181_), .B(ori_ori_n103_), .C(ori_ori_n27_), .Y(ori_ori_n182_));
  NA2        o166(.A(x3), .B(x2), .Y(ori_ori_n183_));
  AOI210     o167(.A0(ori_ori_n183_), .A1(ori_ori_n149_), .B0(ori_ori_n182_), .Y(ori_ori_n184_));
  NAi21      o168(.An(x4), .B(x0), .Y(ori_ori_n185_));
  NO3        o169(.A(ori_ori_n185_), .B(ori_ori_n35_), .C(x2), .Y(ori_ori_n186_));
  NO2        o170(.A(ori_ori_n181_), .B(ori_ori_n281_), .Y(ori_ori_n187_));
  AOI220     o171(.A0(ori_ori_n187_), .A1(ori_ori_n61_), .B0(ori_ori_n18_), .B1(ori_ori_n26_), .Y(ori_ori_n188_));
  NO2        o172(.A(ori_ori_n188_), .B(ori_ori_n22_), .Y(ori_ori_n189_));
  NA3        o173(.A(ori_ori_n30_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n190_));
  INV        o174(.A(ori_ori_n181_), .Y(ori_ori_n191_));
  INV        o175(.A(ori_ori_n136_), .Y(ori_ori_n192_));
  NO2        o176(.A(ori_ori_n153_), .B(ori_ori_n192_), .Y(ori_ori_n193_));
  AO210      o177(.A0(ori_ori_n191_), .A1(ori_ori_n97_), .B0(ori_ori_n193_), .Y(ori_ori_n194_));
  NO4        o178(.A(ori_ori_n194_), .B(ori_ori_n189_), .C(ori_ori_n184_), .D(ori_ori_n180_), .Y(ori_ori_n195_));
  OAI210     o179(.A0(ori_ori_n177_), .A1(ori_ori_n162_), .B0(ori_ori_n195_), .Y(ori04));
  NA2        o180(.A(ori_ori_n43_), .B(ori_ori_n163_), .Y(ori_ori_n197_));
  NA2        o181(.A(x2), .B(ori_ori_n66_), .Y(ori_ori_n198_));
  NA3        o182(.A(ori_ori_n198_), .B(x6), .C(ori_ori_n197_), .Y(ori_ori_n199_));
  NA2        o183(.A(ori_ori_n199_), .B(x6), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n77_), .B(ori_ori_n73_), .Y(ori_ori_n201_));
  NA3        o185(.A(ori_ori_n201_), .B(x6), .C(x3), .Y(ori_ori_n202_));
  NO2        o186(.A(ori_ori_n280_), .B(ori_ori_n190_), .Y(ori_ori_n203_));
  INV        o187(.A(ori_ori_n203_), .Y(ori_ori_n204_));
  NA2        o188(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n205_));
  OAI210     o189(.A0(ori_ori_n73_), .A1(ori_ori_n17_), .B0(ori_ori_n205_), .Y(ori_ori_n206_));
  NA2        o190(.A(ori_ori_n206_), .B(ori_ori_n59_), .Y(ori_ori_n207_));
  NA3        o191(.A(ori_ori_n207_), .B(ori_ori_n204_), .C(ori_ori_n202_), .Y(ori_ori_n208_));
  OAI210     o192(.A0(x1), .A1(x3), .B0(ori_ori_n186_), .Y(ori_ori_n209_));
  NA2        o193(.A(ori_ori_n135_), .B(ori_ori_n62_), .Y(ori_ori_n210_));
  NA3        o194(.A(ori_ori_n210_), .B(ori_ori_n209_), .C(ori_ori_n100_), .Y(ori_ori_n211_));
  AOI210     o195(.A0(ori_ori_n208_), .A1(x4), .B0(ori_ori_n211_), .Y(ori_ori_n212_));
  NA3        o196(.A(ori_ori_n279_), .B(ori_ori_n285_), .C(ori_ori_n66_), .Y(ori_ori_n213_));
  XO2        o197(.A(x4), .B(x0), .Y(ori_ori_n214_));
  AOI210     o198(.A0(ori_ori_n282_), .A1(ori_ori_n213_), .B0(x3), .Y(ori_ori_n215_));
  INV        o199(.A(x4), .Y(ori_ori_n216_));
  NO2        o200(.A(ori_ori_n214_), .B(x2), .Y(ori_ori_n217_));
  INV        o201(.A(ori_ori_n217_), .Y(ori_ori_n218_));
  NA3        o202(.A(ori_ori_n218_), .B(ori_ori_n67_), .C(x6), .Y(ori_ori_n219_));
  NO2        o203(.A(ori_ori_n185_), .B(ori_ori_n65_), .Y(ori_ori_n220_));
  INV        o204(.A(ori_ori_n220_), .Y(ori_ori_n221_));
  NO2        o205(.A(ori_ori_n98_), .B(ori_ori_n60_), .Y(ori_ori_n222_));
  NO2        o206(.A(ori_ori_n29_), .B(x2), .Y(ori_ori_n223_));
  NOi21      o207(.An(ori_ori_n79_), .B(ori_ori_n23_), .Y(ori_ori_n224_));
  AOI210     o208(.A0(ori_ori_n223_), .A1(ori_ori_n222_), .B0(ori_ori_n224_), .Y(ori_ori_n225_));
  NA2        o209(.A(ori_ori_n221_), .B(ori_ori_n225_), .Y(ori_ori_n226_));
  OAI220     o210(.A0(ori_ori_n226_), .A1(x6), .B0(ori_ori_n219_), .B1(ori_ori_n215_), .Y(ori_ori_n227_));
  AO220      o211(.A0(x7), .A1(ori_ori_n227_), .B0(ori_ori_n212_), .B1(ori_ori_n200_), .Y(ori_ori_n228_));
  NA2        o212(.A(ori_ori_n223_), .B(x6), .Y(ori_ori_n229_));
  AOI210     o213(.A0(x6), .A1(x1), .B0(ori_ori_n99_), .Y(ori_ori_n230_));
  NA2        o214(.A(ori_ori_n216_), .B(x0), .Y(ori_ori_n231_));
  NA2        o215(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n232_));
  OAI210     o216(.A0(ori_ori_n231_), .A1(ori_ori_n230_), .B0(ori_ori_n232_), .Y(ori_ori_n233_));
  AOI220     o217(.A0(ori_ori_n233_), .A1(ori_ori_n229_), .B0(ori_ori_n137_), .B1(ori_ori_n39_), .Y(ori_ori_n234_));
  NA2        o218(.A(ori_ori_n234_), .B(ori_ori_n228_), .Y(ori_ori_n235_));
  NA2        o219(.A(ori_ori_n130_), .B(ori_ori_n100_), .Y(ori_ori_n236_));
  OAI210     o220(.A0(ori_ori_n24_), .A1(x1), .B0(ori_ori_n149_), .Y(ori_ori_n237_));
  NO2        o221(.A(ori_ori_n283_), .B(ori_ori_n285_), .Y(ori_ori_n238_));
  AOI210     o222(.A0(ori_ori_n237_), .A1(ori_ori_n78_), .B0(ori_ori_n238_), .Y(ori_ori_n239_));
  AOI210     o223(.A0(ori_ori_n239_), .A1(ori_ori_n236_), .B0(ori_ori_n22_), .Y(ori_ori_n240_));
  OAI210     o224(.A0(ori_ori_n284_), .A1(ori_ori_n240_), .B0(x6), .Y(ori_ori_n241_));
  NO2        o225(.A(x0), .B(ori_ori_n27_), .Y(ori_ori_n242_));
  NA2        o226(.A(ori_ori_n130_), .B(ori_ori_n100_), .Y(ori_ori_n243_));
  INV        o227(.A(x1), .Y(ori_ori_n244_));
  OAI210     o228(.A0(ori_ori_n243_), .A1(x8), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  NAi31      o229(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n246_));
  OAI210     o230(.A0(ori_ori_n246_), .A1(x4), .B0(ori_ori_n105_), .Y(ori_ori_n247_));
  NA2        o231(.A(ori_ori_n247_), .B(ori_ori_n96_), .Y(ori_ori_n248_));
  NA2        o232(.A(ori_ori_n222_), .B(ori_ori_n100_), .Y(ori_ori_n249_));
  NA3        o233(.A(ori_ori_n249_), .B(x1), .C(ori_ori_n248_), .Y(ori_ori_n250_));
  OAI210     o234(.A0(ori_ori_n245_), .A1(ori_ori_n242_), .B0(ori_ori_n250_), .Y(ori_ori_n251_));
  OAI210     o235(.A0(ori_ori_n185_), .A1(ori_ori_n34_), .B0(ori_ori_n214_), .Y(ori_ori_n252_));
  AOI220     o236(.A0(x7), .A1(ori_ori_n66_), .B0(ori_ori_n252_), .B1(ori_ori_n100_), .Y(ori_ori_n253_));
  NO2        o237(.A(ori_ori_n253_), .B(ori_ori_n43_), .Y(ori_ori_n254_));
  INV        o238(.A(ori_ori_n254_), .Y(ori_ori_n255_));
  AOI210     o239(.A0(ori_ori_n255_), .A1(ori_ori_n251_), .B0(ori_ori_n22_), .Y(ori_ori_n256_));
  NA3        o240(.A(ori_ori_n26_), .B(x2), .C(ori_ori_n17_), .Y(ori_ori_n257_));
  NO2        o241(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n258_));
  NA2        o242(.A(ori_ori_n258_), .B(ori_ori_n174_), .Y(ori_ori_n259_));
  INV        o243(.A(ori_ori_n259_), .Y(ori_ori_n260_));
  NO3        o244(.A(ori_ori_n280_), .B(ori_ori_n115_), .C(ori_ori_n31_), .Y(ori_ori_n261_));
  OAI210     o245(.A0(ori_ori_n261_), .A1(ori_ori_n260_), .B0(x7), .Y(ori_ori_n262_));
  NA2        o246(.A(ori_ori_n145_), .B(x7), .Y(ori_ori_n263_));
  NA3        o247(.A(ori_ori_n263_), .B(ori_ori_n99_), .C(ori_ori_n85_), .Y(ori_ori_n264_));
  NA3        o248(.A(ori_ori_n264_), .B(ori_ori_n262_), .C(ori_ori_n257_), .Y(ori_ori_n265_));
  OAI210     o249(.A0(ori_ori_n265_), .A1(ori_ori_n256_), .B0(ori_ori_n30_), .Y(ori_ori_n266_));
  NO4        o250(.A(x0), .B(ori_ori_n58_), .C(x4), .D(ori_ori_n43_), .Y(ori_ori_n267_));
  NA2        o251(.A(x3), .B(ori_ori_n43_), .Y(ori_ori_n268_));
  NO2        o252(.A(x3), .B(ori_ori_n43_), .Y(ori_ori_n269_));
  INV        o253(.A(ori_ori_n269_), .Y(ori_ori_n270_));
  OAI210     o254(.A0(ori_ori_n101_), .A1(ori_ori_n268_), .B0(ori_ori_n270_), .Y(ori_ori_n271_));
  NA2        o255(.A(ori_ori_n271_), .B(x0), .Y(ori_ori_n272_));
  NO2        o256(.A(ori_ori_n272_), .B(ori_ori_n153_), .Y(ori_ori_n273_));
  NO2        o257(.A(ori_ori_n273_), .B(ori_ori_n267_), .Y(ori_ori_n274_));
  NA3        o258(.A(ori_ori_n274_), .B(ori_ori_n266_), .C(ori_ori_n241_), .Y(ori_ori_n275_));
  AOI210     o259(.A0(ori_ori_n235_), .A1(ori_ori_n22_), .B0(ori_ori_n275_), .Y(ori05));
  INV        o260(.A(x2), .Y(ori_ori_n279_));
  INV        o261(.A(x2), .Y(ori_ori_n280_));
  INV        o262(.A(x6), .Y(ori_ori_n281_));
  INV        o263(.A(x4), .Y(ori_ori_n282_));
  INV        o264(.A(x4), .Y(ori_ori_n283_));
  INV        o265(.A(ori_ori_n40_), .Y(ori_ori_n284_));
  INV        o266(.A(x9), .Y(ori_ori_n285_));
  INV        o267(.A(ori_ori_n106_), .Y(ori_ori_n286_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NAi21      m005(.An(mai_mai_n20_), .B(mai_mai_n19_), .Y(mai_mai_n22_));
  NA2        m006(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n23_));
  INV        m007(.A(x5), .Y(mai_mai_n24_));
  NA2        m008(.A(x7), .B(x6), .Y(mai_mai_n25_));
  NA2        m009(.A(x8), .B(x3), .Y(mai_mai_n26_));
  NA2        m010(.A(x4), .B(x2), .Y(mai_mai_n27_));
  NO3        m011(.A(mai_mai_n27_), .B(mai_mai_n25_), .C(mai_mai_n24_), .Y(mai_mai_n28_));
  NO2        m012(.A(mai_mai_n28_), .B(mai_mai_n23_), .Y(mai_mai_n29_));
  NO2        m013(.A(x4), .B(x3), .Y(mai_mai_n30_));
  INV        m014(.A(mai_mai_n30_), .Y(mai_mai_n31_));
  OA210      m015(.A0(mai_mai_n31_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n32_));
  NOi31      m016(.An(mai_mai_n22_), .B(mai_mai_n32_), .C(mai_mai_n29_), .Y(mai00));
  NO2        m017(.A(x1), .B(x0), .Y(mai_mai_n34_));
  INV        m018(.A(x6), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n35_), .B(mai_mai_n24_), .Y(mai_mai_n36_));
  AN2        m020(.A(x8), .B(x7), .Y(mai_mai_n37_));
  NA2        m021(.A(mai_mai_n36_), .B(mai_mai_n34_), .Y(mai_mai_n38_));
  NA2        m022(.A(x4), .B(x3), .Y(mai_mai_n39_));
  AOI210     m023(.A0(mai_mai_n38_), .A1(mai_mai_n22_), .B0(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m024(.A(x2), .B(x0), .Y(mai_mai_n41_));
  INV        m025(.A(x3), .Y(mai_mai_n42_));
  NO2        m026(.A(mai_mai_n42_), .B(mai_mai_n18_), .Y(mai_mai_n43_));
  INV        m027(.A(mai_mai_n43_), .Y(mai_mai_n44_));
  NO2        m028(.A(mai_mai_n36_), .B(x4), .Y(mai_mai_n45_));
  OAI210     m029(.A0(mai_mai_n45_), .A1(mai_mai_n44_), .B0(mai_mai_n41_), .Y(mai_mai_n46_));
  INV        m030(.A(x4), .Y(mai_mai_n47_));
  NO2        m031(.A(mai_mai_n47_), .B(mai_mai_n17_), .Y(mai_mai_n48_));
  NA2        m032(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n49_));
  OAI210     m033(.A0(mai_mai_n49_), .A1(mai_mai_n20_), .B0(mai_mai_n46_), .Y(mai_mai_n50_));
  NA2        m034(.A(mai_mai_n20_), .B(mai_mai_n19_), .Y(mai_mai_n51_));
  INV        m035(.A(x2), .Y(mai_mai_n52_));
  NO2        m036(.A(mai_mai_n52_), .B(mai_mai_n17_), .Y(mai_mai_n53_));
  NA2        m037(.A(mai_mai_n42_), .B(mai_mai_n18_), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n54_), .B(mai_mai_n53_), .Y(mai_mai_n55_));
  OAI210     m039(.A0(mai_mai_n51_), .A1(mai_mai_n31_), .B0(mai_mai_n55_), .Y(mai_mai_n56_));
  NO3        m040(.A(mai_mai_n56_), .B(mai_mai_n50_), .C(mai_mai_n40_), .Y(mai01));
  NA2        m041(.A(x8), .B(x7), .Y(mai_mai_n58_));
  NA2        m042(.A(mai_mai_n42_), .B(x1), .Y(mai_mai_n59_));
  INV        m043(.A(x9), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n60_), .B(mai_mai_n35_), .Y(mai_mai_n61_));
  NO2        m045(.A(mai_mai_n59_), .B(mai_mai_n58_), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n59_), .B(x5), .Y(mai_mai_n63_));
  NO2        m047(.A(x8), .B(x2), .Y(mai_mai_n64_));
  INV        m048(.A(mai_mai_n64_), .Y(mai_mai_n65_));
  OAI210     m049(.A0(mai_mai_n54_), .A1(mai_mai_n20_), .B0(mai_mai_n42_), .Y(mai_mai_n66_));
  NAi21      m050(.An(x1), .B(x5), .Y(mai_mai_n67_));
  NO2        m051(.A(mai_mai_n66_), .B(mai_mai_n63_), .Y(mai_mai_n68_));
  OAI210     m052(.A0(mai_mai_n68_), .A1(mai_mai_n62_), .B0(x4), .Y(mai_mai_n69_));
  NA2        m053(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n70_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n71_));
  NA2        m055(.A(x5), .B(x3), .Y(mai_mai_n72_));
  NO2        m056(.A(x8), .B(x6), .Y(mai_mai_n73_));
  NO2        m057(.A(mai_mai_n72_), .B(mai_mai_n52_), .Y(mai_mai_n74_));
  NAi21      m058(.An(x4), .B(x3), .Y(mai_mai_n75_));
  INV        m059(.A(mai_mai_n75_), .Y(mai_mai_n76_));
  NO2        m060(.A(mai_mai_n76_), .B(mai_mai_n20_), .Y(mai_mai_n77_));
  NO2        m061(.A(x4), .B(x2), .Y(mai_mai_n78_));
  NO2        m062(.A(mai_mai_n78_), .B(x3), .Y(mai_mai_n79_));
  NO3        m063(.A(mai_mai_n79_), .B(mai_mai_n77_), .C(mai_mai_n18_), .Y(mai_mai_n80_));
  NO3        m064(.A(mai_mai_n80_), .B(mai_mai_n74_), .C(mai_mai_n71_), .Y(mai_mai_n81_));
  NA2        m065(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(mai_mai_n24_), .Y(mai_mai_n83_));
  INV        m067(.A(x8), .Y(mai_mai_n84_));
  NA2        m068(.A(x2), .B(x1), .Y(mai_mai_n85_));
  NO2        m069(.A(x2), .B(mai_mai_n83_), .Y(mai_mai_n86_));
  NO2        m070(.A(mai_mai_n86_), .B(mai_mai_n25_), .Y(mai_mai_n87_));
  OAI210     m071(.A0(mai_mai_n44_), .A1(mai_mai_n36_), .B0(mai_mai_n47_), .Y(mai_mai_n88_));
  NO2        m072(.A(mai_mai_n88_), .B(mai_mai_n87_), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n47_), .B(mai_mai_n52_), .Y(mai_mai_n90_));
  OAI210     m074(.A0(mai_mai_n90_), .A1(mai_mai_n42_), .B0(mai_mai_n18_), .Y(mai_mai_n91_));
  INV        m075(.A(mai_mai_n91_), .Y(mai_mai_n92_));
  NO2        m076(.A(x3), .B(x2), .Y(mai_mai_n93_));
  NA3        m077(.A(mai_mai_n93_), .B(mai_mai_n25_), .C(mai_mai_n24_), .Y(mai_mai_n94_));
  AOI210     m078(.A0(x8), .A1(x6), .B0(mai_mai_n94_), .Y(mai_mai_n95_));
  NA2        m079(.A(mai_mai_n52_), .B(x1), .Y(mai_mai_n96_));
  OAI210     m080(.A0(mai_mai_n96_), .A1(mai_mai_n39_), .B0(mai_mai_n17_), .Y(mai_mai_n97_));
  NO4        m081(.A(mai_mai_n97_), .B(mai_mai_n95_), .C(mai_mai_n92_), .D(mai_mai_n89_), .Y(mai_mai_n98_));
  AO210      m082(.A0(mai_mai_n81_), .A1(mai_mai_n69_), .B0(mai_mai_n98_), .Y(mai02));
  NO2        m083(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n100_));
  OAI210     m084(.A0(x4), .A1(x0), .B0(x3), .Y(mai_mai_n101_));
  NA2        m085(.A(mai_mai_n101_), .B(mai_mai_n100_), .Y(mai_mai_n102_));
  NO3        m086(.A(mai_mai_n102_), .B(x7), .C(x5), .Y(mai_mai_n103_));
  NA2        m087(.A(x9), .B(x2), .Y(mai_mai_n104_));
  OR2        m088(.A(x8), .B(x0), .Y(mai_mai_n105_));
  NAi21      m089(.An(x2), .B(x8), .Y(mai_mai_n106_));
  INV        m090(.A(mai_mai_n106_), .Y(mai_mai_n107_));
  NO2        m091(.A(x4), .B(x1), .Y(mai_mai_n108_));
  NO3        m092(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n109_));
  NOi21      m093(.An(x0), .B(x4), .Y(mai_mai_n110_));
  NAi21      m094(.An(x8), .B(x7), .Y(mai_mai_n111_));
  NO2        m095(.A(mai_mai_n111_), .B(mai_mai_n60_), .Y(mai_mai_n112_));
  NA2        m096(.A(mai_mai_n112_), .B(mai_mai_n110_), .Y(mai_mai_n113_));
  NO2        m097(.A(mai_mai_n113_), .B(mai_mai_n72_), .Y(mai_mai_n114_));
  NO2        m098(.A(x5), .B(mai_mai_n47_), .Y(mai_mai_n115_));
  INV        m099(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  NAi21      m100(.An(x0), .B(x4), .Y(mai_mai_n117_));
  NO2        m101(.A(mai_mai_n117_), .B(x1), .Y(mai_mai_n118_));
  NO2        m102(.A(x7), .B(x0), .Y(mai_mai_n119_));
  NO2        m103(.A(mai_mai_n78_), .B(mai_mai_n90_), .Y(mai_mai_n120_));
  NO2        m104(.A(mai_mai_n120_), .B(x3), .Y(mai_mai_n121_));
  OAI210     m105(.A0(mai_mai_n119_), .A1(mai_mai_n118_), .B0(mai_mai_n121_), .Y(mai_mai_n122_));
  NO2        m106(.A(mai_mai_n21_), .B(mai_mai_n42_), .Y(mai_mai_n123_));
  NA2        m107(.A(x5), .B(x0), .Y(mai_mai_n124_));
  NO2        m108(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n125_));
  NA2        m109(.A(mai_mai_n125_), .B(mai_mai_n123_), .Y(mai_mai_n126_));
  NA4        m110(.A(mai_mai_n126_), .B(mai_mai_n122_), .C(mai_mai_n116_), .D(mai_mai_n35_), .Y(mai_mai_n127_));
  NO3        m111(.A(mai_mai_n127_), .B(mai_mai_n114_), .C(mai_mai_n103_), .Y(mai_mai_n128_));
  NO3        m112(.A(mai_mai_n72_), .B(mai_mai_n70_), .C(mai_mai_n23_), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n27_), .B(mai_mai_n24_), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n27_), .B(mai_mai_n58_), .Y(mai_mai_n131_));
  NA2        m115(.A(x7), .B(x3), .Y(mai_mai_n132_));
  NO2        m116(.A(x9), .B(x7), .Y(mai_mai_n133_));
  NOi21      m117(.An(x8), .B(x0), .Y(mai_mai_n134_));
  AN2        m118(.A(x1), .B(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n42_), .B(x2), .Y(mai_mai_n136_));
  INV        m120(.A(x7), .Y(mai_mai_n137_));
  NA2        m121(.A(mai_mai_n137_), .B(mai_mai_n18_), .Y(mai_mai_n138_));
  NA2        m122(.A(mai_mai_n138_), .B(mai_mai_n136_), .Y(mai_mai_n139_));
  NO2        m123(.A(x4), .B(mai_mai_n139_), .Y(mai_mai_n140_));
  AOI210     m124(.A0(mai_mai_n135_), .A1(mai_mai_n42_), .B0(mai_mai_n140_), .Y(mai_mai_n141_));
  OAI210     m125(.A0(mai_mai_n132_), .A1(mai_mai_n49_), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  NA2        m126(.A(x5), .B(x1), .Y(mai_mai_n143_));
  INV        m127(.A(mai_mai_n143_), .Y(mai_mai_n144_));
  AOI210     m128(.A0(mai_mai_n144_), .A1(mai_mai_n110_), .B0(mai_mai_n35_), .Y(mai_mai_n145_));
  NO2        m129(.A(mai_mai_n60_), .B(mai_mai_n84_), .Y(mai_mai_n146_));
  NO2        m130(.A(x2), .B(mai_mai_n146_), .Y(mai_mai_n147_));
  NA2        m131(.A(mai_mai_n147_), .B(mai_mai_n63_), .Y(mai_mai_n148_));
  NAi31      m132(.An(mai_mai_n72_), .B(mai_mai_n37_), .C(mai_mai_n34_), .Y(mai_mai_n149_));
  NA2        m133(.A(mai_mai_n148_), .B(mai_mai_n145_), .Y(mai_mai_n150_));
  NO4        m134(.A(mai_mai_n150_), .B(mai_mai_n142_), .C(mai_mai_n131_), .D(mai_mai_n129_), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n151_), .B(mai_mai_n128_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n124_), .B(mai_mai_n120_), .Y(mai_mai_n153_));
  NA2        m137(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n154_));
  NO2        m138(.A(mai_mai_n137_), .B(mai_mai_n24_), .Y(mai_mai_n155_));
  NA2        m139(.A(x2), .B(x0), .Y(mai_mai_n156_));
  NA2        m140(.A(x4), .B(x1), .Y(mai_mai_n157_));
  NAi21      m141(.An(mai_mai_n108_), .B(mai_mai_n157_), .Y(mai_mai_n158_));
  NOi31      m142(.An(mai_mai_n158_), .B(x5), .C(mai_mai_n156_), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n159_), .B(mai_mai_n153_), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n160_), .B(mai_mai_n42_), .Y(mai_mai_n161_));
  INV        m145(.A(mai_mai_n70_), .Y(mai_mai_n162_));
  INV        m146(.A(mai_mai_n115_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n96_), .B(mai_mai_n17_), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n84_), .B(mai_mai_n164_), .Y(mai_mai_n165_));
  NO3        m149(.A(mai_mai_n165_), .B(mai_mai_n163_), .C(x7), .Y(mai_mai_n166_));
  NA3        m150(.A(mai_mai_n158_), .B(mai_mai_n163_), .C(mai_mai_n41_), .Y(mai_mai_n167_));
  INV        m151(.A(mai_mai_n167_), .Y(mai_mai_n168_));
  NO3        m152(.A(mai_mai_n168_), .B(mai_mai_n166_), .C(mai_mai_n162_), .Y(mai_mai_n169_));
  NO2        m153(.A(mai_mai_n169_), .B(x3), .Y(mai_mai_n170_));
  NO3        m154(.A(mai_mai_n170_), .B(mai_mai_n161_), .C(mai_mai_n152_), .Y(mai03));
  NO2        m155(.A(mai_mai_n47_), .B(x3), .Y(mai_mai_n172_));
  NO2        m156(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n52_), .B(x1), .Y(mai_mai_n174_));
  OAI210     m158(.A0(mai_mai_n174_), .A1(mai_mai_n24_), .B0(mai_mai_n61_), .Y(mai_mai_n175_));
  NO2        m159(.A(mai_mai_n175_), .B(mai_mai_n17_), .Y(mai_mai_n176_));
  NA2        m160(.A(mai_mai_n176_), .B(mai_mai_n172_), .Y(mai_mai_n177_));
  NA2        m161(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n178_));
  NO2        m162(.A(mai_mai_n178_), .B(x4), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n180_));
  NA2        m164(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n181_), .B(mai_mai_n178_), .Y(mai_mai_n182_));
  NA2        m166(.A(x9), .B(mai_mai_n52_), .Y(mai_mai_n183_));
  NA2        m167(.A(mai_mai_n183_), .B(x4), .Y(mai_mai_n184_));
  NA2        m168(.A(mai_mai_n178_), .B(mai_mai_n75_), .Y(mai_mai_n185_));
  AOI210     m169(.A0(mai_mai_n24_), .A1(x3), .B0(mai_mai_n156_), .Y(mai_mai_n186_));
  AOI220     m170(.A0(mai_mai_n186_), .A1(mai_mai_n185_), .B0(mai_mai_n184_), .B1(mai_mai_n182_), .Y(mai_mai_n187_));
  NO2        m171(.A(x5), .B(x1), .Y(mai_mai_n188_));
  AOI220     m172(.A0(mai_mai_n188_), .A1(mai_mai_n17_), .B0(mai_mai_n93_), .B1(x5), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n181_), .B(mai_mai_n154_), .Y(mai_mai_n190_));
  NA2        m174(.A(mai_mai_n370_), .B(mai_mai_n47_), .Y(mai_mai_n191_));
  NA3        m175(.A(mai_mai_n191_), .B(mai_mai_n187_), .C(mai_mai_n177_), .Y(mai_mai_n192_));
  NO2        m176(.A(mai_mai_n47_), .B(mai_mai_n42_), .Y(mai_mai_n193_));
  NA2        m177(.A(mai_mai_n193_), .B(mai_mai_n19_), .Y(mai_mai_n194_));
  NO2        m178(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n195_));
  AO210      m179(.A0(x7), .A1(mai_mai_n194_), .B0(mai_mai_n155_), .Y(mai_mai_n196_));
  NA2        m180(.A(mai_mai_n42_), .B(mai_mai_n52_), .Y(mai_mai_n197_));
  NA2        m181(.A(mai_mai_n125_), .B(mai_mai_n83_), .Y(mai_mai_n198_));
  NA2        m182(.A(x6), .B(mai_mai_n47_), .Y(mai_mai_n199_));
  NA2        m183(.A(mai_mai_n190_), .B(mai_mai_n369_), .Y(mai_mai_n200_));
  NA2        m184(.A(mai_mai_n173_), .B(mai_mai_n118_), .Y(mai_mai_n201_));
  OAI210     m185(.A0(mai_mai_n84_), .A1(mai_mai_n35_), .B0(mai_mai_n63_), .Y(mai_mai_n202_));
  NA3        m186(.A(mai_mai_n202_), .B(mai_mai_n201_), .C(mai_mai_n200_), .Y(mai_mai_n203_));
  NA2        m187(.A(mai_mai_n203_), .B(x2), .Y(mai_mai_n204_));
  NA3        m188(.A(mai_mai_n204_), .B(mai_mai_n198_), .C(mai_mai_n196_), .Y(mai_mai_n205_));
  AOI210     m189(.A0(mai_mai_n192_), .A1(x8), .B0(mai_mai_n205_), .Y(mai_mai_n206_));
  NO2        m190(.A(mai_mai_n84_), .B(x3), .Y(mai_mai_n207_));
  NA2        m191(.A(mai_mai_n207_), .B(mai_mai_n179_), .Y(mai_mai_n208_));
  NO3        m192(.A(mai_mai_n82_), .B(mai_mai_n73_), .C(mai_mai_n24_), .Y(mai_mai_n209_));
  INV        m193(.A(mai_mai_n209_), .Y(mai_mai_n210_));
  AOI210     m194(.A0(mai_mai_n210_), .A1(mai_mai_n208_), .B0(x2), .Y(mai_mai_n211_));
  NO2        m195(.A(x4), .B(mai_mai_n52_), .Y(mai_mai_n212_));
  AOI220     m196(.A0(mai_mai_n179_), .A1(mai_mai_n164_), .B0(mai_mai_n212_), .B1(mai_mai_n63_), .Y(mai_mai_n213_));
  NA2        m197(.A(mai_mai_n60_), .B(x6), .Y(mai_mai_n214_));
  NA3        m198(.A(mai_mai_n24_), .B(x3), .C(x2), .Y(mai_mai_n215_));
  AOI210     m199(.A0(mai_mai_n215_), .A1(mai_mai_n124_), .B0(mai_mai_n214_), .Y(mai_mai_n216_));
  NA2        m200(.A(mai_mai_n42_), .B(mai_mai_n17_), .Y(mai_mai_n217_));
  NO2        m201(.A(mai_mai_n217_), .B(mai_mai_n24_), .Y(mai_mai_n218_));
  OAI210     m202(.A0(mai_mai_n218_), .A1(mai_mai_n216_), .B0(mai_mai_n108_), .Y(mai_mai_n219_));
  NA2        m203(.A(mai_mai_n181_), .B(x6), .Y(mai_mai_n220_));
  NA2        m204(.A(mai_mai_n220_), .B(mai_mai_n130_), .Y(mai_mai_n221_));
  NA4        m205(.A(mai_mai_n221_), .B(mai_mai_n219_), .C(mai_mai_n213_), .D(mai_mai_n137_), .Y(mai_mai_n222_));
  NA2        m206(.A(mai_mai_n173_), .B(mai_mai_n195_), .Y(mai_mai_n223_));
  NO2        m207(.A(x9), .B(x6), .Y(mai_mai_n224_));
  NO2        m208(.A(mai_mai_n124_), .B(mai_mai_n18_), .Y(mai_mai_n225_));
  NAi21      m209(.An(x1), .B(x4), .Y(mai_mai_n226_));
  AOI210     m210(.A0(x3), .A1(x2), .B0(mai_mai_n47_), .Y(mai_mai_n227_));
  OAI210     m211(.A0(mai_mai_n124_), .A1(x3), .B0(mai_mai_n227_), .Y(mai_mai_n228_));
  AOI220     m212(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(mai_mai_n225_), .B1(mai_mai_n224_), .Y(mai_mai_n229_));
  NA2        m213(.A(mai_mai_n229_), .B(mai_mai_n223_), .Y(mai_mai_n230_));
  NO3        m214(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n231_));
  NA2        m215(.A(mai_mai_n96_), .B(mai_mai_n24_), .Y(mai_mai_n232_));
  NA2        m216(.A(x6), .B(x2), .Y(mai_mai_n233_));
  NO2        m217(.A(mai_mai_n233_), .B(mai_mai_n154_), .Y(mai_mai_n234_));
  AOI210     m218(.A0(mai_mai_n232_), .A1(mai_mai_n231_), .B0(mai_mai_n234_), .Y(mai_mai_n235_));
  OAI210     m219(.A0(mai_mai_n235_), .A1(mai_mai_n42_), .B0(mai_mai_n372_), .Y(mai_mai_n236_));
  OAI210     m220(.A0(mai_mai_n236_), .A1(mai_mai_n173_), .B0(mai_mai_n230_), .Y(mai_mai_n237_));
  NO2        m221(.A(x3), .B(mai_mai_n178_), .Y(mai_mai_n238_));
  NA2        m222(.A(x4), .B(x0), .Y(mai_mai_n239_));
  NA2        m223(.A(mai_mai_n238_), .B(mai_mai_n41_), .Y(mai_mai_n240_));
  AOI210     m224(.A0(mai_mai_n240_), .A1(mai_mai_n237_), .B0(x8), .Y(mai_mai_n241_));
  OAI210     m225(.A0(mai_mai_n225_), .A1(mai_mai_n188_), .B0(mai_mai_n60_), .Y(mai_mai_n242_));
  INV        m226(.A(mai_mai_n20_), .Y(mai_mai_n243_));
  AOI210     m227(.A0(mai_mai_n243_), .A1(mai_mai_n242_), .B0(mai_mai_n197_), .Y(mai_mai_n244_));
  NO4        m228(.A(mai_mai_n244_), .B(mai_mai_n241_), .C(mai_mai_n222_), .D(mai_mai_n211_), .Y(mai_mai_n245_));
  NO2        m229(.A(x3), .B(mai_mai_n35_), .Y(mai_mai_n246_));
  NA2        m230(.A(mai_mai_n246_), .B(x2), .Y(mai_mai_n247_));
  NO2        m231(.A(mai_mai_n247_), .B(mai_mai_n163_), .Y(mai_mai_n248_));
  NOi21      m232(.An(mai_mai_n233_), .B(mai_mai_n17_), .Y(mai_mai_n249_));
  NA2        m233(.A(mai_mai_n249_), .B(mai_mai_n188_), .Y(mai_mai_n250_));
  AOI210     m234(.A0(mai_mai_n35_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n251_));
  NA3        m235(.A(mai_mai_n251_), .B(mai_mai_n144_), .C(mai_mai_n31_), .Y(mai_mai_n252_));
  NA2        m236(.A(x3), .B(x2), .Y(mai_mai_n253_));
  AOI220     m237(.A0(mai_mai_n253_), .A1(mai_mai_n197_), .B0(mai_mai_n252_), .B1(mai_mai_n250_), .Y(mai_mai_n254_));
  NAi21      m238(.An(x4), .B(x0), .Y(mai_mai_n255_));
  NO3        m239(.A(mai_mai_n255_), .B(mai_mai_n43_), .C(x2), .Y(mai_mai_n256_));
  NA2        m240(.A(x6), .B(mai_mai_n256_), .Y(mai_mai_n257_));
  OAI210     m241(.A0(mai_mai_n251_), .A1(mai_mai_n249_), .B0(x6), .Y(mai_mai_n258_));
  NA2        m242(.A(mai_mai_n258_), .B(mai_mai_n76_), .Y(mai_mai_n259_));
  AOI210     m243(.A0(mai_mai_n259_), .A1(mai_mai_n257_), .B0(mai_mai_n24_), .Y(mai_mai_n260_));
  INV        m244(.A(mai_mai_n190_), .Y(mai_mai_n261_));
  NA2        m245(.A(mai_mai_n35_), .B(mai_mai_n42_), .Y(mai_mai_n262_));
  OR2        m246(.A(mai_mai_n262_), .B(mai_mai_n239_), .Y(mai_mai_n263_));
  OAI220     m247(.A0(mai_mai_n263_), .A1(mai_mai_n143_), .B0(mai_mai_n199_), .B1(mai_mai_n261_), .Y(mai_mai_n264_));
  NO4        m248(.A(mai_mai_n264_), .B(mai_mai_n260_), .C(mai_mai_n254_), .D(mai_mai_n248_), .Y(mai_mai_n265_));
  OAI210     m249(.A0(mai_mai_n245_), .A1(mai_mai_n206_), .B0(mai_mai_n265_), .Y(mai04));
  OAI210     m250(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n267_));
  NA3        m251(.A(mai_mai_n267_), .B(mai_mai_n231_), .C(mai_mai_n79_), .Y(mai_mai_n268_));
  NO2        m252(.A(x2), .B(x1), .Y(mai_mai_n269_));
  NO2        m253(.A(mai_mai_n269_), .B(mai_mai_n255_), .Y(mai_mai_n270_));
  NO2        m254(.A(x4), .B(x0), .Y(mai_mai_n271_));
  OAI210     m255(.A0(mai_mai_n271_), .A1(mai_mai_n270_), .B0(mai_mai_n207_), .Y(mai_mai_n272_));
  NA3        m256(.A(mai_mai_n82_), .B(x6), .C(mai_mai_n272_), .Y(mai_mai_n273_));
  NA2        m257(.A(mai_mai_n273_), .B(x6), .Y(mai_mai_n274_));
  NO2        m258(.A(mai_mai_n183_), .B(x3), .Y(mai_mai_n275_));
  NO3        m259(.A(mai_mai_n214_), .B(mai_mai_n106_), .C(mai_mai_n18_), .Y(mai_mai_n276_));
  NO2        m260(.A(mai_mai_n276_), .B(mai_mai_n275_), .Y(mai_mai_n277_));
  BUFFER     m261(.A(mai_mai_n134_), .Y(mai_mai_n278_));
  INV        m262(.A(mai_mai_n262_), .Y(mai_mai_n279_));
  AOI210     m263(.A0(mai_mai_n278_), .A1(mai_mai_n61_), .B0(mai_mai_n279_), .Y(mai_mai_n280_));
  NA2        m264(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n281_));
  NA3        m265(.A(mai_mai_n374_), .B(mai_mai_n280_), .C(mai_mai_n277_), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n100_), .A1(x3), .B0(mai_mai_n256_), .Y(mai_mai_n283_));
  NA2        m267(.A(mai_mai_n283_), .B(mai_mai_n137_), .Y(mai_mai_n284_));
  AOI210     m268(.A0(mai_mai_n282_), .A1(x4), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  XO2        m269(.A(x4), .B(x0), .Y(mai_mai_n286_));
  OAI210     m270(.A0(mai_mai_n286_), .A1(mai_mai_n104_), .B0(mai_mai_n226_), .Y(mai_mai_n287_));
  NA2        m271(.A(mai_mai_n287_), .B(x8), .Y(mai_mai_n288_));
  NO2        m272(.A(mai_mai_n288_), .B(x3), .Y(mai_mai_n289_));
  INV        m273(.A(mai_mai_n85_), .Y(mai_mai_n290_));
  NO2        m274(.A(mai_mai_n84_), .B(x4), .Y(mai_mai_n291_));
  AOI220     m275(.A0(mai_mai_n291_), .A1(mai_mai_n43_), .B0(mai_mai_n110_), .B1(mai_mai_n290_), .Y(mai_mai_n292_));
  NA4        m276(.A(mai_mai_n23_), .B(mai_mai_n292_), .C(mai_mai_n194_), .D(x6), .Y(mai_mai_n293_));
  NO2        m277(.A(mai_mai_n42_), .B(x0), .Y(mai_mai_n294_));
  NA2        m278(.A(x0), .B(mai_mai_n291_), .Y(mai_mai_n295_));
  NO2        m279(.A(mai_mai_n134_), .B(mai_mai_n75_), .Y(mai_mai_n296_));
  NA2        m280(.A(mai_mai_n376_), .B(mai_mai_n296_), .Y(mai_mai_n297_));
  NA2        m281(.A(mai_mai_n295_), .B(mai_mai_n297_), .Y(mai_mai_n298_));
  OAI220     m282(.A0(mai_mai_n298_), .A1(x6), .B0(mai_mai_n293_), .B1(mai_mai_n289_), .Y(mai_mai_n299_));
  INV        m283(.A(mai_mai_n41_), .Y(mai_mai_n300_));
  OAI210     m284(.A0(mai_mai_n300_), .A1(mai_mai_n84_), .B0(mai_mai_n263_), .Y(mai_mai_n301_));
  AOI210     m285(.A0(mai_mai_n301_), .A1(mai_mai_n18_), .B0(mai_mai_n137_), .Y(mai_mai_n302_));
  AO220      m286(.A0(mai_mai_n302_), .A1(mai_mai_n299_), .B0(mai_mai_n285_), .B1(mai_mai_n274_), .Y(mai_mai_n303_));
  NA2        m287(.A(mai_mai_n303_), .B(mai_mai_n268_), .Y(mai_mai_n304_));
  AOI210     m288(.A0(mai_mai_n174_), .A1(x8), .B0(mai_mai_n100_), .Y(mai_mai_n305_));
  NA2        m289(.A(mai_mai_n305_), .B(mai_mai_n281_), .Y(mai_mai_n306_));
  NA3        m290(.A(mai_mai_n306_), .B(mai_mai_n172_), .C(mai_mai_n137_), .Y(mai_mai_n307_));
  NA3        m291(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n308_));
  NO2        m292(.A(mai_mai_n308_), .B(mai_mai_n290_), .Y(mai_mai_n309_));
  INV        m293(.A(mai_mai_n309_), .Y(mai_mai_n310_));
  AOI210     m294(.A0(mai_mai_n310_), .A1(mai_mai_n307_), .B0(mai_mai_n24_), .Y(mai_mai_n311_));
  NA3        m295(.A(mai_mai_n107_), .B(mai_mai_n193_), .C(x0), .Y(mai_mai_n312_));
  OAI210     m296(.A0(mai_mai_n172_), .A1(mai_mai_n64_), .B0(mai_mai_n180_), .Y(mai_mai_n313_));
  NA3        m297(.A(mai_mai_n174_), .B(mai_mai_n195_), .C(x8), .Y(mai_mai_n314_));
  AOI210     m298(.A0(mai_mai_n314_), .A1(mai_mai_n313_), .B0(mai_mai_n24_), .Y(mai_mai_n315_));
  AOI210     m299(.A0(mai_mai_n106_), .A1(mai_mai_n105_), .B0(mai_mai_n41_), .Y(mai_mai_n316_));
  NOi31      m300(.An(mai_mai_n316_), .B(mai_mai_n294_), .C(mai_mai_n157_), .Y(mai_mai_n317_));
  OAI210     m301(.A0(mai_mai_n317_), .A1(mai_mai_n315_), .B0(mai_mai_n133_), .Y(mai_mai_n318_));
  NA2        m302(.A(mai_mai_n318_), .B(mai_mai_n312_), .Y(mai_mai_n319_));
  OAI210     m303(.A0(mai_mai_n319_), .A1(mai_mai_n311_), .B0(x6), .Y(mai_mai_n320_));
  INV        m304(.A(mai_mai_n119_), .Y(mai_mai_n321_));
  NA3        m305(.A(mai_mai_n53_), .B(mai_mai_n37_), .C(mai_mai_n30_), .Y(mai_mai_n322_));
  AOI220     m306(.A0(mai_mai_n322_), .A1(mai_mai_n321_), .B0(mai_mai_n39_), .B1(mai_mai_n31_), .Y(mai_mai_n323_));
  AOI220     m307(.A0(mai_mai_n373_), .A1(mai_mai_n193_), .B0(mai_mai_n172_), .B1(mai_mai_n137_), .Y(mai_mai_n324_));
  AOI210     m308(.A0(mai_mai_n112_), .A1(mai_mai_n212_), .B0(x1), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n324_), .A1(x8), .B0(mai_mai_n325_), .Y(mai_mai_n326_));
  NO4        m310(.A(mai_mai_n111_), .B(mai_mai_n255_), .C(x9), .D(x2), .Y(mai_mai_n327_));
  NOi21      m311(.An(mai_mai_n109_), .B(mai_mai_n156_), .Y(mai_mai_n328_));
  NO3        m312(.A(mai_mai_n328_), .B(mai_mai_n327_), .C(mai_mai_n18_), .Y(mai_mai_n329_));
  NA2        m313(.A(mai_mai_n296_), .B(mai_mai_n137_), .Y(mai_mai_n330_));
  NA3        m314(.A(mai_mai_n330_), .B(mai_mai_n329_), .C(mai_mai_n49_), .Y(mai_mai_n331_));
  OAI210     m315(.A0(mai_mai_n326_), .A1(mai_mai_n323_), .B0(mai_mai_n331_), .Y(mai_mai_n332_));
  NOi31      m316(.An(mai_mai_n373_), .B(mai_mai_n31_), .C(x8), .Y(mai_mai_n333_));
  AOI210     m317(.A0(mai_mai_n37_), .A1(x9), .B0(mai_mai_n117_), .Y(mai_mai_n334_));
  NO3        m318(.A(mai_mai_n334_), .B(mai_mai_n109_), .C(mai_mai_n42_), .Y(mai_mai_n335_));
  NO2        m319(.A(mai_mai_n226_), .B(x0), .Y(mai_mai_n336_));
  NO2        m320(.A(mai_mai_n336_), .B(x3), .Y(mai_mai_n337_));
  NO3        m321(.A(mai_mai_n337_), .B(mai_mai_n335_), .C(x2), .Y(mai_mai_n338_));
  NO2        m322(.A(mai_mai_n338_), .B(mai_mai_n333_), .Y(mai_mai_n339_));
  AOI210     m323(.A0(mai_mai_n339_), .A1(mai_mai_n332_), .B0(mai_mai_n24_), .Y(mai_mai_n340_));
  NA2        m324(.A(mai_mai_n371_), .B(mai_mai_n316_), .Y(mai_mai_n341_));
  NO2        m325(.A(mai_mai_n341_), .B(mai_mai_n93_), .Y(mai_mai_n342_));
  NA2        m326(.A(mai_mai_n342_), .B(x7), .Y(mai_mai_n343_));
  NA2        m327(.A(x9), .B(x7), .Y(mai_mai_n344_));
  NA3        m328(.A(mai_mai_n344_), .B(mai_mai_n136_), .C(mai_mai_n118_), .Y(mai_mai_n345_));
  NA2        m329(.A(mai_mai_n345_), .B(mai_mai_n343_), .Y(mai_mai_n346_));
  OAI210     m330(.A0(mai_mai_n346_), .A1(mai_mai_n340_), .B0(mai_mai_n35_), .Y(mai_mai_n347_));
  NA2        m331(.A(mai_mai_n217_), .B(mai_mai_n21_), .Y(mai_mai_n348_));
  NO2        m332(.A(mai_mai_n143_), .B(mai_mai_n119_), .Y(mai_mai_n349_));
  NA2        m333(.A(mai_mai_n349_), .B(mai_mai_n348_), .Y(mai_mai_n350_));
  AOI210     m334(.A0(mai_mai_n350_), .A1(mai_mai_n149_), .B0(mai_mai_n27_), .Y(mai_mai_n351_));
  AOI220     m335(.A0(mai_mai_n294_), .A1(mai_mai_n84_), .B0(mai_mai_n134_), .B1(mai_mai_n174_), .Y(mai_mai_n352_));
  NA2        m336(.A(mai_mai_n352_), .B(mai_mai_n82_), .Y(mai_mai_n353_));
  NA2        m337(.A(mai_mai_n353_), .B(mai_mai_n155_), .Y(mai_mai_n354_));
  OAI220     m338(.A0(x3), .A1(mai_mai_n65_), .B0(mai_mai_n143_), .B1(mai_mai_n42_), .Y(mai_mai_n355_));
  AOI210     m339(.A0(x2), .A1(mai_mai_n26_), .B0(mai_mai_n67_), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n133_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n357_));
  AOI210     m341(.A0(mai_mai_n375_), .A1(mai_mai_n357_), .B0(mai_mai_n356_), .Y(mai_mai_n358_));
  INV        m342(.A(mai_mai_n358_), .Y(mai_mai_n359_));
  AOI220     m343(.A0(mai_mai_n359_), .A1(x0), .B0(mai_mai_n355_), .B1(mai_mai_n119_), .Y(mai_mai_n360_));
  AOI210     m344(.A0(mai_mai_n360_), .A1(mai_mai_n354_), .B0(mai_mai_n199_), .Y(mai_mai_n361_));
  INV        m345(.A(x5), .Y(mai_mai_n362_));
  NO4        m346(.A(mai_mai_n96_), .B(mai_mai_n362_), .C(mai_mai_n58_), .D(mai_mai_n31_), .Y(mai_mai_n363_));
  NO3        m347(.A(mai_mai_n363_), .B(mai_mai_n361_), .C(mai_mai_n351_), .Y(mai_mai_n364_));
  NA3        m348(.A(mai_mai_n364_), .B(mai_mai_n347_), .C(mai_mai_n320_), .Y(mai_mai_n365_));
  AOI210     m349(.A0(mai_mai_n304_), .A1(mai_mai_n24_), .B0(mai_mai_n365_), .Y(mai05));
  INV        m350(.A(x6), .Y(mai_mai_n369_));
  INV        m351(.A(mai_mai_n189_), .Y(mai_mai_n370_));
  INV        m352(.A(x4), .Y(mai_mai_n371_));
  INV        m353(.A(x4), .Y(mai_mai_n372_));
  INV        m354(.A(x0), .Y(mai_mai_n373_));
  INV        m355(.A(mai_mai_n73_), .Y(mai_mai_n374_));
  INV        m356(.A(x1), .Y(mai_mai_n375_));
  INV        m357(.A(x2), .Y(mai_mai_n376_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x8), .B(x3), .Y(men_men_n26_));
  NA2        u010(.A(x4), .B(x2), .Y(men_men_n27_));
  NO2        u011(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n28_));
  NO2        u012(.A(men_men_n28_), .B(men_men_n24_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  NOi21      u015(.An(men_men_n23_), .B(men_men_n29_), .Y(men00));
  NO2        u016(.A(x1), .B(x0), .Y(men_men_n33_));
  INV        u017(.A(x6), .Y(men_men_n34_));
  NO2        u018(.A(men_men_n34_), .B(men_men_n25_), .Y(men_men_n35_));
  AN2        u019(.A(x8), .B(x7), .Y(men_men_n36_));
  NA2        u020(.A(men_men_n36_), .B(men_men_n33_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n23_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  NO2        u026(.A(men_men_n35_), .B(x4), .Y(men_men_n43_));
  NA2        u027(.A(men_men_n41_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u028(.A(x4), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n45_), .B(men_men_n17_), .Y(men_men_n46_));
  NA2        u030(.A(men_men_n46_), .B(x2), .Y(men_men_n47_));
  INV        u031(.A(men_men_n44_), .Y(men_men_n48_));
  NA2        u032(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n49_));
  AOI210     u033(.A0(men_men_n49_), .A1(men_men_n33_), .B0(men_men_n22_), .Y(men_men_n50_));
  INV        u034(.A(x2), .Y(men_men_n51_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n17_), .Y(men_men_n52_));
  NA2        u036(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n53_), .B(men_men_n52_), .Y(men_men_n54_));
  OAI210     u038(.A0(men_men_n50_), .A1(men_men_n31_), .B0(men_men_n54_), .Y(men_men_n55_));
  NO3        u039(.A(men_men_n55_), .B(men_men_n48_), .C(men_men_n39_), .Y(men01));
  NA2        u040(.A(x8), .B(x7), .Y(men_men_n57_));
  NA2        u041(.A(men_men_n41_), .B(x1), .Y(men_men_n58_));
  INV        u042(.A(x9), .Y(men_men_n59_));
  NO2        u043(.A(men_men_n59_), .B(men_men_n34_), .Y(men_men_n60_));
  INV        u044(.A(men_men_n60_), .Y(men_men_n61_));
  NO2        u045(.A(x7), .B(x6), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n58_), .B(x5), .Y(men_men_n63_));
  NO2        u047(.A(x8), .B(x2), .Y(men_men_n64_));
  OA210      u048(.A0(men_men_n64_), .A1(men_men_n63_), .B0(men_men_n62_), .Y(men_men_n65_));
  NA2        u049(.A(men_men_n25_), .B(men_men_n51_), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  NAi31      u051(.An(x1), .B(x9), .C(x5), .Y(men_men_n68_));
  OAI220     u052(.A0(men_men_n68_), .A1(men_men_n41_), .B0(men_men_n67_), .B1(men_men_n65_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n69_), .A1(men_men_n60_), .B0(x4), .Y(men_men_n70_));
  NA2        u054(.A(men_men_n45_), .B(x2), .Y(men_men_n71_));
  NA2        u055(.A(x5), .B(x3), .Y(men_men_n72_));
  NO2        u056(.A(x8), .B(x6), .Y(men_men_n73_));
  NO3        u057(.A(men_men_n73_), .B(men_men_n72_), .C(men_men_n62_), .Y(men_men_n74_));
  NAi21      u058(.An(x4), .B(x3), .Y(men_men_n75_));
  INV        u059(.A(men_men_n75_), .Y(men_men_n76_));
  NO2        u060(.A(men_men_n76_), .B(men_men_n22_), .Y(men_men_n77_));
  NO2        u061(.A(x4), .B(x2), .Y(men_men_n78_));
  NO2        u062(.A(men_men_n78_), .B(x3), .Y(men_men_n79_));
  NO3        u063(.A(men_men_n79_), .B(men_men_n77_), .C(men_men_n18_), .Y(men_men_n80_));
  NO3        u064(.A(men_men_n80_), .B(men_men_n74_), .C(men_men_n414_), .Y(men_men_n81_));
  NO3        u065(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .Y(men_men_n82_));
  NA2        u066(.A(men_men_n59_), .B(men_men_n45_), .Y(men_men_n83_));
  INV        u067(.A(men_men_n83_), .Y(men_men_n84_));
  OAI210     u068(.A0(men_men_n82_), .A1(men_men_n63_), .B0(men_men_n84_), .Y(men_men_n85_));
  NA2        u069(.A(x3), .B(men_men_n18_), .Y(men_men_n86_));
  NO2        u070(.A(men_men_n86_), .B(men_men_n25_), .Y(men_men_n87_));
  INV        u071(.A(x8), .Y(men_men_n88_));
  NA2        u072(.A(x2), .B(x1), .Y(men_men_n89_));
  NO2        u073(.A(men_men_n89_), .B(men_men_n88_), .Y(men_men_n90_));
  NO2        u074(.A(men_men_n90_), .B(men_men_n87_), .Y(men_men_n91_));
  INV        u075(.A(men_men_n91_), .Y(men_men_n92_));
  AOI210     u076(.A0(men_men_n53_), .A1(men_men_n25_), .B0(men_men_n51_), .Y(men_men_n93_));
  NO3        u077(.A(x4), .B(men_men_n93_), .C(men_men_n92_), .Y(men_men_n94_));
  NA2        u078(.A(x4), .B(men_men_n41_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n45_), .B(men_men_n51_), .Y(men_men_n96_));
  OAI210     u080(.A0(men_men_n96_), .A1(men_men_n41_), .B0(men_men_n18_), .Y(men_men_n97_));
  AOI210     u081(.A0(men_men_n95_), .A1(men_men_n49_), .B0(men_men_n97_), .Y(men_men_n98_));
  NO2        u082(.A(x3), .B(x2), .Y(men_men_n99_));
  NA2        u083(.A(men_men_n99_), .B(men_men_n25_), .Y(men_men_n100_));
  AOI210     u084(.A0(x8), .A1(x6), .B0(men_men_n100_), .Y(men_men_n101_));
  NA2        u085(.A(men_men_n51_), .B(x1), .Y(men_men_n102_));
  NO4        u086(.A(x0), .B(men_men_n101_), .C(men_men_n98_), .D(men_men_n94_), .Y(men_men_n103_));
  AO220      u087(.A0(men_men_n103_), .A1(men_men_n85_), .B0(men_men_n81_), .B1(men_men_n70_), .Y(men02));
  NO2        u088(.A(x3), .B(men_men_n51_), .Y(men_men_n105_));
  NA2        u089(.A(men_men_n41_), .B(x0), .Y(men_men_n106_));
  OAI210     u090(.A0(men_men_n83_), .A1(x2), .B0(men_men_n106_), .Y(men_men_n107_));
  NA2        u091(.A(men_men_n107_), .B(x1), .Y(men_men_n108_));
  NO3        u092(.A(men_men_n108_), .B(x7), .C(x5), .Y(men_men_n109_));
  NA2        u093(.A(x9), .B(x2), .Y(men_men_n110_));
  OR2        u094(.A(x8), .B(x0), .Y(men_men_n111_));
  INV        u095(.A(men_men_n111_), .Y(men_men_n112_));
  OAI210     u096(.A0(men_men_n110_), .A1(x7), .B0(men_men_n112_), .Y(men_men_n113_));
  NO2        u097(.A(x4), .B(x1), .Y(men_men_n114_));
  NA3        u098(.A(men_men_n114_), .B(men_men_n113_), .C(men_men_n57_), .Y(men_men_n115_));
  NOi21      u099(.An(x0), .B(x1), .Y(men_men_n116_));
  NO3        u100(.A(x9), .B(x8), .C(x7), .Y(men_men_n117_));
  NOi21      u101(.An(x0), .B(x4), .Y(men_men_n118_));
  NO2        u102(.A(x8), .B(men_men_n59_), .Y(men_men_n119_));
  NA2        u103(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n120_));
  AOI210     u104(.A0(men_men_n120_), .A1(men_men_n115_), .B0(men_men_n72_), .Y(men_men_n121_));
  NO2        u105(.A(x5), .B(men_men_n45_), .Y(men_men_n122_));
  NA2        u106(.A(x2), .B(men_men_n18_), .Y(men_men_n123_));
  AOI210     u107(.A0(men_men_n123_), .A1(men_men_n102_), .B0(men_men_n106_), .Y(men_men_n124_));
  OAI210     u108(.A0(men_men_n124_), .A1(men_men_n33_), .B0(men_men_n122_), .Y(men_men_n125_));
  NO2        u109(.A(x7), .B(x0), .Y(men_men_n126_));
  NO2        u110(.A(men_men_n78_), .B(men_men_n96_), .Y(men_men_n127_));
  NO2        u111(.A(men_men_n21_), .B(men_men_n41_), .Y(men_men_n128_));
  NA2        u112(.A(x5), .B(x0), .Y(men_men_n129_));
  NO2        u113(.A(men_men_n45_), .B(x2), .Y(men_men_n130_));
  NA3        u114(.A(men_men_n130_), .B(men_men_n129_), .C(men_men_n128_), .Y(men_men_n131_));
  NA3        u115(.A(men_men_n131_), .B(men_men_n125_), .C(men_men_n34_), .Y(men_men_n132_));
  NO3        u116(.A(men_men_n132_), .B(men_men_n121_), .C(men_men_n109_), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n27_), .B(men_men_n25_), .Y(men_men_n134_));
  AOI220     u118(.A0(men_men_n116_), .A1(men_men_n134_), .B0(men_men_n63_), .B1(men_men_n17_), .Y(men_men_n135_));
  NO3        u119(.A(men_men_n135_), .B(men_men_n57_), .C(men_men_n59_), .Y(men_men_n136_));
  NA2        u120(.A(x7), .B(x3), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n95_), .B(x5), .Y(men_men_n138_));
  NO2        u122(.A(x9), .B(x7), .Y(men_men_n139_));
  NOi21      u123(.An(x8), .B(x0), .Y(men_men_n140_));
  OA210      u124(.A0(men_men_n139_), .A1(x1), .B0(men_men_n140_), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n41_), .B(x2), .Y(men_men_n142_));
  INV        u126(.A(x7), .Y(men_men_n143_));
  AOI210     u127(.A0(men_men_n105_), .A1(men_men_n36_), .B0(men_men_n142_), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n25_), .B(x4), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n145_), .B(men_men_n118_), .Y(men_men_n146_));
  NO2        u130(.A(men_men_n146_), .B(men_men_n144_), .Y(men_men_n147_));
  AOI210     u131(.A0(men_men_n141_), .A1(men_men_n138_), .B0(men_men_n147_), .Y(men_men_n148_));
  OAI210     u132(.A0(men_men_n137_), .A1(men_men_n47_), .B0(men_men_n148_), .Y(men_men_n149_));
  NA2        u133(.A(x5), .B(x1), .Y(men_men_n150_));
  NO2        u134(.A(men_men_n59_), .B(men_men_n88_), .Y(men_men_n151_));
  NAi21      u135(.An(x2), .B(x7), .Y(men_men_n152_));
  NAi31      u136(.An(men_men_n72_), .B(men_men_n36_), .C(men_men_n33_), .Y(men_men_n153_));
  NA2        u137(.A(men_men_n153_), .B(x6), .Y(men_men_n154_));
  NO3        u138(.A(men_men_n154_), .B(men_men_n149_), .C(men_men_n136_), .Y(men_men_n155_));
  NO2        u139(.A(men_men_n155_), .B(men_men_n133_), .Y(men_men_n156_));
  NA2        u140(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n157_));
  NA2        u141(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n158_));
  NA3        u142(.A(men_men_n158_), .B(men_men_n157_), .C(men_men_n24_), .Y(men_men_n159_));
  AN2        u143(.A(men_men_n159_), .B(men_men_n130_), .Y(men_men_n160_));
  NA2        u144(.A(x8), .B(x0), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n143_), .B(men_men_n25_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n116_), .B(x4), .Y(men_men_n163_));
  NA2        u147(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  INV        u148(.A(men_men_n164_), .Y(men_men_n165_));
  NA2        u149(.A(x2), .B(x0), .Y(men_men_n166_));
  NA2        u150(.A(x4), .B(x1), .Y(men_men_n167_));
  NAi21      u151(.An(men_men_n114_), .B(men_men_n167_), .Y(men_men_n168_));
  NOi31      u152(.An(men_men_n168_), .B(men_men_n145_), .C(men_men_n166_), .Y(men_men_n169_));
  NO3        u153(.A(men_men_n169_), .B(men_men_n165_), .C(men_men_n160_), .Y(men_men_n170_));
  NO2        u154(.A(men_men_n170_), .B(men_men_n41_), .Y(men_men_n171_));
  NO2        u155(.A(men_men_n159_), .B(men_men_n71_), .Y(men_men_n172_));
  INV        u156(.A(men_men_n122_), .Y(men_men_n173_));
  NA3        u157(.A(men_men_n168_), .B(men_men_n173_), .C(men_men_n40_), .Y(men_men_n174_));
  OAI210     u158(.A0(men_men_n158_), .A1(men_men_n127_), .B0(men_men_n174_), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n175_), .B(men_men_n172_), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n176_), .B(x3), .Y(men_men_n177_));
  NO3        u161(.A(men_men_n177_), .B(men_men_n171_), .C(men_men_n156_), .Y(men03));
  NO2        u162(.A(men_men_n51_), .B(x1), .Y(men_men_n179_));
  INV        u163(.A(men_men_n60_), .Y(men_men_n180_));
  OAI220     u164(.A0(men_men_n180_), .A1(men_men_n17_), .B0(men_men_n25_), .B1(men_men_n102_), .Y(men_men_n181_));
  NA2        u165(.A(men_men_n181_), .B(x4), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n72_), .B(x6), .Y(men_men_n183_));
  NA2        u167(.A(x6), .B(men_men_n25_), .Y(men_men_n184_));
  NO2        u168(.A(men_men_n18_), .B(x0), .Y(men_men_n185_));
  AO220      u169(.A0(men_men_n185_), .A1(men_men_n25_), .B0(men_men_n183_), .B1(men_men_n52_), .Y(men_men_n186_));
  NA2        u170(.A(men_men_n186_), .B(men_men_n59_), .Y(men_men_n187_));
  NA2        u171(.A(x3), .B(men_men_n17_), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n188_), .B(men_men_n184_), .Y(men_men_n189_));
  NA2        u173(.A(men_men_n184_), .B(men_men_n75_), .Y(men_men_n190_));
  AOI210     u174(.A0(men_men_n25_), .A1(x3), .B0(men_men_n166_), .Y(men_men_n191_));
  AOI210     u175(.A0(men_men_n191_), .A1(men_men_n190_), .B0(men_men_n189_), .Y(men_men_n192_));
  NO2        u176(.A(x5), .B(x1), .Y(men_men_n193_));
  AOI220     u177(.A0(men_men_n193_), .A1(men_men_n17_), .B0(men_men_n99_), .B1(x5), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n188_), .B(men_men_n157_), .Y(men_men_n195_));
  NO2        u179(.A(men_men_n194_), .B(men_men_n61_), .Y(men_men_n196_));
  INV        u180(.A(men_men_n196_), .Y(men_men_n197_));
  NA4        u181(.A(men_men_n197_), .B(men_men_n192_), .C(men_men_n187_), .D(men_men_n182_), .Y(men_men_n198_));
  NO2        u182(.A(x3), .B(men_men_n17_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n199_), .B(x6), .Y(men_men_n200_));
  NA2        u184(.A(men_men_n59_), .B(men_men_n88_), .Y(men_men_n201_));
  NO2        u185(.A(men_men_n78_), .B(men_men_n143_), .Y(men_men_n202_));
  OR2        u186(.A(men_men_n202_), .B(men_men_n162_), .Y(men_men_n203_));
  NA2        u187(.A(men_men_n41_), .B(men_men_n51_), .Y(men_men_n204_));
  NO3        u188(.A(men_men_n167_), .B(men_men_n59_), .C(x6), .Y(men_men_n205_));
  AOI220     u189(.A0(men_men_n205_), .A1(men_men_n17_), .B0(men_men_n130_), .B1(men_men_n87_), .Y(men_men_n206_));
  NA2        u190(.A(x6), .B(men_men_n45_), .Y(men_men_n207_));
  OAI210     u191(.A0(men_men_n112_), .A1(men_men_n73_), .B0(x4), .Y(men_men_n208_));
  AOI210     u192(.A0(men_men_n208_), .A1(men_men_n207_), .B0(men_men_n72_), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n150_), .B(men_men_n41_), .Y(men_men_n210_));
  OAI210     u194(.A0(men_men_n210_), .A1(men_men_n195_), .B0(x9), .Y(men_men_n211_));
  NA2        u195(.A(men_men_n122_), .B(x6), .Y(men_men_n212_));
  NA2        u196(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n213_));
  OAI210     u197(.A0(men_men_n213_), .A1(men_men_n209_), .B0(x2), .Y(men_men_n214_));
  NA3        u198(.A(men_men_n214_), .B(men_men_n206_), .C(men_men_n203_), .Y(men_men_n215_));
  AOI210     u199(.A0(men_men_n198_), .A1(x8), .B0(men_men_n215_), .Y(men_men_n216_));
  NA2        u200(.A(men_men_n200_), .B(men_men_n145_), .Y(men_men_n217_));
  NO2        u201(.A(men_men_n217_), .B(x2), .Y(men_men_n218_));
  NA2        u202(.A(men_men_n59_), .B(x6), .Y(men_men_n219_));
  NA3        u203(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n220_));
  INV        u204(.A(men_men_n219_), .Y(men_men_n221_));
  NA2        u205(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n222_));
  NA2        u206(.A(men_men_n221_), .B(men_men_n114_), .Y(men_men_n223_));
  NO2        u207(.A(men_men_n188_), .B(x6), .Y(men_men_n224_));
  NA2        u208(.A(men_men_n151_), .B(men_men_n134_), .Y(men_men_n225_));
  NA3        u209(.A(men_men_n225_), .B(men_men_n223_), .C(men_men_n143_), .Y(men_men_n226_));
  NA2        u210(.A(x5), .B(men_men_n199_), .Y(men_men_n227_));
  NO2        u211(.A(x9), .B(x6), .Y(men_men_n228_));
  NO2        u212(.A(men_men_n129_), .B(men_men_n18_), .Y(men_men_n229_));
  NAi21      u213(.An(men_men_n229_), .B(men_men_n220_), .Y(men_men_n230_));
  NAi21      u214(.An(x1), .B(x4), .Y(men_men_n231_));
  AOI210     u215(.A0(x3), .A1(x2), .B0(men_men_n45_), .Y(men_men_n232_));
  OAI210     u216(.A0(men_men_n129_), .A1(x3), .B0(men_men_n232_), .Y(men_men_n233_));
  AOI220     u217(.A0(men_men_n233_), .A1(men_men_n231_), .B0(men_men_n230_), .B1(men_men_n228_), .Y(men_men_n234_));
  NA2        u218(.A(men_men_n234_), .B(men_men_n227_), .Y(men_men_n235_));
  NA2        u219(.A(men_men_n59_), .B(x2), .Y(men_men_n236_));
  NO2        u220(.A(men_men_n236_), .B(men_men_n227_), .Y(men_men_n237_));
  NO3        u221(.A(x9), .B(x6), .C(x0), .Y(men_men_n238_));
  INV        u222(.A(men_men_n238_), .Y(men_men_n239_));
  OAI220     u223(.A0(men_men_n239_), .A1(men_men_n41_), .B0(men_men_n163_), .B1(men_men_n43_), .Y(men_men_n240_));
  OAI210     u224(.A0(men_men_n240_), .A1(men_men_n237_), .B0(men_men_n235_), .Y(men_men_n241_));
  NO2        u225(.A(men_men_n411_), .B(men_men_n184_), .Y(men_men_n242_));
  OR3        u226(.A(men_men_n242_), .B(men_men_n183_), .C(men_men_n138_), .Y(men_men_n243_));
  NA2        u227(.A(x4), .B(x0), .Y(men_men_n244_));
  NO3        u228(.A(men_men_n68_), .B(men_men_n244_), .C(x6), .Y(men_men_n245_));
  AOI210     u229(.A0(men_men_n243_), .A1(men_men_n40_), .B0(men_men_n245_), .Y(men_men_n246_));
  AOI210     u230(.A0(men_men_n246_), .A1(men_men_n241_), .B0(x8), .Y(men_men_n247_));
  INV        u231(.A(men_men_n219_), .Y(men_men_n248_));
  OAI210     u232(.A0(men_men_n229_), .A1(men_men_n193_), .B0(men_men_n248_), .Y(men_men_n249_));
  INV        u233(.A(men_men_n161_), .Y(men_men_n250_));
  OAI210     u234(.A0(men_men_n250_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n251_));
  AOI210     u235(.A0(men_men_n251_), .A1(men_men_n249_), .B0(men_men_n204_), .Y(men_men_n252_));
  NO4        u236(.A(men_men_n252_), .B(men_men_n247_), .C(men_men_n226_), .D(men_men_n218_), .Y(men_men_n253_));
  NO2        u237(.A(men_men_n151_), .B(x1), .Y(men_men_n254_));
  NO3        u238(.A(men_men_n254_), .B(x3), .C(men_men_n34_), .Y(men_men_n255_));
  OAI210     u239(.A0(men_men_n255_), .A1(men_men_n224_), .B0(x2), .Y(men_men_n256_));
  OAI210     u240(.A0(men_men_n250_), .A1(x6), .B0(men_men_n42_), .Y(men_men_n257_));
  AOI210     u241(.A0(men_men_n257_), .A1(men_men_n256_), .B0(men_men_n173_), .Y(men_men_n258_));
  NA3        u242(.A(x0), .B(men_men_n193_), .C(men_men_n38_), .Y(men_men_n259_));
  AOI210     u243(.A0(men_men_n34_), .A1(men_men_n51_), .B0(x0), .Y(men_men_n260_));
  NA2        u244(.A(x3), .B(x2), .Y(men_men_n261_));
  AOI210     u245(.A0(men_men_n261_), .A1(men_men_n204_), .B0(men_men_n259_), .Y(men_men_n262_));
  NAi21      u246(.An(x4), .B(x0), .Y(men_men_n263_));
  NO3        u247(.A(men_men_n263_), .B(men_men_n42_), .C(x2), .Y(men_men_n264_));
  OAI210     u248(.A0(x6), .A1(men_men_n18_), .B0(men_men_n264_), .Y(men_men_n265_));
  OAI220     u249(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n266_));
  NO2        u250(.A(x9), .B(x8), .Y(men_men_n267_));
  NA3        u251(.A(men_men_n267_), .B(men_men_n34_), .C(men_men_n51_), .Y(men_men_n268_));
  OAI210     u252(.A0(men_men_n260_), .A1(x0), .B0(men_men_n268_), .Y(men_men_n269_));
  AOI220     u253(.A0(men_men_n269_), .A1(men_men_n76_), .B0(men_men_n266_), .B1(men_men_n30_), .Y(men_men_n270_));
  AOI210     u254(.A0(men_men_n270_), .A1(men_men_n265_), .B0(men_men_n25_), .Y(men_men_n271_));
  NA3        u255(.A(men_men_n34_), .B(x1), .C(men_men_n17_), .Y(men_men_n272_));
  OAI210     u256(.A0(men_men_n260_), .A1(x0), .B0(men_men_n272_), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n34_), .B(men_men_n41_), .Y(men_men_n274_));
  OR2        u258(.A(men_men_n274_), .B(men_men_n244_), .Y(men_men_n275_));
  NO2        u259(.A(men_men_n275_), .B(men_men_n150_), .Y(men_men_n276_));
  AO210      u260(.A0(men_men_n273_), .A1(men_men_n138_), .B0(men_men_n276_), .Y(men_men_n277_));
  NO4        u261(.A(men_men_n277_), .B(men_men_n271_), .C(men_men_n262_), .D(men_men_n258_), .Y(men_men_n278_));
  OAI210     u262(.A0(men_men_n253_), .A1(men_men_n216_), .B0(men_men_n278_), .Y(men04));
  OAI210     u263(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n280_));
  NA3        u264(.A(men_men_n280_), .B(men_men_n238_), .C(men_men_n79_), .Y(men_men_n281_));
  NO2        u265(.A(x2), .B(x1), .Y(men_men_n282_));
  OAI210     u266(.A0(men_men_n222_), .A1(men_men_n282_), .B0(men_men_n34_), .Y(men_men_n283_));
  NO2        u267(.A(men_men_n282_), .B(men_men_n263_), .Y(men_men_n284_));
  NO2        u268(.A(men_men_n236_), .B(men_men_n86_), .Y(men_men_n285_));
  NO2        u269(.A(men_men_n285_), .B(men_men_n34_), .Y(men_men_n286_));
  NO2        u270(.A(men_men_n261_), .B(men_men_n185_), .Y(men_men_n287_));
  NA2        u271(.A(x9), .B(x0), .Y(men_men_n288_));
  AOI210     u272(.A0(men_men_n86_), .A1(men_men_n71_), .B0(men_men_n288_), .Y(men_men_n289_));
  OAI210     u273(.A0(men_men_n289_), .A1(men_men_n287_), .B0(men_men_n88_), .Y(men_men_n290_));
  NA2        u274(.A(men_men_n290_), .B(men_men_n286_), .Y(men_men_n291_));
  NA2        u275(.A(men_men_n291_), .B(men_men_n283_), .Y(men_men_n292_));
  NO2        u276(.A(x2), .B(men_men_n106_), .Y(men_men_n293_));
  NO3        u277(.A(men_men_n219_), .B(x2), .C(men_men_n18_), .Y(men_men_n294_));
  NO2        u278(.A(men_men_n294_), .B(men_men_n293_), .Y(men_men_n295_));
  OAI210     u279(.A0(men_men_n111_), .A1(men_men_n102_), .B0(men_men_n161_), .Y(men_men_n296_));
  NA3        u280(.A(men_men_n296_), .B(x6), .C(x3), .Y(men_men_n297_));
  NOi21      u281(.An(men_men_n140_), .B(men_men_n123_), .Y(men_men_n298_));
  AOI210     u282(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n299_));
  OAI220     u283(.A0(men_men_n299_), .A1(men_men_n274_), .B0(men_men_n236_), .B1(men_men_n272_), .Y(men_men_n300_));
  AOI210     u284(.A0(men_men_n298_), .A1(men_men_n60_), .B0(men_men_n300_), .Y(men_men_n301_));
  NA2        u285(.A(men_men_n285_), .B(men_men_n88_), .Y(men_men_n302_));
  NA4        u286(.A(men_men_n302_), .B(men_men_n301_), .C(men_men_n297_), .D(men_men_n295_), .Y(men_men_n303_));
  NA3        u287(.A(men_men_n201_), .B(men_men_n412_), .C(men_men_n78_), .Y(men_men_n304_));
  NA2        u288(.A(men_men_n304_), .B(men_men_n143_), .Y(men_men_n305_));
  AOI210     u289(.A0(men_men_n303_), .A1(x4), .B0(men_men_n305_), .Y(men_men_n306_));
  NA2        u290(.A(men_men_n284_), .B(men_men_n88_), .Y(men_men_n307_));
  NOi21      u291(.An(x4), .B(x0), .Y(men_men_n308_));
  XO2        u292(.A(x4), .B(x0), .Y(men_men_n309_));
  OAI210     u293(.A0(men_men_n309_), .A1(men_men_n110_), .B0(men_men_n231_), .Y(men_men_n310_));
  AOI220     u294(.A0(men_men_n310_), .A1(x8), .B0(men_men_n308_), .B1(men_men_n89_), .Y(men_men_n311_));
  AOI210     u295(.A0(men_men_n311_), .A1(men_men_n307_), .B0(x3), .Y(men_men_n312_));
  NO2        u296(.A(men_men_n88_), .B(x4), .Y(men_men_n313_));
  NO3        u297(.A(men_men_n309_), .B(men_men_n151_), .C(x2), .Y(men_men_n314_));
  NO3        u298(.A(men_men_n201_), .B(men_men_n27_), .C(men_men_n24_), .Y(men_men_n315_));
  NO2        u299(.A(men_men_n315_), .B(men_men_n314_), .Y(men_men_n316_));
  NA2        u300(.A(men_men_n316_), .B(x6), .Y(men_men_n317_));
  OR2        u301(.A(men_men_n313_), .B(x3), .Y(men_men_n318_));
  NO2        u302(.A(men_men_n140_), .B(men_men_n102_), .Y(men_men_n319_));
  AOI220     u303(.A0(men_men_n319_), .A1(men_men_n318_), .B0(men_men_n410_), .B1(men_men_n58_), .Y(men_men_n320_));
  NOi21      u304(.An(men_men_n114_), .B(men_men_n26_), .Y(men_men_n321_));
  INV        u305(.A(men_men_n321_), .Y(men_men_n322_));
  OAI210     u306(.A0(men_men_n320_), .A1(men_men_n59_), .B0(men_men_n322_), .Y(men_men_n323_));
  OAI220     u307(.A0(men_men_n323_), .A1(x6), .B0(men_men_n317_), .B1(men_men_n312_), .Y(men_men_n324_));
  OAI210     u308(.A0(men_men_n60_), .A1(men_men_n45_), .B0(men_men_n40_), .Y(men_men_n325_));
  OAI210     u309(.A0(men_men_n325_), .A1(men_men_n88_), .B0(men_men_n275_), .Y(men_men_n326_));
  AOI210     u310(.A0(men_men_n326_), .A1(men_men_n18_), .B0(men_men_n143_), .Y(men_men_n327_));
  AO220      u311(.A0(men_men_n327_), .A1(men_men_n324_), .B0(men_men_n306_), .B1(men_men_n292_), .Y(men_men_n328_));
  AOI210     u312(.A0(x6), .A1(x1), .B0(men_men_n142_), .Y(men_men_n329_));
  NA2        u313(.A(men_men_n313_), .B(x0), .Y(men_men_n330_));
  NO2        u314(.A(men_men_n330_), .B(men_men_n329_), .Y(men_men_n331_));
  INV        u315(.A(men_men_n331_), .Y(men_men_n332_));
  NA3        u316(.A(men_men_n332_), .B(men_men_n328_), .C(men_men_n281_), .Y(men_men_n333_));
  AO220      u317(.A0(x4), .A1(men_men_n139_), .B0(men_men_n105_), .B1(x4), .Y(men_men_n334_));
  NA3        u318(.A(x7), .B(x3), .C(x0), .Y(men_men_n335_));
  NA2        u319(.A(x3), .B(x0), .Y(men_men_n336_));
  NO2        u320(.A(men_men_n336_), .B(x2), .Y(men_men_n337_));
  AOI210     u321(.A0(men_men_n334_), .A1(men_men_n112_), .B0(men_men_n337_), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n338_), .B(men_men_n25_), .Y(men_men_n339_));
  OAI210     u323(.A0(x4), .A1(men_men_n64_), .B0(men_men_n185_), .Y(men_men_n340_));
  NA3        u324(.A(men_men_n179_), .B(men_men_n199_), .C(x8), .Y(men_men_n341_));
  AOI210     u325(.A0(men_men_n341_), .A1(men_men_n340_), .B0(men_men_n25_), .Y(men_men_n342_));
  AOI210     u326(.A0(x2), .A1(men_men_n111_), .B0(men_men_n40_), .Y(men_men_n343_));
  NOi31      u327(.An(men_men_n343_), .B(x3), .C(men_men_n167_), .Y(men_men_n344_));
  OAI210     u328(.A0(men_men_n344_), .A1(men_men_n342_), .B0(men_men_n139_), .Y(men_men_n345_));
  NAi31      u329(.An(men_men_n47_), .B(men_men_n254_), .C(men_men_n162_), .Y(men_men_n346_));
  NA2        u330(.A(men_men_n346_), .B(men_men_n345_), .Y(men_men_n347_));
  OAI210     u331(.A0(men_men_n347_), .A1(men_men_n339_), .B0(x6), .Y(men_men_n348_));
  OAI210     u332(.A0(men_men_n151_), .A1(men_men_n45_), .B0(men_men_n126_), .Y(men_men_n349_));
  NA3        u333(.A(men_men_n52_), .B(men_men_n36_), .C(men_men_n30_), .Y(men_men_n350_));
  AOI220     u334(.A0(men_men_n350_), .A1(men_men_n349_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n351_));
  AOI210     u335(.A0(men_men_n119_), .A1(men_men_n413_), .B0(x1), .Y(men_men_n352_));
  INV        u336(.A(men_men_n352_), .Y(men_men_n353_));
  NAi31      u337(.An(x2), .B(x8), .C(x0), .Y(men_men_n354_));
  OAI210     u338(.A0(men_men_n354_), .A1(x4), .B0(men_men_n152_), .Y(men_men_n355_));
  NA3        u339(.A(men_men_n355_), .B(men_men_n137_), .C(x9), .Y(men_men_n356_));
  NO4        u340(.A(x8), .B(men_men_n263_), .C(x9), .D(x2), .Y(men_men_n357_));
  NOi21      u341(.An(men_men_n117_), .B(men_men_n166_), .Y(men_men_n358_));
  NO3        u342(.A(men_men_n358_), .B(men_men_n357_), .C(men_men_n18_), .Y(men_men_n359_));
  NO3        u343(.A(x9), .B(men_men_n143_), .C(x0), .Y(men_men_n360_));
  NA2        u344(.A(men_men_n360_), .B(x8), .Y(men_men_n361_));
  NA4        u345(.A(men_men_n361_), .B(men_men_n359_), .C(men_men_n356_), .D(men_men_n47_), .Y(men_men_n362_));
  OAI210     u346(.A0(men_men_n353_), .A1(men_men_n351_), .B0(men_men_n362_), .Y(men_men_n363_));
  AOI210     u347(.A0(men_men_n36_), .A1(x9), .B0(x0), .Y(men_men_n364_));
  NO3        u348(.A(men_men_n364_), .B(men_men_n117_), .C(men_men_n41_), .Y(men_men_n365_));
  NOi31      u349(.An(x1), .B(x8), .C(x7), .Y(men_men_n366_));
  AOI220     u350(.A0(men_men_n366_), .A1(men_men_n308_), .B0(men_men_n118_), .B1(x3), .Y(men_men_n367_));
  AOI210     u351(.A0(men_men_n231_), .A1(men_men_n57_), .B0(men_men_n116_), .Y(men_men_n368_));
  OAI210     u352(.A0(men_men_n368_), .A1(x3), .B0(men_men_n367_), .Y(men_men_n369_));
  NO3        u353(.A(men_men_n369_), .B(men_men_n365_), .C(x2), .Y(men_men_n370_));
  OAI220     u354(.A0(men_men_n309_), .A1(men_men_n267_), .B0(men_men_n263_), .B1(men_men_n41_), .Y(men_men_n371_));
  AOI210     u355(.A0(x9), .A1(men_men_n45_), .B0(men_men_n335_), .Y(men_men_n372_));
  AOI220     u356(.A0(men_men_n372_), .A1(men_men_n88_), .B0(men_men_n371_), .B1(men_men_n143_), .Y(men_men_n373_));
  NO2        u357(.A(men_men_n373_), .B(men_men_n51_), .Y(men_men_n374_));
  NO2        u358(.A(men_men_n374_), .B(men_men_n370_), .Y(men_men_n375_));
  AOI210     u359(.A0(men_men_n375_), .A1(men_men_n363_), .B0(men_men_n25_), .Y(men_men_n376_));
  NA4        u360(.A(men_men_n30_), .B(men_men_n88_), .C(x2), .D(men_men_n17_), .Y(men_men_n377_));
  NO3        u361(.A(men_men_n59_), .B(x4), .C(x1), .Y(men_men_n378_));
  NO3        u362(.A(men_men_n64_), .B(men_men_n18_), .C(x0), .Y(men_men_n379_));
  AOI220     u363(.A0(men_men_n379_), .A1(men_men_n232_), .B0(men_men_n378_), .B1(men_men_n343_), .Y(men_men_n380_));
  NO2        u364(.A(men_men_n380_), .B(men_men_n99_), .Y(men_men_n381_));
  NO3        u365(.A(men_men_n236_), .B(men_men_n161_), .C(men_men_n38_), .Y(men_men_n382_));
  OAI210     u366(.A0(men_men_n382_), .A1(men_men_n381_), .B0(x7), .Y(men_men_n383_));
  NA2        u367(.A(men_men_n383_), .B(men_men_n377_), .Y(men_men_n384_));
  OAI210     u368(.A0(men_men_n384_), .A1(men_men_n376_), .B0(men_men_n34_), .Y(men_men_n385_));
  NO2        u369(.A(men_men_n360_), .B(men_men_n185_), .Y(men_men_n386_));
  NO4        u370(.A(men_men_n386_), .B(men_men_n72_), .C(x4), .D(men_men_n51_), .Y(men_men_n387_));
  NA2        u371(.A(men_men_n222_), .B(men_men_n21_), .Y(men_men_n388_));
  NO2        u372(.A(men_men_n150_), .B(men_men_n126_), .Y(men_men_n389_));
  NA2        u373(.A(men_men_n389_), .B(men_men_n388_), .Y(men_men_n390_));
  AOI210     u374(.A0(men_men_n390_), .A1(men_men_n153_), .B0(men_men_n27_), .Y(men_men_n391_));
  AOI220     u375(.A0(x3), .A1(men_men_n88_), .B0(men_men_n140_), .B1(men_men_n179_), .Y(men_men_n392_));
  NA3        u376(.A(men_men_n392_), .B(men_men_n354_), .C(men_men_n86_), .Y(men_men_n393_));
  NA2        u377(.A(men_men_n393_), .B(men_men_n162_), .Y(men_men_n394_));
  OAI220     u378(.A0(men_men_n411_), .A1(x2), .B0(men_men_n150_), .B1(men_men_n41_), .Y(men_men_n395_));
  AOI210     u379(.A0(men_men_n152_), .A1(men_men_n26_), .B0(men_men_n68_), .Y(men_men_n396_));
  OAI210     u380(.A0(men_men_n139_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n397_));
  NO3        u381(.A(men_men_n366_), .B(x3), .C(men_men_n51_), .Y(men_men_n398_));
  AOI210     u382(.A0(men_men_n398_), .A1(men_men_n397_), .B0(men_men_n396_), .Y(men_men_n399_));
  INV        u383(.A(men_men_n399_), .Y(men_men_n400_));
  AOI220     u384(.A0(men_men_n400_), .A1(x0), .B0(men_men_n395_), .B1(men_men_n126_), .Y(men_men_n401_));
  AOI210     u385(.A0(men_men_n401_), .A1(men_men_n394_), .B0(men_men_n207_), .Y(men_men_n402_));
  NA2        u386(.A(x9), .B(x5), .Y(men_men_n403_));
  NO4        u387(.A(men_men_n102_), .B(men_men_n403_), .C(men_men_n57_), .D(men_men_n31_), .Y(men_men_n404_));
  NO4        u388(.A(men_men_n404_), .B(men_men_n402_), .C(men_men_n391_), .D(men_men_n387_), .Y(men_men_n405_));
  NA3        u389(.A(men_men_n405_), .B(men_men_n385_), .C(men_men_n348_), .Y(men_men_n406_));
  AOI210     u390(.A0(men_men_n333_), .A1(men_men_n25_), .B0(men_men_n406_), .Y(men05));
  INV        u391(.A(men_men_n166_), .Y(men_men_n410_));
  INV        u392(.A(x9), .Y(men_men_n411_));
  INV        u393(.A(x0), .Y(men_men_n412_));
  INV        u394(.A(x4), .Y(men_men_n413_));
  INV        u395(.A(x0), .Y(men_men_n414_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule